module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module pg_fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] pg_fa_xor0, output [0:0] pg_fa_and0, output [0:0] pg_fa_xor1);
  xor_gate xor_gate_pg_fa_xor0(.a(a[0]), .b(b[0]), .out(pg_fa_xor0));
  and_gate and_gate_pg_fa_and0(.a(a[0]), .b(b[0]), .out(pg_fa_and0));
  xor_gate xor_gate_pg_fa_xor1(.a(pg_fa_xor0[0]), .b(cin[0]), .out(pg_fa_xor1));
endmodule

module u_pg_rca16(input [15:0] a, input [15:0] b, output [16:0] u_pg_rca16_out);
  wire [0:0] u_pg_rca16_pg_fa0_xor0;
  wire [0:0] u_pg_rca16_pg_fa0_and0;
  wire [0:0] u_pg_rca16_pg_fa1_xor0;
  wire [0:0] u_pg_rca16_pg_fa1_and0;
  wire [0:0] u_pg_rca16_pg_fa1_xor1;
  wire [0:0] u_pg_rca16_and1;
  wire [0:0] u_pg_rca16_or1;
  wire [0:0] u_pg_rca16_pg_fa2_xor0;
  wire [0:0] u_pg_rca16_pg_fa2_and0;
  wire [0:0] u_pg_rca16_pg_fa2_xor1;
  wire [0:0] u_pg_rca16_and2;
  wire [0:0] u_pg_rca16_or2;
  wire [0:0] u_pg_rca16_pg_fa3_xor0;
  wire [0:0] u_pg_rca16_pg_fa3_and0;
  wire [0:0] u_pg_rca16_pg_fa3_xor1;
  wire [0:0] u_pg_rca16_and3;
  wire [0:0] u_pg_rca16_or3;
  wire [0:0] u_pg_rca16_pg_fa4_xor0;
  wire [0:0] u_pg_rca16_pg_fa4_and0;
  wire [0:0] u_pg_rca16_pg_fa4_xor1;
  wire [0:0] u_pg_rca16_and4;
  wire [0:0] u_pg_rca16_or4;
  wire [0:0] u_pg_rca16_pg_fa5_xor0;
  wire [0:0] u_pg_rca16_pg_fa5_and0;
  wire [0:0] u_pg_rca16_pg_fa5_xor1;
  wire [0:0] u_pg_rca16_and5;
  wire [0:0] u_pg_rca16_or5;
  wire [0:0] u_pg_rca16_pg_fa6_xor0;
  wire [0:0] u_pg_rca16_pg_fa6_and0;
  wire [0:0] u_pg_rca16_pg_fa6_xor1;
  wire [0:0] u_pg_rca16_and6;
  wire [0:0] u_pg_rca16_or6;
  wire [0:0] u_pg_rca16_pg_fa7_xor0;
  wire [0:0] u_pg_rca16_pg_fa7_and0;
  wire [0:0] u_pg_rca16_pg_fa7_xor1;
  wire [0:0] u_pg_rca16_and7;
  wire [0:0] u_pg_rca16_or7;
  wire [0:0] u_pg_rca16_pg_fa8_xor0;
  wire [0:0] u_pg_rca16_pg_fa8_and0;
  wire [0:0] u_pg_rca16_pg_fa8_xor1;
  wire [0:0] u_pg_rca16_and8;
  wire [0:0] u_pg_rca16_or8;
  wire [0:0] u_pg_rca16_pg_fa9_xor0;
  wire [0:0] u_pg_rca16_pg_fa9_and0;
  wire [0:0] u_pg_rca16_pg_fa9_xor1;
  wire [0:0] u_pg_rca16_and9;
  wire [0:0] u_pg_rca16_or9;
  wire [0:0] u_pg_rca16_pg_fa10_xor0;
  wire [0:0] u_pg_rca16_pg_fa10_and0;
  wire [0:0] u_pg_rca16_pg_fa10_xor1;
  wire [0:0] u_pg_rca16_and10;
  wire [0:0] u_pg_rca16_or10;
  wire [0:0] u_pg_rca16_pg_fa11_xor0;
  wire [0:0] u_pg_rca16_pg_fa11_and0;
  wire [0:0] u_pg_rca16_pg_fa11_xor1;
  wire [0:0] u_pg_rca16_and11;
  wire [0:0] u_pg_rca16_or11;
  wire [0:0] u_pg_rca16_pg_fa12_xor0;
  wire [0:0] u_pg_rca16_pg_fa12_and0;
  wire [0:0] u_pg_rca16_pg_fa12_xor1;
  wire [0:0] u_pg_rca16_and12;
  wire [0:0] u_pg_rca16_or12;
  wire [0:0] u_pg_rca16_pg_fa13_xor0;
  wire [0:0] u_pg_rca16_pg_fa13_and0;
  wire [0:0] u_pg_rca16_pg_fa13_xor1;
  wire [0:0] u_pg_rca16_and13;
  wire [0:0] u_pg_rca16_or13;
  wire [0:0] u_pg_rca16_pg_fa14_xor0;
  wire [0:0] u_pg_rca16_pg_fa14_and0;
  wire [0:0] u_pg_rca16_pg_fa14_xor1;
  wire [0:0] u_pg_rca16_and14;
  wire [0:0] u_pg_rca16_or14;
  wire [0:0] u_pg_rca16_pg_fa15_xor0;
  wire [0:0] u_pg_rca16_pg_fa15_and0;
  wire [0:0] u_pg_rca16_pg_fa15_xor1;
  wire [0:0] u_pg_rca16_and15;
  wire [0:0] u_pg_rca16_or15;

  pg_fa pg_fa_u_pg_rca16_pg_fa0_out(.a(a[0]), .b(b[0]), .cin(1'b0), .pg_fa_xor0(u_pg_rca16_pg_fa0_xor0), .pg_fa_and0(u_pg_rca16_pg_fa0_and0), .pg_fa_xor1());
  pg_fa pg_fa_u_pg_rca16_pg_fa1_out(.a(a[1]), .b(b[1]), .cin(u_pg_rca16_pg_fa0_and0[0]), .pg_fa_xor0(u_pg_rca16_pg_fa1_xor0), .pg_fa_and0(u_pg_rca16_pg_fa1_and0), .pg_fa_xor1(u_pg_rca16_pg_fa1_xor1));
  and_gate and_gate_u_pg_rca16_and1(.a(u_pg_rca16_pg_fa0_and0[0]), .b(u_pg_rca16_pg_fa1_xor0[0]), .out(u_pg_rca16_and1));
  or_gate or_gate_u_pg_rca16_or1(.a(u_pg_rca16_and1[0]), .b(u_pg_rca16_pg_fa1_and0[0]), .out(u_pg_rca16_or1));
  pg_fa pg_fa_u_pg_rca16_pg_fa2_out(.a(a[2]), .b(b[2]), .cin(u_pg_rca16_or1[0]), .pg_fa_xor0(u_pg_rca16_pg_fa2_xor0), .pg_fa_and0(u_pg_rca16_pg_fa2_and0), .pg_fa_xor1(u_pg_rca16_pg_fa2_xor1));
  and_gate and_gate_u_pg_rca16_and2(.a(u_pg_rca16_or1[0]), .b(u_pg_rca16_pg_fa2_xor0[0]), .out(u_pg_rca16_and2));
  or_gate or_gate_u_pg_rca16_or2(.a(u_pg_rca16_and2[0]), .b(u_pg_rca16_pg_fa2_and0[0]), .out(u_pg_rca16_or2));
  pg_fa pg_fa_u_pg_rca16_pg_fa3_out(.a(a[3]), .b(b[3]), .cin(u_pg_rca16_or2[0]), .pg_fa_xor0(u_pg_rca16_pg_fa3_xor0), .pg_fa_and0(u_pg_rca16_pg_fa3_and0), .pg_fa_xor1(u_pg_rca16_pg_fa3_xor1));
  and_gate and_gate_u_pg_rca16_and3(.a(u_pg_rca16_or2[0]), .b(u_pg_rca16_pg_fa3_xor0[0]), .out(u_pg_rca16_and3));
  or_gate or_gate_u_pg_rca16_or3(.a(u_pg_rca16_and3[0]), .b(u_pg_rca16_pg_fa3_and0[0]), .out(u_pg_rca16_or3));
  pg_fa pg_fa_u_pg_rca16_pg_fa4_out(.a(a[4]), .b(b[4]), .cin(u_pg_rca16_or3[0]), .pg_fa_xor0(u_pg_rca16_pg_fa4_xor0), .pg_fa_and0(u_pg_rca16_pg_fa4_and0), .pg_fa_xor1(u_pg_rca16_pg_fa4_xor1));
  and_gate and_gate_u_pg_rca16_and4(.a(u_pg_rca16_or3[0]), .b(u_pg_rca16_pg_fa4_xor0[0]), .out(u_pg_rca16_and4));
  or_gate or_gate_u_pg_rca16_or4(.a(u_pg_rca16_and4[0]), .b(u_pg_rca16_pg_fa4_and0[0]), .out(u_pg_rca16_or4));
  pg_fa pg_fa_u_pg_rca16_pg_fa5_out(.a(a[5]), .b(b[5]), .cin(u_pg_rca16_or4[0]), .pg_fa_xor0(u_pg_rca16_pg_fa5_xor0), .pg_fa_and0(u_pg_rca16_pg_fa5_and0), .pg_fa_xor1(u_pg_rca16_pg_fa5_xor1));
  and_gate and_gate_u_pg_rca16_and5(.a(u_pg_rca16_or4[0]), .b(u_pg_rca16_pg_fa5_xor0[0]), .out(u_pg_rca16_and5));
  or_gate or_gate_u_pg_rca16_or5(.a(u_pg_rca16_and5[0]), .b(u_pg_rca16_pg_fa5_and0[0]), .out(u_pg_rca16_or5));
  pg_fa pg_fa_u_pg_rca16_pg_fa6_out(.a(a[6]), .b(b[6]), .cin(u_pg_rca16_or5[0]), .pg_fa_xor0(u_pg_rca16_pg_fa6_xor0), .pg_fa_and0(u_pg_rca16_pg_fa6_and0), .pg_fa_xor1(u_pg_rca16_pg_fa6_xor1));
  and_gate and_gate_u_pg_rca16_and6(.a(u_pg_rca16_or5[0]), .b(u_pg_rca16_pg_fa6_xor0[0]), .out(u_pg_rca16_and6));
  or_gate or_gate_u_pg_rca16_or6(.a(u_pg_rca16_and6[0]), .b(u_pg_rca16_pg_fa6_and0[0]), .out(u_pg_rca16_or6));
  pg_fa pg_fa_u_pg_rca16_pg_fa7_out(.a(a[7]), .b(b[7]), .cin(u_pg_rca16_or6[0]), .pg_fa_xor0(u_pg_rca16_pg_fa7_xor0), .pg_fa_and0(u_pg_rca16_pg_fa7_and0), .pg_fa_xor1(u_pg_rca16_pg_fa7_xor1));
  and_gate and_gate_u_pg_rca16_and7(.a(u_pg_rca16_or6[0]), .b(u_pg_rca16_pg_fa7_xor0[0]), .out(u_pg_rca16_and7));
  or_gate or_gate_u_pg_rca16_or7(.a(u_pg_rca16_and7[0]), .b(u_pg_rca16_pg_fa7_and0[0]), .out(u_pg_rca16_or7));
  pg_fa pg_fa_u_pg_rca16_pg_fa8_out(.a(a[8]), .b(b[8]), .cin(u_pg_rca16_or7[0]), .pg_fa_xor0(u_pg_rca16_pg_fa8_xor0), .pg_fa_and0(u_pg_rca16_pg_fa8_and0), .pg_fa_xor1(u_pg_rca16_pg_fa8_xor1));
  and_gate and_gate_u_pg_rca16_and8(.a(u_pg_rca16_or7[0]), .b(u_pg_rca16_pg_fa8_xor0[0]), .out(u_pg_rca16_and8));
  or_gate or_gate_u_pg_rca16_or8(.a(u_pg_rca16_and8[0]), .b(u_pg_rca16_pg_fa8_and0[0]), .out(u_pg_rca16_or8));
  pg_fa pg_fa_u_pg_rca16_pg_fa9_out(.a(a[9]), .b(b[9]), .cin(u_pg_rca16_or8[0]), .pg_fa_xor0(u_pg_rca16_pg_fa9_xor0), .pg_fa_and0(u_pg_rca16_pg_fa9_and0), .pg_fa_xor1(u_pg_rca16_pg_fa9_xor1));
  and_gate and_gate_u_pg_rca16_and9(.a(u_pg_rca16_or8[0]), .b(u_pg_rca16_pg_fa9_xor0[0]), .out(u_pg_rca16_and9));
  or_gate or_gate_u_pg_rca16_or9(.a(u_pg_rca16_and9[0]), .b(u_pg_rca16_pg_fa9_and0[0]), .out(u_pg_rca16_or9));
  pg_fa pg_fa_u_pg_rca16_pg_fa10_out(.a(a[10]), .b(b[10]), .cin(u_pg_rca16_or9[0]), .pg_fa_xor0(u_pg_rca16_pg_fa10_xor0), .pg_fa_and0(u_pg_rca16_pg_fa10_and0), .pg_fa_xor1(u_pg_rca16_pg_fa10_xor1));
  and_gate and_gate_u_pg_rca16_and10(.a(u_pg_rca16_or9[0]), .b(u_pg_rca16_pg_fa10_xor0[0]), .out(u_pg_rca16_and10));
  or_gate or_gate_u_pg_rca16_or10(.a(u_pg_rca16_and10[0]), .b(u_pg_rca16_pg_fa10_and0[0]), .out(u_pg_rca16_or10));
  pg_fa pg_fa_u_pg_rca16_pg_fa11_out(.a(a[11]), .b(b[11]), .cin(u_pg_rca16_or10[0]), .pg_fa_xor0(u_pg_rca16_pg_fa11_xor0), .pg_fa_and0(u_pg_rca16_pg_fa11_and0), .pg_fa_xor1(u_pg_rca16_pg_fa11_xor1));
  and_gate and_gate_u_pg_rca16_and11(.a(u_pg_rca16_or10[0]), .b(u_pg_rca16_pg_fa11_xor0[0]), .out(u_pg_rca16_and11));
  or_gate or_gate_u_pg_rca16_or11(.a(u_pg_rca16_and11[0]), .b(u_pg_rca16_pg_fa11_and0[0]), .out(u_pg_rca16_or11));
  pg_fa pg_fa_u_pg_rca16_pg_fa12_out(.a(a[12]), .b(b[12]), .cin(u_pg_rca16_or11[0]), .pg_fa_xor0(u_pg_rca16_pg_fa12_xor0), .pg_fa_and0(u_pg_rca16_pg_fa12_and0), .pg_fa_xor1(u_pg_rca16_pg_fa12_xor1));
  and_gate and_gate_u_pg_rca16_and12(.a(u_pg_rca16_or11[0]), .b(u_pg_rca16_pg_fa12_xor0[0]), .out(u_pg_rca16_and12));
  or_gate or_gate_u_pg_rca16_or12(.a(u_pg_rca16_and12[0]), .b(u_pg_rca16_pg_fa12_and0[0]), .out(u_pg_rca16_or12));
  pg_fa pg_fa_u_pg_rca16_pg_fa13_out(.a(a[13]), .b(b[13]), .cin(u_pg_rca16_or12[0]), .pg_fa_xor0(u_pg_rca16_pg_fa13_xor0), .pg_fa_and0(u_pg_rca16_pg_fa13_and0), .pg_fa_xor1(u_pg_rca16_pg_fa13_xor1));
  and_gate and_gate_u_pg_rca16_and13(.a(u_pg_rca16_or12[0]), .b(u_pg_rca16_pg_fa13_xor0[0]), .out(u_pg_rca16_and13));
  or_gate or_gate_u_pg_rca16_or13(.a(u_pg_rca16_and13[0]), .b(u_pg_rca16_pg_fa13_and0[0]), .out(u_pg_rca16_or13));
  pg_fa pg_fa_u_pg_rca16_pg_fa14_out(.a(a[14]), .b(b[14]), .cin(u_pg_rca16_or13[0]), .pg_fa_xor0(u_pg_rca16_pg_fa14_xor0), .pg_fa_and0(u_pg_rca16_pg_fa14_and0), .pg_fa_xor1(u_pg_rca16_pg_fa14_xor1));
  and_gate and_gate_u_pg_rca16_and14(.a(u_pg_rca16_or13[0]), .b(u_pg_rca16_pg_fa14_xor0[0]), .out(u_pg_rca16_and14));
  or_gate or_gate_u_pg_rca16_or14(.a(u_pg_rca16_and14[0]), .b(u_pg_rca16_pg_fa14_and0[0]), .out(u_pg_rca16_or14));
  pg_fa pg_fa_u_pg_rca16_pg_fa15_out(.a(a[15]), .b(b[15]), .cin(u_pg_rca16_or14[0]), .pg_fa_xor0(u_pg_rca16_pg_fa15_xor0), .pg_fa_and0(u_pg_rca16_pg_fa15_and0), .pg_fa_xor1(u_pg_rca16_pg_fa15_xor1));
  and_gate and_gate_u_pg_rca16_and15(.a(u_pg_rca16_or14[0]), .b(u_pg_rca16_pg_fa15_xor0[0]), .out(u_pg_rca16_and15));
  or_gate or_gate_u_pg_rca16_or15(.a(u_pg_rca16_and15[0]), .b(u_pg_rca16_pg_fa15_and0[0]), .out(u_pg_rca16_or15));

  assign u_pg_rca16_out[0] = u_pg_rca16_pg_fa0_xor0[0];
  assign u_pg_rca16_out[1] = u_pg_rca16_pg_fa1_xor1[0];
  assign u_pg_rca16_out[2] = u_pg_rca16_pg_fa2_xor1[0];
  assign u_pg_rca16_out[3] = u_pg_rca16_pg_fa3_xor1[0];
  assign u_pg_rca16_out[4] = u_pg_rca16_pg_fa4_xor1[0];
  assign u_pg_rca16_out[5] = u_pg_rca16_pg_fa5_xor1[0];
  assign u_pg_rca16_out[6] = u_pg_rca16_pg_fa6_xor1[0];
  assign u_pg_rca16_out[7] = u_pg_rca16_pg_fa7_xor1[0];
  assign u_pg_rca16_out[8] = u_pg_rca16_pg_fa8_xor1[0];
  assign u_pg_rca16_out[9] = u_pg_rca16_pg_fa9_xor1[0];
  assign u_pg_rca16_out[10] = u_pg_rca16_pg_fa10_xor1[0];
  assign u_pg_rca16_out[11] = u_pg_rca16_pg_fa11_xor1[0];
  assign u_pg_rca16_out[12] = u_pg_rca16_pg_fa12_xor1[0];
  assign u_pg_rca16_out[13] = u_pg_rca16_pg_fa13_xor1[0];
  assign u_pg_rca16_out[14] = u_pg_rca16_pg_fa14_xor1[0];
  assign u_pg_rca16_out[15] = u_pg_rca16_pg_fa15_xor1[0];
  assign u_pg_rca16_out[16] = u_pg_rca16_or15[0];
endmodule