module s_cla16(input [15:0] a, input [15:0] b, output [16:0] s_cla16_out);
  wire s_cla16_pg_logic0_or0;
  wire s_cla16_pg_logic0_and0;
  wire s_cla16_pg_logic0_xor0;
  wire s_cla16_pg_logic1_or0;
  wire s_cla16_pg_logic1_and0;
  wire s_cla16_pg_logic1_xor0;
  wire s_cla16_xor1;
  wire s_cla16_and0;
  wire s_cla16_or0;
  wire s_cla16_pg_logic2_or0;
  wire s_cla16_pg_logic2_and0;
  wire s_cla16_pg_logic2_xor0;
  wire s_cla16_xor2;
  wire s_cla16_and1;
  wire s_cla16_and2;
  wire s_cla16_and3;
  wire s_cla16_and4;
  wire s_cla16_or1;
  wire s_cla16_or2;
  wire s_cla16_pg_logic3_or0;
  wire s_cla16_pg_logic3_and0;
  wire s_cla16_pg_logic3_xor0;
  wire s_cla16_xor3;
  wire s_cla16_and5;
  wire s_cla16_and6;
  wire s_cla16_and7;
  wire s_cla16_and8;
  wire s_cla16_and9;
  wire s_cla16_and10;
  wire s_cla16_and11;
  wire s_cla16_or3;
  wire s_cla16_or4;
  wire s_cla16_or5;
  wire s_cla16_pg_logic4_or0;
  wire s_cla16_pg_logic4_and0;
  wire s_cla16_pg_logic4_xor0;
  wire s_cla16_xor4;
  wire s_cla16_and12;
  wire s_cla16_or6;
  wire s_cla16_pg_logic5_or0;
  wire s_cla16_pg_logic5_and0;
  wire s_cla16_pg_logic5_xor0;
  wire s_cla16_xor5;
  wire s_cla16_and13;
  wire s_cla16_and14;
  wire s_cla16_and15;
  wire s_cla16_or7;
  wire s_cla16_or8;
  wire s_cla16_pg_logic6_or0;
  wire s_cla16_pg_logic6_and0;
  wire s_cla16_pg_logic6_xor0;
  wire s_cla16_xor6;
  wire s_cla16_and16;
  wire s_cla16_and17;
  wire s_cla16_and18;
  wire s_cla16_and19;
  wire s_cla16_and20;
  wire s_cla16_and21;
  wire s_cla16_or9;
  wire s_cla16_or10;
  wire s_cla16_or11;
  wire s_cla16_pg_logic7_or0;
  wire s_cla16_pg_logic7_and0;
  wire s_cla16_pg_logic7_xor0;
  wire s_cla16_xor7;
  wire s_cla16_and22;
  wire s_cla16_and23;
  wire s_cla16_and24;
  wire s_cla16_and25;
  wire s_cla16_and26;
  wire s_cla16_and27;
  wire s_cla16_and28;
  wire s_cla16_and29;
  wire s_cla16_and30;
  wire s_cla16_and31;
  wire s_cla16_or12;
  wire s_cla16_or13;
  wire s_cla16_or14;
  wire s_cla16_or15;
  wire s_cla16_pg_logic8_or0;
  wire s_cla16_pg_logic8_and0;
  wire s_cla16_pg_logic8_xor0;
  wire s_cla16_xor8;
  wire s_cla16_and32;
  wire s_cla16_or16;
  wire s_cla16_pg_logic9_or0;
  wire s_cla16_pg_logic9_and0;
  wire s_cla16_pg_logic9_xor0;
  wire s_cla16_xor9;
  wire s_cla16_and33;
  wire s_cla16_and34;
  wire s_cla16_and35;
  wire s_cla16_or17;
  wire s_cla16_or18;
  wire s_cla16_pg_logic10_or0;
  wire s_cla16_pg_logic10_and0;
  wire s_cla16_pg_logic10_xor0;
  wire s_cla16_xor10;
  wire s_cla16_and36;
  wire s_cla16_and37;
  wire s_cla16_and38;
  wire s_cla16_and39;
  wire s_cla16_and40;
  wire s_cla16_and41;
  wire s_cla16_or19;
  wire s_cla16_or20;
  wire s_cla16_or21;
  wire s_cla16_pg_logic11_or0;
  wire s_cla16_pg_logic11_and0;
  wire s_cla16_pg_logic11_xor0;
  wire s_cla16_xor11;
  wire s_cla16_and42;
  wire s_cla16_and43;
  wire s_cla16_and44;
  wire s_cla16_and45;
  wire s_cla16_and46;
  wire s_cla16_and47;
  wire s_cla16_and48;
  wire s_cla16_and49;
  wire s_cla16_and50;
  wire s_cla16_and51;
  wire s_cla16_or22;
  wire s_cla16_or23;
  wire s_cla16_or24;
  wire s_cla16_or25;
  wire s_cla16_pg_logic12_or0;
  wire s_cla16_pg_logic12_and0;
  wire s_cla16_pg_logic12_xor0;
  wire s_cla16_xor12;
  wire s_cla16_and52;
  wire s_cla16_or26;
  wire s_cla16_pg_logic13_or0;
  wire s_cla16_pg_logic13_and0;
  wire s_cla16_pg_logic13_xor0;
  wire s_cla16_xor13;
  wire s_cla16_and53;
  wire s_cla16_and54;
  wire s_cla16_and55;
  wire s_cla16_or27;
  wire s_cla16_or28;
  wire s_cla16_pg_logic14_or0;
  wire s_cla16_pg_logic14_and0;
  wire s_cla16_pg_logic14_xor0;
  wire s_cla16_xor14;
  wire s_cla16_and56;
  wire s_cla16_and57;
  wire s_cla16_and58;
  wire s_cla16_and59;
  wire s_cla16_and60;
  wire s_cla16_and61;
  wire s_cla16_or29;
  wire s_cla16_or30;
  wire s_cla16_or31;
  wire s_cla16_pg_logic15_or0;
  wire s_cla16_pg_logic15_and0;
  wire s_cla16_pg_logic15_xor0;
  wire s_cla16_xor15;
  wire s_cla16_and62;
  wire s_cla16_and63;
  wire s_cla16_and64;
  wire s_cla16_and65;
  wire s_cla16_and66;
  wire s_cla16_and67;
  wire s_cla16_and68;
  wire s_cla16_and69;
  wire s_cla16_and70;
  wire s_cla16_and71;
  wire s_cla16_or32;
  wire s_cla16_or33;
  wire s_cla16_or34;
  wire s_cla16_or35;
  wire s_cla16_xor16;
  wire s_cla16_xor17;

  assign s_cla16_pg_logic0_or0 = a[0] | b[0];
  assign s_cla16_pg_logic0_and0 = a[0] & b[0];
  assign s_cla16_pg_logic0_xor0 = a[0] ^ b[0];
  assign s_cla16_pg_logic1_or0 = a[1] | b[1];
  assign s_cla16_pg_logic1_and0 = a[1] & b[1];
  assign s_cla16_pg_logic1_xor0 = a[1] ^ b[1];
  assign s_cla16_xor1 = s_cla16_pg_logic1_xor0 ^ s_cla16_pg_logic0_and0;
  assign s_cla16_and0 = s_cla16_pg_logic0_and0 & s_cla16_pg_logic1_or0;
  assign s_cla16_or0 = s_cla16_pg_logic1_and0 | s_cla16_and0;
  assign s_cla16_pg_logic2_or0 = a[2] | b[2];
  assign s_cla16_pg_logic2_and0 = a[2] & b[2];
  assign s_cla16_pg_logic2_xor0 = a[2] ^ b[2];
  assign s_cla16_xor2 = s_cla16_pg_logic2_xor0 ^ s_cla16_or0;
  assign s_cla16_and1 = s_cla16_pg_logic2_or0 & s_cla16_pg_logic0_or0;
  assign s_cla16_and2 = s_cla16_pg_logic0_and0 & s_cla16_pg_logic2_or0;
  assign s_cla16_and3 = s_cla16_and2 & s_cla16_pg_logic1_or0;
  assign s_cla16_and4 = s_cla16_pg_logic1_and0 & s_cla16_pg_logic2_or0;
  assign s_cla16_or1 = s_cla16_and3 | s_cla16_and4;
  assign s_cla16_or2 = s_cla16_pg_logic2_and0 | s_cla16_or1;
  assign s_cla16_pg_logic3_or0 = a[3] | b[3];
  assign s_cla16_pg_logic3_and0 = a[3] & b[3];
  assign s_cla16_pg_logic3_xor0 = a[3] ^ b[3];
  assign s_cla16_xor3 = s_cla16_pg_logic3_xor0 ^ s_cla16_or2;
  assign s_cla16_and5 = s_cla16_pg_logic3_or0 & s_cla16_pg_logic1_or0;
  assign s_cla16_and6 = s_cla16_pg_logic0_and0 & s_cla16_pg_logic2_or0;
  assign s_cla16_and7 = s_cla16_pg_logic3_or0 & s_cla16_pg_logic1_or0;
  assign s_cla16_and8 = s_cla16_and6 & s_cla16_and7;
  assign s_cla16_and9 = s_cla16_pg_logic1_and0 & s_cla16_pg_logic3_or0;
  assign s_cla16_and10 = s_cla16_and9 & s_cla16_pg_logic2_or0;
  assign s_cla16_and11 = s_cla16_pg_logic2_and0 & s_cla16_pg_logic3_or0;
  assign s_cla16_or3 = s_cla16_and8 | s_cla16_and11;
  assign s_cla16_or4 = s_cla16_and10 | s_cla16_or3;
  assign s_cla16_or5 = s_cla16_pg_logic3_and0 | s_cla16_or4;
  assign s_cla16_pg_logic4_or0 = a[4] | b[4];
  assign s_cla16_pg_logic4_and0 = a[4] & b[4];
  assign s_cla16_pg_logic4_xor0 = a[4] ^ b[4];
  assign s_cla16_xor4 = s_cla16_pg_logic4_xor0 ^ s_cla16_or5;
  assign s_cla16_and12 = s_cla16_or5 & s_cla16_pg_logic4_or0;
  assign s_cla16_or6 = s_cla16_pg_logic4_and0 | s_cla16_and12;
  assign s_cla16_pg_logic5_or0 = a[5] | b[5];
  assign s_cla16_pg_logic5_and0 = a[5] & b[5];
  assign s_cla16_pg_logic5_xor0 = a[5] ^ b[5];
  assign s_cla16_xor5 = s_cla16_pg_logic5_xor0 ^ s_cla16_or6;
  assign s_cla16_and13 = s_cla16_or5 & s_cla16_pg_logic5_or0;
  assign s_cla16_and14 = s_cla16_and13 & s_cla16_pg_logic4_or0;
  assign s_cla16_and15 = s_cla16_pg_logic4_and0 & s_cla16_pg_logic5_or0;
  assign s_cla16_or7 = s_cla16_and14 | s_cla16_and15;
  assign s_cla16_or8 = s_cla16_pg_logic5_and0 | s_cla16_or7;
  assign s_cla16_pg_logic6_or0 = a[6] | b[6];
  assign s_cla16_pg_logic6_and0 = a[6] & b[6];
  assign s_cla16_pg_logic6_xor0 = a[6] ^ b[6];
  assign s_cla16_xor6 = s_cla16_pg_logic6_xor0 ^ s_cla16_or8;
  assign s_cla16_and16 = s_cla16_or5 & s_cla16_pg_logic5_or0;
  assign s_cla16_and17 = s_cla16_pg_logic6_or0 & s_cla16_pg_logic4_or0;
  assign s_cla16_and18 = s_cla16_and16 & s_cla16_and17;
  assign s_cla16_and19 = s_cla16_pg_logic4_and0 & s_cla16_pg_logic6_or0;
  assign s_cla16_and20 = s_cla16_and19 & s_cla16_pg_logic5_or0;
  assign s_cla16_and21 = s_cla16_pg_logic5_and0 & s_cla16_pg_logic6_or0;
  assign s_cla16_or9 = s_cla16_and18 | s_cla16_and20;
  assign s_cla16_or10 = s_cla16_or9 | s_cla16_and21;
  assign s_cla16_or11 = s_cla16_pg_logic6_and0 | s_cla16_or10;
  assign s_cla16_pg_logic7_or0 = a[7] | b[7];
  assign s_cla16_pg_logic7_and0 = a[7] & b[7];
  assign s_cla16_pg_logic7_xor0 = a[7] ^ b[7];
  assign s_cla16_xor7 = s_cla16_pg_logic7_xor0 ^ s_cla16_or11;
  assign s_cla16_and22 = s_cla16_or5 & s_cla16_pg_logic6_or0;
  assign s_cla16_and23 = s_cla16_pg_logic7_or0 & s_cla16_pg_logic5_or0;
  assign s_cla16_and24 = s_cla16_and22 & s_cla16_and23;
  assign s_cla16_and25 = s_cla16_and24 & s_cla16_pg_logic4_or0;
  assign s_cla16_and26 = s_cla16_pg_logic4_and0 & s_cla16_pg_logic6_or0;
  assign s_cla16_and27 = s_cla16_pg_logic7_or0 & s_cla16_pg_logic5_or0;
  assign s_cla16_and28 = s_cla16_and26 & s_cla16_and27;
  assign s_cla16_and29 = s_cla16_pg_logic5_and0 & s_cla16_pg_logic7_or0;
  assign s_cla16_and30 = s_cla16_and29 & s_cla16_pg_logic6_or0;
  assign s_cla16_and31 = s_cla16_pg_logic6_and0 & s_cla16_pg_logic7_or0;
  assign s_cla16_or12 = s_cla16_and25 | s_cla16_and30;
  assign s_cla16_or13 = s_cla16_and28 | s_cla16_and31;
  assign s_cla16_or14 = s_cla16_or12 | s_cla16_or13;
  assign s_cla16_or15 = s_cla16_pg_logic7_and0 | s_cla16_or14;
  assign s_cla16_pg_logic8_or0 = a[8] | b[8];
  assign s_cla16_pg_logic8_and0 = a[8] & b[8];
  assign s_cla16_pg_logic8_xor0 = a[8] ^ b[8];
  assign s_cla16_xor8 = s_cla16_pg_logic8_xor0 ^ s_cla16_or15;
  assign s_cla16_and32 = s_cla16_or15 & s_cla16_pg_logic8_or0;
  assign s_cla16_or16 = s_cla16_pg_logic8_and0 | s_cla16_and32;
  assign s_cla16_pg_logic9_or0 = a[9] | b[9];
  assign s_cla16_pg_logic9_and0 = a[9] & b[9];
  assign s_cla16_pg_logic9_xor0 = a[9] ^ b[9];
  assign s_cla16_xor9 = s_cla16_pg_logic9_xor0 ^ s_cla16_or16;
  assign s_cla16_and33 = s_cla16_or15 & s_cla16_pg_logic9_or0;
  assign s_cla16_and34 = s_cla16_and33 & s_cla16_pg_logic8_or0;
  assign s_cla16_and35 = s_cla16_pg_logic8_and0 & s_cla16_pg_logic9_or0;
  assign s_cla16_or17 = s_cla16_and34 | s_cla16_and35;
  assign s_cla16_or18 = s_cla16_pg_logic9_and0 | s_cla16_or17;
  assign s_cla16_pg_logic10_or0 = a[10] | b[10];
  assign s_cla16_pg_logic10_and0 = a[10] & b[10];
  assign s_cla16_pg_logic10_xor0 = a[10] ^ b[10];
  assign s_cla16_xor10 = s_cla16_pg_logic10_xor0 ^ s_cla16_or18;
  assign s_cla16_and36 = s_cla16_or15 & s_cla16_pg_logic9_or0;
  assign s_cla16_and37 = s_cla16_pg_logic10_or0 & s_cla16_pg_logic8_or0;
  assign s_cla16_and38 = s_cla16_and36 & s_cla16_and37;
  assign s_cla16_and39 = s_cla16_pg_logic8_and0 & s_cla16_pg_logic10_or0;
  assign s_cla16_and40 = s_cla16_and39 & s_cla16_pg_logic9_or0;
  assign s_cla16_and41 = s_cla16_pg_logic9_and0 & s_cla16_pg_logic10_or0;
  assign s_cla16_or19 = s_cla16_and38 | s_cla16_and40;
  assign s_cla16_or20 = s_cla16_or19 | s_cla16_and41;
  assign s_cla16_or21 = s_cla16_pg_logic10_and0 | s_cla16_or20;
  assign s_cla16_pg_logic11_or0 = a[11] | b[11];
  assign s_cla16_pg_logic11_and0 = a[11] & b[11];
  assign s_cla16_pg_logic11_xor0 = a[11] ^ b[11];
  assign s_cla16_xor11 = s_cla16_pg_logic11_xor0 ^ s_cla16_or21;
  assign s_cla16_and42 = s_cla16_or15 & s_cla16_pg_logic10_or0;
  assign s_cla16_and43 = s_cla16_pg_logic11_or0 & s_cla16_pg_logic9_or0;
  assign s_cla16_and44 = s_cla16_and42 & s_cla16_and43;
  assign s_cla16_and45 = s_cla16_and44 & s_cla16_pg_logic8_or0;
  assign s_cla16_and46 = s_cla16_pg_logic8_and0 & s_cla16_pg_logic10_or0;
  assign s_cla16_and47 = s_cla16_pg_logic11_or0 & s_cla16_pg_logic9_or0;
  assign s_cla16_and48 = s_cla16_and46 & s_cla16_and47;
  assign s_cla16_and49 = s_cla16_pg_logic9_and0 & s_cla16_pg_logic11_or0;
  assign s_cla16_and50 = s_cla16_and49 & s_cla16_pg_logic10_or0;
  assign s_cla16_and51 = s_cla16_pg_logic10_and0 & s_cla16_pg_logic11_or0;
  assign s_cla16_or22 = s_cla16_and45 | s_cla16_and50;
  assign s_cla16_or23 = s_cla16_and48 | s_cla16_and51;
  assign s_cla16_or24 = s_cla16_or22 | s_cla16_or23;
  assign s_cla16_or25 = s_cla16_pg_logic11_and0 | s_cla16_or24;
  assign s_cla16_pg_logic12_or0 = a[12] | b[12];
  assign s_cla16_pg_logic12_and0 = a[12] & b[12];
  assign s_cla16_pg_logic12_xor0 = a[12] ^ b[12];
  assign s_cla16_xor12 = s_cla16_pg_logic12_xor0 ^ s_cla16_or25;
  assign s_cla16_and52 = s_cla16_or25 & s_cla16_pg_logic12_or0;
  assign s_cla16_or26 = s_cla16_pg_logic12_and0 | s_cla16_and52;
  assign s_cla16_pg_logic13_or0 = a[13] | b[13];
  assign s_cla16_pg_logic13_and0 = a[13] & b[13];
  assign s_cla16_pg_logic13_xor0 = a[13] ^ b[13];
  assign s_cla16_xor13 = s_cla16_pg_logic13_xor0 ^ s_cla16_or26;
  assign s_cla16_and53 = s_cla16_or25 & s_cla16_pg_logic13_or0;
  assign s_cla16_and54 = s_cla16_and53 & s_cla16_pg_logic12_or0;
  assign s_cla16_and55 = s_cla16_pg_logic12_and0 & s_cla16_pg_logic13_or0;
  assign s_cla16_or27 = s_cla16_and54 | s_cla16_and55;
  assign s_cla16_or28 = s_cla16_pg_logic13_and0 | s_cla16_or27;
  assign s_cla16_pg_logic14_or0 = a[14] | b[14];
  assign s_cla16_pg_logic14_and0 = a[14] & b[14];
  assign s_cla16_pg_logic14_xor0 = a[14] ^ b[14];
  assign s_cla16_xor14 = s_cla16_pg_logic14_xor0 ^ s_cla16_or28;
  assign s_cla16_and56 = s_cla16_or25 & s_cla16_pg_logic13_or0;
  assign s_cla16_and57 = s_cla16_pg_logic14_or0 & s_cla16_pg_logic12_or0;
  assign s_cla16_and58 = s_cla16_and56 & s_cla16_and57;
  assign s_cla16_and59 = s_cla16_pg_logic12_and0 & s_cla16_pg_logic14_or0;
  assign s_cla16_and60 = s_cla16_and59 & s_cla16_pg_logic13_or0;
  assign s_cla16_and61 = s_cla16_pg_logic13_and0 & s_cla16_pg_logic14_or0;
  assign s_cla16_or29 = s_cla16_and58 | s_cla16_and60;
  assign s_cla16_or30 = s_cla16_or29 | s_cla16_and61;
  assign s_cla16_or31 = s_cla16_pg_logic14_and0 | s_cla16_or30;
  assign s_cla16_pg_logic15_or0 = a[15] | b[15];
  assign s_cla16_pg_logic15_and0 = a[15] & b[15];
  assign s_cla16_pg_logic15_xor0 = a[15] ^ b[15];
  assign s_cla16_xor15 = s_cla16_pg_logic15_xor0 ^ s_cla16_or31;
  assign s_cla16_and62 = s_cla16_or25 & s_cla16_pg_logic14_or0;
  assign s_cla16_and63 = s_cla16_pg_logic15_or0 & s_cla16_pg_logic13_or0;
  assign s_cla16_and64 = s_cla16_and62 & s_cla16_and63;
  assign s_cla16_and65 = s_cla16_and64 & s_cla16_pg_logic12_or0;
  assign s_cla16_and66 = s_cla16_pg_logic12_and0 & s_cla16_pg_logic14_or0;
  assign s_cla16_and67 = s_cla16_pg_logic15_or0 & s_cla16_pg_logic13_or0;
  assign s_cla16_and68 = s_cla16_and66 & s_cla16_and67;
  assign s_cla16_and69 = s_cla16_pg_logic13_and0 & s_cla16_pg_logic15_or0;
  assign s_cla16_and70 = s_cla16_and69 & s_cla16_pg_logic14_or0;
  assign s_cla16_and71 = s_cla16_pg_logic14_and0 & s_cla16_pg_logic15_or0;
  assign s_cla16_or32 = s_cla16_and65 | s_cla16_and70;
  assign s_cla16_or33 = s_cla16_and68 | s_cla16_and71;
  assign s_cla16_or34 = s_cla16_or32 | s_cla16_or33;
  assign s_cla16_or35 = s_cla16_pg_logic15_and0 | s_cla16_or34;
  assign s_cla16_xor16 = a[15] ^ b[15];
  assign s_cla16_xor17 = s_cla16_xor16 ^ s_cla16_or35;

  assign s_cla16_out[0] = s_cla16_pg_logic0_xor0;
  assign s_cla16_out[1] = s_cla16_xor1;
  assign s_cla16_out[2] = s_cla16_xor2;
  assign s_cla16_out[3] = s_cla16_xor3;
  assign s_cla16_out[4] = s_cla16_xor4;
  assign s_cla16_out[5] = s_cla16_xor5;
  assign s_cla16_out[6] = s_cla16_xor6;
  assign s_cla16_out[7] = s_cla16_xor7;
  assign s_cla16_out[8] = s_cla16_xor8;
  assign s_cla16_out[9] = s_cla16_xor9;
  assign s_cla16_out[10] = s_cla16_xor10;
  assign s_cla16_out[11] = s_cla16_xor11;
  assign s_cla16_out[12] = s_cla16_xor12;
  assign s_cla16_out[13] = s_cla16_xor13;
  assign s_cla16_out[14] = s_cla16_xor14;
  assign s_cla16_out[15] = s_cla16_xor15;
  assign s_cla16_out[16] = s_cla16_xor17;
endmodule