module f_u_rca3(input [2:0] a, input [2:0] b, output [3:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire b_0;
  wire b_1;
  wire b_2;
  wire f_u_rca3_ha_a_0;
  wire f_u_rca3_ha_b_0;
  wire f_u_rca3_ha_y0;
  wire f_u_rca3_ha_y1;
  wire f_u_rca3_fa1_a_1;
  wire f_u_rca3_fa1_b_1;
  wire f_u_rca3_fa1_y0;
  wire f_u_rca3_fa1_y1;
  wire f_u_rca3_fa1_f_u_rca3_ha_y1;
  wire f_u_rca3_fa1_y2;
  wire f_u_rca3_fa1_y3;
  wire f_u_rca3_fa1_y4;
  wire f_u_rca3_fa2_a_2;
  wire f_u_rca3_fa2_b_2;
  wire f_u_rca3_fa2_y0;
  wire f_u_rca3_fa2_y1;
  wire f_u_rca3_fa2_f_u_rca3_fa1_y4;
  wire f_u_rca3_fa2_y2;
  wire f_u_rca3_fa2_y3;
  wire f_u_rca3_fa2_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign f_u_rca3_ha_a_0 = a_0;
  assign f_u_rca3_ha_b_0 = b_0;
  assign f_u_rca3_ha_y0 = f_u_rca3_ha_a_0 ^ f_u_rca3_ha_b_0;
  assign f_u_rca3_ha_y1 = f_u_rca3_ha_a_0 & f_u_rca3_ha_b_0;
  assign f_u_rca3_fa1_a_1 = a_1;
  assign f_u_rca3_fa1_b_1 = b_1;
  assign f_u_rca3_fa1_f_u_rca3_ha_y1 = f_u_rca3_ha_y1;
  assign f_u_rca3_fa1_y0 = f_u_rca3_fa1_a_1 ^ f_u_rca3_fa1_b_1;
  assign f_u_rca3_fa1_y1 = f_u_rca3_fa1_a_1 & f_u_rca3_fa1_b_1;
  assign f_u_rca3_fa1_y2 = f_u_rca3_fa1_y0 ^ f_u_rca3_fa1_f_u_rca3_ha_y1;
  assign f_u_rca3_fa1_y3 = f_u_rca3_fa1_y0 & f_u_rca3_fa1_f_u_rca3_ha_y1;
  assign f_u_rca3_fa1_y4 = f_u_rca3_fa1_y1 | f_u_rca3_fa1_y3;
  assign f_u_rca3_fa2_a_2 = a_2;
  assign f_u_rca3_fa2_b_2 = b_2;
  assign f_u_rca3_fa2_f_u_rca3_fa1_y4 = f_u_rca3_fa1_y4;
  assign f_u_rca3_fa2_y0 = f_u_rca3_fa2_a_2 ^ f_u_rca3_fa2_b_2;
  assign f_u_rca3_fa2_y1 = f_u_rca3_fa2_a_2 & f_u_rca3_fa2_b_2;
  assign f_u_rca3_fa2_y2 = f_u_rca3_fa2_y0 ^ f_u_rca3_fa2_f_u_rca3_fa1_y4;
  assign f_u_rca3_fa2_y3 = f_u_rca3_fa2_y0 & f_u_rca3_fa2_f_u_rca3_fa1_y4;
  assign f_u_rca3_fa2_y4 = f_u_rca3_fa2_y1 | f_u_rca3_fa2_y3;

  assign out[0] = f_u_rca3_ha_y0;
  assign out[1] = f_u_rca3_fa1_y2;
  assign out[2] = f_u_rca3_fa2_y2;
  assign out[3] = f_u_rca3_fa2_y4;
endmodule