module f_u_wallace_pg_rca8(input [7:0] a, input [7:0] b, output [15:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire f_u_wallace_pg_rca8_and_2_0_a_2;
  wire f_u_wallace_pg_rca8_and_2_0_b_0;
  wire f_u_wallace_pg_rca8_and_2_0_y0;
  wire f_u_wallace_pg_rca8_and_1_1_a_1;
  wire f_u_wallace_pg_rca8_and_1_1_b_1;
  wire f_u_wallace_pg_rca8_and_1_1_y0;
  wire f_u_wallace_pg_rca8_ha0_f_u_wallace_pg_rca8_and_2_0_y0;
  wire f_u_wallace_pg_rca8_ha0_f_u_wallace_pg_rca8_and_1_1_y0;
  wire f_u_wallace_pg_rca8_ha0_y0;
  wire f_u_wallace_pg_rca8_ha0_y1;
  wire f_u_wallace_pg_rca8_and_3_0_a_3;
  wire f_u_wallace_pg_rca8_and_3_0_b_0;
  wire f_u_wallace_pg_rca8_and_3_0_y0;
  wire f_u_wallace_pg_rca8_and_2_1_a_2;
  wire f_u_wallace_pg_rca8_and_2_1_b_1;
  wire f_u_wallace_pg_rca8_and_2_1_y0;
  wire f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_ha0_y1;
  wire f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_and_3_0_y0;
  wire f_u_wallace_pg_rca8_fa0_y0;
  wire f_u_wallace_pg_rca8_fa0_y1;
  wire f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_and_2_1_y0;
  wire f_u_wallace_pg_rca8_fa0_y2;
  wire f_u_wallace_pg_rca8_fa0_y3;
  wire f_u_wallace_pg_rca8_fa0_y4;
  wire f_u_wallace_pg_rca8_and_4_0_a_4;
  wire f_u_wallace_pg_rca8_and_4_0_b_0;
  wire f_u_wallace_pg_rca8_and_4_0_y0;
  wire f_u_wallace_pg_rca8_and_3_1_a_3;
  wire f_u_wallace_pg_rca8_and_3_1_b_1;
  wire f_u_wallace_pg_rca8_and_3_1_y0;
  wire f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_fa0_y4;
  wire f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_and_4_0_y0;
  wire f_u_wallace_pg_rca8_fa1_y0;
  wire f_u_wallace_pg_rca8_fa1_y1;
  wire f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_and_3_1_y0;
  wire f_u_wallace_pg_rca8_fa1_y2;
  wire f_u_wallace_pg_rca8_fa1_y3;
  wire f_u_wallace_pg_rca8_fa1_y4;
  wire f_u_wallace_pg_rca8_and_5_0_a_5;
  wire f_u_wallace_pg_rca8_and_5_0_b_0;
  wire f_u_wallace_pg_rca8_and_5_0_y0;
  wire f_u_wallace_pg_rca8_and_4_1_a_4;
  wire f_u_wallace_pg_rca8_and_4_1_b_1;
  wire f_u_wallace_pg_rca8_and_4_1_y0;
  wire f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_fa1_y4;
  wire f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_and_5_0_y0;
  wire f_u_wallace_pg_rca8_fa2_y0;
  wire f_u_wallace_pg_rca8_fa2_y1;
  wire f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_and_4_1_y0;
  wire f_u_wallace_pg_rca8_fa2_y2;
  wire f_u_wallace_pg_rca8_fa2_y3;
  wire f_u_wallace_pg_rca8_fa2_y4;
  wire f_u_wallace_pg_rca8_and_6_0_a_6;
  wire f_u_wallace_pg_rca8_and_6_0_b_0;
  wire f_u_wallace_pg_rca8_and_6_0_y0;
  wire f_u_wallace_pg_rca8_and_5_1_a_5;
  wire f_u_wallace_pg_rca8_and_5_1_b_1;
  wire f_u_wallace_pg_rca8_and_5_1_y0;
  wire f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_fa2_y4;
  wire f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_and_6_0_y0;
  wire f_u_wallace_pg_rca8_fa3_y0;
  wire f_u_wallace_pg_rca8_fa3_y1;
  wire f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_and_5_1_y0;
  wire f_u_wallace_pg_rca8_fa3_y2;
  wire f_u_wallace_pg_rca8_fa3_y3;
  wire f_u_wallace_pg_rca8_fa3_y4;
  wire f_u_wallace_pg_rca8_and_7_0_a_7;
  wire f_u_wallace_pg_rca8_and_7_0_b_0;
  wire f_u_wallace_pg_rca8_and_7_0_y0;
  wire f_u_wallace_pg_rca8_and_6_1_a_6;
  wire f_u_wallace_pg_rca8_and_6_1_b_1;
  wire f_u_wallace_pg_rca8_and_6_1_y0;
  wire f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_fa3_y4;
  wire f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_and_7_0_y0;
  wire f_u_wallace_pg_rca8_fa4_y0;
  wire f_u_wallace_pg_rca8_fa4_y1;
  wire f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_and_6_1_y0;
  wire f_u_wallace_pg_rca8_fa4_y2;
  wire f_u_wallace_pg_rca8_fa4_y3;
  wire f_u_wallace_pg_rca8_fa4_y4;
  wire f_u_wallace_pg_rca8_and_7_1_a_7;
  wire f_u_wallace_pg_rca8_and_7_1_b_1;
  wire f_u_wallace_pg_rca8_and_7_1_y0;
  wire f_u_wallace_pg_rca8_and_6_2_a_6;
  wire f_u_wallace_pg_rca8_and_6_2_b_2;
  wire f_u_wallace_pg_rca8_and_6_2_y0;
  wire f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_fa4_y4;
  wire f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_and_7_1_y0;
  wire f_u_wallace_pg_rca8_fa5_y0;
  wire f_u_wallace_pg_rca8_fa5_y1;
  wire f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_and_6_2_y0;
  wire f_u_wallace_pg_rca8_fa5_y2;
  wire f_u_wallace_pg_rca8_fa5_y3;
  wire f_u_wallace_pg_rca8_fa5_y4;
  wire f_u_wallace_pg_rca8_and_7_2_a_7;
  wire f_u_wallace_pg_rca8_and_7_2_b_2;
  wire f_u_wallace_pg_rca8_and_7_2_y0;
  wire f_u_wallace_pg_rca8_and_6_3_a_6;
  wire f_u_wallace_pg_rca8_and_6_3_b_3;
  wire f_u_wallace_pg_rca8_and_6_3_y0;
  wire f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_fa5_y4;
  wire f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_and_7_2_y0;
  wire f_u_wallace_pg_rca8_fa6_y0;
  wire f_u_wallace_pg_rca8_fa6_y1;
  wire f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_and_6_3_y0;
  wire f_u_wallace_pg_rca8_fa6_y2;
  wire f_u_wallace_pg_rca8_fa6_y3;
  wire f_u_wallace_pg_rca8_fa6_y4;
  wire f_u_wallace_pg_rca8_and_7_3_a_7;
  wire f_u_wallace_pg_rca8_and_7_3_b_3;
  wire f_u_wallace_pg_rca8_and_7_3_y0;
  wire f_u_wallace_pg_rca8_and_6_4_a_6;
  wire f_u_wallace_pg_rca8_and_6_4_b_4;
  wire f_u_wallace_pg_rca8_and_6_4_y0;
  wire f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_fa6_y4;
  wire f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_and_7_3_y0;
  wire f_u_wallace_pg_rca8_fa7_y0;
  wire f_u_wallace_pg_rca8_fa7_y1;
  wire f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_and_6_4_y0;
  wire f_u_wallace_pg_rca8_fa7_y2;
  wire f_u_wallace_pg_rca8_fa7_y3;
  wire f_u_wallace_pg_rca8_fa7_y4;
  wire f_u_wallace_pg_rca8_and_7_4_a_7;
  wire f_u_wallace_pg_rca8_and_7_4_b_4;
  wire f_u_wallace_pg_rca8_and_7_4_y0;
  wire f_u_wallace_pg_rca8_and_6_5_a_6;
  wire f_u_wallace_pg_rca8_and_6_5_b_5;
  wire f_u_wallace_pg_rca8_and_6_5_y0;
  wire f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_fa7_y4;
  wire f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_and_7_4_y0;
  wire f_u_wallace_pg_rca8_fa8_y0;
  wire f_u_wallace_pg_rca8_fa8_y1;
  wire f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_and_6_5_y0;
  wire f_u_wallace_pg_rca8_fa8_y2;
  wire f_u_wallace_pg_rca8_fa8_y3;
  wire f_u_wallace_pg_rca8_fa8_y4;
  wire f_u_wallace_pg_rca8_and_7_5_a_7;
  wire f_u_wallace_pg_rca8_and_7_5_b_5;
  wire f_u_wallace_pg_rca8_and_7_5_y0;
  wire f_u_wallace_pg_rca8_and_6_6_a_6;
  wire f_u_wallace_pg_rca8_and_6_6_b_6;
  wire f_u_wallace_pg_rca8_and_6_6_y0;
  wire f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_fa8_y4;
  wire f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_and_7_5_y0;
  wire f_u_wallace_pg_rca8_fa9_y0;
  wire f_u_wallace_pg_rca8_fa9_y1;
  wire f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_and_6_6_y0;
  wire f_u_wallace_pg_rca8_fa9_y2;
  wire f_u_wallace_pg_rca8_fa9_y3;
  wire f_u_wallace_pg_rca8_fa9_y4;
  wire f_u_wallace_pg_rca8_and_1_2_a_1;
  wire f_u_wallace_pg_rca8_and_1_2_b_2;
  wire f_u_wallace_pg_rca8_and_1_2_y0;
  wire f_u_wallace_pg_rca8_and_0_3_a_0;
  wire f_u_wallace_pg_rca8_and_0_3_b_3;
  wire f_u_wallace_pg_rca8_and_0_3_y0;
  wire f_u_wallace_pg_rca8_ha1_f_u_wallace_pg_rca8_and_1_2_y0;
  wire f_u_wallace_pg_rca8_ha1_f_u_wallace_pg_rca8_and_0_3_y0;
  wire f_u_wallace_pg_rca8_ha1_y0;
  wire f_u_wallace_pg_rca8_ha1_y1;
  wire f_u_wallace_pg_rca8_and_2_2_a_2;
  wire f_u_wallace_pg_rca8_and_2_2_b_2;
  wire f_u_wallace_pg_rca8_and_2_2_y0;
  wire f_u_wallace_pg_rca8_and_1_3_a_1;
  wire f_u_wallace_pg_rca8_and_1_3_b_3;
  wire f_u_wallace_pg_rca8_and_1_3_y0;
  wire f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_ha1_y1;
  wire f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_and_2_2_y0;
  wire f_u_wallace_pg_rca8_fa10_y0;
  wire f_u_wallace_pg_rca8_fa10_y1;
  wire f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_and_1_3_y0;
  wire f_u_wallace_pg_rca8_fa10_y2;
  wire f_u_wallace_pg_rca8_fa10_y3;
  wire f_u_wallace_pg_rca8_fa10_y4;
  wire f_u_wallace_pg_rca8_and_3_2_a_3;
  wire f_u_wallace_pg_rca8_and_3_2_b_2;
  wire f_u_wallace_pg_rca8_and_3_2_y0;
  wire f_u_wallace_pg_rca8_and_2_3_a_2;
  wire f_u_wallace_pg_rca8_and_2_3_b_3;
  wire f_u_wallace_pg_rca8_and_2_3_y0;
  wire f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_fa10_y4;
  wire f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_and_3_2_y0;
  wire f_u_wallace_pg_rca8_fa11_y0;
  wire f_u_wallace_pg_rca8_fa11_y1;
  wire f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_and_2_3_y0;
  wire f_u_wallace_pg_rca8_fa11_y2;
  wire f_u_wallace_pg_rca8_fa11_y3;
  wire f_u_wallace_pg_rca8_fa11_y4;
  wire f_u_wallace_pg_rca8_and_4_2_a_4;
  wire f_u_wallace_pg_rca8_and_4_2_b_2;
  wire f_u_wallace_pg_rca8_and_4_2_y0;
  wire f_u_wallace_pg_rca8_and_3_3_a_3;
  wire f_u_wallace_pg_rca8_and_3_3_b_3;
  wire f_u_wallace_pg_rca8_and_3_3_y0;
  wire f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_fa11_y4;
  wire f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_and_4_2_y0;
  wire f_u_wallace_pg_rca8_fa12_y0;
  wire f_u_wallace_pg_rca8_fa12_y1;
  wire f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_and_3_3_y0;
  wire f_u_wallace_pg_rca8_fa12_y2;
  wire f_u_wallace_pg_rca8_fa12_y3;
  wire f_u_wallace_pg_rca8_fa12_y4;
  wire f_u_wallace_pg_rca8_and_5_2_a_5;
  wire f_u_wallace_pg_rca8_and_5_2_b_2;
  wire f_u_wallace_pg_rca8_and_5_2_y0;
  wire f_u_wallace_pg_rca8_and_4_3_a_4;
  wire f_u_wallace_pg_rca8_and_4_3_b_3;
  wire f_u_wallace_pg_rca8_and_4_3_y0;
  wire f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_fa12_y4;
  wire f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_and_5_2_y0;
  wire f_u_wallace_pg_rca8_fa13_y0;
  wire f_u_wallace_pg_rca8_fa13_y1;
  wire f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_and_4_3_y0;
  wire f_u_wallace_pg_rca8_fa13_y2;
  wire f_u_wallace_pg_rca8_fa13_y3;
  wire f_u_wallace_pg_rca8_fa13_y4;
  wire f_u_wallace_pg_rca8_and_5_3_a_5;
  wire f_u_wallace_pg_rca8_and_5_3_b_3;
  wire f_u_wallace_pg_rca8_and_5_3_y0;
  wire f_u_wallace_pg_rca8_and_4_4_a_4;
  wire f_u_wallace_pg_rca8_and_4_4_b_4;
  wire f_u_wallace_pg_rca8_and_4_4_y0;
  wire f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_fa13_y4;
  wire f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_and_5_3_y0;
  wire f_u_wallace_pg_rca8_fa14_y0;
  wire f_u_wallace_pg_rca8_fa14_y1;
  wire f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_and_4_4_y0;
  wire f_u_wallace_pg_rca8_fa14_y2;
  wire f_u_wallace_pg_rca8_fa14_y3;
  wire f_u_wallace_pg_rca8_fa14_y4;
  wire f_u_wallace_pg_rca8_and_5_4_a_5;
  wire f_u_wallace_pg_rca8_and_5_4_b_4;
  wire f_u_wallace_pg_rca8_and_5_4_y0;
  wire f_u_wallace_pg_rca8_and_4_5_a_4;
  wire f_u_wallace_pg_rca8_and_4_5_b_5;
  wire f_u_wallace_pg_rca8_and_4_5_y0;
  wire f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_fa14_y4;
  wire f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_and_5_4_y0;
  wire f_u_wallace_pg_rca8_fa15_y0;
  wire f_u_wallace_pg_rca8_fa15_y1;
  wire f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_and_4_5_y0;
  wire f_u_wallace_pg_rca8_fa15_y2;
  wire f_u_wallace_pg_rca8_fa15_y3;
  wire f_u_wallace_pg_rca8_fa15_y4;
  wire f_u_wallace_pg_rca8_and_5_5_a_5;
  wire f_u_wallace_pg_rca8_and_5_5_b_5;
  wire f_u_wallace_pg_rca8_and_5_5_y0;
  wire f_u_wallace_pg_rca8_and_4_6_a_4;
  wire f_u_wallace_pg_rca8_and_4_6_b_6;
  wire f_u_wallace_pg_rca8_and_4_6_y0;
  wire f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_fa15_y4;
  wire f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_and_5_5_y0;
  wire f_u_wallace_pg_rca8_fa16_y0;
  wire f_u_wallace_pg_rca8_fa16_y1;
  wire f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_and_4_6_y0;
  wire f_u_wallace_pg_rca8_fa16_y2;
  wire f_u_wallace_pg_rca8_fa16_y3;
  wire f_u_wallace_pg_rca8_fa16_y4;
  wire f_u_wallace_pg_rca8_and_5_6_a_5;
  wire f_u_wallace_pg_rca8_and_5_6_b_6;
  wire f_u_wallace_pg_rca8_and_5_6_y0;
  wire f_u_wallace_pg_rca8_and_4_7_a_4;
  wire f_u_wallace_pg_rca8_and_4_7_b_7;
  wire f_u_wallace_pg_rca8_and_4_7_y0;
  wire f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_fa16_y4;
  wire f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_and_5_6_y0;
  wire f_u_wallace_pg_rca8_fa17_y0;
  wire f_u_wallace_pg_rca8_fa17_y1;
  wire f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_and_4_7_y0;
  wire f_u_wallace_pg_rca8_fa17_y2;
  wire f_u_wallace_pg_rca8_fa17_y3;
  wire f_u_wallace_pg_rca8_fa17_y4;
  wire f_u_wallace_pg_rca8_and_0_4_a_0;
  wire f_u_wallace_pg_rca8_and_0_4_b_4;
  wire f_u_wallace_pg_rca8_and_0_4_y0;
  wire f_u_wallace_pg_rca8_ha2_f_u_wallace_pg_rca8_and_0_4_y0;
  wire f_u_wallace_pg_rca8_ha2_f_u_wallace_pg_rca8_fa1_y2;
  wire f_u_wallace_pg_rca8_ha2_y0;
  wire f_u_wallace_pg_rca8_ha2_y1;
  wire f_u_wallace_pg_rca8_and_1_4_a_1;
  wire f_u_wallace_pg_rca8_and_1_4_b_4;
  wire f_u_wallace_pg_rca8_and_1_4_y0;
  wire f_u_wallace_pg_rca8_and_0_5_a_0;
  wire f_u_wallace_pg_rca8_and_0_5_b_5;
  wire f_u_wallace_pg_rca8_and_0_5_y0;
  wire f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_ha2_y1;
  wire f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_and_1_4_y0;
  wire f_u_wallace_pg_rca8_fa18_y0;
  wire f_u_wallace_pg_rca8_fa18_y1;
  wire f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_and_0_5_y0;
  wire f_u_wallace_pg_rca8_fa18_y2;
  wire f_u_wallace_pg_rca8_fa18_y3;
  wire f_u_wallace_pg_rca8_fa18_y4;
  wire f_u_wallace_pg_rca8_and_2_4_a_2;
  wire f_u_wallace_pg_rca8_and_2_4_b_4;
  wire f_u_wallace_pg_rca8_and_2_4_y0;
  wire f_u_wallace_pg_rca8_and_1_5_a_1;
  wire f_u_wallace_pg_rca8_and_1_5_b_5;
  wire f_u_wallace_pg_rca8_and_1_5_y0;
  wire f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_fa18_y4;
  wire f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_and_2_4_y0;
  wire f_u_wallace_pg_rca8_fa19_y0;
  wire f_u_wallace_pg_rca8_fa19_y1;
  wire f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_and_1_5_y0;
  wire f_u_wallace_pg_rca8_fa19_y2;
  wire f_u_wallace_pg_rca8_fa19_y3;
  wire f_u_wallace_pg_rca8_fa19_y4;
  wire f_u_wallace_pg_rca8_and_3_4_a_3;
  wire f_u_wallace_pg_rca8_and_3_4_b_4;
  wire f_u_wallace_pg_rca8_and_3_4_y0;
  wire f_u_wallace_pg_rca8_and_2_5_a_2;
  wire f_u_wallace_pg_rca8_and_2_5_b_5;
  wire f_u_wallace_pg_rca8_and_2_5_y0;
  wire f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_fa19_y4;
  wire f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_and_3_4_y0;
  wire f_u_wallace_pg_rca8_fa20_y0;
  wire f_u_wallace_pg_rca8_fa20_y1;
  wire f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_and_2_5_y0;
  wire f_u_wallace_pg_rca8_fa20_y2;
  wire f_u_wallace_pg_rca8_fa20_y3;
  wire f_u_wallace_pg_rca8_fa20_y4;
  wire f_u_wallace_pg_rca8_and_3_5_a_3;
  wire f_u_wallace_pg_rca8_and_3_5_b_5;
  wire f_u_wallace_pg_rca8_and_3_5_y0;
  wire f_u_wallace_pg_rca8_and_2_6_a_2;
  wire f_u_wallace_pg_rca8_and_2_6_b_6;
  wire f_u_wallace_pg_rca8_and_2_6_y0;
  wire f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_fa20_y4;
  wire f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_and_3_5_y0;
  wire f_u_wallace_pg_rca8_fa21_y0;
  wire f_u_wallace_pg_rca8_fa21_y1;
  wire f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_and_2_6_y0;
  wire f_u_wallace_pg_rca8_fa21_y2;
  wire f_u_wallace_pg_rca8_fa21_y3;
  wire f_u_wallace_pg_rca8_fa21_y4;
  wire f_u_wallace_pg_rca8_and_3_6_a_3;
  wire f_u_wallace_pg_rca8_and_3_6_b_6;
  wire f_u_wallace_pg_rca8_and_3_6_y0;
  wire f_u_wallace_pg_rca8_and_2_7_a_2;
  wire f_u_wallace_pg_rca8_and_2_7_b_7;
  wire f_u_wallace_pg_rca8_and_2_7_y0;
  wire f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_fa21_y4;
  wire f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_and_3_6_y0;
  wire f_u_wallace_pg_rca8_fa22_y0;
  wire f_u_wallace_pg_rca8_fa22_y1;
  wire f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_and_2_7_y0;
  wire f_u_wallace_pg_rca8_fa22_y2;
  wire f_u_wallace_pg_rca8_fa22_y3;
  wire f_u_wallace_pg_rca8_fa22_y4;
  wire f_u_wallace_pg_rca8_and_3_7_a_3;
  wire f_u_wallace_pg_rca8_and_3_7_b_7;
  wire f_u_wallace_pg_rca8_and_3_7_y0;
  wire f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_fa22_y4;
  wire f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_and_3_7_y0;
  wire f_u_wallace_pg_rca8_fa23_y0;
  wire f_u_wallace_pg_rca8_fa23_y1;
  wire f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_fa7_y2;
  wire f_u_wallace_pg_rca8_fa23_y2;
  wire f_u_wallace_pg_rca8_fa23_y3;
  wire f_u_wallace_pg_rca8_fa23_y4;
  wire f_u_wallace_pg_rca8_ha3_f_u_wallace_pg_rca8_fa2_y2;
  wire f_u_wallace_pg_rca8_ha3_f_u_wallace_pg_rca8_fa11_y2;
  wire f_u_wallace_pg_rca8_ha3_y0;
  wire f_u_wallace_pg_rca8_ha3_y1;
  wire f_u_wallace_pg_rca8_and_0_6_a_0;
  wire f_u_wallace_pg_rca8_and_0_6_b_6;
  wire f_u_wallace_pg_rca8_and_0_6_y0;
  wire f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_ha3_y1;
  wire f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_and_0_6_y0;
  wire f_u_wallace_pg_rca8_fa24_y0;
  wire f_u_wallace_pg_rca8_fa24_y1;
  wire f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_fa3_y2;
  wire f_u_wallace_pg_rca8_fa24_y2;
  wire f_u_wallace_pg_rca8_fa24_y3;
  wire f_u_wallace_pg_rca8_fa24_y4;
  wire f_u_wallace_pg_rca8_and_1_6_a_1;
  wire f_u_wallace_pg_rca8_and_1_6_b_6;
  wire f_u_wallace_pg_rca8_and_1_6_y0;
  wire f_u_wallace_pg_rca8_and_0_7_a_0;
  wire f_u_wallace_pg_rca8_and_0_7_b_7;
  wire f_u_wallace_pg_rca8_and_0_7_y0;
  wire f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_fa24_y4;
  wire f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_and_1_6_y0;
  wire f_u_wallace_pg_rca8_fa25_y0;
  wire f_u_wallace_pg_rca8_fa25_y1;
  wire f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_and_0_7_y0;
  wire f_u_wallace_pg_rca8_fa25_y2;
  wire f_u_wallace_pg_rca8_fa25_y3;
  wire f_u_wallace_pg_rca8_fa25_y4;
  wire f_u_wallace_pg_rca8_and_1_7_a_1;
  wire f_u_wallace_pg_rca8_and_1_7_b_7;
  wire f_u_wallace_pg_rca8_and_1_7_y0;
  wire f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_fa25_y4;
  wire f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_and_1_7_y0;
  wire f_u_wallace_pg_rca8_fa26_y0;
  wire f_u_wallace_pg_rca8_fa26_y1;
  wire f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_fa5_y2;
  wire f_u_wallace_pg_rca8_fa26_y2;
  wire f_u_wallace_pg_rca8_fa26_y3;
  wire f_u_wallace_pg_rca8_fa26_y4;
  wire f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa26_y4;
  wire f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa6_y2;
  wire f_u_wallace_pg_rca8_fa27_y0;
  wire f_u_wallace_pg_rca8_fa27_y1;
  wire f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa15_y2;
  wire f_u_wallace_pg_rca8_fa27_y2;
  wire f_u_wallace_pg_rca8_fa27_y3;
  wire f_u_wallace_pg_rca8_fa27_y4;
  wire f_u_wallace_pg_rca8_ha4_f_u_wallace_pg_rca8_fa12_y2;
  wire f_u_wallace_pg_rca8_ha4_f_u_wallace_pg_rca8_fa19_y2;
  wire f_u_wallace_pg_rca8_ha4_y0;
  wire f_u_wallace_pg_rca8_ha4_y1;
  wire f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_ha4_y1;
  wire f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_fa4_y2;
  wire f_u_wallace_pg_rca8_fa28_y0;
  wire f_u_wallace_pg_rca8_fa28_y1;
  wire f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_fa13_y2;
  wire f_u_wallace_pg_rca8_fa28_y2;
  wire f_u_wallace_pg_rca8_fa28_y3;
  wire f_u_wallace_pg_rca8_fa28_y4;
  wire f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa28_y4;
  wire f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa14_y2;
  wire f_u_wallace_pg_rca8_fa29_y0;
  wire f_u_wallace_pg_rca8_fa29_y1;
  wire f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa21_y2;
  wire f_u_wallace_pg_rca8_fa29_y2;
  wire f_u_wallace_pg_rca8_fa29_y3;
  wire f_u_wallace_pg_rca8_fa29_y4;
  wire f_u_wallace_pg_rca8_ha5_f_u_wallace_pg_rca8_fa20_y2;
  wire f_u_wallace_pg_rca8_ha5_f_u_wallace_pg_rca8_fa25_y2;
  wire f_u_wallace_pg_rca8_ha5_y0;
  wire f_u_wallace_pg_rca8_ha5_y1;
  wire f_u_wallace_pg_rca8_ha6_f_u_wallace_pg_rca8_ha5_y1;
  wire f_u_wallace_pg_rca8_ha6_f_u_wallace_pg_rca8_fa26_y2;
  wire f_u_wallace_pg_rca8_ha6_y0;
  wire f_u_wallace_pg_rca8_ha6_y1;
  wire f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_ha6_y1;
  wire f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_fa29_y4;
  wire f_u_wallace_pg_rca8_fa30_y0;
  wire f_u_wallace_pg_rca8_fa30_y1;
  wire f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_fa22_y2;
  wire f_u_wallace_pg_rca8_fa30_y2;
  wire f_u_wallace_pg_rca8_fa30_y3;
  wire f_u_wallace_pg_rca8_fa30_y4;
  wire f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa30_y4;
  wire f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa27_y4;
  wire f_u_wallace_pg_rca8_fa31_y0;
  wire f_u_wallace_pg_rca8_fa31_y1;
  wire f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa16_y2;
  wire f_u_wallace_pg_rca8_fa31_y2;
  wire f_u_wallace_pg_rca8_fa31_y3;
  wire f_u_wallace_pg_rca8_fa31_y4;
  wire f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa31_y4;
  wire f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa23_y4;
  wire f_u_wallace_pg_rca8_fa32_y0;
  wire f_u_wallace_pg_rca8_fa32_y1;
  wire f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa8_y2;
  wire f_u_wallace_pg_rca8_fa32_y2;
  wire f_u_wallace_pg_rca8_fa32_y3;
  wire f_u_wallace_pg_rca8_fa32_y4;
  wire f_u_wallace_pg_rca8_and_5_7_a_5;
  wire f_u_wallace_pg_rca8_and_5_7_b_7;
  wire f_u_wallace_pg_rca8_and_5_7_y0;
  wire f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_fa32_y4;
  wire f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_fa17_y4;
  wire f_u_wallace_pg_rca8_fa33_y0;
  wire f_u_wallace_pg_rca8_fa33_y1;
  wire f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_and_5_7_y0;
  wire f_u_wallace_pg_rca8_fa33_y2;
  wire f_u_wallace_pg_rca8_fa33_y3;
  wire f_u_wallace_pg_rca8_fa33_y4;
  wire f_u_wallace_pg_rca8_and_7_6_a_7;
  wire f_u_wallace_pg_rca8_and_7_6_b_6;
  wire f_u_wallace_pg_rca8_and_7_6_y0;
  wire f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_fa33_y4;
  wire f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_fa9_y4;
  wire f_u_wallace_pg_rca8_fa34_y0;
  wire f_u_wallace_pg_rca8_fa34_y1;
  wire f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_and_7_6_y0;
  wire f_u_wallace_pg_rca8_fa34_y2;
  wire f_u_wallace_pg_rca8_fa34_y3;
  wire f_u_wallace_pg_rca8_fa34_y4;
  wire f_u_wallace_pg_rca8_and_0_0_a_0;
  wire f_u_wallace_pg_rca8_and_0_0_b_0;
  wire f_u_wallace_pg_rca8_and_0_0_y0;
  wire f_u_wallace_pg_rca8_and_1_0_a_1;
  wire f_u_wallace_pg_rca8_and_1_0_b_0;
  wire f_u_wallace_pg_rca8_and_1_0_y0;
  wire f_u_wallace_pg_rca8_and_0_2_a_0;
  wire f_u_wallace_pg_rca8_and_0_2_b_2;
  wire f_u_wallace_pg_rca8_and_0_2_y0;
  wire f_u_wallace_pg_rca8_and_6_7_a_6;
  wire f_u_wallace_pg_rca8_and_6_7_b_7;
  wire f_u_wallace_pg_rca8_and_6_7_y0;
  wire f_u_wallace_pg_rca8_and_0_1_a_0;
  wire f_u_wallace_pg_rca8_and_0_1_b_1;
  wire f_u_wallace_pg_rca8_and_0_1_y0;
  wire f_u_wallace_pg_rca8_and_7_7_a_7;
  wire f_u_wallace_pg_rca8_and_7_7_b_7;
  wire f_u_wallace_pg_rca8_and_7_7_y0;
  wire constant_wire_value_0_f_u_wallace_pg_rca8_and_1_0_y0;
  wire constant_wire_value_0_f_u_wallace_pg_rca8_and_0_1_y0;
  wire constant_wire_value_0_y0;
  wire constant_wire_value_0_y1;
  wire constant_wire_0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa0_f_u_wallace_pg_rca8_and_1_0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa0_f_u_wallace_pg_rca8_and_0_1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa0_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa0_constant_wire_0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa0_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and0_constant_wire_0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and0_f_u_wallace_pg_rca8_u_pg_rca14_fa0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or0_f_u_wallace_pg_rca8_u_pg_rca14_and0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or0_f_u_wallace_pg_rca8_u_pg_rca14_fa0_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_and_0_2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_ha0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa1_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_u_pg_rca14_or0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa1_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and1_f_u_wallace_pg_rca8_u_pg_rca14_or0_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and1_f_u_wallace_pg_rca8_u_pg_rca14_fa1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or1_f_u_wallace_pg_rca8_u_pg_rca14_and1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or1_f_u_wallace_pg_rca8_u_pg_rca14_fa1_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_fa0_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_ha1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa2_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_u_pg_rca14_or1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa2_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and2_f_u_wallace_pg_rca8_u_pg_rca14_or1_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and2_f_u_wallace_pg_rca8_u_pg_rca14_fa2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or2_f_u_wallace_pg_rca8_u_pg_rca14_and2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or2_f_u_wallace_pg_rca8_u_pg_rca14_fa2_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_fa10_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_ha2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa3_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa3_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_u_pg_rca14_or2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa3_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and3_f_u_wallace_pg_rca8_u_pg_rca14_or2_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and3_f_u_wallace_pg_rca8_u_pg_rca14_fa3_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and3_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or3_f_u_wallace_pg_rca8_u_pg_rca14_and3_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or3_f_u_wallace_pg_rca8_u_pg_rca14_fa3_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or3_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_fa18_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_ha3_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa4_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa4_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_u_pg_rca14_or3_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa4_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and4_f_u_wallace_pg_rca8_u_pg_rca14_or3_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and4_f_u_wallace_pg_rca8_u_pg_rca14_fa4_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and4_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or4_f_u_wallace_pg_rca8_u_pg_rca14_and4_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or4_f_u_wallace_pg_rca8_u_pg_rca14_fa4_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or4_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_fa24_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_ha4_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa5_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa5_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_u_pg_rca14_or4_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa5_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and5_f_u_wallace_pg_rca8_u_pg_rca14_or4_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and5_f_u_wallace_pg_rca8_u_pg_rca14_fa5_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and5_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or5_f_u_wallace_pg_rca8_u_pg_rca14_and5_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or5_f_u_wallace_pg_rca8_u_pg_rca14_fa5_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or5_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_fa28_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_ha5_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa6_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa6_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_u_pg_rca14_or5_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa6_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and6_f_u_wallace_pg_rca8_u_pg_rca14_or5_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and6_f_u_wallace_pg_rca8_u_pg_rca14_fa6_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and6_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or6_f_u_wallace_pg_rca8_u_pg_rca14_and6_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or6_f_u_wallace_pg_rca8_u_pg_rca14_fa6_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or6_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_fa29_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_ha6_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa7_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_u_pg_rca14_or6_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa7_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and7_f_u_wallace_pg_rca8_u_pg_rca14_or6_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and7_f_u_wallace_pg_rca8_u_pg_rca14_fa7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or7_f_u_wallace_pg_rca8_u_pg_rca14_and7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or7_f_u_wallace_pg_rca8_u_pg_rca14_fa7_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_fa27_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_fa30_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa8_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa8_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_u_pg_rca14_or7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa8_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and8_f_u_wallace_pg_rca8_u_pg_rca14_or7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and8_f_u_wallace_pg_rca8_u_pg_rca14_fa8_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and8_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or8_f_u_wallace_pg_rca8_u_pg_rca14_and8_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or8_f_u_wallace_pg_rca8_u_pg_rca14_fa8_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or8_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_fa23_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_fa31_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa9_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa9_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_u_pg_rca14_or8_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa9_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and9_f_u_wallace_pg_rca8_u_pg_rca14_or8_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and9_f_u_wallace_pg_rca8_u_pg_rca14_fa9_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and9_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or9_f_u_wallace_pg_rca8_u_pg_rca14_and9_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or9_f_u_wallace_pg_rca8_u_pg_rca14_fa9_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or9_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_fa17_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_fa32_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa10_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa10_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_u_pg_rca14_or9_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa10_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and10_f_u_wallace_pg_rca8_u_pg_rca14_or9_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and10_f_u_wallace_pg_rca8_u_pg_rca14_fa10_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and10_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or10_f_u_wallace_pg_rca8_u_pg_rca14_and10_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or10_f_u_wallace_pg_rca8_u_pg_rca14_fa10_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or10_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_fa9_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_fa33_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa11_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa11_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_u_pg_rca14_or10_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa11_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and11_f_u_wallace_pg_rca8_u_pg_rca14_or10_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and11_f_u_wallace_pg_rca8_u_pg_rca14_fa11_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and11_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or11_f_u_wallace_pg_rca8_u_pg_rca14_and11_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or11_f_u_wallace_pg_rca8_u_pg_rca14_fa11_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or11_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_and_6_7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_fa34_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa12_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa12_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_u_pg_rca14_or11_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa12_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and12_f_u_wallace_pg_rca8_u_pg_rca14_or11_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and12_f_u_wallace_pg_rca8_u_pg_rca14_fa12_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and12_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or12_f_u_wallace_pg_rca8_u_pg_rca14_and12_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or12_f_u_wallace_pg_rca8_u_pg_rca14_fa12_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or12_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_fa34_y4;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_and_7_7_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa13_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa13_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_u_pg_rca14_or12_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_fa13_y2;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and13_f_u_wallace_pg_rca8_u_pg_rca14_or12_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and13_f_u_wallace_pg_rca8_u_pg_rca14_fa13_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_and13_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or13_f_u_wallace_pg_rca8_u_pg_rca14_and13_y0;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or13_f_u_wallace_pg_rca8_u_pg_rca14_fa13_y1;
  wire f_u_wallace_pg_rca8_u_pg_rca14_or13_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign f_u_wallace_pg_rca8_and_2_0_a_2 = a_2;
  assign f_u_wallace_pg_rca8_and_2_0_b_0 = b_0;
  assign f_u_wallace_pg_rca8_and_2_0_y0 = f_u_wallace_pg_rca8_and_2_0_a_2 & f_u_wallace_pg_rca8_and_2_0_b_0;
  assign f_u_wallace_pg_rca8_and_1_1_a_1 = a_1;
  assign f_u_wallace_pg_rca8_and_1_1_b_1 = b_1;
  assign f_u_wallace_pg_rca8_and_1_1_y0 = f_u_wallace_pg_rca8_and_1_1_a_1 & f_u_wallace_pg_rca8_and_1_1_b_1;
  assign f_u_wallace_pg_rca8_ha0_f_u_wallace_pg_rca8_and_2_0_y0 = f_u_wallace_pg_rca8_and_2_0_y0;
  assign f_u_wallace_pg_rca8_ha0_f_u_wallace_pg_rca8_and_1_1_y0 = f_u_wallace_pg_rca8_and_1_1_y0;
  assign f_u_wallace_pg_rca8_ha0_y0 = f_u_wallace_pg_rca8_ha0_f_u_wallace_pg_rca8_and_2_0_y0 ^ f_u_wallace_pg_rca8_ha0_f_u_wallace_pg_rca8_and_1_1_y0;
  assign f_u_wallace_pg_rca8_ha0_y1 = f_u_wallace_pg_rca8_ha0_f_u_wallace_pg_rca8_and_2_0_y0 & f_u_wallace_pg_rca8_ha0_f_u_wallace_pg_rca8_and_1_1_y0;
  assign f_u_wallace_pg_rca8_and_3_0_a_3 = a_3;
  assign f_u_wallace_pg_rca8_and_3_0_b_0 = b_0;
  assign f_u_wallace_pg_rca8_and_3_0_y0 = f_u_wallace_pg_rca8_and_3_0_a_3 & f_u_wallace_pg_rca8_and_3_0_b_0;
  assign f_u_wallace_pg_rca8_and_2_1_a_2 = a_2;
  assign f_u_wallace_pg_rca8_and_2_1_b_1 = b_1;
  assign f_u_wallace_pg_rca8_and_2_1_y0 = f_u_wallace_pg_rca8_and_2_1_a_2 & f_u_wallace_pg_rca8_and_2_1_b_1;
  assign f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_ha0_y1 = f_u_wallace_pg_rca8_ha0_y1;
  assign f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_and_3_0_y0 = f_u_wallace_pg_rca8_and_3_0_y0;
  assign f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_and_2_1_y0 = f_u_wallace_pg_rca8_and_2_1_y0;
  assign f_u_wallace_pg_rca8_fa0_y0 = f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_ha0_y1 ^ f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_and_3_0_y0;
  assign f_u_wallace_pg_rca8_fa0_y1 = f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_ha0_y1 & f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_and_3_0_y0;
  assign f_u_wallace_pg_rca8_fa0_y2 = f_u_wallace_pg_rca8_fa0_y0 ^ f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_and_2_1_y0;
  assign f_u_wallace_pg_rca8_fa0_y3 = f_u_wallace_pg_rca8_fa0_y0 & f_u_wallace_pg_rca8_fa0_f_u_wallace_pg_rca8_and_2_1_y0;
  assign f_u_wallace_pg_rca8_fa0_y4 = f_u_wallace_pg_rca8_fa0_y1 | f_u_wallace_pg_rca8_fa0_y3;
  assign f_u_wallace_pg_rca8_and_4_0_a_4 = a_4;
  assign f_u_wallace_pg_rca8_and_4_0_b_0 = b_0;
  assign f_u_wallace_pg_rca8_and_4_0_y0 = f_u_wallace_pg_rca8_and_4_0_a_4 & f_u_wallace_pg_rca8_and_4_0_b_0;
  assign f_u_wallace_pg_rca8_and_3_1_a_3 = a_3;
  assign f_u_wallace_pg_rca8_and_3_1_b_1 = b_1;
  assign f_u_wallace_pg_rca8_and_3_1_y0 = f_u_wallace_pg_rca8_and_3_1_a_3 & f_u_wallace_pg_rca8_and_3_1_b_1;
  assign f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_fa0_y4 = f_u_wallace_pg_rca8_fa0_y4;
  assign f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_and_4_0_y0 = f_u_wallace_pg_rca8_and_4_0_y0;
  assign f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_and_3_1_y0 = f_u_wallace_pg_rca8_and_3_1_y0;
  assign f_u_wallace_pg_rca8_fa1_y0 = f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_fa0_y4 ^ f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_and_4_0_y0;
  assign f_u_wallace_pg_rca8_fa1_y1 = f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_fa0_y4 & f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_and_4_0_y0;
  assign f_u_wallace_pg_rca8_fa1_y2 = f_u_wallace_pg_rca8_fa1_y0 ^ f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_and_3_1_y0;
  assign f_u_wallace_pg_rca8_fa1_y3 = f_u_wallace_pg_rca8_fa1_y0 & f_u_wallace_pg_rca8_fa1_f_u_wallace_pg_rca8_and_3_1_y0;
  assign f_u_wallace_pg_rca8_fa1_y4 = f_u_wallace_pg_rca8_fa1_y1 | f_u_wallace_pg_rca8_fa1_y3;
  assign f_u_wallace_pg_rca8_and_5_0_a_5 = a_5;
  assign f_u_wallace_pg_rca8_and_5_0_b_0 = b_0;
  assign f_u_wallace_pg_rca8_and_5_0_y0 = f_u_wallace_pg_rca8_and_5_0_a_5 & f_u_wallace_pg_rca8_and_5_0_b_0;
  assign f_u_wallace_pg_rca8_and_4_1_a_4 = a_4;
  assign f_u_wallace_pg_rca8_and_4_1_b_1 = b_1;
  assign f_u_wallace_pg_rca8_and_4_1_y0 = f_u_wallace_pg_rca8_and_4_1_a_4 & f_u_wallace_pg_rca8_and_4_1_b_1;
  assign f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_fa1_y4 = f_u_wallace_pg_rca8_fa1_y4;
  assign f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_and_5_0_y0 = f_u_wallace_pg_rca8_and_5_0_y0;
  assign f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_and_4_1_y0 = f_u_wallace_pg_rca8_and_4_1_y0;
  assign f_u_wallace_pg_rca8_fa2_y0 = f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_fa1_y4 ^ f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_and_5_0_y0;
  assign f_u_wallace_pg_rca8_fa2_y1 = f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_fa1_y4 & f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_and_5_0_y0;
  assign f_u_wallace_pg_rca8_fa2_y2 = f_u_wallace_pg_rca8_fa2_y0 ^ f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_and_4_1_y0;
  assign f_u_wallace_pg_rca8_fa2_y3 = f_u_wallace_pg_rca8_fa2_y0 & f_u_wallace_pg_rca8_fa2_f_u_wallace_pg_rca8_and_4_1_y0;
  assign f_u_wallace_pg_rca8_fa2_y4 = f_u_wallace_pg_rca8_fa2_y1 | f_u_wallace_pg_rca8_fa2_y3;
  assign f_u_wallace_pg_rca8_and_6_0_a_6 = a_6;
  assign f_u_wallace_pg_rca8_and_6_0_b_0 = b_0;
  assign f_u_wallace_pg_rca8_and_6_0_y0 = f_u_wallace_pg_rca8_and_6_0_a_6 & f_u_wallace_pg_rca8_and_6_0_b_0;
  assign f_u_wallace_pg_rca8_and_5_1_a_5 = a_5;
  assign f_u_wallace_pg_rca8_and_5_1_b_1 = b_1;
  assign f_u_wallace_pg_rca8_and_5_1_y0 = f_u_wallace_pg_rca8_and_5_1_a_5 & f_u_wallace_pg_rca8_and_5_1_b_1;
  assign f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_fa2_y4 = f_u_wallace_pg_rca8_fa2_y4;
  assign f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_and_6_0_y0 = f_u_wallace_pg_rca8_and_6_0_y0;
  assign f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_and_5_1_y0 = f_u_wallace_pg_rca8_and_5_1_y0;
  assign f_u_wallace_pg_rca8_fa3_y0 = f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_fa2_y4 ^ f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_and_6_0_y0;
  assign f_u_wallace_pg_rca8_fa3_y1 = f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_fa2_y4 & f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_and_6_0_y0;
  assign f_u_wallace_pg_rca8_fa3_y2 = f_u_wallace_pg_rca8_fa3_y0 ^ f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_and_5_1_y0;
  assign f_u_wallace_pg_rca8_fa3_y3 = f_u_wallace_pg_rca8_fa3_y0 & f_u_wallace_pg_rca8_fa3_f_u_wallace_pg_rca8_and_5_1_y0;
  assign f_u_wallace_pg_rca8_fa3_y4 = f_u_wallace_pg_rca8_fa3_y1 | f_u_wallace_pg_rca8_fa3_y3;
  assign f_u_wallace_pg_rca8_and_7_0_a_7 = a_7;
  assign f_u_wallace_pg_rca8_and_7_0_b_0 = b_0;
  assign f_u_wallace_pg_rca8_and_7_0_y0 = f_u_wallace_pg_rca8_and_7_0_a_7 & f_u_wallace_pg_rca8_and_7_0_b_0;
  assign f_u_wallace_pg_rca8_and_6_1_a_6 = a_6;
  assign f_u_wallace_pg_rca8_and_6_1_b_1 = b_1;
  assign f_u_wallace_pg_rca8_and_6_1_y0 = f_u_wallace_pg_rca8_and_6_1_a_6 & f_u_wallace_pg_rca8_and_6_1_b_1;
  assign f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_fa3_y4 = f_u_wallace_pg_rca8_fa3_y4;
  assign f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_and_7_0_y0 = f_u_wallace_pg_rca8_and_7_0_y0;
  assign f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_and_6_1_y0 = f_u_wallace_pg_rca8_and_6_1_y0;
  assign f_u_wallace_pg_rca8_fa4_y0 = f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_fa3_y4 ^ f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_and_7_0_y0;
  assign f_u_wallace_pg_rca8_fa4_y1 = f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_fa3_y4 & f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_and_7_0_y0;
  assign f_u_wallace_pg_rca8_fa4_y2 = f_u_wallace_pg_rca8_fa4_y0 ^ f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_and_6_1_y0;
  assign f_u_wallace_pg_rca8_fa4_y3 = f_u_wallace_pg_rca8_fa4_y0 & f_u_wallace_pg_rca8_fa4_f_u_wallace_pg_rca8_and_6_1_y0;
  assign f_u_wallace_pg_rca8_fa4_y4 = f_u_wallace_pg_rca8_fa4_y1 | f_u_wallace_pg_rca8_fa4_y3;
  assign f_u_wallace_pg_rca8_and_7_1_a_7 = a_7;
  assign f_u_wallace_pg_rca8_and_7_1_b_1 = b_1;
  assign f_u_wallace_pg_rca8_and_7_1_y0 = f_u_wallace_pg_rca8_and_7_1_a_7 & f_u_wallace_pg_rca8_and_7_1_b_1;
  assign f_u_wallace_pg_rca8_and_6_2_a_6 = a_6;
  assign f_u_wallace_pg_rca8_and_6_2_b_2 = b_2;
  assign f_u_wallace_pg_rca8_and_6_2_y0 = f_u_wallace_pg_rca8_and_6_2_a_6 & f_u_wallace_pg_rca8_and_6_2_b_2;
  assign f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_fa4_y4 = f_u_wallace_pg_rca8_fa4_y4;
  assign f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_and_7_1_y0 = f_u_wallace_pg_rca8_and_7_1_y0;
  assign f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_and_6_2_y0 = f_u_wallace_pg_rca8_and_6_2_y0;
  assign f_u_wallace_pg_rca8_fa5_y0 = f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_fa4_y4 ^ f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_and_7_1_y0;
  assign f_u_wallace_pg_rca8_fa5_y1 = f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_fa4_y4 & f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_and_7_1_y0;
  assign f_u_wallace_pg_rca8_fa5_y2 = f_u_wallace_pg_rca8_fa5_y0 ^ f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_and_6_2_y0;
  assign f_u_wallace_pg_rca8_fa5_y3 = f_u_wallace_pg_rca8_fa5_y0 & f_u_wallace_pg_rca8_fa5_f_u_wallace_pg_rca8_and_6_2_y0;
  assign f_u_wallace_pg_rca8_fa5_y4 = f_u_wallace_pg_rca8_fa5_y1 | f_u_wallace_pg_rca8_fa5_y3;
  assign f_u_wallace_pg_rca8_and_7_2_a_7 = a_7;
  assign f_u_wallace_pg_rca8_and_7_2_b_2 = b_2;
  assign f_u_wallace_pg_rca8_and_7_2_y0 = f_u_wallace_pg_rca8_and_7_2_a_7 & f_u_wallace_pg_rca8_and_7_2_b_2;
  assign f_u_wallace_pg_rca8_and_6_3_a_6 = a_6;
  assign f_u_wallace_pg_rca8_and_6_3_b_3 = b_3;
  assign f_u_wallace_pg_rca8_and_6_3_y0 = f_u_wallace_pg_rca8_and_6_3_a_6 & f_u_wallace_pg_rca8_and_6_3_b_3;
  assign f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_fa5_y4 = f_u_wallace_pg_rca8_fa5_y4;
  assign f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_and_7_2_y0 = f_u_wallace_pg_rca8_and_7_2_y0;
  assign f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_and_6_3_y0 = f_u_wallace_pg_rca8_and_6_3_y0;
  assign f_u_wallace_pg_rca8_fa6_y0 = f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_fa5_y4 ^ f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_and_7_2_y0;
  assign f_u_wallace_pg_rca8_fa6_y1 = f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_fa5_y4 & f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_and_7_2_y0;
  assign f_u_wallace_pg_rca8_fa6_y2 = f_u_wallace_pg_rca8_fa6_y0 ^ f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_and_6_3_y0;
  assign f_u_wallace_pg_rca8_fa6_y3 = f_u_wallace_pg_rca8_fa6_y0 & f_u_wallace_pg_rca8_fa6_f_u_wallace_pg_rca8_and_6_3_y0;
  assign f_u_wallace_pg_rca8_fa6_y4 = f_u_wallace_pg_rca8_fa6_y1 | f_u_wallace_pg_rca8_fa6_y3;
  assign f_u_wallace_pg_rca8_and_7_3_a_7 = a_7;
  assign f_u_wallace_pg_rca8_and_7_3_b_3 = b_3;
  assign f_u_wallace_pg_rca8_and_7_3_y0 = f_u_wallace_pg_rca8_and_7_3_a_7 & f_u_wallace_pg_rca8_and_7_3_b_3;
  assign f_u_wallace_pg_rca8_and_6_4_a_6 = a_6;
  assign f_u_wallace_pg_rca8_and_6_4_b_4 = b_4;
  assign f_u_wallace_pg_rca8_and_6_4_y0 = f_u_wallace_pg_rca8_and_6_4_a_6 & f_u_wallace_pg_rca8_and_6_4_b_4;
  assign f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_fa6_y4 = f_u_wallace_pg_rca8_fa6_y4;
  assign f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_and_7_3_y0 = f_u_wallace_pg_rca8_and_7_3_y0;
  assign f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_and_6_4_y0 = f_u_wallace_pg_rca8_and_6_4_y0;
  assign f_u_wallace_pg_rca8_fa7_y0 = f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_fa6_y4 ^ f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_and_7_3_y0;
  assign f_u_wallace_pg_rca8_fa7_y1 = f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_fa6_y4 & f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_and_7_3_y0;
  assign f_u_wallace_pg_rca8_fa7_y2 = f_u_wallace_pg_rca8_fa7_y0 ^ f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_and_6_4_y0;
  assign f_u_wallace_pg_rca8_fa7_y3 = f_u_wallace_pg_rca8_fa7_y0 & f_u_wallace_pg_rca8_fa7_f_u_wallace_pg_rca8_and_6_4_y0;
  assign f_u_wallace_pg_rca8_fa7_y4 = f_u_wallace_pg_rca8_fa7_y1 | f_u_wallace_pg_rca8_fa7_y3;
  assign f_u_wallace_pg_rca8_and_7_4_a_7 = a_7;
  assign f_u_wallace_pg_rca8_and_7_4_b_4 = b_4;
  assign f_u_wallace_pg_rca8_and_7_4_y0 = f_u_wallace_pg_rca8_and_7_4_a_7 & f_u_wallace_pg_rca8_and_7_4_b_4;
  assign f_u_wallace_pg_rca8_and_6_5_a_6 = a_6;
  assign f_u_wallace_pg_rca8_and_6_5_b_5 = b_5;
  assign f_u_wallace_pg_rca8_and_6_5_y0 = f_u_wallace_pg_rca8_and_6_5_a_6 & f_u_wallace_pg_rca8_and_6_5_b_5;
  assign f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_fa7_y4 = f_u_wallace_pg_rca8_fa7_y4;
  assign f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_and_7_4_y0 = f_u_wallace_pg_rca8_and_7_4_y0;
  assign f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_and_6_5_y0 = f_u_wallace_pg_rca8_and_6_5_y0;
  assign f_u_wallace_pg_rca8_fa8_y0 = f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_fa7_y4 ^ f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_and_7_4_y0;
  assign f_u_wallace_pg_rca8_fa8_y1 = f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_fa7_y4 & f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_and_7_4_y0;
  assign f_u_wallace_pg_rca8_fa8_y2 = f_u_wallace_pg_rca8_fa8_y0 ^ f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_and_6_5_y0;
  assign f_u_wallace_pg_rca8_fa8_y3 = f_u_wallace_pg_rca8_fa8_y0 & f_u_wallace_pg_rca8_fa8_f_u_wallace_pg_rca8_and_6_5_y0;
  assign f_u_wallace_pg_rca8_fa8_y4 = f_u_wallace_pg_rca8_fa8_y1 | f_u_wallace_pg_rca8_fa8_y3;
  assign f_u_wallace_pg_rca8_and_7_5_a_7 = a_7;
  assign f_u_wallace_pg_rca8_and_7_5_b_5 = b_5;
  assign f_u_wallace_pg_rca8_and_7_5_y0 = f_u_wallace_pg_rca8_and_7_5_a_7 & f_u_wallace_pg_rca8_and_7_5_b_5;
  assign f_u_wallace_pg_rca8_and_6_6_a_6 = a_6;
  assign f_u_wallace_pg_rca8_and_6_6_b_6 = b_6;
  assign f_u_wallace_pg_rca8_and_6_6_y0 = f_u_wallace_pg_rca8_and_6_6_a_6 & f_u_wallace_pg_rca8_and_6_6_b_6;
  assign f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_fa8_y4 = f_u_wallace_pg_rca8_fa8_y4;
  assign f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_and_7_5_y0 = f_u_wallace_pg_rca8_and_7_5_y0;
  assign f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_and_6_6_y0 = f_u_wallace_pg_rca8_and_6_6_y0;
  assign f_u_wallace_pg_rca8_fa9_y0 = f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_fa8_y4 ^ f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_and_7_5_y0;
  assign f_u_wallace_pg_rca8_fa9_y1 = f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_fa8_y4 & f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_and_7_5_y0;
  assign f_u_wallace_pg_rca8_fa9_y2 = f_u_wallace_pg_rca8_fa9_y0 ^ f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_and_6_6_y0;
  assign f_u_wallace_pg_rca8_fa9_y3 = f_u_wallace_pg_rca8_fa9_y0 & f_u_wallace_pg_rca8_fa9_f_u_wallace_pg_rca8_and_6_6_y0;
  assign f_u_wallace_pg_rca8_fa9_y4 = f_u_wallace_pg_rca8_fa9_y1 | f_u_wallace_pg_rca8_fa9_y3;
  assign f_u_wallace_pg_rca8_and_1_2_a_1 = a_1;
  assign f_u_wallace_pg_rca8_and_1_2_b_2 = b_2;
  assign f_u_wallace_pg_rca8_and_1_2_y0 = f_u_wallace_pg_rca8_and_1_2_a_1 & f_u_wallace_pg_rca8_and_1_2_b_2;
  assign f_u_wallace_pg_rca8_and_0_3_a_0 = a_0;
  assign f_u_wallace_pg_rca8_and_0_3_b_3 = b_3;
  assign f_u_wallace_pg_rca8_and_0_3_y0 = f_u_wallace_pg_rca8_and_0_3_a_0 & f_u_wallace_pg_rca8_and_0_3_b_3;
  assign f_u_wallace_pg_rca8_ha1_f_u_wallace_pg_rca8_and_1_2_y0 = f_u_wallace_pg_rca8_and_1_2_y0;
  assign f_u_wallace_pg_rca8_ha1_f_u_wallace_pg_rca8_and_0_3_y0 = f_u_wallace_pg_rca8_and_0_3_y0;
  assign f_u_wallace_pg_rca8_ha1_y0 = f_u_wallace_pg_rca8_ha1_f_u_wallace_pg_rca8_and_1_2_y0 ^ f_u_wallace_pg_rca8_ha1_f_u_wallace_pg_rca8_and_0_3_y0;
  assign f_u_wallace_pg_rca8_ha1_y1 = f_u_wallace_pg_rca8_ha1_f_u_wallace_pg_rca8_and_1_2_y0 & f_u_wallace_pg_rca8_ha1_f_u_wallace_pg_rca8_and_0_3_y0;
  assign f_u_wallace_pg_rca8_and_2_2_a_2 = a_2;
  assign f_u_wallace_pg_rca8_and_2_2_b_2 = b_2;
  assign f_u_wallace_pg_rca8_and_2_2_y0 = f_u_wallace_pg_rca8_and_2_2_a_2 & f_u_wallace_pg_rca8_and_2_2_b_2;
  assign f_u_wallace_pg_rca8_and_1_3_a_1 = a_1;
  assign f_u_wallace_pg_rca8_and_1_3_b_3 = b_3;
  assign f_u_wallace_pg_rca8_and_1_3_y0 = f_u_wallace_pg_rca8_and_1_3_a_1 & f_u_wallace_pg_rca8_and_1_3_b_3;
  assign f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_ha1_y1 = f_u_wallace_pg_rca8_ha1_y1;
  assign f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_and_2_2_y0 = f_u_wallace_pg_rca8_and_2_2_y0;
  assign f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_and_1_3_y0 = f_u_wallace_pg_rca8_and_1_3_y0;
  assign f_u_wallace_pg_rca8_fa10_y0 = f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_ha1_y1 ^ f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_and_2_2_y0;
  assign f_u_wallace_pg_rca8_fa10_y1 = f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_ha1_y1 & f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_and_2_2_y0;
  assign f_u_wallace_pg_rca8_fa10_y2 = f_u_wallace_pg_rca8_fa10_y0 ^ f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_and_1_3_y0;
  assign f_u_wallace_pg_rca8_fa10_y3 = f_u_wallace_pg_rca8_fa10_y0 & f_u_wallace_pg_rca8_fa10_f_u_wallace_pg_rca8_and_1_3_y0;
  assign f_u_wallace_pg_rca8_fa10_y4 = f_u_wallace_pg_rca8_fa10_y1 | f_u_wallace_pg_rca8_fa10_y3;
  assign f_u_wallace_pg_rca8_and_3_2_a_3 = a_3;
  assign f_u_wallace_pg_rca8_and_3_2_b_2 = b_2;
  assign f_u_wallace_pg_rca8_and_3_2_y0 = f_u_wallace_pg_rca8_and_3_2_a_3 & f_u_wallace_pg_rca8_and_3_2_b_2;
  assign f_u_wallace_pg_rca8_and_2_3_a_2 = a_2;
  assign f_u_wallace_pg_rca8_and_2_3_b_3 = b_3;
  assign f_u_wallace_pg_rca8_and_2_3_y0 = f_u_wallace_pg_rca8_and_2_3_a_2 & f_u_wallace_pg_rca8_and_2_3_b_3;
  assign f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_fa10_y4 = f_u_wallace_pg_rca8_fa10_y4;
  assign f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_and_3_2_y0 = f_u_wallace_pg_rca8_and_3_2_y0;
  assign f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_and_2_3_y0 = f_u_wallace_pg_rca8_and_2_3_y0;
  assign f_u_wallace_pg_rca8_fa11_y0 = f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_fa10_y4 ^ f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_and_3_2_y0;
  assign f_u_wallace_pg_rca8_fa11_y1 = f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_fa10_y4 & f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_and_3_2_y0;
  assign f_u_wallace_pg_rca8_fa11_y2 = f_u_wallace_pg_rca8_fa11_y0 ^ f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_and_2_3_y0;
  assign f_u_wallace_pg_rca8_fa11_y3 = f_u_wallace_pg_rca8_fa11_y0 & f_u_wallace_pg_rca8_fa11_f_u_wallace_pg_rca8_and_2_3_y0;
  assign f_u_wallace_pg_rca8_fa11_y4 = f_u_wallace_pg_rca8_fa11_y1 | f_u_wallace_pg_rca8_fa11_y3;
  assign f_u_wallace_pg_rca8_and_4_2_a_4 = a_4;
  assign f_u_wallace_pg_rca8_and_4_2_b_2 = b_2;
  assign f_u_wallace_pg_rca8_and_4_2_y0 = f_u_wallace_pg_rca8_and_4_2_a_4 & f_u_wallace_pg_rca8_and_4_2_b_2;
  assign f_u_wallace_pg_rca8_and_3_3_a_3 = a_3;
  assign f_u_wallace_pg_rca8_and_3_3_b_3 = b_3;
  assign f_u_wallace_pg_rca8_and_3_3_y0 = f_u_wallace_pg_rca8_and_3_3_a_3 & f_u_wallace_pg_rca8_and_3_3_b_3;
  assign f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_fa11_y4 = f_u_wallace_pg_rca8_fa11_y4;
  assign f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_and_4_2_y0 = f_u_wallace_pg_rca8_and_4_2_y0;
  assign f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_and_3_3_y0 = f_u_wallace_pg_rca8_and_3_3_y0;
  assign f_u_wallace_pg_rca8_fa12_y0 = f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_fa11_y4 ^ f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_and_4_2_y0;
  assign f_u_wallace_pg_rca8_fa12_y1 = f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_fa11_y4 & f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_and_4_2_y0;
  assign f_u_wallace_pg_rca8_fa12_y2 = f_u_wallace_pg_rca8_fa12_y0 ^ f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_and_3_3_y0;
  assign f_u_wallace_pg_rca8_fa12_y3 = f_u_wallace_pg_rca8_fa12_y0 & f_u_wallace_pg_rca8_fa12_f_u_wallace_pg_rca8_and_3_3_y0;
  assign f_u_wallace_pg_rca8_fa12_y4 = f_u_wallace_pg_rca8_fa12_y1 | f_u_wallace_pg_rca8_fa12_y3;
  assign f_u_wallace_pg_rca8_and_5_2_a_5 = a_5;
  assign f_u_wallace_pg_rca8_and_5_2_b_2 = b_2;
  assign f_u_wallace_pg_rca8_and_5_2_y0 = f_u_wallace_pg_rca8_and_5_2_a_5 & f_u_wallace_pg_rca8_and_5_2_b_2;
  assign f_u_wallace_pg_rca8_and_4_3_a_4 = a_4;
  assign f_u_wallace_pg_rca8_and_4_3_b_3 = b_3;
  assign f_u_wallace_pg_rca8_and_4_3_y0 = f_u_wallace_pg_rca8_and_4_3_a_4 & f_u_wallace_pg_rca8_and_4_3_b_3;
  assign f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_fa12_y4 = f_u_wallace_pg_rca8_fa12_y4;
  assign f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_and_5_2_y0 = f_u_wallace_pg_rca8_and_5_2_y0;
  assign f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_and_4_3_y0 = f_u_wallace_pg_rca8_and_4_3_y0;
  assign f_u_wallace_pg_rca8_fa13_y0 = f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_fa12_y4 ^ f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_and_5_2_y0;
  assign f_u_wallace_pg_rca8_fa13_y1 = f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_fa12_y4 & f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_and_5_2_y0;
  assign f_u_wallace_pg_rca8_fa13_y2 = f_u_wallace_pg_rca8_fa13_y0 ^ f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_and_4_3_y0;
  assign f_u_wallace_pg_rca8_fa13_y3 = f_u_wallace_pg_rca8_fa13_y0 & f_u_wallace_pg_rca8_fa13_f_u_wallace_pg_rca8_and_4_3_y0;
  assign f_u_wallace_pg_rca8_fa13_y4 = f_u_wallace_pg_rca8_fa13_y1 | f_u_wallace_pg_rca8_fa13_y3;
  assign f_u_wallace_pg_rca8_and_5_3_a_5 = a_5;
  assign f_u_wallace_pg_rca8_and_5_3_b_3 = b_3;
  assign f_u_wallace_pg_rca8_and_5_3_y0 = f_u_wallace_pg_rca8_and_5_3_a_5 & f_u_wallace_pg_rca8_and_5_3_b_3;
  assign f_u_wallace_pg_rca8_and_4_4_a_4 = a_4;
  assign f_u_wallace_pg_rca8_and_4_4_b_4 = b_4;
  assign f_u_wallace_pg_rca8_and_4_4_y0 = f_u_wallace_pg_rca8_and_4_4_a_4 & f_u_wallace_pg_rca8_and_4_4_b_4;
  assign f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_fa13_y4 = f_u_wallace_pg_rca8_fa13_y4;
  assign f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_and_5_3_y0 = f_u_wallace_pg_rca8_and_5_3_y0;
  assign f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_and_4_4_y0 = f_u_wallace_pg_rca8_and_4_4_y0;
  assign f_u_wallace_pg_rca8_fa14_y0 = f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_fa13_y4 ^ f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_and_5_3_y0;
  assign f_u_wallace_pg_rca8_fa14_y1 = f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_fa13_y4 & f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_and_5_3_y0;
  assign f_u_wallace_pg_rca8_fa14_y2 = f_u_wallace_pg_rca8_fa14_y0 ^ f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_and_4_4_y0;
  assign f_u_wallace_pg_rca8_fa14_y3 = f_u_wallace_pg_rca8_fa14_y0 & f_u_wallace_pg_rca8_fa14_f_u_wallace_pg_rca8_and_4_4_y0;
  assign f_u_wallace_pg_rca8_fa14_y4 = f_u_wallace_pg_rca8_fa14_y1 | f_u_wallace_pg_rca8_fa14_y3;
  assign f_u_wallace_pg_rca8_and_5_4_a_5 = a_5;
  assign f_u_wallace_pg_rca8_and_5_4_b_4 = b_4;
  assign f_u_wallace_pg_rca8_and_5_4_y0 = f_u_wallace_pg_rca8_and_5_4_a_5 & f_u_wallace_pg_rca8_and_5_4_b_4;
  assign f_u_wallace_pg_rca8_and_4_5_a_4 = a_4;
  assign f_u_wallace_pg_rca8_and_4_5_b_5 = b_5;
  assign f_u_wallace_pg_rca8_and_4_5_y0 = f_u_wallace_pg_rca8_and_4_5_a_4 & f_u_wallace_pg_rca8_and_4_5_b_5;
  assign f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_fa14_y4 = f_u_wallace_pg_rca8_fa14_y4;
  assign f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_and_5_4_y0 = f_u_wallace_pg_rca8_and_5_4_y0;
  assign f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_and_4_5_y0 = f_u_wallace_pg_rca8_and_4_5_y0;
  assign f_u_wallace_pg_rca8_fa15_y0 = f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_fa14_y4 ^ f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_and_5_4_y0;
  assign f_u_wallace_pg_rca8_fa15_y1 = f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_fa14_y4 & f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_and_5_4_y0;
  assign f_u_wallace_pg_rca8_fa15_y2 = f_u_wallace_pg_rca8_fa15_y0 ^ f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_and_4_5_y0;
  assign f_u_wallace_pg_rca8_fa15_y3 = f_u_wallace_pg_rca8_fa15_y0 & f_u_wallace_pg_rca8_fa15_f_u_wallace_pg_rca8_and_4_5_y0;
  assign f_u_wallace_pg_rca8_fa15_y4 = f_u_wallace_pg_rca8_fa15_y1 | f_u_wallace_pg_rca8_fa15_y3;
  assign f_u_wallace_pg_rca8_and_5_5_a_5 = a_5;
  assign f_u_wallace_pg_rca8_and_5_5_b_5 = b_5;
  assign f_u_wallace_pg_rca8_and_5_5_y0 = f_u_wallace_pg_rca8_and_5_5_a_5 & f_u_wallace_pg_rca8_and_5_5_b_5;
  assign f_u_wallace_pg_rca8_and_4_6_a_4 = a_4;
  assign f_u_wallace_pg_rca8_and_4_6_b_6 = b_6;
  assign f_u_wallace_pg_rca8_and_4_6_y0 = f_u_wallace_pg_rca8_and_4_6_a_4 & f_u_wallace_pg_rca8_and_4_6_b_6;
  assign f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_fa15_y4 = f_u_wallace_pg_rca8_fa15_y4;
  assign f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_and_5_5_y0 = f_u_wallace_pg_rca8_and_5_5_y0;
  assign f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_and_4_6_y0 = f_u_wallace_pg_rca8_and_4_6_y0;
  assign f_u_wallace_pg_rca8_fa16_y0 = f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_fa15_y4 ^ f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_and_5_5_y0;
  assign f_u_wallace_pg_rca8_fa16_y1 = f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_fa15_y4 & f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_and_5_5_y0;
  assign f_u_wallace_pg_rca8_fa16_y2 = f_u_wallace_pg_rca8_fa16_y0 ^ f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_and_4_6_y0;
  assign f_u_wallace_pg_rca8_fa16_y3 = f_u_wallace_pg_rca8_fa16_y0 & f_u_wallace_pg_rca8_fa16_f_u_wallace_pg_rca8_and_4_6_y0;
  assign f_u_wallace_pg_rca8_fa16_y4 = f_u_wallace_pg_rca8_fa16_y1 | f_u_wallace_pg_rca8_fa16_y3;
  assign f_u_wallace_pg_rca8_and_5_6_a_5 = a_5;
  assign f_u_wallace_pg_rca8_and_5_6_b_6 = b_6;
  assign f_u_wallace_pg_rca8_and_5_6_y0 = f_u_wallace_pg_rca8_and_5_6_a_5 & f_u_wallace_pg_rca8_and_5_6_b_6;
  assign f_u_wallace_pg_rca8_and_4_7_a_4 = a_4;
  assign f_u_wallace_pg_rca8_and_4_7_b_7 = b_7;
  assign f_u_wallace_pg_rca8_and_4_7_y0 = f_u_wallace_pg_rca8_and_4_7_a_4 & f_u_wallace_pg_rca8_and_4_7_b_7;
  assign f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_fa16_y4 = f_u_wallace_pg_rca8_fa16_y4;
  assign f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_and_5_6_y0 = f_u_wallace_pg_rca8_and_5_6_y0;
  assign f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_and_4_7_y0 = f_u_wallace_pg_rca8_and_4_7_y0;
  assign f_u_wallace_pg_rca8_fa17_y0 = f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_fa16_y4 ^ f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_and_5_6_y0;
  assign f_u_wallace_pg_rca8_fa17_y1 = f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_fa16_y4 & f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_and_5_6_y0;
  assign f_u_wallace_pg_rca8_fa17_y2 = f_u_wallace_pg_rca8_fa17_y0 ^ f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_and_4_7_y0;
  assign f_u_wallace_pg_rca8_fa17_y3 = f_u_wallace_pg_rca8_fa17_y0 & f_u_wallace_pg_rca8_fa17_f_u_wallace_pg_rca8_and_4_7_y0;
  assign f_u_wallace_pg_rca8_fa17_y4 = f_u_wallace_pg_rca8_fa17_y1 | f_u_wallace_pg_rca8_fa17_y3;
  assign f_u_wallace_pg_rca8_and_0_4_a_0 = a_0;
  assign f_u_wallace_pg_rca8_and_0_4_b_4 = b_4;
  assign f_u_wallace_pg_rca8_and_0_4_y0 = f_u_wallace_pg_rca8_and_0_4_a_0 & f_u_wallace_pg_rca8_and_0_4_b_4;
  assign f_u_wallace_pg_rca8_ha2_f_u_wallace_pg_rca8_and_0_4_y0 = f_u_wallace_pg_rca8_and_0_4_y0;
  assign f_u_wallace_pg_rca8_ha2_f_u_wallace_pg_rca8_fa1_y2 = f_u_wallace_pg_rca8_fa1_y2;
  assign f_u_wallace_pg_rca8_ha2_y0 = f_u_wallace_pg_rca8_ha2_f_u_wallace_pg_rca8_and_0_4_y0 ^ f_u_wallace_pg_rca8_ha2_f_u_wallace_pg_rca8_fa1_y2;
  assign f_u_wallace_pg_rca8_ha2_y1 = f_u_wallace_pg_rca8_ha2_f_u_wallace_pg_rca8_and_0_4_y0 & f_u_wallace_pg_rca8_ha2_f_u_wallace_pg_rca8_fa1_y2;
  assign f_u_wallace_pg_rca8_and_1_4_a_1 = a_1;
  assign f_u_wallace_pg_rca8_and_1_4_b_4 = b_4;
  assign f_u_wallace_pg_rca8_and_1_4_y0 = f_u_wallace_pg_rca8_and_1_4_a_1 & f_u_wallace_pg_rca8_and_1_4_b_4;
  assign f_u_wallace_pg_rca8_and_0_5_a_0 = a_0;
  assign f_u_wallace_pg_rca8_and_0_5_b_5 = b_5;
  assign f_u_wallace_pg_rca8_and_0_5_y0 = f_u_wallace_pg_rca8_and_0_5_a_0 & f_u_wallace_pg_rca8_and_0_5_b_5;
  assign f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_ha2_y1 = f_u_wallace_pg_rca8_ha2_y1;
  assign f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_and_1_4_y0 = f_u_wallace_pg_rca8_and_1_4_y0;
  assign f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_and_0_5_y0 = f_u_wallace_pg_rca8_and_0_5_y0;
  assign f_u_wallace_pg_rca8_fa18_y0 = f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_ha2_y1 ^ f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_and_1_4_y0;
  assign f_u_wallace_pg_rca8_fa18_y1 = f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_ha2_y1 & f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_and_1_4_y0;
  assign f_u_wallace_pg_rca8_fa18_y2 = f_u_wallace_pg_rca8_fa18_y0 ^ f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_and_0_5_y0;
  assign f_u_wallace_pg_rca8_fa18_y3 = f_u_wallace_pg_rca8_fa18_y0 & f_u_wallace_pg_rca8_fa18_f_u_wallace_pg_rca8_and_0_5_y0;
  assign f_u_wallace_pg_rca8_fa18_y4 = f_u_wallace_pg_rca8_fa18_y1 | f_u_wallace_pg_rca8_fa18_y3;
  assign f_u_wallace_pg_rca8_and_2_4_a_2 = a_2;
  assign f_u_wallace_pg_rca8_and_2_4_b_4 = b_4;
  assign f_u_wallace_pg_rca8_and_2_4_y0 = f_u_wallace_pg_rca8_and_2_4_a_2 & f_u_wallace_pg_rca8_and_2_4_b_4;
  assign f_u_wallace_pg_rca8_and_1_5_a_1 = a_1;
  assign f_u_wallace_pg_rca8_and_1_5_b_5 = b_5;
  assign f_u_wallace_pg_rca8_and_1_5_y0 = f_u_wallace_pg_rca8_and_1_5_a_1 & f_u_wallace_pg_rca8_and_1_5_b_5;
  assign f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_fa18_y4 = f_u_wallace_pg_rca8_fa18_y4;
  assign f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_and_2_4_y0 = f_u_wallace_pg_rca8_and_2_4_y0;
  assign f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_and_1_5_y0 = f_u_wallace_pg_rca8_and_1_5_y0;
  assign f_u_wallace_pg_rca8_fa19_y0 = f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_fa18_y4 ^ f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_and_2_4_y0;
  assign f_u_wallace_pg_rca8_fa19_y1 = f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_fa18_y4 & f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_and_2_4_y0;
  assign f_u_wallace_pg_rca8_fa19_y2 = f_u_wallace_pg_rca8_fa19_y0 ^ f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_and_1_5_y0;
  assign f_u_wallace_pg_rca8_fa19_y3 = f_u_wallace_pg_rca8_fa19_y0 & f_u_wallace_pg_rca8_fa19_f_u_wallace_pg_rca8_and_1_5_y0;
  assign f_u_wallace_pg_rca8_fa19_y4 = f_u_wallace_pg_rca8_fa19_y1 | f_u_wallace_pg_rca8_fa19_y3;
  assign f_u_wallace_pg_rca8_and_3_4_a_3 = a_3;
  assign f_u_wallace_pg_rca8_and_3_4_b_4 = b_4;
  assign f_u_wallace_pg_rca8_and_3_4_y0 = f_u_wallace_pg_rca8_and_3_4_a_3 & f_u_wallace_pg_rca8_and_3_4_b_4;
  assign f_u_wallace_pg_rca8_and_2_5_a_2 = a_2;
  assign f_u_wallace_pg_rca8_and_2_5_b_5 = b_5;
  assign f_u_wallace_pg_rca8_and_2_5_y0 = f_u_wallace_pg_rca8_and_2_5_a_2 & f_u_wallace_pg_rca8_and_2_5_b_5;
  assign f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_fa19_y4 = f_u_wallace_pg_rca8_fa19_y4;
  assign f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_and_3_4_y0 = f_u_wallace_pg_rca8_and_3_4_y0;
  assign f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_and_2_5_y0 = f_u_wallace_pg_rca8_and_2_5_y0;
  assign f_u_wallace_pg_rca8_fa20_y0 = f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_fa19_y4 ^ f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_and_3_4_y0;
  assign f_u_wallace_pg_rca8_fa20_y1 = f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_fa19_y4 & f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_and_3_4_y0;
  assign f_u_wallace_pg_rca8_fa20_y2 = f_u_wallace_pg_rca8_fa20_y0 ^ f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_and_2_5_y0;
  assign f_u_wallace_pg_rca8_fa20_y3 = f_u_wallace_pg_rca8_fa20_y0 & f_u_wallace_pg_rca8_fa20_f_u_wallace_pg_rca8_and_2_5_y0;
  assign f_u_wallace_pg_rca8_fa20_y4 = f_u_wallace_pg_rca8_fa20_y1 | f_u_wallace_pg_rca8_fa20_y3;
  assign f_u_wallace_pg_rca8_and_3_5_a_3 = a_3;
  assign f_u_wallace_pg_rca8_and_3_5_b_5 = b_5;
  assign f_u_wallace_pg_rca8_and_3_5_y0 = f_u_wallace_pg_rca8_and_3_5_a_3 & f_u_wallace_pg_rca8_and_3_5_b_5;
  assign f_u_wallace_pg_rca8_and_2_6_a_2 = a_2;
  assign f_u_wallace_pg_rca8_and_2_6_b_6 = b_6;
  assign f_u_wallace_pg_rca8_and_2_6_y0 = f_u_wallace_pg_rca8_and_2_6_a_2 & f_u_wallace_pg_rca8_and_2_6_b_6;
  assign f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_fa20_y4 = f_u_wallace_pg_rca8_fa20_y4;
  assign f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_and_3_5_y0 = f_u_wallace_pg_rca8_and_3_5_y0;
  assign f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_and_2_6_y0 = f_u_wallace_pg_rca8_and_2_6_y0;
  assign f_u_wallace_pg_rca8_fa21_y0 = f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_fa20_y4 ^ f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_and_3_5_y0;
  assign f_u_wallace_pg_rca8_fa21_y1 = f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_fa20_y4 & f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_and_3_5_y0;
  assign f_u_wallace_pg_rca8_fa21_y2 = f_u_wallace_pg_rca8_fa21_y0 ^ f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_and_2_6_y0;
  assign f_u_wallace_pg_rca8_fa21_y3 = f_u_wallace_pg_rca8_fa21_y0 & f_u_wallace_pg_rca8_fa21_f_u_wallace_pg_rca8_and_2_6_y0;
  assign f_u_wallace_pg_rca8_fa21_y4 = f_u_wallace_pg_rca8_fa21_y1 | f_u_wallace_pg_rca8_fa21_y3;
  assign f_u_wallace_pg_rca8_and_3_6_a_3 = a_3;
  assign f_u_wallace_pg_rca8_and_3_6_b_6 = b_6;
  assign f_u_wallace_pg_rca8_and_3_6_y0 = f_u_wallace_pg_rca8_and_3_6_a_3 & f_u_wallace_pg_rca8_and_3_6_b_6;
  assign f_u_wallace_pg_rca8_and_2_7_a_2 = a_2;
  assign f_u_wallace_pg_rca8_and_2_7_b_7 = b_7;
  assign f_u_wallace_pg_rca8_and_2_7_y0 = f_u_wallace_pg_rca8_and_2_7_a_2 & f_u_wallace_pg_rca8_and_2_7_b_7;
  assign f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_fa21_y4 = f_u_wallace_pg_rca8_fa21_y4;
  assign f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_and_3_6_y0 = f_u_wallace_pg_rca8_and_3_6_y0;
  assign f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_and_2_7_y0 = f_u_wallace_pg_rca8_and_2_7_y0;
  assign f_u_wallace_pg_rca8_fa22_y0 = f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_fa21_y4 ^ f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_and_3_6_y0;
  assign f_u_wallace_pg_rca8_fa22_y1 = f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_fa21_y4 & f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_and_3_6_y0;
  assign f_u_wallace_pg_rca8_fa22_y2 = f_u_wallace_pg_rca8_fa22_y0 ^ f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_and_2_7_y0;
  assign f_u_wallace_pg_rca8_fa22_y3 = f_u_wallace_pg_rca8_fa22_y0 & f_u_wallace_pg_rca8_fa22_f_u_wallace_pg_rca8_and_2_7_y0;
  assign f_u_wallace_pg_rca8_fa22_y4 = f_u_wallace_pg_rca8_fa22_y1 | f_u_wallace_pg_rca8_fa22_y3;
  assign f_u_wallace_pg_rca8_and_3_7_a_3 = a_3;
  assign f_u_wallace_pg_rca8_and_3_7_b_7 = b_7;
  assign f_u_wallace_pg_rca8_and_3_7_y0 = f_u_wallace_pg_rca8_and_3_7_a_3 & f_u_wallace_pg_rca8_and_3_7_b_7;
  assign f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_fa22_y4 = f_u_wallace_pg_rca8_fa22_y4;
  assign f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_and_3_7_y0 = f_u_wallace_pg_rca8_and_3_7_y0;
  assign f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_fa7_y2 = f_u_wallace_pg_rca8_fa7_y2;
  assign f_u_wallace_pg_rca8_fa23_y0 = f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_fa22_y4 ^ f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_and_3_7_y0;
  assign f_u_wallace_pg_rca8_fa23_y1 = f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_fa22_y4 & f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_and_3_7_y0;
  assign f_u_wallace_pg_rca8_fa23_y2 = f_u_wallace_pg_rca8_fa23_y0 ^ f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_fa7_y2;
  assign f_u_wallace_pg_rca8_fa23_y3 = f_u_wallace_pg_rca8_fa23_y0 & f_u_wallace_pg_rca8_fa23_f_u_wallace_pg_rca8_fa7_y2;
  assign f_u_wallace_pg_rca8_fa23_y4 = f_u_wallace_pg_rca8_fa23_y1 | f_u_wallace_pg_rca8_fa23_y3;
  assign f_u_wallace_pg_rca8_ha3_f_u_wallace_pg_rca8_fa2_y2 = f_u_wallace_pg_rca8_fa2_y2;
  assign f_u_wallace_pg_rca8_ha3_f_u_wallace_pg_rca8_fa11_y2 = f_u_wallace_pg_rca8_fa11_y2;
  assign f_u_wallace_pg_rca8_ha3_y0 = f_u_wallace_pg_rca8_ha3_f_u_wallace_pg_rca8_fa2_y2 ^ f_u_wallace_pg_rca8_ha3_f_u_wallace_pg_rca8_fa11_y2;
  assign f_u_wallace_pg_rca8_ha3_y1 = f_u_wallace_pg_rca8_ha3_f_u_wallace_pg_rca8_fa2_y2 & f_u_wallace_pg_rca8_ha3_f_u_wallace_pg_rca8_fa11_y2;
  assign f_u_wallace_pg_rca8_and_0_6_a_0 = a_0;
  assign f_u_wallace_pg_rca8_and_0_6_b_6 = b_6;
  assign f_u_wallace_pg_rca8_and_0_6_y0 = f_u_wallace_pg_rca8_and_0_6_a_0 & f_u_wallace_pg_rca8_and_0_6_b_6;
  assign f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_ha3_y1 = f_u_wallace_pg_rca8_ha3_y1;
  assign f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_and_0_6_y0 = f_u_wallace_pg_rca8_and_0_6_y0;
  assign f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_fa3_y2 = f_u_wallace_pg_rca8_fa3_y2;
  assign f_u_wallace_pg_rca8_fa24_y0 = f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_ha3_y1 ^ f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_and_0_6_y0;
  assign f_u_wallace_pg_rca8_fa24_y1 = f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_ha3_y1 & f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_and_0_6_y0;
  assign f_u_wallace_pg_rca8_fa24_y2 = f_u_wallace_pg_rca8_fa24_y0 ^ f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_fa3_y2;
  assign f_u_wallace_pg_rca8_fa24_y3 = f_u_wallace_pg_rca8_fa24_y0 & f_u_wallace_pg_rca8_fa24_f_u_wallace_pg_rca8_fa3_y2;
  assign f_u_wallace_pg_rca8_fa24_y4 = f_u_wallace_pg_rca8_fa24_y1 | f_u_wallace_pg_rca8_fa24_y3;
  assign f_u_wallace_pg_rca8_and_1_6_a_1 = a_1;
  assign f_u_wallace_pg_rca8_and_1_6_b_6 = b_6;
  assign f_u_wallace_pg_rca8_and_1_6_y0 = f_u_wallace_pg_rca8_and_1_6_a_1 & f_u_wallace_pg_rca8_and_1_6_b_6;
  assign f_u_wallace_pg_rca8_and_0_7_a_0 = a_0;
  assign f_u_wallace_pg_rca8_and_0_7_b_7 = b_7;
  assign f_u_wallace_pg_rca8_and_0_7_y0 = f_u_wallace_pg_rca8_and_0_7_a_0 & f_u_wallace_pg_rca8_and_0_7_b_7;
  assign f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_fa24_y4 = f_u_wallace_pg_rca8_fa24_y4;
  assign f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_and_1_6_y0 = f_u_wallace_pg_rca8_and_1_6_y0;
  assign f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_and_0_7_y0 = f_u_wallace_pg_rca8_and_0_7_y0;
  assign f_u_wallace_pg_rca8_fa25_y0 = f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_fa24_y4 ^ f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_and_1_6_y0;
  assign f_u_wallace_pg_rca8_fa25_y1 = f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_fa24_y4 & f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_and_1_6_y0;
  assign f_u_wallace_pg_rca8_fa25_y2 = f_u_wallace_pg_rca8_fa25_y0 ^ f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_and_0_7_y0;
  assign f_u_wallace_pg_rca8_fa25_y3 = f_u_wallace_pg_rca8_fa25_y0 & f_u_wallace_pg_rca8_fa25_f_u_wallace_pg_rca8_and_0_7_y0;
  assign f_u_wallace_pg_rca8_fa25_y4 = f_u_wallace_pg_rca8_fa25_y1 | f_u_wallace_pg_rca8_fa25_y3;
  assign f_u_wallace_pg_rca8_and_1_7_a_1 = a_1;
  assign f_u_wallace_pg_rca8_and_1_7_b_7 = b_7;
  assign f_u_wallace_pg_rca8_and_1_7_y0 = f_u_wallace_pg_rca8_and_1_7_a_1 & f_u_wallace_pg_rca8_and_1_7_b_7;
  assign f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_fa25_y4 = f_u_wallace_pg_rca8_fa25_y4;
  assign f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_and_1_7_y0 = f_u_wallace_pg_rca8_and_1_7_y0;
  assign f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_fa5_y2 = f_u_wallace_pg_rca8_fa5_y2;
  assign f_u_wallace_pg_rca8_fa26_y0 = f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_fa25_y4 ^ f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_and_1_7_y0;
  assign f_u_wallace_pg_rca8_fa26_y1 = f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_fa25_y4 & f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_and_1_7_y0;
  assign f_u_wallace_pg_rca8_fa26_y2 = f_u_wallace_pg_rca8_fa26_y0 ^ f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_fa5_y2;
  assign f_u_wallace_pg_rca8_fa26_y3 = f_u_wallace_pg_rca8_fa26_y0 & f_u_wallace_pg_rca8_fa26_f_u_wallace_pg_rca8_fa5_y2;
  assign f_u_wallace_pg_rca8_fa26_y4 = f_u_wallace_pg_rca8_fa26_y1 | f_u_wallace_pg_rca8_fa26_y3;
  assign f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa26_y4 = f_u_wallace_pg_rca8_fa26_y4;
  assign f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa6_y2 = f_u_wallace_pg_rca8_fa6_y2;
  assign f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa15_y2 = f_u_wallace_pg_rca8_fa15_y2;
  assign f_u_wallace_pg_rca8_fa27_y0 = f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa26_y4 ^ f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa6_y2;
  assign f_u_wallace_pg_rca8_fa27_y1 = f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa26_y4 & f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa6_y2;
  assign f_u_wallace_pg_rca8_fa27_y2 = f_u_wallace_pg_rca8_fa27_y0 ^ f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa15_y2;
  assign f_u_wallace_pg_rca8_fa27_y3 = f_u_wallace_pg_rca8_fa27_y0 & f_u_wallace_pg_rca8_fa27_f_u_wallace_pg_rca8_fa15_y2;
  assign f_u_wallace_pg_rca8_fa27_y4 = f_u_wallace_pg_rca8_fa27_y1 | f_u_wallace_pg_rca8_fa27_y3;
  assign f_u_wallace_pg_rca8_ha4_f_u_wallace_pg_rca8_fa12_y2 = f_u_wallace_pg_rca8_fa12_y2;
  assign f_u_wallace_pg_rca8_ha4_f_u_wallace_pg_rca8_fa19_y2 = f_u_wallace_pg_rca8_fa19_y2;
  assign f_u_wallace_pg_rca8_ha4_y0 = f_u_wallace_pg_rca8_ha4_f_u_wallace_pg_rca8_fa12_y2 ^ f_u_wallace_pg_rca8_ha4_f_u_wallace_pg_rca8_fa19_y2;
  assign f_u_wallace_pg_rca8_ha4_y1 = f_u_wallace_pg_rca8_ha4_f_u_wallace_pg_rca8_fa12_y2 & f_u_wallace_pg_rca8_ha4_f_u_wallace_pg_rca8_fa19_y2;
  assign f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_ha4_y1 = f_u_wallace_pg_rca8_ha4_y1;
  assign f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_fa4_y2 = f_u_wallace_pg_rca8_fa4_y2;
  assign f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_fa13_y2 = f_u_wallace_pg_rca8_fa13_y2;
  assign f_u_wallace_pg_rca8_fa28_y0 = f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_ha4_y1 ^ f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_fa4_y2;
  assign f_u_wallace_pg_rca8_fa28_y1 = f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_ha4_y1 & f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_fa4_y2;
  assign f_u_wallace_pg_rca8_fa28_y2 = f_u_wallace_pg_rca8_fa28_y0 ^ f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_fa13_y2;
  assign f_u_wallace_pg_rca8_fa28_y3 = f_u_wallace_pg_rca8_fa28_y0 & f_u_wallace_pg_rca8_fa28_f_u_wallace_pg_rca8_fa13_y2;
  assign f_u_wallace_pg_rca8_fa28_y4 = f_u_wallace_pg_rca8_fa28_y1 | f_u_wallace_pg_rca8_fa28_y3;
  assign f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa28_y4 = f_u_wallace_pg_rca8_fa28_y4;
  assign f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa14_y2 = f_u_wallace_pg_rca8_fa14_y2;
  assign f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa21_y2 = f_u_wallace_pg_rca8_fa21_y2;
  assign f_u_wallace_pg_rca8_fa29_y0 = f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa28_y4 ^ f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa14_y2;
  assign f_u_wallace_pg_rca8_fa29_y1 = f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa28_y4 & f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa14_y2;
  assign f_u_wallace_pg_rca8_fa29_y2 = f_u_wallace_pg_rca8_fa29_y0 ^ f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa21_y2;
  assign f_u_wallace_pg_rca8_fa29_y3 = f_u_wallace_pg_rca8_fa29_y0 & f_u_wallace_pg_rca8_fa29_f_u_wallace_pg_rca8_fa21_y2;
  assign f_u_wallace_pg_rca8_fa29_y4 = f_u_wallace_pg_rca8_fa29_y1 | f_u_wallace_pg_rca8_fa29_y3;
  assign f_u_wallace_pg_rca8_ha5_f_u_wallace_pg_rca8_fa20_y2 = f_u_wallace_pg_rca8_fa20_y2;
  assign f_u_wallace_pg_rca8_ha5_f_u_wallace_pg_rca8_fa25_y2 = f_u_wallace_pg_rca8_fa25_y2;
  assign f_u_wallace_pg_rca8_ha5_y0 = f_u_wallace_pg_rca8_ha5_f_u_wallace_pg_rca8_fa20_y2 ^ f_u_wallace_pg_rca8_ha5_f_u_wallace_pg_rca8_fa25_y2;
  assign f_u_wallace_pg_rca8_ha5_y1 = f_u_wallace_pg_rca8_ha5_f_u_wallace_pg_rca8_fa20_y2 & f_u_wallace_pg_rca8_ha5_f_u_wallace_pg_rca8_fa25_y2;
  assign f_u_wallace_pg_rca8_ha6_f_u_wallace_pg_rca8_ha5_y1 = f_u_wallace_pg_rca8_ha5_y1;
  assign f_u_wallace_pg_rca8_ha6_f_u_wallace_pg_rca8_fa26_y2 = f_u_wallace_pg_rca8_fa26_y2;
  assign f_u_wallace_pg_rca8_ha6_y0 = f_u_wallace_pg_rca8_ha6_f_u_wallace_pg_rca8_ha5_y1 ^ f_u_wallace_pg_rca8_ha6_f_u_wallace_pg_rca8_fa26_y2;
  assign f_u_wallace_pg_rca8_ha6_y1 = f_u_wallace_pg_rca8_ha6_f_u_wallace_pg_rca8_ha5_y1 & f_u_wallace_pg_rca8_ha6_f_u_wallace_pg_rca8_fa26_y2;
  assign f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_ha6_y1 = f_u_wallace_pg_rca8_ha6_y1;
  assign f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_fa29_y4 = f_u_wallace_pg_rca8_fa29_y4;
  assign f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_fa22_y2 = f_u_wallace_pg_rca8_fa22_y2;
  assign f_u_wallace_pg_rca8_fa30_y0 = f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_ha6_y1 ^ f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_fa29_y4;
  assign f_u_wallace_pg_rca8_fa30_y1 = f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_ha6_y1 & f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_fa29_y4;
  assign f_u_wallace_pg_rca8_fa30_y2 = f_u_wallace_pg_rca8_fa30_y0 ^ f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_fa22_y2;
  assign f_u_wallace_pg_rca8_fa30_y3 = f_u_wallace_pg_rca8_fa30_y0 & f_u_wallace_pg_rca8_fa30_f_u_wallace_pg_rca8_fa22_y2;
  assign f_u_wallace_pg_rca8_fa30_y4 = f_u_wallace_pg_rca8_fa30_y1 | f_u_wallace_pg_rca8_fa30_y3;
  assign f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa30_y4 = f_u_wallace_pg_rca8_fa30_y4;
  assign f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa27_y4 = f_u_wallace_pg_rca8_fa27_y4;
  assign f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa16_y2 = f_u_wallace_pg_rca8_fa16_y2;
  assign f_u_wallace_pg_rca8_fa31_y0 = f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa30_y4 ^ f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa27_y4;
  assign f_u_wallace_pg_rca8_fa31_y1 = f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa30_y4 & f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa27_y4;
  assign f_u_wallace_pg_rca8_fa31_y2 = f_u_wallace_pg_rca8_fa31_y0 ^ f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa16_y2;
  assign f_u_wallace_pg_rca8_fa31_y3 = f_u_wallace_pg_rca8_fa31_y0 & f_u_wallace_pg_rca8_fa31_f_u_wallace_pg_rca8_fa16_y2;
  assign f_u_wallace_pg_rca8_fa31_y4 = f_u_wallace_pg_rca8_fa31_y1 | f_u_wallace_pg_rca8_fa31_y3;
  assign f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa31_y4 = f_u_wallace_pg_rca8_fa31_y4;
  assign f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa23_y4 = f_u_wallace_pg_rca8_fa23_y4;
  assign f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa8_y2 = f_u_wallace_pg_rca8_fa8_y2;
  assign f_u_wallace_pg_rca8_fa32_y0 = f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa31_y4 ^ f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa23_y4;
  assign f_u_wallace_pg_rca8_fa32_y1 = f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa31_y4 & f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa23_y4;
  assign f_u_wallace_pg_rca8_fa32_y2 = f_u_wallace_pg_rca8_fa32_y0 ^ f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa8_y2;
  assign f_u_wallace_pg_rca8_fa32_y3 = f_u_wallace_pg_rca8_fa32_y0 & f_u_wallace_pg_rca8_fa32_f_u_wallace_pg_rca8_fa8_y2;
  assign f_u_wallace_pg_rca8_fa32_y4 = f_u_wallace_pg_rca8_fa32_y1 | f_u_wallace_pg_rca8_fa32_y3;
  assign f_u_wallace_pg_rca8_and_5_7_a_5 = a_5;
  assign f_u_wallace_pg_rca8_and_5_7_b_7 = b_7;
  assign f_u_wallace_pg_rca8_and_5_7_y0 = f_u_wallace_pg_rca8_and_5_7_a_5 & f_u_wallace_pg_rca8_and_5_7_b_7;
  assign f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_fa32_y4 = f_u_wallace_pg_rca8_fa32_y4;
  assign f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_fa17_y4 = f_u_wallace_pg_rca8_fa17_y4;
  assign f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_and_5_7_y0 = f_u_wallace_pg_rca8_and_5_7_y0;
  assign f_u_wallace_pg_rca8_fa33_y0 = f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_fa32_y4 ^ f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_fa17_y4;
  assign f_u_wallace_pg_rca8_fa33_y1 = f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_fa32_y4 & f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_fa17_y4;
  assign f_u_wallace_pg_rca8_fa33_y2 = f_u_wallace_pg_rca8_fa33_y0 ^ f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_and_5_7_y0;
  assign f_u_wallace_pg_rca8_fa33_y3 = f_u_wallace_pg_rca8_fa33_y0 & f_u_wallace_pg_rca8_fa33_f_u_wallace_pg_rca8_and_5_7_y0;
  assign f_u_wallace_pg_rca8_fa33_y4 = f_u_wallace_pg_rca8_fa33_y1 | f_u_wallace_pg_rca8_fa33_y3;
  assign f_u_wallace_pg_rca8_and_7_6_a_7 = a_7;
  assign f_u_wallace_pg_rca8_and_7_6_b_6 = b_6;
  assign f_u_wallace_pg_rca8_and_7_6_y0 = f_u_wallace_pg_rca8_and_7_6_a_7 & f_u_wallace_pg_rca8_and_7_6_b_6;
  assign f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_fa33_y4 = f_u_wallace_pg_rca8_fa33_y4;
  assign f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_fa9_y4 = f_u_wallace_pg_rca8_fa9_y4;
  assign f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_and_7_6_y0 = f_u_wallace_pg_rca8_and_7_6_y0;
  assign f_u_wallace_pg_rca8_fa34_y0 = f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_fa33_y4 ^ f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_fa9_y4;
  assign f_u_wallace_pg_rca8_fa34_y1 = f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_fa33_y4 & f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_fa9_y4;
  assign f_u_wallace_pg_rca8_fa34_y2 = f_u_wallace_pg_rca8_fa34_y0 ^ f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_and_7_6_y0;
  assign f_u_wallace_pg_rca8_fa34_y3 = f_u_wallace_pg_rca8_fa34_y0 & f_u_wallace_pg_rca8_fa34_f_u_wallace_pg_rca8_and_7_6_y0;
  assign f_u_wallace_pg_rca8_fa34_y4 = f_u_wallace_pg_rca8_fa34_y1 | f_u_wallace_pg_rca8_fa34_y3;
  assign f_u_wallace_pg_rca8_and_0_0_a_0 = a_0;
  assign f_u_wallace_pg_rca8_and_0_0_b_0 = b_0;
  assign f_u_wallace_pg_rca8_and_0_0_y0 = f_u_wallace_pg_rca8_and_0_0_a_0 & f_u_wallace_pg_rca8_and_0_0_b_0;
  assign f_u_wallace_pg_rca8_and_1_0_a_1 = a_1;
  assign f_u_wallace_pg_rca8_and_1_0_b_0 = b_0;
  assign f_u_wallace_pg_rca8_and_1_0_y0 = f_u_wallace_pg_rca8_and_1_0_a_1 & f_u_wallace_pg_rca8_and_1_0_b_0;
  assign f_u_wallace_pg_rca8_and_0_2_a_0 = a_0;
  assign f_u_wallace_pg_rca8_and_0_2_b_2 = b_2;
  assign f_u_wallace_pg_rca8_and_0_2_y0 = f_u_wallace_pg_rca8_and_0_2_a_0 & f_u_wallace_pg_rca8_and_0_2_b_2;
  assign f_u_wallace_pg_rca8_and_6_7_a_6 = a_6;
  assign f_u_wallace_pg_rca8_and_6_7_b_7 = b_7;
  assign f_u_wallace_pg_rca8_and_6_7_y0 = f_u_wallace_pg_rca8_and_6_7_a_6 & f_u_wallace_pg_rca8_and_6_7_b_7;
  assign f_u_wallace_pg_rca8_and_0_1_a_0 = a_0;
  assign f_u_wallace_pg_rca8_and_0_1_b_1 = b_1;
  assign f_u_wallace_pg_rca8_and_0_1_y0 = f_u_wallace_pg_rca8_and_0_1_a_0 & f_u_wallace_pg_rca8_and_0_1_b_1;
  assign f_u_wallace_pg_rca8_and_7_7_a_7 = a_7;
  assign f_u_wallace_pg_rca8_and_7_7_b_7 = b_7;
  assign f_u_wallace_pg_rca8_and_7_7_y0 = f_u_wallace_pg_rca8_and_7_7_a_7 & f_u_wallace_pg_rca8_and_7_7_b_7;
  assign constant_wire_value_0_f_u_wallace_pg_rca8_and_1_0_y0 = f_u_wallace_pg_rca8_and_1_0_y0;
  assign constant_wire_value_0_f_u_wallace_pg_rca8_and_0_1_y0 = f_u_wallace_pg_rca8_and_0_1_y0;
  assign constant_wire_value_0_y0 = constant_wire_value_0_f_u_wallace_pg_rca8_and_1_0_y0 ^ constant_wire_value_0_f_u_wallace_pg_rca8_and_0_1_y0;
  assign constant_wire_value_0_y1 = ~(constant_wire_value_0_f_u_wallace_pg_rca8_and_1_0_y0 ^ constant_wire_value_0_f_u_wallace_pg_rca8_and_0_1_y0);
  assign constant_wire_0 = ~(constant_wire_value_0_y0 | constant_wire_value_0_y1);
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa0_f_u_wallace_pg_rca8_and_1_0_y0 = f_u_wallace_pg_rca8_and_1_0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa0_f_u_wallace_pg_rca8_and_0_1_y0 = f_u_wallace_pg_rca8_and_0_1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa0_constant_wire_0 = constant_wire_0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa0_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa0_f_u_wallace_pg_rca8_and_1_0_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa0_f_u_wallace_pg_rca8_and_0_1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa0_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa0_f_u_wallace_pg_rca8_and_1_0_y0 & f_u_wallace_pg_rca8_u_pg_rca14_fa0_f_u_wallace_pg_rca8_and_0_1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa0_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa0_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa0_constant_wire_0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and0_constant_wire_0 = constant_wire_0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and0_f_u_wallace_pg_rca8_u_pg_rca14_fa0_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and0_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and0_constant_wire_0 & f_u_wallace_pg_rca8_u_pg_rca14_and0_f_u_wallace_pg_rca8_u_pg_rca14_fa0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or0_f_u_wallace_pg_rca8_u_pg_rca14_and0_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or0_f_u_wallace_pg_rca8_u_pg_rca14_fa0_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa0_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or0_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or0_f_u_wallace_pg_rca8_u_pg_rca14_and0_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or0_f_u_wallace_pg_rca8_u_pg_rca14_fa0_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_and_0_2_y0 = f_u_wallace_pg_rca8_and_0_2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_ha0_y0 = f_u_wallace_pg_rca8_ha0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_u_pg_rca14_or0_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa1_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_and_0_2_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_ha0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa1_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_and_0_2_y0 & f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_ha0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa1_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa1_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa1_f_u_wallace_pg_rca8_u_pg_rca14_or0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and1_f_u_wallace_pg_rca8_u_pg_rca14_or0_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or0_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and1_f_u_wallace_pg_rca8_u_pg_rca14_fa1_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and1_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and1_f_u_wallace_pg_rca8_u_pg_rca14_or0_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and1_f_u_wallace_pg_rca8_u_pg_rca14_fa1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or1_f_u_wallace_pg_rca8_u_pg_rca14_and1_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or1_f_u_wallace_pg_rca8_u_pg_rca14_fa1_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa1_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or1_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or1_f_u_wallace_pg_rca8_u_pg_rca14_and1_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or1_f_u_wallace_pg_rca8_u_pg_rca14_fa1_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_fa0_y2 = f_u_wallace_pg_rca8_fa0_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_ha1_y0 = f_u_wallace_pg_rca8_ha1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_u_pg_rca14_or1_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa2_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_fa0_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_ha1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa2_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_fa0_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_ha1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa2_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa2_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa2_f_u_wallace_pg_rca8_u_pg_rca14_or1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and2_f_u_wallace_pg_rca8_u_pg_rca14_or1_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or1_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and2_f_u_wallace_pg_rca8_u_pg_rca14_fa2_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and2_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and2_f_u_wallace_pg_rca8_u_pg_rca14_or1_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and2_f_u_wallace_pg_rca8_u_pg_rca14_fa2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or2_f_u_wallace_pg_rca8_u_pg_rca14_and2_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or2_f_u_wallace_pg_rca8_u_pg_rca14_fa2_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa2_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or2_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or2_f_u_wallace_pg_rca8_u_pg_rca14_and2_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or2_f_u_wallace_pg_rca8_u_pg_rca14_fa2_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_fa10_y2 = f_u_wallace_pg_rca8_fa10_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_ha2_y0 = f_u_wallace_pg_rca8_ha2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_u_pg_rca14_or2_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa3_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_fa10_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_ha2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa3_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_fa10_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_ha2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa3_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa3_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa3_f_u_wallace_pg_rca8_u_pg_rca14_or2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and3_f_u_wallace_pg_rca8_u_pg_rca14_or2_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or2_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and3_f_u_wallace_pg_rca8_u_pg_rca14_fa3_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and3_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and3_f_u_wallace_pg_rca8_u_pg_rca14_or2_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and3_f_u_wallace_pg_rca8_u_pg_rca14_fa3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or3_f_u_wallace_pg_rca8_u_pg_rca14_and3_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or3_f_u_wallace_pg_rca8_u_pg_rca14_fa3_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa3_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or3_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or3_f_u_wallace_pg_rca8_u_pg_rca14_and3_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or3_f_u_wallace_pg_rca8_u_pg_rca14_fa3_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_fa18_y2 = f_u_wallace_pg_rca8_fa18_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_ha3_y0 = f_u_wallace_pg_rca8_ha3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_u_pg_rca14_or3_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa4_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_fa18_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_ha3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa4_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_fa18_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_ha3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa4_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa4_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa4_f_u_wallace_pg_rca8_u_pg_rca14_or3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and4_f_u_wallace_pg_rca8_u_pg_rca14_or3_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or3_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and4_f_u_wallace_pg_rca8_u_pg_rca14_fa4_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and4_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and4_f_u_wallace_pg_rca8_u_pg_rca14_or3_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and4_f_u_wallace_pg_rca8_u_pg_rca14_fa4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or4_f_u_wallace_pg_rca8_u_pg_rca14_and4_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or4_f_u_wallace_pg_rca8_u_pg_rca14_fa4_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa4_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or4_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or4_f_u_wallace_pg_rca8_u_pg_rca14_and4_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or4_f_u_wallace_pg_rca8_u_pg_rca14_fa4_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_fa24_y2 = f_u_wallace_pg_rca8_fa24_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_ha4_y0 = f_u_wallace_pg_rca8_ha4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_u_pg_rca14_or4_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa5_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_fa24_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_ha4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa5_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_fa24_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_ha4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa5_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa5_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa5_f_u_wallace_pg_rca8_u_pg_rca14_or4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and5_f_u_wallace_pg_rca8_u_pg_rca14_or4_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or4_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and5_f_u_wallace_pg_rca8_u_pg_rca14_fa5_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and5_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and5_f_u_wallace_pg_rca8_u_pg_rca14_or4_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and5_f_u_wallace_pg_rca8_u_pg_rca14_fa5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or5_f_u_wallace_pg_rca8_u_pg_rca14_and5_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or5_f_u_wallace_pg_rca8_u_pg_rca14_fa5_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa5_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or5_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or5_f_u_wallace_pg_rca8_u_pg_rca14_and5_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or5_f_u_wallace_pg_rca8_u_pg_rca14_fa5_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_fa28_y2 = f_u_wallace_pg_rca8_fa28_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_ha5_y0 = f_u_wallace_pg_rca8_ha5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_u_pg_rca14_or5_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa6_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_fa28_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_ha5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa6_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_fa28_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_ha5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa6_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa6_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa6_f_u_wallace_pg_rca8_u_pg_rca14_or5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and6_f_u_wallace_pg_rca8_u_pg_rca14_or5_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or5_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and6_f_u_wallace_pg_rca8_u_pg_rca14_fa6_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and6_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and6_f_u_wallace_pg_rca8_u_pg_rca14_or5_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and6_f_u_wallace_pg_rca8_u_pg_rca14_fa6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or6_f_u_wallace_pg_rca8_u_pg_rca14_and6_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or6_f_u_wallace_pg_rca8_u_pg_rca14_fa6_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa6_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or6_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or6_f_u_wallace_pg_rca8_u_pg_rca14_and6_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or6_f_u_wallace_pg_rca8_u_pg_rca14_fa6_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_fa29_y2 = f_u_wallace_pg_rca8_fa29_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_ha6_y0 = f_u_wallace_pg_rca8_ha6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_u_pg_rca14_or6_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa7_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_fa29_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_ha6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa7_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_fa29_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_ha6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa7_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa7_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa7_f_u_wallace_pg_rca8_u_pg_rca14_or6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and7_f_u_wallace_pg_rca8_u_pg_rca14_or6_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or6_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and7_f_u_wallace_pg_rca8_u_pg_rca14_fa7_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and7_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and7_f_u_wallace_pg_rca8_u_pg_rca14_or6_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and7_f_u_wallace_pg_rca8_u_pg_rca14_fa7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or7_f_u_wallace_pg_rca8_u_pg_rca14_and7_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or7_f_u_wallace_pg_rca8_u_pg_rca14_fa7_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa7_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or7_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or7_f_u_wallace_pg_rca8_u_pg_rca14_and7_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or7_f_u_wallace_pg_rca8_u_pg_rca14_fa7_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_fa27_y2 = f_u_wallace_pg_rca8_fa27_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_fa30_y2 = f_u_wallace_pg_rca8_fa30_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_u_pg_rca14_or7_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa8_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_fa27_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_fa30_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa8_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_fa27_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_fa30_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa8_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa8_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa8_f_u_wallace_pg_rca8_u_pg_rca14_or7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and8_f_u_wallace_pg_rca8_u_pg_rca14_or7_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and8_f_u_wallace_pg_rca8_u_pg_rca14_fa8_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa8_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and8_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and8_f_u_wallace_pg_rca8_u_pg_rca14_or7_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and8_f_u_wallace_pg_rca8_u_pg_rca14_fa8_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or8_f_u_wallace_pg_rca8_u_pg_rca14_and8_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and8_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or8_f_u_wallace_pg_rca8_u_pg_rca14_fa8_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa8_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or8_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or8_f_u_wallace_pg_rca8_u_pg_rca14_and8_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or8_f_u_wallace_pg_rca8_u_pg_rca14_fa8_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_fa23_y2 = f_u_wallace_pg_rca8_fa23_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_fa31_y2 = f_u_wallace_pg_rca8_fa31_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_u_pg_rca14_or8_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or8_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa9_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_fa23_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_fa31_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa9_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_fa23_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_fa31_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa9_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa9_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa9_f_u_wallace_pg_rca8_u_pg_rca14_or8_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and9_f_u_wallace_pg_rca8_u_pg_rca14_or8_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or8_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and9_f_u_wallace_pg_rca8_u_pg_rca14_fa9_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa9_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and9_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and9_f_u_wallace_pg_rca8_u_pg_rca14_or8_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and9_f_u_wallace_pg_rca8_u_pg_rca14_fa9_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or9_f_u_wallace_pg_rca8_u_pg_rca14_and9_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and9_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or9_f_u_wallace_pg_rca8_u_pg_rca14_fa9_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa9_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or9_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or9_f_u_wallace_pg_rca8_u_pg_rca14_and9_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or9_f_u_wallace_pg_rca8_u_pg_rca14_fa9_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_fa17_y2 = f_u_wallace_pg_rca8_fa17_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_fa32_y2 = f_u_wallace_pg_rca8_fa32_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_u_pg_rca14_or9_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or9_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa10_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_fa17_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_fa32_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa10_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_fa17_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_fa32_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa10_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa10_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa10_f_u_wallace_pg_rca8_u_pg_rca14_or9_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and10_f_u_wallace_pg_rca8_u_pg_rca14_or9_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or9_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and10_f_u_wallace_pg_rca8_u_pg_rca14_fa10_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa10_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and10_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and10_f_u_wallace_pg_rca8_u_pg_rca14_or9_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and10_f_u_wallace_pg_rca8_u_pg_rca14_fa10_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or10_f_u_wallace_pg_rca8_u_pg_rca14_and10_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and10_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or10_f_u_wallace_pg_rca8_u_pg_rca14_fa10_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa10_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or10_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or10_f_u_wallace_pg_rca8_u_pg_rca14_and10_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or10_f_u_wallace_pg_rca8_u_pg_rca14_fa10_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_fa9_y2 = f_u_wallace_pg_rca8_fa9_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_fa33_y2 = f_u_wallace_pg_rca8_fa33_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_u_pg_rca14_or10_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or10_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa11_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_fa9_y2 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_fa33_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa11_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_fa9_y2 & f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_fa33_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa11_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa11_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa11_f_u_wallace_pg_rca8_u_pg_rca14_or10_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and11_f_u_wallace_pg_rca8_u_pg_rca14_or10_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or10_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and11_f_u_wallace_pg_rca8_u_pg_rca14_fa11_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa11_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and11_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and11_f_u_wallace_pg_rca8_u_pg_rca14_or10_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and11_f_u_wallace_pg_rca8_u_pg_rca14_fa11_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or11_f_u_wallace_pg_rca8_u_pg_rca14_and11_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and11_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or11_f_u_wallace_pg_rca8_u_pg_rca14_fa11_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa11_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or11_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or11_f_u_wallace_pg_rca8_u_pg_rca14_and11_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or11_f_u_wallace_pg_rca8_u_pg_rca14_fa11_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_and_6_7_y0 = f_u_wallace_pg_rca8_and_6_7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_fa34_y2 = f_u_wallace_pg_rca8_fa34_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_u_pg_rca14_or11_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or11_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa12_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_and_6_7_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_fa34_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa12_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_and_6_7_y0 & f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_fa34_y2;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa12_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa12_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa12_f_u_wallace_pg_rca8_u_pg_rca14_or11_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and12_f_u_wallace_pg_rca8_u_pg_rca14_or11_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or11_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and12_f_u_wallace_pg_rca8_u_pg_rca14_fa12_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa12_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and12_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and12_f_u_wallace_pg_rca8_u_pg_rca14_or11_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and12_f_u_wallace_pg_rca8_u_pg_rca14_fa12_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or12_f_u_wallace_pg_rca8_u_pg_rca14_and12_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and12_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or12_f_u_wallace_pg_rca8_u_pg_rca14_fa12_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa12_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or12_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or12_f_u_wallace_pg_rca8_u_pg_rca14_and12_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or12_f_u_wallace_pg_rca8_u_pg_rca14_fa12_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_fa34_y4 = f_u_wallace_pg_rca8_fa34_y4;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_and_7_7_y0 = f_u_wallace_pg_rca8_and_7_7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_u_pg_rca14_or12_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or12_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa13_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_fa34_y4 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_and_7_7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa13_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_fa34_y4 & f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_and_7_7_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_fa13_y2 = f_u_wallace_pg_rca8_u_pg_rca14_fa13_y0 ^ f_u_wallace_pg_rca8_u_pg_rca14_fa13_f_u_wallace_pg_rca8_u_pg_rca14_or12_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and13_f_u_wallace_pg_rca8_u_pg_rca14_or12_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or12_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and13_f_u_wallace_pg_rca8_u_pg_rca14_fa13_y0 = f_u_wallace_pg_rca8_u_pg_rca14_fa13_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_and13_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and13_f_u_wallace_pg_rca8_u_pg_rca14_or12_y0 & f_u_wallace_pg_rca8_u_pg_rca14_and13_f_u_wallace_pg_rca8_u_pg_rca14_fa13_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or13_f_u_wallace_pg_rca8_u_pg_rca14_and13_y0 = f_u_wallace_pg_rca8_u_pg_rca14_and13_y0;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or13_f_u_wallace_pg_rca8_u_pg_rca14_fa13_y1 = f_u_wallace_pg_rca8_u_pg_rca14_fa13_y1;
  assign f_u_wallace_pg_rca8_u_pg_rca14_or13_y0 = f_u_wallace_pg_rca8_u_pg_rca14_or13_f_u_wallace_pg_rca8_u_pg_rca14_and13_y0 | f_u_wallace_pg_rca8_u_pg_rca14_or13_f_u_wallace_pg_rca8_u_pg_rca14_fa13_y1;

  assign out[0] = f_u_wallace_pg_rca8_and_0_0_y0;
  assign out[1] = f_u_wallace_pg_rca8_u_pg_rca14_fa0_y2;
  assign out[2] = f_u_wallace_pg_rca8_u_pg_rca14_fa1_y2;
  assign out[3] = f_u_wallace_pg_rca8_u_pg_rca14_fa2_y2;
  assign out[4] = f_u_wallace_pg_rca8_u_pg_rca14_fa3_y2;
  assign out[5] = f_u_wallace_pg_rca8_u_pg_rca14_fa4_y2;
  assign out[6] = f_u_wallace_pg_rca8_u_pg_rca14_fa5_y2;
  assign out[7] = f_u_wallace_pg_rca8_u_pg_rca14_fa6_y2;
  assign out[8] = f_u_wallace_pg_rca8_u_pg_rca14_fa7_y2;
  assign out[9] = f_u_wallace_pg_rca8_u_pg_rca14_fa8_y2;
  assign out[10] = f_u_wallace_pg_rca8_u_pg_rca14_fa9_y2;
  assign out[11] = f_u_wallace_pg_rca8_u_pg_rca14_fa10_y2;
  assign out[12] = f_u_wallace_pg_rca8_u_pg_rca14_fa11_y2;
  assign out[13] = f_u_wallace_pg_rca8_u_pg_rca14_fa12_y2;
  assign out[14] = f_u_wallace_pg_rca8_u_pg_rca14_fa13_y2;
  assign out[15] = f_u_wallace_pg_rca8_u_pg_rca14_or13_y0;
endmodule