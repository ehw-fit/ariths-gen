module f_s_wallace_cla8(input [7:0] a, input [7:0] b, output [15:0] f_s_wallace_cla8_out);
  wire f_s_wallace_cla8_and_2_0;
  wire f_s_wallace_cla8_and_1_1;
  wire f_s_wallace_cla8_ha0_xor0;
  wire f_s_wallace_cla8_ha0_and0;
  wire f_s_wallace_cla8_and_3_0;
  wire f_s_wallace_cla8_and_2_1;
  wire f_s_wallace_cla8_fa0_xor0;
  wire f_s_wallace_cla8_fa0_and0;
  wire f_s_wallace_cla8_fa0_xor1;
  wire f_s_wallace_cla8_fa0_and1;
  wire f_s_wallace_cla8_fa0_or0;
  wire f_s_wallace_cla8_and_4_0;
  wire f_s_wallace_cla8_and_3_1;
  wire f_s_wallace_cla8_fa1_xor0;
  wire f_s_wallace_cla8_fa1_and0;
  wire f_s_wallace_cla8_fa1_xor1;
  wire f_s_wallace_cla8_fa1_and1;
  wire f_s_wallace_cla8_fa1_or0;
  wire f_s_wallace_cla8_and_5_0;
  wire f_s_wallace_cla8_and_4_1;
  wire f_s_wallace_cla8_fa2_xor0;
  wire f_s_wallace_cla8_fa2_and0;
  wire f_s_wallace_cla8_fa2_xor1;
  wire f_s_wallace_cla8_fa2_and1;
  wire f_s_wallace_cla8_fa2_or0;
  wire f_s_wallace_cla8_and_6_0;
  wire f_s_wallace_cla8_and_5_1;
  wire f_s_wallace_cla8_fa3_xor0;
  wire f_s_wallace_cla8_fa3_and0;
  wire f_s_wallace_cla8_fa3_xor1;
  wire f_s_wallace_cla8_fa3_and1;
  wire f_s_wallace_cla8_fa3_or0;
  wire f_s_wallace_cla8_nand_7_0;
  wire f_s_wallace_cla8_and_6_1;
  wire f_s_wallace_cla8_fa4_xor0;
  wire f_s_wallace_cla8_fa4_and0;
  wire f_s_wallace_cla8_fa4_xor1;
  wire f_s_wallace_cla8_fa4_and1;
  wire f_s_wallace_cla8_fa4_or0;
  wire f_s_wallace_cla8_nand_7_1;
  wire f_s_wallace_cla8_fa5_xor0;
  wire f_s_wallace_cla8_fa5_xor1;
  wire f_s_wallace_cla8_fa5_and1;
  wire f_s_wallace_cla8_fa5_or0;
  wire f_s_wallace_cla8_nand_7_2;
  wire f_s_wallace_cla8_and_6_3;
  wire f_s_wallace_cla8_fa6_xor0;
  wire f_s_wallace_cla8_fa6_and0;
  wire f_s_wallace_cla8_fa6_xor1;
  wire f_s_wallace_cla8_fa6_and1;
  wire f_s_wallace_cla8_fa6_or0;
  wire f_s_wallace_cla8_nand_7_3;
  wire f_s_wallace_cla8_and_6_4;
  wire f_s_wallace_cla8_fa7_xor0;
  wire f_s_wallace_cla8_fa7_and0;
  wire f_s_wallace_cla8_fa7_xor1;
  wire f_s_wallace_cla8_fa7_and1;
  wire f_s_wallace_cla8_fa7_or0;
  wire f_s_wallace_cla8_nand_7_4;
  wire f_s_wallace_cla8_and_6_5;
  wire f_s_wallace_cla8_fa8_xor0;
  wire f_s_wallace_cla8_fa8_and0;
  wire f_s_wallace_cla8_fa8_xor1;
  wire f_s_wallace_cla8_fa8_and1;
  wire f_s_wallace_cla8_fa8_or0;
  wire f_s_wallace_cla8_nand_7_5;
  wire f_s_wallace_cla8_and_6_6;
  wire f_s_wallace_cla8_fa9_xor0;
  wire f_s_wallace_cla8_fa9_and0;
  wire f_s_wallace_cla8_fa9_xor1;
  wire f_s_wallace_cla8_fa9_and1;
  wire f_s_wallace_cla8_fa9_or0;
  wire f_s_wallace_cla8_and_1_2;
  wire f_s_wallace_cla8_and_0_3;
  wire f_s_wallace_cla8_ha1_xor0;
  wire f_s_wallace_cla8_ha1_and0;
  wire f_s_wallace_cla8_and_2_2;
  wire f_s_wallace_cla8_and_1_3;
  wire f_s_wallace_cla8_fa10_xor0;
  wire f_s_wallace_cla8_fa10_and0;
  wire f_s_wallace_cla8_fa10_xor1;
  wire f_s_wallace_cla8_fa10_and1;
  wire f_s_wallace_cla8_fa10_or0;
  wire f_s_wallace_cla8_and_3_2;
  wire f_s_wallace_cla8_and_2_3;
  wire f_s_wallace_cla8_fa11_xor0;
  wire f_s_wallace_cla8_fa11_and0;
  wire f_s_wallace_cla8_fa11_xor1;
  wire f_s_wallace_cla8_fa11_and1;
  wire f_s_wallace_cla8_fa11_or0;
  wire f_s_wallace_cla8_and_4_2;
  wire f_s_wallace_cla8_and_3_3;
  wire f_s_wallace_cla8_fa12_xor0;
  wire f_s_wallace_cla8_fa12_and0;
  wire f_s_wallace_cla8_fa12_xor1;
  wire f_s_wallace_cla8_fa12_and1;
  wire f_s_wallace_cla8_fa12_or0;
  wire f_s_wallace_cla8_and_5_2;
  wire f_s_wallace_cla8_and_4_3;
  wire f_s_wallace_cla8_fa13_xor0;
  wire f_s_wallace_cla8_fa13_and0;
  wire f_s_wallace_cla8_fa13_xor1;
  wire f_s_wallace_cla8_fa13_and1;
  wire f_s_wallace_cla8_fa13_or0;
  wire f_s_wallace_cla8_and_6_2;
  wire f_s_wallace_cla8_and_5_3;
  wire f_s_wallace_cla8_fa14_xor0;
  wire f_s_wallace_cla8_fa14_and0;
  wire f_s_wallace_cla8_fa14_xor1;
  wire f_s_wallace_cla8_fa14_and1;
  wire f_s_wallace_cla8_fa14_or0;
  wire f_s_wallace_cla8_and_5_4;
  wire f_s_wallace_cla8_and_4_5;
  wire f_s_wallace_cla8_fa15_xor0;
  wire f_s_wallace_cla8_fa15_and0;
  wire f_s_wallace_cla8_fa15_xor1;
  wire f_s_wallace_cla8_fa15_and1;
  wire f_s_wallace_cla8_fa15_or0;
  wire f_s_wallace_cla8_and_5_5;
  wire f_s_wallace_cla8_and_4_6;
  wire f_s_wallace_cla8_fa16_xor0;
  wire f_s_wallace_cla8_fa16_and0;
  wire f_s_wallace_cla8_fa16_xor1;
  wire f_s_wallace_cla8_fa16_and1;
  wire f_s_wallace_cla8_fa16_or0;
  wire f_s_wallace_cla8_and_5_6;
  wire f_s_wallace_cla8_nand_4_7;
  wire f_s_wallace_cla8_fa17_xor0;
  wire f_s_wallace_cla8_fa17_and0;
  wire f_s_wallace_cla8_fa17_xor1;
  wire f_s_wallace_cla8_fa17_and1;
  wire f_s_wallace_cla8_fa17_or0;
  wire f_s_wallace_cla8_and_0_4;
  wire f_s_wallace_cla8_ha2_xor0;
  wire f_s_wallace_cla8_ha2_and0;
  wire f_s_wallace_cla8_and_1_4;
  wire f_s_wallace_cla8_and_0_5;
  wire f_s_wallace_cla8_fa18_xor0;
  wire f_s_wallace_cla8_fa18_and0;
  wire f_s_wallace_cla8_fa18_xor1;
  wire f_s_wallace_cla8_fa18_and1;
  wire f_s_wallace_cla8_fa18_or0;
  wire f_s_wallace_cla8_and_2_4;
  wire f_s_wallace_cla8_and_1_5;
  wire f_s_wallace_cla8_fa19_xor0;
  wire f_s_wallace_cla8_fa19_and0;
  wire f_s_wallace_cla8_fa19_xor1;
  wire f_s_wallace_cla8_fa19_and1;
  wire f_s_wallace_cla8_fa19_or0;
  wire f_s_wallace_cla8_and_3_4;
  wire f_s_wallace_cla8_and_2_5;
  wire f_s_wallace_cla8_fa20_xor0;
  wire f_s_wallace_cla8_fa20_and0;
  wire f_s_wallace_cla8_fa20_xor1;
  wire f_s_wallace_cla8_fa20_and1;
  wire f_s_wallace_cla8_fa20_or0;
  wire f_s_wallace_cla8_and_4_4;
  wire f_s_wallace_cla8_and_3_5;
  wire f_s_wallace_cla8_fa21_xor0;
  wire f_s_wallace_cla8_fa21_and0;
  wire f_s_wallace_cla8_fa21_xor1;
  wire f_s_wallace_cla8_fa21_and1;
  wire f_s_wallace_cla8_fa21_or0;
  wire f_s_wallace_cla8_and_3_6;
  wire f_s_wallace_cla8_nand_2_7;
  wire f_s_wallace_cla8_fa22_xor0;
  wire f_s_wallace_cla8_fa22_and0;
  wire f_s_wallace_cla8_fa22_xor1;
  wire f_s_wallace_cla8_fa22_and1;
  wire f_s_wallace_cla8_fa22_or0;
  wire f_s_wallace_cla8_nand_3_7;
  wire f_s_wallace_cla8_fa23_xor0;
  wire f_s_wallace_cla8_fa23_and0;
  wire f_s_wallace_cla8_fa23_xor1;
  wire f_s_wallace_cla8_fa23_and1;
  wire f_s_wallace_cla8_fa23_or0;
  wire f_s_wallace_cla8_ha3_xor0;
  wire f_s_wallace_cla8_ha3_and0;
  wire f_s_wallace_cla8_and_0_6;
  wire f_s_wallace_cla8_fa24_xor0;
  wire f_s_wallace_cla8_fa24_and0;
  wire f_s_wallace_cla8_fa24_xor1;
  wire f_s_wallace_cla8_fa24_and1;
  wire f_s_wallace_cla8_fa24_or0;
  wire f_s_wallace_cla8_and_1_6;
  wire f_s_wallace_cla8_nand_0_7;
  wire f_s_wallace_cla8_fa25_xor0;
  wire f_s_wallace_cla8_fa25_and0;
  wire f_s_wallace_cla8_fa25_xor1;
  wire f_s_wallace_cla8_fa25_and1;
  wire f_s_wallace_cla8_fa25_or0;
  wire f_s_wallace_cla8_and_2_6;
  wire f_s_wallace_cla8_nand_1_7;
  wire f_s_wallace_cla8_fa26_xor0;
  wire f_s_wallace_cla8_fa26_and0;
  wire f_s_wallace_cla8_fa26_xor1;
  wire f_s_wallace_cla8_fa26_and1;
  wire f_s_wallace_cla8_fa26_or0;
  wire f_s_wallace_cla8_fa27_xor0;
  wire f_s_wallace_cla8_fa27_and0;
  wire f_s_wallace_cla8_fa27_xor1;
  wire f_s_wallace_cla8_fa27_and1;
  wire f_s_wallace_cla8_fa27_or0;
  wire f_s_wallace_cla8_ha4_xor0;
  wire f_s_wallace_cla8_ha4_and0;
  wire f_s_wallace_cla8_fa28_xor0;
  wire f_s_wallace_cla8_fa28_and0;
  wire f_s_wallace_cla8_fa28_xor1;
  wire f_s_wallace_cla8_fa28_and1;
  wire f_s_wallace_cla8_fa28_or0;
  wire f_s_wallace_cla8_fa29_xor0;
  wire f_s_wallace_cla8_fa29_and0;
  wire f_s_wallace_cla8_fa29_xor1;
  wire f_s_wallace_cla8_fa29_and1;
  wire f_s_wallace_cla8_fa29_or0;
  wire f_s_wallace_cla8_ha5_xor0;
  wire f_s_wallace_cla8_ha5_and0;
  wire f_s_wallace_cla8_fa30_xor0;
  wire f_s_wallace_cla8_fa30_and0;
  wire f_s_wallace_cla8_fa30_xor1;
  wire f_s_wallace_cla8_fa30_and1;
  wire f_s_wallace_cla8_fa30_or0;
  wire f_s_wallace_cla8_fa31_xor0;
  wire f_s_wallace_cla8_fa31_and0;
  wire f_s_wallace_cla8_fa31_xor1;
  wire f_s_wallace_cla8_fa31_and1;
  wire f_s_wallace_cla8_fa31_or0;
  wire f_s_wallace_cla8_fa32_xor0;
  wire f_s_wallace_cla8_fa32_and0;
  wire f_s_wallace_cla8_fa32_xor1;
  wire f_s_wallace_cla8_fa32_and1;
  wire f_s_wallace_cla8_fa32_or0;
  wire f_s_wallace_cla8_fa33_xor0;
  wire f_s_wallace_cla8_fa33_and0;
  wire f_s_wallace_cla8_fa33_xor1;
  wire f_s_wallace_cla8_fa33_and1;
  wire f_s_wallace_cla8_fa33_or0;
  wire f_s_wallace_cla8_nand_5_7;
  wire f_s_wallace_cla8_fa34_xor0;
  wire f_s_wallace_cla8_fa34_and0;
  wire f_s_wallace_cla8_fa34_xor1;
  wire f_s_wallace_cla8_fa34_and1;
  wire f_s_wallace_cla8_fa34_or0;
  wire f_s_wallace_cla8_nand_7_6;
  wire f_s_wallace_cla8_fa35_xor0;
  wire f_s_wallace_cla8_fa35_and0;
  wire f_s_wallace_cla8_fa35_xor1;
  wire f_s_wallace_cla8_fa35_and1;
  wire f_s_wallace_cla8_fa35_or0;
  wire f_s_wallace_cla8_and_0_0;
  wire f_s_wallace_cla8_and_1_0;
  wire f_s_wallace_cla8_and_0_2;
  wire f_s_wallace_cla8_nand_6_7;
  wire f_s_wallace_cla8_and_0_1;
  wire f_s_wallace_cla8_and_7_7;
  wire f_s_wallace_cla8_u_cla14_pg_logic0_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic0_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic0_xor0;
  wire f_s_wallace_cla8_u_cla14_pg_logic1_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic1_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic1_xor0;
  wire f_s_wallace_cla8_u_cla14_xor1;
  wire f_s_wallace_cla8_u_cla14_and0;
  wire f_s_wallace_cla8_u_cla14_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic2_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic2_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic2_xor0;
  wire f_s_wallace_cla8_u_cla14_xor2;
  wire f_s_wallace_cla8_u_cla14_and1;
  wire f_s_wallace_cla8_u_cla14_and2;
  wire f_s_wallace_cla8_u_cla14_and3;
  wire f_s_wallace_cla8_u_cla14_and4;
  wire f_s_wallace_cla8_u_cla14_or1;
  wire f_s_wallace_cla8_u_cla14_or2;
  wire f_s_wallace_cla8_u_cla14_pg_logic3_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic3_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic3_xor0;
  wire f_s_wallace_cla8_u_cla14_xor3;
  wire f_s_wallace_cla8_u_cla14_and5;
  wire f_s_wallace_cla8_u_cla14_and6;
  wire f_s_wallace_cla8_u_cla14_and7;
  wire f_s_wallace_cla8_u_cla14_and8;
  wire f_s_wallace_cla8_u_cla14_and9;
  wire f_s_wallace_cla8_u_cla14_and10;
  wire f_s_wallace_cla8_u_cla14_and11;
  wire f_s_wallace_cla8_u_cla14_or3;
  wire f_s_wallace_cla8_u_cla14_or4;
  wire f_s_wallace_cla8_u_cla14_or5;
  wire f_s_wallace_cla8_u_cla14_pg_logic4_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic4_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic4_xor0;
  wire f_s_wallace_cla8_u_cla14_xor4;
  wire f_s_wallace_cla8_u_cla14_and12;
  wire f_s_wallace_cla8_u_cla14_or6;
  wire f_s_wallace_cla8_u_cla14_pg_logic5_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic5_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic5_xor0;
  wire f_s_wallace_cla8_u_cla14_xor5;
  wire f_s_wallace_cla8_u_cla14_and13;
  wire f_s_wallace_cla8_u_cla14_and14;
  wire f_s_wallace_cla8_u_cla14_and15;
  wire f_s_wallace_cla8_u_cla14_or7;
  wire f_s_wallace_cla8_u_cla14_or8;
  wire f_s_wallace_cla8_u_cla14_pg_logic6_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic6_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic6_xor0;
  wire f_s_wallace_cla8_u_cla14_xor6;
  wire f_s_wallace_cla8_u_cla14_and16;
  wire f_s_wallace_cla8_u_cla14_and17;
  wire f_s_wallace_cla8_u_cla14_and18;
  wire f_s_wallace_cla8_u_cla14_and19;
  wire f_s_wallace_cla8_u_cla14_and20;
  wire f_s_wallace_cla8_u_cla14_and21;
  wire f_s_wallace_cla8_u_cla14_or9;
  wire f_s_wallace_cla8_u_cla14_or10;
  wire f_s_wallace_cla8_u_cla14_or11;
  wire f_s_wallace_cla8_u_cla14_pg_logic7_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic7_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic7_xor0;
  wire f_s_wallace_cla8_u_cla14_xor7;
  wire f_s_wallace_cla8_u_cla14_and22;
  wire f_s_wallace_cla8_u_cla14_and23;
  wire f_s_wallace_cla8_u_cla14_and24;
  wire f_s_wallace_cla8_u_cla14_and25;
  wire f_s_wallace_cla8_u_cla14_and26;
  wire f_s_wallace_cla8_u_cla14_and27;
  wire f_s_wallace_cla8_u_cla14_and28;
  wire f_s_wallace_cla8_u_cla14_and29;
  wire f_s_wallace_cla8_u_cla14_and30;
  wire f_s_wallace_cla8_u_cla14_and31;
  wire f_s_wallace_cla8_u_cla14_or12;
  wire f_s_wallace_cla8_u_cla14_or13;
  wire f_s_wallace_cla8_u_cla14_or14;
  wire f_s_wallace_cla8_u_cla14_or15;
  wire f_s_wallace_cla8_u_cla14_pg_logic8_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic8_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic8_xor0;
  wire f_s_wallace_cla8_u_cla14_xor8;
  wire f_s_wallace_cla8_u_cla14_and32;
  wire f_s_wallace_cla8_u_cla14_or16;
  wire f_s_wallace_cla8_u_cla14_pg_logic9_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic9_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic9_xor0;
  wire f_s_wallace_cla8_u_cla14_xor9;
  wire f_s_wallace_cla8_u_cla14_and33;
  wire f_s_wallace_cla8_u_cla14_and34;
  wire f_s_wallace_cla8_u_cla14_and35;
  wire f_s_wallace_cla8_u_cla14_or17;
  wire f_s_wallace_cla8_u_cla14_or18;
  wire f_s_wallace_cla8_u_cla14_pg_logic10_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic10_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic10_xor0;
  wire f_s_wallace_cla8_u_cla14_xor10;
  wire f_s_wallace_cla8_u_cla14_and36;
  wire f_s_wallace_cla8_u_cla14_and37;
  wire f_s_wallace_cla8_u_cla14_and38;
  wire f_s_wallace_cla8_u_cla14_and39;
  wire f_s_wallace_cla8_u_cla14_and40;
  wire f_s_wallace_cla8_u_cla14_and41;
  wire f_s_wallace_cla8_u_cla14_or19;
  wire f_s_wallace_cla8_u_cla14_or20;
  wire f_s_wallace_cla8_u_cla14_or21;
  wire f_s_wallace_cla8_u_cla14_pg_logic11_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic11_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic11_xor0;
  wire f_s_wallace_cla8_u_cla14_xor11;
  wire f_s_wallace_cla8_u_cla14_and42;
  wire f_s_wallace_cla8_u_cla14_and43;
  wire f_s_wallace_cla8_u_cla14_and44;
  wire f_s_wallace_cla8_u_cla14_and45;
  wire f_s_wallace_cla8_u_cla14_and46;
  wire f_s_wallace_cla8_u_cla14_and47;
  wire f_s_wallace_cla8_u_cla14_and48;
  wire f_s_wallace_cla8_u_cla14_and49;
  wire f_s_wallace_cla8_u_cla14_and50;
  wire f_s_wallace_cla8_u_cla14_and51;
  wire f_s_wallace_cla8_u_cla14_or22;
  wire f_s_wallace_cla8_u_cla14_or23;
  wire f_s_wallace_cla8_u_cla14_or24;
  wire f_s_wallace_cla8_u_cla14_or25;
  wire f_s_wallace_cla8_u_cla14_pg_logic12_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic12_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic12_xor0;
  wire f_s_wallace_cla8_u_cla14_xor12;
  wire f_s_wallace_cla8_u_cla14_and52;
  wire f_s_wallace_cla8_u_cla14_or26;
  wire f_s_wallace_cla8_u_cla14_pg_logic13_or0;
  wire f_s_wallace_cla8_u_cla14_pg_logic13_and0;
  wire f_s_wallace_cla8_u_cla14_pg_logic13_xor0;
  wire f_s_wallace_cla8_u_cla14_xor13;
  wire f_s_wallace_cla8_u_cla14_and53;
  wire f_s_wallace_cla8_u_cla14_and54;
  wire f_s_wallace_cla8_u_cla14_and55;
  wire f_s_wallace_cla8_u_cla14_or27;
  wire f_s_wallace_cla8_u_cla14_or28;
  wire f_s_wallace_cla8_xor0;

  assign f_s_wallace_cla8_and_2_0 = a[2] & b[0];
  assign f_s_wallace_cla8_and_1_1 = a[1] & b[1];
  assign f_s_wallace_cla8_ha0_xor0 = f_s_wallace_cla8_and_2_0 ^ f_s_wallace_cla8_and_1_1;
  assign f_s_wallace_cla8_ha0_and0 = f_s_wallace_cla8_and_2_0 & f_s_wallace_cla8_and_1_1;
  assign f_s_wallace_cla8_and_3_0 = a[3] & b[0];
  assign f_s_wallace_cla8_and_2_1 = a[2] & b[1];
  assign f_s_wallace_cla8_fa0_xor0 = f_s_wallace_cla8_ha0_and0 ^ f_s_wallace_cla8_and_3_0;
  assign f_s_wallace_cla8_fa0_and0 = f_s_wallace_cla8_ha0_and0 & f_s_wallace_cla8_and_3_0;
  assign f_s_wallace_cla8_fa0_xor1 = f_s_wallace_cla8_fa0_xor0 ^ f_s_wallace_cla8_and_2_1;
  assign f_s_wallace_cla8_fa0_and1 = f_s_wallace_cla8_fa0_xor0 & f_s_wallace_cla8_and_2_1;
  assign f_s_wallace_cla8_fa0_or0 = f_s_wallace_cla8_fa0_and0 | f_s_wallace_cla8_fa0_and1;
  assign f_s_wallace_cla8_and_4_0 = a[4] & b[0];
  assign f_s_wallace_cla8_and_3_1 = a[3] & b[1];
  assign f_s_wallace_cla8_fa1_xor0 = f_s_wallace_cla8_fa0_or0 ^ f_s_wallace_cla8_and_4_0;
  assign f_s_wallace_cla8_fa1_and0 = f_s_wallace_cla8_fa0_or0 & f_s_wallace_cla8_and_4_0;
  assign f_s_wallace_cla8_fa1_xor1 = f_s_wallace_cla8_fa1_xor0 ^ f_s_wallace_cla8_and_3_1;
  assign f_s_wallace_cla8_fa1_and1 = f_s_wallace_cla8_fa1_xor0 & f_s_wallace_cla8_and_3_1;
  assign f_s_wallace_cla8_fa1_or0 = f_s_wallace_cla8_fa1_and0 | f_s_wallace_cla8_fa1_and1;
  assign f_s_wallace_cla8_and_5_0 = a[5] & b[0];
  assign f_s_wallace_cla8_and_4_1 = a[4] & b[1];
  assign f_s_wallace_cla8_fa2_xor0 = f_s_wallace_cla8_fa1_or0 ^ f_s_wallace_cla8_and_5_0;
  assign f_s_wallace_cla8_fa2_and0 = f_s_wallace_cla8_fa1_or0 & f_s_wallace_cla8_and_5_0;
  assign f_s_wallace_cla8_fa2_xor1 = f_s_wallace_cla8_fa2_xor0 ^ f_s_wallace_cla8_and_4_1;
  assign f_s_wallace_cla8_fa2_and1 = f_s_wallace_cla8_fa2_xor0 & f_s_wallace_cla8_and_4_1;
  assign f_s_wallace_cla8_fa2_or0 = f_s_wallace_cla8_fa2_and0 | f_s_wallace_cla8_fa2_and1;
  assign f_s_wallace_cla8_and_6_0 = a[6] & b[0];
  assign f_s_wallace_cla8_and_5_1 = a[5] & b[1];
  assign f_s_wallace_cla8_fa3_xor0 = f_s_wallace_cla8_fa2_or0 ^ f_s_wallace_cla8_and_6_0;
  assign f_s_wallace_cla8_fa3_and0 = f_s_wallace_cla8_fa2_or0 & f_s_wallace_cla8_and_6_0;
  assign f_s_wallace_cla8_fa3_xor1 = f_s_wallace_cla8_fa3_xor0 ^ f_s_wallace_cla8_and_5_1;
  assign f_s_wallace_cla8_fa3_and1 = f_s_wallace_cla8_fa3_xor0 & f_s_wallace_cla8_and_5_1;
  assign f_s_wallace_cla8_fa3_or0 = f_s_wallace_cla8_fa3_and0 | f_s_wallace_cla8_fa3_and1;
  assign f_s_wallace_cla8_nand_7_0 = ~(a[7] & b[0]);
  assign f_s_wallace_cla8_and_6_1 = a[6] & b[1];
  assign f_s_wallace_cla8_fa4_xor0 = f_s_wallace_cla8_fa3_or0 ^ f_s_wallace_cla8_nand_7_0;
  assign f_s_wallace_cla8_fa4_and0 = f_s_wallace_cla8_fa3_or0 & f_s_wallace_cla8_nand_7_0;
  assign f_s_wallace_cla8_fa4_xor1 = f_s_wallace_cla8_fa4_xor0 ^ f_s_wallace_cla8_and_6_1;
  assign f_s_wallace_cla8_fa4_and1 = f_s_wallace_cla8_fa4_xor0 & f_s_wallace_cla8_and_6_1;
  assign f_s_wallace_cla8_fa4_or0 = f_s_wallace_cla8_fa4_and0 | f_s_wallace_cla8_fa4_and1;
  assign f_s_wallace_cla8_nand_7_1 = ~(a[7] & b[1]);
  assign f_s_wallace_cla8_fa5_xor0 = ~f_s_wallace_cla8_fa4_or0;
  assign f_s_wallace_cla8_fa5_xor1 = f_s_wallace_cla8_fa5_xor0 ^ f_s_wallace_cla8_nand_7_1;
  assign f_s_wallace_cla8_fa5_and1 = f_s_wallace_cla8_fa5_xor0 & f_s_wallace_cla8_nand_7_1;
  assign f_s_wallace_cla8_fa5_or0 = f_s_wallace_cla8_fa4_or0 | f_s_wallace_cla8_fa5_and1;
  assign f_s_wallace_cla8_nand_7_2 = ~(a[7] & b[2]);
  assign f_s_wallace_cla8_and_6_3 = a[6] & b[3];
  assign f_s_wallace_cla8_fa6_xor0 = f_s_wallace_cla8_fa5_or0 ^ f_s_wallace_cla8_nand_7_2;
  assign f_s_wallace_cla8_fa6_and0 = f_s_wallace_cla8_fa5_or0 & f_s_wallace_cla8_nand_7_2;
  assign f_s_wallace_cla8_fa6_xor1 = f_s_wallace_cla8_fa6_xor0 ^ f_s_wallace_cla8_and_6_3;
  assign f_s_wallace_cla8_fa6_and1 = f_s_wallace_cla8_fa6_xor0 & f_s_wallace_cla8_and_6_3;
  assign f_s_wallace_cla8_fa6_or0 = f_s_wallace_cla8_fa6_and0 | f_s_wallace_cla8_fa6_and1;
  assign f_s_wallace_cla8_nand_7_3 = ~(a[7] & b[3]);
  assign f_s_wallace_cla8_and_6_4 = a[6] & b[4];
  assign f_s_wallace_cla8_fa7_xor0 = f_s_wallace_cla8_fa6_or0 ^ f_s_wallace_cla8_nand_7_3;
  assign f_s_wallace_cla8_fa7_and0 = f_s_wallace_cla8_fa6_or0 & f_s_wallace_cla8_nand_7_3;
  assign f_s_wallace_cla8_fa7_xor1 = f_s_wallace_cla8_fa7_xor0 ^ f_s_wallace_cla8_and_6_4;
  assign f_s_wallace_cla8_fa7_and1 = f_s_wallace_cla8_fa7_xor0 & f_s_wallace_cla8_and_6_4;
  assign f_s_wallace_cla8_fa7_or0 = f_s_wallace_cla8_fa7_and0 | f_s_wallace_cla8_fa7_and1;
  assign f_s_wallace_cla8_nand_7_4 = ~(a[7] & b[4]);
  assign f_s_wallace_cla8_and_6_5 = a[6] & b[5];
  assign f_s_wallace_cla8_fa8_xor0 = f_s_wallace_cla8_fa7_or0 ^ f_s_wallace_cla8_nand_7_4;
  assign f_s_wallace_cla8_fa8_and0 = f_s_wallace_cla8_fa7_or0 & f_s_wallace_cla8_nand_7_4;
  assign f_s_wallace_cla8_fa8_xor1 = f_s_wallace_cla8_fa8_xor0 ^ f_s_wallace_cla8_and_6_5;
  assign f_s_wallace_cla8_fa8_and1 = f_s_wallace_cla8_fa8_xor0 & f_s_wallace_cla8_and_6_5;
  assign f_s_wallace_cla8_fa8_or0 = f_s_wallace_cla8_fa8_and0 | f_s_wallace_cla8_fa8_and1;
  assign f_s_wallace_cla8_nand_7_5 = ~(a[7] & b[5]);
  assign f_s_wallace_cla8_and_6_6 = a[6] & b[6];
  assign f_s_wallace_cla8_fa9_xor0 = f_s_wallace_cla8_fa8_or0 ^ f_s_wallace_cla8_nand_7_5;
  assign f_s_wallace_cla8_fa9_and0 = f_s_wallace_cla8_fa8_or0 & f_s_wallace_cla8_nand_7_5;
  assign f_s_wallace_cla8_fa9_xor1 = f_s_wallace_cla8_fa9_xor0 ^ f_s_wallace_cla8_and_6_6;
  assign f_s_wallace_cla8_fa9_and1 = f_s_wallace_cla8_fa9_xor0 & f_s_wallace_cla8_and_6_6;
  assign f_s_wallace_cla8_fa9_or0 = f_s_wallace_cla8_fa9_and0 | f_s_wallace_cla8_fa9_and1;
  assign f_s_wallace_cla8_and_1_2 = a[1] & b[2];
  assign f_s_wallace_cla8_and_0_3 = a[0] & b[3];
  assign f_s_wallace_cla8_ha1_xor0 = f_s_wallace_cla8_and_1_2 ^ f_s_wallace_cla8_and_0_3;
  assign f_s_wallace_cla8_ha1_and0 = f_s_wallace_cla8_and_1_2 & f_s_wallace_cla8_and_0_3;
  assign f_s_wallace_cla8_and_2_2 = a[2] & b[2];
  assign f_s_wallace_cla8_and_1_3 = a[1] & b[3];
  assign f_s_wallace_cla8_fa10_xor0 = f_s_wallace_cla8_ha1_and0 ^ f_s_wallace_cla8_and_2_2;
  assign f_s_wallace_cla8_fa10_and0 = f_s_wallace_cla8_ha1_and0 & f_s_wallace_cla8_and_2_2;
  assign f_s_wallace_cla8_fa10_xor1 = f_s_wallace_cla8_fa10_xor0 ^ f_s_wallace_cla8_and_1_3;
  assign f_s_wallace_cla8_fa10_and1 = f_s_wallace_cla8_fa10_xor0 & f_s_wallace_cla8_and_1_3;
  assign f_s_wallace_cla8_fa10_or0 = f_s_wallace_cla8_fa10_and0 | f_s_wallace_cla8_fa10_and1;
  assign f_s_wallace_cla8_and_3_2 = a[3] & b[2];
  assign f_s_wallace_cla8_and_2_3 = a[2] & b[3];
  assign f_s_wallace_cla8_fa11_xor0 = f_s_wallace_cla8_fa10_or0 ^ f_s_wallace_cla8_and_3_2;
  assign f_s_wallace_cla8_fa11_and0 = f_s_wallace_cla8_fa10_or0 & f_s_wallace_cla8_and_3_2;
  assign f_s_wallace_cla8_fa11_xor1 = f_s_wallace_cla8_fa11_xor0 ^ f_s_wallace_cla8_and_2_3;
  assign f_s_wallace_cla8_fa11_and1 = f_s_wallace_cla8_fa11_xor0 & f_s_wallace_cla8_and_2_3;
  assign f_s_wallace_cla8_fa11_or0 = f_s_wallace_cla8_fa11_and0 | f_s_wallace_cla8_fa11_and1;
  assign f_s_wallace_cla8_and_4_2 = a[4] & b[2];
  assign f_s_wallace_cla8_and_3_3 = a[3] & b[3];
  assign f_s_wallace_cla8_fa12_xor0 = f_s_wallace_cla8_fa11_or0 ^ f_s_wallace_cla8_and_4_2;
  assign f_s_wallace_cla8_fa12_and0 = f_s_wallace_cla8_fa11_or0 & f_s_wallace_cla8_and_4_2;
  assign f_s_wallace_cla8_fa12_xor1 = f_s_wallace_cla8_fa12_xor0 ^ f_s_wallace_cla8_and_3_3;
  assign f_s_wallace_cla8_fa12_and1 = f_s_wallace_cla8_fa12_xor0 & f_s_wallace_cla8_and_3_3;
  assign f_s_wallace_cla8_fa12_or0 = f_s_wallace_cla8_fa12_and0 | f_s_wallace_cla8_fa12_and1;
  assign f_s_wallace_cla8_and_5_2 = a[5] & b[2];
  assign f_s_wallace_cla8_and_4_3 = a[4] & b[3];
  assign f_s_wallace_cla8_fa13_xor0 = f_s_wallace_cla8_fa12_or0 ^ f_s_wallace_cla8_and_5_2;
  assign f_s_wallace_cla8_fa13_and0 = f_s_wallace_cla8_fa12_or0 & f_s_wallace_cla8_and_5_2;
  assign f_s_wallace_cla8_fa13_xor1 = f_s_wallace_cla8_fa13_xor0 ^ f_s_wallace_cla8_and_4_3;
  assign f_s_wallace_cla8_fa13_and1 = f_s_wallace_cla8_fa13_xor0 & f_s_wallace_cla8_and_4_3;
  assign f_s_wallace_cla8_fa13_or0 = f_s_wallace_cla8_fa13_and0 | f_s_wallace_cla8_fa13_and1;
  assign f_s_wallace_cla8_and_6_2 = a[6] & b[2];
  assign f_s_wallace_cla8_and_5_3 = a[5] & b[3];
  assign f_s_wallace_cla8_fa14_xor0 = f_s_wallace_cla8_fa13_or0 ^ f_s_wallace_cla8_and_6_2;
  assign f_s_wallace_cla8_fa14_and0 = f_s_wallace_cla8_fa13_or0 & f_s_wallace_cla8_and_6_2;
  assign f_s_wallace_cla8_fa14_xor1 = f_s_wallace_cla8_fa14_xor0 ^ f_s_wallace_cla8_and_5_3;
  assign f_s_wallace_cla8_fa14_and1 = f_s_wallace_cla8_fa14_xor0 & f_s_wallace_cla8_and_5_3;
  assign f_s_wallace_cla8_fa14_or0 = f_s_wallace_cla8_fa14_and0 | f_s_wallace_cla8_fa14_and1;
  assign f_s_wallace_cla8_and_5_4 = a[5] & b[4];
  assign f_s_wallace_cla8_and_4_5 = a[4] & b[5];
  assign f_s_wallace_cla8_fa15_xor0 = f_s_wallace_cla8_fa14_or0 ^ f_s_wallace_cla8_and_5_4;
  assign f_s_wallace_cla8_fa15_and0 = f_s_wallace_cla8_fa14_or0 & f_s_wallace_cla8_and_5_4;
  assign f_s_wallace_cla8_fa15_xor1 = f_s_wallace_cla8_fa15_xor0 ^ f_s_wallace_cla8_and_4_5;
  assign f_s_wallace_cla8_fa15_and1 = f_s_wallace_cla8_fa15_xor0 & f_s_wallace_cla8_and_4_5;
  assign f_s_wallace_cla8_fa15_or0 = f_s_wallace_cla8_fa15_and0 | f_s_wallace_cla8_fa15_and1;
  assign f_s_wallace_cla8_and_5_5 = a[5] & b[5];
  assign f_s_wallace_cla8_and_4_6 = a[4] & b[6];
  assign f_s_wallace_cla8_fa16_xor0 = f_s_wallace_cla8_fa15_or0 ^ f_s_wallace_cla8_and_5_5;
  assign f_s_wallace_cla8_fa16_and0 = f_s_wallace_cla8_fa15_or0 & f_s_wallace_cla8_and_5_5;
  assign f_s_wallace_cla8_fa16_xor1 = f_s_wallace_cla8_fa16_xor0 ^ f_s_wallace_cla8_and_4_6;
  assign f_s_wallace_cla8_fa16_and1 = f_s_wallace_cla8_fa16_xor0 & f_s_wallace_cla8_and_4_6;
  assign f_s_wallace_cla8_fa16_or0 = f_s_wallace_cla8_fa16_and0 | f_s_wallace_cla8_fa16_and1;
  assign f_s_wallace_cla8_and_5_6 = a[5] & b[6];
  assign f_s_wallace_cla8_nand_4_7 = ~(a[4] & b[7]);
  assign f_s_wallace_cla8_fa17_xor0 = f_s_wallace_cla8_fa16_or0 ^ f_s_wallace_cla8_and_5_6;
  assign f_s_wallace_cla8_fa17_and0 = f_s_wallace_cla8_fa16_or0 & f_s_wallace_cla8_and_5_6;
  assign f_s_wallace_cla8_fa17_xor1 = f_s_wallace_cla8_fa17_xor0 ^ f_s_wallace_cla8_nand_4_7;
  assign f_s_wallace_cla8_fa17_and1 = f_s_wallace_cla8_fa17_xor0 & f_s_wallace_cla8_nand_4_7;
  assign f_s_wallace_cla8_fa17_or0 = f_s_wallace_cla8_fa17_and0 | f_s_wallace_cla8_fa17_and1;
  assign f_s_wallace_cla8_and_0_4 = a[0] & b[4];
  assign f_s_wallace_cla8_ha2_xor0 = f_s_wallace_cla8_and_0_4 ^ f_s_wallace_cla8_fa1_xor1;
  assign f_s_wallace_cla8_ha2_and0 = f_s_wallace_cla8_and_0_4 & f_s_wallace_cla8_fa1_xor1;
  assign f_s_wallace_cla8_and_1_4 = a[1] & b[4];
  assign f_s_wallace_cla8_and_0_5 = a[0] & b[5];
  assign f_s_wallace_cla8_fa18_xor0 = f_s_wallace_cla8_ha2_and0 ^ f_s_wallace_cla8_and_1_4;
  assign f_s_wallace_cla8_fa18_and0 = f_s_wallace_cla8_ha2_and0 & f_s_wallace_cla8_and_1_4;
  assign f_s_wallace_cla8_fa18_xor1 = f_s_wallace_cla8_fa18_xor0 ^ f_s_wallace_cla8_and_0_5;
  assign f_s_wallace_cla8_fa18_and1 = f_s_wallace_cla8_fa18_xor0 & f_s_wallace_cla8_and_0_5;
  assign f_s_wallace_cla8_fa18_or0 = f_s_wallace_cla8_fa18_and0 | f_s_wallace_cla8_fa18_and1;
  assign f_s_wallace_cla8_and_2_4 = a[2] & b[4];
  assign f_s_wallace_cla8_and_1_5 = a[1] & b[5];
  assign f_s_wallace_cla8_fa19_xor0 = f_s_wallace_cla8_fa18_or0 ^ f_s_wallace_cla8_and_2_4;
  assign f_s_wallace_cla8_fa19_and0 = f_s_wallace_cla8_fa18_or0 & f_s_wallace_cla8_and_2_4;
  assign f_s_wallace_cla8_fa19_xor1 = f_s_wallace_cla8_fa19_xor0 ^ f_s_wallace_cla8_and_1_5;
  assign f_s_wallace_cla8_fa19_and1 = f_s_wallace_cla8_fa19_xor0 & f_s_wallace_cla8_and_1_5;
  assign f_s_wallace_cla8_fa19_or0 = f_s_wallace_cla8_fa19_and0 | f_s_wallace_cla8_fa19_and1;
  assign f_s_wallace_cla8_and_3_4 = a[3] & b[4];
  assign f_s_wallace_cla8_and_2_5 = a[2] & b[5];
  assign f_s_wallace_cla8_fa20_xor0 = f_s_wallace_cla8_fa19_or0 ^ f_s_wallace_cla8_and_3_4;
  assign f_s_wallace_cla8_fa20_and0 = f_s_wallace_cla8_fa19_or0 & f_s_wallace_cla8_and_3_4;
  assign f_s_wallace_cla8_fa20_xor1 = f_s_wallace_cla8_fa20_xor0 ^ f_s_wallace_cla8_and_2_5;
  assign f_s_wallace_cla8_fa20_and1 = f_s_wallace_cla8_fa20_xor0 & f_s_wallace_cla8_and_2_5;
  assign f_s_wallace_cla8_fa20_or0 = f_s_wallace_cla8_fa20_and0 | f_s_wallace_cla8_fa20_and1;
  assign f_s_wallace_cla8_and_4_4 = a[4] & b[4];
  assign f_s_wallace_cla8_and_3_5 = a[3] & b[5];
  assign f_s_wallace_cla8_fa21_xor0 = f_s_wallace_cla8_fa20_or0 ^ f_s_wallace_cla8_and_4_4;
  assign f_s_wallace_cla8_fa21_and0 = f_s_wallace_cla8_fa20_or0 & f_s_wallace_cla8_and_4_4;
  assign f_s_wallace_cla8_fa21_xor1 = f_s_wallace_cla8_fa21_xor0 ^ f_s_wallace_cla8_and_3_5;
  assign f_s_wallace_cla8_fa21_and1 = f_s_wallace_cla8_fa21_xor0 & f_s_wallace_cla8_and_3_5;
  assign f_s_wallace_cla8_fa21_or0 = f_s_wallace_cla8_fa21_and0 | f_s_wallace_cla8_fa21_and1;
  assign f_s_wallace_cla8_and_3_6 = a[3] & b[6];
  assign f_s_wallace_cla8_nand_2_7 = ~(a[2] & b[7]);
  assign f_s_wallace_cla8_fa22_xor0 = f_s_wallace_cla8_fa21_or0 ^ f_s_wallace_cla8_and_3_6;
  assign f_s_wallace_cla8_fa22_and0 = f_s_wallace_cla8_fa21_or0 & f_s_wallace_cla8_and_3_6;
  assign f_s_wallace_cla8_fa22_xor1 = f_s_wallace_cla8_fa22_xor0 ^ f_s_wallace_cla8_nand_2_7;
  assign f_s_wallace_cla8_fa22_and1 = f_s_wallace_cla8_fa22_xor0 & f_s_wallace_cla8_nand_2_7;
  assign f_s_wallace_cla8_fa22_or0 = f_s_wallace_cla8_fa22_and0 | f_s_wallace_cla8_fa22_and1;
  assign f_s_wallace_cla8_nand_3_7 = ~(a[3] & b[7]);
  assign f_s_wallace_cla8_fa23_xor0 = f_s_wallace_cla8_fa22_or0 ^ f_s_wallace_cla8_nand_3_7;
  assign f_s_wallace_cla8_fa23_and0 = f_s_wallace_cla8_fa22_or0 & f_s_wallace_cla8_nand_3_7;
  assign f_s_wallace_cla8_fa23_xor1 = f_s_wallace_cla8_fa23_xor0 ^ f_s_wallace_cla8_fa7_xor1;
  assign f_s_wallace_cla8_fa23_and1 = f_s_wallace_cla8_fa23_xor0 & f_s_wallace_cla8_fa7_xor1;
  assign f_s_wallace_cla8_fa23_or0 = f_s_wallace_cla8_fa23_and0 | f_s_wallace_cla8_fa23_and1;
  assign f_s_wallace_cla8_ha3_xor0 = f_s_wallace_cla8_fa2_xor1 ^ f_s_wallace_cla8_fa11_xor1;
  assign f_s_wallace_cla8_ha3_and0 = f_s_wallace_cla8_fa2_xor1 & f_s_wallace_cla8_fa11_xor1;
  assign f_s_wallace_cla8_and_0_6 = a[0] & b[6];
  assign f_s_wallace_cla8_fa24_xor0 = f_s_wallace_cla8_ha3_and0 ^ f_s_wallace_cla8_and_0_6;
  assign f_s_wallace_cla8_fa24_and0 = f_s_wallace_cla8_ha3_and0 & f_s_wallace_cla8_and_0_6;
  assign f_s_wallace_cla8_fa24_xor1 = f_s_wallace_cla8_fa24_xor0 ^ f_s_wallace_cla8_fa3_xor1;
  assign f_s_wallace_cla8_fa24_and1 = f_s_wallace_cla8_fa24_xor0 & f_s_wallace_cla8_fa3_xor1;
  assign f_s_wallace_cla8_fa24_or0 = f_s_wallace_cla8_fa24_and0 | f_s_wallace_cla8_fa24_and1;
  assign f_s_wallace_cla8_and_1_6 = a[1] & b[6];
  assign f_s_wallace_cla8_nand_0_7 = ~(a[0] & b[7]);
  assign f_s_wallace_cla8_fa25_xor0 = f_s_wallace_cla8_fa24_or0 ^ f_s_wallace_cla8_and_1_6;
  assign f_s_wallace_cla8_fa25_and0 = f_s_wallace_cla8_fa24_or0 & f_s_wallace_cla8_and_1_6;
  assign f_s_wallace_cla8_fa25_xor1 = f_s_wallace_cla8_fa25_xor0 ^ f_s_wallace_cla8_nand_0_7;
  assign f_s_wallace_cla8_fa25_and1 = f_s_wallace_cla8_fa25_xor0 & f_s_wallace_cla8_nand_0_7;
  assign f_s_wallace_cla8_fa25_or0 = f_s_wallace_cla8_fa25_and0 | f_s_wallace_cla8_fa25_and1;
  assign f_s_wallace_cla8_and_2_6 = a[2] & b[6];
  assign f_s_wallace_cla8_nand_1_7 = ~(a[1] & b[7]);
  assign f_s_wallace_cla8_fa26_xor0 = f_s_wallace_cla8_fa25_or0 ^ f_s_wallace_cla8_and_2_6;
  assign f_s_wallace_cla8_fa26_and0 = f_s_wallace_cla8_fa25_or0 & f_s_wallace_cla8_and_2_6;
  assign f_s_wallace_cla8_fa26_xor1 = f_s_wallace_cla8_fa26_xor0 ^ f_s_wallace_cla8_nand_1_7;
  assign f_s_wallace_cla8_fa26_and1 = f_s_wallace_cla8_fa26_xor0 & f_s_wallace_cla8_nand_1_7;
  assign f_s_wallace_cla8_fa26_or0 = f_s_wallace_cla8_fa26_and0 | f_s_wallace_cla8_fa26_and1;
  assign f_s_wallace_cla8_fa27_xor0 = f_s_wallace_cla8_fa26_or0 ^ f_s_wallace_cla8_fa6_xor1;
  assign f_s_wallace_cla8_fa27_and0 = f_s_wallace_cla8_fa26_or0 & f_s_wallace_cla8_fa6_xor1;
  assign f_s_wallace_cla8_fa27_xor1 = f_s_wallace_cla8_fa27_xor0 ^ f_s_wallace_cla8_fa15_xor1;
  assign f_s_wallace_cla8_fa27_and1 = f_s_wallace_cla8_fa27_xor0 & f_s_wallace_cla8_fa15_xor1;
  assign f_s_wallace_cla8_fa27_or0 = f_s_wallace_cla8_fa27_and0 | f_s_wallace_cla8_fa27_and1;
  assign f_s_wallace_cla8_ha4_xor0 = f_s_wallace_cla8_fa12_xor1 ^ f_s_wallace_cla8_fa19_xor1;
  assign f_s_wallace_cla8_ha4_and0 = f_s_wallace_cla8_fa12_xor1 & f_s_wallace_cla8_fa19_xor1;
  assign f_s_wallace_cla8_fa28_xor0 = f_s_wallace_cla8_ha4_and0 ^ f_s_wallace_cla8_fa4_xor1;
  assign f_s_wallace_cla8_fa28_and0 = f_s_wallace_cla8_ha4_and0 & f_s_wallace_cla8_fa4_xor1;
  assign f_s_wallace_cla8_fa28_xor1 = f_s_wallace_cla8_fa28_xor0 ^ f_s_wallace_cla8_fa13_xor1;
  assign f_s_wallace_cla8_fa28_and1 = f_s_wallace_cla8_fa28_xor0 & f_s_wallace_cla8_fa13_xor1;
  assign f_s_wallace_cla8_fa28_or0 = f_s_wallace_cla8_fa28_and0 | f_s_wallace_cla8_fa28_and1;
  assign f_s_wallace_cla8_fa29_xor0 = f_s_wallace_cla8_fa28_or0 ^ f_s_wallace_cla8_fa5_xor1;
  assign f_s_wallace_cla8_fa29_and0 = f_s_wallace_cla8_fa28_or0 & f_s_wallace_cla8_fa5_xor1;
  assign f_s_wallace_cla8_fa29_xor1 = f_s_wallace_cla8_fa29_xor0 ^ f_s_wallace_cla8_fa14_xor1;
  assign f_s_wallace_cla8_fa29_and1 = f_s_wallace_cla8_fa29_xor0 & f_s_wallace_cla8_fa14_xor1;
  assign f_s_wallace_cla8_fa29_or0 = f_s_wallace_cla8_fa29_and0 | f_s_wallace_cla8_fa29_and1;
  assign f_s_wallace_cla8_ha5_xor0 = f_s_wallace_cla8_fa20_xor1 ^ f_s_wallace_cla8_fa25_xor1;
  assign f_s_wallace_cla8_ha5_and0 = f_s_wallace_cla8_fa20_xor1 & f_s_wallace_cla8_fa25_xor1;
  assign f_s_wallace_cla8_fa30_xor0 = f_s_wallace_cla8_ha5_and0 ^ f_s_wallace_cla8_fa21_xor1;
  assign f_s_wallace_cla8_fa30_and0 = f_s_wallace_cla8_ha5_and0 & f_s_wallace_cla8_fa21_xor1;
  assign f_s_wallace_cla8_fa30_xor1 = f_s_wallace_cla8_fa30_xor0 ^ f_s_wallace_cla8_fa26_xor1;
  assign f_s_wallace_cla8_fa30_and1 = f_s_wallace_cla8_fa30_xor0 & f_s_wallace_cla8_fa26_xor1;
  assign f_s_wallace_cla8_fa30_or0 = f_s_wallace_cla8_fa30_and0 | f_s_wallace_cla8_fa30_and1;
  assign f_s_wallace_cla8_fa31_xor0 = f_s_wallace_cla8_fa30_or0 ^ f_s_wallace_cla8_fa29_or0;
  assign f_s_wallace_cla8_fa31_and0 = f_s_wallace_cla8_fa30_or0 & f_s_wallace_cla8_fa29_or0;
  assign f_s_wallace_cla8_fa31_xor1 = f_s_wallace_cla8_fa31_xor0 ^ f_s_wallace_cla8_fa22_xor1;
  assign f_s_wallace_cla8_fa31_and1 = f_s_wallace_cla8_fa31_xor0 & f_s_wallace_cla8_fa22_xor1;
  assign f_s_wallace_cla8_fa31_or0 = f_s_wallace_cla8_fa31_and0 | f_s_wallace_cla8_fa31_and1;
  assign f_s_wallace_cla8_fa32_xor0 = f_s_wallace_cla8_fa31_or0 ^ f_s_wallace_cla8_fa27_or0;
  assign f_s_wallace_cla8_fa32_and0 = f_s_wallace_cla8_fa31_or0 & f_s_wallace_cla8_fa27_or0;
  assign f_s_wallace_cla8_fa32_xor1 = f_s_wallace_cla8_fa32_xor0 ^ f_s_wallace_cla8_fa16_xor1;
  assign f_s_wallace_cla8_fa32_and1 = f_s_wallace_cla8_fa32_xor0 & f_s_wallace_cla8_fa16_xor1;
  assign f_s_wallace_cla8_fa32_or0 = f_s_wallace_cla8_fa32_and0 | f_s_wallace_cla8_fa32_and1;
  assign f_s_wallace_cla8_fa33_xor0 = f_s_wallace_cla8_fa32_or0 ^ f_s_wallace_cla8_fa23_or0;
  assign f_s_wallace_cla8_fa33_and0 = f_s_wallace_cla8_fa32_or0 & f_s_wallace_cla8_fa23_or0;
  assign f_s_wallace_cla8_fa33_xor1 = f_s_wallace_cla8_fa33_xor0 ^ f_s_wallace_cla8_fa8_xor1;
  assign f_s_wallace_cla8_fa33_and1 = f_s_wallace_cla8_fa33_xor0 & f_s_wallace_cla8_fa8_xor1;
  assign f_s_wallace_cla8_fa33_or0 = f_s_wallace_cla8_fa33_and0 | f_s_wallace_cla8_fa33_and1;
  assign f_s_wallace_cla8_nand_5_7 = ~(a[5] & b[7]);
  assign f_s_wallace_cla8_fa34_xor0 = f_s_wallace_cla8_fa33_or0 ^ f_s_wallace_cla8_fa17_or0;
  assign f_s_wallace_cla8_fa34_and0 = f_s_wallace_cla8_fa33_or0 & f_s_wallace_cla8_fa17_or0;
  assign f_s_wallace_cla8_fa34_xor1 = f_s_wallace_cla8_fa34_xor0 ^ f_s_wallace_cla8_nand_5_7;
  assign f_s_wallace_cla8_fa34_and1 = f_s_wallace_cla8_fa34_xor0 & f_s_wallace_cla8_nand_5_7;
  assign f_s_wallace_cla8_fa34_or0 = f_s_wallace_cla8_fa34_and0 | f_s_wallace_cla8_fa34_and1;
  assign f_s_wallace_cla8_nand_7_6 = ~(a[7] & b[6]);
  assign f_s_wallace_cla8_fa35_xor0 = f_s_wallace_cla8_fa34_or0 ^ f_s_wallace_cla8_fa9_or0;
  assign f_s_wallace_cla8_fa35_and0 = f_s_wallace_cla8_fa34_or0 & f_s_wallace_cla8_fa9_or0;
  assign f_s_wallace_cla8_fa35_xor1 = f_s_wallace_cla8_fa35_xor0 ^ f_s_wallace_cla8_nand_7_6;
  assign f_s_wallace_cla8_fa35_and1 = f_s_wallace_cla8_fa35_xor0 & f_s_wallace_cla8_nand_7_6;
  assign f_s_wallace_cla8_fa35_or0 = f_s_wallace_cla8_fa35_and0 | f_s_wallace_cla8_fa35_and1;
  assign f_s_wallace_cla8_and_0_0 = a[0] & b[0];
  assign f_s_wallace_cla8_and_1_0 = a[1] & b[0];
  assign f_s_wallace_cla8_and_0_2 = a[0] & b[2];
  assign f_s_wallace_cla8_nand_6_7 = ~(a[6] & b[7]);
  assign f_s_wallace_cla8_and_0_1 = a[0] & b[1];
  assign f_s_wallace_cla8_and_7_7 = a[7] & b[7];
  assign f_s_wallace_cla8_u_cla14_pg_logic0_or0 = f_s_wallace_cla8_and_1_0 | f_s_wallace_cla8_and_0_1;
  assign f_s_wallace_cla8_u_cla14_pg_logic0_and0 = f_s_wallace_cla8_and_1_0 & f_s_wallace_cla8_and_0_1;
  assign f_s_wallace_cla8_u_cla14_pg_logic0_xor0 = f_s_wallace_cla8_and_1_0 ^ f_s_wallace_cla8_and_0_1;
  assign f_s_wallace_cla8_u_cla14_pg_logic1_or0 = f_s_wallace_cla8_and_0_2 | f_s_wallace_cla8_ha0_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic1_and0 = f_s_wallace_cla8_and_0_2 & f_s_wallace_cla8_ha0_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic1_xor0 = f_s_wallace_cla8_and_0_2 ^ f_s_wallace_cla8_ha0_xor0;
  assign f_s_wallace_cla8_u_cla14_xor1 = f_s_wallace_cla8_u_cla14_pg_logic1_xor0 ^ f_s_wallace_cla8_u_cla14_pg_logic0_and0;
  assign f_s_wallace_cla8_u_cla14_and0 = f_s_wallace_cla8_u_cla14_pg_logic0_and0 & f_s_wallace_cla8_u_cla14_pg_logic1_or0;
  assign f_s_wallace_cla8_u_cla14_or0 = f_s_wallace_cla8_u_cla14_pg_logic1_and0 | f_s_wallace_cla8_u_cla14_and0;
  assign f_s_wallace_cla8_u_cla14_pg_logic2_or0 = f_s_wallace_cla8_fa0_xor1 | f_s_wallace_cla8_ha1_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic2_and0 = f_s_wallace_cla8_fa0_xor1 & f_s_wallace_cla8_ha1_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic2_xor0 = f_s_wallace_cla8_fa0_xor1 ^ f_s_wallace_cla8_ha1_xor0;
  assign f_s_wallace_cla8_u_cla14_xor2 = f_s_wallace_cla8_u_cla14_pg_logic2_xor0 ^ f_s_wallace_cla8_u_cla14_or0;
  assign f_s_wallace_cla8_u_cla14_and1 = f_s_wallace_cla8_u_cla14_pg_logic2_or0 & f_s_wallace_cla8_u_cla14_pg_logic0_or0;
  assign f_s_wallace_cla8_u_cla14_and2 = f_s_wallace_cla8_u_cla14_pg_logic0_and0 & f_s_wallace_cla8_u_cla14_pg_logic2_or0;
  assign f_s_wallace_cla8_u_cla14_and3 = f_s_wallace_cla8_u_cla14_and2 & f_s_wallace_cla8_u_cla14_pg_logic1_or0;
  assign f_s_wallace_cla8_u_cla14_and4 = f_s_wallace_cla8_u_cla14_pg_logic1_and0 & f_s_wallace_cla8_u_cla14_pg_logic2_or0;
  assign f_s_wallace_cla8_u_cla14_or1 = f_s_wallace_cla8_u_cla14_and3 | f_s_wallace_cla8_u_cla14_and4;
  assign f_s_wallace_cla8_u_cla14_or2 = f_s_wallace_cla8_u_cla14_pg_logic2_and0 | f_s_wallace_cla8_u_cla14_or1;
  assign f_s_wallace_cla8_u_cla14_pg_logic3_or0 = f_s_wallace_cla8_fa10_xor1 | f_s_wallace_cla8_ha2_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic3_and0 = f_s_wallace_cla8_fa10_xor1 & f_s_wallace_cla8_ha2_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic3_xor0 = f_s_wallace_cla8_fa10_xor1 ^ f_s_wallace_cla8_ha2_xor0;
  assign f_s_wallace_cla8_u_cla14_xor3 = f_s_wallace_cla8_u_cla14_pg_logic3_xor0 ^ f_s_wallace_cla8_u_cla14_or2;
  assign f_s_wallace_cla8_u_cla14_and5 = f_s_wallace_cla8_u_cla14_pg_logic3_or0 & f_s_wallace_cla8_u_cla14_pg_logic1_or0;
  assign f_s_wallace_cla8_u_cla14_and6 = f_s_wallace_cla8_u_cla14_pg_logic0_and0 & f_s_wallace_cla8_u_cla14_pg_logic2_or0;
  assign f_s_wallace_cla8_u_cla14_and7 = f_s_wallace_cla8_u_cla14_pg_logic3_or0 & f_s_wallace_cla8_u_cla14_pg_logic1_or0;
  assign f_s_wallace_cla8_u_cla14_and8 = f_s_wallace_cla8_u_cla14_and6 & f_s_wallace_cla8_u_cla14_and7;
  assign f_s_wallace_cla8_u_cla14_and9 = f_s_wallace_cla8_u_cla14_pg_logic1_and0 & f_s_wallace_cla8_u_cla14_pg_logic3_or0;
  assign f_s_wallace_cla8_u_cla14_and10 = f_s_wallace_cla8_u_cla14_and9 & f_s_wallace_cla8_u_cla14_pg_logic2_or0;
  assign f_s_wallace_cla8_u_cla14_and11 = f_s_wallace_cla8_u_cla14_pg_logic2_and0 & f_s_wallace_cla8_u_cla14_pg_logic3_or0;
  assign f_s_wallace_cla8_u_cla14_or3 = f_s_wallace_cla8_u_cla14_and8 | f_s_wallace_cla8_u_cla14_and11;
  assign f_s_wallace_cla8_u_cla14_or4 = f_s_wallace_cla8_u_cla14_and10 | f_s_wallace_cla8_u_cla14_or3;
  assign f_s_wallace_cla8_u_cla14_or5 = f_s_wallace_cla8_u_cla14_pg_logic3_and0 | f_s_wallace_cla8_u_cla14_or4;
  assign f_s_wallace_cla8_u_cla14_pg_logic4_or0 = f_s_wallace_cla8_fa18_xor1 | f_s_wallace_cla8_ha3_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic4_and0 = f_s_wallace_cla8_fa18_xor1 & f_s_wallace_cla8_ha3_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic4_xor0 = f_s_wallace_cla8_fa18_xor1 ^ f_s_wallace_cla8_ha3_xor0;
  assign f_s_wallace_cla8_u_cla14_xor4 = f_s_wallace_cla8_u_cla14_pg_logic4_xor0 ^ f_s_wallace_cla8_u_cla14_or5;
  assign f_s_wallace_cla8_u_cla14_and12 = f_s_wallace_cla8_u_cla14_or5 & f_s_wallace_cla8_u_cla14_pg_logic4_or0;
  assign f_s_wallace_cla8_u_cla14_or6 = f_s_wallace_cla8_u_cla14_pg_logic4_and0 | f_s_wallace_cla8_u_cla14_and12;
  assign f_s_wallace_cla8_u_cla14_pg_logic5_or0 = f_s_wallace_cla8_fa24_xor1 | f_s_wallace_cla8_ha4_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic5_and0 = f_s_wallace_cla8_fa24_xor1 & f_s_wallace_cla8_ha4_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic5_xor0 = f_s_wallace_cla8_fa24_xor1 ^ f_s_wallace_cla8_ha4_xor0;
  assign f_s_wallace_cla8_u_cla14_xor5 = f_s_wallace_cla8_u_cla14_pg_logic5_xor0 ^ f_s_wallace_cla8_u_cla14_or6;
  assign f_s_wallace_cla8_u_cla14_and13 = f_s_wallace_cla8_u_cla14_or5 & f_s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign f_s_wallace_cla8_u_cla14_and14 = f_s_wallace_cla8_u_cla14_and13 & f_s_wallace_cla8_u_cla14_pg_logic4_or0;
  assign f_s_wallace_cla8_u_cla14_and15 = f_s_wallace_cla8_u_cla14_pg_logic4_and0 & f_s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign f_s_wallace_cla8_u_cla14_or7 = f_s_wallace_cla8_u_cla14_and14 | f_s_wallace_cla8_u_cla14_and15;
  assign f_s_wallace_cla8_u_cla14_or8 = f_s_wallace_cla8_u_cla14_pg_logic5_and0 | f_s_wallace_cla8_u_cla14_or7;
  assign f_s_wallace_cla8_u_cla14_pg_logic6_or0 = f_s_wallace_cla8_fa28_xor1 | f_s_wallace_cla8_ha5_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic6_and0 = f_s_wallace_cla8_fa28_xor1 & f_s_wallace_cla8_ha5_xor0;
  assign f_s_wallace_cla8_u_cla14_pg_logic6_xor0 = f_s_wallace_cla8_fa28_xor1 ^ f_s_wallace_cla8_ha5_xor0;
  assign f_s_wallace_cla8_u_cla14_xor6 = f_s_wallace_cla8_u_cla14_pg_logic6_xor0 ^ f_s_wallace_cla8_u_cla14_or8;
  assign f_s_wallace_cla8_u_cla14_and16 = f_s_wallace_cla8_u_cla14_or5 & f_s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign f_s_wallace_cla8_u_cla14_and17 = f_s_wallace_cla8_u_cla14_pg_logic6_or0 & f_s_wallace_cla8_u_cla14_pg_logic4_or0;
  assign f_s_wallace_cla8_u_cla14_and18 = f_s_wallace_cla8_u_cla14_and16 & f_s_wallace_cla8_u_cla14_and17;
  assign f_s_wallace_cla8_u_cla14_and19 = f_s_wallace_cla8_u_cla14_pg_logic4_and0 & f_s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign f_s_wallace_cla8_u_cla14_and20 = f_s_wallace_cla8_u_cla14_and19 & f_s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign f_s_wallace_cla8_u_cla14_and21 = f_s_wallace_cla8_u_cla14_pg_logic5_and0 & f_s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign f_s_wallace_cla8_u_cla14_or9 = f_s_wallace_cla8_u_cla14_and18 | f_s_wallace_cla8_u_cla14_and20;
  assign f_s_wallace_cla8_u_cla14_or10 = f_s_wallace_cla8_u_cla14_or9 | f_s_wallace_cla8_u_cla14_and21;
  assign f_s_wallace_cla8_u_cla14_or11 = f_s_wallace_cla8_u_cla14_pg_logic6_and0 | f_s_wallace_cla8_u_cla14_or10;
  assign f_s_wallace_cla8_u_cla14_pg_logic7_or0 = f_s_wallace_cla8_fa29_xor1 | f_s_wallace_cla8_fa30_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic7_and0 = f_s_wallace_cla8_fa29_xor1 & f_s_wallace_cla8_fa30_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic7_xor0 = f_s_wallace_cla8_fa29_xor1 ^ f_s_wallace_cla8_fa30_xor1;
  assign f_s_wallace_cla8_u_cla14_xor7 = f_s_wallace_cla8_u_cla14_pg_logic7_xor0 ^ f_s_wallace_cla8_u_cla14_or11;
  assign f_s_wallace_cla8_u_cla14_and22 = f_s_wallace_cla8_u_cla14_or5 & f_s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign f_s_wallace_cla8_u_cla14_and23 = f_s_wallace_cla8_u_cla14_pg_logic7_or0 & f_s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign f_s_wallace_cla8_u_cla14_and24 = f_s_wallace_cla8_u_cla14_and22 & f_s_wallace_cla8_u_cla14_and23;
  assign f_s_wallace_cla8_u_cla14_and25 = f_s_wallace_cla8_u_cla14_and24 & f_s_wallace_cla8_u_cla14_pg_logic4_or0;
  assign f_s_wallace_cla8_u_cla14_and26 = f_s_wallace_cla8_u_cla14_pg_logic4_and0 & f_s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign f_s_wallace_cla8_u_cla14_and27 = f_s_wallace_cla8_u_cla14_pg_logic7_or0 & f_s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign f_s_wallace_cla8_u_cla14_and28 = f_s_wallace_cla8_u_cla14_and26 & f_s_wallace_cla8_u_cla14_and27;
  assign f_s_wallace_cla8_u_cla14_and29 = f_s_wallace_cla8_u_cla14_pg_logic5_and0 & f_s_wallace_cla8_u_cla14_pg_logic7_or0;
  assign f_s_wallace_cla8_u_cla14_and30 = f_s_wallace_cla8_u_cla14_and29 & f_s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign f_s_wallace_cla8_u_cla14_and31 = f_s_wallace_cla8_u_cla14_pg_logic6_and0 & f_s_wallace_cla8_u_cla14_pg_logic7_or0;
  assign f_s_wallace_cla8_u_cla14_or12 = f_s_wallace_cla8_u_cla14_and25 | f_s_wallace_cla8_u_cla14_and30;
  assign f_s_wallace_cla8_u_cla14_or13 = f_s_wallace_cla8_u_cla14_and28 | f_s_wallace_cla8_u_cla14_and31;
  assign f_s_wallace_cla8_u_cla14_or14 = f_s_wallace_cla8_u_cla14_or12 | f_s_wallace_cla8_u_cla14_or13;
  assign f_s_wallace_cla8_u_cla14_or15 = f_s_wallace_cla8_u_cla14_pg_logic7_and0 | f_s_wallace_cla8_u_cla14_or14;
  assign f_s_wallace_cla8_u_cla14_pg_logic8_or0 = f_s_wallace_cla8_fa27_xor1 | f_s_wallace_cla8_fa31_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic8_and0 = f_s_wallace_cla8_fa27_xor1 & f_s_wallace_cla8_fa31_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic8_xor0 = f_s_wallace_cla8_fa27_xor1 ^ f_s_wallace_cla8_fa31_xor1;
  assign f_s_wallace_cla8_u_cla14_xor8 = f_s_wallace_cla8_u_cla14_pg_logic8_xor0 ^ f_s_wallace_cla8_u_cla14_or15;
  assign f_s_wallace_cla8_u_cla14_and32 = f_s_wallace_cla8_u_cla14_or15 & f_s_wallace_cla8_u_cla14_pg_logic8_or0;
  assign f_s_wallace_cla8_u_cla14_or16 = f_s_wallace_cla8_u_cla14_pg_logic8_and0 | f_s_wallace_cla8_u_cla14_and32;
  assign f_s_wallace_cla8_u_cla14_pg_logic9_or0 = f_s_wallace_cla8_fa23_xor1 | f_s_wallace_cla8_fa32_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic9_and0 = f_s_wallace_cla8_fa23_xor1 & f_s_wallace_cla8_fa32_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic9_xor0 = f_s_wallace_cla8_fa23_xor1 ^ f_s_wallace_cla8_fa32_xor1;
  assign f_s_wallace_cla8_u_cla14_xor9 = f_s_wallace_cla8_u_cla14_pg_logic9_xor0 ^ f_s_wallace_cla8_u_cla14_or16;
  assign f_s_wallace_cla8_u_cla14_and33 = f_s_wallace_cla8_u_cla14_or15 & f_s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign f_s_wallace_cla8_u_cla14_and34 = f_s_wallace_cla8_u_cla14_and33 & f_s_wallace_cla8_u_cla14_pg_logic8_or0;
  assign f_s_wallace_cla8_u_cla14_and35 = f_s_wallace_cla8_u_cla14_pg_logic8_and0 & f_s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign f_s_wallace_cla8_u_cla14_or17 = f_s_wallace_cla8_u_cla14_and34 | f_s_wallace_cla8_u_cla14_and35;
  assign f_s_wallace_cla8_u_cla14_or18 = f_s_wallace_cla8_u_cla14_pg_logic9_and0 | f_s_wallace_cla8_u_cla14_or17;
  assign f_s_wallace_cla8_u_cla14_pg_logic10_or0 = f_s_wallace_cla8_fa17_xor1 | f_s_wallace_cla8_fa33_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic10_and0 = f_s_wallace_cla8_fa17_xor1 & f_s_wallace_cla8_fa33_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic10_xor0 = f_s_wallace_cla8_fa17_xor1 ^ f_s_wallace_cla8_fa33_xor1;
  assign f_s_wallace_cla8_u_cla14_xor10 = f_s_wallace_cla8_u_cla14_pg_logic10_xor0 ^ f_s_wallace_cla8_u_cla14_or18;
  assign f_s_wallace_cla8_u_cla14_and36 = f_s_wallace_cla8_u_cla14_or15 & f_s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign f_s_wallace_cla8_u_cla14_and37 = f_s_wallace_cla8_u_cla14_pg_logic10_or0 & f_s_wallace_cla8_u_cla14_pg_logic8_or0;
  assign f_s_wallace_cla8_u_cla14_and38 = f_s_wallace_cla8_u_cla14_and36 & f_s_wallace_cla8_u_cla14_and37;
  assign f_s_wallace_cla8_u_cla14_and39 = f_s_wallace_cla8_u_cla14_pg_logic8_and0 & f_s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign f_s_wallace_cla8_u_cla14_and40 = f_s_wallace_cla8_u_cla14_and39 & f_s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign f_s_wallace_cla8_u_cla14_and41 = f_s_wallace_cla8_u_cla14_pg_logic9_and0 & f_s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign f_s_wallace_cla8_u_cla14_or19 = f_s_wallace_cla8_u_cla14_and38 | f_s_wallace_cla8_u_cla14_and40;
  assign f_s_wallace_cla8_u_cla14_or20 = f_s_wallace_cla8_u_cla14_or19 | f_s_wallace_cla8_u_cla14_and41;
  assign f_s_wallace_cla8_u_cla14_or21 = f_s_wallace_cla8_u_cla14_pg_logic10_and0 | f_s_wallace_cla8_u_cla14_or20;
  assign f_s_wallace_cla8_u_cla14_pg_logic11_or0 = f_s_wallace_cla8_fa9_xor1 | f_s_wallace_cla8_fa34_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic11_and0 = f_s_wallace_cla8_fa9_xor1 & f_s_wallace_cla8_fa34_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic11_xor0 = f_s_wallace_cla8_fa9_xor1 ^ f_s_wallace_cla8_fa34_xor1;
  assign f_s_wallace_cla8_u_cla14_xor11 = f_s_wallace_cla8_u_cla14_pg_logic11_xor0 ^ f_s_wallace_cla8_u_cla14_or21;
  assign f_s_wallace_cla8_u_cla14_and42 = f_s_wallace_cla8_u_cla14_or15 & f_s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign f_s_wallace_cla8_u_cla14_and43 = f_s_wallace_cla8_u_cla14_pg_logic11_or0 & f_s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign f_s_wallace_cla8_u_cla14_and44 = f_s_wallace_cla8_u_cla14_and42 & f_s_wallace_cla8_u_cla14_and43;
  assign f_s_wallace_cla8_u_cla14_and45 = f_s_wallace_cla8_u_cla14_and44 & f_s_wallace_cla8_u_cla14_pg_logic8_or0;
  assign f_s_wallace_cla8_u_cla14_and46 = f_s_wallace_cla8_u_cla14_pg_logic8_and0 & f_s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign f_s_wallace_cla8_u_cla14_and47 = f_s_wallace_cla8_u_cla14_pg_logic11_or0 & f_s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign f_s_wallace_cla8_u_cla14_and48 = f_s_wallace_cla8_u_cla14_and46 & f_s_wallace_cla8_u_cla14_and47;
  assign f_s_wallace_cla8_u_cla14_and49 = f_s_wallace_cla8_u_cla14_pg_logic9_and0 & f_s_wallace_cla8_u_cla14_pg_logic11_or0;
  assign f_s_wallace_cla8_u_cla14_and50 = f_s_wallace_cla8_u_cla14_and49 & f_s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign f_s_wallace_cla8_u_cla14_and51 = f_s_wallace_cla8_u_cla14_pg_logic10_and0 & f_s_wallace_cla8_u_cla14_pg_logic11_or0;
  assign f_s_wallace_cla8_u_cla14_or22 = f_s_wallace_cla8_u_cla14_and45 | f_s_wallace_cla8_u_cla14_and50;
  assign f_s_wallace_cla8_u_cla14_or23 = f_s_wallace_cla8_u_cla14_and48 | f_s_wallace_cla8_u_cla14_and51;
  assign f_s_wallace_cla8_u_cla14_or24 = f_s_wallace_cla8_u_cla14_or22 | f_s_wallace_cla8_u_cla14_or23;
  assign f_s_wallace_cla8_u_cla14_or25 = f_s_wallace_cla8_u_cla14_pg_logic11_and0 | f_s_wallace_cla8_u_cla14_or24;
  assign f_s_wallace_cla8_u_cla14_pg_logic12_or0 = f_s_wallace_cla8_nand_6_7 | f_s_wallace_cla8_fa35_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic12_and0 = f_s_wallace_cla8_nand_6_7 & f_s_wallace_cla8_fa35_xor1;
  assign f_s_wallace_cla8_u_cla14_pg_logic12_xor0 = f_s_wallace_cla8_nand_6_7 ^ f_s_wallace_cla8_fa35_xor1;
  assign f_s_wallace_cla8_u_cla14_xor12 = f_s_wallace_cla8_u_cla14_pg_logic12_xor0 ^ f_s_wallace_cla8_u_cla14_or25;
  assign f_s_wallace_cla8_u_cla14_and52 = f_s_wallace_cla8_u_cla14_or25 & f_s_wallace_cla8_u_cla14_pg_logic12_or0;
  assign f_s_wallace_cla8_u_cla14_or26 = f_s_wallace_cla8_u_cla14_pg_logic12_and0 | f_s_wallace_cla8_u_cla14_and52;
  assign f_s_wallace_cla8_u_cla14_pg_logic13_or0 = f_s_wallace_cla8_fa35_or0 | f_s_wallace_cla8_and_7_7;
  assign f_s_wallace_cla8_u_cla14_pg_logic13_and0 = f_s_wallace_cla8_fa35_or0 & f_s_wallace_cla8_and_7_7;
  assign f_s_wallace_cla8_u_cla14_pg_logic13_xor0 = f_s_wallace_cla8_fa35_or0 ^ f_s_wallace_cla8_and_7_7;
  assign f_s_wallace_cla8_u_cla14_xor13 = f_s_wallace_cla8_u_cla14_pg_logic13_xor0 ^ f_s_wallace_cla8_u_cla14_or26;
  assign f_s_wallace_cla8_u_cla14_and53 = f_s_wallace_cla8_u_cla14_or25 & f_s_wallace_cla8_u_cla14_pg_logic13_or0;
  assign f_s_wallace_cla8_u_cla14_and54 = f_s_wallace_cla8_u_cla14_and53 & f_s_wallace_cla8_u_cla14_pg_logic12_or0;
  assign f_s_wallace_cla8_u_cla14_and55 = f_s_wallace_cla8_u_cla14_pg_logic12_and0 & f_s_wallace_cla8_u_cla14_pg_logic13_or0;
  assign f_s_wallace_cla8_u_cla14_or27 = f_s_wallace_cla8_u_cla14_and54 | f_s_wallace_cla8_u_cla14_and55;
  assign f_s_wallace_cla8_u_cla14_or28 = f_s_wallace_cla8_u_cla14_pg_logic13_and0 | f_s_wallace_cla8_u_cla14_or27;
  assign f_s_wallace_cla8_xor0 = ~f_s_wallace_cla8_u_cla14_or28;

  assign f_s_wallace_cla8_out[0] = f_s_wallace_cla8_and_0_0;
  assign f_s_wallace_cla8_out[1] = f_s_wallace_cla8_u_cla14_pg_logic0_xor0;
  assign f_s_wallace_cla8_out[2] = f_s_wallace_cla8_u_cla14_xor1;
  assign f_s_wallace_cla8_out[3] = f_s_wallace_cla8_u_cla14_xor2;
  assign f_s_wallace_cla8_out[4] = f_s_wallace_cla8_u_cla14_xor3;
  assign f_s_wallace_cla8_out[5] = f_s_wallace_cla8_u_cla14_xor4;
  assign f_s_wallace_cla8_out[6] = f_s_wallace_cla8_u_cla14_xor5;
  assign f_s_wallace_cla8_out[7] = f_s_wallace_cla8_u_cla14_xor6;
  assign f_s_wallace_cla8_out[8] = f_s_wallace_cla8_u_cla14_xor7;
  assign f_s_wallace_cla8_out[9] = f_s_wallace_cla8_u_cla14_xor8;
  assign f_s_wallace_cla8_out[10] = f_s_wallace_cla8_u_cla14_xor9;
  assign f_s_wallace_cla8_out[11] = f_s_wallace_cla8_u_cla14_xor10;
  assign f_s_wallace_cla8_out[12] = f_s_wallace_cla8_u_cla14_xor11;
  assign f_s_wallace_cla8_out[13] = f_s_wallace_cla8_u_cla14_xor12;
  assign f_s_wallace_cla8_out[14] = f_s_wallace_cla8_u_cla14_xor13;
  assign f_s_wallace_cla8_out[15] = f_s_wallace_cla8_xor0;
endmodule