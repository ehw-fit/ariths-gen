module u_CSAwallace_cska32(input [31:0] a, input [31:0] b, output [63:0] u_CSAwallace_cska32_out);
  wire u_CSAwallace_cska32_and_0_0;
  wire u_CSAwallace_cska32_and_1_0;
  wire u_CSAwallace_cska32_and_2_0;
  wire u_CSAwallace_cska32_and_3_0;
  wire u_CSAwallace_cska32_and_4_0;
  wire u_CSAwallace_cska32_and_5_0;
  wire u_CSAwallace_cska32_and_6_0;
  wire u_CSAwallace_cska32_and_7_0;
  wire u_CSAwallace_cska32_and_8_0;
  wire u_CSAwallace_cska32_and_9_0;
  wire u_CSAwallace_cska32_and_10_0;
  wire u_CSAwallace_cska32_and_11_0;
  wire u_CSAwallace_cska32_and_12_0;
  wire u_CSAwallace_cska32_and_13_0;
  wire u_CSAwallace_cska32_and_14_0;
  wire u_CSAwallace_cska32_and_15_0;
  wire u_CSAwallace_cska32_and_16_0;
  wire u_CSAwallace_cska32_and_17_0;
  wire u_CSAwallace_cska32_and_18_0;
  wire u_CSAwallace_cska32_and_19_0;
  wire u_CSAwallace_cska32_and_20_0;
  wire u_CSAwallace_cska32_and_21_0;
  wire u_CSAwallace_cska32_and_22_0;
  wire u_CSAwallace_cska32_and_23_0;
  wire u_CSAwallace_cska32_and_24_0;
  wire u_CSAwallace_cska32_and_25_0;
  wire u_CSAwallace_cska32_and_26_0;
  wire u_CSAwallace_cska32_and_27_0;
  wire u_CSAwallace_cska32_and_28_0;
  wire u_CSAwallace_cska32_and_29_0;
  wire u_CSAwallace_cska32_and_30_0;
  wire u_CSAwallace_cska32_and_31_0;
  wire u_CSAwallace_cska32_and_0_1;
  wire u_CSAwallace_cska32_and_1_1;
  wire u_CSAwallace_cska32_and_2_1;
  wire u_CSAwallace_cska32_and_3_1;
  wire u_CSAwallace_cska32_and_4_1;
  wire u_CSAwallace_cska32_and_5_1;
  wire u_CSAwallace_cska32_and_6_1;
  wire u_CSAwallace_cska32_and_7_1;
  wire u_CSAwallace_cska32_and_8_1;
  wire u_CSAwallace_cska32_and_9_1;
  wire u_CSAwallace_cska32_and_10_1;
  wire u_CSAwallace_cska32_and_11_1;
  wire u_CSAwallace_cska32_and_12_1;
  wire u_CSAwallace_cska32_and_13_1;
  wire u_CSAwallace_cska32_and_14_1;
  wire u_CSAwallace_cska32_and_15_1;
  wire u_CSAwallace_cska32_and_16_1;
  wire u_CSAwallace_cska32_and_17_1;
  wire u_CSAwallace_cska32_and_18_1;
  wire u_CSAwallace_cska32_and_19_1;
  wire u_CSAwallace_cska32_and_20_1;
  wire u_CSAwallace_cska32_and_21_1;
  wire u_CSAwallace_cska32_and_22_1;
  wire u_CSAwallace_cska32_and_23_1;
  wire u_CSAwallace_cska32_and_24_1;
  wire u_CSAwallace_cska32_and_25_1;
  wire u_CSAwallace_cska32_and_26_1;
  wire u_CSAwallace_cska32_and_27_1;
  wire u_CSAwallace_cska32_and_28_1;
  wire u_CSAwallace_cska32_and_29_1;
  wire u_CSAwallace_cska32_and_30_1;
  wire u_CSAwallace_cska32_and_31_1;
  wire u_CSAwallace_cska32_and_0_2;
  wire u_CSAwallace_cska32_and_1_2;
  wire u_CSAwallace_cska32_and_2_2;
  wire u_CSAwallace_cska32_and_3_2;
  wire u_CSAwallace_cska32_and_4_2;
  wire u_CSAwallace_cska32_and_5_2;
  wire u_CSAwallace_cska32_and_6_2;
  wire u_CSAwallace_cska32_and_7_2;
  wire u_CSAwallace_cska32_and_8_2;
  wire u_CSAwallace_cska32_and_9_2;
  wire u_CSAwallace_cska32_and_10_2;
  wire u_CSAwallace_cska32_and_11_2;
  wire u_CSAwallace_cska32_and_12_2;
  wire u_CSAwallace_cska32_and_13_2;
  wire u_CSAwallace_cska32_and_14_2;
  wire u_CSAwallace_cska32_and_15_2;
  wire u_CSAwallace_cska32_and_16_2;
  wire u_CSAwallace_cska32_and_17_2;
  wire u_CSAwallace_cska32_and_18_2;
  wire u_CSAwallace_cska32_and_19_2;
  wire u_CSAwallace_cska32_and_20_2;
  wire u_CSAwallace_cska32_and_21_2;
  wire u_CSAwallace_cska32_and_22_2;
  wire u_CSAwallace_cska32_and_23_2;
  wire u_CSAwallace_cska32_and_24_2;
  wire u_CSAwallace_cska32_and_25_2;
  wire u_CSAwallace_cska32_and_26_2;
  wire u_CSAwallace_cska32_and_27_2;
  wire u_CSAwallace_cska32_and_28_2;
  wire u_CSAwallace_cska32_and_29_2;
  wire u_CSAwallace_cska32_and_30_2;
  wire u_CSAwallace_cska32_and_31_2;
  wire u_CSAwallace_cska32_and_0_3;
  wire u_CSAwallace_cska32_and_1_3;
  wire u_CSAwallace_cska32_and_2_3;
  wire u_CSAwallace_cska32_and_3_3;
  wire u_CSAwallace_cska32_and_4_3;
  wire u_CSAwallace_cska32_and_5_3;
  wire u_CSAwallace_cska32_and_6_3;
  wire u_CSAwallace_cska32_and_7_3;
  wire u_CSAwallace_cska32_and_8_3;
  wire u_CSAwallace_cska32_and_9_3;
  wire u_CSAwallace_cska32_and_10_3;
  wire u_CSAwallace_cska32_and_11_3;
  wire u_CSAwallace_cska32_and_12_3;
  wire u_CSAwallace_cska32_and_13_3;
  wire u_CSAwallace_cska32_and_14_3;
  wire u_CSAwallace_cska32_and_15_3;
  wire u_CSAwallace_cska32_and_16_3;
  wire u_CSAwallace_cska32_and_17_3;
  wire u_CSAwallace_cska32_and_18_3;
  wire u_CSAwallace_cska32_and_19_3;
  wire u_CSAwallace_cska32_and_20_3;
  wire u_CSAwallace_cska32_and_21_3;
  wire u_CSAwallace_cska32_and_22_3;
  wire u_CSAwallace_cska32_and_23_3;
  wire u_CSAwallace_cska32_and_24_3;
  wire u_CSAwallace_cska32_and_25_3;
  wire u_CSAwallace_cska32_and_26_3;
  wire u_CSAwallace_cska32_and_27_3;
  wire u_CSAwallace_cska32_and_28_3;
  wire u_CSAwallace_cska32_and_29_3;
  wire u_CSAwallace_cska32_and_30_3;
  wire u_CSAwallace_cska32_and_31_3;
  wire u_CSAwallace_cska32_and_0_4;
  wire u_CSAwallace_cska32_and_1_4;
  wire u_CSAwallace_cska32_and_2_4;
  wire u_CSAwallace_cska32_and_3_4;
  wire u_CSAwallace_cska32_and_4_4;
  wire u_CSAwallace_cska32_and_5_4;
  wire u_CSAwallace_cska32_and_6_4;
  wire u_CSAwallace_cska32_and_7_4;
  wire u_CSAwallace_cska32_and_8_4;
  wire u_CSAwallace_cska32_and_9_4;
  wire u_CSAwallace_cska32_and_10_4;
  wire u_CSAwallace_cska32_and_11_4;
  wire u_CSAwallace_cska32_and_12_4;
  wire u_CSAwallace_cska32_and_13_4;
  wire u_CSAwallace_cska32_and_14_4;
  wire u_CSAwallace_cska32_and_15_4;
  wire u_CSAwallace_cska32_and_16_4;
  wire u_CSAwallace_cska32_and_17_4;
  wire u_CSAwallace_cska32_and_18_4;
  wire u_CSAwallace_cska32_and_19_4;
  wire u_CSAwallace_cska32_and_20_4;
  wire u_CSAwallace_cska32_and_21_4;
  wire u_CSAwallace_cska32_and_22_4;
  wire u_CSAwallace_cska32_and_23_4;
  wire u_CSAwallace_cska32_and_24_4;
  wire u_CSAwallace_cska32_and_25_4;
  wire u_CSAwallace_cska32_and_26_4;
  wire u_CSAwallace_cska32_and_27_4;
  wire u_CSAwallace_cska32_and_28_4;
  wire u_CSAwallace_cska32_and_29_4;
  wire u_CSAwallace_cska32_and_30_4;
  wire u_CSAwallace_cska32_and_31_4;
  wire u_CSAwallace_cska32_and_0_5;
  wire u_CSAwallace_cska32_and_1_5;
  wire u_CSAwallace_cska32_and_2_5;
  wire u_CSAwallace_cska32_and_3_5;
  wire u_CSAwallace_cska32_and_4_5;
  wire u_CSAwallace_cska32_and_5_5;
  wire u_CSAwallace_cska32_and_6_5;
  wire u_CSAwallace_cska32_and_7_5;
  wire u_CSAwallace_cska32_and_8_5;
  wire u_CSAwallace_cska32_and_9_5;
  wire u_CSAwallace_cska32_and_10_5;
  wire u_CSAwallace_cska32_and_11_5;
  wire u_CSAwallace_cska32_and_12_5;
  wire u_CSAwallace_cska32_and_13_5;
  wire u_CSAwallace_cska32_and_14_5;
  wire u_CSAwallace_cska32_and_15_5;
  wire u_CSAwallace_cska32_and_16_5;
  wire u_CSAwallace_cska32_and_17_5;
  wire u_CSAwallace_cska32_and_18_5;
  wire u_CSAwallace_cska32_and_19_5;
  wire u_CSAwallace_cska32_and_20_5;
  wire u_CSAwallace_cska32_and_21_5;
  wire u_CSAwallace_cska32_and_22_5;
  wire u_CSAwallace_cska32_and_23_5;
  wire u_CSAwallace_cska32_and_24_5;
  wire u_CSAwallace_cska32_and_25_5;
  wire u_CSAwallace_cska32_and_26_5;
  wire u_CSAwallace_cska32_and_27_5;
  wire u_CSAwallace_cska32_and_28_5;
  wire u_CSAwallace_cska32_and_29_5;
  wire u_CSAwallace_cska32_and_30_5;
  wire u_CSAwallace_cska32_and_31_5;
  wire u_CSAwallace_cska32_and_0_6;
  wire u_CSAwallace_cska32_and_1_6;
  wire u_CSAwallace_cska32_and_2_6;
  wire u_CSAwallace_cska32_and_3_6;
  wire u_CSAwallace_cska32_and_4_6;
  wire u_CSAwallace_cska32_and_5_6;
  wire u_CSAwallace_cska32_and_6_6;
  wire u_CSAwallace_cska32_and_7_6;
  wire u_CSAwallace_cska32_and_8_6;
  wire u_CSAwallace_cska32_and_9_6;
  wire u_CSAwallace_cska32_and_10_6;
  wire u_CSAwallace_cska32_and_11_6;
  wire u_CSAwallace_cska32_and_12_6;
  wire u_CSAwallace_cska32_and_13_6;
  wire u_CSAwallace_cska32_and_14_6;
  wire u_CSAwallace_cska32_and_15_6;
  wire u_CSAwallace_cska32_and_16_6;
  wire u_CSAwallace_cska32_and_17_6;
  wire u_CSAwallace_cska32_and_18_6;
  wire u_CSAwallace_cska32_and_19_6;
  wire u_CSAwallace_cska32_and_20_6;
  wire u_CSAwallace_cska32_and_21_6;
  wire u_CSAwallace_cska32_and_22_6;
  wire u_CSAwallace_cska32_and_23_6;
  wire u_CSAwallace_cska32_and_24_6;
  wire u_CSAwallace_cska32_and_25_6;
  wire u_CSAwallace_cska32_and_26_6;
  wire u_CSAwallace_cska32_and_27_6;
  wire u_CSAwallace_cska32_and_28_6;
  wire u_CSAwallace_cska32_and_29_6;
  wire u_CSAwallace_cska32_and_30_6;
  wire u_CSAwallace_cska32_and_31_6;
  wire u_CSAwallace_cska32_and_0_7;
  wire u_CSAwallace_cska32_and_1_7;
  wire u_CSAwallace_cska32_and_2_7;
  wire u_CSAwallace_cska32_and_3_7;
  wire u_CSAwallace_cska32_and_4_7;
  wire u_CSAwallace_cska32_and_5_7;
  wire u_CSAwallace_cska32_and_6_7;
  wire u_CSAwallace_cska32_and_7_7;
  wire u_CSAwallace_cska32_and_8_7;
  wire u_CSAwallace_cska32_and_9_7;
  wire u_CSAwallace_cska32_and_10_7;
  wire u_CSAwallace_cska32_and_11_7;
  wire u_CSAwallace_cska32_and_12_7;
  wire u_CSAwallace_cska32_and_13_7;
  wire u_CSAwallace_cska32_and_14_7;
  wire u_CSAwallace_cska32_and_15_7;
  wire u_CSAwallace_cska32_and_16_7;
  wire u_CSAwallace_cska32_and_17_7;
  wire u_CSAwallace_cska32_and_18_7;
  wire u_CSAwallace_cska32_and_19_7;
  wire u_CSAwallace_cska32_and_20_7;
  wire u_CSAwallace_cska32_and_21_7;
  wire u_CSAwallace_cska32_and_22_7;
  wire u_CSAwallace_cska32_and_23_7;
  wire u_CSAwallace_cska32_and_24_7;
  wire u_CSAwallace_cska32_and_25_7;
  wire u_CSAwallace_cska32_and_26_7;
  wire u_CSAwallace_cska32_and_27_7;
  wire u_CSAwallace_cska32_and_28_7;
  wire u_CSAwallace_cska32_and_29_7;
  wire u_CSAwallace_cska32_and_30_7;
  wire u_CSAwallace_cska32_and_31_7;
  wire u_CSAwallace_cska32_and_0_8;
  wire u_CSAwallace_cska32_and_1_8;
  wire u_CSAwallace_cska32_and_2_8;
  wire u_CSAwallace_cska32_and_3_8;
  wire u_CSAwallace_cska32_and_4_8;
  wire u_CSAwallace_cska32_and_5_8;
  wire u_CSAwallace_cska32_and_6_8;
  wire u_CSAwallace_cska32_and_7_8;
  wire u_CSAwallace_cska32_and_8_8;
  wire u_CSAwallace_cska32_and_9_8;
  wire u_CSAwallace_cska32_and_10_8;
  wire u_CSAwallace_cska32_and_11_8;
  wire u_CSAwallace_cska32_and_12_8;
  wire u_CSAwallace_cska32_and_13_8;
  wire u_CSAwallace_cska32_and_14_8;
  wire u_CSAwallace_cska32_and_15_8;
  wire u_CSAwallace_cska32_and_16_8;
  wire u_CSAwallace_cska32_and_17_8;
  wire u_CSAwallace_cska32_and_18_8;
  wire u_CSAwallace_cska32_and_19_8;
  wire u_CSAwallace_cska32_and_20_8;
  wire u_CSAwallace_cska32_and_21_8;
  wire u_CSAwallace_cska32_and_22_8;
  wire u_CSAwallace_cska32_and_23_8;
  wire u_CSAwallace_cska32_and_24_8;
  wire u_CSAwallace_cska32_and_25_8;
  wire u_CSAwallace_cska32_and_26_8;
  wire u_CSAwallace_cska32_and_27_8;
  wire u_CSAwallace_cska32_and_28_8;
  wire u_CSAwallace_cska32_and_29_8;
  wire u_CSAwallace_cska32_and_30_8;
  wire u_CSAwallace_cska32_and_31_8;
  wire u_CSAwallace_cska32_and_0_9;
  wire u_CSAwallace_cska32_and_1_9;
  wire u_CSAwallace_cska32_and_2_9;
  wire u_CSAwallace_cska32_and_3_9;
  wire u_CSAwallace_cska32_and_4_9;
  wire u_CSAwallace_cska32_and_5_9;
  wire u_CSAwallace_cska32_and_6_9;
  wire u_CSAwallace_cska32_and_7_9;
  wire u_CSAwallace_cska32_and_8_9;
  wire u_CSAwallace_cska32_and_9_9;
  wire u_CSAwallace_cska32_and_10_9;
  wire u_CSAwallace_cska32_and_11_9;
  wire u_CSAwallace_cska32_and_12_9;
  wire u_CSAwallace_cska32_and_13_9;
  wire u_CSAwallace_cska32_and_14_9;
  wire u_CSAwallace_cska32_and_15_9;
  wire u_CSAwallace_cska32_and_16_9;
  wire u_CSAwallace_cska32_and_17_9;
  wire u_CSAwallace_cska32_and_18_9;
  wire u_CSAwallace_cska32_and_19_9;
  wire u_CSAwallace_cska32_and_20_9;
  wire u_CSAwallace_cska32_and_21_9;
  wire u_CSAwallace_cska32_and_22_9;
  wire u_CSAwallace_cska32_and_23_9;
  wire u_CSAwallace_cska32_and_24_9;
  wire u_CSAwallace_cska32_and_25_9;
  wire u_CSAwallace_cska32_and_26_9;
  wire u_CSAwallace_cska32_and_27_9;
  wire u_CSAwallace_cska32_and_28_9;
  wire u_CSAwallace_cska32_and_29_9;
  wire u_CSAwallace_cska32_and_30_9;
  wire u_CSAwallace_cska32_and_31_9;
  wire u_CSAwallace_cska32_and_0_10;
  wire u_CSAwallace_cska32_and_1_10;
  wire u_CSAwallace_cska32_and_2_10;
  wire u_CSAwallace_cska32_and_3_10;
  wire u_CSAwallace_cska32_and_4_10;
  wire u_CSAwallace_cska32_and_5_10;
  wire u_CSAwallace_cska32_and_6_10;
  wire u_CSAwallace_cska32_and_7_10;
  wire u_CSAwallace_cska32_and_8_10;
  wire u_CSAwallace_cska32_and_9_10;
  wire u_CSAwallace_cska32_and_10_10;
  wire u_CSAwallace_cska32_and_11_10;
  wire u_CSAwallace_cska32_and_12_10;
  wire u_CSAwallace_cska32_and_13_10;
  wire u_CSAwallace_cska32_and_14_10;
  wire u_CSAwallace_cska32_and_15_10;
  wire u_CSAwallace_cska32_and_16_10;
  wire u_CSAwallace_cska32_and_17_10;
  wire u_CSAwallace_cska32_and_18_10;
  wire u_CSAwallace_cska32_and_19_10;
  wire u_CSAwallace_cska32_and_20_10;
  wire u_CSAwallace_cska32_and_21_10;
  wire u_CSAwallace_cska32_and_22_10;
  wire u_CSAwallace_cska32_and_23_10;
  wire u_CSAwallace_cska32_and_24_10;
  wire u_CSAwallace_cska32_and_25_10;
  wire u_CSAwallace_cska32_and_26_10;
  wire u_CSAwallace_cska32_and_27_10;
  wire u_CSAwallace_cska32_and_28_10;
  wire u_CSAwallace_cska32_and_29_10;
  wire u_CSAwallace_cska32_and_30_10;
  wire u_CSAwallace_cska32_and_31_10;
  wire u_CSAwallace_cska32_and_0_11;
  wire u_CSAwallace_cska32_and_1_11;
  wire u_CSAwallace_cska32_and_2_11;
  wire u_CSAwallace_cska32_and_3_11;
  wire u_CSAwallace_cska32_and_4_11;
  wire u_CSAwallace_cska32_and_5_11;
  wire u_CSAwallace_cska32_and_6_11;
  wire u_CSAwallace_cska32_and_7_11;
  wire u_CSAwallace_cska32_and_8_11;
  wire u_CSAwallace_cska32_and_9_11;
  wire u_CSAwallace_cska32_and_10_11;
  wire u_CSAwallace_cska32_and_11_11;
  wire u_CSAwallace_cska32_and_12_11;
  wire u_CSAwallace_cska32_and_13_11;
  wire u_CSAwallace_cska32_and_14_11;
  wire u_CSAwallace_cska32_and_15_11;
  wire u_CSAwallace_cska32_and_16_11;
  wire u_CSAwallace_cska32_and_17_11;
  wire u_CSAwallace_cska32_and_18_11;
  wire u_CSAwallace_cska32_and_19_11;
  wire u_CSAwallace_cska32_and_20_11;
  wire u_CSAwallace_cska32_and_21_11;
  wire u_CSAwallace_cska32_and_22_11;
  wire u_CSAwallace_cska32_and_23_11;
  wire u_CSAwallace_cska32_and_24_11;
  wire u_CSAwallace_cska32_and_25_11;
  wire u_CSAwallace_cska32_and_26_11;
  wire u_CSAwallace_cska32_and_27_11;
  wire u_CSAwallace_cska32_and_28_11;
  wire u_CSAwallace_cska32_and_29_11;
  wire u_CSAwallace_cska32_and_30_11;
  wire u_CSAwallace_cska32_and_31_11;
  wire u_CSAwallace_cska32_and_0_12;
  wire u_CSAwallace_cska32_and_1_12;
  wire u_CSAwallace_cska32_and_2_12;
  wire u_CSAwallace_cska32_and_3_12;
  wire u_CSAwallace_cska32_and_4_12;
  wire u_CSAwallace_cska32_and_5_12;
  wire u_CSAwallace_cska32_and_6_12;
  wire u_CSAwallace_cska32_and_7_12;
  wire u_CSAwallace_cska32_and_8_12;
  wire u_CSAwallace_cska32_and_9_12;
  wire u_CSAwallace_cska32_and_10_12;
  wire u_CSAwallace_cska32_and_11_12;
  wire u_CSAwallace_cska32_and_12_12;
  wire u_CSAwallace_cska32_and_13_12;
  wire u_CSAwallace_cska32_and_14_12;
  wire u_CSAwallace_cska32_and_15_12;
  wire u_CSAwallace_cska32_and_16_12;
  wire u_CSAwallace_cska32_and_17_12;
  wire u_CSAwallace_cska32_and_18_12;
  wire u_CSAwallace_cska32_and_19_12;
  wire u_CSAwallace_cska32_and_20_12;
  wire u_CSAwallace_cska32_and_21_12;
  wire u_CSAwallace_cska32_and_22_12;
  wire u_CSAwallace_cska32_and_23_12;
  wire u_CSAwallace_cska32_and_24_12;
  wire u_CSAwallace_cska32_and_25_12;
  wire u_CSAwallace_cska32_and_26_12;
  wire u_CSAwallace_cska32_and_27_12;
  wire u_CSAwallace_cska32_and_28_12;
  wire u_CSAwallace_cska32_and_29_12;
  wire u_CSAwallace_cska32_and_30_12;
  wire u_CSAwallace_cska32_and_31_12;
  wire u_CSAwallace_cska32_and_0_13;
  wire u_CSAwallace_cska32_and_1_13;
  wire u_CSAwallace_cska32_and_2_13;
  wire u_CSAwallace_cska32_and_3_13;
  wire u_CSAwallace_cska32_and_4_13;
  wire u_CSAwallace_cska32_and_5_13;
  wire u_CSAwallace_cska32_and_6_13;
  wire u_CSAwallace_cska32_and_7_13;
  wire u_CSAwallace_cska32_and_8_13;
  wire u_CSAwallace_cska32_and_9_13;
  wire u_CSAwallace_cska32_and_10_13;
  wire u_CSAwallace_cska32_and_11_13;
  wire u_CSAwallace_cska32_and_12_13;
  wire u_CSAwallace_cska32_and_13_13;
  wire u_CSAwallace_cska32_and_14_13;
  wire u_CSAwallace_cska32_and_15_13;
  wire u_CSAwallace_cska32_and_16_13;
  wire u_CSAwallace_cska32_and_17_13;
  wire u_CSAwallace_cska32_and_18_13;
  wire u_CSAwallace_cska32_and_19_13;
  wire u_CSAwallace_cska32_and_20_13;
  wire u_CSAwallace_cska32_and_21_13;
  wire u_CSAwallace_cska32_and_22_13;
  wire u_CSAwallace_cska32_and_23_13;
  wire u_CSAwallace_cska32_and_24_13;
  wire u_CSAwallace_cska32_and_25_13;
  wire u_CSAwallace_cska32_and_26_13;
  wire u_CSAwallace_cska32_and_27_13;
  wire u_CSAwallace_cska32_and_28_13;
  wire u_CSAwallace_cska32_and_29_13;
  wire u_CSAwallace_cska32_and_30_13;
  wire u_CSAwallace_cska32_and_31_13;
  wire u_CSAwallace_cska32_and_0_14;
  wire u_CSAwallace_cska32_and_1_14;
  wire u_CSAwallace_cska32_and_2_14;
  wire u_CSAwallace_cska32_and_3_14;
  wire u_CSAwallace_cska32_and_4_14;
  wire u_CSAwallace_cska32_and_5_14;
  wire u_CSAwallace_cska32_and_6_14;
  wire u_CSAwallace_cska32_and_7_14;
  wire u_CSAwallace_cska32_and_8_14;
  wire u_CSAwallace_cska32_and_9_14;
  wire u_CSAwallace_cska32_and_10_14;
  wire u_CSAwallace_cska32_and_11_14;
  wire u_CSAwallace_cska32_and_12_14;
  wire u_CSAwallace_cska32_and_13_14;
  wire u_CSAwallace_cska32_and_14_14;
  wire u_CSAwallace_cska32_and_15_14;
  wire u_CSAwallace_cska32_and_16_14;
  wire u_CSAwallace_cska32_and_17_14;
  wire u_CSAwallace_cska32_and_18_14;
  wire u_CSAwallace_cska32_and_19_14;
  wire u_CSAwallace_cska32_and_20_14;
  wire u_CSAwallace_cska32_and_21_14;
  wire u_CSAwallace_cska32_and_22_14;
  wire u_CSAwallace_cska32_and_23_14;
  wire u_CSAwallace_cska32_and_24_14;
  wire u_CSAwallace_cska32_and_25_14;
  wire u_CSAwallace_cska32_and_26_14;
  wire u_CSAwallace_cska32_and_27_14;
  wire u_CSAwallace_cska32_and_28_14;
  wire u_CSAwallace_cska32_and_29_14;
  wire u_CSAwallace_cska32_and_30_14;
  wire u_CSAwallace_cska32_and_31_14;
  wire u_CSAwallace_cska32_and_0_15;
  wire u_CSAwallace_cska32_and_1_15;
  wire u_CSAwallace_cska32_and_2_15;
  wire u_CSAwallace_cska32_and_3_15;
  wire u_CSAwallace_cska32_and_4_15;
  wire u_CSAwallace_cska32_and_5_15;
  wire u_CSAwallace_cska32_and_6_15;
  wire u_CSAwallace_cska32_and_7_15;
  wire u_CSAwallace_cska32_and_8_15;
  wire u_CSAwallace_cska32_and_9_15;
  wire u_CSAwallace_cska32_and_10_15;
  wire u_CSAwallace_cska32_and_11_15;
  wire u_CSAwallace_cska32_and_12_15;
  wire u_CSAwallace_cska32_and_13_15;
  wire u_CSAwallace_cska32_and_14_15;
  wire u_CSAwallace_cska32_and_15_15;
  wire u_CSAwallace_cska32_and_16_15;
  wire u_CSAwallace_cska32_and_17_15;
  wire u_CSAwallace_cska32_and_18_15;
  wire u_CSAwallace_cska32_and_19_15;
  wire u_CSAwallace_cska32_and_20_15;
  wire u_CSAwallace_cska32_and_21_15;
  wire u_CSAwallace_cska32_and_22_15;
  wire u_CSAwallace_cska32_and_23_15;
  wire u_CSAwallace_cska32_and_24_15;
  wire u_CSAwallace_cska32_and_25_15;
  wire u_CSAwallace_cska32_and_26_15;
  wire u_CSAwallace_cska32_and_27_15;
  wire u_CSAwallace_cska32_and_28_15;
  wire u_CSAwallace_cska32_and_29_15;
  wire u_CSAwallace_cska32_and_30_15;
  wire u_CSAwallace_cska32_and_31_15;
  wire u_CSAwallace_cska32_and_0_16;
  wire u_CSAwallace_cska32_and_1_16;
  wire u_CSAwallace_cska32_and_2_16;
  wire u_CSAwallace_cska32_and_3_16;
  wire u_CSAwallace_cska32_and_4_16;
  wire u_CSAwallace_cska32_and_5_16;
  wire u_CSAwallace_cska32_and_6_16;
  wire u_CSAwallace_cska32_and_7_16;
  wire u_CSAwallace_cska32_and_8_16;
  wire u_CSAwallace_cska32_and_9_16;
  wire u_CSAwallace_cska32_and_10_16;
  wire u_CSAwallace_cska32_and_11_16;
  wire u_CSAwallace_cska32_and_12_16;
  wire u_CSAwallace_cska32_and_13_16;
  wire u_CSAwallace_cska32_and_14_16;
  wire u_CSAwallace_cska32_and_15_16;
  wire u_CSAwallace_cska32_and_16_16;
  wire u_CSAwallace_cska32_and_17_16;
  wire u_CSAwallace_cska32_and_18_16;
  wire u_CSAwallace_cska32_and_19_16;
  wire u_CSAwallace_cska32_and_20_16;
  wire u_CSAwallace_cska32_and_21_16;
  wire u_CSAwallace_cska32_and_22_16;
  wire u_CSAwallace_cska32_and_23_16;
  wire u_CSAwallace_cska32_and_24_16;
  wire u_CSAwallace_cska32_and_25_16;
  wire u_CSAwallace_cska32_and_26_16;
  wire u_CSAwallace_cska32_and_27_16;
  wire u_CSAwallace_cska32_and_28_16;
  wire u_CSAwallace_cska32_and_29_16;
  wire u_CSAwallace_cska32_and_30_16;
  wire u_CSAwallace_cska32_and_31_16;
  wire u_CSAwallace_cska32_and_0_17;
  wire u_CSAwallace_cska32_and_1_17;
  wire u_CSAwallace_cska32_and_2_17;
  wire u_CSAwallace_cska32_and_3_17;
  wire u_CSAwallace_cska32_and_4_17;
  wire u_CSAwallace_cska32_and_5_17;
  wire u_CSAwallace_cska32_and_6_17;
  wire u_CSAwallace_cska32_and_7_17;
  wire u_CSAwallace_cska32_and_8_17;
  wire u_CSAwallace_cska32_and_9_17;
  wire u_CSAwallace_cska32_and_10_17;
  wire u_CSAwallace_cska32_and_11_17;
  wire u_CSAwallace_cska32_and_12_17;
  wire u_CSAwallace_cska32_and_13_17;
  wire u_CSAwallace_cska32_and_14_17;
  wire u_CSAwallace_cska32_and_15_17;
  wire u_CSAwallace_cska32_and_16_17;
  wire u_CSAwallace_cska32_and_17_17;
  wire u_CSAwallace_cska32_and_18_17;
  wire u_CSAwallace_cska32_and_19_17;
  wire u_CSAwallace_cska32_and_20_17;
  wire u_CSAwallace_cska32_and_21_17;
  wire u_CSAwallace_cska32_and_22_17;
  wire u_CSAwallace_cska32_and_23_17;
  wire u_CSAwallace_cska32_and_24_17;
  wire u_CSAwallace_cska32_and_25_17;
  wire u_CSAwallace_cska32_and_26_17;
  wire u_CSAwallace_cska32_and_27_17;
  wire u_CSAwallace_cska32_and_28_17;
  wire u_CSAwallace_cska32_and_29_17;
  wire u_CSAwallace_cska32_and_30_17;
  wire u_CSAwallace_cska32_and_31_17;
  wire u_CSAwallace_cska32_and_0_18;
  wire u_CSAwallace_cska32_and_1_18;
  wire u_CSAwallace_cska32_and_2_18;
  wire u_CSAwallace_cska32_and_3_18;
  wire u_CSAwallace_cska32_and_4_18;
  wire u_CSAwallace_cska32_and_5_18;
  wire u_CSAwallace_cska32_and_6_18;
  wire u_CSAwallace_cska32_and_7_18;
  wire u_CSAwallace_cska32_and_8_18;
  wire u_CSAwallace_cska32_and_9_18;
  wire u_CSAwallace_cska32_and_10_18;
  wire u_CSAwallace_cska32_and_11_18;
  wire u_CSAwallace_cska32_and_12_18;
  wire u_CSAwallace_cska32_and_13_18;
  wire u_CSAwallace_cska32_and_14_18;
  wire u_CSAwallace_cska32_and_15_18;
  wire u_CSAwallace_cska32_and_16_18;
  wire u_CSAwallace_cska32_and_17_18;
  wire u_CSAwallace_cska32_and_18_18;
  wire u_CSAwallace_cska32_and_19_18;
  wire u_CSAwallace_cska32_and_20_18;
  wire u_CSAwallace_cska32_and_21_18;
  wire u_CSAwallace_cska32_and_22_18;
  wire u_CSAwallace_cska32_and_23_18;
  wire u_CSAwallace_cska32_and_24_18;
  wire u_CSAwallace_cska32_and_25_18;
  wire u_CSAwallace_cska32_and_26_18;
  wire u_CSAwallace_cska32_and_27_18;
  wire u_CSAwallace_cska32_and_28_18;
  wire u_CSAwallace_cska32_and_29_18;
  wire u_CSAwallace_cska32_and_30_18;
  wire u_CSAwallace_cska32_and_31_18;
  wire u_CSAwallace_cska32_and_0_19;
  wire u_CSAwallace_cska32_and_1_19;
  wire u_CSAwallace_cska32_and_2_19;
  wire u_CSAwallace_cska32_and_3_19;
  wire u_CSAwallace_cska32_and_4_19;
  wire u_CSAwallace_cska32_and_5_19;
  wire u_CSAwallace_cska32_and_6_19;
  wire u_CSAwallace_cska32_and_7_19;
  wire u_CSAwallace_cska32_and_8_19;
  wire u_CSAwallace_cska32_and_9_19;
  wire u_CSAwallace_cska32_and_10_19;
  wire u_CSAwallace_cska32_and_11_19;
  wire u_CSAwallace_cska32_and_12_19;
  wire u_CSAwallace_cska32_and_13_19;
  wire u_CSAwallace_cska32_and_14_19;
  wire u_CSAwallace_cska32_and_15_19;
  wire u_CSAwallace_cska32_and_16_19;
  wire u_CSAwallace_cska32_and_17_19;
  wire u_CSAwallace_cska32_and_18_19;
  wire u_CSAwallace_cska32_and_19_19;
  wire u_CSAwallace_cska32_and_20_19;
  wire u_CSAwallace_cska32_and_21_19;
  wire u_CSAwallace_cska32_and_22_19;
  wire u_CSAwallace_cska32_and_23_19;
  wire u_CSAwallace_cska32_and_24_19;
  wire u_CSAwallace_cska32_and_25_19;
  wire u_CSAwallace_cska32_and_26_19;
  wire u_CSAwallace_cska32_and_27_19;
  wire u_CSAwallace_cska32_and_28_19;
  wire u_CSAwallace_cska32_and_29_19;
  wire u_CSAwallace_cska32_and_30_19;
  wire u_CSAwallace_cska32_and_31_19;
  wire u_CSAwallace_cska32_and_0_20;
  wire u_CSAwallace_cska32_and_1_20;
  wire u_CSAwallace_cska32_and_2_20;
  wire u_CSAwallace_cska32_and_3_20;
  wire u_CSAwallace_cska32_and_4_20;
  wire u_CSAwallace_cska32_and_5_20;
  wire u_CSAwallace_cska32_and_6_20;
  wire u_CSAwallace_cska32_and_7_20;
  wire u_CSAwallace_cska32_and_8_20;
  wire u_CSAwallace_cska32_and_9_20;
  wire u_CSAwallace_cska32_and_10_20;
  wire u_CSAwallace_cska32_and_11_20;
  wire u_CSAwallace_cska32_and_12_20;
  wire u_CSAwallace_cska32_and_13_20;
  wire u_CSAwallace_cska32_and_14_20;
  wire u_CSAwallace_cska32_and_15_20;
  wire u_CSAwallace_cska32_and_16_20;
  wire u_CSAwallace_cska32_and_17_20;
  wire u_CSAwallace_cska32_and_18_20;
  wire u_CSAwallace_cska32_and_19_20;
  wire u_CSAwallace_cska32_and_20_20;
  wire u_CSAwallace_cska32_and_21_20;
  wire u_CSAwallace_cska32_and_22_20;
  wire u_CSAwallace_cska32_and_23_20;
  wire u_CSAwallace_cska32_and_24_20;
  wire u_CSAwallace_cska32_and_25_20;
  wire u_CSAwallace_cska32_and_26_20;
  wire u_CSAwallace_cska32_and_27_20;
  wire u_CSAwallace_cska32_and_28_20;
  wire u_CSAwallace_cska32_and_29_20;
  wire u_CSAwallace_cska32_and_30_20;
  wire u_CSAwallace_cska32_and_31_20;
  wire u_CSAwallace_cska32_and_0_21;
  wire u_CSAwallace_cska32_and_1_21;
  wire u_CSAwallace_cska32_and_2_21;
  wire u_CSAwallace_cska32_and_3_21;
  wire u_CSAwallace_cska32_and_4_21;
  wire u_CSAwallace_cska32_and_5_21;
  wire u_CSAwallace_cska32_and_6_21;
  wire u_CSAwallace_cska32_and_7_21;
  wire u_CSAwallace_cska32_and_8_21;
  wire u_CSAwallace_cska32_and_9_21;
  wire u_CSAwallace_cska32_and_10_21;
  wire u_CSAwallace_cska32_and_11_21;
  wire u_CSAwallace_cska32_and_12_21;
  wire u_CSAwallace_cska32_and_13_21;
  wire u_CSAwallace_cska32_and_14_21;
  wire u_CSAwallace_cska32_and_15_21;
  wire u_CSAwallace_cska32_and_16_21;
  wire u_CSAwallace_cska32_and_17_21;
  wire u_CSAwallace_cska32_and_18_21;
  wire u_CSAwallace_cska32_and_19_21;
  wire u_CSAwallace_cska32_and_20_21;
  wire u_CSAwallace_cska32_and_21_21;
  wire u_CSAwallace_cska32_and_22_21;
  wire u_CSAwallace_cska32_and_23_21;
  wire u_CSAwallace_cska32_and_24_21;
  wire u_CSAwallace_cska32_and_25_21;
  wire u_CSAwallace_cska32_and_26_21;
  wire u_CSAwallace_cska32_and_27_21;
  wire u_CSAwallace_cska32_and_28_21;
  wire u_CSAwallace_cska32_and_29_21;
  wire u_CSAwallace_cska32_and_30_21;
  wire u_CSAwallace_cska32_and_31_21;
  wire u_CSAwallace_cska32_and_0_22;
  wire u_CSAwallace_cska32_and_1_22;
  wire u_CSAwallace_cska32_and_2_22;
  wire u_CSAwallace_cska32_and_3_22;
  wire u_CSAwallace_cska32_and_4_22;
  wire u_CSAwallace_cska32_and_5_22;
  wire u_CSAwallace_cska32_and_6_22;
  wire u_CSAwallace_cska32_and_7_22;
  wire u_CSAwallace_cska32_and_8_22;
  wire u_CSAwallace_cska32_and_9_22;
  wire u_CSAwallace_cska32_and_10_22;
  wire u_CSAwallace_cska32_and_11_22;
  wire u_CSAwallace_cska32_and_12_22;
  wire u_CSAwallace_cska32_and_13_22;
  wire u_CSAwallace_cska32_and_14_22;
  wire u_CSAwallace_cska32_and_15_22;
  wire u_CSAwallace_cska32_and_16_22;
  wire u_CSAwallace_cska32_and_17_22;
  wire u_CSAwallace_cska32_and_18_22;
  wire u_CSAwallace_cska32_and_19_22;
  wire u_CSAwallace_cska32_and_20_22;
  wire u_CSAwallace_cska32_and_21_22;
  wire u_CSAwallace_cska32_and_22_22;
  wire u_CSAwallace_cska32_and_23_22;
  wire u_CSAwallace_cska32_and_24_22;
  wire u_CSAwallace_cska32_and_25_22;
  wire u_CSAwallace_cska32_and_26_22;
  wire u_CSAwallace_cska32_and_27_22;
  wire u_CSAwallace_cska32_and_28_22;
  wire u_CSAwallace_cska32_and_29_22;
  wire u_CSAwallace_cska32_and_30_22;
  wire u_CSAwallace_cska32_and_31_22;
  wire u_CSAwallace_cska32_and_0_23;
  wire u_CSAwallace_cska32_and_1_23;
  wire u_CSAwallace_cska32_and_2_23;
  wire u_CSAwallace_cska32_and_3_23;
  wire u_CSAwallace_cska32_and_4_23;
  wire u_CSAwallace_cska32_and_5_23;
  wire u_CSAwallace_cska32_and_6_23;
  wire u_CSAwallace_cska32_and_7_23;
  wire u_CSAwallace_cska32_and_8_23;
  wire u_CSAwallace_cska32_and_9_23;
  wire u_CSAwallace_cska32_and_10_23;
  wire u_CSAwallace_cska32_and_11_23;
  wire u_CSAwallace_cska32_and_12_23;
  wire u_CSAwallace_cska32_and_13_23;
  wire u_CSAwallace_cska32_and_14_23;
  wire u_CSAwallace_cska32_and_15_23;
  wire u_CSAwallace_cska32_and_16_23;
  wire u_CSAwallace_cska32_and_17_23;
  wire u_CSAwallace_cska32_and_18_23;
  wire u_CSAwallace_cska32_and_19_23;
  wire u_CSAwallace_cska32_and_20_23;
  wire u_CSAwallace_cska32_and_21_23;
  wire u_CSAwallace_cska32_and_22_23;
  wire u_CSAwallace_cska32_and_23_23;
  wire u_CSAwallace_cska32_and_24_23;
  wire u_CSAwallace_cska32_and_25_23;
  wire u_CSAwallace_cska32_and_26_23;
  wire u_CSAwallace_cska32_and_27_23;
  wire u_CSAwallace_cska32_and_28_23;
  wire u_CSAwallace_cska32_and_29_23;
  wire u_CSAwallace_cska32_and_30_23;
  wire u_CSAwallace_cska32_and_31_23;
  wire u_CSAwallace_cska32_and_0_24;
  wire u_CSAwallace_cska32_and_1_24;
  wire u_CSAwallace_cska32_and_2_24;
  wire u_CSAwallace_cska32_and_3_24;
  wire u_CSAwallace_cska32_and_4_24;
  wire u_CSAwallace_cska32_and_5_24;
  wire u_CSAwallace_cska32_and_6_24;
  wire u_CSAwallace_cska32_and_7_24;
  wire u_CSAwallace_cska32_and_8_24;
  wire u_CSAwallace_cska32_and_9_24;
  wire u_CSAwallace_cska32_and_10_24;
  wire u_CSAwallace_cska32_and_11_24;
  wire u_CSAwallace_cska32_and_12_24;
  wire u_CSAwallace_cska32_and_13_24;
  wire u_CSAwallace_cska32_and_14_24;
  wire u_CSAwallace_cska32_and_15_24;
  wire u_CSAwallace_cska32_and_16_24;
  wire u_CSAwallace_cska32_and_17_24;
  wire u_CSAwallace_cska32_and_18_24;
  wire u_CSAwallace_cska32_and_19_24;
  wire u_CSAwallace_cska32_and_20_24;
  wire u_CSAwallace_cska32_and_21_24;
  wire u_CSAwallace_cska32_and_22_24;
  wire u_CSAwallace_cska32_and_23_24;
  wire u_CSAwallace_cska32_and_24_24;
  wire u_CSAwallace_cska32_and_25_24;
  wire u_CSAwallace_cska32_and_26_24;
  wire u_CSAwallace_cska32_and_27_24;
  wire u_CSAwallace_cska32_and_28_24;
  wire u_CSAwallace_cska32_and_29_24;
  wire u_CSAwallace_cska32_and_30_24;
  wire u_CSAwallace_cska32_and_31_24;
  wire u_CSAwallace_cska32_and_0_25;
  wire u_CSAwallace_cska32_and_1_25;
  wire u_CSAwallace_cska32_and_2_25;
  wire u_CSAwallace_cska32_and_3_25;
  wire u_CSAwallace_cska32_and_4_25;
  wire u_CSAwallace_cska32_and_5_25;
  wire u_CSAwallace_cska32_and_6_25;
  wire u_CSAwallace_cska32_and_7_25;
  wire u_CSAwallace_cska32_and_8_25;
  wire u_CSAwallace_cska32_and_9_25;
  wire u_CSAwallace_cska32_and_10_25;
  wire u_CSAwallace_cska32_and_11_25;
  wire u_CSAwallace_cska32_and_12_25;
  wire u_CSAwallace_cska32_and_13_25;
  wire u_CSAwallace_cska32_and_14_25;
  wire u_CSAwallace_cska32_and_15_25;
  wire u_CSAwallace_cska32_and_16_25;
  wire u_CSAwallace_cska32_and_17_25;
  wire u_CSAwallace_cska32_and_18_25;
  wire u_CSAwallace_cska32_and_19_25;
  wire u_CSAwallace_cska32_and_20_25;
  wire u_CSAwallace_cska32_and_21_25;
  wire u_CSAwallace_cska32_and_22_25;
  wire u_CSAwallace_cska32_and_23_25;
  wire u_CSAwallace_cska32_and_24_25;
  wire u_CSAwallace_cska32_and_25_25;
  wire u_CSAwallace_cska32_and_26_25;
  wire u_CSAwallace_cska32_and_27_25;
  wire u_CSAwallace_cska32_and_28_25;
  wire u_CSAwallace_cska32_and_29_25;
  wire u_CSAwallace_cska32_and_30_25;
  wire u_CSAwallace_cska32_and_31_25;
  wire u_CSAwallace_cska32_and_0_26;
  wire u_CSAwallace_cska32_and_1_26;
  wire u_CSAwallace_cska32_and_2_26;
  wire u_CSAwallace_cska32_and_3_26;
  wire u_CSAwallace_cska32_and_4_26;
  wire u_CSAwallace_cska32_and_5_26;
  wire u_CSAwallace_cska32_and_6_26;
  wire u_CSAwallace_cska32_and_7_26;
  wire u_CSAwallace_cska32_and_8_26;
  wire u_CSAwallace_cska32_and_9_26;
  wire u_CSAwallace_cska32_and_10_26;
  wire u_CSAwallace_cska32_and_11_26;
  wire u_CSAwallace_cska32_and_12_26;
  wire u_CSAwallace_cska32_and_13_26;
  wire u_CSAwallace_cska32_and_14_26;
  wire u_CSAwallace_cska32_and_15_26;
  wire u_CSAwallace_cska32_and_16_26;
  wire u_CSAwallace_cska32_and_17_26;
  wire u_CSAwallace_cska32_and_18_26;
  wire u_CSAwallace_cska32_and_19_26;
  wire u_CSAwallace_cska32_and_20_26;
  wire u_CSAwallace_cska32_and_21_26;
  wire u_CSAwallace_cska32_and_22_26;
  wire u_CSAwallace_cska32_and_23_26;
  wire u_CSAwallace_cska32_and_24_26;
  wire u_CSAwallace_cska32_and_25_26;
  wire u_CSAwallace_cska32_and_26_26;
  wire u_CSAwallace_cska32_and_27_26;
  wire u_CSAwallace_cska32_and_28_26;
  wire u_CSAwallace_cska32_and_29_26;
  wire u_CSAwallace_cska32_and_30_26;
  wire u_CSAwallace_cska32_and_31_26;
  wire u_CSAwallace_cska32_and_0_27;
  wire u_CSAwallace_cska32_and_1_27;
  wire u_CSAwallace_cska32_and_2_27;
  wire u_CSAwallace_cska32_and_3_27;
  wire u_CSAwallace_cska32_and_4_27;
  wire u_CSAwallace_cska32_and_5_27;
  wire u_CSAwallace_cska32_and_6_27;
  wire u_CSAwallace_cska32_and_7_27;
  wire u_CSAwallace_cska32_and_8_27;
  wire u_CSAwallace_cska32_and_9_27;
  wire u_CSAwallace_cska32_and_10_27;
  wire u_CSAwallace_cska32_and_11_27;
  wire u_CSAwallace_cska32_and_12_27;
  wire u_CSAwallace_cska32_and_13_27;
  wire u_CSAwallace_cska32_and_14_27;
  wire u_CSAwallace_cska32_and_15_27;
  wire u_CSAwallace_cska32_and_16_27;
  wire u_CSAwallace_cska32_and_17_27;
  wire u_CSAwallace_cska32_and_18_27;
  wire u_CSAwallace_cska32_and_19_27;
  wire u_CSAwallace_cska32_and_20_27;
  wire u_CSAwallace_cska32_and_21_27;
  wire u_CSAwallace_cska32_and_22_27;
  wire u_CSAwallace_cska32_and_23_27;
  wire u_CSAwallace_cska32_and_24_27;
  wire u_CSAwallace_cska32_and_25_27;
  wire u_CSAwallace_cska32_and_26_27;
  wire u_CSAwallace_cska32_and_27_27;
  wire u_CSAwallace_cska32_and_28_27;
  wire u_CSAwallace_cska32_and_29_27;
  wire u_CSAwallace_cska32_and_30_27;
  wire u_CSAwallace_cska32_and_31_27;
  wire u_CSAwallace_cska32_and_0_28;
  wire u_CSAwallace_cska32_and_1_28;
  wire u_CSAwallace_cska32_and_2_28;
  wire u_CSAwallace_cska32_and_3_28;
  wire u_CSAwallace_cska32_and_4_28;
  wire u_CSAwallace_cska32_and_5_28;
  wire u_CSAwallace_cska32_and_6_28;
  wire u_CSAwallace_cska32_and_7_28;
  wire u_CSAwallace_cska32_and_8_28;
  wire u_CSAwallace_cska32_and_9_28;
  wire u_CSAwallace_cska32_and_10_28;
  wire u_CSAwallace_cska32_and_11_28;
  wire u_CSAwallace_cska32_and_12_28;
  wire u_CSAwallace_cska32_and_13_28;
  wire u_CSAwallace_cska32_and_14_28;
  wire u_CSAwallace_cska32_and_15_28;
  wire u_CSAwallace_cska32_and_16_28;
  wire u_CSAwallace_cska32_and_17_28;
  wire u_CSAwallace_cska32_and_18_28;
  wire u_CSAwallace_cska32_and_19_28;
  wire u_CSAwallace_cska32_and_20_28;
  wire u_CSAwallace_cska32_and_21_28;
  wire u_CSAwallace_cska32_and_22_28;
  wire u_CSAwallace_cska32_and_23_28;
  wire u_CSAwallace_cska32_and_24_28;
  wire u_CSAwallace_cska32_and_25_28;
  wire u_CSAwallace_cska32_and_26_28;
  wire u_CSAwallace_cska32_and_27_28;
  wire u_CSAwallace_cska32_and_28_28;
  wire u_CSAwallace_cska32_and_29_28;
  wire u_CSAwallace_cska32_and_30_28;
  wire u_CSAwallace_cska32_and_31_28;
  wire u_CSAwallace_cska32_and_0_29;
  wire u_CSAwallace_cska32_and_1_29;
  wire u_CSAwallace_cska32_and_2_29;
  wire u_CSAwallace_cska32_and_3_29;
  wire u_CSAwallace_cska32_and_4_29;
  wire u_CSAwallace_cska32_and_5_29;
  wire u_CSAwallace_cska32_and_6_29;
  wire u_CSAwallace_cska32_and_7_29;
  wire u_CSAwallace_cska32_and_8_29;
  wire u_CSAwallace_cska32_and_9_29;
  wire u_CSAwallace_cska32_and_10_29;
  wire u_CSAwallace_cska32_and_11_29;
  wire u_CSAwallace_cska32_and_12_29;
  wire u_CSAwallace_cska32_and_13_29;
  wire u_CSAwallace_cska32_and_14_29;
  wire u_CSAwallace_cska32_and_15_29;
  wire u_CSAwallace_cska32_and_16_29;
  wire u_CSAwallace_cska32_and_17_29;
  wire u_CSAwallace_cska32_and_18_29;
  wire u_CSAwallace_cska32_and_19_29;
  wire u_CSAwallace_cska32_and_20_29;
  wire u_CSAwallace_cska32_and_21_29;
  wire u_CSAwallace_cska32_and_22_29;
  wire u_CSAwallace_cska32_and_23_29;
  wire u_CSAwallace_cska32_and_24_29;
  wire u_CSAwallace_cska32_and_25_29;
  wire u_CSAwallace_cska32_and_26_29;
  wire u_CSAwallace_cska32_and_27_29;
  wire u_CSAwallace_cska32_and_28_29;
  wire u_CSAwallace_cska32_and_29_29;
  wire u_CSAwallace_cska32_and_30_29;
  wire u_CSAwallace_cska32_and_31_29;
  wire u_CSAwallace_cska32_and_0_30;
  wire u_CSAwallace_cska32_and_1_30;
  wire u_CSAwallace_cska32_and_2_30;
  wire u_CSAwallace_cska32_and_3_30;
  wire u_CSAwallace_cska32_and_4_30;
  wire u_CSAwallace_cska32_and_5_30;
  wire u_CSAwallace_cska32_and_6_30;
  wire u_CSAwallace_cska32_and_7_30;
  wire u_CSAwallace_cska32_and_8_30;
  wire u_CSAwallace_cska32_and_9_30;
  wire u_CSAwallace_cska32_and_10_30;
  wire u_CSAwallace_cska32_and_11_30;
  wire u_CSAwallace_cska32_and_12_30;
  wire u_CSAwallace_cska32_and_13_30;
  wire u_CSAwallace_cska32_and_14_30;
  wire u_CSAwallace_cska32_and_15_30;
  wire u_CSAwallace_cska32_and_16_30;
  wire u_CSAwallace_cska32_and_17_30;
  wire u_CSAwallace_cska32_and_18_30;
  wire u_CSAwallace_cska32_and_19_30;
  wire u_CSAwallace_cska32_and_20_30;
  wire u_CSAwallace_cska32_and_21_30;
  wire u_CSAwallace_cska32_and_22_30;
  wire u_CSAwallace_cska32_and_23_30;
  wire u_CSAwallace_cska32_and_24_30;
  wire u_CSAwallace_cska32_and_25_30;
  wire u_CSAwallace_cska32_and_26_30;
  wire u_CSAwallace_cska32_and_27_30;
  wire u_CSAwallace_cska32_and_28_30;
  wire u_CSAwallace_cska32_and_29_30;
  wire u_CSAwallace_cska32_and_30_30;
  wire u_CSAwallace_cska32_and_31_30;
  wire u_CSAwallace_cska32_and_0_31;
  wire u_CSAwallace_cska32_and_1_31;
  wire u_CSAwallace_cska32_and_2_31;
  wire u_CSAwallace_cska32_and_3_31;
  wire u_CSAwallace_cska32_and_4_31;
  wire u_CSAwallace_cska32_and_5_31;
  wire u_CSAwallace_cska32_and_6_31;
  wire u_CSAwallace_cska32_and_7_31;
  wire u_CSAwallace_cska32_and_8_31;
  wire u_CSAwallace_cska32_and_9_31;
  wire u_CSAwallace_cska32_and_10_31;
  wire u_CSAwallace_cska32_and_11_31;
  wire u_CSAwallace_cska32_and_12_31;
  wire u_CSAwallace_cska32_and_13_31;
  wire u_CSAwallace_cska32_and_14_31;
  wire u_CSAwallace_cska32_and_15_31;
  wire u_CSAwallace_cska32_and_16_31;
  wire u_CSAwallace_cska32_and_17_31;
  wire u_CSAwallace_cska32_and_18_31;
  wire u_CSAwallace_cska32_and_19_31;
  wire u_CSAwallace_cska32_and_20_31;
  wire u_CSAwallace_cska32_and_21_31;
  wire u_CSAwallace_cska32_and_22_31;
  wire u_CSAwallace_cska32_and_23_31;
  wire u_CSAwallace_cska32_and_24_31;
  wire u_CSAwallace_cska32_and_25_31;
  wire u_CSAwallace_cska32_and_26_31;
  wire u_CSAwallace_cska32_and_27_31;
  wire u_CSAwallace_cska32_and_28_31;
  wire u_CSAwallace_cska32_and_29_31;
  wire u_CSAwallace_cska32_and_30_31;
  wire u_CSAwallace_cska32_and_31_31;
  wire u_CSAwallace_cska32_csa0_csa_component_fa1_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa1_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa2_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa2_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa2_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa2_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa2_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa3_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa3_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa3_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa3_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa3_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa4_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa4_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa4_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa4_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa4_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa5_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa5_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa5_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa5_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa5_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa6_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa6_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa6_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa6_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa6_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa7_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa7_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa7_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa8_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa8_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa8_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa9_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa9_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa9_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa10_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa10_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa10_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa0_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa0_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa4_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa4_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa5_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa5_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa5_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa5_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa5_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa6_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa6_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa6_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa6_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa6_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa7_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa7_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa7_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa8_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa8_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa8_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa9_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa9_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa9_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa10_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa10_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa10_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa1_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa1_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa8_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa8_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa8_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa9_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa9_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa9_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa10_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa10_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa10_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa2_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa2_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa3_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa3_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa4_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa4_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa5_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa5_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa6_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa6_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa7_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa7_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa53_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa53_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa53_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa54_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa54_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa54_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa55_xor0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa55_and0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa55_or0;
  wire u_CSAwallace_cska32_csa8_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa8_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa53_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa53_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa53_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa54_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa54_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa54_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa55_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa55_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa55_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa56_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa56_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa56_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa57_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa57_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa57_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa58_xor0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa58_and0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa58_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa58_and1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa58_or0;
  wire u_CSAwallace_cska32_csa9_csa_component_fa59_xor1;
  wire u_CSAwallace_cska32_csa9_csa_component_fa59_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa2_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa2_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa3_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa3_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa3_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa3_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa3_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa4_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa4_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa4_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa4_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa4_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa5_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa5_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa5_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa5_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa5_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa6_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa6_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa6_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa6_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa6_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa7_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa7_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa7_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa8_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa8_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa8_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa9_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa9_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa9_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa10_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa10_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa10_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa10_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa10_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa6_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa6_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa8_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa8_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa8_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa9_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa9_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa9_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa10_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa10_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa10_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa11_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa11_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa12_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa12_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa13_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa13_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa14_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa14_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa53_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa53_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa53_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa54_xor0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa54_and0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa54_or0;
  wire u_CSAwallace_cska32_csa15_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa15_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa53_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa53_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa53_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa54_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa54_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa54_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa55_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa55_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa55_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa56_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa56_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa56_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa57_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa57_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa57_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa58_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa58_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa58_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa58_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa58_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa59_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa59_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa59_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa59_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa59_or0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa60_xor0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa60_and0;
  wire u_CSAwallace_cska32_csa16_csa_component_fa60_xor1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa60_and1;
  wire u_CSAwallace_cska32_csa16_csa_component_fa60_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa3_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa3_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa4_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa4_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa5_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa5_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa5_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa5_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa5_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa6_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa6_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa6_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa6_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa6_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa7_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa7_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa7_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa8_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa8_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa8_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa9_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa9_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa9_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa10_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa10_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa10_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa17_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa17_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa18_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa18_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa19_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa19_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa20_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa20_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa53_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa53_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa53_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa54_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa54_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa54_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa55_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa55_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa55_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa56_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa56_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa56_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa57_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa57_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa57_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa58_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa58_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa58_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa58_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa58_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa59_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa59_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa59_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa59_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa59_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa60_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa60_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa60_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa60_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa60_or0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa61_xor0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa61_and0;
  wire u_CSAwallace_cska32_csa21_csa_component_fa61_xor1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa61_and1;
  wire u_CSAwallace_cska32_csa21_csa_component_fa61_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa4_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa4_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa5_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa5_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa6_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa6_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa7_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa7_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa7_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa8_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa8_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa8_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa9_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa9_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa9_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa10_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa10_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa10_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa22_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa22_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa23_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa23_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa53_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa53_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa53_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa54_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa54_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa54_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa55_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa55_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa55_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa56_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa56_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa56_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa57_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa57_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa57_or0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa58_xor0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa58_and0;
  wire u_CSAwallace_cska32_csa24_csa_component_fa58_xor1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa58_and1;
  wire u_CSAwallace_cska32_csa24_csa_component_fa58_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa5_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa5_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa6_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa6_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa10_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa10_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa10_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa11_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa11_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa11_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa12_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa12_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa12_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa13_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa13_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa13_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa14_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa14_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa14_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa25_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa25_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa26_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa58_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa58_and1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa59_xor1;
  wire u_CSAwallace_cska32_csa26_csa_component_fa59_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa6_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa6_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa15_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa15_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa15_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa16_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa16_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa16_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa17_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa17_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa17_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa18_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa18_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa18_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa19_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa19_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa19_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa20_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa20_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa20_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa21_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa21_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa21_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa27_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa27_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa7_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa7_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa22_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa22_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa22_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa23_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa23_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa23_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa24_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa24_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa24_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa25_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa25_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa25_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa26_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa26_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa26_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa27_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa27_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa27_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa28_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa28_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa28_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa29_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa29_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa29_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa30_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa30_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa30_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa53_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa53_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa53_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa54_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa54_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa54_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa55_xor0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa55_and0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa55_or0;
  wire u_CSAwallace_cska32_csa28_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa58_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa58_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa59_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa59_and1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa60_xor1;
  wire u_CSAwallace_cska32_csa28_csa_component_fa60_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa8_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa8_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa9_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa9_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa10_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa10_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa11_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa11_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa12_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa12_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa13_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa13_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa14_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa14_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa15_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa15_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa16_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa16_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa17_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa17_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa18_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa18_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa19_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa19_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa20_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa20_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa21_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa21_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa22_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa22_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa23_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa23_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa24_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa24_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa25_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa25_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa26_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa26_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa27_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa27_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa28_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa28_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa29_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa29_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa30_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa30_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa31_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa31_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa31_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa31_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa31_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa32_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa32_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa32_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa32_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa32_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa33_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa33_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa33_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa33_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa33_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa34_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa34_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa34_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa34_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa34_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa35_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa35_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa35_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa35_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa35_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa36_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa36_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa36_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa36_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa36_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa37_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa37_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa37_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa37_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa37_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa38_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa38_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa38_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa38_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa38_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa39_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa39_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa39_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa39_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa39_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa40_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa40_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa40_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa40_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa40_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa41_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa41_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa41_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa41_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa41_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa42_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa42_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa42_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa42_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa42_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa43_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa43_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa43_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa43_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa43_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa44_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa44_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa44_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa44_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa44_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa45_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa45_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa45_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa45_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa45_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa46_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa46_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa46_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa46_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa46_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa47_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa47_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa47_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa47_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa47_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa48_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa48_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa48_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa48_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa48_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa49_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa49_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa49_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa49_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa49_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa50_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa50_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa50_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa50_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa50_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa51_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa51_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa51_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa51_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa51_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa52_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa52_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa52_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa52_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa52_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa53_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa53_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa53_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa53_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa53_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa54_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa54_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa54_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa54_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa54_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa55_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa55_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa55_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa55_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa55_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa56_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa56_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa56_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa56_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa56_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa57_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa57_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa57_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa57_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa57_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa58_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa58_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa58_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa58_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa58_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa59_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa59_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa59_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa59_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa59_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa60_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa60_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa60_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa60_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa60_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa61_xor0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa61_and0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa61_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa61_and1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa61_or0;
  wire u_CSAwallace_cska32_csa29_csa_component_fa62_xor1;
  wire u_CSAwallace_cska32_csa29_csa_component_fa62_and1;
  wire u_CSAwallace_cska32_u_cska64_and_propagate00;
  wire u_CSAwallace_cska32_u_cska64_and_propagate01;
  wire u_CSAwallace_cska32_u_cska64_and_propagate02;
  wire u_CSAwallace_cska32_u_cska64_mux2to10_not0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate13;
  wire u_CSAwallace_cska32_u_cska64_and_propagate14;
  wire u_CSAwallace_cska32_u_cska64_and_propagate15;
  wire u_CSAwallace_cska32_u_cska64_mux2to11_not0;
  wire u_CSAwallace_cska32_u_cska64_xor9;
  wire u_CSAwallace_cska32_u_cska64_fa8_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa8_and0;
  wire u_CSAwallace_cska32_u_cska64_xor10;
  wire u_CSAwallace_cska32_u_cska64_fa9_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa9_and0;
  wire u_CSAwallace_cska32_u_cska64_fa9_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa9_and1;
  wire u_CSAwallace_cska32_u_cska64_fa9_or0;
  wire u_CSAwallace_cska32_u_cska64_xor11;
  wire u_CSAwallace_cska32_u_cska64_fa10_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa10_and0;
  wire u_CSAwallace_cska32_u_cska64_fa10_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa10_and1;
  wire u_CSAwallace_cska32_u_cska64_fa10_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate26;
  wire u_CSAwallace_cska32_u_cska64_and_propagate27;
  wire u_CSAwallace_cska32_u_cska64_and_propagate28;
  wire u_CSAwallace_cska32_u_cska64_mux2to12_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to12_and1;
  wire u_CSAwallace_cska32_u_cska64_xor12;
  wire u_CSAwallace_cska32_u_cska64_fa11_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa11_and0;
  wire u_CSAwallace_cska32_u_cska64_fa11_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa11_and1;
  wire u_CSAwallace_cska32_u_cska64_fa11_or0;
  wire u_CSAwallace_cska32_u_cska64_xor13;
  wire u_CSAwallace_cska32_u_cska64_fa12_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa12_and0;
  wire u_CSAwallace_cska32_u_cska64_fa12_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa12_and1;
  wire u_CSAwallace_cska32_u_cska64_fa12_or0;
  wire u_CSAwallace_cska32_u_cska64_xor14;
  wire u_CSAwallace_cska32_u_cska64_fa13_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa13_and0;
  wire u_CSAwallace_cska32_u_cska64_fa13_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa13_and1;
  wire u_CSAwallace_cska32_u_cska64_fa13_or0;
  wire u_CSAwallace_cska32_u_cska64_xor15;
  wire u_CSAwallace_cska32_u_cska64_fa14_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa14_and0;
  wire u_CSAwallace_cska32_u_cska64_fa14_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa14_and1;
  wire u_CSAwallace_cska32_u_cska64_fa14_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate39;
  wire u_CSAwallace_cska32_u_cska64_and_propagate310;
  wire u_CSAwallace_cska32_u_cska64_and_propagate311;
  wire u_CSAwallace_cska32_u_cska64_mux2to13_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to13_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to13_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to13_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor16;
  wire u_CSAwallace_cska32_u_cska64_fa15_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa15_and0;
  wire u_CSAwallace_cska32_u_cska64_fa15_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa15_and1;
  wire u_CSAwallace_cska32_u_cska64_fa15_or0;
  wire u_CSAwallace_cska32_u_cska64_xor17;
  wire u_CSAwallace_cska32_u_cska64_fa16_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa16_and0;
  wire u_CSAwallace_cska32_u_cska64_fa16_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa16_and1;
  wire u_CSAwallace_cska32_u_cska64_fa16_or0;
  wire u_CSAwallace_cska32_u_cska64_xor18;
  wire u_CSAwallace_cska32_u_cska64_fa17_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa17_and0;
  wire u_CSAwallace_cska32_u_cska64_fa17_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa17_and1;
  wire u_CSAwallace_cska32_u_cska64_fa17_or0;
  wire u_CSAwallace_cska32_u_cska64_xor19;
  wire u_CSAwallace_cska32_u_cska64_fa18_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa18_and0;
  wire u_CSAwallace_cska32_u_cska64_fa18_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa18_and1;
  wire u_CSAwallace_cska32_u_cska64_fa18_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate412;
  wire u_CSAwallace_cska32_u_cska64_and_propagate413;
  wire u_CSAwallace_cska32_u_cska64_and_propagate414;
  wire u_CSAwallace_cska32_u_cska64_mux2to14_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to14_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to14_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to14_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor20;
  wire u_CSAwallace_cska32_u_cska64_fa19_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa19_and0;
  wire u_CSAwallace_cska32_u_cska64_fa19_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa19_and1;
  wire u_CSAwallace_cska32_u_cska64_fa19_or0;
  wire u_CSAwallace_cska32_u_cska64_xor21;
  wire u_CSAwallace_cska32_u_cska64_fa20_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa20_and0;
  wire u_CSAwallace_cska32_u_cska64_fa20_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa20_and1;
  wire u_CSAwallace_cska32_u_cska64_fa20_or0;
  wire u_CSAwallace_cska32_u_cska64_xor22;
  wire u_CSAwallace_cska32_u_cska64_fa21_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa21_and0;
  wire u_CSAwallace_cska32_u_cska64_fa21_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa21_and1;
  wire u_CSAwallace_cska32_u_cska64_fa21_or0;
  wire u_CSAwallace_cska32_u_cska64_xor23;
  wire u_CSAwallace_cska32_u_cska64_fa22_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa22_and0;
  wire u_CSAwallace_cska32_u_cska64_fa22_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa22_and1;
  wire u_CSAwallace_cska32_u_cska64_fa22_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate515;
  wire u_CSAwallace_cska32_u_cska64_and_propagate516;
  wire u_CSAwallace_cska32_u_cska64_and_propagate517;
  wire u_CSAwallace_cska32_u_cska64_mux2to15_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to15_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to15_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to15_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor24;
  wire u_CSAwallace_cska32_u_cska64_fa23_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa23_and0;
  wire u_CSAwallace_cska32_u_cska64_fa23_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa23_and1;
  wire u_CSAwallace_cska32_u_cska64_fa23_or0;
  wire u_CSAwallace_cska32_u_cska64_xor25;
  wire u_CSAwallace_cska32_u_cska64_fa24_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa24_and0;
  wire u_CSAwallace_cska32_u_cska64_fa24_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa24_and1;
  wire u_CSAwallace_cska32_u_cska64_fa24_or0;
  wire u_CSAwallace_cska32_u_cska64_xor26;
  wire u_CSAwallace_cska32_u_cska64_fa25_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa25_and0;
  wire u_CSAwallace_cska32_u_cska64_fa25_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa25_and1;
  wire u_CSAwallace_cska32_u_cska64_fa25_or0;
  wire u_CSAwallace_cska32_u_cska64_xor27;
  wire u_CSAwallace_cska32_u_cska64_fa26_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa26_and0;
  wire u_CSAwallace_cska32_u_cska64_fa26_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa26_and1;
  wire u_CSAwallace_cska32_u_cska64_fa26_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate618;
  wire u_CSAwallace_cska32_u_cska64_and_propagate619;
  wire u_CSAwallace_cska32_u_cska64_and_propagate620;
  wire u_CSAwallace_cska32_u_cska64_mux2to16_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to16_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to16_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to16_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor28;
  wire u_CSAwallace_cska32_u_cska64_fa27_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa27_and0;
  wire u_CSAwallace_cska32_u_cska64_fa27_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa27_and1;
  wire u_CSAwallace_cska32_u_cska64_fa27_or0;
  wire u_CSAwallace_cska32_u_cska64_xor29;
  wire u_CSAwallace_cska32_u_cska64_fa28_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa28_and0;
  wire u_CSAwallace_cska32_u_cska64_fa28_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa28_and1;
  wire u_CSAwallace_cska32_u_cska64_fa28_or0;
  wire u_CSAwallace_cska32_u_cska64_xor30;
  wire u_CSAwallace_cska32_u_cska64_fa29_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa29_and0;
  wire u_CSAwallace_cska32_u_cska64_fa29_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa29_and1;
  wire u_CSAwallace_cska32_u_cska64_fa29_or0;
  wire u_CSAwallace_cska32_u_cska64_xor31;
  wire u_CSAwallace_cska32_u_cska64_fa30_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa30_and0;
  wire u_CSAwallace_cska32_u_cska64_fa30_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa30_and1;
  wire u_CSAwallace_cska32_u_cska64_fa30_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate721;
  wire u_CSAwallace_cska32_u_cska64_and_propagate722;
  wire u_CSAwallace_cska32_u_cska64_and_propagate723;
  wire u_CSAwallace_cska32_u_cska64_mux2to17_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to17_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to17_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to17_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor32;
  wire u_CSAwallace_cska32_u_cska64_fa31_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa31_and0;
  wire u_CSAwallace_cska32_u_cska64_fa31_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa31_and1;
  wire u_CSAwallace_cska32_u_cska64_fa31_or0;
  wire u_CSAwallace_cska32_u_cska64_xor33;
  wire u_CSAwallace_cska32_u_cska64_fa32_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa32_and0;
  wire u_CSAwallace_cska32_u_cska64_fa32_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa32_and1;
  wire u_CSAwallace_cska32_u_cska64_fa32_or0;
  wire u_CSAwallace_cska32_u_cska64_xor34;
  wire u_CSAwallace_cska32_u_cska64_fa33_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa33_and0;
  wire u_CSAwallace_cska32_u_cska64_fa33_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa33_and1;
  wire u_CSAwallace_cska32_u_cska64_fa33_or0;
  wire u_CSAwallace_cska32_u_cska64_xor35;
  wire u_CSAwallace_cska32_u_cska64_fa34_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa34_and0;
  wire u_CSAwallace_cska32_u_cska64_fa34_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa34_and1;
  wire u_CSAwallace_cska32_u_cska64_fa34_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate824;
  wire u_CSAwallace_cska32_u_cska64_and_propagate825;
  wire u_CSAwallace_cska32_u_cska64_and_propagate826;
  wire u_CSAwallace_cska32_u_cska64_mux2to18_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to18_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to18_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to18_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor36;
  wire u_CSAwallace_cska32_u_cska64_fa35_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa35_and0;
  wire u_CSAwallace_cska32_u_cska64_fa35_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa35_and1;
  wire u_CSAwallace_cska32_u_cska64_fa35_or0;
  wire u_CSAwallace_cska32_u_cska64_xor37;
  wire u_CSAwallace_cska32_u_cska64_fa36_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa36_and0;
  wire u_CSAwallace_cska32_u_cska64_fa36_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa36_and1;
  wire u_CSAwallace_cska32_u_cska64_fa36_or0;
  wire u_CSAwallace_cska32_u_cska64_xor38;
  wire u_CSAwallace_cska32_u_cska64_fa37_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa37_and0;
  wire u_CSAwallace_cska32_u_cska64_fa37_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa37_and1;
  wire u_CSAwallace_cska32_u_cska64_fa37_or0;
  wire u_CSAwallace_cska32_u_cska64_xor39;
  wire u_CSAwallace_cska32_u_cska64_fa38_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa38_and0;
  wire u_CSAwallace_cska32_u_cska64_fa38_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa38_and1;
  wire u_CSAwallace_cska32_u_cska64_fa38_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate927;
  wire u_CSAwallace_cska32_u_cska64_and_propagate928;
  wire u_CSAwallace_cska32_u_cska64_and_propagate929;
  wire u_CSAwallace_cska32_u_cska64_mux2to19_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to19_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to19_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to19_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor40;
  wire u_CSAwallace_cska32_u_cska64_fa39_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa39_and0;
  wire u_CSAwallace_cska32_u_cska64_fa39_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa39_and1;
  wire u_CSAwallace_cska32_u_cska64_fa39_or0;
  wire u_CSAwallace_cska32_u_cska64_xor41;
  wire u_CSAwallace_cska32_u_cska64_fa40_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa40_and0;
  wire u_CSAwallace_cska32_u_cska64_fa40_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa40_and1;
  wire u_CSAwallace_cska32_u_cska64_fa40_or0;
  wire u_CSAwallace_cska32_u_cska64_xor42;
  wire u_CSAwallace_cska32_u_cska64_fa41_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa41_and0;
  wire u_CSAwallace_cska32_u_cska64_fa41_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa41_and1;
  wire u_CSAwallace_cska32_u_cska64_fa41_or0;
  wire u_CSAwallace_cska32_u_cska64_xor43;
  wire u_CSAwallace_cska32_u_cska64_fa42_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa42_and0;
  wire u_CSAwallace_cska32_u_cska64_fa42_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa42_and1;
  wire u_CSAwallace_cska32_u_cska64_fa42_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1030;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1031;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1032;
  wire u_CSAwallace_cska32_u_cska64_mux2to110_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to110_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to110_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to110_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor44;
  wire u_CSAwallace_cska32_u_cska64_fa43_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa43_and0;
  wire u_CSAwallace_cska32_u_cska64_fa43_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa43_and1;
  wire u_CSAwallace_cska32_u_cska64_fa43_or0;
  wire u_CSAwallace_cska32_u_cska64_xor45;
  wire u_CSAwallace_cska32_u_cska64_fa44_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa44_and0;
  wire u_CSAwallace_cska32_u_cska64_fa44_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa44_and1;
  wire u_CSAwallace_cska32_u_cska64_fa44_or0;
  wire u_CSAwallace_cska32_u_cska64_xor46;
  wire u_CSAwallace_cska32_u_cska64_fa45_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa45_and0;
  wire u_CSAwallace_cska32_u_cska64_fa45_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa45_and1;
  wire u_CSAwallace_cska32_u_cska64_fa45_or0;
  wire u_CSAwallace_cska32_u_cska64_xor47;
  wire u_CSAwallace_cska32_u_cska64_fa46_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa46_and0;
  wire u_CSAwallace_cska32_u_cska64_fa46_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa46_and1;
  wire u_CSAwallace_cska32_u_cska64_fa46_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1133;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1134;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1135;
  wire u_CSAwallace_cska32_u_cska64_mux2to111_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to111_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to111_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to111_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor48;
  wire u_CSAwallace_cska32_u_cska64_fa47_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa47_and0;
  wire u_CSAwallace_cska32_u_cska64_fa47_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa47_and1;
  wire u_CSAwallace_cska32_u_cska64_fa47_or0;
  wire u_CSAwallace_cska32_u_cska64_xor49;
  wire u_CSAwallace_cska32_u_cska64_fa48_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa48_and0;
  wire u_CSAwallace_cska32_u_cska64_fa48_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa48_and1;
  wire u_CSAwallace_cska32_u_cska64_fa48_or0;
  wire u_CSAwallace_cska32_u_cska64_xor50;
  wire u_CSAwallace_cska32_u_cska64_fa49_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa49_and0;
  wire u_CSAwallace_cska32_u_cska64_fa49_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa49_and1;
  wire u_CSAwallace_cska32_u_cska64_fa49_or0;
  wire u_CSAwallace_cska32_u_cska64_xor51;
  wire u_CSAwallace_cska32_u_cska64_fa50_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa50_and0;
  wire u_CSAwallace_cska32_u_cska64_fa50_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa50_and1;
  wire u_CSAwallace_cska32_u_cska64_fa50_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1236;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1237;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1238;
  wire u_CSAwallace_cska32_u_cska64_mux2to112_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to112_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to112_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to112_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor52;
  wire u_CSAwallace_cska32_u_cska64_fa51_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa51_and0;
  wire u_CSAwallace_cska32_u_cska64_fa51_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa51_and1;
  wire u_CSAwallace_cska32_u_cska64_fa51_or0;
  wire u_CSAwallace_cska32_u_cska64_xor53;
  wire u_CSAwallace_cska32_u_cska64_fa52_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa52_and0;
  wire u_CSAwallace_cska32_u_cska64_fa52_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa52_and1;
  wire u_CSAwallace_cska32_u_cska64_fa52_or0;
  wire u_CSAwallace_cska32_u_cska64_xor54;
  wire u_CSAwallace_cska32_u_cska64_fa53_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa53_and0;
  wire u_CSAwallace_cska32_u_cska64_fa53_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa53_and1;
  wire u_CSAwallace_cska32_u_cska64_fa53_or0;
  wire u_CSAwallace_cska32_u_cska64_xor55;
  wire u_CSAwallace_cska32_u_cska64_fa54_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa54_and0;
  wire u_CSAwallace_cska32_u_cska64_fa54_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa54_and1;
  wire u_CSAwallace_cska32_u_cska64_fa54_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1339;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1340;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1341;
  wire u_CSAwallace_cska32_u_cska64_mux2to113_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to113_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to113_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to113_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor56;
  wire u_CSAwallace_cska32_u_cska64_fa55_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa55_and0;
  wire u_CSAwallace_cska32_u_cska64_fa55_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa55_and1;
  wire u_CSAwallace_cska32_u_cska64_fa55_or0;
  wire u_CSAwallace_cska32_u_cska64_xor57;
  wire u_CSAwallace_cska32_u_cska64_fa56_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa56_and0;
  wire u_CSAwallace_cska32_u_cska64_fa56_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa56_and1;
  wire u_CSAwallace_cska32_u_cska64_fa56_or0;
  wire u_CSAwallace_cska32_u_cska64_xor58;
  wire u_CSAwallace_cska32_u_cska64_fa57_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa57_and0;
  wire u_CSAwallace_cska32_u_cska64_fa57_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa57_and1;
  wire u_CSAwallace_cska32_u_cska64_fa57_or0;
  wire u_CSAwallace_cska32_u_cska64_xor59;
  wire u_CSAwallace_cska32_u_cska64_fa58_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa58_and0;
  wire u_CSAwallace_cska32_u_cska64_fa58_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa58_and1;
  wire u_CSAwallace_cska32_u_cska64_fa58_or0;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1442;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1443;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1444;
  wire u_CSAwallace_cska32_u_cska64_mux2to114_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to114_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to114_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to114_xor0;
  wire u_CSAwallace_cska32_u_cska64_xor60;
  wire u_CSAwallace_cska32_u_cska64_fa59_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa59_and0;
  wire u_CSAwallace_cska32_u_cska64_fa59_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa59_and1;
  wire u_CSAwallace_cska32_u_cska64_fa59_or0;
  wire u_CSAwallace_cska32_u_cska64_xor61;
  wire u_CSAwallace_cska32_u_cska64_fa60_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa60_and0;
  wire u_CSAwallace_cska32_u_cska64_fa60_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa60_and1;
  wire u_CSAwallace_cska32_u_cska64_fa60_or0;
  wire u_CSAwallace_cska32_u_cska64_xor62;
  wire u_CSAwallace_cska32_u_cska64_fa61_xor0;
  wire u_CSAwallace_cska32_u_cska64_fa61_and0;
  wire u_CSAwallace_cska32_u_cska64_fa61_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa61_and1;
  wire u_CSAwallace_cska32_u_cska64_fa61_or0;
  wire u_CSAwallace_cska32_u_cska64_fa62_xor1;
  wire u_CSAwallace_cska32_u_cska64_fa62_and1;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1545;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1546;
  wire u_CSAwallace_cska32_u_cska64_and_propagate1547;
  wire u_CSAwallace_cska32_u_cska64_mux2to115_and0;
  wire u_CSAwallace_cska32_u_cska64_mux2to115_not0;
  wire u_CSAwallace_cska32_u_cska64_mux2to115_and1;
  wire u_CSAwallace_cska32_u_cska64_mux2to115_xor0;

  assign u_CSAwallace_cska32_and_0_0 = a[0] & b[0];
  assign u_CSAwallace_cska32_and_1_0 = a[1] & b[0];
  assign u_CSAwallace_cska32_and_2_0 = a[2] & b[0];
  assign u_CSAwallace_cska32_and_3_0 = a[3] & b[0];
  assign u_CSAwallace_cska32_and_4_0 = a[4] & b[0];
  assign u_CSAwallace_cska32_and_5_0 = a[5] & b[0];
  assign u_CSAwallace_cska32_and_6_0 = a[6] & b[0];
  assign u_CSAwallace_cska32_and_7_0 = a[7] & b[0];
  assign u_CSAwallace_cska32_and_8_0 = a[8] & b[0];
  assign u_CSAwallace_cska32_and_9_0 = a[9] & b[0];
  assign u_CSAwallace_cska32_and_10_0 = a[10] & b[0];
  assign u_CSAwallace_cska32_and_11_0 = a[11] & b[0];
  assign u_CSAwallace_cska32_and_12_0 = a[12] & b[0];
  assign u_CSAwallace_cska32_and_13_0 = a[13] & b[0];
  assign u_CSAwallace_cska32_and_14_0 = a[14] & b[0];
  assign u_CSAwallace_cska32_and_15_0 = a[15] & b[0];
  assign u_CSAwallace_cska32_and_16_0 = a[16] & b[0];
  assign u_CSAwallace_cska32_and_17_0 = a[17] & b[0];
  assign u_CSAwallace_cska32_and_18_0 = a[18] & b[0];
  assign u_CSAwallace_cska32_and_19_0 = a[19] & b[0];
  assign u_CSAwallace_cska32_and_20_0 = a[20] & b[0];
  assign u_CSAwallace_cska32_and_21_0 = a[21] & b[0];
  assign u_CSAwallace_cska32_and_22_0 = a[22] & b[0];
  assign u_CSAwallace_cska32_and_23_0 = a[23] & b[0];
  assign u_CSAwallace_cska32_and_24_0 = a[24] & b[0];
  assign u_CSAwallace_cska32_and_25_0 = a[25] & b[0];
  assign u_CSAwallace_cska32_and_26_0 = a[26] & b[0];
  assign u_CSAwallace_cska32_and_27_0 = a[27] & b[0];
  assign u_CSAwallace_cska32_and_28_0 = a[28] & b[0];
  assign u_CSAwallace_cska32_and_29_0 = a[29] & b[0];
  assign u_CSAwallace_cska32_and_30_0 = a[30] & b[0];
  assign u_CSAwallace_cska32_and_31_0 = a[31] & b[0];
  assign u_CSAwallace_cska32_and_0_1 = a[0] & b[1];
  assign u_CSAwallace_cska32_and_1_1 = a[1] & b[1];
  assign u_CSAwallace_cska32_and_2_1 = a[2] & b[1];
  assign u_CSAwallace_cska32_and_3_1 = a[3] & b[1];
  assign u_CSAwallace_cska32_and_4_1 = a[4] & b[1];
  assign u_CSAwallace_cska32_and_5_1 = a[5] & b[1];
  assign u_CSAwallace_cska32_and_6_1 = a[6] & b[1];
  assign u_CSAwallace_cska32_and_7_1 = a[7] & b[1];
  assign u_CSAwallace_cska32_and_8_1 = a[8] & b[1];
  assign u_CSAwallace_cska32_and_9_1 = a[9] & b[1];
  assign u_CSAwallace_cska32_and_10_1 = a[10] & b[1];
  assign u_CSAwallace_cska32_and_11_1 = a[11] & b[1];
  assign u_CSAwallace_cska32_and_12_1 = a[12] & b[1];
  assign u_CSAwallace_cska32_and_13_1 = a[13] & b[1];
  assign u_CSAwallace_cska32_and_14_1 = a[14] & b[1];
  assign u_CSAwallace_cska32_and_15_1 = a[15] & b[1];
  assign u_CSAwallace_cska32_and_16_1 = a[16] & b[1];
  assign u_CSAwallace_cska32_and_17_1 = a[17] & b[1];
  assign u_CSAwallace_cska32_and_18_1 = a[18] & b[1];
  assign u_CSAwallace_cska32_and_19_1 = a[19] & b[1];
  assign u_CSAwallace_cska32_and_20_1 = a[20] & b[1];
  assign u_CSAwallace_cska32_and_21_1 = a[21] & b[1];
  assign u_CSAwallace_cska32_and_22_1 = a[22] & b[1];
  assign u_CSAwallace_cska32_and_23_1 = a[23] & b[1];
  assign u_CSAwallace_cska32_and_24_1 = a[24] & b[1];
  assign u_CSAwallace_cska32_and_25_1 = a[25] & b[1];
  assign u_CSAwallace_cska32_and_26_1 = a[26] & b[1];
  assign u_CSAwallace_cska32_and_27_1 = a[27] & b[1];
  assign u_CSAwallace_cska32_and_28_1 = a[28] & b[1];
  assign u_CSAwallace_cska32_and_29_1 = a[29] & b[1];
  assign u_CSAwallace_cska32_and_30_1 = a[30] & b[1];
  assign u_CSAwallace_cska32_and_31_1 = a[31] & b[1];
  assign u_CSAwallace_cska32_and_0_2 = a[0] & b[2];
  assign u_CSAwallace_cska32_and_1_2 = a[1] & b[2];
  assign u_CSAwallace_cska32_and_2_2 = a[2] & b[2];
  assign u_CSAwallace_cska32_and_3_2 = a[3] & b[2];
  assign u_CSAwallace_cska32_and_4_2 = a[4] & b[2];
  assign u_CSAwallace_cska32_and_5_2 = a[5] & b[2];
  assign u_CSAwallace_cska32_and_6_2 = a[6] & b[2];
  assign u_CSAwallace_cska32_and_7_2 = a[7] & b[2];
  assign u_CSAwallace_cska32_and_8_2 = a[8] & b[2];
  assign u_CSAwallace_cska32_and_9_2 = a[9] & b[2];
  assign u_CSAwallace_cska32_and_10_2 = a[10] & b[2];
  assign u_CSAwallace_cska32_and_11_2 = a[11] & b[2];
  assign u_CSAwallace_cska32_and_12_2 = a[12] & b[2];
  assign u_CSAwallace_cska32_and_13_2 = a[13] & b[2];
  assign u_CSAwallace_cska32_and_14_2 = a[14] & b[2];
  assign u_CSAwallace_cska32_and_15_2 = a[15] & b[2];
  assign u_CSAwallace_cska32_and_16_2 = a[16] & b[2];
  assign u_CSAwallace_cska32_and_17_2 = a[17] & b[2];
  assign u_CSAwallace_cska32_and_18_2 = a[18] & b[2];
  assign u_CSAwallace_cska32_and_19_2 = a[19] & b[2];
  assign u_CSAwallace_cska32_and_20_2 = a[20] & b[2];
  assign u_CSAwallace_cska32_and_21_2 = a[21] & b[2];
  assign u_CSAwallace_cska32_and_22_2 = a[22] & b[2];
  assign u_CSAwallace_cska32_and_23_2 = a[23] & b[2];
  assign u_CSAwallace_cska32_and_24_2 = a[24] & b[2];
  assign u_CSAwallace_cska32_and_25_2 = a[25] & b[2];
  assign u_CSAwallace_cska32_and_26_2 = a[26] & b[2];
  assign u_CSAwallace_cska32_and_27_2 = a[27] & b[2];
  assign u_CSAwallace_cska32_and_28_2 = a[28] & b[2];
  assign u_CSAwallace_cska32_and_29_2 = a[29] & b[2];
  assign u_CSAwallace_cska32_and_30_2 = a[30] & b[2];
  assign u_CSAwallace_cska32_and_31_2 = a[31] & b[2];
  assign u_CSAwallace_cska32_and_0_3 = a[0] & b[3];
  assign u_CSAwallace_cska32_and_1_3 = a[1] & b[3];
  assign u_CSAwallace_cska32_and_2_3 = a[2] & b[3];
  assign u_CSAwallace_cska32_and_3_3 = a[3] & b[3];
  assign u_CSAwallace_cska32_and_4_3 = a[4] & b[3];
  assign u_CSAwallace_cska32_and_5_3 = a[5] & b[3];
  assign u_CSAwallace_cska32_and_6_3 = a[6] & b[3];
  assign u_CSAwallace_cska32_and_7_3 = a[7] & b[3];
  assign u_CSAwallace_cska32_and_8_3 = a[8] & b[3];
  assign u_CSAwallace_cska32_and_9_3 = a[9] & b[3];
  assign u_CSAwallace_cska32_and_10_3 = a[10] & b[3];
  assign u_CSAwallace_cska32_and_11_3 = a[11] & b[3];
  assign u_CSAwallace_cska32_and_12_3 = a[12] & b[3];
  assign u_CSAwallace_cska32_and_13_3 = a[13] & b[3];
  assign u_CSAwallace_cska32_and_14_3 = a[14] & b[3];
  assign u_CSAwallace_cska32_and_15_3 = a[15] & b[3];
  assign u_CSAwallace_cska32_and_16_3 = a[16] & b[3];
  assign u_CSAwallace_cska32_and_17_3 = a[17] & b[3];
  assign u_CSAwallace_cska32_and_18_3 = a[18] & b[3];
  assign u_CSAwallace_cska32_and_19_3 = a[19] & b[3];
  assign u_CSAwallace_cska32_and_20_3 = a[20] & b[3];
  assign u_CSAwallace_cska32_and_21_3 = a[21] & b[3];
  assign u_CSAwallace_cska32_and_22_3 = a[22] & b[3];
  assign u_CSAwallace_cska32_and_23_3 = a[23] & b[3];
  assign u_CSAwallace_cska32_and_24_3 = a[24] & b[3];
  assign u_CSAwallace_cska32_and_25_3 = a[25] & b[3];
  assign u_CSAwallace_cska32_and_26_3 = a[26] & b[3];
  assign u_CSAwallace_cska32_and_27_3 = a[27] & b[3];
  assign u_CSAwallace_cska32_and_28_3 = a[28] & b[3];
  assign u_CSAwallace_cska32_and_29_3 = a[29] & b[3];
  assign u_CSAwallace_cska32_and_30_3 = a[30] & b[3];
  assign u_CSAwallace_cska32_and_31_3 = a[31] & b[3];
  assign u_CSAwallace_cska32_and_0_4 = a[0] & b[4];
  assign u_CSAwallace_cska32_and_1_4 = a[1] & b[4];
  assign u_CSAwallace_cska32_and_2_4 = a[2] & b[4];
  assign u_CSAwallace_cska32_and_3_4 = a[3] & b[4];
  assign u_CSAwallace_cska32_and_4_4 = a[4] & b[4];
  assign u_CSAwallace_cska32_and_5_4 = a[5] & b[4];
  assign u_CSAwallace_cska32_and_6_4 = a[6] & b[4];
  assign u_CSAwallace_cska32_and_7_4 = a[7] & b[4];
  assign u_CSAwallace_cska32_and_8_4 = a[8] & b[4];
  assign u_CSAwallace_cska32_and_9_4 = a[9] & b[4];
  assign u_CSAwallace_cska32_and_10_4 = a[10] & b[4];
  assign u_CSAwallace_cska32_and_11_4 = a[11] & b[4];
  assign u_CSAwallace_cska32_and_12_4 = a[12] & b[4];
  assign u_CSAwallace_cska32_and_13_4 = a[13] & b[4];
  assign u_CSAwallace_cska32_and_14_4 = a[14] & b[4];
  assign u_CSAwallace_cska32_and_15_4 = a[15] & b[4];
  assign u_CSAwallace_cska32_and_16_4 = a[16] & b[4];
  assign u_CSAwallace_cska32_and_17_4 = a[17] & b[4];
  assign u_CSAwallace_cska32_and_18_4 = a[18] & b[4];
  assign u_CSAwallace_cska32_and_19_4 = a[19] & b[4];
  assign u_CSAwallace_cska32_and_20_4 = a[20] & b[4];
  assign u_CSAwallace_cska32_and_21_4 = a[21] & b[4];
  assign u_CSAwallace_cska32_and_22_4 = a[22] & b[4];
  assign u_CSAwallace_cska32_and_23_4 = a[23] & b[4];
  assign u_CSAwallace_cska32_and_24_4 = a[24] & b[4];
  assign u_CSAwallace_cska32_and_25_4 = a[25] & b[4];
  assign u_CSAwallace_cska32_and_26_4 = a[26] & b[4];
  assign u_CSAwallace_cska32_and_27_4 = a[27] & b[4];
  assign u_CSAwallace_cska32_and_28_4 = a[28] & b[4];
  assign u_CSAwallace_cska32_and_29_4 = a[29] & b[4];
  assign u_CSAwallace_cska32_and_30_4 = a[30] & b[4];
  assign u_CSAwallace_cska32_and_31_4 = a[31] & b[4];
  assign u_CSAwallace_cska32_and_0_5 = a[0] & b[5];
  assign u_CSAwallace_cska32_and_1_5 = a[1] & b[5];
  assign u_CSAwallace_cska32_and_2_5 = a[2] & b[5];
  assign u_CSAwallace_cska32_and_3_5 = a[3] & b[5];
  assign u_CSAwallace_cska32_and_4_5 = a[4] & b[5];
  assign u_CSAwallace_cska32_and_5_5 = a[5] & b[5];
  assign u_CSAwallace_cska32_and_6_5 = a[6] & b[5];
  assign u_CSAwallace_cska32_and_7_5 = a[7] & b[5];
  assign u_CSAwallace_cska32_and_8_5 = a[8] & b[5];
  assign u_CSAwallace_cska32_and_9_5 = a[9] & b[5];
  assign u_CSAwallace_cska32_and_10_5 = a[10] & b[5];
  assign u_CSAwallace_cska32_and_11_5 = a[11] & b[5];
  assign u_CSAwallace_cska32_and_12_5 = a[12] & b[5];
  assign u_CSAwallace_cska32_and_13_5 = a[13] & b[5];
  assign u_CSAwallace_cska32_and_14_5 = a[14] & b[5];
  assign u_CSAwallace_cska32_and_15_5 = a[15] & b[5];
  assign u_CSAwallace_cska32_and_16_5 = a[16] & b[5];
  assign u_CSAwallace_cska32_and_17_5 = a[17] & b[5];
  assign u_CSAwallace_cska32_and_18_5 = a[18] & b[5];
  assign u_CSAwallace_cska32_and_19_5 = a[19] & b[5];
  assign u_CSAwallace_cska32_and_20_5 = a[20] & b[5];
  assign u_CSAwallace_cska32_and_21_5 = a[21] & b[5];
  assign u_CSAwallace_cska32_and_22_5 = a[22] & b[5];
  assign u_CSAwallace_cska32_and_23_5 = a[23] & b[5];
  assign u_CSAwallace_cska32_and_24_5 = a[24] & b[5];
  assign u_CSAwallace_cska32_and_25_5 = a[25] & b[5];
  assign u_CSAwallace_cska32_and_26_5 = a[26] & b[5];
  assign u_CSAwallace_cska32_and_27_5 = a[27] & b[5];
  assign u_CSAwallace_cska32_and_28_5 = a[28] & b[5];
  assign u_CSAwallace_cska32_and_29_5 = a[29] & b[5];
  assign u_CSAwallace_cska32_and_30_5 = a[30] & b[5];
  assign u_CSAwallace_cska32_and_31_5 = a[31] & b[5];
  assign u_CSAwallace_cska32_and_0_6 = a[0] & b[6];
  assign u_CSAwallace_cska32_and_1_6 = a[1] & b[6];
  assign u_CSAwallace_cska32_and_2_6 = a[2] & b[6];
  assign u_CSAwallace_cska32_and_3_6 = a[3] & b[6];
  assign u_CSAwallace_cska32_and_4_6 = a[4] & b[6];
  assign u_CSAwallace_cska32_and_5_6 = a[5] & b[6];
  assign u_CSAwallace_cska32_and_6_6 = a[6] & b[6];
  assign u_CSAwallace_cska32_and_7_6 = a[7] & b[6];
  assign u_CSAwallace_cska32_and_8_6 = a[8] & b[6];
  assign u_CSAwallace_cska32_and_9_6 = a[9] & b[6];
  assign u_CSAwallace_cska32_and_10_6 = a[10] & b[6];
  assign u_CSAwallace_cska32_and_11_6 = a[11] & b[6];
  assign u_CSAwallace_cska32_and_12_6 = a[12] & b[6];
  assign u_CSAwallace_cska32_and_13_6 = a[13] & b[6];
  assign u_CSAwallace_cska32_and_14_6 = a[14] & b[6];
  assign u_CSAwallace_cska32_and_15_6 = a[15] & b[6];
  assign u_CSAwallace_cska32_and_16_6 = a[16] & b[6];
  assign u_CSAwallace_cska32_and_17_6 = a[17] & b[6];
  assign u_CSAwallace_cska32_and_18_6 = a[18] & b[6];
  assign u_CSAwallace_cska32_and_19_6 = a[19] & b[6];
  assign u_CSAwallace_cska32_and_20_6 = a[20] & b[6];
  assign u_CSAwallace_cska32_and_21_6 = a[21] & b[6];
  assign u_CSAwallace_cska32_and_22_6 = a[22] & b[6];
  assign u_CSAwallace_cska32_and_23_6 = a[23] & b[6];
  assign u_CSAwallace_cska32_and_24_6 = a[24] & b[6];
  assign u_CSAwallace_cska32_and_25_6 = a[25] & b[6];
  assign u_CSAwallace_cska32_and_26_6 = a[26] & b[6];
  assign u_CSAwallace_cska32_and_27_6 = a[27] & b[6];
  assign u_CSAwallace_cska32_and_28_6 = a[28] & b[6];
  assign u_CSAwallace_cska32_and_29_6 = a[29] & b[6];
  assign u_CSAwallace_cska32_and_30_6 = a[30] & b[6];
  assign u_CSAwallace_cska32_and_31_6 = a[31] & b[6];
  assign u_CSAwallace_cska32_and_0_7 = a[0] & b[7];
  assign u_CSAwallace_cska32_and_1_7 = a[1] & b[7];
  assign u_CSAwallace_cska32_and_2_7 = a[2] & b[7];
  assign u_CSAwallace_cska32_and_3_7 = a[3] & b[7];
  assign u_CSAwallace_cska32_and_4_7 = a[4] & b[7];
  assign u_CSAwallace_cska32_and_5_7 = a[5] & b[7];
  assign u_CSAwallace_cska32_and_6_7 = a[6] & b[7];
  assign u_CSAwallace_cska32_and_7_7 = a[7] & b[7];
  assign u_CSAwallace_cska32_and_8_7 = a[8] & b[7];
  assign u_CSAwallace_cska32_and_9_7 = a[9] & b[7];
  assign u_CSAwallace_cska32_and_10_7 = a[10] & b[7];
  assign u_CSAwallace_cska32_and_11_7 = a[11] & b[7];
  assign u_CSAwallace_cska32_and_12_7 = a[12] & b[7];
  assign u_CSAwallace_cska32_and_13_7 = a[13] & b[7];
  assign u_CSAwallace_cska32_and_14_7 = a[14] & b[7];
  assign u_CSAwallace_cska32_and_15_7 = a[15] & b[7];
  assign u_CSAwallace_cska32_and_16_7 = a[16] & b[7];
  assign u_CSAwallace_cska32_and_17_7 = a[17] & b[7];
  assign u_CSAwallace_cska32_and_18_7 = a[18] & b[7];
  assign u_CSAwallace_cska32_and_19_7 = a[19] & b[7];
  assign u_CSAwallace_cska32_and_20_7 = a[20] & b[7];
  assign u_CSAwallace_cska32_and_21_7 = a[21] & b[7];
  assign u_CSAwallace_cska32_and_22_7 = a[22] & b[7];
  assign u_CSAwallace_cska32_and_23_7 = a[23] & b[7];
  assign u_CSAwallace_cska32_and_24_7 = a[24] & b[7];
  assign u_CSAwallace_cska32_and_25_7 = a[25] & b[7];
  assign u_CSAwallace_cska32_and_26_7 = a[26] & b[7];
  assign u_CSAwallace_cska32_and_27_7 = a[27] & b[7];
  assign u_CSAwallace_cska32_and_28_7 = a[28] & b[7];
  assign u_CSAwallace_cska32_and_29_7 = a[29] & b[7];
  assign u_CSAwallace_cska32_and_30_7 = a[30] & b[7];
  assign u_CSAwallace_cska32_and_31_7 = a[31] & b[7];
  assign u_CSAwallace_cska32_and_0_8 = a[0] & b[8];
  assign u_CSAwallace_cska32_and_1_8 = a[1] & b[8];
  assign u_CSAwallace_cska32_and_2_8 = a[2] & b[8];
  assign u_CSAwallace_cska32_and_3_8 = a[3] & b[8];
  assign u_CSAwallace_cska32_and_4_8 = a[4] & b[8];
  assign u_CSAwallace_cska32_and_5_8 = a[5] & b[8];
  assign u_CSAwallace_cska32_and_6_8 = a[6] & b[8];
  assign u_CSAwallace_cska32_and_7_8 = a[7] & b[8];
  assign u_CSAwallace_cska32_and_8_8 = a[8] & b[8];
  assign u_CSAwallace_cska32_and_9_8 = a[9] & b[8];
  assign u_CSAwallace_cska32_and_10_8 = a[10] & b[8];
  assign u_CSAwallace_cska32_and_11_8 = a[11] & b[8];
  assign u_CSAwallace_cska32_and_12_8 = a[12] & b[8];
  assign u_CSAwallace_cska32_and_13_8 = a[13] & b[8];
  assign u_CSAwallace_cska32_and_14_8 = a[14] & b[8];
  assign u_CSAwallace_cska32_and_15_8 = a[15] & b[8];
  assign u_CSAwallace_cska32_and_16_8 = a[16] & b[8];
  assign u_CSAwallace_cska32_and_17_8 = a[17] & b[8];
  assign u_CSAwallace_cska32_and_18_8 = a[18] & b[8];
  assign u_CSAwallace_cska32_and_19_8 = a[19] & b[8];
  assign u_CSAwallace_cska32_and_20_8 = a[20] & b[8];
  assign u_CSAwallace_cska32_and_21_8 = a[21] & b[8];
  assign u_CSAwallace_cska32_and_22_8 = a[22] & b[8];
  assign u_CSAwallace_cska32_and_23_8 = a[23] & b[8];
  assign u_CSAwallace_cska32_and_24_8 = a[24] & b[8];
  assign u_CSAwallace_cska32_and_25_8 = a[25] & b[8];
  assign u_CSAwallace_cska32_and_26_8 = a[26] & b[8];
  assign u_CSAwallace_cska32_and_27_8 = a[27] & b[8];
  assign u_CSAwallace_cska32_and_28_8 = a[28] & b[8];
  assign u_CSAwallace_cska32_and_29_8 = a[29] & b[8];
  assign u_CSAwallace_cska32_and_30_8 = a[30] & b[8];
  assign u_CSAwallace_cska32_and_31_8 = a[31] & b[8];
  assign u_CSAwallace_cska32_and_0_9 = a[0] & b[9];
  assign u_CSAwallace_cska32_and_1_9 = a[1] & b[9];
  assign u_CSAwallace_cska32_and_2_9 = a[2] & b[9];
  assign u_CSAwallace_cska32_and_3_9 = a[3] & b[9];
  assign u_CSAwallace_cska32_and_4_9 = a[4] & b[9];
  assign u_CSAwallace_cska32_and_5_9 = a[5] & b[9];
  assign u_CSAwallace_cska32_and_6_9 = a[6] & b[9];
  assign u_CSAwallace_cska32_and_7_9 = a[7] & b[9];
  assign u_CSAwallace_cska32_and_8_9 = a[8] & b[9];
  assign u_CSAwallace_cska32_and_9_9 = a[9] & b[9];
  assign u_CSAwallace_cska32_and_10_9 = a[10] & b[9];
  assign u_CSAwallace_cska32_and_11_9 = a[11] & b[9];
  assign u_CSAwallace_cska32_and_12_9 = a[12] & b[9];
  assign u_CSAwallace_cska32_and_13_9 = a[13] & b[9];
  assign u_CSAwallace_cska32_and_14_9 = a[14] & b[9];
  assign u_CSAwallace_cska32_and_15_9 = a[15] & b[9];
  assign u_CSAwallace_cska32_and_16_9 = a[16] & b[9];
  assign u_CSAwallace_cska32_and_17_9 = a[17] & b[9];
  assign u_CSAwallace_cska32_and_18_9 = a[18] & b[9];
  assign u_CSAwallace_cska32_and_19_9 = a[19] & b[9];
  assign u_CSAwallace_cska32_and_20_9 = a[20] & b[9];
  assign u_CSAwallace_cska32_and_21_9 = a[21] & b[9];
  assign u_CSAwallace_cska32_and_22_9 = a[22] & b[9];
  assign u_CSAwallace_cska32_and_23_9 = a[23] & b[9];
  assign u_CSAwallace_cska32_and_24_9 = a[24] & b[9];
  assign u_CSAwallace_cska32_and_25_9 = a[25] & b[9];
  assign u_CSAwallace_cska32_and_26_9 = a[26] & b[9];
  assign u_CSAwallace_cska32_and_27_9 = a[27] & b[9];
  assign u_CSAwallace_cska32_and_28_9 = a[28] & b[9];
  assign u_CSAwallace_cska32_and_29_9 = a[29] & b[9];
  assign u_CSAwallace_cska32_and_30_9 = a[30] & b[9];
  assign u_CSAwallace_cska32_and_31_9 = a[31] & b[9];
  assign u_CSAwallace_cska32_and_0_10 = a[0] & b[10];
  assign u_CSAwallace_cska32_and_1_10 = a[1] & b[10];
  assign u_CSAwallace_cska32_and_2_10 = a[2] & b[10];
  assign u_CSAwallace_cska32_and_3_10 = a[3] & b[10];
  assign u_CSAwallace_cska32_and_4_10 = a[4] & b[10];
  assign u_CSAwallace_cska32_and_5_10 = a[5] & b[10];
  assign u_CSAwallace_cska32_and_6_10 = a[6] & b[10];
  assign u_CSAwallace_cska32_and_7_10 = a[7] & b[10];
  assign u_CSAwallace_cska32_and_8_10 = a[8] & b[10];
  assign u_CSAwallace_cska32_and_9_10 = a[9] & b[10];
  assign u_CSAwallace_cska32_and_10_10 = a[10] & b[10];
  assign u_CSAwallace_cska32_and_11_10 = a[11] & b[10];
  assign u_CSAwallace_cska32_and_12_10 = a[12] & b[10];
  assign u_CSAwallace_cska32_and_13_10 = a[13] & b[10];
  assign u_CSAwallace_cska32_and_14_10 = a[14] & b[10];
  assign u_CSAwallace_cska32_and_15_10 = a[15] & b[10];
  assign u_CSAwallace_cska32_and_16_10 = a[16] & b[10];
  assign u_CSAwallace_cska32_and_17_10 = a[17] & b[10];
  assign u_CSAwallace_cska32_and_18_10 = a[18] & b[10];
  assign u_CSAwallace_cska32_and_19_10 = a[19] & b[10];
  assign u_CSAwallace_cska32_and_20_10 = a[20] & b[10];
  assign u_CSAwallace_cska32_and_21_10 = a[21] & b[10];
  assign u_CSAwallace_cska32_and_22_10 = a[22] & b[10];
  assign u_CSAwallace_cska32_and_23_10 = a[23] & b[10];
  assign u_CSAwallace_cska32_and_24_10 = a[24] & b[10];
  assign u_CSAwallace_cska32_and_25_10 = a[25] & b[10];
  assign u_CSAwallace_cska32_and_26_10 = a[26] & b[10];
  assign u_CSAwallace_cska32_and_27_10 = a[27] & b[10];
  assign u_CSAwallace_cska32_and_28_10 = a[28] & b[10];
  assign u_CSAwallace_cska32_and_29_10 = a[29] & b[10];
  assign u_CSAwallace_cska32_and_30_10 = a[30] & b[10];
  assign u_CSAwallace_cska32_and_31_10 = a[31] & b[10];
  assign u_CSAwallace_cska32_and_0_11 = a[0] & b[11];
  assign u_CSAwallace_cska32_and_1_11 = a[1] & b[11];
  assign u_CSAwallace_cska32_and_2_11 = a[2] & b[11];
  assign u_CSAwallace_cska32_and_3_11 = a[3] & b[11];
  assign u_CSAwallace_cska32_and_4_11 = a[4] & b[11];
  assign u_CSAwallace_cska32_and_5_11 = a[5] & b[11];
  assign u_CSAwallace_cska32_and_6_11 = a[6] & b[11];
  assign u_CSAwallace_cska32_and_7_11 = a[7] & b[11];
  assign u_CSAwallace_cska32_and_8_11 = a[8] & b[11];
  assign u_CSAwallace_cska32_and_9_11 = a[9] & b[11];
  assign u_CSAwallace_cska32_and_10_11 = a[10] & b[11];
  assign u_CSAwallace_cska32_and_11_11 = a[11] & b[11];
  assign u_CSAwallace_cska32_and_12_11 = a[12] & b[11];
  assign u_CSAwallace_cska32_and_13_11 = a[13] & b[11];
  assign u_CSAwallace_cska32_and_14_11 = a[14] & b[11];
  assign u_CSAwallace_cska32_and_15_11 = a[15] & b[11];
  assign u_CSAwallace_cska32_and_16_11 = a[16] & b[11];
  assign u_CSAwallace_cska32_and_17_11 = a[17] & b[11];
  assign u_CSAwallace_cska32_and_18_11 = a[18] & b[11];
  assign u_CSAwallace_cska32_and_19_11 = a[19] & b[11];
  assign u_CSAwallace_cska32_and_20_11 = a[20] & b[11];
  assign u_CSAwallace_cska32_and_21_11 = a[21] & b[11];
  assign u_CSAwallace_cska32_and_22_11 = a[22] & b[11];
  assign u_CSAwallace_cska32_and_23_11 = a[23] & b[11];
  assign u_CSAwallace_cska32_and_24_11 = a[24] & b[11];
  assign u_CSAwallace_cska32_and_25_11 = a[25] & b[11];
  assign u_CSAwallace_cska32_and_26_11 = a[26] & b[11];
  assign u_CSAwallace_cska32_and_27_11 = a[27] & b[11];
  assign u_CSAwallace_cska32_and_28_11 = a[28] & b[11];
  assign u_CSAwallace_cska32_and_29_11 = a[29] & b[11];
  assign u_CSAwallace_cska32_and_30_11 = a[30] & b[11];
  assign u_CSAwallace_cska32_and_31_11 = a[31] & b[11];
  assign u_CSAwallace_cska32_and_0_12 = a[0] & b[12];
  assign u_CSAwallace_cska32_and_1_12 = a[1] & b[12];
  assign u_CSAwallace_cska32_and_2_12 = a[2] & b[12];
  assign u_CSAwallace_cska32_and_3_12 = a[3] & b[12];
  assign u_CSAwallace_cska32_and_4_12 = a[4] & b[12];
  assign u_CSAwallace_cska32_and_5_12 = a[5] & b[12];
  assign u_CSAwallace_cska32_and_6_12 = a[6] & b[12];
  assign u_CSAwallace_cska32_and_7_12 = a[7] & b[12];
  assign u_CSAwallace_cska32_and_8_12 = a[8] & b[12];
  assign u_CSAwallace_cska32_and_9_12 = a[9] & b[12];
  assign u_CSAwallace_cska32_and_10_12 = a[10] & b[12];
  assign u_CSAwallace_cska32_and_11_12 = a[11] & b[12];
  assign u_CSAwallace_cska32_and_12_12 = a[12] & b[12];
  assign u_CSAwallace_cska32_and_13_12 = a[13] & b[12];
  assign u_CSAwallace_cska32_and_14_12 = a[14] & b[12];
  assign u_CSAwallace_cska32_and_15_12 = a[15] & b[12];
  assign u_CSAwallace_cska32_and_16_12 = a[16] & b[12];
  assign u_CSAwallace_cska32_and_17_12 = a[17] & b[12];
  assign u_CSAwallace_cska32_and_18_12 = a[18] & b[12];
  assign u_CSAwallace_cska32_and_19_12 = a[19] & b[12];
  assign u_CSAwallace_cska32_and_20_12 = a[20] & b[12];
  assign u_CSAwallace_cska32_and_21_12 = a[21] & b[12];
  assign u_CSAwallace_cska32_and_22_12 = a[22] & b[12];
  assign u_CSAwallace_cska32_and_23_12 = a[23] & b[12];
  assign u_CSAwallace_cska32_and_24_12 = a[24] & b[12];
  assign u_CSAwallace_cska32_and_25_12 = a[25] & b[12];
  assign u_CSAwallace_cska32_and_26_12 = a[26] & b[12];
  assign u_CSAwallace_cska32_and_27_12 = a[27] & b[12];
  assign u_CSAwallace_cska32_and_28_12 = a[28] & b[12];
  assign u_CSAwallace_cska32_and_29_12 = a[29] & b[12];
  assign u_CSAwallace_cska32_and_30_12 = a[30] & b[12];
  assign u_CSAwallace_cska32_and_31_12 = a[31] & b[12];
  assign u_CSAwallace_cska32_and_0_13 = a[0] & b[13];
  assign u_CSAwallace_cska32_and_1_13 = a[1] & b[13];
  assign u_CSAwallace_cska32_and_2_13 = a[2] & b[13];
  assign u_CSAwallace_cska32_and_3_13 = a[3] & b[13];
  assign u_CSAwallace_cska32_and_4_13 = a[4] & b[13];
  assign u_CSAwallace_cska32_and_5_13 = a[5] & b[13];
  assign u_CSAwallace_cska32_and_6_13 = a[6] & b[13];
  assign u_CSAwallace_cska32_and_7_13 = a[7] & b[13];
  assign u_CSAwallace_cska32_and_8_13 = a[8] & b[13];
  assign u_CSAwallace_cska32_and_9_13 = a[9] & b[13];
  assign u_CSAwallace_cska32_and_10_13 = a[10] & b[13];
  assign u_CSAwallace_cska32_and_11_13 = a[11] & b[13];
  assign u_CSAwallace_cska32_and_12_13 = a[12] & b[13];
  assign u_CSAwallace_cska32_and_13_13 = a[13] & b[13];
  assign u_CSAwallace_cska32_and_14_13 = a[14] & b[13];
  assign u_CSAwallace_cska32_and_15_13 = a[15] & b[13];
  assign u_CSAwallace_cska32_and_16_13 = a[16] & b[13];
  assign u_CSAwallace_cska32_and_17_13 = a[17] & b[13];
  assign u_CSAwallace_cska32_and_18_13 = a[18] & b[13];
  assign u_CSAwallace_cska32_and_19_13 = a[19] & b[13];
  assign u_CSAwallace_cska32_and_20_13 = a[20] & b[13];
  assign u_CSAwallace_cska32_and_21_13 = a[21] & b[13];
  assign u_CSAwallace_cska32_and_22_13 = a[22] & b[13];
  assign u_CSAwallace_cska32_and_23_13 = a[23] & b[13];
  assign u_CSAwallace_cska32_and_24_13 = a[24] & b[13];
  assign u_CSAwallace_cska32_and_25_13 = a[25] & b[13];
  assign u_CSAwallace_cska32_and_26_13 = a[26] & b[13];
  assign u_CSAwallace_cska32_and_27_13 = a[27] & b[13];
  assign u_CSAwallace_cska32_and_28_13 = a[28] & b[13];
  assign u_CSAwallace_cska32_and_29_13 = a[29] & b[13];
  assign u_CSAwallace_cska32_and_30_13 = a[30] & b[13];
  assign u_CSAwallace_cska32_and_31_13 = a[31] & b[13];
  assign u_CSAwallace_cska32_and_0_14 = a[0] & b[14];
  assign u_CSAwallace_cska32_and_1_14 = a[1] & b[14];
  assign u_CSAwallace_cska32_and_2_14 = a[2] & b[14];
  assign u_CSAwallace_cska32_and_3_14 = a[3] & b[14];
  assign u_CSAwallace_cska32_and_4_14 = a[4] & b[14];
  assign u_CSAwallace_cska32_and_5_14 = a[5] & b[14];
  assign u_CSAwallace_cska32_and_6_14 = a[6] & b[14];
  assign u_CSAwallace_cska32_and_7_14 = a[7] & b[14];
  assign u_CSAwallace_cska32_and_8_14 = a[8] & b[14];
  assign u_CSAwallace_cska32_and_9_14 = a[9] & b[14];
  assign u_CSAwallace_cska32_and_10_14 = a[10] & b[14];
  assign u_CSAwallace_cska32_and_11_14 = a[11] & b[14];
  assign u_CSAwallace_cska32_and_12_14 = a[12] & b[14];
  assign u_CSAwallace_cska32_and_13_14 = a[13] & b[14];
  assign u_CSAwallace_cska32_and_14_14 = a[14] & b[14];
  assign u_CSAwallace_cska32_and_15_14 = a[15] & b[14];
  assign u_CSAwallace_cska32_and_16_14 = a[16] & b[14];
  assign u_CSAwallace_cska32_and_17_14 = a[17] & b[14];
  assign u_CSAwallace_cska32_and_18_14 = a[18] & b[14];
  assign u_CSAwallace_cska32_and_19_14 = a[19] & b[14];
  assign u_CSAwallace_cska32_and_20_14 = a[20] & b[14];
  assign u_CSAwallace_cska32_and_21_14 = a[21] & b[14];
  assign u_CSAwallace_cska32_and_22_14 = a[22] & b[14];
  assign u_CSAwallace_cska32_and_23_14 = a[23] & b[14];
  assign u_CSAwallace_cska32_and_24_14 = a[24] & b[14];
  assign u_CSAwallace_cska32_and_25_14 = a[25] & b[14];
  assign u_CSAwallace_cska32_and_26_14 = a[26] & b[14];
  assign u_CSAwallace_cska32_and_27_14 = a[27] & b[14];
  assign u_CSAwallace_cska32_and_28_14 = a[28] & b[14];
  assign u_CSAwallace_cska32_and_29_14 = a[29] & b[14];
  assign u_CSAwallace_cska32_and_30_14 = a[30] & b[14];
  assign u_CSAwallace_cska32_and_31_14 = a[31] & b[14];
  assign u_CSAwallace_cska32_and_0_15 = a[0] & b[15];
  assign u_CSAwallace_cska32_and_1_15 = a[1] & b[15];
  assign u_CSAwallace_cska32_and_2_15 = a[2] & b[15];
  assign u_CSAwallace_cska32_and_3_15 = a[3] & b[15];
  assign u_CSAwallace_cska32_and_4_15 = a[4] & b[15];
  assign u_CSAwallace_cska32_and_5_15 = a[5] & b[15];
  assign u_CSAwallace_cska32_and_6_15 = a[6] & b[15];
  assign u_CSAwallace_cska32_and_7_15 = a[7] & b[15];
  assign u_CSAwallace_cska32_and_8_15 = a[8] & b[15];
  assign u_CSAwallace_cska32_and_9_15 = a[9] & b[15];
  assign u_CSAwallace_cska32_and_10_15 = a[10] & b[15];
  assign u_CSAwallace_cska32_and_11_15 = a[11] & b[15];
  assign u_CSAwallace_cska32_and_12_15 = a[12] & b[15];
  assign u_CSAwallace_cska32_and_13_15 = a[13] & b[15];
  assign u_CSAwallace_cska32_and_14_15 = a[14] & b[15];
  assign u_CSAwallace_cska32_and_15_15 = a[15] & b[15];
  assign u_CSAwallace_cska32_and_16_15 = a[16] & b[15];
  assign u_CSAwallace_cska32_and_17_15 = a[17] & b[15];
  assign u_CSAwallace_cska32_and_18_15 = a[18] & b[15];
  assign u_CSAwallace_cska32_and_19_15 = a[19] & b[15];
  assign u_CSAwallace_cska32_and_20_15 = a[20] & b[15];
  assign u_CSAwallace_cska32_and_21_15 = a[21] & b[15];
  assign u_CSAwallace_cska32_and_22_15 = a[22] & b[15];
  assign u_CSAwallace_cska32_and_23_15 = a[23] & b[15];
  assign u_CSAwallace_cska32_and_24_15 = a[24] & b[15];
  assign u_CSAwallace_cska32_and_25_15 = a[25] & b[15];
  assign u_CSAwallace_cska32_and_26_15 = a[26] & b[15];
  assign u_CSAwallace_cska32_and_27_15 = a[27] & b[15];
  assign u_CSAwallace_cska32_and_28_15 = a[28] & b[15];
  assign u_CSAwallace_cska32_and_29_15 = a[29] & b[15];
  assign u_CSAwallace_cska32_and_30_15 = a[30] & b[15];
  assign u_CSAwallace_cska32_and_31_15 = a[31] & b[15];
  assign u_CSAwallace_cska32_and_0_16 = a[0] & b[16];
  assign u_CSAwallace_cska32_and_1_16 = a[1] & b[16];
  assign u_CSAwallace_cska32_and_2_16 = a[2] & b[16];
  assign u_CSAwallace_cska32_and_3_16 = a[3] & b[16];
  assign u_CSAwallace_cska32_and_4_16 = a[4] & b[16];
  assign u_CSAwallace_cska32_and_5_16 = a[5] & b[16];
  assign u_CSAwallace_cska32_and_6_16 = a[6] & b[16];
  assign u_CSAwallace_cska32_and_7_16 = a[7] & b[16];
  assign u_CSAwallace_cska32_and_8_16 = a[8] & b[16];
  assign u_CSAwallace_cska32_and_9_16 = a[9] & b[16];
  assign u_CSAwallace_cska32_and_10_16 = a[10] & b[16];
  assign u_CSAwallace_cska32_and_11_16 = a[11] & b[16];
  assign u_CSAwallace_cska32_and_12_16 = a[12] & b[16];
  assign u_CSAwallace_cska32_and_13_16 = a[13] & b[16];
  assign u_CSAwallace_cska32_and_14_16 = a[14] & b[16];
  assign u_CSAwallace_cska32_and_15_16 = a[15] & b[16];
  assign u_CSAwallace_cska32_and_16_16 = a[16] & b[16];
  assign u_CSAwallace_cska32_and_17_16 = a[17] & b[16];
  assign u_CSAwallace_cska32_and_18_16 = a[18] & b[16];
  assign u_CSAwallace_cska32_and_19_16 = a[19] & b[16];
  assign u_CSAwallace_cska32_and_20_16 = a[20] & b[16];
  assign u_CSAwallace_cska32_and_21_16 = a[21] & b[16];
  assign u_CSAwallace_cska32_and_22_16 = a[22] & b[16];
  assign u_CSAwallace_cska32_and_23_16 = a[23] & b[16];
  assign u_CSAwallace_cska32_and_24_16 = a[24] & b[16];
  assign u_CSAwallace_cska32_and_25_16 = a[25] & b[16];
  assign u_CSAwallace_cska32_and_26_16 = a[26] & b[16];
  assign u_CSAwallace_cska32_and_27_16 = a[27] & b[16];
  assign u_CSAwallace_cska32_and_28_16 = a[28] & b[16];
  assign u_CSAwallace_cska32_and_29_16 = a[29] & b[16];
  assign u_CSAwallace_cska32_and_30_16 = a[30] & b[16];
  assign u_CSAwallace_cska32_and_31_16 = a[31] & b[16];
  assign u_CSAwallace_cska32_and_0_17 = a[0] & b[17];
  assign u_CSAwallace_cska32_and_1_17 = a[1] & b[17];
  assign u_CSAwallace_cska32_and_2_17 = a[2] & b[17];
  assign u_CSAwallace_cska32_and_3_17 = a[3] & b[17];
  assign u_CSAwallace_cska32_and_4_17 = a[4] & b[17];
  assign u_CSAwallace_cska32_and_5_17 = a[5] & b[17];
  assign u_CSAwallace_cska32_and_6_17 = a[6] & b[17];
  assign u_CSAwallace_cska32_and_7_17 = a[7] & b[17];
  assign u_CSAwallace_cska32_and_8_17 = a[8] & b[17];
  assign u_CSAwallace_cska32_and_9_17 = a[9] & b[17];
  assign u_CSAwallace_cska32_and_10_17 = a[10] & b[17];
  assign u_CSAwallace_cska32_and_11_17 = a[11] & b[17];
  assign u_CSAwallace_cska32_and_12_17 = a[12] & b[17];
  assign u_CSAwallace_cska32_and_13_17 = a[13] & b[17];
  assign u_CSAwallace_cska32_and_14_17 = a[14] & b[17];
  assign u_CSAwallace_cska32_and_15_17 = a[15] & b[17];
  assign u_CSAwallace_cska32_and_16_17 = a[16] & b[17];
  assign u_CSAwallace_cska32_and_17_17 = a[17] & b[17];
  assign u_CSAwallace_cska32_and_18_17 = a[18] & b[17];
  assign u_CSAwallace_cska32_and_19_17 = a[19] & b[17];
  assign u_CSAwallace_cska32_and_20_17 = a[20] & b[17];
  assign u_CSAwallace_cska32_and_21_17 = a[21] & b[17];
  assign u_CSAwallace_cska32_and_22_17 = a[22] & b[17];
  assign u_CSAwallace_cska32_and_23_17 = a[23] & b[17];
  assign u_CSAwallace_cska32_and_24_17 = a[24] & b[17];
  assign u_CSAwallace_cska32_and_25_17 = a[25] & b[17];
  assign u_CSAwallace_cska32_and_26_17 = a[26] & b[17];
  assign u_CSAwallace_cska32_and_27_17 = a[27] & b[17];
  assign u_CSAwallace_cska32_and_28_17 = a[28] & b[17];
  assign u_CSAwallace_cska32_and_29_17 = a[29] & b[17];
  assign u_CSAwallace_cska32_and_30_17 = a[30] & b[17];
  assign u_CSAwallace_cska32_and_31_17 = a[31] & b[17];
  assign u_CSAwallace_cska32_and_0_18 = a[0] & b[18];
  assign u_CSAwallace_cska32_and_1_18 = a[1] & b[18];
  assign u_CSAwallace_cska32_and_2_18 = a[2] & b[18];
  assign u_CSAwallace_cska32_and_3_18 = a[3] & b[18];
  assign u_CSAwallace_cska32_and_4_18 = a[4] & b[18];
  assign u_CSAwallace_cska32_and_5_18 = a[5] & b[18];
  assign u_CSAwallace_cska32_and_6_18 = a[6] & b[18];
  assign u_CSAwallace_cska32_and_7_18 = a[7] & b[18];
  assign u_CSAwallace_cska32_and_8_18 = a[8] & b[18];
  assign u_CSAwallace_cska32_and_9_18 = a[9] & b[18];
  assign u_CSAwallace_cska32_and_10_18 = a[10] & b[18];
  assign u_CSAwallace_cska32_and_11_18 = a[11] & b[18];
  assign u_CSAwallace_cska32_and_12_18 = a[12] & b[18];
  assign u_CSAwallace_cska32_and_13_18 = a[13] & b[18];
  assign u_CSAwallace_cska32_and_14_18 = a[14] & b[18];
  assign u_CSAwallace_cska32_and_15_18 = a[15] & b[18];
  assign u_CSAwallace_cska32_and_16_18 = a[16] & b[18];
  assign u_CSAwallace_cska32_and_17_18 = a[17] & b[18];
  assign u_CSAwallace_cska32_and_18_18 = a[18] & b[18];
  assign u_CSAwallace_cska32_and_19_18 = a[19] & b[18];
  assign u_CSAwallace_cska32_and_20_18 = a[20] & b[18];
  assign u_CSAwallace_cska32_and_21_18 = a[21] & b[18];
  assign u_CSAwallace_cska32_and_22_18 = a[22] & b[18];
  assign u_CSAwallace_cska32_and_23_18 = a[23] & b[18];
  assign u_CSAwallace_cska32_and_24_18 = a[24] & b[18];
  assign u_CSAwallace_cska32_and_25_18 = a[25] & b[18];
  assign u_CSAwallace_cska32_and_26_18 = a[26] & b[18];
  assign u_CSAwallace_cska32_and_27_18 = a[27] & b[18];
  assign u_CSAwallace_cska32_and_28_18 = a[28] & b[18];
  assign u_CSAwallace_cska32_and_29_18 = a[29] & b[18];
  assign u_CSAwallace_cska32_and_30_18 = a[30] & b[18];
  assign u_CSAwallace_cska32_and_31_18 = a[31] & b[18];
  assign u_CSAwallace_cska32_and_0_19 = a[0] & b[19];
  assign u_CSAwallace_cska32_and_1_19 = a[1] & b[19];
  assign u_CSAwallace_cska32_and_2_19 = a[2] & b[19];
  assign u_CSAwallace_cska32_and_3_19 = a[3] & b[19];
  assign u_CSAwallace_cska32_and_4_19 = a[4] & b[19];
  assign u_CSAwallace_cska32_and_5_19 = a[5] & b[19];
  assign u_CSAwallace_cska32_and_6_19 = a[6] & b[19];
  assign u_CSAwallace_cska32_and_7_19 = a[7] & b[19];
  assign u_CSAwallace_cska32_and_8_19 = a[8] & b[19];
  assign u_CSAwallace_cska32_and_9_19 = a[9] & b[19];
  assign u_CSAwallace_cska32_and_10_19 = a[10] & b[19];
  assign u_CSAwallace_cska32_and_11_19 = a[11] & b[19];
  assign u_CSAwallace_cska32_and_12_19 = a[12] & b[19];
  assign u_CSAwallace_cska32_and_13_19 = a[13] & b[19];
  assign u_CSAwallace_cska32_and_14_19 = a[14] & b[19];
  assign u_CSAwallace_cska32_and_15_19 = a[15] & b[19];
  assign u_CSAwallace_cska32_and_16_19 = a[16] & b[19];
  assign u_CSAwallace_cska32_and_17_19 = a[17] & b[19];
  assign u_CSAwallace_cska32_and_18_19 = a[18] & b[19];
  assign u_CSAwallace_cska32_and_19_19 = a[19] & b[19];
  assign u_CSAwallace_cska32_and_20_19 = a[20] & b[19];
  assign u_CSAwallace_cska32_and_21_19 = a[21] & b[19];
  assign u_CSAwallace_cska32_and_22_19 = a[22] & b[19];
  assign u_CSAwallace_cska32_and_23_19 = a[23] & b[19];
  assign u_CSAwallace_cska32_and_24_19 = a[24] & b[19];
  assign u_CSAwallace_cska32_and_25_19 = a[25] & b[19];
  assign u_CSAwallace_cska32_and_26_19 = a[26] & b[19];
  assign u_CSAwallace_cska32_and_27_19 = a[27] & b[19];
  assign u_CSAwallace_cska32_and_28_19 = a[28] & b[19];
  assign u_CSAwallace_cska32_and_29_19 = a[29] & b[19];
  assign u_CSAwallace_cska32_and_30_19 = a[30] & b[19];
  assign u_CSAwallace_cska32_and_31_19 = a[31] & b[19];
  assign u_CSAwallace_cska32_and_0_20 = a[0] & b[20];
  assign u_CSAwallace_cska32_and_1_20 = a[1] & b[20];
  assign u_CSAwallace_cska32_and_2_20 = a[2] & b[20];
  assign u_CSAwallace_cska32_and_3_20 = a[3] & b[20];
  assign u_CSAwallace_cska32_and_4_20 = a[4] & b[20];
  assign u_CSAwallace_cska32_and_5_20 = a[5] & b[20];
  assign u_CSAwallace_cska32_and_6_20 = a[6] & b[20];
  assign u_CSAwallace_cska32_and_7_20 = a[7] & b[20];
  assign u_CSAwallace_cska32_and_8_20 = a[8] & b[20];
  assign u_CSAwallace_cska32_and_9_20 = a[9] & b[20];
  assign u_CSAwallace_cska32_and_10_20 = a[10] & b[20];
  assign u_CSAwallace_cska32_and_11_20 = a[11] & b[20];
  assign u_CSAwallace_cska32_and_12_20 = a[12] & b[20];
  assign u_CSAwallace_cska32_and_13_20 = a[13] & b[20];
  assign u_CSAwallace_cska32_and_14_20 = a[14] & b[20];
  assign u_CSAwallace_cska32_and_15_20 = a[15] & b[20];
  assign u_CSAwallace_cska32_and_16_20 = a[16] & b[20];
  assign u_CSAwallace_cska32_and_17_20 = a[17] & b[20];
  assign u_CSAwallace_cska32_and_18_20 = a[18] & b[20];
  assign u_CSAwallace_cska32_and_19_20 = a[19] & b[20];
  assign u_CSAwallace_cska32_and_20_20 = a[20] & b[20];
  assign u_CSAwallace_cska32_and_21_20 = a[21] & b[20];
  assign u_CSAwallace_cska32_and_22_20 = a[22] & b[20];
  assign u_CSAwallace_cska32_and_23_20 = a[23] & b[20];
  assign u_CSAwallace_cska32_and_24_20 = a[24] & b[20];
  assign u_CSAwallace_cska32_and_25_20 = a[25] & b[20];
  assign u_CSAwallace_cska32_and_26_20 = a[26] & b[20];
  assign u_CSAwallace_cska32_and_27_20 = a[27] & b[20];
  assign u_CSAwallace_cska32_and_28_20 = a[28] & b[20];
  assign u_CSAwallace_cska32_and_29_20 = a[29] & b[20];
  assign u_CSAwallace_cska32_and_30_20 = a[30] & b[20];
  assign u_CSAwallace_cska32_and_31_20 = a[31] & b[20];
  assign u_CSAwallace_cska32_and_0_21 = a[0] & b[21];
  assign u_CSAwallace_cska32_and_1_21 = a[1] & b[21];
  assign u_CSAwallace_cska32_and_2_21 = a[2] & b[21];
  assign u_CSAwallace_cska32_and_3_21 = a[3] & b[21];
  assign u_CSAwallace_cska32_and_4_21 = a[4] & b[21];
  assign u_CSAwallace_cska32_and_5_21 = a[5] & b[21];
  assign u_CSAwallace_cska32_and_6_21 = a[6] & b[21];
  assign u_CSAwallace_cska32_and_7_21 = a[7] & b[21];
  assign u_CSAwallace_cska32_and_8_21 = a[8] & b[21];
  assign u_CSAwallace_cska32_and_9_21 = a[9] & b[21];
  assign u_CSAwallace_cska32_and_10_21 = a[10] & b[21];
  assign u_CSAwallace_cska32_and_11_21 = a[11] & b[21];
  assign u_CSAwallace_cska32_and_12_21 = a[12] & b[21];
  assign u_CSAwallace_cska32_and_13_21 = a[13] & b[21];
  assign u_CSAwallace_cska32_and_14_21 = a[14] & b[21];
  assign u_CSAwallace_cska32_and_15_21 = a[15] & b[21];
  assign u_CSAwallace_cska32_and_16_21 = a[16] & b[21];
  assign u_CSAwallace_cska32_and_17_21 = a[17] & b[21];
  assign u_CSAwallace_cska32_and_18_21 = a[18] & b[21];
  assign u_CSAwallace_cska32_and_19_21 = a[19] & b[21];
  assign u_CSAwallace_cska32_and_20_21 = a[20] & b[21];
  assign u_CSAwallace_cska32_and_21_21 = a[21] & b[21];
  assign u_CSAwallace_cska32_and_22_21 = a[22] & b[21];
  assign u_CSAwallace_cska32_and_23_21 = a[23] & b[21];
  assign u_CSAwallace_cska32_and_24_21 = a[24] & b[21];
  assign u_CSAwallace_cska32_and_25_21 = a[25] & b[21];
  assign u_CSAwallace_cska32_and_26_21 = a[26] & b[21];
  assign u_CSAwallace_cska32_and_27_21 = a[27] & b[21];
  assign u_CSAwallace_cska32_and_28_21 = a[28] & b[21];
  assign u_CSAwallace_cska32_and_29_21 = a[29] & b[21];
  assign u_CSAwallace_cska32_and_30_21 = a[30] & b[21];
  assign u_CSAwallace_cska32_and_31_21 = a[31] & b[21];
  assign u_CSAwallace_cska32_and_0_22 = a[0] & b[22];
  assign u_CSAwallace_cska32_and_1_22 = a[1] & b[22];
  assign u_CSAwallace_cska32_and_2_22 = a[2] & b[22];
  assign u_CSAwallace_cska32_and_3_22 = a[3] & b[22];
  assign u_CSAwallace_cska32_and_4_22 = a[4] & b[22];
  assign u_CSAwallace_cska32_and_5_22 = a[5] & b[22];
  assign u_CSAwallace_cska32_and_6_22 = a[6] & b[22];
  assign u_CSAwallace_cska32_and_7_22 = a[7] & b[22];
  assign u_CSAwallace_cska32_and_8_22 = a[8] & b[22];
  assign u_CSAwallace_cska32_and_9_22 = a[9] & b[22];
  assign u_CSAwallace_cska32_and_10_22 = a[10] & b[22];
  assign u_CSAwallace_cska32_and_11_22 = a[11] & b[22];
  assign u_CSAwallace_cska32_and_12_22 = a[12] & b[22];
  assign u_CSAwallace_cska32_and_13_22 = a[13] & b[22];
  assign u_CSAwallace_cska32_and_14_22 = a[14] & b[22];
  assign u_CSAwallace_cska32_and_15_22 = a[15] & b[22];
  assign u_CSAwallace_cska32_and_16_22 = a[16] & b[22];
  assign u_CSAwallace_cska32_and_17_22 = a[17] & b[22];
  assign u_CSAwallace_cska32_and_18_22 = a[18] & b[22];
  assign u_CSAwallace_cska32_and_19_22 = a[19] & b[22];
  assign u_CSAwallace_cska32_and_20_22 = a[20] & b[22];
  assign u_CSAwallace_cska32_and_21_22 = a[21] & b[22];
  assign u_CSAwallace_cska32_and_22_22 = a[22] & b[22];
  assign u_CSAwallace_cska32_and_23_22 = a[23] & b[22];
  assign u_CSAwallace_cska32_and_24_22 = a[24] & b[22];
  assign u_CSAwallace_cska32_and_25_22 = a[25] & b[22];
  assign u_CSAwallace_cska32_and_26_22 = a[26] & b[22];
  assign u_CSAwallace_cska32_and_27_22 = a[27] & b[22];
  assign u_CSAwallace_cska32_and_28_22 = a[28] & b[22];
  assign u_CSAwallace_cska32_and_29_22 = a[29] & b[22];
  assign u_CSAwallace_cska32_and_30_22 = a[30] & b[22];
  assign u_CSAwallace_cska32_and_31_22 = a[31] & b[22];
  assign u_CSAwallace_cska32_and_0_23 = a[0] & b[23];
  assign u_CSAwallace_cska32_and_1_23 = a[1] & b[23];
  assign u_CSAwallace_cska32_and_2_23 = a[2] & b[23];
  assign u_CSAwallace_cska32_and_3_23 = a[3] & b[23];
  assign u_CSAwallace_cska32_and_4_23 = a[4] & b[23];
  assign u_CSAwallace_cska32_and_5_23 = a[5] & b[23];
  assign u_CSAwallace_cska32_and_6_23 = a[6] & b[23];
  assign u_CSAwallace_cska32_and_7_23 = a[7] & b[23];
  assign u_CSAwallace_cska32_and_8_23 = a[8] & b[23];
  assign u_CSAwallace_cska32_and_9_23 = a[9] & b[23];
  assign u_CSAwallace_cska32_and_10_23 = a[10] & b[23];
  assign u_CSAwallace_cska32_and_11_23 = a[11] & b[23];
  assign u_CSAwallace_cska32_and_12_23 = a[12] & b[23];
  assign u_CSAwallace_cska32_and_13_23 = a[13] & b[23];
  assign u_CSAwallace_cska32_and_14_23 = a[14] & b[23];
  assign u_CSAwallace_cska32_and_15_23 = a[15] & b[23];
  assign u_CSAwallace_cska32_and_16_23 = a[16] & b[23];
  assign u_CSAwallace_cska32_and_17_23 = a[17] & b[23];
  assign u_CSAwallace_cska32_and_18_23 = a[18] & b[23];
  assign u_CSAwallace_cska32_and_19_23 = a[19] & b[23];
  assign u_CSAwallace_cska32_and_20_23 = a[20] & b[23];
  assign u_CSAwallace_cska32_and_21_23 = a[21] & b[23];
  assign u_CSAwallace_cska32_and_22_23 = a[22] & b[23];
  assign u_CSAwallace_cska32_and_23_23 = a[23] & b[23];
  assign u_CSAwallace_cska32_and_24_23 = a[24] & b[23];
  assign u_CSAwallace_cska32_and_25_23 = a[25] & b[23];
  assign u_CSAwallace_cska32_and_26_23 = a[26] & b[23];
  assign u_CSAwallace_cska32_and_27_23 = a[27] & b[23];
  assign u_CSAwallace_cska32_and_28_23 = a[28] & b[23];
  assign u_CSAwallace_cska32_and_29_23 = a[29] & b[23];
  assign u_CSAwallace_cska32_and_30_23 = a[30] & b[23];
  assign u_CSAwallace_cska32_and_31_23 = a[31] & b[23];
  assign u_CSAwallace_cska32_and_0_24 = a[0] & b[24];
  assign u_CSAwallace_cska32_and_1_24 = a[1] & b[24];
  assign u_CSAwallace_cska32_and_2_24 = a[2] & b[24];
  assign u_CSAwallace_cska32_and_3_24 = a[3] & b[24];
  assign u_CSAwallace_cska32_and_4_24 = a[4] & b[24];
  assign u_CSAwallace_cska32_and_5_24 = a[5] & b[24];
  assign u_CSAwallace_cska32_and_6_24 = a[6] & b[24];
  assign u_CSAwallace_cska32_and_7_24 = a[7] & b[24];
  assign u_CSAwallace_cska32_and_8_24 = a[8] & b[24];
  assign u_CSAwallace_cska32_and_9_24 = a[9] & b[24];
  assign u_CSAwallace_cska32_and_10_24 = a[10] & b[24];
  assign u_CSAwallace_cska32_and_11_24 = a[11] & b[24];
  assign u_CSAwallace_cska32_and_12_24 = a[12] & b[24];
  assign u_CSAwallace_cska32_and_13_24 = a[13] & b[24];
  assign u_CSAwallace_cska32_and_14_24 = a[14] & b[24];
  assign u_CSAwallace_cska32_and_15_24 = a[15] & b[24];
  assign u_CSAwallace_cska32_and_16_24 = a[16] & b[24];
  assign u_CSAwallace_cska32_and_17_24 = a[17] & b[24];
  assign u_CSAwallace_cska32_and_18_24 = a[18] & b[24];
  assign u_CSAwallace_cska32_and_19_24 = a[19] & b[24];
  assign u_CSAwallace_cska32_and_20_24 = a[20] & b[24];
  assign u_CSAwallace_cska32_and_21_24 = a[21] & b[24];
  assign u_CSAwallace_cska32_and_22_24 = a[22] & b[24];
  assign u_CSAwallace_cska32_and_23_24 = a[23] & b[24];
  assign u_CSAwallace_cska32_and_24_24 = a[24] & b[24];
  assign u_CSAwallace_cska32_and_25_24 = a[25] & b[24];
  assign u_CSAwallace_cska32_and_26_24 = a[26] & b[24];
  assign u_CSAwallace_cska32_and_27_24 = a[27] & b[24];
  assign u_CSAwallace_cska32_and_28_24 = a[28] & b[24];
  assign u_CSAwallace_cska32_and_29_24 = a[29] & b[24];
  assign u_CSAwallace_cska32_and_30_24 = a[30] & b[24];
  assign u_CSAwallace_cska32_and_31_24 = a[31] & b[24];
  assign u_CSAwallace_cska32_and_0_25 = a[0] & b[25];
  assign u_CSAwallace_cska32_and_1_25 = a[1] & b[25];
  assign u_CSAwallace_cska32_and_2_25 = a[2] & b[25];
  assign u_CSAwallace_cska32_and_3_25 = a[3] & b[25];
  assign u_CSAwallace_cska32_and_4_25 = a[4] & b[25];
  assign u_CSAwallace_cska32_and_5_25 = a[5] & b[25];
  assign u_CSAwallace_cska32_and_6_25 = a[6] & b[25];
  assign u_CSAwallace_cska32_and_7_25 = a[7] & b[25];
  assign u_CSAwallace_cska32_and_8_25 = a[8] & b[25];
  assign u_CSAwallace_cska32_and_9_25 = a[9] & b[25];
  assign u_CSAwallace_cska32_and_10_25 = a[10] & b[25];
  assign u_CSAwallace_cska32_and_11_25 = a[11] & b[25];
  assign u_CSAwallace_cska32_and_12_25 = a[12] & b[25];
  assign u_CSAwallace_cska32_and_13_25 = a[13] & b[25];
  assign u_CSAwallace_cska32_and_14_25 = a[14] & b[25];
  assign u_CSAwallace_cska32_and_15_25 = a[15] & b[25];
  assign u_CSAwallace_cska32_and_16_25 = a[16] & b[25];
  assign u_CSAwallace_cska32_and_17_25 = a[17] & b[25];
  assign u_CSAwallace_cska32_and_18_25 = a[18] & b[25];
  assign u_CSAwallace_cska32_and_19_25 = a[19] & b[25];
  assign u_CSAwallace_cska32_and_20_25 = a[20] & b[25];
  assign u_CSAwallace_cska32_and_21_25 = a[21] & b[25];
  assign u_CSAwallace_cska32_and_22_25 = a[22] & b[25];
  assign u_CSAwallace_cska32_and_23_25 = a[23] & b[25];
  assign u_CSAwallace_cska32_and_24_25 = a[24] & b[25];
  assign u_CSAwallace_cska32_and_25_25 = a[25] & b[25];
  assign u_CSAwallace_cska32_and_26_25 = a[26] & b[25];
  assign u_CSAwallace_cska32_and_27_25 = a[27] & b[25];
  assign u_CSAwallace_cska32_and_28_25 = a[28] & b[25];
  assign u_CSAwallace_cska32_and_29_25 = a[29] & b[25];
  assign u_CSAwallace_cska32_and_30_25 = a[30] & b[25];
  assign u_CSAwallace_cska32_and_31_25 = a[31] & b[25];
  assign u_CSAwallace_cska32_and_0_26 = a[0] & b[26];
  assign u_CSAwallace_cska32_and_1_26 = a[1] & b[26];
  assign u_CSAwallace_cska32_and_2_26 = a[2] & b[26];
  assign u_CSAwallace_cska32_and_3_26 = a[3] & b[26];
  assign u_CSAwallace_cska32_and_4_26 = a[4] & b[26];
  assign u_CSAwallace_cska32_and_5_26 = a[5] & b[26];
  assign u_CSAwallace_cska32_and_6_26 = a[6] & b[26];
  assign u_CSAwallace_cska32_and_7_26 = a[7] & b[26];
  assign u_CSAwallace_cska32_and_8_26 = a[8] & b[26];
  assign u_CSAwallace_cska32_and_9_26 = a[9] & b[26];
  assign u_CSAwallace_cska32_and_10_26 = a[10] & b[26];
  assign u_CSAwallace_cska32_and_11_26 = a[11] & b[26];
  assign u_CSAwallace_cska32_and_12_26 = a[12] & b[26];
  assign u_CSAwallace_cska32_and_13_26 = a[13] & b[26];
  assign u_CSAwallace_cska32_and_14_26 = a[14] & b[26];
  assign u_CSAwallace_cska32_and_15_26 = a[15] & b[26];
  assign u_CSAwallace_cska32_and_16_26 = a[16] & b[26];
  assign u_CSAwallace_cska32_and_17_26 = a[17] & b[26];
  assign u_CSAwallace_cska32_and_18_26 = a[18] & b[26];
  assign u_CSAwallace_cska32_and_19_26 = a[19] & b[26];
  assign u_CSAwallace_cska32_and_20_26 = a[20] & b[26];
  assign u_CSAwallace_cska32_and_21_26 = a[21] & b[26];
  assign u_CSAwallace_cska32_and_22_26 = a[22] & b[26];
  assign u_CSAwallace_cska32_and_23_26 = a[23] & b[26];
  assign u_CSAwallace_cska32_and_24_26 = a[24] & b[26];
  assign u_CSAwallace_cska32_and_25_26 = a[25] & b[26];
  assign u_CSAwallace_cska32_and_26_26 = a[26] & b[26];
  assign u_CSAwallace_cska32_and_27_26 = a[27] & b[26];
  assign u_CSAwallace_cska32_and_28_26 = a[28] & b[26];
  assign u_CSAwallace_cska32_and_29_26 = a[29] & b[26];
  assign u_CSAwallace_cska32_and_30_26 = a[30] & b[26];
  assign u_CSAwallace_cska32_and_31_26 = a[31] & b[26];
  assign u_CSAwallace_cska32_and_0_27 = a[0] & b[27];
  assign u_CSAwallace_cska32_and_1_27 = a[1] & b[27];
  assign u_CSAwallace_cska32_and_2_27 = a[2] & b[27];
  assign u_CSAwallace_cska32_and_3_27 = a[3] & b[27];
  assign u_CSAwallace_cska32_and_4_27 = a[4] & b[27];
  assign u_CSAwallace_cska32_and_5_27 = a[5] & b[27];
  assign u_CSAwallace_cska32_and_6_27 = a[6] & b[27];
  assign u_CSAwallace_cska32_and_7_27 = a[7] & b[27];
  assign u_CSAwallace_cska32_and_8_27 = a[8] & b[27];
  assign u_CSAwallace_cska32_and_9_27 = a[9] & b[27];
  assign u_CSAwallace_cska32_and_10_27 = a[10] & b[27];
  assign u_CSAwallace_cska32_and_11_27 = a[11] & b[27];
  assign u_CSAwallace_cska32_and_12_27 = a[12] & b[27];
  assign u_CSAwallace_cska32_and_13_27 = a[13] & b[27];
  assign u_CSAwallace_cska32_and_14_27 = a[14] & b[27];
  assign u_CSAwallace_cska32_and_15_27 = a[15] & b[27];
  assign u_CSAwallace_cska32_and_16_27 = a[16] & b[27];
  assign u_CSAwallace_cska32_and_17_27 = a[17] & b[27];
  assign u_CSAwallace_cska32_and_18_27 = a[18] & b[27];
  assign u_CSAwallace_cska32_and_19_27 = a[19] & b[27];
  assign u_CSAwallace_cska32_and_20_27 = a[20] & b[27];
  assign u_CSAwallace_cska32_and_21_27 = a[21] & b[27];
  assign u_CSAwallace_cska32_and_22_27 = a[22] & b[27];
  assign u_CSAwallace_cska32_and_23_27 = a[23] & b[27];
  assign u_CSAwallace_cska32_and_24_27 = a[24] & b[27];
  assign u_CSAwallace_cska32_and_25_27 = a[25] & b[27];
  assign u_CSAwallace_cska32_and_26_27 = a[26] & b[27];
  assign u_CSAwallace_cska32_and_27_27 = a[27] & b[27];
  assign u_CSAwallace_cska32_and_28_27 = a[28] & b[27];
  assign u_CSAwallace_cska32_and_29_27 = a[29] & b[27];
  assign u_CSAwallace_cska32_and_30_27 = a[30] & b[27];
  assign u_CSAwallace_cska32_and_31_27 = a[31] & b[27];
  assign u_CSAwallace_cska32_and_0_28 = a[0] & b[28];
  assign u_CSAwallace_cska32_and_1_28 = a[1] & b[28];
  assign u_CSAwallace_cska32_and_2_28 = a[2] & b[28];
  assign u_CSAwallace_cska32_and_3_28 = a[3] & b[28];
  assign u_CSAwallace_cska32_and_4_28 = a[4] & b[28];
  assign u_CSAwallace_cska32_and_5_28 = a[5] & b[28];
  assign u_CSAwallace_cska32_and_6_28 = a[6] & b[28];
  assign u_CSAwallace_cska32_and_7_28 = a[7] & b[28];
  assign u_CSAwallace_cska32_and_8_28 = a[8] & b[28];
  assign u_CSAwallace_cska32_and_9_28 = a[9] & b[28];
  assign u_CSAwallace_cska32_and_10_28 = a[10] & b[28];
  assign u_CSAwallace_cska32_and_11_28 = a[11] & b[28];
  assign u_CSAwallace_cska32_and_12_28 = a[12] & b[28];
  assign u_CSAwallace_cska32_and_13_28 = a[13] & b[28];
  assign u_CSAwallace_cska32_and_14_28 = a[14] & b[28];
  assign u_CSAwallace_cska32_and_15_28 = a[15] & b[28];
  assign u_CSAwallace_cska32_and_16_28 = a[16] & b[28];
  assign u_CSAwallace_cska32_and_17_28 = a[17] & b[28];
  assign u_CSAwallace_cska32_and_18_28 = a[18] & b[28];
  assign u_CSAwallace_cska32_and_19_28 = a[19] & b[28];
  assign u_CSAwallace_cska32_and_20_28 = a[20] & b[28];
  assign u_CSAwallace_cska32_and_21_28 = a[21] & b[28];
  assign u_CSAwallace_cska32_and_22_28 = a[22] & b[28];
  assign u_CSAwallace_cska32_and_23_28 = a[23] & b[28];
  assign u_CSAwallace_cska32_and_24_28 = a[24] & b[28];
  assign u_CSAwallace_cska32_and_25_28 = a[25] & b[28];
  assign u_CSAwallace_cska32_and_26_28 = a[26] & b[28];
  assign u_CSAwallace_cska32_and_27_28 = a[27] & b[28];
  assign u_CSAwallace_cska32_and_28_28 = a[28] & b[28];
  assign u_CSAwallace_cska32_and_29_28 = a[29] & b[28];
  assign u_CSAwallace_cska32_and_30_28 = a[30] & b[28];
  assign u_CSAwallace_cska32_and_31_28 = a[31] & b[28];
  assign u_CSAwallace_cska32_and_0_29 = a[0] & b[29];
  assign u_CSAwallace_cska32_and_1_29 = a[1] & b[29];
  assign u_CSAwallace_cska32_and_2_29 = a[2] & b[29];
  assign u_CSAwallace_cska32_and_3_29 = a[3] & b[29];
  assign u_CSAwallace_cska32_and_4_29 = a[4] & b[29];
  assign u_CSAwallace_cska32_and_5_29 = a[5] & b[29];
  assign u_CSAwallace_cska32_and_6_29 = a[6] & b[29];
  assign u_CSAwallace_cska32_and_7_29 = a[7] & b[29];
  assign u_CSAwallace_cska32_and_8_29 = a[8] & b[29];
  assign u_CSAwallace_cska32_and_9_29 = a[9] & b[29];
  assign u_CSAwallace_cska32_and_10_29 = a[10] & b[29];
  assign u_CSAwallace_cska32_and_11_29 = a[11] & b[29];
  assign u_CSAwallace_cska32_and_12_29 = a[12] & b[29];
  assign u_CSAwallace_cska32_and_13_29 = a[13] & b[29];
  assign u_CSAwallace_cska32_and_14_29 = a[14] & b[29];
  assign u_CSAwallace_cska32_and_15_29 = a[15] & b[29];
  assign u_CSAwallace_cska32_and_16_29 = a[16] & b[29];
  assign u_CSAwallace_cska32_and_17_29 = a[17] & b[29];
  assign u_CSAwallace_cska32_and_18_29 = a[18] & b[29];
  assign u_CSAwallace_cska32_and_19_29 = a[19] & b[29];
  assign u_CSAwallace_cska32_and_20_29 = a[20] & b[29];
  assign u_CSAwallace_cska32_and_21_29 = a[21] & b[29];
  assign u_CSAwallace_cska32_and_22_29 = a[22] & b[29];
  assign u_CSAwallace_cska32_and_23_29 = a[23] & b[29];
  assign u_CSAwallace_cska32_and_24_29 = a[24] & b[29];
  assign u_CSAwallace_cska32_and_25_29 = a[25] & b[29];
  assign u_CSAwallace_cska32_and_26_29 = a[26] & b[29];
  assign u_CSAwallace_cska32_and_27_29 = a[27] & b[29];
  assign u_CSAwallace_cska32_and_28_29 = a[28] & b[29];
  assign u_CSAwallace_cska32_and_29_29 = a[29] & b[29];
  assign u_CSAwallace_cska32_and_30_29 = a[30] & b[29];
  assign u_CSAwallace_cska32_and_31_29 = a[31] & b[29];
  assign u_CSAwallace_cska32_and_0_30 = a[0] & b[30];
  assign u_CSAwallace_cska32_and_1_30 = a[1] & b[30];
  assign u_CSAwallace_cska32_and_2_30 = a[2] & b[30];
  assign u_CSAwallace_cska32_and_3_30 = a[3] & b[30];
  assign u_CSAwallace_cska32_and_4_30 = a[4] & b[30];
  assign u_CSAwallace_cska32_and_5_30 = a[5] & b[30];
  assign u_CSAwallace_cska32_and_6_30 = a[6] & b[30];
  assign u_CSAwallace_cska32_and_7_30 = a[7] & b[30];
  assign u_CSAwallace_cska32_and_8_30 = a[8] & b[30];
  assign u_CSAwallace_cska32_and_9_30 = a[9] & b[30];
  assign u_CSAwallace_cska32_and_10_30 = a[10] & b[30];
  assign u_CSAwallace_cska32_and_11_30 = a[11] & b[30];
  assign u_CSAwallace_cska32_and_12_30 = a[12] & b[30];
  assign u_CSAwallace_cska32_and_13_30 = a[13] & b[30];
  assign u_CSAwallace_cska32_and_14_30 = a[14] & b[30];
  assign u_CSAwallace_cska32_and_15_30 = a[15] & b[30];
  assign u_CSAwallace_cska32_and_16_30 = a[16] & b[30];
  assign u_CSAwallace_cska32_and_17_30 = a[17] & b[30];
  assign u_CSAwallace_cska32_and_18_30 = a[18] & b[30];
  assign u_CSAwallace_cska32_and_19_30 = a[19] & b[30];
  assign u_CSAwallace_cska32_and_20_30 = a[20] & b[30];
  assign u_CSAwallace_cska32_and_21_30 = a[21] & b[30];
  assign u_CSAwallace_cska32_and_22_30 = a[22] & b[30];
  assign u_CSAwallace_cska32_and_23_30 = a[23] & b[30];
  assign u_CSAwallace_cska32_and_24_30 = a[24] & b[30];
  assign u_CSAwallace_cska32_and_25_30 = a[25] & b[30];
  assign u_CSAwallace_cska32_and_26_30 = a[26] & b[30];
  assign u_CSAwallace_cska32_and_27_30 = a[27] & b[30];
  assign u_CSAwallace_cska32_and_28_30 = a[28] & b[30];
  assign u_CSAwallace_cska32_and_29_30 = a[29] & b[30];
  assign u_CSAwallace_cska32_and_30_30 = a[30] & b[30];
  assign u_CSAwallace_cska32_and_31_30 = a[31] & b[30];
  assign u_CSAwallace_cska32_and_0_31 = a[0] & b[31];
  assign u_CSAwallace_cska32_and_1_31 = a[1] & b[31];
  assign u_CSAwallace_cska32_and_2_31 = a[2] & b[31];
  assign u_CSAwallace_cska32_and_3_31 = a[3] & b[31];
  assign u_CSAwallace_cska32_and_4_31 = a[4] & b[31];
  assign u_CSAwallace_cska32_and_5_31 = a[5] & b[31];
  assign u_CSAwallace_cska32_and_6_31 = a[6] & b[31];
  assign u_CSAwallace_cska32_and_7_31 = a[7] & b[31];
  assign u_CSAwallace_cska32_and_8_31 = a[8] & b[31];
  assign u_CSAwallace_cska32_and_9_31 = a[9] & b[31];
  assign u_CSAwallace_cska32_and_10_31 = a[10] & b[31];
  assign u_CSAwallace_cska32_and_11_31 = a[11] & b[31];
  assign u_CSAwallace_cska32_and_12_31 = a[12] & b[31];
  assign u_CSAwallace_cska32_and_13_31 = a[13] & b[31];
  assign u_CSAwallace_cska32_and_14_31 = a[14] & b[31];
  assign u_CSAwallace_cska32_and_15_31 = a[15] & b[31];
  assign u_CSAwallace_cska32_and_16_31 = a[16] & b[31];
  assign u_CSAwallace_cska32_and_17_31 = a[17] & b[31];
  assign u_CSAwallace_cska32_and_18_31 = a[18] & b[31];
  assign u_CSAwallace_cska32_and_19_31 = a[19] & b[31];
  assign u_CSAwallace_cska32_and_20_31 = a[20] & b[31];
  assign u_CSAwallace_cska32_and_21_31 = a[21] & b[31];
  assign u_CSAwallace_cska32_and_22_31 = a[22] & b[31];
  assign u_CSAwallace_cska32_and_23_31 = a[23] & b[31];
  assign u_CSAwallace_cska32_and_24_31 = a[24] & b[31];
  assign u_CSAwallace_cska32_and_25_31 = a[25] & b[31];
  assign u_CSAwallace_cska32_and_26_31 = a[26] & b[31];
  assign u_CSAwallace_cska32_and_27_31 = a[27] & b[31];
  assign u_CSAwallace_cska32_and_28_31 = a[28] & b[31];
  assign u_CSAwallace_cska32_and_29_31 = a[29] & b[31];
  assign u_CSAwallace_cska32_and_30_31 = a[30] & b[31];
  assign u_CSAwallace_cska32_and_31_31 = a[31] & b[31];
  assign u_CSAwallace_cska32_csa0_csa_component_fa1_xor0 = u_CSAwallace_cska32_and_1_0 ^ u_CSAwallace_cska32_and_0_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa1_and0 = u_CSAwallace_cska32_and_1_0 & u_CSAwallace_cska32_and_0_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa2_xor0 = u_CSAwallace_cska32_and_2_0 ^ u_CSAwallace_cska32_and_1_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa2_and0 = u_CSAwallace_cska32_and_2_0 & u_CSAwallace_cska32_and_1_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa2_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa2_xor0 ^ u_CSAwallace_cska32_and_0_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa2_and1 = u_CSAwallace_cska32_csa0_csa_component_fa2_xor0 & u_CSAwallace_cska32_and_0_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa2_or0 = u_CSAwallace_cska32_csa0_csa_component_fa2_and0 | u_CSAwallace_cska32_csa0_csa_component_fa2_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa3_xor0 = u_CSAwallace_cska32_and_3_0 ^ u_CSAwallace_cska32_and_2_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa3_and0 = u_CSAwallace_cska32_and_3_0 & u_CSAwallace_cska32_and_2_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa3_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa3_xor0 ^ u_CSAwallace_cska32_and_1_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa3_and1 = u_CSAwallace_cska32_csa0_csa_component_fa3_xor0 & u_CSAwallace_cska32_and_1_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa3_or0 = u_CSAwallace_cska32_csa0_csa_component_fa3_and0 | u_CSAwallace_cska32_csa0_csa_component_fa3_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa4_xor0 = u_CSAwallace_cska32_and_4_0 ^ u_CSAwallace_cska32_and_3_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa4_and0 = u_CSAwallace_cska32_and_4_0 & u_CSAwallace_cska32_and_3_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa4_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa4_xor0 ^ u_CSAwallace_cska32_and_2_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa4_and1 = u_CSAwallace_cska32_csa0_csa_component_fa4_xor0 & u_CSAwallace_cska32_and_2_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa4_or0 = u_CSAwallace_cska32_csa0_csa_component_fa4_and0 | u_CSAwallace_cska32_csa0_csa_component_fa4_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa5_xor0 = u_CSAwallace_cska32_and_5_0 ^ u_CSAwallace_cska32_and_4_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa5_and0 = u_CSAwallace_cska32_and_5_0 & u_CSAwallace_cska32_and_4_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa5_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa5_xor0 ^ u_CSAwallace_cska32_and_3_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa5_and1 = u_CSAwallace_cska32_csa0_csa_component_fa5_xor0 & u_CSAwallace_cska32_and_3_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa5_or0 = u_CSAwallace_cska32_csa0_csa_component_fa5_and0 | u_CSAwallace_cska32_csa0_csa_component_fa5_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa6_xor0 = u_CSAwallace_cska32_and_6_0 ^ u_CSAwallace_cska32_and_5_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa6_and0 = u_CSAwallace_cska32_and_6_0 & u_CSAwallace_cska32_and_5_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa6_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa6_xor0 ^ u_CSAwallace_cska32_and_4_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa6_and1 = u_CSAwallace_cska32_csa0_csa_component_fa6_xor0 & u_CSAwallace_cska32_and_4_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa6_or0 = u_CSAwallace_cska32_csa0_csa_component_fa6_and0 | u_CSAwallace_cska32_csa0_csa_component_fa6_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa7_xor0 = u_CSAwallace_cska32_and_7_0 ^ u_CSAwallace_cska32_and_6_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa7_and0 = u_CSAwallace_cska32_and_7_0 & u_CSAwallace_cska32_and_6_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa7_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa7_xor0 ^ u_CSAwallace_cska32_and_5_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa7_and1 = u_CSAwallace_cska32_csa0_csa_component_fa7_xor0 & u_CSAwallace_cska32_and_5_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa7_or0 = u_CSAwallace_cska32_csa0_csa_component_fa7_and0 | u_CSAwallace_cska32_csa0_csa_component_fa7_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa8_xor0 = u_CSAwallace_cska32_and_8_0 ^ u_CSAwallace_cska32_and_7_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa8_and0 = u_CSAwallace_cska32_and_8_0 & u_CSAwallace_cska32_and_7_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa8_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_and_6_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa8_and1 = u_CSAwallace_cska32_csa0_csa_component_fa8_xor0 & u_CSAwallace_cska32_and_6_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa8_or0 = u_CSAwallace_cska32_csa0_csa_component_fa8_and0 | u_CSAwallace_cska32_csa0_csa_component_fa8_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa9_xor0 = u_CSAwallace_cska32_and_9_0 ^ u_CSAwallace_cska32_and_8_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa9_and0 = u_CSAwallace_cska32_and_9_0 & u_CSAwallace_cska32_and_8_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa9_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_and_7_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa9_and1 = u_CSAwallace_cska32_csa0_csa_component_fa9_xor0 & u_CSAwallace_cska32_and_7_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa9_or0 = u_CSAwallace_cska32_csa0_csa_component_fa9_and0 | u_CSAwallace_cska32_csa0_csa_component_fa9_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa10_xor0 = u_CSAwallace_cska32_and_10_0 ^ u_CSAwallace_cska32_and_9_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa10_and0 = u_CSAwallace_cska32_and_10_0 & u_CSAwallace_cska32_and_9_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa10_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_and_8_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa10_and1 = u_CSAwallace_cska32_csa0_csa_component_fa10_xor0 & u_CSAwallace_cska32_and_8_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa10_or0 = u_CSAwallace_cska32_csa0_csa_component_fa10_and0 | u_CSAwallace_cska32_csa0_csa_component_fa10_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa11_xor0 = u_CSAwallace_cska32_and_11_0 ^ u_CSAwallace_cska32_and_10_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa11_and0 = u_CSAwallace_cska32_and_11_0 & u_CSAwallace_cska32_and_10_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_and_9_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa11_and1 = u_CSAwallace_cska32_csa0_csa_component_fa11_xor0 & u_CSAwallace_cska32_and_9_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa11_or0 = u_CSAwallace_cska32_csa0_csa_component_fa11_and0 | u_CSAwallace_cska32_csa0_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa12_xor0 = u_CSAwallace_cska32_and_12_0 ^ u_CSAwallace_cska32_and_11_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa12_and0 = u_CSAwallace_cska32_and_12_0 & u_CSAwallace_cska32_and_11_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_and_10_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa12_and1 = u_CSAwallace_cska32_csa0_csa_component_fa12_xor0 & u_CSAwallace_cska32_and_10_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa12_or0 = u_CSAwallace_cska32_csa0_csa_component_fa12_and0 | u_CSAwallace_cska32_csa0_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa13_xor0 = u_CSAwallace_cska32_and_13_0 ^ u_CSAwallace_cska32_and_12_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa13_and0 = u_CSAwallace_cska32_and_13_0 & u_CSAwallace_cska32_and_12_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_and_11_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa13_and1 = u_CSAwallace_cska32_csa0_csa_component_fa13_xor0 & u_CSAwallace_cska32_and_11_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa13_or0 = u_CSAwallace_cska32_csa0_csa_component_fa13_and0 | u_CSAwallace_cska32_csa0_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa14_xor0 = u_CSAwallace_cska32_and_14_0 ^ u_CSAwallace_cska32_and_13_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa14_and0 = u_CSAwallace_cska32_and_14_0 & u_CSAwallace_cska32_and_13_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_and_12_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa14_and1 = u_CSAwallace_cska32_csa0_csa_component_fa14_xor0 & u_CSAwallace_cska32_and_12_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa14_or0 = u_CSAwallace_cska32_csa0_csa_component_fa14_and0 | u_CSAwallace_cska32_csa0_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa15_xor0 = u_CSAwallace_cska32_and_15_0 ^ u_CSAwallace_cska32_and_14_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa15_and0 = u_CSAwallace_cska32_and_15_0 & u_CSAwallace_cska32_and_14_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_and_13_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa15_and1 = u_CSAwallace_cska32_csa0_csa_component_fa15_xor0 & u_CSAwallace_cska32_and_13_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa15_or0 = u_CSAwallace_cska32_csa0_csa_component_fa15_and0 | u_CSAwallace_cska32_csa0_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa16_xor0 = u_CSAwallace_cska32_and_16_0 ^ u_CSAwallace_cska32_and_15_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa16_and0 = u_CSAwallace_cska32_and_16_0 & u_CSAwallace_cska32_and_15_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_and_14_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa16_and1 = u_CSAwallace_cska32_csa0_csa_component_fa16_xor0 & u_CSAwallace_cska32_and_14_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa16_or0 = u_CSAwallace_cska32_csa0_csa_component_fa16_and0 | u_CSAwallace_cska32_csa0_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa17_xor0 = u_CSAwallace_cska32_and_17_0 ^ u_CSAwallace_cska32_and_16_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa17_and0 = u_CSAwallace_cska32_and_17_0 & u_CSAwallace_cska32_and_16_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_and_15_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa17_and1 = u_CSAwallace_cska32_csa0_csa_component_fa17_xor0 & u_CSAwallace_cska32_and_15_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa17_or0 = u_CSAwallace_cska32_csa0_csa_component_fa17_and0 | u_CSAwallace_cska32_csa0_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa18_xor0 = u_CSAwallace_cska32_and_18_0 ^ u_CSAwallace_cska32_and_17_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa18_and0 = u_CSAwallace_cska32_and_18_0 & u_CSAwallace_cska32_and_17_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_and_16_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa18_and1 = u_CSAwallace_cska32_csa0_csa_component_fa18_xor0 & u_CSAwallace_cska32_and_16_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa18_or0 = u_CSAwallace_cska32_csa0_csa_component_fa18_and0 | u_CSAwallace_cska32_csa0_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa19_xor0 = u_CSAwallace_cska32_and_19_0 ^ u_CSAwallace_cska32_and_18_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa19_and0 = u_CSAwallace_cska32_and_19_0 & u_CSAwallace_cska32_and_18_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_and_17_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa19_and1 = u_CSAwallace_cska32_csa0_csa_component_fa19_xor0 & u_CSAwallace_cska32_and_17_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa19_or0 = u_CSAwallace_cska32_csa0_csa_component_fa19_and0 | u_CSAwallace_cska32_csa0_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa20_xor0 = u_CSAwallace_cska32_and_20_0 ^ u_CSAwallace_cska32_and_19_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa20_and0 = u_CSAwallace_cska32_and_20_0 & u_CSAwallace_cska32_and_19_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_and_18_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa20_and1 = u_CSAwallace_cska32_csa0_csa_component_fa20_xor0 & u_CSAwallace_cska32_and_18_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa20_or0 = u_CSAwallace_cska32_csa0_csa_component_fa20_and0 | u_CSAwallace_cska32_csa0_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa21_xor0 = u_CSAwallace_cska32_and_21_0 ^ u_CSAwallace_cska32_and_20_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa21_and0 = u_CSAwallace_cska32_and_21_0 & u_CSAwallace_cska32_and_20_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_and_19_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa21_and1 = u_CSAwallace_cska32_csa0_csa_component_fa21_xor0 & u_CSAwallace_cska32_and_19_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa21_or0 = u_CSAwallace_cska32_csa0_csa_component_fa21_and0 | u_CSAwallace_cska32_csa0_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa22_xor0 = u_CSAwallace_cska32_and_22_0 ^ u_CSAwallace_cska32_and_21_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa22_and0 = u_CSAwallace_cska32_and_22_0 & u_CSAwallace_cska32_and_21_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_and_20_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa22_and1 = u_CSAwallace_cska32_csa0_csa_component_fa22_xor0 & u_CSAwallace_cska32_and_20_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa22_or0 = u_CSAwallace_cska32_csa0_csa_component_fa22_and0 | u_CSAwallace_cska32_csa0_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa23_xor0 = u_CSAwallace_cska32_and_23_0 ^ u_CSAwallace_cska32_and_22_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa23_and0 = u_CSAwallace_cska32_and_23_0 & u_CSAwallace_cska32_and_22_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_and_21_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa23_and1 = u_CSAwallace_cska32_csa0_csa_component_fa23_xor0 & u_CSAwallace_cska32_and_21_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa23_or0 = u_CSAwallace_cska32_csa0_csa_component_fa23_and0 | u_CSAwallace_cska32_csa0_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa24_xor0 = u_CSAwallace_cska32_and_24_0 ^ u_CSAwallace_cska32_and_23_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa24_and0 = u_CSAwallace_cska32_and_24_0 & u_CSAwallace_cska32_and_23_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_and_22_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa24_and1 = u_CSAwallace_cska32_csa0_csa_component_fa24_xor0 & u_CSAwallace_cska32_and_22_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa24_or0 = u_CSAwallace_cska32_csa0_csa_component_fa24_and0 | u_CSAwallace_cska32_csa0_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_25_0 ^ u_CSAwallace_cska32_and_24_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa25_and0 = u_CSAwallace_cska32_and_25_0 & u_CSAwallace_cska32_and_24_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_and_23_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa25_and1 = u_CSAwallace_cska32_csa0_csa_component_fa25_xor0 & u_CSAwallace_cska32_and_23_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa25_or0 = u_CSAwallace_cska32_csa0_csa_component_fa25_and0 | u_CSAwallace_cska32_csa0_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_26_0 ^ u_CSAwallace_cska32_and_25_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa26_and0 = u_CSAwallace_cska32_and_26_0 & u_CSAwallace_cska32_and_25_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_24_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa26_and1 = u_CSAwallace_cska32_csa0_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_24_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa26_or0 = u_CSAwallace_cska32_csa0_csa_component_fa26_and0 | u_CSAwallace_cska32_csa0_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_27_0 ^ u_CSAwallace_cska32_and_26_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa27_and0 = u_CSAwallace_cska32_and_27_0 & u_CSAwallace_cska32_and_26_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_25_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa27_and1 = u_CSAwallace_cska32_csa0_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_25_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa27_or0 = u_CSAwallace_cska32_csa0_csa_component_fa27_and0 | u_CSAwallace_cska32_csa0_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_28_0 ^ u_CSAwallace_cska32_and_27_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa28_and0 = u_CSAwallace_cska32_and_28_0 & u_CSAwallace_cska32_and_27_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_26_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa28_and1 = u_CSAwallace_cska32_csa0_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_26_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa28_or0 = u_CSAwallace_cska32_csa0_csa_component_fa28_and0 | u_CSAwallace_cska32_csa0_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_29_0 ^ u_CSAwallace_cska32_and_28_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa29_and0 = u_CSAwallace_cska32_and_29_0 & u_CSAwallace_cska32_and_28_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_27_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa29_and1 = u_CSAwallace_cska32_csa0_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_27_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa29_or0 = u_CSAwallace_cska32_csa0_csa_component_fa29_and0 | u_CSAwallace_cska32_csa0_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_30_0 ^ u_CSAwallace_cska32_and_29_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa30_and0 = u_CSAwallace_cska32_and_30_0 & u_CSAwallace_cska32_and_29_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_28_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa30_and1 = u_CSAwallace_cska32_csa0_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_28_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa30_or0 = u_CSAwallace_cska32_csa0_csa_component_fa30_and0 | u_CSAwallace_cska32_csa0_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_31_0 ^ u_CSAwallace_cska32_and_30_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa31_and0 = u_CSAwallace_cska32_and_31_0 & u_CSAwallace_cska32_and_30_1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa0_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_29_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa31_and1 = u_CSAwallace_cska32_csa0_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_29_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa31_or0 = u_CSAwallace_cska32_csa0_csa_component_fa31_and0 | u_CSAwallace_cska32_csa0_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa0_csa_component_fa32_xor1 = u_CSAwallace_cska32_and_31_1 ^ u_CSAwallace_cska32_and_30_2;
  assign u_CSAwallace_cska32_csa0_csa_component_fa32_and1 = u_CSAwallace_cska32_and_31_1 & u_CSAwallace_cska32_and_30_2;
  assign u_CSAwallace_cska32_csa1_csa_component_fa4_xor0 = u_CSAwallace_cska32_and_1_3 ^ u_CSAwallace_cska32_and_0_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa4_and0 = u_CSAwallace_cska32_and_1_3 & u_CSAwallace_cska32_and_0_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa5_xor0 = u_CSAwallace_cska32_and_2_3 ^ u_CSAwallace_cska32_and_1_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa5_and0 = u_CSAwallace_cska32_and_2_3 & u_CSAwallace_cska32_and_1_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa5_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa5_xor0 ^ u_CSAwallace_cska32_and_0_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa5_and1 = u_CSAwallace_cska32_csa1_csa_component_fa5_xor0 & u_CSAwallace_cska32_and_0_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa5_or0 = u_CSAwallace_cska32_csa1_csa_component_fa5_and0 | u_CSAwallace_cska32_csa1_csa_component_fa5_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa6_xor0 = u_CSAwallace_cska32_and_3_3 ^ u_CSAwallace_cska32_and_2_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa6_and0 = u_CSAwallace_cska32_and_3_3 & u_CSAwallace_cska32_and_2_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa6_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa6_xor0 ^ u_CSAwallace_cska32_and_1_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa6_and1 = u_CSAwallace_cska32_csa1_csa_component_fa6_xor0 & u_CSAwallace_cska32_and_1_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa6_or0 = u_CSAwallace_cska32_csa1_csa_component_fa6_and0 | u_CSAwallace_cska32_csa1_csa_component_fa6_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa7_xor0 = u_CSAwallace_cska32_and_4_3 ^ u_CSAwallace_cska32_and_3_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa7_and0 = u_CSAwallace_cska32_and_4_3 & u_CSAwallace_cska32_and_3_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa7_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa7_xor0 ^ u_CSAwallace_cska32_and_2_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa7_and1 = u_CSAwallace_cska32_csa1_csa_component_fa7_xor0 & u_CSAwallace_cska32_and_2_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa7_or0 = u_CSAwallace_cska32_csa1_csa_component_fa7_and0 | u_CSAwallace_cska32_csa1_csa_component_fa7_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa8_xor0 = u_CSAwallace_cska32_and_5_3 ^ u_CSAwallace_cska32_and_4_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa8_and0 = u_CSAwallace_cska32_and_5_3 & u_CSAwallace_cska32_and_4_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa8_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_and_3_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa8_and1 = u_CSAwallace_cska32_csa1_csa_component_fa8_xor0 & u_CSAwallace_cska32_and_3_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa8_or0 = u_CSAwallace_cska32_csa1_csa_component_fa8_and0 | u_CSAwallace_cska32_csa1_csa_component_fa8_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa9_xor0 = u_CSAwallace_cska32_and_6_3 ^ u_CSAwallace_cska32_and_5_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa9_and0 = u_CSAwallace_cska32_and_6_3 & u_CSAwallace_cska32_and_5_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa9_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_and_4_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa9_and1 = u_CSAwallace_cska32_csa1_csa_component_fa9_xor0 & u_CSAwallace_cska32_and_4_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa9_or0 = u_CSAwallace_cska32_csa1_csa_component_fa9_and0 | u_CSAwallace_cska32_csa1_csa_component_fa9_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa10_xor0 = u_CSAwallace_cska32_and_7_3 ^ u_CSAwallace_cska32_and_6_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa10_and0 = u_CSAwallace_cska32_and_7_3 & u_CSAwallace_cska32_and_6_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa10_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_and_5_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa10_and1 = u_CSAwallace_cska32_csa1_csa_component_fa10_xor0 & u_CSAwallace_cska32_and_5_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa10_or0 = u_CSAwallace_cska32_csa1_csa_component_fa10_and0 | u_CSAwallace_cska32_csa1_csa_component_fa10_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa11_xor0 = u_CSAwallace_cska32_and_8_3 ^ u_CSAwallace_cska32_and_7_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa11_and0 = u_CSAwallace_cska32_and_8_3 & u_CSAwallace_cska32_and_7_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_and_6_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa11_and1 = u_CSAwallace_cska32_csa1_csa_component_fa11_xor0 & u_CSAwallace_cska32_and_6_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa11_or0 = u_CSAwallace_cska32_csa1_csa_component_fa11_and0 | u_CSAwallace_cska32_csa1_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa12_xor0 = u_CSAwallace_cska32_and_9_3 ^ u_CSAwallace_cska32_and_8_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa12_and0 = u_CSAwallace_cska32_and_9_3 & u_CSAwallace_cska32_and_8_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_and_7_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa12_and1 = u_CSAwallace_cska32_csa1_csa_component_fa12_xor0 & u_CSAwallace_cska32_and_7_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa12_or0 = u_CSAwallace_cska32_csa1_csa_component_fa12_and0 | u_CSAwallace_cska32_csa1_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa13_xor0 = u_CSAwallace_cska32_and_10_3 ^ u_CSAwallace_cska32_and_9_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa13_and0 = u_CSAwallace_cska32_and_10_3 & u_CSAwallace_cska32_and_9_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_and_8_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa13_and1 = u_CSAwallace_cska32_csa1_csa_component_fa13_xor0 & u_CSAwallace_cska32_and_8_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa13_or0 = u_CSAwallace_cska32_csa1_csa_component_fa13_and0 | u_CSAwallace_cska32_csa1_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa14_xor0 = u_CSAwallace_cska32_and_11_3 ^ u_CSAwallace_cska32_and_10_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa14_and0 = u_CSAwallace_cska32_and_11_3 & u_CSAwallace_cska32_and_10_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_and_9_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa14_and1 = u_CSAwallace_cska32_csa1_csa_component_fa14_xor0 & u_CSAwallace_cska32_and_9_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa14_or0 = u_CSAwallace_cska32_csa1_csa_component_fa14_and0 | u_CSAwallace_cska32_csa1_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa15_xor0 = u_CSAwallace_cska32_and_12_3 ^ u_CSAwallace_cska32_and_11_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa15_and0 = u_CSAwallace_cska32_and_12_3 & u_CSAwallace_cska32_and_11_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_and_10_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa15_and1 = u_CSAwallace_cska32_csa1_csa_component_fa15_xor0 & u_CSAwallace_cska32_and_10_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa15_or0 = u_CSAwallace_cska32_csa1_csa_component_fa15_and0 | u_CSAwallace_cska32_csa1_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa16_xor0 = u_CSAwallace_cska32_and_13_3 ^ u_CSAwallace_cska32_and_12_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa16_and0 = u_CSAwallace_cska32_and_13_3 & u_CSAwallace_cska32_and_12_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_and_11_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa16_and1 = u_CSAwallace_cska32_csa1_csa_component_fa16_xor0 & u_CSAwallace_cska32_and_11_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa16_or0 = u_CSAwallace_cska32_csa1_csa_component_fa16_and0 | u_CSAwallace_cska32_csa1_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa17_xor0 = u_CSAwallace_cska32_and_14_3 ^ u_CSAwallace_cska32_and_13_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa17_and0 = u_CSAwallace_cska32_and_14_3 & u_CSAwallace_cska32_and_13_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_and_12_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa17_and1 = u_CSAwallace_cska32_csa1_csa_component_fa17_xor0 & u_CSAwallace_cska32_and_12_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa17_or0 = u_CSAwallace_cska32_csa1_csa_component_fa17_and0 | u_CSAwallace_cska32_csa1_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa18_xor0 = u_CSAwallace_cska32_and_15_3 ^ u_CSAwallace_cska32_and_14_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa18_and0 = u_CSAwallace_cska32_and_15_3 & u_CSAwallace_cska32_and_14_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_and_13_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa18_and1 = u_CSAwallace_cska32_csa1_csa_component_fa18_xor0 & u_CSAwallace_cska32_and_13_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa18_or0 = u_CSAwallace_cska32_csa1_csa_component_fa18_and0 | u_CSAwallace_cska32_csa1_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa19_xor0 = u_CSAwallace_cska32_and_16_3 ^ u_CSAwallace_cska32_and_15_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa19_and0 = u_CSAwallace_cska32_and_16_3 & u_CSAwallace_cska32_and_15_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_and_14_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa19_and1 = u_CSAwallace_cska32_csa1_csa_component_fa19_xor0 & u_CSAwallace_cska32_and_14_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa19_or0 = u_CSAwallace_cska32_csa1_csa_component_fa19_and0 | u_CSAwallace_cska32_csa1_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa20_xor0 = u_CSAwallace_cska32_and_17_3 ^ u_CSAwallace_cska32_and_16_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa20_and0 = u_CSAwallace_cska32_and_17_3 & u_CSAwallace_cska32_and_16_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_and_15_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa20_and1 = u_CSAwallace_cska32_csa1_csa_component_fa20_xor0 & u_CSAwallace_cska32_and_15_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa20_or0 = u_CSAwallace_cska32_csa1_csa_component_fa20_and0 | u_CSAwallace_cska32_csa1_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa21_xor0 = u_CSAwallace_cska32_and_18_3 ^ u_CSAwallace_cska32_and_17_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa21_and0 = u_CSAwallace_cska32_and_18_3 & u_CSAwallace_cska32_and_17_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_and_16_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa21_and1 = u_CSAwallace_cska32_csa1_csa_component_fa21_xor0 & u_CSAwallace_cska32_and_16_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa21_or0 = u_CSAwallace_cska32_csa1_csa_component_fa21_and0 | u_CSAwallace_cska32_csa1_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa22_xor0 = u_CSAwallace_cska32_and_19_3 ^ u_CSAwallace_cska32_and_18_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa22_and0 = u_CSAwallace_cska32_and_19_3 & u_CSAwallace_cska32_and_18_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_and_17_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa22_and1 = u_CSAwallace_cska32_csa1_csa_component_fa22_xor0 & u_CSAwallace_cska32_and_17_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa22_or0 = u_CSAwallace_cska32_csa1_csa_component_fa22_and0 | u_CSAwallace_cska32_csa1_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa23_xor0 = u_CSAwallace_cska32_and_20_3 ^ u_CSAwallace_cska32_and_19_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa23_and0 = u_CSAwallace_cska32_and_20_3 & u_CSAwallace_cska32_and_19_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_and_18_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa23_and1 = u_CSAwallace_cska32_csa1_csa_component_fa23_xor0 & u_CSAwallace_cska32_and_18_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa23_or0 = u_CSAwallace_cska32_csa1_csa_component_fa23_and0 | u_CSAwallace_cska32_csa1_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa24_xor0 = u_CSAwallace_cska32_and_21_3 ^ u_CSAwallace_cska32_and_20_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa24_and0 = u_CSAwallace_cska32_and_21_3 & u_CSAwallace_cska32_and_20_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_and_19_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa24_and1 = u_CSAwallace_cska32_csa1_csa_component_fa24_xor0 & u_CSAwallace_cska32_and_19_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa24_or0 = u_CSAwallace_cska32_csa1_csa_component_fa24_and0 | u_CSAwallace_cska32_csa1_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_22_3 ^ u_CSAwallace_cska32_and_21_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa25_and0 = u_CSAwallace_cska32_and_22_3 & u_CSAwallace_cska32_and_21_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_and_20_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa25_and1 = u_CSAwallace_cska32_csa1_csa_component_fa25_xor0 & u_CSAwallace_cska32_and_20_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa25_or0 = u_CSAwallace_cska32_csa1_csa_component_fa25_and0 | u_CSAwallace_cska32_csa1_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_23_3 ^ u_CSAwallace_cska32_and_22_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa26_and0 = u_CSAwallace_cska32_and_23_3 & u_CSAwallace_cska32_and_22_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_21_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa26_and1 = u_CSAwallace_cska32_csa1_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_21_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa26_or0 = u_CSAwallace_cska32_csa1_csa_component_fa26_and0 | u_CSAwallace_cska32_csa1_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_24_3 ^ u_CSAwallace_cska32_and_23_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa27_and0 = u_CSAwallace_cska32_and_24_3 & u_CSAwallace_cska32_and_23_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_22_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa27_and1 = u_CSAwallace_cska32_csa1_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_22_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa27_or0 = u_CSAwallace_cska32_csa1_csa_component_fa27_and0 | u_CSAwallace_cska32_csa1_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_25_3 ^ u_CSAwallace_cska32_and_24_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa28_and0 = u_CSAwallace_cska32_and_25_3 & u_CSAwallace_cska32_and_24_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_23_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa28_and1 = u_CSAwallace_cska32_csa1_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_23_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa28_or0 = u_CSAwallace_cska32_csa1_csa_component_fa28_and0 | u_CSAwallace_cska32_csa1_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_26_3 ^ u_CSAwallace_cska32_and_25_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa29_and0 = u_CSAwallace_cska32_and_26_3 & u_CSAwallace_cska32_and_25_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_24_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa29_and1 = u_CSAwallace_cska32_csa1_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_24_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa29_or0 = u_CSAwallace_cska32_csa1_csa_component_fa29_and0 | u_CSAwallace_cska32_csa1_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_27_3 ^ u_CSAwallace_cska32_and_26_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa30_and0 = u_CSAwallace_cska32_and_27_3 & u_CSAwallace_cska32_and_26_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_25_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa30_and1 = u_CSAwallace_cska32_csa1_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_25_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa30_or0 = u_CSAwallace_cska32_csa1_csa_component_fa30_and0 | u_CSAwallace_cska32_csa1_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_28_3 ^ u_CSAwallace_cska32_and_27_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa31_and0 = u_CSAwallace_cska32_and_28_3 & u_CSAwallace_cska32_and_27_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_26_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa31_and1 = u_CSAwallace_cska32_csa1_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_26_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa31_or0 = u_CSAwallace_cska32_csa1_csa_component_fa31_and0 | u_CSAwallace_cska32_csa1_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_29_3 ^ u_CSAwallace_cska32_and_28_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa32_and0 = u_CSAwallace_cska32_and_29_3 & u_CSAwallace_cska32_and_28_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_27_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa32_and1 = u_CSAwallace_cska32_csa1_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_27_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa32_or0 = u_CSAwallace_cska32_csa1_csa_component_fa32_and0 | u_CSAwallace_cska32_csa1_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_30_3 ^ u_CSAwallace_cska32_and_29_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa33_and0 = u_CSAwallace_cska32_and_30_3 & u_CSAwallace_cska32_and_29_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_28_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa33_and1 = u_CSAwallace_cska32_csa1_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_28_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa33_or0 = u_CSAwallace_cska32_csa1_csa_component_fa33_and0 | u_CSAwallace_cska32_csa1_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_31_3 ^ u_CSAwallace_cska32_and_30_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa34_and0 = u_CSAwallace_cska32_and_31_3 & u_CSAwallace_cska32_and_30_4;
  assign u_CSAwallace_cska32_csa1_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_29_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa34_and1 = u_CSAwallace_cska32_csa1_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_29_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa34_or0 = u_CSAwallace_cska32_csa1_csa_component_fa34_and0 | u_CSAwallace_cska32_csa1_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa1_csa_component_fa35_xor1 = u_CSAwallace_cska32_and_31_4 ^ u_CSAwallace_cska32_and_30_5;
  assign u_CSAwallace_cska32_csa1_csa_component_fa35_and1 = u_CSAwallace_cska32_and_31_4 & u_CSAwallace_cska32_and_30_5;
  assign u_CSAwallace_cska32_csa2_csa_component_fa7_xor0 = u_CSAwallace_cska32_and_1_6 ^ u_CSAwallace_cska32_and_0_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa7_and0 = u_CSAwallace_cska32_and_1_6 & u_CSAwallace_cska32_and_0_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa8_xor0 = u_CSAwallace_cska32_and_2_6 ^ u_CSAwallace_cska32_and_1_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa8_and0 = u_CSAwallace_cska32_and_2_6 & u_CSAwallace_cska32_and_1_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa8_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_and_0_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa8_and1 = u_CSAwallace_cska32_csa2_csa_component_fa8_xor0 & u_CSAwallace_cska32_and_0_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa8_or0 = u_CSAwallace_cska32_csa2_csa_component_fa8_and0 | u_CSAwallace_cska32_csa2_csa_component_fa8_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa9_xor0 = u_CSAwallace_cska32_and_3_6 ^ u_CSAwallace_cska32_and_2_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa9_and0 = u_CSAwallace_cska32_and_3_6 & u_CSAwallace_cska32_and_2_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa9_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_and_1_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa9_and1 = u_CSAwallace_cska32_csa2_csa_component_fa9_xor0 & u_CSAwallace_cska32_and_1_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa9_or0 = u_CSAwallace_cska32_csa2_csa_component_fa9_and0 | u_CSAwallace_cska32_csa2_csa_component_fa9_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa10_xor0 = u_CSAwallace_cska32_and_4_6 ^ u_CSAwallace_cska32_and_3_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa10_and0 = u_CSAwallace_cska32_and_4_6 & u_CSAwallace_cska32_and_3_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa10_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_and_2_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa10_and1 = u_CSAwallace_cska32_csa2_csa_component_fa10_xor0 & u_CSAwallace_cska32_and_2_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa10_or0 = u_CSAwallace_cska32_csa2_csa_component_fa10_and0 | u_CSAwallace_cska32_csa2_csa_component_fa10_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa11_xor0 = u_CSAwallace_cska32_and_5_6 ^ u_CSAwallace_cska32_and_4_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa11_and0 = u_CSAwallace_cska32_and_5_6 & u_CSAwallace_cska32_and_4_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_and_3_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa11_and1 = u_CSAwallace_cska32_csa2_csa_component_fa11_xor0 & u_CSAwallace_cska32_and_3_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa11_or0 = u_CSAwallace_cska32_csa2_csa_component_fa11_and0 | u_CSAwallace_cska32_csa2_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa12_xor0 = u_CSAwallace_cska32_and_6_6 ^ u_CSAwallace_cska32_and_5_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa12_and0 = u_CSAwallace_cska32_and_6_6 & u_CSAwallace_cska32_and_5_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_and_4_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa12_and1 = u_CSAwallace_cska32_csa2_csa_component_fa12_xor0 & u_CSAwallace_cska32_and_4_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa12_or0 = u_CSAwallace_cska32_csa2_csa_component_fa12_and0 | u_CSAwallace_cska32_csa2_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa13_xor0 = u_CSAwallace_cska32_and_7_6 ^ u_CSAwallace_cska32_and_6_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa13_and0 = u_CSAwallace_cska32_and_7_6 & u_CSAwallace_cska32_and_6_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_and_5_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa13_and1 = u_CSAwallace_cska32_csa2_csa_component_fa13_xor0 & u_CSAwallace_cska32_and_5_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa13_or0 = u_CSAwallace_cska32_csa2_csa_component_fa13_and0 | u_CSAwallace_cska32_csa2_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa14_xor0 = u_CSAwallace_cska32_and_8_6 ^ u_CSAwallace_cska32_and_7_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa14_and0 = u_CSAwallace_cska32_and_8_6 & u_CSAwallace_cska32_and_7_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_and_6_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa14_and1 = u_CSAwallace_cska32_csa2_csa_component_fa14_xor0 & u_CSAwallace_cska32_and_6_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa14_or0 = u_CSAwallace_cska32_csa2_csa_component_fa14_and0 | u_CSAwallace_cska32_csa2_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa15_xor0 = u_CSAwallace_cska32_and_9_6 ^ u_CSAwallace_cska32_and_8_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa15_and0 = u_CSAwallace_cska32_and_9_6 & u_CSAwallace_cska32_and_8_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_and_7_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa15_and1 = u_CSAwallace_cska32_csa2_csa_component_fa15_xor0 & u_CSAwallace_cska32_and_7_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa15_or0 = u_CSAwallace_cska32_csa2_csa_component_fa15_and0 | u_CSAwallace_cska32_csa2_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa16_xor0 = u_CSAwallace_cska32_and_10_6 ^ u_CSAwallace_cska32_and_9_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa16_and0 = u_CSAwallace_cska32_and_10_6 & u_CSAwallace_cska32_and_9_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_and_8_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa16_and1 = u_CSAwallace_cska32_csa2_csa_component_fa16_xor0 & u_CSAwallace_cska32_and_8_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa16_or0 = u_CSAwallace_cska32_csa2_csa_component_fa16_and0 | u_CSAwallace_cska32_csa2_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa17_xor0 = u_CSAwallace_cska32_and_11_6 ^ u_CSAwallace_cska32_and_10_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa17_and0 = u_CSAwallace_cska32_and_11_6 & u_CSAwallace_cska32_and_10_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_and_9_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa17_and1 = u_CSAwallace_cska32_csa2_csa_component_fa17_xor0 & u_CSAwallace_cska32_and_9_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa17_or0 = u_CSAwallace_cska32_csa2_csa_component_fa17_and0 | u_CSAwallace_cska32_csa2_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa18_xor0 = u_CSAwallace_cska32_and_12_6 ^ u_CSAwallace_cska32_and_11_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa18_and0 = u_CSAwallace_cska32_and_12_6 & u_CSAwallace_cska32_and_11_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_and_10_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa18_and1 = u_CSAwallace_cska32_csa2_csa_component_fa18_xor0 & u_CSAwallace_cska32_and_10_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa18_or0 = u_CSAwallace_cska32_csa2_csa_component_fa18_and0 | u_CSAwallace_cska32_csa2_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa19_xor0 = u_CSAwallace_cska32_and_13_6 ^ u_CSAwallace_cska32_and_12_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa19_and0 = u_CSAwallace_cska32_and_13_6 & u_CSAwallace_cska32_and_12_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_and_11_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa19_and1 = u_CSAwallace_cska32_csa2_csa_component_fa19_xor0 & u_CSAwallace_cska32_and_11_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa19_or0 = u_CSAwallace_cska32_csa2_csa_component_fa19_and0 | u_CSAwallace_cska32_csa2_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa20_xor0 = u_CSAwallace_cska32_and_14_6 ^ u_CSAwallace_cska32_and_13_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa20_and0 = u_CSAwallace_cska32_and_14_6 & u_CSAwallace_cska32_and_13_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_and_12_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa20_and1 = u_CSAwallace_cska32_csa2_csa_component_fa20_xor0 & u_CSAwallace_cska32_and_12_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa20_or0 = u_CSAwallace_cska32_csa2_csa_component_fa20_and0 | u_CSAwallace_cska32_csa2_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa21_xor0 = u_CSAwallace_cska32_and_15_6 ^ u_CSAwallace_cska32_and_14_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa21_and0 = u_CSAwallace_cska32_and_15_6 & u_CSAwallace_cska32_and_14_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_and_13_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa21_and1 = u_CSAwallace_cska32_csa2_csa_component_fa21_xor0 & u_CSAwallace_cska32_and_13_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa21_or0 = u_CSAwallace_cska32_csa2_csa_component_fa21_and0 | u_CSAwallace_cska32_csa2_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa22_xor0 = u_CSAwallace_cska32_and_16_6 ^ u_CSAwallace_cska32_and_15_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa22_and0 = u_CSAwallace_cska32_and_16_6 & u_CSAwallace_cska32_and_15_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_and_14_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa22_and1 = u_CSAwallace_cska32_csa2_csa_component_fa22_xor0 & u_CSAwallace_cska32_and_14_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa22_or0 = u_CSAwallace_cska32_csa2_csa_component_fa22_and0 | u_CSAwallace_cska32_csa2_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa23_xor0 = u_CSAwallace_cska32_and_17_6 ^ u_CSAwallace_cska32_and_16_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa23_and0 = u_CSAwallace_cska32_and_17_6 & u_CSAwallace_cska32_and_16_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_and_15_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa23_and1 = u_CSAwallace_cska32_csa2_csa_component_fa23_xor0 & u_CSAwallace_cska32_and_15_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa23_or0 = u_CSAwallace_cska32_csa2_csa_component_fa23_and0 | u_CSAwallace_cska32_csa2_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa24_xor0 = u_CSAwallace_cska32_and_18_6 ^ u_CSAwallace_cska32_and_17_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa24_and0 = u_CSAwallace_cska32_and_18_6 & u_CSAwallace_cska32_and_17_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_and_16_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa24_and1 = u_CSAwallace_cska32_csa2_csa_component_fa24_xor0 & u_CSAwallace_cska32_and_16_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa24_or0 = u_CSAwallace_cska32_csa2_csa_component_fa24_and0 | u_CSAwallace_cska32_csa2_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_19_6 ^ u_CSAwallace_cska32_and_18_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa25_and0 = u_CSAwallace_cska32_and_19_6 & u_CSAwallace_cska32_and_18_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_and_17_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa25_and1 = u_CSAwallace_cska32_csa2_csa_component_fa25_xor0 & u_CSAwallace_cska32_and_17_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa25_or0 = u_CSAwallace_cska32_csa2_csa_component_fa25_and0 | u_CSAwallace_cska32_csa2_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_20_6 ^ u_CSAwallace_cska32_and_19_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa26_and0 = u_CSAwallace_cska32_and_20_6 & u_CSAwallace_cska32_and_19_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_18_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa26_and1 = u_CSAwallace_cska32_csa2_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_18_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa26_or0 = u_CSAwallace_cska32_csa2_csa_component_fa26_and0 | u_CSAwallace_cska32_csa2_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_21_6 ^ u_CSAwallace_cska32_and_20_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa27_and0 = u_CSAwallace_cska32_and_21_6 & u_CSAwallace_cska32_and_20_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_19_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa27_and1 = u_CSAwallace_cska32_csa2_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_19_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa27_or0 = u_CSAwallace_cska32_csa2_csa_component_fa27_and0 | u_CSAwallace_cska32_csa2_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_22_6 ^ u_CSAwallace_cska32_and_21_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa28_and0 = u_CSAwallace_cska32_and_22_6 & u_CSAwallace_cska32_and_21_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_20_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa28_and1 = u_CSAwallace_cska32_csa2_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_20_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa28_or0 = u_CSAwallace_cska32_csa2_csa_component_fa28_and0 | u_CSAwallace_cska32_csa2_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_23_6 ^ u_CSAwallace_cska32_and_22_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa29_and0 = u_CSAwallace_cska32_and_23_6 & u_CSAwallace_cska32_and_22_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_21_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa29_and1 = u_CSAwallace_cska32_csa2_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_21_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa29_or0 = u_CSAwallace_cska32_csa2_csa_component_fa29_and0 | u_CSAwallace_cska32_csa2_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_24_6 ^ u_CSAwallace_cska32_and_23_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa30_and0 = u_CSAwallace_cska32_and_24_6 & u_CSAwallace_cska32_and_23_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_22_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa30_and1 = u_CSAwallace_cska32_csa2_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_22_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa30_or0 = u_CSAwallace_cska32_csa2_csa_component_fa30_and0 | u_CSAwallace_cska32_csa2_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_25_6 ^ u_CSAwallace_cska32_and_24_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa31_and0 = u_CSAwallace_cska32_and_25_6 & u_CSAwallace_cska32_and_24_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_23_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa31_and1 = u_CSAwallace_cska32_csa2_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_23_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa31_or0 = u_CSAwallace_cska32_csa2_csa_component_fa31_and0 | u_CSAwallace_cska32_csa2_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_26_6 ^ u_CSAwallace_cska32_and_25_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa32_and0 = u_CSAwallace_cska32_and_26_6 & u_CSAwallace_cska32_and_25_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_24_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa32_and1 = u_CSAwallace_cska32_csa2_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_24_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa32_or0 = u_CSAwallace_cska32_csa2_csa_component_fa32_and0 | u_CSAwallace_cska32_csa2_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_27_6 ^ u_CSAwallace_cska32_and_26_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa33_and0 = u_CSAwallace_cska32_and_27_6 & u_CSAwallace_cska32_and_26_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_25_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa33_and1 = u_CSAwallace_cska32_csa2_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_25_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa33_or0 = u_CSAwallace_cska32_csa2_csa_component_fa33_and0 | u_CSAwallace_cska32_csa2_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_28_6 ^ u_CSAwallace_cska32_and_27_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa34_and0 = u_CSAwallace_cska32_and_28_6 & u_CSAwallace_cska32_and_27_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_26_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa34_and1 = u_CSAwallace_cska32_csa2_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_26_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa34_or0 = u_CSAwallace_cska32_csa2_csa_component_fa34_and0 | u_CSAwallace_cska32_csa2_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa35_xor0 = u_CSAwallace_cska32_and_29_6 ^ u_CSAwallace_cska32_and_28_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa35_and0 = u_CSAwallace_cska32_and_29_6 & u_CSAwallace_cska32_and_28_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_27_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa35_and1 = u_CSAwallace_cska32_csa2_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_27_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa35_or0 = u_CSAwallace_cska32_csa2_csa_component_fa35_and0 | u_CSAwallace_cska32_csa2_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa36_xor0 = u_CSAwallace_cska32_and_30_6 ^ u_CSAwallace_cska32_and_29_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa36_and0 = u_CSAwallace_cska32_and_30_6 & u_CSAwallace_cska32_and_29_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_28_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa36_and1 = u_CSAwallace_cska32_csa2_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_28_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa36_or0 = u_CSAwallace_cska32_csa2_csa_component_fa36_and0 | u_CSAwallace_cska32_csa2_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa37_xor0 = u_CSAwallace_cska32_and_31_6 ^ u_CSAwallace_cska32_and_30_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa37_and0 = u_CSAwallace_cska32_and_31_6 & u_CSAwallace_cska32_and_30_7;
  assign u_CSAwallace_cska32_csa2_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_29_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa37_and1 = u_CSAwallace_cska32_csa2_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_29_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa37_or0 = u_CSAwallace_cska32_csa2_csa_component_fa37_and0 | u_CSAwallace_cska32_csa2_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa2_csa_component_fa38_xor1 = u_CSAwallace_cska32_and_31_7 ^ u_CSAwallace_cska32_and_30_8;
  assign u_CSAwallace_cska32_csa2_csa_component_fa38_and1 = u_CSAwallace_cska32_and_31_7 & u_CSAwallace_cska32_and_30_8;
  assign u_CSAwallace_cska32_csa3_csa_component_fa10_xor0 = u_CSAwallace_cska32_and_1_9 ^ u_CSAwallace_cska32_and_0_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa10_and0 = u_CSAwallace_cska32_and_1_9 & u_CSAwallace_cska32_and_0_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa11_xor0 = u_CSAwallace_cska32_and_2_9 ^ u_CSAwallace_cska32_and_1_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa11_and0 = u_CSAwallace_cska32_and_2_9 & u_CSAwallace_cska32_and_1_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_and_0_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa11_and1 = u_CSAwallace_cska32_csa3_csa_component_fa11_xor0 & u_CSAwallace_cska32_and_0_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa11_or0 = u_CSAwallace_cska32_csa3_csa_component_fa11_and0 | u_CSAwallace_cska32_csa3_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa12_xor0 = u_CSAwallace_cska32_and_3_9 ^ u_CSAwallace_cska32_and_2_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa12_and0 = u_CSAwallace_cska32_and_3_9 & u_CSAwallace_cska32_and_2_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_and_1_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa12_and1 = u_CSAwallace_cska32_csa3_csa_component_fa12_xor0 & u_CSAwallace_cska32_and_1_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa12_or0 = u_CSAwallace_cska32_csa3_csa_component_fa12_and0 | u_CSAwallace_cska32_csa3_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa13_xor0 = u_CSAwallace_cska32_and_4_9 ^ u_CSAwallace_cska32_and_3_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa13_and0 = u_CSAwallace_cska32_and_4_9 & u_CSAwallace_cska32_and_3_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_and_2_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa13_and1 = u_CSAwallace_cska32_csa3_csa_component_fa13_xor0 & u_CSAwallace_cska32_and_2_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa13_or0 = u_CSAwallace_cska32_csa3_csa_component_fa13_and0 | u_CSAwallace_cska32_csa3_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa14_xor0 = u_CSAwallace_cska32_and_5_9 ^ u_CSAwallace_cska32_and_4_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa14_and0 = u_CSAwallace_cska32_and_5_9 & u_CSAwallace_cska32_and_4_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_and_3_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa14_and1 = u_CSAwallace_cska32_csa3_csa_component_fa14_xor0 & u_CSAwallace_cska32_and_3_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa14_or0 = u_CSAwallace_cska32_csa3_csa_component_fa14_and0 | u_CSAwallace_cska32_csa3_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa15_xor0 = u_CSAwallace_cska32_and_6_9 ^ u_CSAwallace_cska32_and_5_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa15_and0 = u_CSAwallace_cska32_and_6_9 & u_CSAwallace_cska32_and_5_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_and_4_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa15_and1 = u_CSAwallace_cska32_csa3_csa_component_fa15_xor0 & u_CSAwallace_cska32_and_4_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa15_or0 = u_CSAwallace_cska32_csa3_csa_component_fa15_and0 | u_CSAwallace_cska32_csa3_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa16_xor0 = u_CSAwallace_cska32_and_7_9 ^ u_CSAwallace_cska32_and_6_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa16_and0 = u_CSAwallace_cska32_and_7_9 & u_CSAwallace_cska32_and_6_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_and_5_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa16_and1 = u_CSAwallace_cska32_csa3_csa_component_fa16_xor0 & u_CSAwallace_cska32_and_5_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa16_or0 = u_CSAwallace_cska32_csa3_csa_component_fa16_and0 | u_CSAwallace_cska32_csa3_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa17_xor0 = u_CSAwallace_cska32_and_8_9 ^ u_CSAwallace_cska32_and_7_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa17_and0 = u_CSAwallace_cska32_and_8_9 & u_CSAwallace_cska32_and_7_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_and_6_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa17_and1 = u_CSAwallace_cska32_csa3_csa_component_fa17_xor0 & u_CSAwallace_cska32_and_6_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa17_or0 = u_CSAwallace_cska32_csa3_csa_component_fa17_and0 | u_CSAwallace_cska32_csa3_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa18_xor0 = u_CSAwallace_cska32_and_9_9 ^ u_CSAwallace_cska32_and_8_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa18_and0 = u_CSAwallace_cska32_and_9_9 & u_CSAwallace_cska32_and_8_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_and_7_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa18_and1 = u_CSAwallace_cska32_csa3_csa_component_fa18_xor0 & u_CSAwallace_cska32_and_7_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa18_or0 = u_CSAwallace_cska32_csa3_csa_component_fa18_and0 | u_CSAwallace_cska32_csa3_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa19_xor0 = u_CSAwallace_cska32_and_10_9 ^ u_CSAwallace_cska32_and_9_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa19_and0 = u_CSAwallace_cska32_and_10_9 & u_CSAwallace_cska32_and_9_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_and_8_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa19_and1 = u_CSAwallace_cska32_csa3_csa_component_fa19_xor0 & u_CSAwallace_cska32_and_8_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa19_or0 = u_CSAwallace_cska32_csa3_csa_component_fa19_and0 | u_CSAwallace_cska32_csa3_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa20_xor0 = u_CSAwallace_cska32_and_11_9 ^ u_CSAwallace_cska32_and_10_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa20_and0 = u_CSAwallace_cska32_and_11_9 & u_CSAwallace_cska32_and_10_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_and_9_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa20_and1 = u_CSAwallace_cska32_csa3_csa_component_fa20_xor0 & u_CSAwallace_cska32_and_9_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa20_or0 = u_CSAwallace_cska32_csa3_csa_component_fa20_and0 | u_CSAwallace_cska32_csa3_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa21_xor0 = u_CSAwallace_cska32_and_12_9 ^ u_CSAwallace_cska32_and_11_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa21_and0 = u_CSAwallace_cska32_and_12_9 & u_CSAwallace_cska32_and_11_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_and_10_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa21_and1 = u_CSAwallace_cska32_csa3_csa_component_fa21_xor0 & u_CSAwallace_cska32_and_10_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa21_or0 = u_CSAwallace_cska32_csa3_csa_component_fa21_and0 | u_CSAwallace_cska32_csa3_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa22_xor0 = u_CSAwallace_cska32_and_13_9 ^ u_CSAwallace_cska32_and_12_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa22_and0 = u_CSAwallace_cska32_and_13_9 & u_CSAwallace_cska32_and_12_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_and_11_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa22_and1 = u_CSAwallace_cska32_csa3_csa_component_fa22_xor0 & u_CSAwallace_cska32_and_11_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa22_or0 = u_CSAwallace_cska32_csa3_csa_component_fa22_and0 | u_CSAwallace_cska32_csa3_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa23_xor0 = u_CSAwallace_cska32_and_14_9 ^ u_CSAwallace_cska32_and_13_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa23_and0 = u_CSAwallace_cska32_and_14_9 & u_CSAwallace_cska32_and_13_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_and_12_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa23_and1 = u_CSAwallace_cska32_csa3_csa_component_fa23_xor0 & u_CSAwallace_cska32_and_12_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa23_or0 = u_CSAwallace_cska32_csa3_csa_component_fa23_and0 | u_CSAwallace_cska32_csa3_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa24_xor0 = u_CSAwallace_cska32_and_15_9 ^ u_CSAwallace_cska32_and_14_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa24_and0 = u_CSAwallace_cska32_and_15_9 & u_CSAwallace_cska32_and_14_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_and_13_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa24_and1 = u_CSAwallace_cska32_csa3_csa_component_fa24_xor0 & u_CSAwallace_cska32_and_13_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa24_or0 = u_CSAwallace_cska32_csa3_csa_component_fa24_and0 | u_CSAwallace_cska32_csa3_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_16_9 ^ u_CSAwallace_cska32_and_15_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa25_and0 = u_CSAwallace_cska32_and_16_9 & u_CSAwallace_cska32_and_15_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_and_14_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa25_and1 = u_CSAwallace_cska32_csa3_csa_component_fa25_xor0 & u_CSAwallace_cska32_and_14_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa25_or0 = u_CSAwallace_cska32_csa3_csa_component_fa25_and0 | u_CSAwallace_cska32_csa3_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_17_9 ^ u_CSAwallace_cska32_and_16_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa26_and0 = u_CSAwallace_cska32_and_17_9 & u_CSAwallace_cska32_and_16_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_15_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa26_and1 = u_CSAwallace_cska32_csa3_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_15_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa26_or0 = u_CSAwallace_cska32_csa3_csa_component_fa26_and0 | u_CSAwallace_cska32_csa3_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_18_9 ^ u_CSAwallace_cska32_and_17_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa27_and0 = u_CSAwallace_cska32_and_18_9 & u_CSAwallace_cska32_and_17_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_16_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa27_and1 = u_CSAwallace_cska32_csa3_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_16_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa27_or0 = u_CSAwallace_cska32_csa3_csa_component_fa27_and0 | u_CSAwallace_cska32_csa3_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_19_9 ^ u_CSAwallace_cska32_and_18_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa28_and0 = u_CSAwallace_cska32_and_19_9 & u_CSAwallace_cska32_and_18_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_17_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa28_and1 = u_CSAwallace_cska32_csa3_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_17_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa28_or0 = u_CSAwallace_cska32_csa3_csa_component_fa28_and0 | u_CSAwallace_cska32_csa3_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_20_9 ^ u_CSAwallace_cska32_and_19_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa29_and0 = u_CSAwallace_cska32_and_20_9 & u_CSAwallace_cska32_and_19_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_18_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa29_and1 = u_CSAwallace_cska32_csa3_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_18_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa29_or0 = u_CSAwallace_cska32_csa3_csa_component_fa29_and0 | u_CSAwallace_cska32_csa3_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_21_9 ^ u_CSAwallace_cska32_and_20_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa30_and0 = u_CSAwallace_cska32_and_21_9 & u_CSAwallace_cska32_and_20_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_19_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa30_and1 = u_CSAwallace_cska32_csa3_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_19_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa30_or0 = u_CSAwallace_cska32_csa3_csa_component_fa30_and0 | u_CSAwallace_cska32_csa3_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_22_9 ^ u_CSAwallace_cska32_and_21_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa31_and0 = u_CSAwallace_cska32_and_22_9 & u_CSAwallace_cska32_and_21_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_20_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa31_and1 = u_CSAwallace_cska32_csa3_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_20_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa31_or0 = u_CSAwallace_cska32_csa3_csa_component_fa31_and0 | u_CSAwallace_cska32_csa3_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_23_9 ^ u_CSAwallace_cska32_and_22_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa32_and0 = u_CSAwallace_cska32_and_23_9 & u_CSAwallace_cska32_and_22_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_21_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa32_and1 = u_CSAwallace_cska32_csa3_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_21_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa32_or0 = u_CSAwallace_cska32_csa3_csa_component_fa32_and0 | u_CSAwallace_cska32_csa3_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_24_9 ^ u_CSAwallace_cska32_and_23_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa33_and0 = u_CSAwallace_cska32_and_24_9 & u_CSAwallace_cska32_and_23_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_22_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa33_and1 = u_CSAwallace_cska32_csa3_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_22_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa33_or0 = u_CSAwallace_cska32_csa3_csa_component_fa33_and0 | u_CSAwallace_cska32_csa3_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_25_9 ^ u_CSAwallace_cska32_and_24_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa34_and0 = u_CSAwallace_cska32_and_25_9 & u_CSAwallace_cska32_and_24_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_23_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa34_and1 = u_CSAwallace_cska32_csa3_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_23_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa34_or0 = u_CSAwallace_cska32_csa3_csa_component_fa34_and0 | u_CSAwallace_cska32_csa3_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa35_xor0 = u_CSAwallace_cska32_and_26_9 ^ u_CSAwallace_cska32_and_25_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa35_and0 = u_CSAwallace_cska32_and_26_9 & u_CSAwallace_cska32_and_25_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_24_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa35_and1 = u_CSAwallace_cska32_csa3_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_24_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa35_or0 = u_CSAwallace_cska32_csa3_csa_component_fa35_and0 | u_CSAwallace_cska32_csa3_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa36_xor0 = u_CSAwallace_cska32_and_27_9 ^ u_CSAwallace_cska32_and_26_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa36_and0 = u_CSAwallace_cska32_and_27_9 & u_CSAwallace_cska32_and_26_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_25_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa36_and1 = u_CSAwallace_cska32_csa3_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_25_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa36_or0 = u_CSAwallace_cska32_csa3_csa_component_fa36_and0 | u_CSAwallace_cska32_csa3_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa37_xor0 = u_CSAwallace_cska32_and_28_9 ^ u_CSAwallace_cska32_and_27_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa37_and0 = u_CSAwallace_cska32_and_28_9 & u_CSAwallace_cska32_and_27_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_26_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa37_and1 = u_CSAwallace_cska32_csa3_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_26_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa37_or0 = u_CSAwallace_cska32_csa3_csa_component_fa37_and0 | u_CSAwallace_cska32_csa3_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa38_xor0 = u_CSAwallace_cska32_and_29_9 ^ u_CSAwallace_cska32_and_28_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa38_and0 = u_CSAwallace_cska32_and_29_9 & u_CSAwallace_cska32_and_28_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_27_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa38_and1 = u_CSAwallace_cska32_csa3_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_27_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa38_or0 = u_CSAwallace_cska32_csa3_csa_component_fa38_and0 | u_CSAwallace_cska32_csa3_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa39_xor0 = u_CSAwallace_cska32_and_30_9 ^ u_CSAwallace_cska32_and_29_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa39_and0 = u_CSAwallace_cska32_and_30_9 & u_CSAwallace_cska32_and_29_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_28_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa39_and1 = u_CSAwallace_cska32_csa3_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_28_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa39_or0 = u_CSAwallace_cska32_csa3_csa_component_fa39_and0 | u_CSAwallace_cska32_csa3_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa40_xor0 = u_CSAwallace_cska32_and_31_9 ^ u_CSAwallace_cska32_and_30_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa40_and0 = u_CSAwallace_cska32_and_31_9 & u_CSAwallace_cska32_and_30_10;
  assign u_CSAwallace_cska32_csa3_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa3_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_29_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa40_and1 = u_CSAwallace_cska32_csa3_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_29_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa40_or0 = u_CSAwallace_cska32_csa3_csa_component_fa40_and0 | u_CSAwallace_cska32_csa3_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa3_csa_component_fa41_xor1 = u_CSAwallace_cska32_and_31_10 ^ u_CSAwallace_cska32_and_30_11;
  assign u_CSAwallace_cska32_csa3_csa_component_fa41_and1 = u_CSAwallace_cska32_and_31_10 & u_CSAwallace_cska32_and_30_11;
  assign u_CSAwallace_cska32_csa4_csa_component_fa13_xor0 = u_CSAwallace_cska32_and_1_12 ^ u_CSAwallace_cska32_and_0_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa13_and0 = u_CSAwallace_cska32_and_1_12 & u_CSAwallace_cska32_and_0_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa14_xor0 = u_CSAwallace_cska32_and_2_12 ^ u_CSAwallace_cska32_and_1_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa14_and0 = u_CSAwallace_cska32_and_2_12 & u_CSAwallace_cska32_and_1_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_and_0_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa14_and1 = u_CSAwallace_cska32_csa4_csa_component_fa14_xor0 & u_CSAwallace_cska32_and_0_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa14_or0 = u_CSAwallace_cska32_csa4_csa_component_fa14_and0 | u_CSAwallace_cska32_csa4_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa15_xor0 = u_CSAwallace_cska32_and_3_12 ^ u_CSAwallace_cska32_and_2_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa15_and0 = u_CSAwallace_cska32_and_3_12 & u_CSAwallace_cska32_and_2_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_and_1_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa15_and1 = u_CSAwallace_cska32_csa4_csa_component_fa15_xor0 & u_CSAwallace_cska32_and_1_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa15_or0 = u_CSAwallace_cska32_csa4_csa_component_fa15_and0 | u_CSAwallace_cska32_csa4_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa16_xor0 = u_CSAwallace_cska32_and_4_12 ^ u_CSAwallace_cska32_and_3_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa16_and0 = u_CSAwallace_cska32_and_4_12 & u_CSAwallace_cska32_and_3_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_and_2_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa16_and1 = u_CSAwallace_cska32_csa4_csa_component_fa16_xor0 & u_CSAwallace_cska32_and_2_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa16_or0 = u_CSAwallace_cska32_csa4_csa_component_fa16_and0 | u_CSAwallace_cska32_csa4_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa17_xor0 = u_CSAwallace_cska32_and_5_12 ^ u_CSAwallace_cska32_and_4_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa17_and0 = u_CSAwallace_cska32_and_5_12 & u_CSAwallace_cska32_and_4_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_and_3_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa17_and1 = u_CSAwallace_cska32_csa4_csa_component_fa17_xor0 & u_CSAwallace_cska32_and_3_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa17_or0 = u_CSAwallace_cska32_csa4_csa_component_fa17_and0 | u_CSAwallace_cska32_csa4_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa18_xor0 = u_CSAwallace_cska32_and_6_12 ^ u_CSAwallace_cska32_and_5_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa18_and0 = u_CSAwallace_cska32_and_6_12 & u_CSAwallace_cska32_and_5_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_and_4_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa18_and1 = u_CSAwallace_cska32_csa4_csa_component_fa18_xor0 & u_CSAwallace_cska32_and_4_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa18_or0 = u_CSAwallace_cska32_csa4_csa_component_fa18_and0 | u_CSAwallace_cska32_csa4_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa19_xor0 = u_CSAwallace_cska32_and_7_12 ^ u_CSAwallace_cska32_and_6_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa19_and0 = u_CSAwallace_cska32_and_7_12 & u_CSAwallace_cska32_and_6_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_and_5_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa19_and1 = u_CSAwallace_cska32_csa4_csa_component_fa19_xor0 & u_CSAwallace_cska32_and_5_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa19_or0 = u_CSAwallace_cska32_csa4_csa_component_fa19_and0 | u_CSAwallace_cska32_csa4_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa20_xor0 = u_CSAwallace_cska32_and_8_12 ^ u_CSAwallace_cska32_and_7_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa20_and0 = u_CSAwallace_cska32_and_8_12 & u_CSAwallace_cska32_and_7_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_and_6_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa20_and1 = u_CSAwallace_cska32_csa4_csa_component_fa20_xor0 & u_CSAwallace_cska32_and_6_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa20_or0 = u_CSAwallace_cska32_csa4_csa_component_fa20_and0 | u_CSAwallace_cska32_csa4_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa21_xor0 = u_CSAwallace_cska32_and_9_12 ^ u_CSAwallace_cska32_and_8_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa21_and0 = u_CSAwallace_cska32_and_9_12 & u_CSAwallace_cska32_and_8_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_and_7_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa21_and1 = u_CSAwallace_cska32_csa4_csa_component_fa21_xor0 & u_CSAwallace_cska32_and_7_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa21_or0 = u_CSAwallace_cska32_csa4_csa_component_fa21_and0 | u_CSAwallace_cska32_csa4_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa22_xor0 = u_CSAwallace_cska32_and_10_12 ^ u_CSAwallace_cska32_and_9_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa22_and0 = u_CSAwallace_cska32_and_10_12 & u_CSAwallace_cska32_and_9_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_and_8_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa22_and1 = u_CSAwallace_cska32_csa4_csa_component_fa22_xor0 & u_CSAwallace_cska32_and_8_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa22_or0 = u_CSAwallace_cska32_csa4_csa_component_fa22_and0 | u_CSAwallace_cska32_csa4_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa23_xor0 = u_CSAwallace_cska32_and_11_12 ^ u_CSAwallace_cska32_and_10_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa23_and0 = u_CSAwallace_cska32_and_11_12 & u_CSAwallace_cska32_and_10_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_and_9_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa23_and1 = u_CSAwallace_cska32_csa4_csa_component_fa23_xor0 & u_CSAwallace_cska32_and_9_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa23_or0 = u_CSAwallace_cska32_csa4_csa_component_fa23_and0 | u_CSAwallace_cska32_csa4_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa24_xor0 = u_CSAwallace_cska32_and_12_12 ^ u_CSAwallace_cska32_and_11_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa24_and0 = u_CSAwallace_cska32_and_12_12 & u_CSAwallace_cska32_and_11_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_and_10_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa24_and1 = u_CSAwallace_cska32_csa4_csa_component_fa24_xor0 & u_CSAwallace_cska32_and_10_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa24_or0 = u_CSAwallace_cska32_csa4_csa_component_fa24_and0 | u_CSAwallace_cska32_csa4_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_13_12 ^ u_CSAwallace_cska32_and_12_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa25_and0 = u_CSAwallace_cska32_and_13_12 & u_CSAwallace_cska32_and_12_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_and_11_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa25_and1 = u_CSAwallace_cska32_csa4_csa_component_fa25_xor0 & u_CSAwallace_cska32_and_11_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa25_or0 = u_CSAwallace_cska32_csa4_csa_component_fa25_and0 | u_CSAwallace_cska32_csa4_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_14_12 ^ u_CSAwallace_cska32_and_13_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa26_and0 = u_CSAwallace_cska32_and_14_12 & u_CSAwallace_cska32_and_13_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_12_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa26_and1 = u_CSAwallace_cska32_csa4_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_12_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa26_or0 = u_CSAwallace_cska32_csa4_csa_component_fa26_and0 | u_CSAwallace_cska32_csa4_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_15_12 ^ u_CSAwallace_cska32_and_14_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa27_and0 = u_CSAwallace_cska32_and_15_12 & u_CSAwallace_cska32_and_14_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_13_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa27_and1 = u_CSAwallace_cska32_csa4_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_13_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa27_or0 = u_CSAwallace_cska32_csa4_csa_component_fa27_and0 | u_CSAwallace_cska32_csa4_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_16_12 ^ u_CSAwallace_cska32_and_15_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa28_and0 = u_CSAwallace_cska32_and_16_12 & u_CSAwallace_cska32_and_15_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_14_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa28_and1 = u_CSAwallace_cska32_csa4_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_14_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa28_or0 = u_CSAwallace_cska32_csa4_csa_component_fa28_and0 | u_CSAwallace_cska32_csa4_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_17_12 ^ u_CSAwallace_cska32_and_16_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa29_and0 = u_CSAwallace_cska32_and_17_12 & u_CSAwallace_cska32_and_16_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_15_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa29_and1 = u_CSAwallace_cska32_csa4_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_15_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa29_or0 = u_CSAwallace_cska32_csa4_csa_component_fa29_and0 | u_CSAwallace_cska32_csa4_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_18_12 ^ u_CSAwallace_cska32_and_17_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa30_and0 = u_CSAwallace_cska32_and_18_12 & u_CSAwallace_cska32_and_17_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_16_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa30_and1 = u_CSAwallace_cska32_csa4_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_16_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa30_or0 = u_CSAwallace_cska32_csa4_csa_component_fa30_and0 | u_CSAwallace_cska32_csa4_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_19_12 ^ u_CSAwallace_cska32_and_18_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa31_and0 = u_CSAwallace_cska32_and_19_12 & u_CSAwallace_cska32_and_18_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_17_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa31_and1 = u_CSAwallace_cska32_csa4_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_17_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa31_or0 = u_CSAwallace_cska32_csa4_csa_component_fa31_and0 | u_CSAwallace_cska32_csa4_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_20_12 ^ u_CSAwallace_cska32_and_19_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa32_and0 = u_CSAwallace_cska32_and_20_12 & u_CSAwallace_cska32_and_19_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_18_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa32_and1 = u_CSAwallace_cska32_csa4_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_18_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa32_or0 = u_CSAwallace_cska32_csa4_csa_component_fa32_and0 | u_CSAwallace_cska32_csa4_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_21_12 ^ u_CSAwallace_cska32_and_20_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa33_and0 = u_CSAwallace_cska32_and_21_12 & u_CSAwallace_cska32_and_20_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_19_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa33_and1 = u_CSAwallace_cska32_csa4_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_19_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa33_or0 = u_CSAwallace_cska32_csa4_csa_component_fa33_and0 | u_CSAwallace_cska32_csa4_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_22_12 ^ u_CSAwallace_cska32_and_21_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa34_and0 = u_CSAwallace_cska32_and_22_12 & u_CSAwallace_cska32_and_21_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_20_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa34_and1 = u_CSAwallace_cska32_csa4_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_20_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa34_or0 = u_CSAwallace_cska32_csa4_csa_component_fa34_and0 | u_CSAwallace_cska32_csa4_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa35_xor0 = u_CSAwallace_cska32_and_23_12 ^ u_CSAwallace_cska32_and_22_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa35_and0 = u_CSAwallace_cska32_and_23_12 & u_CSAwallace_cska32_and_22_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_21_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa35_and1 = u_CSAwallace_cska32_csa4_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_21_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa35_or0 = u_CSAwallace_cska32_csa4_csa_component_fa35_and0 | u_CSAwallace_cska32_csa4_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa36_xor0 = u_CSAwallace_cska32_and_24_12 ^ u_CSAwallace_cska32_and_23_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa36_and0 = u_CSAwallace_cska32_and_24_12 & u_CSAwallace_cska32_and_23_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_22_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa36_and1 = u_CSAwallace_cska32_csa4_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_22_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa36_or0 = u_CSAwallace_cska32_csa4_csa_component_fa36_and0 | u_CSAwallace_cska32_csa4_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa37_xor0 = u_CSAwallace_cska32_and_25_12 ^ u_CSAwallace_cska32_and_24_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa37_and0 = u_CSAwallace_cska32_and_25_12 & u_CSAwallace_cska32_and_24_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_23_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa37_and1 = u_CSAwallace_cska32_csa4_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_23_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa37_or0 = u_CSAwallace_cska32_csa4_csa_component_fa37_and0 | u_CSAwallace_cska32_csa4_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa38_xor0 = u_CSAwallace_cska32_and_26_12 ^ u_CSAwallace_cska32_and_25_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa38_and0 = u_CSAwallace_cska32_and_26_12 & u_CSAwallace_cska32_and_25_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_24_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa38_and1 = u_CSAwallace_cska32_csa4_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_24_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa38_or0 = u_CSAwallace_cska32_csa4_csa_component_fa38_and0 | u_CSAwallace_cska32_csa4_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa39_xor0 = u_CSAwallace_cska32_and_27_12 ^ u_CSAwallace_cska32_and_26_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa39_and0 = u_CSAwallace_cska32_and_27_12 & u_CSAwallace_cska32_and_26_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_25_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa39_and1 = u_CSAwallace_cska32_csa4_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_25_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa39_or0 = u_CSAwallace_cska32_csa4_csa_component_fa39_and0 | u_CSAwallace_cska32_csa4_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa40_xor0 = u_CSAwallace_cska32_and_28_12 ^ u_CSAwallace_cska32_and_27_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa40_and0 = u_CSAwallace_cska32_and_28_12 & u_CSAwallace_cska32_and_27_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_26_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa40_and1 = u_CSAwallace_cska32_csa4_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_26_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa40_or0 = u_CSAwallace_cska32_csa4_csa_component_fa40_and0 | u_CSAwallace_cska32_csa4_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa41_xor0 = u_CSAwallace_cska32_and_29_12 ^ u_CSAwallace_cska32_and_28_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa41_and0 = u_CSAwallace_cska32_and_29_12 & u_CSAwallace_cska32_and_28_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_and_27_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa41_and1 = u_CSAwallace_cska32_csa4_csa_component_fa41_xor0 & u_CSAwallace_cska32_and_27_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa41_or0 = u_CSAwallace_cska32_csa4_csa_component_fa41_and0 | u_CSAwallace_cska32_csa4_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa42_xor0 = u_CSAwallace_cska32_and_30_12 ^ u_CSAwallace_cska32_and_29_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa42_and0 = u_CSAwallace_cska32_and_30_12 & u_CSAwallace_cska32_and_29_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_and_28_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa42_and1 = u_CSAwallace_cska32_csa4_csa_component_fa42_xor0 & u_CSAwallace_cska32_and_28_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa42_or0 = u_CSAwallace_cska32_csa4_csa_component_fa42_and0 | u_CSAwallace_cska32_csa4_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa43_xor0 = u_CSAwallace_cska32_and_31_12 ^ u_CSAwallace_cska32_and_30_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa43_and0 = u_CSAwallace_cska32_and_31_12 & u_CSAwallace_cska32_and_30_13;
  assign u_CSAwallace_cska32_csa4_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_and_29_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa43_and1 = u_CSAwallace_cska32_csa4_csa_component_fa43_xor0 & u_CSAwallace_cska32_and_29_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa43_or0 = u_CSAwallace_cska32_csa4_csa_component_fa43_and0 | u_CSAwallace_cska32_csa4_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa4_csa_component_fa44_xor1 = u_CSAwallace_cska32_and_31_13 ^ u_CSAwallace_cska32_and_30_14;
  assign u_CSAwallace_cska32_csa4_csa_component_fa44_and1 = u_CSAwallace_cska32_and_31_13 & u_CSAwallace_cska32_and_30_14;
  assign u_CSAwallace_cska32_csa5_csa_component_fa16_xor0 = u_CSAwallace_cska32_and_1_15 ^ u_CSAwallace_cska32_and_0_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa16_and0 = u_CSAwallace_cska32_and_1_15 & u_CSAwallace_cska32_and_0_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa17_xor0 = u_CSAwallace_cska32_and_2_15 ^ u_CSAwallace_cska32_and_1_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa17_and0 = u_CSAwallace_cska32_and_2_15 & u_CSAwallace_cska32_and_1_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_and_0_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa17_and1 = u_CSAwallace_cska32_csa5_csa_component_fa17_xor0 & u_CSAwallace_cska32_and_0_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa17_or0 = u_CSAwallace_cska32_csa5_csa_component_fa17_and0 | u_CSAwallace_cska32_csa5_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa18_xor0 = u_CSAwallace_cska32_and_3_15 ^ u_CSAwallace_cska32_and_2_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa18_and0 = u_CSAwallace_cska32_and_3_15 & u_CSAwallace_cska32_and_2_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_and_1_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa18_and1 = u_CSAwallace_cska32_csa5_csa_component_fa18_xor0 & u_CSAwallace_cska32_and_1_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa18_or0 = u_CSAwallace_cska32_csa5_csa_component_fa18_and0 | u_CSAwallace_cska32_csa5_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa19_xor0 = u_CSAwallace_cska32_and_4_15 ^ u_CSAwallace_cska32_and_3_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa19_and0 = u_CSAwallace_cska32_and_4_15 & u_CSAwallace_cska32_and_3_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_and_2_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa19_and1 = u_CSAwallace_cska32_csa5_csa_component_fa19_xor0 & u_CSAwallace_cska32_and_2_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa19_or0 = u_CSAwallace_cska32_csa5_csa_component_fa19_and0 | u_CSAwallace_cska32_csa5_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa20_xor0 = u_CSAwallace_cska32_and_5_15 ^ u_CSAwallace_cska32_and_4_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa20_and0 = u_CSAwallace_cska32_and_5_15 & u_CSAwallace_cska32_and_4_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_and_3_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa20_and1 = u_CSAwallace_cska32_csa5_csa_component_fa20_xor0 & u_CSAwallace_cska32_and_3_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa20_or0 = u_CSAwallace_cska32_csa5_csa_component_fa20_and0 | u_CSAwallace_cska32_csa5_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa21_xor0 = u_CSAwallace_cska32_and_6_15 ^ u_CSAwallace_cska32_and_5_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa21_and0 = u_CSAwallace_cska32_and_6_15 & u_CSAwallace_cska32_and_5_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_and_4_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa21_and1 = u_CSAwallace_cska32_csa5_csa_component_fa21_xor0 & u_CSAwallace_cska32_and_4_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa21_or0 = u_CSAwallace_cska32_csa5_csa_component_fa21_and0 | u_CSAwallace_cska32_csa5_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa22_xor0 = u_CSAwallace_cska32_and_7_15 ^ u_CSAwallace_cska32_and_6_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa22_and0 = u_CSAwallace_cska32_and_7_15 & u_CSAwallace_cska32_and_6_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_and_5_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa22_and1 = u_CSAwallace_cska32_csa5_csa_component_fa22_xor0 & u_CSAwallace_cska32_and_5_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa22_or0 = u_CSAwallace_cska32_csa5_csa_component_fa22_and0 | u_CSAwallace_cska32_csa5_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa23_xor0 = u_CSAwallace_cska32_and_8_15 ^ u_CSAwallace_cska32_and_7_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa23_and0 = u_CSAwallace_cska32_and_8_15 & u_CSAwallace_cska32_and_7_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_and_6_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa23_and1 = u_CSAwallace_cska32_csa5_csa_component_fa23_xor0 & u_CSAwallace_cska32_and_6_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa23_or0 = u_CSAwallace_cska32_csa5_csa_component_fa23_and0 | u_CSAwallace_cska32_csa5_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa24_xor0 = u_CSAwallace_cska32_and_9_15 ^ u_CSAwallace_cska32_and_8_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa24_and0 = u_CSAwallace_cska32_and_9_15 & u_CSAwallace_cska32_and_8_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_and_7_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa24_and1 = u_CSAwallace_cska32_csa5_csa_component_fa24_xor0 & u_CSAwallace_cska32_and_7_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa24_or0 = u_CSAwallace_cska32_csa5_csa_component_fa24_and0 | u_CSAwallace_cska32_csa5_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_10_15 ^ u_CSAwallace_cska32_and_9_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa25_and0 = u_CSAwallace_cska32_and_10_15 & u_CSAwallace_cska32_and_9_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_and_8_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa25_and1 = u_CSAwallace_cska32_csa5_csa_component_fa25_xor0 & u_CSAwallace_cska32_and_8_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa25_or0 = u_CSAwallace_cska32_csa5_csa_component_fa25_and0 | u_CSAwallace_cska32_csa5_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_11_15 ^ u_CSAwallace_cska32_and_10_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa26_and0 = u_CSAwallace_cska32_and_11_15 & u_CSAwallace_cska32_and_10_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_9_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa26_and1 = u_CSAwallace_cska32_csa5_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_9_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa26_or0 = u_CSAwallace_cska32_csa5_csa_component_fa26_and0 | u_CSAwallace_cska32_csa5_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_12_15 ^ u_CSAwallace_cska32_and_11_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa27_and0 = u_CSAwallace_cska32_and_12_15 & u_CSAwallace_cska32_and_11_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_10_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa27_and1 = u_CSAwallace_cska32_csa5_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_10_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa27_or0 = u_CSAwallace_cska32_csa5_csa_component_fa27_and0 | u_CSAwallace_cska32_csa5_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_13_15 ^ u_CSAwallace_cska32_and_12_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa28_and0 = u_CSAwallace_cska32_and_13_15 & u_CSAwallace_cska32_and_12_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_11_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa28_and1 = u_CSAwallace_cska32_csa5_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_11_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa28_or0 = u_CSAwallace_cska32_csa5_csa_component_fa28_and0 | u_CSAwallace_cska32_csa5_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_14_15 ^ u_CSAwallace_cska32_and_13_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa29_and0 = u_CSAwallace_cska32_and_14_15 & u_CSAwallace_cska32_and_13_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_12_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa29_and1 = u_CSAwallace_cska32_csa5_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_12_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa29_or0 = u_CSAwallace_cska32_csa5_csa_component_fa29_and0 | u_CSAwallace_cska32_csa5_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_15_15 ^ u_CSAwallace_cska32_and_14_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa30_and0 = u_CSAwallace_cska32_and_15_15 & u_CSAwallace_cska32_and_14_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_13_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa30_and1 = u_CSAwallace_cska32_csa5_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_13_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa30_or0 = u_CSAwallace_cska32_csa5_csa_component_fa30_and0 | u_CSAwallace_cska32_csa5_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_16_15 ^ u_CSAwallace_cska32_and_15_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa31_and0 = u_CSAwallace_cska32_and_16_15 & u_CSAwallace_cska32_and_15_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_14_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa31_and1 = u_CSAwallace_cska32_csa5_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_14_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa31_or0 = u_CSAwallace_cska32_csa5_csa_component_fa31_and0 | u_CSAwallace_cska32_csa5_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_17_15 ^ u_CSAwallace_cska32_and_16_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa32_and0 = u_CSAwallace_cska32_and_17_15 & u_CSAwallace_cska32_and_16_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_15_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa32_and1 = u_CSAwallace_cska32_csa5_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_15_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa32_or0 = u_CSAwallace_cska32_csa5_csa_component_fa32_and0 | u_CSAwallace_cska32_csa5_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_18_15 ^ u_CSAwallace_cska32_and_17_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa33_and0 = u_CSAwallace_cska32_and_18_15 & u_CSAwallace_cska32_and_17_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_16_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa33_and1 = u_CSAwallace_cska32_csa5_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_16_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa33_or0 = u_CSAwallace_cska32_csa5_csa_component_fa33_and0 | u_CSAwallace_cska32_csa5_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_19_15 ^ u_CSAwallace_cska32_and_18_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa34_and0 = u_CSAwallace_cska32_and_19_15 & u_CSAwallace_cska32_and_18_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_17_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa34_and1 = u_CSAwallace_cska32_csa5_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_17_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa34_or0 = u_CSAwallace_cska32_csa5_csa_component_fa34_and0 | u_CSAwallace_cska32_csa5_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa35_xor0 = u_CSAwallace_cska32_and_20_15 ^ u_CSAwallace_cska32_and_19_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa35_and0 = u_CSAwallace_cska32_and_20_15 & u_CSAwallace_cska32_and_19_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_18_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa35_and1 = u_CSAwallace_cska32_csa5_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_18_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa35_or0 = u_CSAwallace_cska32_csa5_csa_component_fa35_and0 | u_CSAwallace_cska32_csa5_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa36_xor0 = u_CSAwallace_cska32_and_21_15 ^ u_CSAwallace_cska32_and_20_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa36_and0 = u_CSAwallace_cska32_and_21_15 & u_CSAwallace_cska32_and_20_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_19_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa36_and1 = u_CSAwallace_cska32_csa5_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_19_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa36_or0 = u_CSAwallace_cska32_csa5_csa_component_fa36_and0 | u_CSAwallace_cska32_csa5_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa37_xor0 = u_CSAwallace_cska32_and_22_15 ^ u_CSAwallace_cska32_and_21_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa37_and0 = u_CSAwallace_cska32_and_22_15 & u_CSAwallace_cska32_and_21_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_20_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa37_and1 = u_CSAwallace_cska32_csa5_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_20_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa37_or0 = u_CSAwallace_cska32_csa5_csa_component_fa37_and0 | u_CSAwallace_cska32_csa5_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa38_xor0 = u_CSAwallace_cska32_and_23_15 ^ u_CSAwallace_cska32_and_22_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa38_and0 = u_CSAwallace_cska32_and_23_15 & u_CSAwallace_cska32_and_22_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_21_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa38_and1 = u_CSAwallace_cska32_csa5_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_21_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa38_or0 = u_CSAwallace_cska32_csa5_csa_component_fa38_and0 | u_CSAwallace_cska32_csa5_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa39_xor0 = u_CSAwallace_cska32_and_24_15 ^ u_CSAwallace_cska32_and_23_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa39_and0 = u_CSAwallace_cska32_and_24_15 & u_CSAwallace_cska32_and_23_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_22_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa39_and1 = u_CSAwallace_cska32_csa5_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_22_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa39_or0 = u_CSAwallace_cska32_csa5_csa_component_fa39_and0 | u_CSAwallace_cska32_csa5_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa40_xor0 = u_CSAwallace_cska32_and_25_15 ^ u_CSAwallace_cska32_and_24_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa40_and0 = u_CSAwallace_cska32_and_25_15 & u_CSAwallace_cska32_and_24_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_23_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa40_and1 = u_CSAwallace_cska32_csa5_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_23_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa40_or0 = u_CSAwallace_cska32_csa5_csa_component_fa40_and0 | u_CSAwallace_cska32_csa5_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa41_xor0 = u_CSAwallace_cska32_and_26_15 ^ u_CSAwallace_cska32_and_25_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa41_and0 = u_CSAwallace_cska32_and_26_15 & u_CSAwallace_cska32_and_25_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_and_24_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa41_and1 = u_CSAwallace_cska32_csa5_csa_component_fa41_xor0 & u_CSAwallace_cska32_and_24_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa41_or0 = u_CSAwallace_cska32_csa5_csa_component_fa41_and0 | u_CSAwallace_cska32_csa5_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa42_xor0 = u_CSAwallace_cska32_and_27_15 ^ u_CSAwallace_cska32_and_26_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa42_and0 = u_CSAwallace_cska32_and_27_15 & u_CSAwallace_cska32_and_26_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_and_25_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa42_and1 = u_CSAwallace_cska32_csa5_csa_component_fa42_xor0 & u_CSAwallace_cska32_and_25_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa42_or0 = u_CSAwallace_cska32_csa5_csa_component_fa42_and0 | u_CSAwallace_cska32_csa5_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa43_xor0 = u_CSAwallace_cska32_and_28_15 ^ u_CSAwallace_cska32_and_27_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa43_and0 = u_CSAwallace_cska32_and_28_15 & u_CSAwallace_cska32_and_27_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_and_26_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa43_and1 = u_CSAwallace_cska32_csa5_csa_component_fa43_xor0 & u_CSAwallace_cska32_and_26_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa43_or0 = u_CSAwallace_cska32_csa5_csa_component_fa43_and0 | u_CSAwallace_cska32_csa5_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa44_xor0 = u_CSAwallace_cska32_and_29_15 ^ u_CSAwallace_cska32_and_28_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa44_and0 = u_CSAwallace_cska32_and_29_15 & u_CSAwallace_cska32_and_28_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_and_27_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa44_and1 = u_CSAwallace_cska32_csa5_csa_component_fa44_xor0 & u_CSAwallace_cska32_and_27_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa44_or0 = u_CSAwallace_cska32_csa5_csa_component_fa44_and0 | u_CSAwallace_cska32_csa5_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa45_xor0 = u_CSAwallace_cska32_and_30_15 ^ u_CSAwallace_cska32_and_29_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa45_and0 = u_CSAwallace_cska32_and_30_15 & u_CSAwallace_cska32_and_29_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_and_28_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa45_and1 = u_CSAwallace_cska32_csa5_csa_component_fa45_xor0 & u_CSAwallace_cska32_and_28_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa45_or0 = u_CSAwallace_cska32_csa5_csa_component_fa45_and0 | u_CSAwallace_cska32_csa5_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa46_xor0 = u_CSAwallace_cska32_and_31_15 ^ u_CSAwallace_cska32_and_30_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa46_and0 = u_CSAwallace_cska32_and_31_15 & u_CSAwallace_cska32_and_30_16;
  assign u_CSAwallace_cska32_csa5_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_and_29_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa46_and1 = u_CSAwallace_cska32_csa5_csa_component_fa46_xor0 & u_CSAwallace_cska32_and_29_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa46_or0 = u_CSAwallace_cska32_csa5_csa_component_fa46_and0 | u_CSAwallace_cska32_csa5_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa5_csa_component_fa47_xor1 = u_CSAwallace_cska32_and_31_16 ^ u_CSAwallace_cska32_and_30_17;
  assign u_CSAwallace_cska32_csa5_csa_component_fa47_and1 = u_CSAwallace_cska32_and_31_16 & u_CSAwallace_cska32_and_30_17;
  assign u_CSAwallace_cska32_csa6_csa_component_fa19_xor0 = u_CSAwallace_cska32_and_1_18 ^ u_CSAwallace_cska32_and_0_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa19_and0 = u_CSAwallace_cska32_and_1_18 & u_CSAwallace_cska32_and_0_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa20_xor0 = u_CSAwallace_cska32_and_2_18 ^ u_CSAwallace_cska32_and_1_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa20_and0 = u_CSAwallace_cska32_and_2_18 & u_CSAwallace_cska32_and_1_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_and_0_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa20_and1 = u_CSAwallace_cska32_csa6_csa_component_fa20_xor0 & u_CSAwallace_cska32_and_0_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa20_or0 = u_CSAwallace_cska32_csa6_csa_component_fa20_and0 | u_CSAwallace_cska32_csa6_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa21_xor0 = u_CSAwallace_cska32_and_3_18 ^ u_CSAwallace_cska32_and_2_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa21_and0 = u_CSAwallace_cska32_and_3_18 & u_CSAwallace_cska32_and_2_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_and_1_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa21_and1 = u_CSAwallace_cska32_csa6_csa_component_fa21_xor0 & u_CSAwallace_cska32_and_1_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa21_or0 = u_CSAwallace_cska32_csa6_csa_component_fa21_and0 | u_CSAwallace_cska32_csa6_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa22_xor0 = u_CSAwallace_cska32_and_4_18 ^ u_CSAwallace_cska32_and_3_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa22_and0 = u_CSAwallace_cska32_and_4_18 & u_CSAwallace_cska32_and_3_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_and_2_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa22_and1 = u_CSAwallace_cska32_csa6_csa_component_fa22_xor0 & u_CSAwallace_cska32_and_2_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa22_or0 = u_CSAwallace_cska32_csa6_csa_component_fa22_and0 | u_CSAwallace_cska32_csa6_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa23_xor0 = u_CSAwallace_cska32_and_5_18 ^ u_CSAwallace_cska32_and_4_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa23_and0 = u_CSAwallace_cska32_and_5_18 & u_CSAwallace_cska32_and_4_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_and_3_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa23_and1 = u_CSAwallace_cska32_csa6_csa_component_fa23_xor0 & u_CSAwallace_cska32_and_3_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa23_or0 = u_CSAwallace_cska32_csa6_csa_component_fa23_and0 | u_CSAwallace_cska32_csa6_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa24_xor0 = u_CSAwallace_cska32_and_6_18 ^ u_CSAwallace_cska32_and_5_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa24_and0 = u_CSAwallace_cska32_and_6_18 & u_CSAwallace_cska32_and_5_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_and_4_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa24_and1 = u_CSAwallace_cska32_csa6_csa_component_fa24_xor0 & u_CSAwallace_cska32_and_4_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa24_or0 = u_CSAwallace_cska32_csa6_csa_component_fa24_and0 | u_CSAwallace_cska32_csa6_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_7_18 ^ u_CSAwallace_cska32_and_6_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa25_and0 = u_CSAwallace_cska32_and_7_18 & u_CSAwallace_cska32_and_6_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_and_5_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa25_and1 = u_CSAwallace_cska32_csa6_csa_component_fa25_xor0 & u_CSAwallace_cska32_and_5_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa25_or0 = u_CSAwallace_cska32_csa6_csa_component_fa25_and0 | u_CSAwallace_cska32_csa6_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_8_18 ^ u_CSAwallace_cska32_and_7_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa26_and0 = u_CSAwallace_cska32_and_8_18 & u_CSAwallace_cska32_and_7_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_6_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa26_and1 = u_CSAwallace_cska32_csa6_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_6_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa26_or0 = u_CSAwallace_cska32_csa6_csa_component_fa26_and0 | u_CSAwallace_cska32_csa6_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_9_18 ^ u_CSAwallace_cska32_and_8_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa27_and0 = u_CSAwallace_cska32_and_9_18 & u_CSAwallace_cska32_and_8_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_7_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa27_and1 = u_CSAwallace_cska32_csa6_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_7_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa27_or0 = u_CSAwallace_cska32_csa6_csa_component_fa27_and0 | u_CSAwallace_cska32_csa6_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_10_18 ^ u_CSAwallace_cska32_and_9_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa28_and0 = u_CSAwallace_cska32_and_10_18 & u_CSAwallace_cska32_and_9_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_8_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa28_and1 = u_CSAwallace_cska32_csa6_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_8_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa28_or0 = u_CSAwallace_cska32_csa6_csa_component_fa28_and0 | u_CSAwallace_cska32_csa6_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_11_18 ^ u_CSAwallace_cska32_and_10_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa29_and0 = u_CSAwallace_cska32_and_11_18 & u_CSAwallace_cska32_and_10_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_9_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa29_and1 = u_CSAwallace_cska32_csa6_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_9_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa29_or0 = u_CSAwallace_cska32_csa6_csa_component_fa29_and0 | u_CSAwallace_cska32_csa6_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_12_18 ^ u_CSAwallace_cska32_and_11_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa30_and0 = u_CSAwallace_cska32_and_12_18 & u_CSAwallace_cska32_and_11_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_10_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa30_and1 = u_CSAwallace_cska32_csa6_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_10_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa30_or0 = u_CSAwallace_cska32_csa6_csa_component_fa30_and0 | u_CSAwallace_cska32_csa6_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_13_18 ^ u_CSAwallace_cska32_and_12_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa31_and0 = u_CSAwallace_cska32_and_13_18 & u_CSAwallace_cska32_and_12_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_11_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa31_and1 = u_CSAwallace_cska32_csa6_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_11_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa31_or0 = u_CSAwallace_cska32_csa6_csa_component_fa31_and0 | u_CSAwallace_cska32_csa6_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_14_18 ^ u_CSAwallace_cska32_and_13_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa32_and0 = u_CSAwallace_cska32_and_14_18 & u_CSAwallace_cska32_and_13_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_12_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa32_and1 = u_CSAwallace_cska32_csa6_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_12_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa32_or0 = u_CSAwallace_cska32_csa6_csa_component_fa32_and0 | u_CSAwallace_cska32_csa6_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_15_18 ^ u_CSAwallace_cska32_and_14_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa33_and0 = u_CSAwallace_cska32_and_15_18 & u_CSAwallace_cska32_and_14_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_13_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa33_and1 = u_CSAwallace_cska32_csa6_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_13_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa33_or0 = u_CSAwallace_cska32_csa6_csa_component_fa33_and0 | u_CSAwallace_cska32_csa6_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_16_18 ^ u_CSAwallace_cska32_and_15_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa34_and0 = u_CSAwallace_cska32_and_16_18 & u_CSAwallace_cska32_and_15_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_14_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa34_and1 = u_CSAwallace_cska32_csa6_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_14_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa34_or0 = u_CSAwallace_cska32_csa6_csa_component_fa34_and0 | u_CSAwallace_cska32_csa6_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa35_xor0 = u_CSAwallace_cska32_and_17_18 ^ u_CSAwallace_cska32_and_16_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa35_and0 = u_CSAwallace_cska32_and_17_18 & u_CSAwallace_cska32_and_16_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_15_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa35_and1 = u_CSAwallace_cska32_csa6_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_15_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa35_or0 = u_CSAwallace_cska32_csa6_csa_component_fa35_and0 | u_CSAwallace_cska32_csa6_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa36_xor0 = u_CSAwallace_cska32_and_18_18 ^ u_CSAwallace_cska32_and_17_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa36_and0 = u_CSAwallace_cska32_and_18_18 & u_CSAwallace_cska32_and_17_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_16_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa36_and1 = u_CSAwallace_cska32_csa6_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_16_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa36_or0 = u_CSAwallace_cska32_csa6_csa_component_fa36_and0 | u_CSAwallace_cska32_csa6_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa37_xor0 = u_CSAwallace_cska32_and_19_18 ^ u_CSAwallace_cska32_and_18_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa37_and0 = u_CSAwallace_cska32_and_19_18 & u_CSAwallace_cska32_and_18_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_17_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa37_and1 = u_CSAwallace_cska32_csa6_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_17_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa37_or0 = u_CSAwallace_cska32_csa6_csa_component_fa37_and0 | u_CSAwallace_cska32_csa6_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa38_xor0 = u_CSAwallace_cska32_and_20_18 ^ u_CSAwallace_cska32_and_19_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa38_and0 = u_CSAwallace_cska32_and_20_18 & u_CSAwallace_cska32_and_19_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_18_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa38_and1 = u_CSAwallace_cska32_csa6_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_18_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa38_or0 = u_CSAwallace_cska32_csa6_csa_component_fa38_and0 | u_CSAwallace_cska32_csa6_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa39_xor0 = u_CSAwallace_cska32_and_21_18 ^ u_CSAwallace_cska32_and_20_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa39_and0 = u_CSAwallace_cska32_and_21_18 & u_CSAwallace_cska32_and_20_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_19_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa39_and1 = u_CSAwallace_cska32_csa6_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_19_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa39_or0 = u_CSAwallace_cska32_csa6_csa_component_fa39_and0 | u_CSAwallace_cska32_csa6_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa40_xor0 = u_CSAwallace_cska32_and_22_18 ^ u_CSAwallace_cska32_and_21_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa40_and0 = u_CSAwallace_cska32_and_22_18 & u_CSAwallace_cska32_and_21_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_20_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa40_and1 = u_CSAwallace_cska32_csa6_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_20_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa40_or0 = u_CSAwallace_cska32_csa6_csa_component_fa40_and0 | u_CSAwallace_cska32_csa6_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa41_xor0 = u_CSAwallace_cska32_and_23_18 ^ u_CSAwallace_cska32_and_22_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa41_and0 = u_CSAwallace_cska32_and_23_18 & u_CSAwallace_cska32_and_22_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_and_21_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa41_and1 = u_CSAwallace_cska32_csa6_csa_component_fa41_xor0 & u_CSAwallace_cska32_and_21_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa41_or0 = u_CSAwallace_cska32_csa6_csa_component_fa41_and0 | u_CSAwallace_cska32_csa6_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa42_xor0 = u_CSAwallace_cska32_and_24_18 ^ u_CSAwallace_cska32_and_23_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa42_and0 = u_CSAwallace_cska32_and_24_18 & u_CSAwallace_cska32_and_23_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_and_22_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa42_and1 = u_CSAwallace_cska32_csa6_csa_component_fa42_xor0 & u_CSAwallace_cska32_and_22_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa42_or0 = u_CSAwallace_cska32_csa6_csa_component_fa42_and0 | u_CSAwallace_cska32_csa6_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa43_xor0 = u_CSAwallace_cska32_and_25_18 ^ u_CSAwallace_cska32_and_24_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa43_and0 = u_CSAwallace_cska32_and_25_18 & u_CSAwallace_cska32_and_24_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_and_23_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa43_and1 = u_CSAwallace_cska32_csa6_csa_component_fa43_xor0 & u_CSAwallace_cska32_and_23_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa43_or0 = u_CSAwallace_cska32_csa6_csa_component_fa43_and0 | u_CSAwallace_cska32_csa6_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa44_xor0 = u_CSAwallace_cska32_and_26_18 ^ u_CSAwallace_cska32_and_25_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa44_and0 = u_CSAwallace_cska32_and_26_18 & u_CSAwallace_cska32_and_25_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_and_24_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa44_and1 = u_CSAwallace_cska32_csa6_csa_component_fa44_xor0 & u_CSAwallace_cska32_and_24_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa44_or0 = u_CSAwallace_cska32_csa6_csa_component_fa44_and0 | u_CSAwallace_cska32_csa6_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa45_xor0 = u_CSAwallace_cska32_and_27_18 ^ u_CSAwallace_cska32_and_26_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa45_and0 = u_CSAwallace_cska32_and_27_18 & u_CSAwallace_cska32_and_26_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_and_25_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa45_and1 = u_CSAwallace_cska32_csa6_csa_component_fa45_xor0 & u_CSAwallace_cska32_and_25_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa45_or0 = u_CSAwallace_cska32_csa6_csa_component_fa45_and0 | u_CSAwallace_cska32_csa6_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa46_xor0 = u_CSAwallace_cska32_and_28_18 ^ u_CSAwallace_cska32_and_27_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa46_and0 = u_CSAwallace_cska32_and_28_18 & u_CSAwallace_cska32_and_27_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_and_26_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa46_and1 = u_CSAwallace_cska32_csa6_csa_component_fa46_xor0 & u_CSAwallace_cska32_and_26_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa46_or0 = u_CSAwallace_cska32_csa6_csa_component_fa46_and0 | u_CSAwallace_cska32_csa6_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa47_xor0 = u_CSAwallace_cska32_and_29_18 ^ u_CSAwallace_cska32_and_28_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa47_and0 = u_CSAwallace_cska32_and_29_18 & u_CSAwallace_cska32_and_28_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_and_27_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa47_and1 = u_CSAwallace_cska32_csa6_csa_component_fa47_xor0 & u_CSAwallace_cska32_and_27_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa47_or0 = u_CSAwallace_cska32_csa6_csa_component_fa47_and0 | u_CSAwallace_cska32_csa6_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa48_xor0 = u_CSAwallace_cska32_and_30_18 ^ u_CSAwallace_cska32_and_29_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa48_and0 = u_CSAwallace_cska32_and_30_18 & u_CSAwallace_cska32_and_29_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_and_28_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa48_and1 = u_CSAwallace_cska32_csa6_csa_component_fa48_xor0 & u_CSAwallace_cska32_and_28_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa48_or0 = u_CSAwallace_cska32_csa6_csa_component_fa48_and0 | u_CSAwallace_cska32_csa6_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa49_xor0 = u_CSAwallace_cska32_and_31_18 ^ u_CSAwallace_cska32_and_30_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa49_and0 = u_CSAwallace_cska32_and_31_18 & u_CSAwallace_cska32_and_30_19;
  assign u_CSAwallace_cska32_csa6_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa6_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_and_29_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa49_and1 = u_CSAwallace_cska32_csa6_csa_component_fa49_xor0 & u_CSAwallace_cska32_and_29_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa49_or0 = u_CSAwallace_cska32_csa6_csa_component_fa49_and0 | u_CSAwallace_cska32_csa6_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa6_csa_component_fa50_xor1 = u_CSAwallace_cska32_and_31_19 ^ u_CSAwallace_cska32_and_30_20;
  assign u_CSAwallace_cska32_csa6_csa_component_fa50_and1 = u_CSAwallace_cska32_and_31_19 & u_CSAwallace_cska32_and_30_20;
  assign u_CSAwallace_cska32_csa7_csa_component_fa22_xor0 = u_CSAwallace_cska32_and_1_21 ^ u_CSAwallace_cska32_and_0_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa22_and0 = u_CSAwallace_cska32_and_1_21 & u_CSAwallace_cska32_and_0_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa23_xor0 = u_CSAwallace_cska32_and_2_21 ^ u_CSAwallace_cska32_and_1_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa23_and0 = u_CSAwallace_cska32_and_2_21 & u_CSAwallace_cska32_and_1_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_and_0_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa23_and1 = u_CSAwallace_cska32_csa7_csa_component_fa23_xor0 & u_CSAwallace_cska32_and_0_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa23_or0 = u_CSAwallace_cska32_csa7_csa_component_fa23_and0 | u_CSAwallace_cska32_csa7_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa24_xor0 = u_CSAwallace_cska32_and_3_21 ^ u_CSAwallace_cska32_and_2_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa24_and0 = u_CSAwallace_cska32_and_3_21 & u_CSAwallace_cska32_and_2_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_and_1_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa24_and1 = u_CSAwallace_cska32_csa7_csa_component_fa24_xor0 & u_CSAwallace_cska32_and_1_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa24_or0 = u_CSAwallace_cska32_csa7_csa_component_fa24_and0 | u_CSAwallace_cska32_csa7_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_4_21 ^ u_CSAwallace_cska32_and_3_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa25_and0 = u_CSAwallace_cska32_and_4_21 & u_CSAwallace_cska32_and_3_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_and_2_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa25_and1 = u_CSAwallace_cska32_csa7_csa_component_fa25_xor0 & u_CSAwallace_cska32_and_2_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa25_or0 = u_CSAwallace_cska32_csa7_csa_component_fa25_and0 | u_CSAwallace_cska32_csa7_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_5_21 ^ u_CSAwallace_cska32_and_4_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa26_and0 = u_CSAwallace_cska32_and_5_21 & u_CSAwallace_cska32_and_4_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_3_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa26_and1 = u_CSAwallace_cska32_csa7_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_3_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa26_or0 = u_CSAwallace_cska32_csa7_csa_component_fa26_and0 | u_CSAwallace_cska32_csa7_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_6_21 ^ u_CSAwallace_cska32_and_5_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa27_and0 = u_CSAwallace_cska32_and_6_21 & u_CSAwallace_cska32_and_5_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_4_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa27_and1 = u_CSAwallace_cska32_csa7_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_4_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa27_or0 = u_CSAwallace_cska32_csa7_csa_component_fa27_and0 | u_CSAwallace_cska32_csa7_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_7_21 ^ u_CSAwallace_cska32_and_6_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa28_and0 = u_CSAwallace_cska32_and_7_21 & u_CSAwallace_cska32_and_6_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_5_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa28_and1 = u_CSAwallace_cska32_csa7_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_5_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa28_or0 = u_CSAwallace_cska32_csa7_csa_component_fa28_and0 | u_CSAwallace_cska32_csa7_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_8_21 ^ u_CSAwallace_cska32_and_7_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa29_and0 = u_CSAwallace_cska32_and_8_21 & u_CSAwallace_cska32_and_7_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_6_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa29_and1 = u_CSAwallace_cska32_csa7_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_6_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa29_or0 = u_CSAwallace_cska32_csa7_csa_component_fa29_and0 | u_CSAwallace_cska32_csa7_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_9_21 ^ u_CSAwallace_cska32_and_8_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa30_and0 = u_CSAwallace_cska32_and_9_21 & u_CSAwallace_cska32_and_8_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_7_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa30_and1 = u_CSAwallace_cska32_csa7_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_7_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa30_or0 = u_CSAwallace_cska32_csa7_csa_component_fa30_and0 | u_CSAwallace_cska32_csa7_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_10_21 ^ u_CSAwallace_cska32_and_9_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa31_and0 = u_CSAwallace_cska32_and_10_21 & u_CSAwallace_cska32_and_9_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_8_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa31_and1 = u_CSAwallace_cska32_csa7_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_8_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa31_or0 = u_CSAwallace_cska32_csa7_csa_component_fa31_and0 | u_CSAwallace_cska32_csa7_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_11_21 ^ u_CSAwallace_cska32_and_10_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa32_and0 = u_CSAwallace_cska32_and_11_21 & u_CSAwallace_cska32_and_10_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_9_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa32_and1 = u_CSAwallace_cska32_csa7_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_9_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa32_or0 = u_CSAwallace_cska32_csa7_csa_component_fa32_and0 | u_CSAwallace_cska32_csa7_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_12_21 ^ u_CSAwallace_cska32_and_11_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa33_and0 = u_CSAwallace_cska32_and_12_21 & u_CSAwallace_cska32_and_11_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_10_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa33_and1 = u_CSAwallace_cska32_csa7_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_10_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa33_or0 = u_CSAwallace_cska32_csa7_csa_component_fa33_and0 | u_CSAwallace_cska32_csa7_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_13_21 ^ u_CSAwallace_cska32_and_12_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa34_and0 = u_CSAwallace_cska32_and_13_21 & u_CSAwallace_cska32_and_12_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_11_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa34_and1 = u_CSAwallace_cska32_csa7_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_11_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa34_or0 = u_CSAwallace_cska32_csa7_csa_component_fa34_and0 | u_CSAwallace_cska32_csa7_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa35_xor0 = u_CSAwallace_cska32_and_14_21 ^ u_CSAwallace_cska32_and_13_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa35_and0 = u_CSAwallace_cska32_and_14_21 & u_CSAwallace_cska32_and_13_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_12_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa35_and1 = u_CSAwallace_cska32_csa7_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_12_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa35_or0 = u_CSAwallace_cska32_csa7_csa_component_fa35_and0 | u_CSAwallace_cska32_csa7_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa36_xor0 = u_CSAwallace_cska32_and_15_21 ^ u_CSAwallace_cska32_and_14_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa36_and0 = u_CSAwallace_cska32_and_15_21 & u_CSAwallace_cska32_and_14_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_13_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa36_and1 = u_CSAwallace_cska32_csa7_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_13_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa36_or0 = u_CSAwallace_cska32_csa7_csa_component_fa36_and0 | u_CSAwallace_cska32_csa7_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa37_xor0 = u_CSAwallace_cska32_and_16_21 ^ u_CSAwallace_cska32_and_15_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa37_and0 = u_CSAwallace_cska32_and_16_21 & u_CSAwallace_cska32_and_15_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_14_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa37_and1 = u_CSAwallace_cska32_csa7_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_14_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa37_or0 = u_CSAwallace_cska32_csa7_csa_component_fa37_and0 | u_CSAwallace_cska32_csa7_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa38_xor0 = u_CSAwallace_cska32_and_17_21 ^ u_CSAwallace_cska32_and_16_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa38_and0 = u_CSAwallace_cska32_and_17_21 & u_CSAwallace_cska32_and_16_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_15_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa38_and1 = u_CSAwallace_cska32_csa7_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_15_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa38_or0 = u_CSAwallace_cska32_csa7_csa_component_fa38_and0 | u_CSAwallace_cska32_csa7_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa39_xor0 = u_CSAwallace_cska32_and_18_21 ^ u_CSAwallace_cska32_and_17_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa39_and0 = u_CSAwallace_cska32_and_18_21 & u_CSAwallace_cska32_and_17_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_16_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa39_and1 = u_CSAwallace_cska32_csa7_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_16_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa39_or0 = u_CSAwallace_cska32_csa7_csa_component_fa39_and0 | u_CSAwallace_cska32_csa7_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa40_xor0 = u_CSAwallace_cska32_and_19_21 ^ u_CSAwallace_cska32_and_18_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa40_and0 = u_CSAwallace_cska32_and_19_21 & u_CSAwallace_cska32_and_18_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_17_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa40_and1 = u_CSAwallace_cska32_csa7_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_17_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa40_or0 = u_CSAwallace_cska32_csa7_csa_component_fa40_and0 | u_CSAwallace_cska32_csa7_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa41_xor0 = u_CSAwallace_cska32_and_20_21 ^ u_CSAwallace_cska32_and_19_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa41_and0 = u_CSAwallace_cska32_and_20_21 & u_CSAwallace_cska32_and_19_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_and_18_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa41_and1 = u_CSAwallace_cska32_csa7_csa_component_fa41_xor0 & u_CSAwallace_cska32_and_18_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa41_or0 = u_CSAwallace_cska32_csa7_csa_component_fa41_and0 | u_CSAwallace_cska32_csa7_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa42_xor0 = u_CSAwallace_cska32_and_21_21 ^ u_CSAwallace_cska32_and_20_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa42_and0 = u_CSAwallace_cska32_and_21_21 & u_CSAwallace_cska32_and_20_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_and_19_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa42_and1 = u_CSAwallace_cska32_csa7_csa_component_fa42_xor0 & u_CSAwallace_cska32_and_19_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa42_or0 = u_CSAwallace_cska32_csa7_csa_component_fa42_and0 | u_CSAwallace_cska32_csa7_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa43_xor0 = u_CSAwallace_cska32_and_22_21 ^ u_CSAwallace_cska32_and_21_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa43_and0 = u_CSAwallace_cska32_and_22_21 & u_CSAwallace_cska32_and_21_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_and_20_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa43_and1 = u_CSAwallace_cska32_csa7_csa_component_fa43_xor0 & u_CSAwallace_cska32_and_20_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa43_or0 = u_CSAwallace_cska32_csa7_csa_component_fa43_and0 | u_CSAwallace_cska32_csa7_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa44_xor0 = u_CSAwallace_cska32_and_23_21 ^ u_CSAwallace_cska32_and_22_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa44_and0 = u_CSAwallace_cska32_and_23_21 & u_CSAwallace_cska32_and_22_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_and_21_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa44_and1 = u_CSAwallace_cska32_csa7_csa_component_fa44_xor0 & u_CSAwallace_cska32_and_21_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa44_or0 = u_CSAwallace_cska32_csa7_csa_component_fa44_and0 | u_CSAwallace_cska32_csa7_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa45_xor0 = u_CSAwallace_cska32_and_24_21 ^ u_CSAwallace_cska32_and_23_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa45_and0 = u_CSAwallace_cska32_and_24_21 & u_CSAwallace_cska32_and_23_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_and_22_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa45_and1 = u_CSAwallace_cska32_csa7_csa_component_fa45_xor0 & u_CSAwallace_cska32_and_22_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa45_or0 = u_CSAwallace_cska32_csa7_csa_component_fa45_and0 | u_CSAwallace_cska32_csa7_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa46_xor0 = u_CSAwallace_cska32_and_25_21 ^ u_CSAwallace_cska32_and_24_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa46_and0 = u_CSAwallace_cska32_and_25_21 & u_CSAwallace_cska32_and_24_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_and_23_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa46_and1 = u_CSAwallace_cska32_csa7_csa_component_fa46_xor0 & u_CSAwallace_cska32_and_23_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa46_or0 = u_CSAwallace_cska32_csa7_csa_component_fa46_and0 | u_CSAwallace_cska32_csa7_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa47_xor0 = u_CSAwallace_cska32_and_26_21 ^ u_CSAwallace_cska32_and_25_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa47_and0 = u_CSAwallace_cska32_and_26_21 & u_CSAwallace_cska32_and_25_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_and_24_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa47_and1 = u_CSAwallace_cska32_csa7_csa_component_fa47_xor0 & u_CSAwallace_cska32_and_24_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa47_or0 = u_CSAwallace_cska32_csa7_csa_component_fa47_and0 | u_CSAwallace_cska32_csa7_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa48_xor0 = u_CSAwallace_cska32_and_27_21 ^ u_CSAwallace_cska32_and_26_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa48_and0 = u_CSAwallace_cska32_and_27_21 & u_CSAwallace_cska32_and_26_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_and_25_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa48_and1 = u_CSAwallace_cska32_csa7_csa_component_fa48_xor0 & u_CSAwallace_cska32_and_25_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa48_or0 = u_CSAwallace_cska32_csa7_csa_component_fa48_and0 | u_CSAwallace_cska32_csa7_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa49_xor0 = u_CSAwallace_cska32_and_28_21 ^ u_CSAwallace_cska32_and_27_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa49_and0 = u_CSAwallace_cska32_and_28_21 & u_CSAwallace_cska32_and_27_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_and_26_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa49_and1 = u_CSAwallace_cska32_csa7_csa_component_fa49_xor0 & u_CSAwallace_cska32_and_26_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa49_or0 = u_CSAwallace_cska32_csa7_csa_component_fa49_and0 | u_CSAwallace_cska32_csa7_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa50_xor0 = u_CSAwallace_cska32_and_29_21 ^ u_CSAwallace_cska32_and_28_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa50_and0 = u_CSAwallace_cska32_and_29_21 & u_CSAwallace_cska32_and_28_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_and_27_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa50_and1 = u_CSAwallace_cska32_csa7_csa_component_fa50_xor0 & u_CSAwallace_cska32_and_27_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa50_or0 = u_CSAwallace_cska32_csa7_csa_component_fa50_and0 | u_CSAwallace_cska32_csa7_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa51_xor0 = u_CSAwallace_cska32_and_30_21 ^ u_CSAwallace_cska32_and_29_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa51_and0 = u_CSAwallace_cska32_and_30_21 & u_CSAwallace_cska32_and_29_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_and_28_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa51_and1 = u_CSAwallace_cska32_csa7_csa_component_fa51_xor0 & u_CSAwallace_cska32_and_28_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa51_or0 = u_CSAwallace_cska32_csa7_csa_component_fa51_and0 | u_CSAwallace_cska32_csa7_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa52_xor0 = u_CSAwallace_cska32_and_31_21 ^ u_CSAwallace_cska32_and_30_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa52_and0 = u_CSAwallace_cska32_and_31_21 & u_CSAwallace_cska32_and_30_22;
  assign u_CSAwallace_cska32_csa7_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_and_29_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa52_and1 = u_CSAwallace_cska32_csa7_csa_component_fa52_xor0 & u_CSAwallace_cska32_and_29_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa52_or0 = u_CSAwallace_cska32_csa7_csa_component_fa52_and0 | u_CSAwallace_cska32_csa7_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa7_csa_component_fa53_xor1 = u_CSAwallace_cska32_and_31_22 ^ u_CSAwallace_cska32_and_30_23;
  assign u_CSAwallace_cska32_csa7_csa_component_fa53_and1 = u_CSAwallace_cska32_and_31_22 & u_CSAwallace_cska32_and_30_23;
  assign u_CSAwallace_cska32_csa8_csa_component_fa25_xor0 = u_CSAwallace_cska32_and_1_24 ^ u_CSAwallace_cska32_and_0_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa25_and0 = u_CSAwallace_cska32_and_1_24 & u_CSAwallace_cska32_and_0_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa26_xor0 = u_CSAwallace_cska32_and_2_24 ^ u_CSAwallace_cska32_and_1_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa26_and0 = u_CSAwallace_cska32_and_2_24 & u_CSAwallace_cska32_and_1_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_and_0_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa26_and1 = u_CSAwallace_cska32_csa8_csa_component_fa26_xor0 & u_CSAwallace_cska32_and_0_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa26_or0 = u_CSAwallace_cska32_csa8_csa_component_fa26_and0 | u_CSAwallace_cska32_csa8_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa27_xor0 = u_CSAwallace_cska32_and_3_24 ^ u_CSAwallace_cska32_and_2_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa27_and0 = u_CSAwallace_cska32_and_3_24 & u_CSAwallace_cska32_and_2_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_1_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa27_and1 = u_CSAwallace_cska32_csa8_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_1_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa27_or0 = u_CSAwallace_cska32_csa8_csa_component_fa27_and0 | u_CSAwallace_cska32_csa8_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_4_24 ^ u_CSAwallace_cska32_and_3_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa28_and0 = u_CSAwallace_cska32_and_4_24 & u_CSAwallace_cska32_and_3_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_and_2_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa28_and1 = u_CSAwallace_cska32_csa8_csa_component_fa28_xor0 & u_CSAwallace_cska32_and_2_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa28_or0 = u_CSAwallace_cska32_csa8_csa_component_fa28_and0 | u_CSAwallace_cska32_csa8_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_5_24 ^ u_CSAwallace_cska32_and_4_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa29_and0 = u_CSAwallace_cska32_and_5_24 & u_CSAwallace_cska32_and_4_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_3_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa29_and1 = u_CSAwallace_cska32_csa8_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_3_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa29_or0 = u_CSAwallace_cska32_csa8_csa_component_fa29_and0 | u_CSAwallace_cska32_csa8_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_6_24 ^ u_CSAwallace_cska32_and_5_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa30_and0 = u_CSAwallace_cska32_and_6_24 & u_CSAwallace_cska32_and_5_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_4_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa30_and1 = u_CSAwallace_cska32_csa8_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_4_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa30_or0 = u_CSAwallace_cska32_csa8_csa_component_fa30_and0 | u_CSAwallace_cska32_csa8_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_7_24 ^ u_CSAwallace_cska32_and_6_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa31_and0 = u_CSAwallace_cska32_and_7_24 & u_CSAwallace_cska32_and_6_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_5_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa31_and1 = u_CSAwallace_cska32_csa8_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_5_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa31_or0 = u_CSAwallace_cska32_csa8_csa_component_fa31_and0 | u_CSAwallace_cska32_csa8_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_8_24 ^ u_CSAwallace_cska32_and_7_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa32_and0 = u_CSAwallace_cska32_and_8_24 & u_CSAwallace_cska32_and_7_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_6_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa32_and1 = u_CSAwallace_cska32_csa8_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_6_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa32_or0 = u_CSAwallace_cska32_csa8_csa_component_fa32_and0 | u_CSAwallace_cska32_csa8_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_9_24 ^ u_CSAwallace_cska32_and_8_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa33_and0 = u_CSAwallace_cska32_and_9_24 & u_CSAwallace_cska32_and_8_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_7_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa33_and1 = u_CSAwallace_cska32_csa8_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_7_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa33_or0 = u_CSAwallace_cska32_csa8_csa_component_fa33_and0 | u_CSAwallace_cska32_csa8_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_10_24 ^ u_CSAwallace_cska32_and_9_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa34_and0 = u_CSAwallace_cska32_and_10_24 & u_CSAwallace_cska32_and_9_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_8_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa34_and1 = u_CSAwallace_cska32_csa8_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_8_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa34_or0 = u_CSAwallace_cska32_csa8_csa_component_fa34_and0 | u_CSAwallace_cska32_csa8_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa35_xor0 = u_CSAwallace_cska32_and_11_24 ^ u_CSAwallace_cska32_and_10_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa35_and0 = u_CSAwallace_cska32_and_11_24 & u_CSAwallace_cska32_and_10_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_9_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa35_and1 = u_CSAwallace_cska32_csa8_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_9_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa35_or0 = u_CSAwallace_cska32_csa8_csa_component_fa35_and0 | u_CSAwallace_cska32_csa8_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa36_xor0 = u_CSAwallace_cska32_and_12_24 ^ u_CSAwallace_cska32_and_11_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa36_and0 = u_CSAwallace_cska32_and_12_24 & u_CSAwallace_cska32_and_11_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_10_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa36_and1 = u_CSAwallace_cska32_csa8_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_10_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa36_or0 = u_CSAwallace_cska32_csa8_csa_component_fa36_and0 | u_CSAwallace_cska32_csa8_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa37_xor0 = u_CSAwallace_cska32_and_13_24 ^ u_CSAwallace_cska32_and_12_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa37_and0 = u_CSAwallace_cska32_and_13_24 & u_CSAwallace_cska32_and_12_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_11_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa37_and1 = u_CSAwallace_cska32_csa8_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_11_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa37_or0 = u_CSAwallace_cska32_csa8_csa_component_fa37_and0 | u_CSAwallace_cska32_csa8_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa38_xor0 = u_CSAwallace_cska32_and_14_24 ^ u_CSAwallace_cska32_and_13_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa38_and0 = u_CSAwallace_cska32_and_14_24 & u_CSAwallace_cska32_and_13_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_12_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa38_and1 = u_CSAwallace_cska32_csa8_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_12_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa38_or0 = u_CSAwallace_cska32_csa8_csa_component_fa38_and0 | u_CSAwallace_cska32_csa8_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa39_xor0 = u_CSAwallace_cska32_and_15_24 ^ u_CSAwallace_cska32_and_14_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa39_and0 = u_CSAwallace_cska32_and_15_24 & u_CSAwallace_cska32_and_14_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_13_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa39_and1 = u_CSAwallace_cska32_csa8_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_13_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa39_or0 = u_CSAwallace_cska32_csa8_csa_component_fa39_and0 | u_CSAwallace_cska32_csa8_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa40_xor0 = u_CSAwallace_cska32_and_16_24 ^ u_CSAwallace_cska32_and_15_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa40_and0 = u_CSAwallace_cska32_and_16_24 & u_CSAwallace_cska32_and_15_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_14_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa40_and1 = u_CSAwallace_cska32_csa8_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_14_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa40_or0 = u_CSAwallace_cska32_csa8_csa_component_fa40_and0 | u_CSAwallace_cska32_csa8_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa41_xor0 = u_CSAwallace_cska32_and_17_24 ^ u_CSAwallace_cska32_and_16_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa41_and0 = u_CSAwallace_cska32_and_17_24 & u_CSAwallace_cska32_and_16_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_and_15_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa41_and1 = u_CSAwallace_cska32_csa8_csa_component_fa41_xor0 & u_CSAwallace_cska32_and_15_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa41_or0 = u_CSAwallace_cska32_csa8_csa_component_fa41_and0 | u_CSAwallace_cska32_csa8_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa42_xor0 = u_CSAwallace_cska32_and_18_24 ^ u_CSAwallace_cska32_and_17_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa42_and0 = u_CSAwallace_cska32_and_18_24 & u_CSAwallace_cska32_and_17_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_and_16_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa42_and1 = u_CSAwallace_cska32_csa8_csa_component_fa42_xor0 & u_CSAwallace_cska32_and_16_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa42_or0 = u_CSAwallace_cska32_csa8_csa_component_fa42_and0 | u_CSAwallace_cska32_csa8_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa43_xor0 = u_CSAwallace_cska32_and_19_24 ^ u_CSAwallace_cska32_and_18_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa43_and0 = u_CSAwallace_cska32_and_19_24 & u_CSAwallace_cska32_and_18_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_and_17_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa43_and1 = u_CSAwallace_cska32_csa8_csa_component_fa43_xor0 & u_CSAwallace_cska32_and_17_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa43_or0 = u_CSAwallace_cska32_csa8_csa_component_fa43_and0 | u_CSAwallace_cska32_csa8_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa44_xor0 = u_CSAwallace_cska32_and_20_24 ^ u_CSAwallace_cska32_and_19_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa44_and0 = u_CSAwallace_cska32_and_20_24 & u_CSAwallace_cska32_and_19_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_and_18_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa44_and1 = u_CSAwallace_cska32_csa8_csa_component_fa44_xor0 & u_CSAwallace_cska32_and_18_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa44_or0 = u_CSAwallace_cska32_csa8_csa_component_fa44_and0 | u_CSAwallace_cska32_csa8_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa45_xor0 = u_CSAwallace_cska32_and_21_24 ^ u_CSAwallace_cska32_and_20_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa45_and0 = u_CSAwallace_cska32_and_21_24 & u_CSAwallace_cska32_and_20_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_and_19_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa45_and1 = u_CSAwallace_cska32_csa8_csa_component_fa45_xor0 & u_CSAwallace_cska32_and_19_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa45_or0 = u_CSAwallace_cska32_csa8_csa_component_fa45_and0 | u_CSAwallace_cska32_csa8_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa46_xor0 = u_CSAwallace_cska32_and_22_24 ^ u_CSAwallace_cska32_and_21_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa46_and0 = u_CSAwallace_cska32_and_22_24 & u_CSAwallace_cska32_and_21_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_and_20_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa46_and1 = u_CSAwallace_cska32_csa8_csa_component_fa46_xor0 & u_CSAwallace_cska32_and_20_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa46_or0 = u_CSAwallace_cska32_csa8_csa_component_fa46_and0 | u_CSAwallace_cska32_csa8_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa47_xor0 = u_CSAwallace_cska32_and_23_24 ^ u_CSAwallace_cska32_and_22_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa47_and0 = u_CSAwallace_cska32_and_23_24 & u_CSAwallace_cska32_and_22_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_and_21_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa47_and1 = u_CSAwallace_cska32_csa8_csa_component_fa47_xor0 & u_CSAwallace_cska32_and_21_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa47_or0 = u_CSAwallace_cska32_csa8_csa_component_fa47_and0 | u_CSAwallace_cska32_csa8_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa48_xor0 = u_CSAwallace_cska32_and_24_24 ^ u_CSAwallace_cska32_and_23_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa48_and0 = u_CSAwallace_cska32_and_24_24 & u_CSAwallace_cska32_and_23_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_and_22_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa48_and1 = u_CSAwallace_cska32_csa8_csa_component_fa48_xor0 & u_CSAwallace_cska32_and_22_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa48_or0 = u_CSAwallace_cska32_csa8_csa_component_fa48_and0 | u_CSAwallace_cska32_csa8_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa49_xor0 = u_CSAwallace_cska32_and_25_24 ^ u_CSAwallace_cska32_and_24_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa49_and0 = u_CSAwallace_cska32_and_25_24 & u_CSAwallace_cska32_and_24_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_and_23_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa49_and1 = u_CSAwallace_cska32_csa8_csa_component_fa49_xor0 & u_CSAwallace_cska32_and_23_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa49_or0 = u_CSAwallace_cska32_csa8_csa_component_fa49_and0 | u_CSAwallace_cska32_csa8_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa50_xor0 = u_CSAwallace_cska32_and_26_24 ^ u_CSAwallace_cska32_and_25_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa50_and0 = u_CSAwallace_cska32_and_26_24 & u_CSAwallace_cska32_and_25_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_and_24_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa50_and1 = u_CSAwallace_cska32_csa8_csa_component_fa50_xor0 & u_CSAwallace_cska32_and_24_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa50_or0 = u_CSAwallace_cska32_csa8_csa_component_fa50_and0 | u_CSAwallace_cska32_csa8_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa51_xor0 = u_CSAwallace_cska32_and_27_24 ^ u_CSAwallace_cska32_and_26_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa51_and0 = u_CSAwallace_cska32_and_27_24 & u_CSAwallace_cska32_and_26_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_and_25_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa51_and1 = u_CSAwallace_cska32_csa8_csa_component_fa51_xor0 & u_CSAwallace_cska32_and_25_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa51_or0 = u_CSAwallace_cska32_csa8_csa_component_fa51_and0 | u_CSAwallace_cska32_csa8_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa52_xor0 = u_CSAwallace_cska32_and_28_24 ^ u_CSAwallace_cska32_and_27_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa52_and0 = u_CSAwallace_cska32_and_28_24 & u_CSAwallace_cska32_and_27_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_and_26_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa52_and1 = u_CSAwallace_cska32_csa8_csa_component_fa52_xor0 & u_CSAwallace_cska32_and_26_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa52_or0 = u_CSAwallace_cska32_csa8_csa_component_fa52_and0 | u_CSAwallace_cska32_csa8_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa53_xor0 = u_CSAwallace_cska32_and_29_24 ^ u_CSAwallace_cska32_and_28_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa53_and0 = u_CSAwallace_cska32_and_29_24 & u_CSAwallace_cska32_and_28_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa53_xor0 ^ u_CSAwallace_cska32_and_27_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa53_and1 = u_CSAwallace_cska32_csa8_csa_component_fa53_xor0 & u_CSAwallace_cska32_and_27_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa53_or0 = u_CSAwallace_cska32_csa8_csa_component_fa53_and0 | u_CSAwallace_cska32_csa8_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa54_xor0 = u_CSAwallace_cska32_and_30_24 ^ u_CSAwallace_cska32_and_29_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa54_and0 = u_CSAwallace_cska32_and_30_24 & u_CSAwallace_cska32_and_29_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa54_xor0 ^ u_CSAwallace_cska32_and_28_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa54_and1 = u_CSAwallace_cska32_csa8_csa_component_fa54_xor0 & u_CSAwallace_cska32_and_28_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa54_or0 = u_CSAwallace_cska32_csa8_csa_component_fa54_and0 | u_CSAwallace_cska32_csa8_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa55_xor0 = u_CSAwallace_cska32_and_31_24 ^ u_CSAwallace_cska32_and_30_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa55_and0 = u_CSAwallace_cska32_and_31_24 & u_CSAwallace_cska32_and_30_25;
  assign u_CSAwallace_cska32_csa8_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa55_xor0 ^ u_CSAwallace_cska32_and_29_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa55_and1 = u_CSAwallace_cska32_csa8_csa_component_fa55_xor0 & u_CSAwallace_cska32_and_29_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa55_or0 = u_CSAwallace_cska32_csa8_csa_component_fa55_and0 | u_CSAwallace_cska32_csa8_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa8_csa_component_fa56_xor1 = u_CSAwallace_cska32_and_31_25 ^ u_CSAwallace_cska32_and_30_26;
  assign u_CSAwallace_cska32_csa8_csa_component_fa56_and1 = u_CSAwallace_cska32_and_31_25 & u_CSAwallace_cska32_and_30_26;
  assign u_CSAwallace_cska32_csa9_csa_component_fa28_xor0 = u_CSAwallace_cska32_and_1_27 ^ u_CSAwallace_cska32_and_0_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa28_and0 = u_CSAwallace_cska32_and_1_27 & u_CSAwallace_cska32_and_0_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa29_xor0 = u_CSAwallace_cska32_and_2_27 ^ u_CSAwallace_cska32_and_1_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa29_and0 = u_CSAwallace_cska32_and_2_27 & u_CSAwallace_cska32_and_1_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_and_0_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa29_and1 = u_CSAwallace_cska32_csa9_csa_component_fa29_xor0 & u_CSAwallace_cska32_and_0_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa29_or0 = u_CSAwallace_cska32_csa9_csa_component_fa29_and0 | u_CSAwallace_cska32_csa9_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa30_xor0 = u_CSAwallace_cska32_and_3_27 ^ u_CSAwallace_cska32_and_2_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa30_and0 = u_CSAwallace_cska32_and_3_27 & u_CSAwallace_cska32_and_2_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_1_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa30_and1 = u_CSAwallace_cska32_csa9_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_1_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa30_or0 = u_CSAwallace_cska32_csa9_csa_component_fa30_and0 | u_CSAwallace_cska32_csa9_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa31_xor0 = u_CSAwallace_cska32_and_4_27 ^ u_CSAwallace_cska32_and_3_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa31_and0 = u_CSAwallace_cska32_and_4_27 & u_CSAwallace_cska32_and_3_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_2_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa31_and1 = u_CSAwallace_cska32_csa9_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_2_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa31_or0 = u_CSAwallace_cska32_csa9_csa_component_fa31_and0 | u_CSAwallace_cska32_csa9_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa32_xor0 = u_CSAwallace_cska32_and_5_27 ^ u_CSAwallace_cska32_and_4_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa32_and0 = u_CSAwallace_cska32_and_5_27 & u_CSAwallace_cska32_and_4_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_3_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa32_and1 = u_CSAwallace_cska32_csa9_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_3_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa32_or0 = u_CSAwallace_cska32_csa9_csa_component_fa32_and0 | u_CSAwallace_cska32_csa9_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_6_27 ^ u_CSAwallace_cska32_and_5_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa33_and0 = u_CSAwallace_cska32_and_6_27 & u_CSAwallace_cska32_and_5_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_4_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa33_and1 = u_CSAwallace_cska32_csa9_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_4_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa33_or0 = u_CSAwallace_cska32_csa9_csa_component_fa33_and0 | u_CSAwallace_cska32_csa9_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa34_xor0 = u_CSAwallace_cska32_and_7_27 ^ u_CSAwallace_cska32_and_6_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa34_and0 = u_CSAwallace_cska32_and_7_27 & u_CSAwallace_cska32_and_6_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_5_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa34_and1 = u_CSAwallace_cska32_csa9_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_5_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa34_or0 = u_CSAwallace_cska32_csa9_csa_component_fa34_and0 | u_CSAwallace_cska32_csa9_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa35_xor0 = u_CSAwallace_cska32_and_8_27 ^ u_CSAwallace_cska32_and_7_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa35_and0 = u_CSAwallace_cska32_and_8_27 & u_CSAwallace_cska32_and_7_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_6_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa35_and1 = u_CSAwallace_cska32_csa9_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_6_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa35_or0 = u_CSAwallace_cska32_csa9_csa_component_fa35_and0 | u_CSAwallace_cska32_csa9_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa36_xor0 = u_CSAwallace_cska32_and_9_27 ^ u_CSAwallace_cska32_and_8_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa36_and0 = u_CSAwallace_cska32_and_9_27 & u_CSAwallace_cska32_and_8_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_7_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa36_and1 = u_CSAwallace_cska32_csa9_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_7_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa36_or0 = u_CSAwallace_cska32_csa9_csa_component_fa36_and0 | u_CSAwallace_cska32_csa9_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa37_xor0 = u_CSAwallace_cska32_and_10_27 ^ u_CSAwallace_cska32_and_9_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa37_and0 = u_CSAwallace_cska32_and_10_27 & u_CSAwallace_cska32_and_9_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_8_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa37_and1 = u_CSAwallace_cska32_csa9_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_8_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa37_or0 = u_CSAwallace_cska32_csa9_csa_component_fa37_and0 | u_CSAwallace_cska32_csa9_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa38_xor0 = u_CSAwallace_cska32_and_11_27 ^ u_CSAwallace_cska32_and_10_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa38_and0 = u_CSAwallace_cska32_and_11_27 & u_CSAwallace_cska32_and_10_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_9_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa38_and1 = u_CSAwallace_cska32_csa9_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_9_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa38_or0 = u_CSAwallace_cska32_csa9_csa_component_fa38_and0 | u_CSAwallace_cska32_csa9_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa39_xor0 = u_CSAwallace_cska32_and_12_27 ^ u_CSAwallace_cska32_and_11_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa39_and0 = u_CSAwallace_cska32_and_12_27 & u_CSAwallace_cska32_and_11_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_10_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa39_and1 = u_CSAwallace_cska32_csa9_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_10_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa39_or0 = u_CSAwallace_cska32_csa9_csa_component_fa39_and0 | u_CSAwallace_cska32_csa9_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa40_xor0 = u_CSAwallace_cska32_and_13_27 ^ u_CSAwallace_cska32_and_12_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa40_and0 = u_CSAwallace_cska32_and_13_27 & u_CSAwallace_cska32_and_12_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_11_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa40_and1 = u_CSAwallace_cska32_csa9_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_11_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa40_or0 = u_CSAwallace_cska32_csa9_csa_component_fa40_and0 | u_CSAwallace_cska32_csa9_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa41_xor0 = u_CSAwallace_cska32_and_14_27 ^ u_CSAwallace_cska32_and_13_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa41_and0 = u_CSAwallace_cska32_and_14_27 & u_CSAwallace_cska32_and_13_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_and_12_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa41_and1 = u_CSAwallace_cska32_csa9_csa_component_fa41_xor0 & u_CSAwallace_cska32_and_12_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa41_or0 = u_CSAwallace_cska32_csa9_csa_component_fa41_and0 | u_CSAwallace_cska32_csa9_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa42_xor0 = u_CSAwallace_cska32_and_15_27 ^ u_CSAwallace_cska32_and_14_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa42_and0 = u_CSAwallace_cska32_and_15_27 & u_CSAwallace_cska32_and_14_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_and_13_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa42_and1 = u_CSAwallace_cska32_csa9_csa_component_fa42_xor0 & u_CSAwallace_cska32_and_13_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa42_or0 = u_CSAwallace_cska32_csa9_csa_component_fa42_and0 | u_CSAwallace_cska32_csa9_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa43_xor0 = u_CSAwallace_cska32_and_16_27 ^ u_CSAwallace_cska32_and_15_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa43_and0 = u_CSAwallace_cska32_and_16_27 & u_CSAwallace_cska32_and_15_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_and_14_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa43_and1 = u_CSAwallace_cska32_csa9_csa_component_fa43_xor0 & u_CSAwallace_cska32_and_14_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa43_or0 = u_CSAwallace_cska32_csa9_csa_component_fa43_and0 | u_CSAwallace_cska32_csa9_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa44_xor0 = u_CSAwallace_cska32_and_17_27 ^ u_CSAwallace_cska32_and_16_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa44_and0 = u_CSAwallace_cska32_and_17_27 & u_CSAwallace_cska32_and_16_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_and_15_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa44_and1 = u_CSAwallace_cska32_csa9_csa_component_fa44_xor0 & u_CSAwallace_cska32_and_15_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa44_or0 = u_CSAwallace_cska32_csa9_csa_component_fa44_and0 | u_CSAwallace_cska32_csa9_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa45_xor0 = u_CSAwallace_cska32_and_18_27 ^ u_CSAwallace_cska32_and_17_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa45_and0 = u_CSAwallace_cska32_and_18_27 & u_CSAwallace_cska32_and_17_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_and_16_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa45_and1 = u_CSAwallace_cska32_csa9_csa_component_fa45_xor0 & u_CSAwallace_cska32_and_16_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa45_or0 = u_CSAwallace_cska32_csa9_csa_component_fa45_and0 | u_CSAwallace_cska32_csa9_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa46_xor0 = u_CSAwallace_cska32_and_19_27 ^ u_CSAwallace_cska32_and_18_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa46_and0 = u_CSAwallace_cska32_and_19_27 & u_CSAwallace_cska32_and_18_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_and_17_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa46_and1 = u_CSAwallace_cska32_csa9_csa_component_fa46_xor0 & u_CSAwallace_cska32_and_17_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa46_or0 = u_CSAwallace_cska32_csa9_csa_component_fa46_and0 | u_CSAwallace_cska32_csa9_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa47_xor0 = u_CSAwallace_cska32_and_20_27 ^ u_CSAwallace_cska32_and_19_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa47_and0 = u_CSAwallace_cska32_and_20_27 & u_CSAwallace_cska32_and_19_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_and_18_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa47_and1 = u_CSAwallace_cska32_csa9_csa_component_fa47_xor0 & u_CSAwallace_cska32_and_18_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa47_or0 = u_CSAwallace_cska32_csa9_csa_component_fa47_and0 | u_CSAwallace_cska32_csa9_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa48_xor0 = u_CSAwallace_cska32_and_21_27 ^ u_CSAwallace_cska32_and_20_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa48_and0 = u_CSAwallace_cska32_and_21_27 & u_CSAwallace_cska32_and_20_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_and_19_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa48_and1 = u_CSAwallace_cska32_csa9_csa_component_fa48_xor0 & u_CSAwallace_cska32_and_19_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa48_or0 = u_CSAwallace_cska32_csa9_csa_component_fa48_and0 | u_CSAwallace_cska32_csa9_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa49_xor0 = u_CSAwallace_cska32_and_22_27 ^ u_CSAwallace_cska32_and_21_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa49_and0 = u_CSAwallace_cska32_and_22_27 & u_CSAwallace_cska32_and_21_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_and_20_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa49_and1 = u_CSAwallace_cska32_csa9_csa_component_fa49_xor0 & u_CSAwallace_cska32_and_20_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa49_or0 = u_CSAwallace_cska32_csa9_csa_component_fa49_and0 | u_CSAwallace_cska32_csa9_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa50_xor0 = u_CSAwallace_cska32_and_23_27 ^ u_CSAwallace_cska32_and_22_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa50_and0 = u_CSAwallace_cska32_and_23_27 & u_CSAwallace_cska32_and_22_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_and_21_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa50_and1 = u_CSAwallace_cska32_csa9_csa_component_fa50_xor0 & u_CSAwallace_cska32_and_21_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa50_or0 = u_CSAwallace_cska32_csa9_csa_component_fa50_and0 | u_CSAwallace_cska32_csa9_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa51_xor0 = u_CSAwallace_cska32_and_24_27 ^ u_CSAwallace_cska32_and_23_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa51_and0 = u_CSAwallace_cska32_and_24_27 & u_CSAwallace_cska32_and_23_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_and_22_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa51_and1 = u_CSAwallace_cska32_csa9_csa_component_fa51_xor0 & u_CSAwallace_cska32_and_22_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa51_or0 = u_CSAwallace_cska32_csa9_csa_component_fa51_and0 | u_CSAwallace_cska32_csa9_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa52_xor0 = u_CSAwallace_cska32_and_25_27 ^ u_CSAwallace_cska32_and_24_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa52_and0 = u_CSAwallace_cska32_and_25_27 & u_CSAwallace_cska32_and_24_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_and_23_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa52_and1 = u_CSAwallace_cska32_csa9_csa_component_fa52_xor0 & u_CSAwallace_cska32_and_23_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa52_or0 = u_CSAwallace_cska32_csa9_csa_component_fa52_and0 | u_CSAwallace_cska32_csa9_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa53_xor0 = u_CSAwallace_cska32_and_26_27 ^ u_CSAwallace_cska32_and_25_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa53_and0 = u_CSAwallace_cska32_and_26_27 & u_CSAwallace_cska32_and_25_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa53_xor0 ^ u_CSAwallace_cska32_and_24_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa53_and1 = u_CSAwallace_cska32_csa9_csa_component_fa53_xor0 & u_CSAwallace_cska32_and_24_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa53_or0 = u_CSAwallace_cska32_csa9_csa_component_fa53_and0 | u_CSAwallace_cska32_csa9_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa54_xor0 = u_CSAwallace_cska32_and_27_27 ^ u_CSAwallace_cska32_and_26_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa54_and0 = u_CSAwallace_cska32_and_27_27 & u_CSAwallace_cska32_and_26_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa54_xor0 ^ u_CSAwallace_cska32_and_25_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa54_and1 = u_CSAwallace_cska32_csa9_csa_component_fa54_xor0 & u_CSAwallace_cska32_and_25_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa54_or0 = u_CSAwallace_cska32_csa9_csa_component_fa54_and0 | u_CSAwallace_cska32_csa9_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa55_xor0 = u_CSAwallace_cska32_and_28_27 ^ u_CSAwallace_cska32_and_27_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa55_and0 = u_CSAwallace_cska32_and_28_27 & u_CSAwallace_cska32_and_27_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa55_xor0 ^ u_CSAwallace_cska32_and_26_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa55_and1 = u_CSAwallace_cska32_csa9_csa_component_fa55_xor0 & u_CSAwallace_cska32_and_26_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa55_or0 = u_CSAwallace_cska32_csa9_csa_component_fa55_and0 | u_CSAwallace_cska32_csa9_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa56_xor0 = u_CSAwallace_cska32_and_29_27 ^ u_CSAwallace_cska32_and_28_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa56_and0 = u_CSAwallace_cska32_and_29_27 & u_CSAwallace_cska32_and_28_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa56_xor0 ^ u_CSAwallace_cska32_and_27_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa56_and1 = u_CSAwallace_cska32_csa9_csa_component_fa56_xor0 & u_CSAwallace_cska32_and_27_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa56_or0 = u_CSAwallace_cska32_csa9_csa_component_fa56_and0 | u_CSAwallace_cska32_csa9_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa57_xor0 = u_CSAwallace_cska32_and_30_27 ^ u_CSAwallace_cska32_and_29_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa57_and0 = u_CSAwallace_cska32_and_30_27 & u_CSAwallace_cska32_and_29_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa57_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa57_xor0 ^ u_CSAwallace_cska32_and_28_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa57_and1 = u_CSAwallace_cska32_csa9_csa_component_fa57_xor0 & u_CSAwallace_cska32_and_28_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa57_or0 = u_CSAwallace_cska32_csa9_csa_component_fa57_and0 | u_CSAwallace_cska32_csa9_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa58_xor0 = u_CSAwallace_cska32_and_31_27 ^ u_CSAwallace_cska32_and_30_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa58_and0 = u_CSAwallace_cska32_and_31_27 & u_CSAwallace_cska32_and_30_28;
  assign u_CSAwallace_cska32_csa9_csa_component_fa58_xor1 = u_CSAwallace_cska32_csa9_csa_component_fa58_xor0 ^ u_CSAwallace_cska32_and_29_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa58_and1 = u_CSAwallace_cska32_csa9_csa_component_fa58_xor0 & u_CSAwallace_cska32_and_29_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa58_or0 = u_CSAwallace_cska32_csa9_csa_component_fa58_and0 | u_CSAwallace_cska32_csa9_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa9_csa_component_fa59_xor1 = u_CSAwallace_cska32_and_31_28 ^ u_CSAwallace_cska32_and_30_29;
  assign u_CSAwallace_cska32_csa9_csa_component_fa59_and1 = u_CSAwallace_cska32_and_31_28 & u_CSAwallace_cska32_and_30_29;
  assign u_CSAwallace_cska32_csa10_csa_component_fa2_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa2_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa2_and0 = u_CSAwallace_cska32_csa0_csa_component_fa2_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa3_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa3_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa3_and0 = u_CSAwallace_cska32_csa0_csa_component_fa3_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa3_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa3_xor0 ^ u_CSAwallace_cska32_and_0_3;
  assign u_CSAwallace_cska32_csa10_csa_component_fa3_and1 = u_CSAwallace_cska32_csa10_csa_component_fa3_xor0 & u_CSAwallace_cska32_and_0_3;
  assign u_CSAwallace_cska32_csa10_csa_component_fa3_or0 = u_CSAwallace_cska32_csa10_csa_component_fa3_and0 | u_CSAwallace_cska32_csa10_csa_component_fa3_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa4_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa4_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa4_and0 = u_CSAwallace_cska32_csa0_csa_component_fa4_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa4_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa4_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa4_xor0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa4_and1 = u_CSAwallace_cska32_csa10_csa_component_fa4_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa4_xor0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa4_or0 = u_CSAwallace_cska32_csa10_csa_component_fa4_and0 | u_CSAwallace_cska32_csa10_csa_component_fa4_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa5_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa5_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa4_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa5_and0 = u_CSAwallace_cska32_csa0_csa_component_fa5_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa4_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa5_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa5_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa5_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa5_and1 = u_CSAwallace_cska32_csa10_csa_component_fa5_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa5_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa5_or0 = u_CSAwallace_cska32_csa10_csa_component_fa5_and0 | u_CSAwallace_cska32_csa10_csa_component_fa5_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa6_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa6_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa5_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa6_and0 = u_CSAwallace_cska32_csa0_csa_component_fa6_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa5_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa6_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa6_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa6_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa6_and1 = u_CSAwallace_cska32_csa10_csa_component_fa6_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa6_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa6_or0 = u_CSAwallace_cska32_csa10_csa_component_fa6_and0 | u_CSAwallace_cska32_csa10_csa_component_fa6_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa7_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa7_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa6_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa7_and0 = u_CSAwallace_cska32_csa0_csa_component_fa7_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa6_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa7_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa7_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa7_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa7_and1 = u_CSAwallace_cska32_csa10_csa_component_fa7_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa7_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa7_or0 = u_CSAwallace_cska32_csa10_csa_component_fa7_and0 | u_CSAwallace_cska32_csa10_csa_component_fa7_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa8_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa8_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa7_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa8_and0 = u_CSAwallace_cska32_csa0_csa_component_fa8_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa7_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa8_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa8_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa8_and1 = u_CSAwallace_cska32_csa10_csa_component_fa8_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa8_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa8_or0 = u_CSAwallace_cska32_csa10_csa_component_fa8_and0 | u_CSAwallace_cska32_csa10_csa_component_fa8_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa9_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa9_and0 = u_CSAwallace_cska32_csa0_csa_component_fa9_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa9_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa9_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa9_and1 = u_CSAwallace_cska32_csa10_csa_component_fa9_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa9_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa9_or0 = u_CSAwallace_cska32_csa10_csa_component_fa9_and0 | u_CSAwallace_cska32_csa10_csa_component_fa9_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa10_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa10_and0 = u_CSAwallace_cska32_csa0_csa_component_fa10_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa10_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa10_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa10_and1 = u_CSAwallace_cska32_csa10_csa_component_fa10_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa10_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa10_or0 = u_CSAwallace_cska32_csa10_csa_component_fa10_and0 | u_CSAwallace_cska32_csa10_csa_component_fa10_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa11_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa11_and0 = u_CSAwallace_cska32_csa0_csa_component_fa11_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa11_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa11_and1 = u_CSAwallace_cska32_csa10_csa_component_fa11_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa11_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa11_or0 = u_CSAwallace_cska32_csa10_csa_component_fa11_and0 | u_CSAwallace_cska32_csa10_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa12_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa12_and0 = u_CSAwallace_cska32_csa0_csa_component_fa12_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa12_and1 = u_CSAwallace_cska32_csa10_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa12_or0 = u_CSAwallace_cska32_csa10_csa_component_fa12_and0 | u_CSAwallace_cska32_csa10_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa13_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa13_and0 = u_CSAwallace_cska32_csa0_csa_component_fa13_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa13_and1 = u_CSAwallace_cska32_csa10_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa13_or0 = u_CSAwallace_cska32_csa10_csa_component_fa13_and0 | u_CSAwallace_cska32_csa10_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa14_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa14_and0 = u_CSAwallace_cska32_csa0_csa_component_fa14_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa14_and1 = u_CSAwallace_cska32_csa10_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa14_or0 = u_CSAwallace_cska32_csa10_csa_component_fa14_and0 | u_CSAwallace_cska32_csa10_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa15_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa15_and0 = u_CSAwallace_cska32_csa0_csa_component_fa15_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa15_and1 = u_CSAwallace_cska32_csa10_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa15_or0 = u_CSAwallace_cska32_csa10_csa_component_fa15_and0 | u_CSAwallace_cska32_csa10_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa16_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa16_and0 = u_CSAwallace_cska32_csa0_csa_component_fa16_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa16_and1 = u_CSAwallace_cska32_csa10_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa16_or0 = u_CSAwallace_cska32_csa10_csa_component_fa16_and0 | u_CSAwallace_cska32_csa10_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa17_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa17_and0 = u_CSAwallace_cska32_csa0_csa_component_fa17_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa17_and1 = u_CSAwallace_cska32_csa10_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa17_or0 = u_CSAwallace_cska32_csa10_csa_component_fa17_and0 | u_CSAwallace_cska32_csa10_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa18_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa18_and0 = u_CSAwallace_cska32_csa0_csa_component_fa18_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa18_and1 = u_CSAwallace_cska32_csa10_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa18_or0 = u_CSAwallace_cska32_csa10_csa_component_fa18_and0 | u_CSAwallace_cska32_csa10_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa19_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa19_and0 = u_CSAwallace_cska32_csa0_csa_component_fa19_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa19_and1 = u_CSAwallace_cska32_csa10_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa19_or0 = u_CSAwallace_cska32_csa10_csa_component_fa19_and0 | u_CSAwallace_cska32_csa10_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa20_and0 = u_CSAwallace_cska32_csa0_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa20_and1 = u_CSAwallace_cska32_csa10_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa20_or0 = u_CSAwallace_cska32_csa10_csa_component_fa20_and0 | u_CSAwallace_cska32_csa10_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa21_and0 = u_CSAwallace_cska32_csa0_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa21_and1 = u_CSAwallace_cska32_csa10_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa21_or0 = u_CSAwallace_cska32_csa10_csa_component_fa21_and0 | u_CSAwallace_cska32_csa10_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa22_and0 = u_CSAwallace_cska32_csa0_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa22_and1 = u_CSAwallace_cska32_csa10_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa22_or0 = u_CSAwallace_cska32_csa10_csa_component_fa22_and0 | u_CSAwallace_cska32_csa10_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa23_and0 = u_CSAwallace_cska32_csa0_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa23_and1 = u_CSAwallace_cska32_csa10_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa23_or0 = u_CSAwallace_cska32_csa10_csa_component_fa23_and0 | u_CSAwallace_cska32_csa10_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa24_and0 = u_CSAwallace_cska32_csa0_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa24_and1 = u_CSAwallace_cska32_csa10_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa24_or0 = u_CSAwallace_cska32_csa10_csa_component_fa24_and0 | u_CSAwallace_cska32_csa10_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa25_and0 = u_CSAwallace_cska32_csa0_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa25_and1 = u_CSAwallace_cska32_csa10_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa25_or0 = u_CSAwallace_cska32_csa10_csa_component_fa25_and0 | u_CSAwallace_cska32_csa10_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa26_and0 = u_CSAwallace_cska32_csa0_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa26_and1 = u_CSAwallace_cska32_csa10_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa26_or0 = u_CSAwallace_cska32_csa10_csa_component_fa26_and0 | u_CSAwallace_cska32_csa10_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa27_and0 = u_CSAwallace_cska32_csa0_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa27_and1 = u_CSAwallace_cska32_csa10_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa27_or0 = u_CSAwallace_cska32_csa10_csa_component_fa27_and0 | u_CSAwallace_cska32_csa10_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa28_and0 = u_CSAwallace_cska32_csa0_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa28_and1 = u_CSAwallace_cska32_csa10_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa28_or0 = u_CSAwallace_cska32_csa10_csa_component_fa28_and0 | u_CSAwallace_cska32_csa10_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa29_and0 = u_CSAwallace_cska32_csa0_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa29_and1 = u_CSAwallace_cska32_csa10_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa29_or0 = u_CSAwallace_cska32_csa10_csa_component_fa29_and0 | u_CSAwallace_cska32_csa10_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa30_and0 = u_CSAwallace_cska32_csa0_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa30_and1 = u_CSAwallace_cska32_csa10_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa30_or0 = u_CSAwallace_cska32_csa10_csa_component_fa30_and0 | u_CSAwallace_cska32_csa10_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa31_and0 = u_CSAwallace_cska32_csa0_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa31_and1 = u_CSAwallace_cska32_csa10_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa31_or0 = u_CSAwallace_cska32_csa10_csa_component_fa31_and0 | u_CSAwallace_cska32_csa10_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa0_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa0_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa32_and0 = u_CSAwallace_cska32_csa0_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa0_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa10_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa32_and1 = u_CSAwallace_cska32_csa10_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa32_or0 = u_CSAwallace_cska32_csa10_csa_component_fa32_and0 | u_CSAwallace_cska32_csa10_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa33_xor0 = u_CSAwallace_cska32_and_31_2 ^ u_CSAwallace_cska32_csa0_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa33_and0 = u_CSAwallace_cska32_and_31_2 & u_CSAwallace_cska32_csa0_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa10_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa33_and1 = u_CSAwallace_cska32_csa10_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa10_csa_component_fa33_or0 = u_CSAwallace_cska32_csa10_csa_component_fa33_and0 | u_CSAwallace_cska32_csa10_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa6_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa5_or0 ^ u_CSAwallace_cska32_and_0_6;
  assign u_CSAwallace_cska32_csa11_csa_component_fa6_and0 = u_CSAwallace_cska32_csa1_csa_component_fa5_or0 & u_CSAwallace_cska32_and_0_6;
  assign u_CSAwallace_cska32_csa11_csa_component_fa7_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa6_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa7_xor0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa7_and0 = u_CSAwallace_cska32_csa1_csa_component_fa6_or0 & u_CSAwallace_cska32_csa2_csa_component_fa7_xor0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa8_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa7_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa8_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa8_and0 = u_CSAwallace_cska32_csa1_csa_component_fa7_or0 & u_CSAwallace_cska32_csa2_csa_component_fa8_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa8_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa8_and1 = u_CSAwallace_cska32_csa11_csa_component_fa8_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa8_or0 = u_CSAwallace_cska32_csa11_csa_component_fa8_and0 | u_CSAwallace_cska32_csa11_csa_component_fa8_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa8_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa9_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa9_and0 = u_CSAwallace_cska32_csa1_csa_component_fa8_or0 & u_CSAwallace_cska32_csa2_csa_component_fa9_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa9_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa9_and1 = u_CSAwallace_cska32_csa11_csa_component_fa9_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa9_or0 = u_CSAwallace_cska32_csa11_csa_component_fa9_and0 | u_CSAwallace_cska32_csa11_csa_component_fa9_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa9_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa10_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa10_and0 = u_CSAwallace_cska32_csa1_csa_component_fa9_or0 & u_CSAwallace_cska32_csa2_csa_component_fa10_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa10_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa10_and1 = u_CSAwallace_cska32_csa11_csa_component_fa10_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa10_or0 = u_CSAwallace_cska32_csa11_csa_component_fa10_and0 | u_CSAwallace_cska32_csa11_csa_component_fa10_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa10_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa11_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa11_and0 = u_CSAwallace_cska32_csa1_csa_component_fa10_or0 & u_CSAwallace_cska32_csa2_csa_component_fa11_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa11_and1 = u_CSAwallace_cska32_csa11_csa_component_fa11_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa11_or0 = u_CSAwallace_cska32_csa11_csa_component_fa11_and0 | u_CSAwallace_cska32_csa11_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa11_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa12_and0 = u_CSAwallace_cska32_csa1_csa_component_fa11_or0 & u_CSAwallace_cska32_csa2_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa12_and1 = u_CSAwallace_cska32_csa11_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa12_or0 = u_CSAwallace_cska32_csa11_csa_component_fa12_and0 | u_CSAwallace_cska32_csa11_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa12_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa13_and0 = u_CSAwallace_cska32_csa1_csa_component_fa12_or0 & u_CSAwallace_cska32_csa2_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa13_and1 = u_CSAwallace_cska32_csa11_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa13_or0 = u_CSAwallace_cska32_csa11_csa_component_fa13_and0 | u_CSAwallace_cska32_csa11_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa13_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa14_and0 = u_CSAwallace_cska32_csa1_csa_component_fa13_or0 & u_CSAwallace_cska32_csa2_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa14_and1 = u_CSAwallace_cska32_csa11_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa14_or0 = u_CSAwallace_cska32_csa11_csa_component_fa14_and0 | u_CSAwallace_cska32_csa11_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa14_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa15_and0 = u_CSAwallace_cska32_csa1_csa_component_fa14_or0 & u_CSAwallace_cska32_csa2_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa15_and1 = u_CSAwallace_cska32_csa11_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa15_or0 = u_CSAwallace_cska32_csa11_csa_component_fa15_and0 | u_CSAwallace_cska32_csa11_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa15_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa16_and0 = u_CSAwallace_cska32_csa1_csa_component_fa15_or0 & u_CSAwallace_cska32_csa2_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa16_and1 = u_CSAwallace_cska32_csa11_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa16_or0 = u_CSAwallace_cska32_csa11_csa_component_fa16_and0 | u_CSAwallace_cska32_csa11_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa16_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa17_and0 = u_CSAwallace_cska32_csa1_csa_component_fa16_or0 & u_CSAwallace_cska32_csa2_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa17_and1 = u_CSAwallace_cska32_csa11_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa17_or0 = u_CSAwallace_cska32_csa11_csa_component_fa17_and0 | u_CSAwallace_cska32_csa11_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa17_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa18_and0 = u_CSAwallace_cska32_csa1_csa_component_fa17_or0 & u_CSAwallace_cska32_csa2_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa18_and1 = u_CSAwallace_cska32_csa11_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa18_or0 = u_CSAwallace_cska32_csa11_csa_component_fa18_and0 | u_CSAwallace_cska32_csa11_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa18_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa19_and0 = u_CSAwallace_cska32_csa1_csa_component_fa18_or0 & u_CSAwallace_cska32_csa2_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa19_and1 = u_CSAwallace_cska32_csa11_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa19_or0 = u_CSAwallace_cska32_csa11_csa_component_fa19_and0 | u_CSAwallace_cska32_csa11_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa19_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa20_and0 = u_CSAwallace_cska32_csa1_csa_component_fa19_or0 & u_CSAwallace_cska32_csa2_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa20_and1 = u_CSAwallace_cska32_csa11_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa20_or0 = u_CSAwallace_cska32_csa11_csa_component_fa20_and0 | u_CSAwallace_cska32_csa11_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa20_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa21_and0 = u_CSAwallace_cska32_csa1_csa_component_fa20_or0 & u_CSAwallace_cska32_csa2_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa21_and1 = u_CSAwallace_cska32_csa11_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa21_or0 = u_CSAwallace_cska32_csa11_csa_component_fa21_and0 | u_CSAwallace_cska32_csa11_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa21_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa22_and0 = u_CSAwallace_cska32_csa1_csa_component_fa21_or0 & u_CSAwallace_cska32_csa2_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa22_and1 = u_CSAwallace_cska32_csa11_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa22_or0 = u_CSAwallace_cska32_csa11_csa_component_fa22_and0 | u_CSAwallace_cska32_csa11_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa22_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa23_and0 = u_CSAwallace_cska32_csa1_csa_component_fa22_or0 & u_CSAwallace_cska32_csa2_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa23_and1 = u_CSAwallace_cska32_csa11_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa23_or0 = u_CSAwallace_cska32_csa11_csa_component_fa23_and0 | u_CSAwallace_cska32_csa11_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa23_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa24_and0 = u_CSAwallace_cska32_csa1_csa_component_fa23_or0 & u_CSAwallace_cska32_csa2_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa24_and1 = u_CSAwallace_cska32_csa11_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa24_or0 = u_CSAwallace_cska32_csa11_csa_component_fa24_and0 | u_CSAwallace_cska32_csa11_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa24_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa25_and0 = u_CSAwallace_cska32_csa1_csa_component_fa24_or0 & u_CSAwallace_cska32_csa2_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa25_and1 = u_CSAwallace_cska32_csa11_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa25_or0 = u_CSAwallace_cska32_csa11_csa_component_fa25_and0 | u_CSAwallace_cska32_csa11_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa25_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa26_and0 = u_CSAwallace_cska32_csa1_csa_component_fa25_or0 & u_CSAwallace_cska32_csa2_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa26_and1 = u_CSAwallace_cska32_csa11_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa26_or0 = u_CSAwallace_cska32_csa11_csa_component_fa26_and0 | u_CSAwallace_cska32_csa11_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa26_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa27_and0 = u_CSAwallace_cska32_csa1_csa_component_fa26_or0 & u_CSAwallace_cska32_csa2_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa27_and1 = u_CSAwallace_cska32_csa11_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa27_or0 = u_CSAwallace_cska32_csa11_csa_component_fa27_and0 | u_CSAwallace_cska32_csa11_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa27_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa28_and0 = u_CSAwallace_cska32_csa1_csa_component_fa27_or0 & u_CSAwallace_cska32_csa2_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa28_and1 = u_CSAwallace_cska32_csa11_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa28_or0 = u_CSAwallace_cska32_csa11_csa_component_fa28_and0 | u_CSAwallace_cska32_csa11_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa28_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa29_and0 = u_CSAwallace_cska32_csa1_csa_component_fa28_or0 & u_CSAwallace_cska32_csa2_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa29_and1 = u_CSAwallace_cska32_csa11_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa29_or0 = u_CSAwallace_cska32_csa11_csa_component_fa29_and0 | u_CSAwallace_cska32_csa11_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa29_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa30_and0 = u_CSAwallace_cska32_csa1_csa_component_fa29_or0 & u_CSAwallace_cska32_csa2_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa30_and1 = u_CSAwallace_cska32_csa11_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa30_or0 = u_CSAwallace_cska32_csa11_csa_component_fa30_and0 | u_CSAwallace_cska32_csa11_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa30_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa31_and0 = u_CSAwallace_cska32_csa1_csa_component_fa30_or0 & u_CSAwallace_cska32_csa2_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa31_and1 = u_CSAwallace_cska32_csa11_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa31_or0 = u_CSAwallace_cska32_csa11_csa_component_fa31_and0 | u_CSAwallace_cska32_csa11_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa31_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa32_and0 = u_CSAwallace_cska32_csa1_csa_component_fa31_or0 & u_CSAwallace_cska32_csa2_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa32_and1 = u_CSAwallace_cska32_csa11_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa32_or0 = u_CSAwallace_cska32_csa11_csa_component_fa32_and0 | u_CSAwallace_cska32_csa11_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa32_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa33_and0 = u_CSAwallace_cska32_csa1_csa_component_fa32_or0 & u_CSAwallace_cska32_csa2_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa33_and1 = u_CSAwallace_cska32_csa11_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa33_or0 = u_CSAwallace_cska32_csa11_csa_component_fa33_and0 | u_CSAwallace_cska32_csa11_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa33_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa34_and0 = u_CSAwallace_cska32_csa1_csa_component_fa33_or0 & u_CSAwallace_cska32_csa2_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa34_and1 = u_CSAwallace_cska32_csa11_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa34_or0 = u_CSAwallace_cska32_csa11_csa_component_fa34_and0 | u_CSAwallace_cska32_csa11_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa34_or0 ^ u_CSAwallace_cska32_csa2_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa35_and0 = u_CSAwallace_cska32_csa1_csa_component_fa34_or0 & u_CSAwallace_cska32_csa2_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa35_and1 = u_CSAwallace_cska32_csa11_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa35_or0 = u_CSAwallace_cska32_csa11_csa_component_fa35_and0 | u_CSAwallace_cska32_csa11_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa35_and1 ^ u_CSAwallace_cska32_csa2_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa36_and0 = u_CSAwallace_cska32_csa1_csa_component_fa35_and1 & u_CSAwallace_cska32_csa2_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa2_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa36_and1 = u_CSAwallace_cska32_csa11_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa2_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa36_or0 = u_CSAwallace_cska32_csa11_csa_component_fa36_and0 | u_CSAwallace_cska32_csa11_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa2_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa37_and1 = u_CSAwallace_cska32_csa2_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa2_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa2_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa2_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa38_and1 = u_CSAwallace_cska32_csa2_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa2_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa11_csa_component_fa39_xor1 = u_CSAwallace_cska32_and_31_8 ^ u_CSAwallace_cska32_csa2_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa11_csa_component_fa39_and1 = u_CSAwallace_cska32_and_31_8 & u_CSAwallace_cska32_csa2_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa11_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa11_and0 = u_CSAwallace_cska32_csa3_csa_component_fa11_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa12_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa12_and0 = u_CSAwallace_cska32_csa3_csa_component_fa12_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_and_0_12;
  assign u_CSAwallace_cska32_csa12_csa_component_fa12_and1 = u_CSAwallace_cska32_csa12_csa_component_fa12_xor0 & u_CSAwallace_cska32_and_0_12;
  assign u_CSAwallace_cska32_csa12_csa_component_fa12_or0 = u_CSAwallace_cska32_csa12_csa_component_fa12_and0 | u_CSAwallace_cska32_csa12_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa13_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa13_and0 = u_CSAwallace_cska32_csa3_csa_component_fa13_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa13_xor0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa13_and1 = u_CSAwallace_cska32_csa12_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa13_xor0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa13_or0 = u_CSAwallace_cska32_csa12_csa_component_fa13_and0 | u_CSAwallace_cska32_csa12_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa14_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa14_and0 = u_CSAwallace_cska32_csa3_csa_component_fa14_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa14_and1 = u_CSAwallace_cska32_csa12_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa14_or0 = u_CSAwallace_cska32_csa12_csa_component_fa14_and0 | u_CSAwallace_cska32_csa12_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa15_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa15_and0 = u_CSAwallace_cska32_csa3_csa_component_fa15_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa15_and1 = u_CSAwallace_cska32_csa12_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa15_or0 = u_CSAwallace_cska32_csa12_csa_component_fa15_and0 | u_CSAwallace_cska32_csa12_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa16_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa16_and0 = u_CSAwallace_cska32_csa3_csa_component_fa16_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa16_and1 = u_CSAwallace_cska32_csa12_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa16_or0 = u_CSAwallace_cska32_csa12_csa_component_fa16_and0 | u_CSAwallace_cska32_csa12_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa17_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa17_and0 = u_CSAwallace_cska32_csa3_csa_component_fa17_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa17_and1 = u_CSAwallace_cska32_csa12_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa17_or0 = u_CSAwallace_cska32_csa12_csa_component_fa17_and0 | u_CSAwallace_cska32_csa12_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa18_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa18_and0 = u_CSAwallace_cska32_csa3_csa_component_fa18_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa18_and1 = u_CSAwallace_cska32_csa12_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa18_or0 = u_CSAwallace_cska32_csa12_csa_component_fa18_and0 | u_CSAwallace_cska32_csa12_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa19_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa19_and0 = u_CSAwallace_cska32_csa3_csa_component_fa19_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa19_and1 = u_CSAwallace_cska32_csa12_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa19_or0 = u_CSAwallace_cska32_csa12_csa_component_fa19_and0 | u_CSAwallace_cska32_csa12_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa20_and0 = u_CSAwallace_cska32_csa3_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa20_and1 = u_CSAwallace_cska32_csa12_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa20_or0 = u_CSAwallace_cska32_csa12_csa_component_fa20_and0 | u_CSAwallace_cska32_csa12_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa21_and0 = u_CSAwallace_cska32_csa3_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa21_and1 = u_CSAwallace_cska32_csa12_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa21_or0 = u_CSAwallace_cska32_csa12_csa_component_fa21_and0 | u_CSAwallace_cska32_csa12_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa22_and0 = u_CSAwallace_cska32_csa3_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa22_and1 = u_CSAwallace_cska32_csa12_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa22_or0 = u_CSAwallace_cska32_csa12_csa_component_fa22_and0 | u_CSAwallace_cska32_csa12_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa23_and0 = u_CSAwallace_cska32_csa3_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa23_and1 = u_CSAwallace_cska32_csa12_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa23_or0 = u_CSAwallace_cska32_csa12_csa_component_fa23_and0 | u_CSAwallace_cska32_csa12_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa24_and0 = u_CSAwallace_cska32_csa3_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa24_and1 = u_CSAwallace_cska32_csa12_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa24_or0 = u_CSAwallace_cska32_csa12_csa_component_fa24_and0 | u_CSAwallace_cska32_csa12_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa25_and0 = u_CSAwallace_cska32_csa3_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa25_and1 = u_CSAwallace_cska32_csa12_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa25_or0 = u_CSAwallace_cska32_csa12_csa_component_fa25_and0 | u_CSAwallace_cska32_csa12_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa26_and0 = u_CSAwallace_cska32_csa3_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa26_and1 = u_CSAwallace_cska32_csa12_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa26_or0 = u_CSAwallace_cska32_csa12_csa_component_fa26_and0 | u_CSAwallace_cska32_csa12_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa27_and0 = u_CSAwallace_cska32_csa3_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa27_and1 = u_CSAwallace_cska32_csa12_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa27_or0 = u_CSAwallace_cska32_csa12_csa_component_fa27_and0 | u_CSAwallace_cska32_csa12_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa28_and0 = u_CSAwallace_cska32_csa3_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa28_and1 = u_CSAwallace_cska32_csa12_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa28_or0 = u_CSAwallace_cska32_csa12_csa_component_fa28_and0 | u_CSAwallace_cska32_csa12_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa29_and0 = u_CSAwallace_cska32_csa3_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa29_and1 = u_CSAwallace_cska32_csa12_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa29_or0 = u_CSAwallace_cska32_csa12_csa_component_fa29_and0 | u_CSAwallace_cska32_csa12_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa30_and0 = u_CSAwallace_cska32_csa3_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa30_and1 = u_CSAwallace_cska32_csa12_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa30_or0 = u_CSAwallace_cska32_csa12_csa_component_fa30_and0 | u_CSAwallace_cska32_csa12_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa31_and0 = u_CSAwallace_cska32_csa3_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa31_and1 = u_CSAwallace_cska32_csa12_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa31_or0 = u_CSAwallace_cska32_csa12_csa_component_fa31_and0 | u_CSAwallace_cska32_csa12_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa32_and0 = u_CSAwallace_cska32_csa3_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa32_and1 = u_CSAwallace_cska32_csa12_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa32_or0 = u_CSAwallace_cska32_csa12_csa_component_fa32_and0 | u_CSAwallace_cska32_csa12_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa33_and0 = u_CSAwallace_cska32_csa3_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa33_and1 = u_CSAwallace_cska32_csa12_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa33_or0 = u_CSAwallace_cska32_csa12_csa_component_fa33_and0 | u_CSAwallace_cska32_csa12_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa34_and0 = u_CSAwallace_cska32_csa3_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa34_and1 = u_CSAwallace_cska32_csa12_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa34_or0 = u_CSAwallace_cska32_csa12_csa_component_fa34_and0 | u_CSAwallace_cska32_csa12_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa35_and0 = u_CSAwallace_cska32_csa3_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa35_and1 = u_CSAwallace_cska32_csa12_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa35_or0 = u_CSAwallace_cska32_csa12_csa_component_fa35_and0 | u_CSAwallace_cska32_csa12_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa36_and0 = u_CSAwallace_cska32_csa3_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa36_and1 = u_CSAwallace_cska32_csa12_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa36_or0 = u_CSAwallace_cska32_csa12_csa_component_fa36_and0 | u_CSAwallace_cska32_csa12_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa37_and0 = u_CSAwallace_cska32_csa3_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa37_and1 = u_CSAwallace_cska32_csa12_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa37_or0 = u_CSAwallace_cska32_csa12_csa_component_fa37_and0 | u_CSAwallace_cska32_csa12_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa38_and0 = u_CSAwallace_cska32_csa3_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa38_and1 = u_CSAwallace_cska32_csa12_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa38_or0 = u_CSAwallace_cska32_csa12_csa_component_fa38_and0 | u_CSAwallace_cska32_csa12_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa39_and0 = u_CSAwallace_cska32_csa3_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa39_and1 = u_CSAwallace_cska32_csa12_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa39_or0 = u_CSAwallace_cska32_csa12_csa_component_fa39_and0 | u_CSAwallace_cska32_csa12_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa40_and0 = u_CSAwallace_cska32_csa3_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa40_and1 = u_CSAwallace_cska32_csa12_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa40_or0 = u_CSAwallace_cska32_csa12_csa_component_fa40_and0 | u_CSAwallace_cska32_csa12_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa3_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa3_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa41_and0 = u_CSAwallace_cska32_csa3_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa3_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa12_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa41_and1 = u_CSAwallace_cska32_csa12_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa41_or0 = u_CSAwallace_cska32_csa12_csa_component_fa41_and0 | u_CSAwallace_cska32_csa12_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa42_xor0 = u_CSAwallace_cska32_and_31_11 ^ u_CSAwallace_cska32_csa3_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa42_and0 = u_CSAwallace_cska32_and_31_11 & u_CSAwallace_cska32_csa3_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa4_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa42_and1 = u_CSAwallace_cska32_csa12_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa4_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa12_csa_component_fa42_or0 = u_CSAwallace_cska32_csa12_csa_component_fa42_and0 | u_CSAwallace_cska32_csa12_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa14_or0 ^ u_CSAwallace_cska32_and_0_15;
  assign u_CSAwallace_cska32_csa13_csa_component_fa15_and0 = u_CSAwallace_cska32_csa4_csa_component_fa14_or0 & u_CSAwallace_cska32_and_0_15;
  assign u_CSAwallace_cska32_csa13_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa15_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa16_xor0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa16_and0 = u_CSAwallace_cska32_csa4_csa_component_fa15_or0 & u_CSAwallace_cska32_csa5_csa_component_fa16_xor0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa16_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa17_and0 = u_CSAwallace_cska32_csa4_csa_component_fa16_or0 & u_CSAwallace_cska32_csa5_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa17_and1 = u_CSAwallace_cska32_csa13_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa17_or0 = u_CSAwallace_cska32_csa13_csa_component_fa17_and0 | u_CSAwallace_cska32_csa13_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa17_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa18_and0 = u_CSAwallace_cska32_csa4_csa_component_fa17_or0 & u_CSAwallace_cska32_csa5_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa18_and1 = u_CSAwallace_cska32_csa13_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa18_or0 = u_CSAwallace_cska32_csa13_csa_component_fa18_and0 | u_CSAwallace_cska32_csa13_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa18_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa19_and0 = u_CSAwallace_cska32_csa4_csa_component_fa18_or0 & u_CSAwallace_cska32_csa5_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa19_and1 = u_CSAwallace_cska32_csa13_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa19_or0 = u_CSAwallace_cska32_csa13_csa_component_fa19_and0 | u_CSAwallace_cska32_csa13_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa19_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa20_and0 = u_CSAwallace_cska32_csa4_csa_component_fa19_or0 & u_CSAwallace_cska32_csa5_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa20_and1 = u_CSAwallace_cska32_csa13_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa20_or0 = u_CSAwallace_cska32_csa13_csa_component_fa20_and0 | u_CSAwallace_cska32_csa13_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa20_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa21_and0 = u_CSAwallace_cska32_csa4_csa_component_fa20_or0 & u_CSAwallace_cska32_csa5_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa21_and1 = u_CSAwallace_cska32_csa13_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa21_or0 = u_CSAwallace_cska32_csa13_csa_component_fa21_and0 | u_CSAwallace_cska32_csa13_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa21_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa22_and0 = u_CSAwallace_cska32_csa4_csa_component_fa21_or0 & u_CSAwallace_cska32_csa5_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa22_and1 = u_CSAwallace_cska32_csa13_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa22_or0 = u_CSAwallace_cska32_csa13_csa_component_fa22_and0 | u_CSAwallace_cska32_csa13_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa22_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa23_and0 = u_CSAwallace_cska32_csa4_csa_component_fa22_or0 & u_CSAwallace_cska32_csa5_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa23_and1 = u_CSAwallace_cska32_csa13_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa23_or0 = u_CSAwallace_cska32_csa13_csa_component_fa23_and0 | u_CSAwallace_cska32_csa13_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa23_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa24_and0 = u_CSAwallace_cska32_csa4_csa_component_fa23_or0 & u_CSAwallace_cska32_csa5_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa24_and1 = u_CSAwallace_cska32_csa13_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa24_or0 = u_CSAwallace_cska32_csa13_csa_component_fa24_and0 | u_CSAwallace_cska32_csa13_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa24_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa25_and0 = u_CSAwallace_cska32_csa4_csa_component_fa24_or0 & u_CSAwallace_cska32_csa5_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa25_and1 = u_CSAwallace_cska32_csa13_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa25_or0 = u_CSAwallace_cska32_csa13_csa_component_fa25_and0 | u_CSAwallace_cska32_csa13_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa25_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa26_and0 = u_CSAwallace_cska32_csa4_csa_component_fa25_or0 & u_CSAwallace_cska32_csa5_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa26_and1 = u_CSAwallace_cska32_csa13_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa26_or0 = u_CSAwallace_cska32_csa13_csa_component_fa26_and0 | u_CSAwallace_cska32_csa13_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa26_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa27_and0 = u_CSAwallace_cska32_csa4_csa_component_fa26_or0 & u_CSAwallace_cska32_csa5_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa27_and1 = u_CSAwallace_cska32_csa13_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa27_or0 = u_CSAwallace_cska32_csa13_csa_component_fa27_and0 | u_CSAwallace_cska32_csa13_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa27_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa28_and0 = u_CSAwallace_cska32_csa4_csa_component_fa27_or0 & u_CSAwallace_cska32_csa5_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa28_and1 = u_CSAwallace_cska32_csa13_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa28_or0 = u_CSAwallace_cska32_csa13_csa_component_fa28_and0 | u_CSAwallace_cska32_csa13_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa28_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa29_and0 = u_CSAwallace_cska32_csa4_csa_component_fa28_or0 & u_CSAwallace_cska32_csa5_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa29_and1 = u_CSAwallace_cska32_csa13_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa29_or0 = u_CSAwallace_cska32_csa13_csa_component_fa29_and0 | u_CSAwallace_cska32_csa13_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa29_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa30_and0 = u_CSAwallace_cska32_csa4_csa_component_fa29_or0 & u_CSAwallace_cska32_csa5_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa30_and1 = u_CSAwallace_cska32_csa13_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa30_or0 = u_CSAwallace_cska32_csa13_csa_component_fa30_and0 | u_CSAwallace_cska32_csa13_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa30_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa31_and0 = u_CSAwallace_cska32_csa4_csa_component_fa30_or0 & u_CSAwallace_cska32_csa5_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa31_and1 = u_CSAwallace_cska32_csa13_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa31_or0 = u_CSAwallace_cska32_csa13_csa_component_fa31_and0 | u_CSAwallace_cska32_csa13_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa31_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa32_and0 = u_CSAwallace_cska32_csa4_csa_component_fa31_or0 & u_CSAwallace_cska32_csa5_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa32_and1 = u_CSAwallace_cska32_csa13_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa32_or0 = u_CSAwallace_cska32_csa13_csa_component_fa32_and0 | u_CSAwallace_cska32_csa13_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa32_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa33_and0 = u_CSAwallace_cska32_csa4_csa_component_fa32_or0 & u_CSAwallace_cska32_csa5_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa33_and1 = u_CSAwallace_cska32_csa13_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa33_or0 = u_CSAwallace_cska32_csa13_csa_component_fa33_and0 | u_CSAwallace_cska32_csa13_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa33_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa34_and0 = u_CSAwallace_cska32_csa4_csa_component_fa33_or0 & u_CSAwallace_cska32_csa5_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa34_and1 = u_CSAwallace_cska32_csa13_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa34_or0 = u_CSAwallace_cska32_csa13_csa_component_fa34_and0 | u_CSAwallace_cska32_csa13_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa34_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa35_and0 = u_CSAwallace_cska32_csa4_csa_component_fa34_or0 & u_CSAwallace_cska32_csa5_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa35_and1 = u_CSAwallace_cska32_csa13_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa35_or0 = u_CSAwallace_cska32_csa13_csa_component_fa35_and0 | u_CSAwallace_cska32_csa13_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa35_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa36_and0 = u_CSAwallace_cska32_csa4_csa_component_fa35_or0 & u_CSAwallace_cska32_csa5_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa36_and1 = u_CSAwallace_cska32_csa13_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa36_or0 = u_CSAwallace_cska32_csa13_csa_component_fa36_and0 | u_CSAwallace_cska32_csa13_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa36_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa37_and0 = u_CSAwallace_cska32_csa4_csa_component_fa36_or0 & u_CSAwallace_cska32_csa5_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa37_and1 = u_CSAwallace_cska32_csa13_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa37_or0 = u_CSAwallace_cska32_csa13_csa_component_fa37_and0 | u_CSAwallace_cska32_csa13_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa37_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa38_and0 = u_CSAwallace_cska32_csa4_csa_component_fa37_or0 & u_CSAwallace_cska32_csa5_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa38_and1 = u_CSAwallace_cska32_csa13_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa38_or0 = u_CSAwallace_cska32_csa13_csa_component_fa38_and0 | u_CSAwallace_cska32_csa13_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa38_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa39_and0 = u_CSAwallace_cska32_csa4_csa_component_fa38_or0 & u_CSAwallace_cska32_csa5_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa39_and1 = u_CSAwallace_cska32_csa13_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa39_or0 = u_CSAwallace_cska32_csa13_csa_component_fa39_and0 | u_CSAwallace_cska32_csa13_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa39_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa40_and0 = u_CSAwallace_cska32_csa4_csa_component_fa39_or0 & u_CSAwallace_cska32_csa5_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa40_and1 = u_CSAwallace_cska32_csa13_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa40_or0 = u_CSAwallace_cska32_csa13_csa_component_fa40_and0 | u_CSAwallace_cska32_csa13_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa40_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa41_and0 = u_CSAwallace_cska32_csa4_csa_component_fa40_or0 & u_CSAwallace_cska32_csa5_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa41_and1 = u_CSAwallace_cska32_csa13_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa41_or0 = u_CSAwallace_cska32_csa13_csa_component_fa41_and0 | u_CSAwallace_cska32_csa13_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa41_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa42_and0 = u_CSAwallace_cska32_csa4_csa_component_fa41_or0 & u_CSAwallace_cska32_csa5_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa42_and1 = u_CSAwallace_cska32_csa13_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa42_or0 = u_CSAwallace_cska32_csa13_csa_component_fa42_and0 | u_CSAwallace_cska32_csa13_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa42_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa43_and0 = u_CSAwallace_cska32_csa4_csa_component_fa42_or0 & u_CSAwallace_cska32_csa5_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa43_and1 = u_CSAwallace_cska32_csa13_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa43_or0 = u_CSAwallace_cska32_csa13_csa_component_fa43_and0 | u_CSAwallace_cska32_csa13_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa43_or0 ^ u_CSAwallace_cska32_csa5_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa44_and0 = u_CSAwallace_cska32_csa4_csa_component_fa43_or0 & u_CSAwallace_cska32_csa5_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa44_and1 = u_CSAwallace_cska32_csa13_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa44_or0 = u_CSAwallace_cska32_csa13_csa_component_fa44_and0 | u_CSAwallace_cska32_csa13_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa4_csa_component_fa44_and1 ^ u_CSAwallace_cska32_csa5_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa45_and0 = u_CSAwallace_cska32_csa4_csa_component_fa44_and1 & u_CSAwallace_cska32_csa5_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa5_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa45_and1 = u_CSAwallace_cska32_csa13_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa5_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa45_or0 = u_CSAwallace_cska32_csa13_csa_component_fa45_and0 | u_CSAwallace_cska32_csa13_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa5_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa46_and1 = u_CSAwallace_cska32_csa5_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa5_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa5_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa5_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa47_and1 = u_CSAwallace_cska32_csa5_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa5_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa13_csa_component_fa48_xor1 = u_CSAwallace_cska32_and_31_17 ^ u_CSAwallace_cska32_csa5_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa13_csa_component_fa48_and1 = u_CSAwallace_cska32_and_31_17 & u_CSAwallace_cska32_csa5_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa19_and0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa20_and0 = u_CSAwallace_cska32_csa6_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa19_and0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa21_and0 = u_CSAwallace_cska32_csa6_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_and_0_21;
  assign u_CSAwallace_cska32_csa14_csa_component_fa21_and1 = u_CSAwallace_cska32_csa14_csa_component_fa21_xor0 & u_CSAwallace_cska32_and_0_21;
  assign u_CSAwallace_cska32_csa14_csa_component_fa21_or0 = u_CSAwallace_cska32_csa14_csa_component_fa21_and0 | u_CSAwallace_cska32_csa14_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa22_and0 = u_CSAwallace_cska32_csa6_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa22_xor0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa22_and1 = u_CSAwallace_cska32_csa14_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa22_xor0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa22_or0 = u_CSAwallace_cska32_csa14_csa_component_fa22_and0 | u_CSAwallace_cska32_csa14_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa23_and0 = u_CSAwallace_cska32_csa6_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa23_and1 = u_CSAwallace_cska32_csa14_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa23_or0 = u_CSAwallace_cska32_csa14_csa_component_fa23_and0 | u_CSAwallace_cska32_csa14_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa24_and0 = u_CSAwallace_cska32_csa6_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa24_and1 = u_CSAwallace_cska32_csa14_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa24_or0 = u_CSAwallace_cska32_csa14_csa_component_fa24_and0 | u_CSAwallace_cska32_csa14_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa25_and0 = u_CSAwallace_cska32_csa6_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa25_and1 = u_CSAwallace_cska32_csa14_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa25_or0 = u_CSAwallace_cska32_csa14_csa_component_fa25_and0 | u_CSAwallace_cska32_csa14_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa26_and0 = u_CSAwallace_cska32_csa6_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa26_and1 = u_CSAwallace_cska32_csa14_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa26_or0 = u_CSAwallace_cska32_csa14_csa_component_fa26_and0 | u_CSAwallace_cska32_csa14_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa27_and0 = u_CSAwallace_cska32_csa6_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa27_and1 = u_CSAwallace_cska32_csa14_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa27_or0 = u_CSAwallace_cska32_csa14_csa_component_fa27_and0 | u_CSAwallace_cska32_csa14_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa28_and0 = u_CSAwallace_cska32_csa6_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa28_and1 = u_CSAwallace_cska32_csa14_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa28_or0 = u_CSAwallace_cska32_csa14_csa_component_fa28_and0 | u_CSAwallace_cska32_csa14_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa29_and0 = u_CSAwallace_cska32_csa6_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa29_and1 = u_CSAwallace_cska32_csa14_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa29_or0 = u_CSAwallace_cska32_csa14_csa_component_fa29_and0 | u_CSAwallace_cska32_csa14_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa30_and0 = u_CSAwallace_cska32_csa6_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa30_and1 = u_CSAwallace_cska32_csa14_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa30_or0 = u_CSAwallace_cska32_csa14_csa_component_fa30_and0 | u_CSAwallace_cska32_csa14_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa31_and0 = u_CSAwallace_cska32_csa6_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa31_and1 = u_CSAwallace_cska32_csa14_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa31_or0 = u_CSAwallace_cska32_csa14_csa_component_fa31_and0 | u_CSAwallace_cska32_csa14_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa32_and0 = u_CSAwallace_cska32_csa6_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa32_and1 = u_CSAwallace_cska32_csa14_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa32_or0 = u_CSAwallace_cska32_csa14_csa_component_fa32_and0 | u_CSAwallace_cska32_csa14_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa33_and0 = u_CSAwallace_cska32_csa6_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa33_and1 = u_CSAwallace_cska32_csa14_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa33_or0 = u_CSAwallace_cska32_csa14_csa_component_fa33_and0 | u_CSAwallace_cska32_csa14_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa34_and0 = u_CSAwallace_cska32_csa6_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa34_and1 = u_CSAwallace_cska32_csa14_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa34_or0 = u_CSAwallace_cska32_csa14_csa_component_fa34_and0 | u_CSAwallace_cska32_csa14_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa35_and0 = u_CSAwallace_cska32_csa6_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa35_and1 = u_CSAwallace_cska32_csa14_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa35_or0 = u_CSAwallace_cska32_csa14_csa_component_fa35_and0 | u_CSAwallace_cska32_csa14_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa36_and0 = u_CSAwallace_cska32_csa6_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa36_and1 = u_CSAwallace_cska32_csa14_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa36_or0 = u_CSAwallace_cska32_csa14_csa_component_fa36_and0 | u_CSAwallace_cska32_csa14_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa37_and0 = u_CSAwallace_cska32_csa6_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa37_and1 = u_CSAwallace_cska32_csa14_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa37_or0 = u_CSAwallace_cska32_csa14_csa_component_fa37_and0 | u_CSAwallace_cska32_csa14_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa38_and0 = u_CSAwallace_cska32_csa6_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa38_and1 = u_CSAwallace_cska32_csa14_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa38_or0 = u_CSAwallace_cska32_csa14_csa_component_fa38_and0 | u_CSAwallace_cska32_csa14_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa39_and0 = u_CSAwallace_cska32_csa6_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa39_and1 = u_CSAwallace_cska32_csa14_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa39_or0 = u_CSAwallace_cska32_csa14_csa_component_fa39_and0 | u_CSAwallace_cska32_csa14_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa40_and0 = u_CSAwallace_cska32_csa6_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa40_and1 = u_CSAwallace_cska32_csa14_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa40_or0 = u_CSAwallace_cska32_csa14_csa_component_fa40_and0 | u_CSAwallace_cska32_csa14_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa41_and0 = u_CSAwallace_cska32_csa6_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa41_and1 = u_CSAwallace_cska32_csa14_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa41_or0 = u_CSAwallace_cska32_csa14_csa_component_fa41_and0 | u_CSAwallace_cska32_csa14_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa42_and0 = u_CSAwallace_cska32_csa6_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa42_and1 = u_CSAwallace_cska32_csa14_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa42_or0 = u_CSAwallace_cska32_csa14_csa_component_fa42_and0 | u_CSAwallace_cska32_csa14_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa43_and0 = u_CSAwallace_cska32_csa6_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa43_and1 = u_CSAwallace_cska32_csa14_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa43_or0 = u_CSAwallace_cska32_csa14_csa_component_fa43_and0 | u_CSAwallace_cska32_csa14_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa44_and0 = u_CSAwallace_cska32_csa6_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa44_and1 = u_CSAwallace_cska32_csa14_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa44_or0 = u_CSAwallace_cska32_csa14_csa_component_fa44_and0 | u_CSAwallace_cska32_csa14_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa45_and0 = u_CSAwallace_cska32_csa6_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa45_and1 = u_CSAwallace_cska32_csa14_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa45_or0 = u_CSAwallace_cska32_csa14_csa_component_fa45_and0 | u_CSAwallace_cska32_csa14_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa46_and0 = u_CSAwallace_cska32_csa6_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa46_and1 = u_CSAwallace_cska32_csa14_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa46_or0 = u_CSAwallace_cska32_csa14_csa_component_fa46_and0 | u_CSAwallace_cska32_csa14_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa47_and0 = u_CSAwallace_cska32_csa6_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa47_and1 = u_CSAwallace_cska32_csa14_csa_component_fa47_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa47_or0 = u_CSAwallace_cska32_csa14_csa_component_fa47_and0 | u_CSAwallace_cska32_csa14_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa48_and0 = u_CSAwallace_cska32_csa6_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa48_and1 = u_CSAwallace_cska32_csa14_csa_component_fa48_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa48_or0 = u_CSAwallace_cska32_csa14_csa_component_fa48_and0 | u_CSAwallace_cska32_csa14_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa49_and0 = u_CSAwallace_cska32_csa6_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa49_and1 = u_CSAwallace_cska32_csa14_csa_component_fa49_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa49_or0 = u_CSAwallace_cska32_csa14_csa_component_fa49_and0 | u_CSAwallace_cska32_csa14_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa6_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa6_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa50_and0 = u_CSAwallace_cska32_csa6_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa6_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa14_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa50_and1 = u_CSAwallace_cska32_csa14_csa_component_fa50_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa50_or0 = u_CSAwallace_cska32_csa14_csa_component_fa50_and0 | u_CSAwallace_cska32_csa14_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa51_xor0 = u_CSAwallace_cska32_and_31_20 ^ u_CSAwallace_cska32_csa6_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa51_and0 = u_CSAwallace_cska32_and_31_20 & u_CSAwallace_cska32_csa6_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_csa7_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa51_and1 = u_CSAwallace_cska32_csa14_csa_component_fa51_xor0 & u_CSAwallace_cska32_csa7_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa14_csa_component_fa51_or0 = u_CSAwallace_cska32_csa14_csa_component_fa51_and0 | u_CSAwallace_cska32_csa14_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa23_or0 ^ u_CSAwallace_cska32_and_0_24;
  assign u_CSAwallace_cska32_csa15_csa_component_fa24_and0 = u_CSAwallace_cska32_csa7_csa_component_fa23_or0 & u_CSAwallace_cska32_and_0_24;
  assign u_CSAwallace_cska32_csa15_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa24_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa25_xor0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa25_and0 = u_CSAwallace_cska32_csa7_csa_component_fa24_or0 & u_CSAwallace_cska32_csa8_csa_component_fa25_xor0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa25_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa26_and0 = u_CSAwallace_cska32_csa7_csa_component_fa25_or0 & u_CSAwallace_cska32_csa8_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa26_and1 = u_CSAwallace_cska32_csa15_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa26_or0 = u_CSAwallace_cska32_csa15_csa_component_fa26_and0 | u_CSAwallace_cska32_csa15_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa26_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa27_and0 = u_CSAwallace_cska32_csa7_csa_component_fa26_or0 & u_CSAwallace_cska32_csa8_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa27_and1 = u_CSAwallace_cska32_csa15_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa27_or0 = u_CSAwallace_cska32_csa15_csa_component_fa27_and0 | u_CSAwallace_cska32_csa15_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa27_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa28_and0 = u_CSAwallace_cska32_csa7_csa_component_fa27_or0 & u_CSAwallace_cska32_csa8_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa28_and1 = u_CSAwallace_cska32_csa15_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa28_or0 = u_CSAwallace_cska32_csa15_csa_component_fa28_and0 | u_CSAwallace_cska32_csa15_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa28_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa29_and0 = u_CSAwallace_cska32_csa7_csa_component_fa28_or0 & u_CSAwallace_cska32_csa8_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa29_and1 = u_CSAwallace_cska32_csa15_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa29_or0 = u_CSAwallace_cska32_csa15_csa_component_fa29_and0 | u_CSAwallace_cska32_csa15_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa29_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa30_and0 = u_CSAwallace_cska32_csa7_csa_component_fa29_or0 & u_CSAwallace_cska32_csa8_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa30_and1 = u_CSAwallace_cska32_csa15_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa30_or0 = u_CSAwallace_cska32_csa15_csa_component_fa30_and0 | u_CSAwallace_cska32_csa15_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa30_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa31_and0 = u_CSAwallace_cska32_csa7_csa_component_fa30_or0 & u_CSAwallace_cska32_csa8_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa31_and1 = u_CSAwallace_cska32_csa15_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa31_or0 = u_CSAwallace_cska32_csa15_csa_component_fa31_and0 | u_CSAwallace_cska32_csa15_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa31_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa32_and0 = u_CSAwallace_cska32_csa7_csa_component_fa31_or0 & u_CSAwallace_cska32_csa8_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa32_and1 = u_CSAwallace_cska32_csa15_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa32_or0 = u_CSAwallace_cska32_csa15_csa_component_fa32_and0 | u_CSAwallace_cska32_csa15_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa32_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa33_and0 = u_CSAwallace_cska32_csa7_csa_component_fa32_or0 & u_CSAwallace_cska32_csa8_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa33_and1 = u_CSAwallace_cska32_csa15_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa33_or0 = u_CSAwallace_cska32_csa15_csa_component_fa33_and0 | u_CSAwallace_cska32_csa15_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa33_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa34_and0 = u_CSAwallace_cska32_csa7_csa_component_fa33_or0 & u_CSAwallace_cska32_csa8_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa34_and1 = u_CSAwallace_cska32_csa15_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa34_or0 = u_CSAwallace_cska32_csa15_csa_component_fa34_and0 | u_CSAwallace_cska32_csa15_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa34_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa35_and0 = u_CSAwallace_cska32_csa7_csa_component_fa34_or0 & u_CSAwallace_cska32_csa8_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa35_and1 = u_CSAwallace_cska32_csa15_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa35_or0 = u_CSAwallace_cska32_csa15_csa_component_fa35_and0 | u_CSAwallace_cska32_csa15_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa35_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa36_and0 = u_CSAwallace_cska32_csa7_csa_component_fa35_or0 & u_CSAwallace_cska32_csa8_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa36_and1 = u_CSAwallace_cska32_csa15_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa36_or0 = u_CSAwallace_cska32_csa15_csa_component_fa36_and0 | u_CSAwallace_cska32_csa15_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa36_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa37_and0 = u_CSAwallace_cska32_csa7_csa_component_fa36_or0 & u_CSAwallace_cska32_csa8_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa37_and1 = u_CSAwallace_cska32_csa15_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa37_or0 = u_CSAwallace_cska32_csa15_csa_component_fa37_and0 | u_CSAwallace_cska32_csa15_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa37_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa38_and0 = u_CSAwallace_cska32_csa7_csa_component_fa37_or0 & u_CSAwallace_cska32_csa8_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa38_and1 = u_CSAwallace_cska32_csa15_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa38_or0 = u_CSAwallace_cska32_csa15_csa_component_fa38_and0 | u_CSAwallace_cska32_csa15_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa38_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa39_and0 = u_CSAwallace_cska32_csa7_csa_component_fa38_or0 & u_CSAwallace_cska32_csa8_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa39_and1 = u_CSAwallace_cska32_csa15_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa39_or0 = u_CSAwallace_cska32_csa15_csa_component_fa39_and0 | u_CSAwallace_cska32_csa15_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa39_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa40_and0 = u_CSAwallace_cska32_csa7_csa_component_fa39_or0 & u_CSAwallace_cska32_csa8_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa40_and1 = u_CSAwallace_cska32_csa15_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa40_or0 = u_CSAwallace_cska32_csa15_csa_component_fa40_and0 | u_CSAwallace_cska32_csa15_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa40_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa41_and0 = u_CSAwallace_cska32_csa7_csa_component_fa40_or0 & u_CSAwallace_cska32_csa8_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa41_and1 = u_CSAwallace_cska32_csa15_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa41_or0 = u_CSAwallace_cska32_csa15_csa_component_fa41_and0 | u_CSAwallace_cska32_csa15_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa41_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa42_and0 = u_CSAwallace_cska32_csa7_csa_component_fa41_or0 & u_CSAwallace_cska32_csa8_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa42_and1 = u_CSAwallace_cska32_csa15_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa42_or0 = u_CSAwallace_cska32_csa15_csa_component_fa42_and0 | u_CSAwallace_cska32_csa15_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa42_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa43_and0 = u_CSAwallace_cska32_csa7_csa_component_fa42_or0 & u_CSAwallace_cska32_csa8_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa43_and1 = u_CSAwallace_cska32_csa15_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa43_or0 = u_CSAwallace_cska32_csa15_csa_component_fa43_and0 | u_CSAwallace_cska32_csa15_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa43_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa44_and0 = u_CSAwallace_cska32_csa7_csa_component_fa43_or0 & u_CSAwallace_cska32_csa8_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa44_and1 = u_CSAwallace_cska32_csa15_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa44_or0 = u_CSAwallace_cska32_csa15_csa_component_fa44_and0 | u_CSAwallace_cska32_csa15_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa44_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa45_and0 = u_CSAwallace_cska32_csa7_csa_component_fa44_or0 & u_CSAwallace_cska32_csa8_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa45_and1 = u_CSAwallace_cska32_csa15_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa45_or0 = u_CSAwallace_cska32_csa15_csa_component_fa45_and0 | u_CSAwallace_cska32_csa15_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa45_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa46_and0 = u_CSAwallace_cska32_csa7_csa_component_fa45_or0 & u_CSAwallace_cska32_csa8_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa46_and1 = u_CSAwallace_cska32_csa15_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa46_or0 = u_CSAwallace_cska32_csa15_csa_component_fa46_and0 | u_CSAwallace_cska32_csa15_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa46_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa47_and0 = u_CSAwallace_cska32_csa7_csa_component_fa46_or0 & u_CSAwallace_cska32_csa8_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa47_and1 = u_CSAwallace_cska32_csa15_csa_component_fa47_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa47_or0 = u_CSAwallace_cska32_csa15_csa_component_fa47_and0 | u_CSAwallace_cska32_csa15_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa47_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa48_and0 = u_CSAwallace_cska32_csa7_csa_component_fa47_or0 & u_CSAwallace_cska32_csa8_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa48_and1 = u_CSAwallace_cska32_csa15_csa_component_fa48_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa48_or0 = u_CSAwallace_cska32_csa15_csa_component_fa48_and0 | u_CSAwallace_cska32_csa15_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa48_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa49_and0 = u_CSAwallace_cska32_csa7_csa_component_fa48_or0 & u_CSAwallace_cska32_csa8_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa49_and1 = u_CSAwallace_cska32_csa15_csa_component_fa49_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa49_or0 = u_CSAwallace_cska32_csa15_csa_component_fa49_and0 | u_CSAwallace_cska32_csa15_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa49_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa50_and0 = u_CSAwallace_cska32_csa7_csa_component_fa49_or0 & u_CSAwallace_cska32_csa8_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa50_and1 = u_CSAwallace_cska32_csa15_csa_component_fa50_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa50_or0 = u_CSAwallace_cska32_csa15_csa_component_fa50_and0 | u_CSAwallace_cska32_csa15_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa51_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa50_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa51_and0 = u_CSAwallace_cska32_csa7_csa_component_fa50_or0 & u_CSAwallace_cska32_csa8_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa51_and1 = u_CSAwallace_cska32_csa15_csa_component_fa51_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa51_or0 = u_CSAwallace_cska32_csa15_csa_component_fa51_and0 | u_CSAwallace_cska32_csa15_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa52_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa51_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa52_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa52_and0 = u_CSAwallace_cska32_csa7_csa_component_fa51_or0 & u_CSAwallace_cska32_csa8_csa_component_fa52_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa52_and1 = u_CSAwallace_cska32_csa15_csa_component_fa52_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa52_or0 = u_CSAwallace_cska32_csa15_csa_component_fa52_and0 | u_CSAwallace_cska32_csa15_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa53_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa52_or0 ^ u_CSAwallace_cska32_csa8_csa_component_fa53_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa53_and0 = u_CSAwallace_cska32_csa7_csa_component_fa52_or0 & u_CSAwallace_cska32_csa8_csa_component_fa53_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa53_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa53_and1 = u_CSAwallace_cska32_csa15_csa_component_fa53_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa53_or0 = u_CSAwallace_cska32_csa15_csa_component_fa53_and0 | u_CSAwallace_cska32_csa15_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa54_xor0 = u_CSAwallace_cska32_csa7_csa_component_fa53_and1 ^ u_CSAwallace_cska32_csa8_csa_component_fa54_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa54_and0 = u_CSAwallace_cska32_csa7_csa_component_fa53_and1 & u_CSAwallace_cska32_csa8_csa_component_fa54_xor1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa54_xor0 ^ u_CSAwallace_cska32_csa8_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa54_and1 = u_CSAwallace_cska32_csa15_csa_component_fa54_xor0 & u_CSAwallace_cska32_csa8_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa54_or0 = u_CSAwallace_cska32_csa15_csa_component_fa54_and0 | u_CSAwallace_cska32_csa15_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa8_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa55_and1 = u_CSAwallace_cska32_csa8_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa8_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa8_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa8_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa56_and1 = u_CSAwallace_cska32_csa8_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa8_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa15_csa_component_fa57_xor1 = u_CSAwallace_cska32_and_31_26 ^ u_CSAwallace_cska32_csa8_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa15_csa_component_fa57_and1 = u_CSAwallace_cska32_and_31_26 & u_CSAwallace_cska32_csa8_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa28_and0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa29_and0 = u_CSAwallace_cska32_csa9_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa28_and0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa30_and0 = u_CSAwallace_cska32_csa9_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_and_0_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa30_and1 = u_CSAwallace_cska32_csa16_csa_component_fa30_xor0 & u_CSAwallace_cska32_and_0_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa30_or0 = u_CSAwallace_cska32_csa16_csa_component_fa30_and0 | u_CSAwallace_cska32_csa16_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa31_and0 = u_CSAwallace_cska32_csa9_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_1_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa31_and1 = u_CSAwallace_cska32_csa16_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_1_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa31_or0 = u_CSAwallace_cska32_csa16_csa_component_fa31_and0 | u_CSAwallace_cska32_csa16_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa32_and0 = u_CSAwallace_cska32_csa9_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_2_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa32_and1 = u_CSAwallace_cska32_csa16_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_2_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa32_or0 = u_CSAwallace_cska32_csa16_csa_component_fa32_and0 | u_CSAwallace_cska32_csa16_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa33_and0 = u_CSAwallace_cska32_csa9_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_3_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa33_and1 = u_CSAwallace_cska32_csa16_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_3_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa33_or0 = u_CSAwallace_cska32_csa16_csa_component_fa33_and0 | u_CSAwallace_cska32_csa16_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa34_and0 = u_CSAwallace_cska32_csa9_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_4_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa34_and1 = u_CSAwallace_cska32_csa16_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_4_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa34_or0 = u_CSAwallace_cska32_csa16_csa_component_fa34_and0 | u_CSAwallace_cska32_csa16_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa35_and0 = u_CSAwallace_cska32_csa9_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_5_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa35_and1 = u_CSAwallace_cska32_csa16_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_5_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa35_or0 = u_CSAwallace_cska32_csa16_csa_component_fa35_and0 | u_CSAwallace_cska32_csa16_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa36_and0 = u_CSAwallace_cska32_csa9_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_6_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa36_and1 = u_CSAwallace_cska32_csa16_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_6_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa36_or0 = u_CSAwallace_cska32_csa16_csa_component_fa36_and0 | u_CSAwallace_cska32_csa16_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa37_and0 = u_CSAwallace_cska32_csa9_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_7_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa37_and1 = u_CSAwallace_cska32_csa16_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_7_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa37_or0 = u_CSAwallace_cska32_csa16_csa_component_fa37_and0 | u_CSAwallace_cska32_csa16_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa38_and0 = u_CSAwallace_cska32_csa9_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_8_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa38_and1 = u_CSAwallace_cska32_csa16_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_8_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa38_or0 = u_CSAwallace_cska32_csa16_csa_component_fa38_and0 | u_CSAwallace_cska32_csa16_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa39_and0 = u_CSAwallace_cska32_csa9_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_9_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa39_and1 = u_CSAwallace_cska32_csa16_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_9_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa39_or0 = u_CSAwallace_cska32_csa16_csa_component_fa39_and0 | u_CSAwallace_cska32_csa16_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa40_and0 = u_CSAwallace_cska32_csa9_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_10_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa40_and1 = u_CSAwallace_cska32_csa16_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_10_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa40_or0 = u_CSAwallace_cska32_csa16_csa_component_fa40_and0 | u_CSAwallace_cska32_csa16_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa41_and0 = u_CSAwallace_cska32_csa9_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_and_11_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa41_and1 = u_CSAwallace_cska32_csa16_csa_component_fa41_xor0 & u_CSAwallace_cska32_and_11_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa41_or0 = u_CSAwallace_cska32_csa16_csa_component_fa41_and0 | u_CSAwallace_cska32_csa16_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa42_and0 = u_CSAwallace_cska32_csa9_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_and_12_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa42_and1 = u_CSAwallace_cska32_csa16_csa_component_fa42_xor0 & u_CSAwallace_cska32_and_12_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa42_or0 = u_CSAwallace_cska32_csa16_csa_component_fa42_and0 | u_CSAwallace_cska32_csa16_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa43_and0 = u_CSAwallace_cska32_csa9_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_and_13_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa43_and1 = u_CSAwallace_cska32_csa16_csa_component_fa43_xor0 & u_CSAwallace_cska32_and_13_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa43_or0 = u_CSAwallace_cska32_csa16_csa_component_fa43_and0 | u_CSAwallace_cska32_csa16_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa44_and0 = u_CSAwallace_cska32_csa9_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_and_14_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa44_and1 = u_CSAwallace_cska32_csa16_csa_component_fa44_xor0 & u_CSAwallace_cska32_and_14_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa44_or0 = u_CSAwallace_cska32_csa16_csa_component_fa44_and0 | u_CSAwallace_cska32_csa16_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa45_and0 = u_CSAwallace_cska32_csa9_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_and_15_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa45_and1 = u_CSAwallace_cska32_csa16_csa_component_fa45_xor0 & u_CSAwallace_cska32_and_15_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa45_or0 = u_CSAwallace_cska32_csa16_csa_component_fa45_and0 | u_CSAwallace_cska32_csa16_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa46_and0 = u_CSAwallace_cska32_csa9_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_and_16_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa46_and1 = u_CSAwallace_cska32_csa16_csa_component_fa46_xor0 & u_CSAwallace_cska32_and_16_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa46_or0 = u_CSAwallace_cska32_csa16_csa_component_fa46_and0 | u_CSAwallace_cska32_csa16_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa47_and0 = u_CSAwallace_cska32_csa9_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_and_17_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa47_and1 = u_CSAwallace_cska32_csa16_csa_component_fa47_xor0 & u_CSAwallace_cska32_and_17_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa47_or0 = u_CSAwallace_cska32_csa16_csa_component_fa47_and0 | u_CSAwallace_cska32_csa16_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa48_and0 = u_CSAwallace_cska32_csa9_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_and_18_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa48_and1 = u_CSAwallace_cska32_csa16_csa_component_fa48_xor0 & u_CSAwallace_cska32_and_18_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa48_or0 = u_CSAwallace_cska32_csa16_csa_component_fa48_and0 | u_CSAwallace_cska32_csa16_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa49_and0 = u_CSAwallace_cska32_csa9_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_and_19_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa49_and1 = u_CSAwallace_cska32_csa16_csa_component_fa49_xor0 & u_CSAwallace_cska32_and_19_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa49_or0 = u_CSAwallace_cska32_csa16_csa_component_fa49_and0 | u_CSAwallace_cska32_csa16_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa50_and0 = u_CSAwallace_cska32_csa9_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_and_20_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa50_and1 = u_CSAwallace_cska32_csa16_csa_component_fa50_xor0 & u_CSAwallace_cska32_and_20_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa50_or0 = u_CSAwallace_cska32_csa16_csa_component_fa50_and0 | u_CSAwallace_cska32_csa16_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa51_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa51_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa51_and0 = u_CSAwallace_cska32_csa9_csa_component_fa51_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_and_21_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa51_and1 = u_CSAwallace_cska32_csa16_csa_component_fa51_xor0 & u_CSAwallace_cska32_and_21_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa51_or0 = u_CSAwallace_cska32_csa16_csa_component_fa51_and0 | u_CSAwallace_cska32_csa16_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa52_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa52_and0 = u_CSAwallace_cska32_csa9_csa_component_fa52_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_and_22_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa52_and1 = u_CSAwallace_cska32_csa16_csa_component_fa52_xor0 & u_CSAwallace_cska32_and_22_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa52_or0 = u_CSAwallace_cska32_csa16_csa_component_fa52_and0 | u_CSAwallace_cska32_csa16_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa53_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa53_and0 = u_CSAwallace_cska32_csa9_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa53_xor0 ^ u_CSAwallace_cska32_and_23_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa53_and1 = u_CSAwallace_cska32_csa16_csa_component_fa53_xor0 & u_CSAwallace_cska32_and_23_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa53_or0 = u_CSAwallace_cska32_csa16_csa_component_fa53_and0 | u_CSAwallace_cska32_csa16_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa54_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa54_and0 = u_CSAwallace_cska32_csa9_csa_component_fa54_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa54_xor0 ^ u_CSAwallace_cska32_and_24_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa54_and1 = u_CSAwallace_cska32_csa16_csa_component_fa54_xor0 & u_CSAwallace_cska32_and_24_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa54_or0 = u_CSAwallace_cska32_csa16_csa_component_fa54_and0 | u_CSAwallace_cska32_csa16_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa55_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa55_and0 = u_CSAwallace_cska32_csa9_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa55_xor0 ^ u_CSAwallace_cska32_and_25_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa55_and1 = u_CSAwallace_cska32_csa16_csa_component_fa55_xor0 & u_CSAwallace_cska32_and_25_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa55_or0 = u_CSAwallace_cska32_csa16_csa_component_fa55_and0 | u_CSAwallace_cska32_csa16_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa56_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa56_and0 = u_CSAwallace_cska32_csa9_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa56_xor0 ^ u_CSAwallace_cska32_and_26_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa56_and1 = u_CSAwallace_cska32_csa16_csa_component_fa56_xor0 & u_CSAwallace_cska32_and_26_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa56_or0 = u_CSAwallace_cska32_csa16_csa_component_fa56_and0 | u_CSAwallace_cska32_csa16_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa57_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa57_and0 = u_CSAwallace_cska32_csa9_csa_component_fa57_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa57_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa57_xor0 ^ u_CSAwallace_cska32_and_27_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa57_and1 = u_CSAwallace_cska32_csa16_csa_component_fa57_xor0 & u_CSAwallace_cska32_and_27_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa57_or0 = u_CSAwallace_cska32_csa16_csa_component_fa57_and0 | u_CSAwallace_cska32_csa16_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa58_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa58_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa58_and0 = u_CSAwallace_cska32_csa9_csa_component_fa58_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa58_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa58_xor0 ^ u_CSAwallace_cska32_and_28_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa58_and1 = u_CSAwallace_cska32_csa16_csa_component_fa58_xor0 & u_CSAwallace_cska32_and_28_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa58_or0 = u_CSAwallace_cska32_csa16_csa_component_fa58_and0 | u_CSAwallace_cska32_csa16_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa59_xor0 = u_CSAwallace_cska32_csa9_csa_component_fa59_xor1 ^ u_CSAwallace_cska32_csa9_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa59_and0 = u_CSAwallace_cska32_csa9_csa_component_fa59_xor1 & u_CSAwallace_cska32_csa9_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_csa16_csa_component_fa59_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa59_xor0 ^ u_CSAwallace_cska32_and_29_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa59_and1 = u_CSAwallace_cska32_csa16_csa_component_fa59_xor0 & u_CSAwallace_cska32_and_29_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa59_or0 = u_CSAwallace_cska32_csa16_csa_component_fa59_and0 | u_CSAwallace_cska32_csa16_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa60_xor0 = u_CSAwallace_cska32_and_31_29 ^ u_CSAwallace_cska32_csa9_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa60_and0 = u_CSAwallace_cska32_and_31_29 & u_CSAwallace_cska32_csa9_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa16_csa_component_fa60_xor1 = u_CSAwallace_cska32_csa16_csa_component_fa60_xor0 ^ u_CSAwallace_cska32_and_30_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa60_and1 = u_CSAwallace_cska32_csa16_csa_component_fa60_xor0 & u_CSAwallace_cska32_and_30_30;
  assign u_CSAwallace_cska32_csa16_csa_component_fa60_or0 = u_CSAwallace_cska32_csa16_csa_component_fa60_and0 | u_CSAwallace_cska32_csa16_csa_component_fa60_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa3_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa3_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa2_and0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa3_and0 = u_CSAwallace_cska32_csa10_csa_component_fa3_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa2_and0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa4_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa4_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa3_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa4_and0 = u_CSAwallace_cska32_csa10_csa_component_fa4_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa3_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa5_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa5_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa4_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa5_and0 = u_CSAwallace_cska32_csa10_csa_component_fa5_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa4_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa5_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa5_xor0 ^ u_CSAwallace_cska32_csa1_csa_component_fa4_and0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa5_and1 = u_CSAwallace_cska32_csa17_csa_component_fa5_xor0 & u_CSAwallace_cska32_csa1_csa_component_fa4_and0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa5_or0 = u_CSAwallace_cska32_csa17_csa_component_fa5_and0 | u_CSAwallace_cska32_csa17_csa_component_fa5_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa6_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa6_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa5_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa6_and0 = u_CSAwallace_cska32_csa10_csa_component_fa6_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa5_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa6_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa6_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa6_xor0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa6_and1 = u_CSAwallace_cska32_csa17_csa_component_fa6_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa6_xor0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa6_or0 = u_CSAwallace_cska32_csa17_csa_component_fa6_and0 | u_CSAwallace_cska32_csa17_csa_component_fa6_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa7_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa7_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa6_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa7_and0 = u_CSAwallace_cska32_csa10_csa_component_fa7_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa6_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa7_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa7_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa7_xor0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa7_and1 = u_CSAwallace_cska32_csa17_csa_component_fa7_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa7_xor0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa7_or0 = u_CSAwallace_cska32_csa17_csa_component_fa7_and0 | u_CSAwallace_cska32_csa17_csa_component_fa7_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa8_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa8_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa7_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa8_and0 = u_CSAwallace_cska32_csa10_csa_component_fa8_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa7_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa8_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa8_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa8_and1 = u_CSAwallace_cska32_csa17_csa_component_fa8_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa8_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa8_or0 = u_CSAwallace_cska32_csa17_csa_component_fa8_and0 | u_CSAwallace_cska32_csa17_csa_component_fa8_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa9_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa9_and0 = u_CSAwallace_cska32_csa10_csa_component_fa9_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa9_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa9_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa9_and1 = u_CSAwallace_cska32_csa17_csa_component_fa9_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa9_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa9_or0 = u_CSAwallace_cska32_csa17_csa_component_fa9_and0 | u_CSAwallace_cska32_csa17_csa_component_fa9_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa10_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa10_and0 = u_CSAwallace_cska32_csa10_csa_component_fa10_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa10_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa10_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa10_and1 = u_CSAwallace_cska32_csa17_csa_component_fa10_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa10_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa10_or0 = u_CSAwallace_cska32_csa17_csa_component_fa10_and0 | u_CSAwallace_cska32_csa17_csa_component_fa10_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa11_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa11_and0 = u_CSAwallace_cska32_csa10_csa_component_fa11_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa11_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa11_and1 = u_CSAwallace_cska32_csa17_csa_component_fa11_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa11_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa11_or0 = u_CSAwallace_cska32_csa17_csa_component_fa11_and0 | u_CSAwallace_cska32_csa17_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa12_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa12_and0 = u_CSAwallace_cska32_csa10_csa_component_fa12_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa12_and1 = u_CSAwallace_cska32_csa17_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa12_or0 = u_CSAwallace_cska32_csa17_csa_component_fa12_and0 | u_CSAwallace_cska32_csa17_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa13_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa13_and0 = u_CSAwallace_cska32_csa10_csa_component_fa13_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa13_and1 = u_CSAwallace_cska32_csa17_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa13_or0 = u_CSAwallace_cska32_csa17_csa_component_fa13_and0 | u_CSAwallace_cska32_csa17_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa14_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa14_and0 = u_CSAwallace_cska32_csa10_csa_component_fa14_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa14_and1 = u_CSAwallace_cska32_csa17_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa14_or0 = u_CSAwallace_cska32_csa17_csa_component_fa14_and0 | u_CSAwallace_cska32_csa17_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa15_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa15_and0 = u_CSAwallace_cska32_csa10_csa_component_fa15_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa15_and1 = u_CSAwallace_cska32_csa17_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa15_or0 = u_CSAwallace_cska32_csa17_csa_component_fa15_and0 | u_CSAwallace_cska32_csa17_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa16_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa16_and0 = u_CSAwallace_cska32_csa10_csa_component_fa16_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa16_and1 = u_CSAwallace_cska32_csa17_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa16_or0 = u_CSAwallace_cska32_csa17_csa_component_fa16_and0 | u_CSAwallace_cska32_csa17_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa17_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa17_and0 = u_CSAwallace_cska32_csa10_csa_component_fa17_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa17_and1 = u_CSAwallace_cska32_csa17_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa17_or0 = u_CSAwallace_cska32_csa17_csa_component_fa17_and0 | u_CSAwallace_cska32_csa17_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa18_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa18_and0 = u_CSAwallace_cska32_csa10_csa_component_fa18_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa18_and1 = u_CSAwallace_cska32_csa17_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa18_or0 = u_CSAwallace_cska32_csa17_csa_component_fa18_and0 | u_CSAwallace_cska32_csa17_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa19_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa19_and0 = u_CSAwallace_cska32_csa10_csa_component_fa19_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa19_and1 = u_CSAwallace_cska32_csa17_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa19_or0 = u_CSAwallace_cska32_csa17_csa_component_fa19_and0 | u_CSAwallace_cska32_csa17_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa20_and0 = u_CSAwallace_cska32_csa10_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa20_and1 = u_CSAwallace_cska32_csa17_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa20_or0 = u_CSAwallace_cska32_csa17_csa_component_fa20_and0 | u_CSAwallace_cska32_csa17_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa21_and0 = u_CSAwallace_cska32_csa10_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa21_and1 = u_CSAwallace_cska32_csa17_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa21_or0 = u_CSAwallace_cska32_csa17_csa_component_fa21_and0 | u_CSAwallace_cska32_csa17_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa22_and0 = u_CSAwallace_cska32_csa10_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa22_and1 = u_CSAwallace_cska32_csa17_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa22_or0 = u_CSAwallace_cska32_csa17_csa_component_fa22_and0 | u_CSAwallace_cska32_csa17_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa23_and0 = u_CSAwallace_cska32_csa10_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa23_and1 = u_CSAwallace_cska32_csa17_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa23_or0 = u_CSAwallace_cska32_csa17_csa_component_fa23_and0 | u_CSAwallace_cska32_csa17_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa24_and0 = u_CSAwallace_cska32_csa10_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa24_and1 = u_CSAwallace_cska32_csa17_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa24_or0 = u_CSAwallace_cska32_csa17_csa_component_fa24_and0 | u_CSAwallace_cska32_csa17_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa25_and0 = u_CSAwallace_cska32_csa10_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa25_and1 = u_CSAwallace_cska32_csa17_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa25_or0 = u_CSAwallace_cska32_csa17_csa_component_fa25_and0 | u_CSAwallace_cska32_csa17_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa26_and0 = u_CSAwallace_cska32_csa10_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa26_and1 = u_CSAwallace_cska32_csa17_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa26_or0 = u_CSAwallace_cska32_csa17_csa_component_fa26_and0 | u_CSAwallace_cska32_csa17_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa27_and0 = u_CSAwallace_cska32_csa10_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa27_and1 = u_CSAwallace_cska32_csa17_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa27_or0 = u_CSAwallace_cska32_csa17_csa_component_fa27_and0 | u_CSAwallace_cska32_csa17_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa28_and0 = u_CSAwallace_cska32_csa10_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa28_and1 = u_CSAwallace_cska32_csa17_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa28_or0 = u_CSAwallace_cska32_csa17_csa_component_fa28_and0 | u_CSAwallace_cska32_csa17_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa29_and0 = u_CSAwallace_cska32_csa10_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa29_and1 = u_CSAwallace_cska32_csa17_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa29_or0 = u_CSAwallace_cska32_csa17_csa_component_fa29_and0 | u_CSAwallace_cska32_csa17_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa30_and0 = u_CSAwallace_cska32_csa10_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa30_and1 = u_CSAwallace_cska32_csa17_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa30_or0 = u_CSAwallace_cska32_csa17_csa_component_fa30_and0 | u_CSAwallace_cska32_csa17_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa31_and0 = u_CSAwallace_cska32_csa10_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa31_and1 = u_CSAwallace_cska32_csa17_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa31_or0 = u_CSAwallace_cska32_csa17_csa_component_fa31_and0 | u_CSAwallace_cska32_csa17_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa32_and0 = u_CSAwallace_cska32_csa10_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa32_and1 = u_CSAwallace_cska32_csa17_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa32_or0 = u_CSAwallace_cska32_csa17_csa_component_fa32_and0 | u_CSAwallace_cska32_csa17_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa10_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa33_and0 = u_CSAwallace_cska32_csa10_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa33_and1 = u_CSAwallace_cska32_csa17_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa33_or0 = u_CSAwallace_cska32_csa17_csa_component_fa33_and0 | u_CSAwallace_cska32_csa17_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa1_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa10_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa34_and0 = u_CSAwallace_cska32_csa1_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa10_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa17_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa17_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa34_and1 = u_CSAwallace_cska32_csa17_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa34_or0 = u_CSAwallace_cska32_csa17_csa_component_fa34_and0 | u_CSAwallace_cska32_csa17_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa1_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa11_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa35_and1 = u_CSAwallace_cska32_csa1_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa11_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa36_xor1 = u_CSAwallace_cska32_and_31_5 ^ u_CSAwallace_cska32_csa11_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa17_csa_component_fa36_and1 = u_CSAwallace_cska32_and_31_5 & u_CSAwallace_cska32_csa11_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa8_or0 ^ u_CSAwallace_cska32_and_0_9;
  assign u_CSAwallace_cska32_csa18_csa_component_fa9_and0 = u_CSAwallace_cska32_csa11_csa_component_fa8_or0 & u_CSAwallace_cska32_and_0_9;
  assign u_CSAwallace_cska32_csa18_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa9_or0 ^ u_CSAwallace_cska32_csa3_csa_component_fa10_xor0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa10_and0 = u_CSAwallace_cska32_csa11_csa_component_fa9_or0 & u_CSAwallace_cska32_csa3_csa_component_fa10_xor0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa10_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa11_xor0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa11_and0 = u_CSAwallace_cska32_csa11_csa_component_fa10_or0 & u_CSAwallace_cska32_csa12_csa_component_fa11_xor0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa11_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa12_and0 = u_CSAwallace_cska32_csa11_csa_component_fa11_or0 & u_CSAwallace_cska32_csa12_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa12_and1 = u_CSAwallace_cska32_csa18_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa12_or0 = u_CSAwallace_cska32_csa18_csa_component_fa12_and0 | u_CSAwallace_cska32_csa18_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa12_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa13_and0 = u_CSAwallace_cska32_csa11_csa_component_fa12_or0 & u_CSAwallace_cska32_csa12_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa13_and1 = u_CSAwallace_cska32_csa18_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa13_or0 = u_CSAwallace_cska32_csa18_csa_component_fa13_and0 | u_CSAwallace_cska32_csa18_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa13_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa14_and0 = u_CSAwallace_cska32_csa11_csa_component_fa13_or0 & u_CSAwallace_cska32_csa12_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa14_and1 = u_CSAwallace_cska32_csa18_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa14_or0 = u_CSAwallace_cska32_csa18_csa_component_fa14_and0 | u_CSAwallace_cska32_csa18_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa14_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa15_and0 = u_CSAwallace_cska32_csa11_csa_component_fa14_or0 & u_CSAwallace_cska32_csa12_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa15_and1 = u_CSAwallace_cska32_csa18_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa15_or0 = u_CSAwallace_cska32_csa18_csa_component_fa15_and0 | u_CSAwallace_cska32_csa18_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa15_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa16_and0 = u_CSAwallace_cska32_csa11_csa_component_fa15_or0 & u_CSAwallace_cska32_csa12_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa16_and1 = u_CSAwallace_cska32_csa18_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa16_or0 = u_CSAwallace_cska32_csa18_csa_component_fa16_and0 | u_CSAwallace_cska32_csa18_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa16_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa17_and0 = u_CSAwallace_cska32_csa11_csa_component_fa16_or0 & u_CSAwallace_cska32_csa12_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa17_and1 = u_CSAwallace_cska32_csa18_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa17_or0 = u_CSAwallace_cska32_csa18_csa_component_fa17_and0 | u_CSAwallace_cska32_csa18_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa17_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa18_and0 = u_CSAwallace_cska32_csa11_csa_component_fa17_or0 & u_CSAwallace_cska32_csa12_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa18_and1 = u_CSAwallace_cska32_csa18_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa18_or0 = u_CSAwallace_cska32_csa18_csa_component_fa18_and0 | u_CSAwallace_cska32_csa18_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa18_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa19_and0 = u_CSAwallace_cska32_csa11_csa_component_fa18_or0 & u_CSAwallace_cska32_csa12_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa19_and1 = u_CSAwallace_cska32_csa18_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa19_or0 = u_CSAwallace_cska32_csa18_csa_component_fa19_and0 | u_CSAwallace_cska32_csa18_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa19_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa20_and0 = u_CSAwallace_cska32_csa11_csa_component_fa19_or0 & u_CSAwallace_cska32_csa12_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa20_and1 = u_CSAwallace_cska32_csa18_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa20_or0 = u_CSAwallace_cska32_csa18_csa_component_fa20_and0 | u_CSAwallace_cska32_csa18_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa20_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa21_and0 = u_CSAwallace_cska32_csa11_csa_component_fa20_or0 & u_CSAwallace_cska32_csa12_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa21_and1 = u_CSAwallace_cska32_csa18_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa21_or0 = u_CSAwallace_cska32_csa18_csa_component_fa21_and0 | u_CSAwallace_cska32_csa18_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa21_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa22_and0 = u_CSAwallace_cska32_csa11_csa_component_fa21_or0 & u_CSAwallace_cska32_csa12_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa22_and1 = u_CSAwallace_cska32_csa18_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa22_or0 = u_CSAwallace_cska32_csa18_csa_component_fa22_and0 | u_CSAwallace_cska32_csa18_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa22_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa23_and0 = u_CSAwallace_cska32_csa11_csa_component_fa22_or0 & u_CSAwallace_cska32_csa12_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa23_and1 = u_CSAwallace_cska32_csa18_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa23_or0 = u_CSAwallace_cska32_csa18_csa_component_fa23_and0 | u_CSAwallace_cska32_csa18_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa23_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa24_and0 = u_CSAwallace_cska32_csa11_csa_component_fa23_or0 & u_CSAwallace_cska32_csa12_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa24_and1 = u_CSAwallace_cska32_csa18_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa24_or0 = u_CSAwallace_cska32_csa18_csa_component_fa24_and0 | u_CSAwallace_cska32_csa18_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa24_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa25_and0 = u_CSAwallace_cska32_csa11_csa_component_fa24_or0 & u_CSAwallace_cska32_csa12_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa25_and1 = u_CSAwallace_cska32_csa18_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa25_or0 = u_CSAwallace_cska32_csa18_csa_component_fa25_and0 | u_CSAwallace_cska32_csa18_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa25_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa26_and0 = u_CSAwallace_cska32_csa11_csa_component_fa25_or0 & u_CSAwallace_cska32_csa12_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa26_and1 = u_CSAwallace_cska32_csa18_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa26_or0 = u_CSAwallace_cska32_csa18_csa_component_fa26_and0 | u_CSAwallace_cska32_csa18_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa26_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa27_and0 = u_CSAwallace_cska32_csa11_csa_component_fa26_or0 & u_CSAwallace_cska32_csa12_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa27_and1 = u_CSAwallace_cska32_csa18_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa27_or0 = u_CSAwallace_cska32_csa18_csa_component_fa27_and0 | u_CSAwallace_cska32_csa18_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa27_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa28_and0 = u_CSAwallace_cska32_csa11_csa_component_fa27_or0 & u_CSAwallace_cska32_csa12_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa28_and1 = u_CSAwallace_cska32_csa18_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa28_or0 = u_CSAwallace_cska32_csa18_csa_component_fa28_and0 | u_CSAwallace_cska32_csa18_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa28_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa29_and0 = u_CSAwallace_cska32_csa11_csa_component_fa28_or0 & u_CSAwallace_cska32_csa12_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa29_and1 = u_CSAwallace_cska32_csa18_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa29_or0 = u_CSAwallace_cska32_csa18_csa_component_fa29_and0 | u_CSAwallace_cska32_csa18_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa29_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa30_and0 = u_CSAwallace_cska32_csa11_csa_component_fa29_or0 & u_CSAwallace_cska32_csa12_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa30_and1 = u_CSAwallace_cska32_csa18_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa30_or0 = u_CSAwallace_cska32_csa18_csa_component_fa30_and0 | u_CSAwallace_cska32_csa18_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa30_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa31_and0 = u_CSAwallace_cska32_csa11_csa_component_fa30_or0 & u_CSAwallace_cska32_csa12_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa31_and1 = u_CSAwallace_cska32_csa18_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa31_or0 = u_CSAwallace_cska32_csa18_csa_component_fa31_and0 | u_CSAwallace_cska32_csa18_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa31_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa32_and0 = u_CSAwallace_cska32_csa11_csa_component_fa31_or0 & u_CSAwallace_cska32_csa12_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa32_and1 = u_CSAwallace_cska32_csa18_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa32_or0 = u_CSAwallace_cska32_csa18_csa_component_fa32_and0 | u_CSAwallace_cska32_csa18_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa32_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa33_and0 = u_CSAwallace_cska32_csa11_csa_component_fa32_or0 & u_CSAwallace_cska32_csa12_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa33_and1 = u_CSAwallace_cska32_csa18_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa33_or0 = u_CSAwallace_cska32_csa18_csa_component_fa33_and0 | u_CSAwallace_cska32_csa18_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa33_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa34_and0 = u_CSAwallace_cska32_csa11_csa_component_fa33_or0 & u_CSAwallace_cska32_csa12_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa34_and1 = u_CSAwallace_cska32_csa18_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa34_or0 = u_CSAwallace_cska32_csa18_csa_component_fa34_and0 | u_CSAwallace_cska32_csa18_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa34_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa35_and0 = u_CSAwallace_cska32_csa11_csa_component_fa34_or0 & u_CSAwallace_cska32_csa12_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa35_and1 = u_CSAwallace_cska32_csa18_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa35_or0 = u_CSAwallace_cska32_csa18_csa_component_fa35_and0 | u_CSAwallace_cska32_csa18_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa35_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa36_and0 = u_CSAwallace_cska32_csa11_csa_component_fa35_or0 & u_CSAwallace_cska32_csa12_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa36_and1 = u_CSAwallace_cska32_csa18_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa36_or0 = u_CSAwallace_cska32_csa18_csa_component_fa36_and0 | u_CSAwallace_cska32_csa18_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa36_or0 ^ u_CSAwallace_cska32_csa12_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa37_and0 = u_CSAwallace_cska32_csa11_csa_component_fa36_or0 & u_CSAwallace_cska32_csa12_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa37_and1 = u_CSAwallace_cska32_csa18_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa37_or0 = u_CSAwallace_cska32_csa18_csa_component_fa37_and0 | u_CSAwallace_cska32_csa18_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa37_and1 ^ u_CSAwallace_cska32_csa12_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa38_and0 = u_CSAwallace_cska32_csa11_csa_component_fa37_and1 & u_CSAwallace_cska32_csa12_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa38_and1 = u_CSAwallace_cska32_csa18_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa38_or0 = u_CSAwallace_cska32_csa18_csa_component_fa38_and0 | u_CSAwallace_cska32_csa18_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa38_and1 ^ u_CSAwallace_cska32_csa12_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa39_and0 = u_CSAwallace_cska32_csa11_csa_component_fa38_and1 & u_CSAwallace_cska32_csa12_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa39_and1 = u_CSAwallace_cska32_csa18_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa39_or0 = u_CSAwallace_cska32_csa18_csa_component_fa39_and0 | u_CSAwallace_cska32_csa18_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa39_and1 ^ u_CSAwallace_cska32_csa12_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa40_and0 = u_CSAwallace_cska32_csa11_csa_component_fa39_and1 & u_CSAwallace_cska32_csa12_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa12_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa40_and1 = u_CSAwallace_cska32_csa18_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa12_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa40_or0 = u_CSAwallace_cska32_csa18_csa_component_fa40_and0 | u_CSAwallace_cska32_csa18_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa18_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa12_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa41_and1 = u_CSAwallace_cska32_csa12_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa12_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa12_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa12_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa42_and1 = u_CSAwallace_cska32_csa12_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa12_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa12_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa18_csa_component_fa43_and1 = u_CSAwallace_cska32_csa4_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa12_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa13_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa16_and0 = u_CSAwallace_cska32_csa13_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa13_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa17_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa17_and0 = u_CSAwallace_cska32_csa13_csa_component_fa17_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa18_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa18_and0 = u_CSAwallace_cska32_csa13_csa_component_fa18_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_and_0_18;
  assign u_CSAwallace_cska32_csa19_csa_component_fa18_and1 = u_CSAwallace_cska32_csa19_csa_component_fa18_xor0 & u_CSAwallace_cska32_and_0_18;
  assign u_CSAwallace_cska32_csa19_csa_component_fa18_or0 = u_CSAwallace_cska32_csa19_csa_component_fa18_and0 | u_CSAwallace_cska32_csa19_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa19_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa19_and0 = u_CSAwallace_cska32_csa13_csa_component_fa19_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa6_csa_component_fa19_xor0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa19_and1 = u_CSAwallace_cska32_csa19_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa6_csa_component_fa19_xor0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa19_or0 = u_CSAwallace_cska32_csa19_csa_component_fa19_and0 | u_CSAwallace_cska32_csa19_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa20_and0 = u_CSAwallace_cska32_csa13_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa20_xor0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa20_and1 = u_CSAwallace_cska32_csa19_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa20_xor0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa20_or0 = u_CSAwallace_cska32_csa19_csa_component_fa20_and0 | u_CSAwallace_cska32_csa19_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa21_and0 = u_CSAwallace_cska32_csa13_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa21_and1 = u_CSAwallace_cska32_csa19_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa21_or0 = u_CSAwallace_cska32_csa19_csa_component_fa21_and0 | u_CSAwallace_cska32_csa19_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa22_and0 = u_CSAwallace_cska32_csa13_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa22_and1 = u_CSAwallace_cska32_csa19_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa22_or0 = u_CSAwallace_cska32_csa19_csa_component_fa22_and0 | u_CSAwallace_cska32_csa19_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa23_and0 = u_CSAwallace_cska32_csa13_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa23_and1 = u_CSAwallace_cska32_csa19_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa23_or0 = u_CSAwallace_cska32_csa19_csa_component_fa23_and0 | u_CSAwallace_cska32_csa19_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa24_and0 = u_CSAwallace_cska32_csa13_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa24_and1 = u_CSAwallace_cska32_csa19_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa24_or0 = u_CSAwallace_cska32_csa19_csa_component_fa24_and0 | u_CSAwallace_cska32_csa19_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa25_and0 = u_CSAwallace_cska32_csa13_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa25_and1 = u_CSAwallace_cska32_csa19_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa25_or0 = u_CSAwallace_cska32_csa19_csa_component_fa25_and0 | u_CSAwallace_cska32_csa19_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa26_and0 = u_CSAwallace_cska32_csa13_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa26_and1 = u_CSAwallace_cska32_csa19_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa26_or0 = u_CSAwallace_cska32_csa19_csa_component_fa26_and0 | u_CSAwallace_cska32_csa19_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa27_and0 = u_CSAwallace_cska32_csa13_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa27_and1 = u_CSAwallace_cska32_csa19_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa27_or0 = u_CSAwallace_cska32_csa19_csa_component_fa27_and0 | u_CSAwallace_cska32_csa19_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa28_and0 = u_CSAwallace_cska32_csa13_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa28_and1 = u_CSAwallace_cska32_csa19_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa28_or0 = u_CSAwallace_cska32_csa19_csa_component_fa28_and0 | u_CSAwallace_cska32_csa19_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa29_and0 = u_CSAwallace_cska32_csa13_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa29_and1 = u_CSAwallace_cska32_csa19_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa29_or0 = u_CSAwallace_cska32_csa19_csa_component_fa29_and0 | u_CSAwallace_cska32_csa19_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa30_and0 = u_CSAwallace_cska32_csa13_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa30_and1 = u_CSAwallace_cska32_csa19_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa30_or0 = u_CSAwallace_cska32_csa19_csa_component_fa30_and0 | u_CSAwallace_cska32_csa19_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa31_and0 = u_CSAwallace_cska32_csa13_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa31_and1 = u_CSAwallace_cska32_csa19_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa31_or0 = u_CSAwallace_cska32_csa19_csa_component_fa31_and0 | u_CSAwallace_cska32_csa19_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa32_and0 = u_CSAwallace_cska32_csa13_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa32_and1 = u_CSAwallace_cska32_csa19_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa32_or0 = u_CSAwallace_cska32_csa19_csa_component_fa32_and0 | u_CSAwallace_cska32_csa19_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa33_and0 = u_CSAwallace_cska32_csa13_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa33_and1 = u_CSAwallace_cska32_csa19_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa33_or0 = u_CSAwallace_cska32_csa19_csa_component_fa33_and0 | u_CSAwallace_cska32_csa19_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa34_and0 = u_CSAwallace_cska32_csa13_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa34_and1 = u_CSAwallace_cska32_csa19_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa34_or0 = u_CSAwallace_cska32_csa19_csa_component_fa34_and0 | u_CSAwallace_cska32_csa19_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa35_and0 = u_CSAwallace_cska32_csa13_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa35_and1 = u_CSAwallace_cska32_csa19_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa35_or0 = u_CSAwallace_cska32_csa19_csa_component_fa35_and0 | u_CSAwallace_cska32_csa19_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa36_and0 = u_CSAwallace_cska32_csa13_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa36_and1 = u_CSAwallace_cska32_csa19_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa36_or0 = u_CSAwallace_cska32_csa19_csa_component_fa36_and0 | u_CSAwallace_cska32_csa19_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa37_and0 = u_CSAwallace_cska32_csa13_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa37_and1 = u_CSAwallace_cska32_csa19_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa37_or0 = u_CSAwallace_cska32_csa19_csa_component_fa37_and0 | u_CSAwallace_cska32_csa19_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa38_and0 = u_CSAwallace_cska32_csa13_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa38_and1 = u_CSAwallace_cska32_csa19_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa38_or0 = u_CSAwallace_cska32_csa19_csa_component_fa38_and0 | u_CSAwallace_cska32_csa19_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa39_and0 = u_CSAwallace_cska32_csa13_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa39_and1 = u_CSAwallace_cska32_csa19_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa39_or0 = u_CSAwallace_cska32_csa19_csa_component_fa39_and0 | u_CSAwallace_cska32_csa19_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa40_and0 = u_CSAwallace_cska32_csa13_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa40_and1 = u_CSAwallace_cska32_csa19_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa40_or0 = u_CSAwallace_cska32_csa19_csa_component_fa40_and0 | u_CSAwallace_cska32_csa19_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa41_and0 = u_CSAwallace_cska32_csa13_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa41_and1 = u_CSAwallace_cska32_csa19_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa41_or0 = u_CSAwallace_cska32_csa19_csa_component_fa41_and0 | u_CSAwallace_cska32_csa19_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa42_and0 = u_CSAwallace_cska32_csa13_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa42_and1 = u_CSAwallace_cska32_csa19_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa42_or0 = u_CSAwallace_cska32_csa19_csa_component_fa42_and0 | u_CSAwallace_cska32_csa19_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa43_and0 = u_CSAwallace_cska32_csa13_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa43_and1 = u_CSAwallace_cska32_csa19_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa43_or0 = u_CSAwallace_cska32_csa19_csa_component_fa43_and0 | u_CSAwallace_cska32_csa19_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa44_and0 = u_CSAwallace_cska32_csa13_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa44_and1 = u_CSAwallace_cska32_csa19_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa44_or0 = u_CSAwallace_cska32_csa19_csa_component_fa44_and0 | u_CSAwallace_cska32_csa19_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa45_and0 = u_CSAwallace_cska32_csa13_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa45_and1 = u_CSAwallace_cska32_csa19_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa45_or0 = u_CSAwallace_cska32_csa19_csa_component_fa45_and0 | u_CSAwallace_cska32_csa19_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa46_and0 = u_CSAwallace_cska32_csa13_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa19_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa46_and1 = u_CSAwallace_cska32_csa19_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa46_or0 = u_CSAwallace_cska32_csa19_csa_component_fa46_and0 | u_CSAwallace_cska32_csa19_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa47_and0 = u_CSAwallace_cska32_csa13_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa47_and1 = u_CSAwallace_cska32_csa19_csa_component_fa47_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa47_or0 = u_CSAwallace_cska32_csa19_csa_component_fa47_and0 | u_CSAwallace_cska32_csa19_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa13_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa13_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa48_and0 = u_CSAwallace_cska32_csa13_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa13_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_csa14_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa48_and1 = u_CSAwallace_cska32_csa19_csa_component_fa48_xor0 & u_CSAwallace_cska32_csa14_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa48_or0 = u_CSAwallace_cska32_csa19_csa_component_fa48_and0 | u_CSAwallace_cska32_csa19_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa13_csa_component_fa48_and1 ^ u_CSAwallace_cska32_csa14_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa19_csa_component_fa49_and1 = u_CSAwallace_cska32_csa13_csa_component_fa48_and1 & u_CSAwallace_cska32_csa14_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa22_or0 ^ u_CSAwallace_cska32_csa7_csa_component_fa22_and0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa23_and0 = u_CSAwallace_cska32_csa14_csa_component_fa22_or0 & u_CSAwallace_cska32_csa7_csa_component_fa22_and0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa23_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa24_xor0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa24_and0 = u_CSAwallace_cska32_csa14_csa_component_fa23_or0 & u_CSAwallace_cska32_csa15_csa_component_fa24_xor0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa24_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa25_xor0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa25_and0 = u_CSAwallace_cska32_csa14_csa_component_fa24_or0 & u_CSAwallace_cska32_csa15_csa_component_fa25_xor0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa25_and1 = u_CSAwallace_cska32_csa20_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa25_or0 = u_CSAwallace_cska32_csa20_csa_component_fa25_and0 | u_CSAwallace_cska32_csa20_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa25_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa26_and0 = u_CSAwallace_cska32_csa14_csa_component_fa25_or0 & u_CSAwallace_cska32_csa15_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa26_and1 = u_CSAwallace_cska32_csa20_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa26_or0 = u_CSAwallace_cska32_csa20_csa_component_fa26_and0 | u_CSAwallace_cska32_csa20_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa26_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa27_and0 = u_CSAwallace_cska32_csa14_csa_component_fa26_or0 & u_CSAwallace_cska32_csa15_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa27_and1 = u_CSAwallace_cska32_csa20_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa27_or0 = u_CSAwallace_cska32_csa20_csa_component_fa27_and0 | u_CSAwallace_cska32_csa20_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa27_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa28_and0 = u_CSAwallace_cska32_csa14_csa_component_fa27_or0 & u_CSAwallace_cska32_csa15_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa28_and1 = u_CSAwallace_cska32_csa20_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa28_or0 = u_CSAwallace_cska32_csa20_csa_component_fa28_and0 | u_CSAwallace_cska32_csa20_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa28_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa29_and0 = u_CSAwallace_cska32_csa14_csa_component_fa28_or0 & u_CSAwallace_cska32_csa15_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa29_and1 = u_CSAwallace_cska32_csa20_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa29_or0 = u_CSAwallace_cska32_csa20_csa_component_fa29_and0 | u_CSAwallace_cska32_csa20_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa29_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa30_and0 = u_CSAwallace_cska32_csa14_csa_component_fa29_or0 & u_CSAwallace_cska32_csa15_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa30_and1 = u_CSAwallace_cska32_csa20_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa30_or0 = u_CSAwallace_cska32_csa20_csa_component_fa30_and0 | u_CSAwallace_cska32_csa20_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa30_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa31_and0 = u_CSAwallace_cska32_csa14_csa_component_fa30_or0 & u_CSAwallace_cska32_csa15_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa31_and1 = u_CSAwallace_cska32_csa20_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa31_or0 = u_CSAwallace_cska32_csa20_csa_component_fa31_and0 | u_CSAwallace_cska32_csa20_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa31_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa32_and0 = u_CSAwallace_cska32_csa14_csa_component_fa31_or0 & u_CSAwallace_cska32_csa15_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa32_and1 = u_CSAwallace_cska32_csa20_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa32_or0 = u_CSAwallace_cska32_csa20_csa_component_fa32_and0 | u_CSAwallace_cska32_csa20_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa32_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa33_and0 = u_CSAwallace_cska32_csa14_csa_component_fa32_or0 & u_CSAwallace_cska32_csa15_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa33_and1 = u_CSAwallace_cska32_csa20_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa33_or0 = u_CSAwallace_cska32_csa20_csa_component_fa33_and0 | u_CSAwallace_cska32_csa20_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa33_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa34_and0 = u_CSAwallace_cska32_csa14_csa_component_fa33_or0 & u_CSAwallace_cska32_csa15_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa34_and1 = u_CSAwallace_cska32_csa20_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa34_or0 = u_CSAwallace_cska32_csa20_csa_component_fa34_and0 | u_CSAwallace_cska32_csa20_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa34_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa35_and0 = u_CSAwallace_cska32_csa14_csa_component_fa34_or0 & u_CSAwallace_cska32_csa15_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa35_and1 = u_CSAwallace_cska32_csa20_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa35_or0 = u_CSAwallace_cska32_csa20_csa_component_fa35_and0 | u_CSAwallace_cska32_csa20_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa35_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa36_and0 = u_CSAwallace_cska32_csa14_csa_component_fa35_or0 & u_CSAwallace_cska32_csa15_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa36_and1 = u_CSAwallace_cska32_csa20_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa36_or0 = u_CSAwallace_cska32_csa20_csa_component_fa36_and0 | u_CSAwallace_cska32_csa20_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa36_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa37_and0 = u_CSAwallace_cska32_csa14_csa_component_fa36_or0 & u_CSAwallace_cska32_csa15_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa37_and1 = u_CSAwallace_cska32_csa20_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa37_or0 = u_CSAwallace_cska32_csa20_csa_component_fa37_and0 | u_CSAwallace_cska32_csa20_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa37_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa38_and0 = u_CSAwallace_cska32_csa14_csa_component_fa37_or0 & u_CSAwallace_cska32_csa15_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa38_and1 = u_CSAwallace_cska32_csa20_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa38_or0 = u_CSAwallace_cska32_csa20_csa_component_fa38_and0 | u_CSAwallace_cska32_csa20_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa38_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa39_and0 = u_CSAwallace_cska32_csa14_csa_component_fa38_or0 & u_CSAwallace_cska32_csa15_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa39_and1 = u_CSAwallace_cska32_csa20_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa39_or0 = u_CSAwallace_cska32_csa20_csa_component_fa39_and0 | u_CSAwallace_cska32_csa20_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa39_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa40_and0 = u_CSAwallace_cska32_csa14_csa_component_fa39_or0 & u_CSAwallace_cska32_csa15_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa40_and1 = u_CSAwallace_cska32_csa20_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa40_or0 = u_CSAwallace_cska32_csa20_csa_component_fa40_and0 | u_CSAwallace_cska32_csa20_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa40_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa41_and0 = u_CSAwallace_cska32_csa14_csa_component_fa40_or0 & u_CSAwallace_cska32_csa15_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa41_and1 = u_CSAwallace_cska32_csa20_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa41_or0 = u_CSAwallace_cska32_csa20_csa_component_fa41_and0 | u_CSAwallace_cska32_csa20_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa41_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa42_and0 = u_CSAwallace_cska32_csa14_csa_component_fa41_or0 & u_CSAwallace_cska32_csa15_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa42_and1 = u_CSAwallace_cska32_csa20_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa42_or0 = u_CSAwallace_cska32_csa20_csa_component_fa42_and0 | u_CSAwallace_cska32_csa20_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa42_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa43_and0 = u_CSAwallace_cska32_csa14_csa_component_fa42_or0 & u_CSAwallace_cska32_csa15_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa43_and1 = u_CSAwallace_cska32_csa20_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa43_or0 = u_CSAwallace_cska32_csa20_csa_component_fa43_and0 | u_CSAwallace_cska32_csa20_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa43_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa44_and0 = u_CSAwallace_cska32_csa14_csa_component_fa43_or0 & u_CSAwallace_cska32_csa15_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa44_and1 = u_CSAwallace_cska32_csa20_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa44_or0 = u_CSAwallace_cska32_csa20_csa_component_fa44_and0 | u_CSAwallace_cska32_csa20_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa44_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa45_and0 = u_CSAwallace_cska32_csa14_csa_component_fa44_or0 & u_CSAwallace_cska32_csa15_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa45_and1 = u_CSAwallace_cska32_csa20_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa45_or0 = u_CSAwallace_cska32_csa20_csa_component_fa45_and0 | u_CSAwallace_cska32_csa20_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa45_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa46_and0 = u_CSAwallace_cska32_csa14_csa_component_fa45_or0 & u_CSAwallace_cska32_csa15_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa46_and1 = u_CSAwallace_cska32_csa20_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa46_or0 = u_CSAwallace_cska32_csa20_csa_component_fa46_and0 | u_CSAwallace_cska32_csa20_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa46_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa47_and0 = u_CSAwallace_cska32_csa14_csa_component_fa46_or0 & u_CSAwallace_cska32_csa15_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa47_and1 = u_CSAwallace_cska32_csa20_csa_component_fa47_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa47_or0 = u_CSAwallace_cska32_csa20_csa_component_fa47_and0 | u_CSAwallace_cska32_csa20_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa47_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa48_and0 = u_CSAwallace_cska32_csa14_csa_component_fa47_or0 & u_CSAwallace_cska32_csa15_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa48_and1 = u_CSAwallace_cska32_csa20_csa_component_fa48_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa48_or0 = u_CSAwallace_cska32_csa20_csa_component_fa48_and0 | u_CSAwallace_cska32_csa20_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa48_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa49_and0 = u_CSAwallace_cska32_csa14_csa_component_fa48_or0 & u_CSAwallace_cska32_csa15_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa49_and1 = u_CSAwallace_cska32_csa20_csa_component_fa49_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa49_or0 = u_CSAwallace_cska32_csa20_csa_component_fa49_and0 | u_CSAwallace_cska32_csa20_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa49_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa50_and0 = u_CSAwallace_cska32_csa14_csa_component_fa49_or0 & u_CSAwallace_cska32_csa15_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa50_and1 = u_CSAwallace_cska32_csa20_csa_component_fa50_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa50_or0 = u_CSAwallace_cska32_csa20_csa_component_fa50_and0 | u_CSAwallace_cska32_csa20_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa51_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa50_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa51_and0 = u_CSAwallace_cska32_csa14_csa_component_fa50_or0 & u_CSAwallace_cska32_csa15_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa51_and1 = u_CSAwallace_cska32_csa20_csa_component_fa51_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa51_or0 = u_CSAwallace_cska32_csa20_csa_component_fa51_and0 | u_CSAwallace_cska32_csa20_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa52_xor0 = u_CSAwallace_cska32_csa14_csa_component_fa51_or0 ^ u_CSAwallace_cska32_csa15_csa_component_fa52_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa52_and0 = u_CSAwallace_cska32_csa14_csa_component_fa51_or0 & u_CSAwallace_cska32_csa15_csa_component_fa52_xor1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa20_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_csa15_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa52_and1 = u_CSAwallace_cska32_csa20_csa_component_fa52_xor0 & u_CSAwallace_cska32_csa15_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa52_or0 = u_CSAwallace_cska32_csa20_csa_component_fa52_and0 | u_CSAwallace_cska32_csa20_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa15_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa53_and1 = u_CSAwallace_cska32_csa15_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa15_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa15_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa54_and1 = u_CSAwallace_cska32_csa15_csa_component_fa54_xor1 & u_CSAwallace_cska32_csa15_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa15_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa55_and1 = u_CSAwallace_cska32_csa15_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa15_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa20_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa15_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa56_and1 = u_CSAwallace_cska32_csa15_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa15_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa57_xor1 = u_CSAwallace_cska32_csa15_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa15_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa20_csa_component_fa57_and1 = u_CSAwallace_cska32_csa15_csa_component_fa57_xor1 & u_CSAwallace_cska32_csa15_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa29_and0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa30_and0 = u_CSAwallace_cska32_csa16_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa29_and0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa31_and0 = u_CSAwallace_cska32_csa16_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_and_0_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa31_and1 = u_CSAwallace_cska32_csa21_csa_component_fa31_xor0 & u_CSAwallace_cska32_and_0_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa31_or0 = u_CSAwallace_cska32_csa21_csa_component_fa31_and0 | u_CSAwallace_cska32_csa21_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa32_and0 = u_CSAwallace_cska32_csa16_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_and_1_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa32_and1 = u_CSAwallace_cska32_csa21_csa_component_fa32_xor0 & u_CSAwallace_cska32_and_1_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa32_or0 = u_CSAwallace_cska32_csa21_csa_component_fa32_and0 | u_CSAwallace_cska32_csa21_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa33_and0 = u_CSAwallace_cska32_csa16_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_and_2_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa33_and1 = u_CSAwallace_cska32_csa21_csa_component_fa33_xor0 & u_CSAwallace_cska32_and_2_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa33_or0 = u_CSAwallace_cska32_csa21_csa_component_fa33_and0 | u_CSAwallace_cska32_csa21_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa34_and0 = u_CSAwallace_cska32_csa16_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_and_3_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa34_and1 = u_CSAwallace_cska32_csa21_csa_component_fa34_xor0 & u_CSAwallace_cska32_and_3_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa34_or0 = u_CSAwallace_cska32_csa21_csa_component_fa34_and0 | u_CSAwallace_cska32_csa21_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa35_and0 = u_CSAwallace_cska32_csa16_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_and_4_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa35_and1 = u_CSAwallace_cska32_csa21_csa_component_fa35_xor0 & u_CSAwallace_cska32_and_4_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa35_or0 = u_CSAwallace_cska32_csa21_csa_component_fa35_and0 | u_CSAwallace_cska32_csa21_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa36_and0 = u_CSAwallace_cska32_csa16_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_and_5_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa36_and1 = u_CSAwallace_cska32_csa21_csa_component_fa36_xor0 & u_CSAwallace_cska32_and_5_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa36_or0 = u_CSAwallace_cska32_csa21_csa_component_fa36_and0 | u_CSAwallace_cska32_csa21_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa37_and0 = u_CSAwallace_cska32_csa16_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_and_6_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa37_and1 = u_CSAwallace_cska32_csa21_csa_component_fa37_xor0 & u_CSAwallace_cska32_and_6_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa37_or0 = u_CSAwallace_cska32_csa21_csa_component_fa37_and0 | u_CSAwallace_cska32_csa21_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa38_and0 = u_CSAwallace_cska32_csa16_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_and_7_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa38_and1 = u_CSAwallace_cska32_csa21_csa_component_fa38_xor0 & u_CSAwallace_cska32_and_7_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa38_or0 = u_CSAwallace_cska32_csa21_csa_component_fa38_and0 | u_CSAwallace_cska32_csa21_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa39_and0 = u_CSAwallace_cska32_csa16_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_and_8_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa39_and1 = u_CSAwallace_cska32_csa21_csa_component_fa39_xor0 & u_CSAwallace_cska32_and_8_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa39_or0 = u_CSAwallace_cska32_csa21_csa_component_fa39_and0 | u_CSAwallace_cska32_csa21_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa40_and0 = u_CSAwallace_cska32_csa16_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_and_9_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa40_and1 = u_CSAwallace_cska32_csa21_csa_component_fa40_xor0 & u_CSAwallace_cska32_and_9_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa40_or0 = u_CSAwallace_cska32_csa21_csa_component_fa40_and0 | u_CSAwallace_cska32_csa21_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa41_and0 = u_CSAwallace_cska32_csa16_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_and_10_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa41_and1 = u_CSAwallace_cska32_csa21_csa_component_fa41_xor0 & u_CSAwallace_cska32_and_10_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa41_or0 = u_CSAwallace_cska32_csa21_csa_component_fa41_and0 | u_CSAwallace_cska32_csa21_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa42_and0 = u_CSAwallace_cska32_csa16_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_and_11_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa42_and1 = u_CSAwallace_cska32_csa21_csa_component_fa42_xor0 & u_CSAwallace_cska32_and_11_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa42_or0 = u_CSAwallace_cska32_csa21_csa_component_fa42_and0 | u_CSAwallace_cska32_csa21_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa43_and0 = u_CSAwallace_cska32_csa16_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_and_12_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa43_and1 = u_CSAwallace_cska32_csa21_csa_component_fa43_xor0 & u_CSAwallace_cska32_and_12_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa43_or0 = u_CSAwallace_cska32_csa21_csa_component_fa43_and0 | u_CSAwallace_cska32_csa21_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa44_and0 = u_CSAwallace_cska32_csa16_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_and_13_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa44_and1 = u_CSAwallace_cska32_csa21_csa_component_fa44_xor0 & u_CSAwallace_cska32_and_13_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa44_or0 = u_CSAwallace_cska32_csa21_csa_component_fa44_and0 | u_CSAwallace_cska32_csa21_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa45_and0 = u_CSAwallace_cska32_csa16_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_and_14_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa45_and1 = u_CSAwallace_cska32_csa21_csa_component_fa45_xor0 & u_CSAwallace_cska32_and_14_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa45_or0 = u_CSAwallace_cska32_csa21_csa_component_fa45_and0 | u_CSAwallace_cska32_csa21_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa46_and0 = u_CSAwallace_cska32_csa16_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_and_15_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa46_and1 = u_CSAwallace_cska32_csa21_csa_component_fa46_xor0 & u_CSAwallace_cska32_and_15_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa46_or0 = u_CSAwallace_cska32_csa21_csa_component_fa46_and0 | u_CSAwallace_cska32_csa21_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa47_and0 = u_CSAwallace_cska32_csa16_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_and_16_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa47_and1 = u_CSAwallace_cska32_csa21_csa_component_fa47_xor0 & u_CSAwallace_cska32_and_16_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa47_or0 = u_CSAwallace_cska32_csa21_csa_component_fa47_and0 | u_CSAwallace_cska32_csa21_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa48_and0 = u_CSAwallace_cska32_csa16_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_and_17_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa48_and1 = u_CSAwallace_cska32_csa21_csa_component_fa48_xor0 & u_CSAwallace_cska32_and_17_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa48_or0 = u_CSAwallace_cska32_csa21_csa_component_fa48_and0 | u_CSAwallace_cska32_csa21_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa49_and0 = u_CSAwallace_cska32_csa16_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_and_18_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa49_and1 = u_CSAwallace_cska32_csa21_csa_component_fa49_xor0 & u_CSAwallace_cska32_and_18_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa49_or0 = u_CSAwallace_cska32_csa21_csa_component_fa49_and0 | u_CSAwallace_cska32_csa21_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa50_and0 = u_CSAwallace_cska32_csa16_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_and_19_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa50_and1 = u_CSAwallace_cska32_csa21_csa_component_fa50_xor0 & u_CSAwallace_cska32_and_19_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa50_or0 = u_CSAwallace_cska32_csa21_csa_component_fa50_and0 | u_CSAwallace_cska32_csa21_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa51_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa51_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa51_and0 = u_CSAwallace_cska32_csa16_csa_component_fa51_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_and_20_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa51_and1 = u_CSAwallace_cska32_csa21_csa_component_fa51_xor0 & u_CSAwallace_cska32_and_20_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa51_or0 = u_CSAwallace_cska32_csa21_csa_component_fa51_and0 | u_CSAwallace_cska32_csa21_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa52_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa52_and0 = u_CSAwallace_cska32_csa16_csa_component_fa52_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_and_21_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa52_and1 = u_CSAwallace_cska32_csa21_csa_component_fa52_xor0 & u_CSAwallace_cska32_and_21_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa52_or0 = u_CSAwallace_cska32_csa21_csa_component_fa52_and0 | u_CSAwallace_cska32_csa21_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa53_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa53_and0 = u_CSAwallace_cska32_csa16_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa53_xor0 ^ u_CSAwallace_cska32_and_22_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa53_and1 = u_CSAwallace_cska32_csa21_csa_component_fa53_xor0 & u_CSAwallace_cska32_and_22_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa53_or0 = u_CSAwallace_cska32_csa21_csa_component_fa53_and0 | u_CSAwallace_cska32_csa21_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa54_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa54_and0 = u_CSAwallace_cska32_csa16_csa_component_fa54_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa54_xor0 ^ u_CSAwallace_cska32_and_23_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa54_and1 = u_CSAwallace_cska32_csa21_csa_component_fa54_xor0 & u_CSAwallace_cska32_and_23_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa54_or0 = u_CSAwallace_cska32_csa21_csa_component_fa54_and0 | u_CSAwallace_cska32_csa21_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa55_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa55_and0 = u_CSAwallace_cska32_csa16_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa55_xor0 ^ u_CSAwallace_cska32_and_24_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa55_and1 = u_CSAwallace_cska32_csa21_csa_component_fa55_xor0 & u_CSAwallace_cska32_and_24_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa55_or0 = u_CSAwallace_cska32_csa21_csa_component_fa55_and0 | u_CSAwallace_cska32_csa21_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa56_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa56_and0 = u_CSAwallace_cska32_csa16_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa56_xor0 ^ u_CSAwallace_cska32_and_25_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa56_and1 = u_CSAwallace_cska32_csa21_csa_component_fa56_xor0 & u_CSAwallace_cska32_and_25_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa56_or0 = u_CSAwallace_cska32_csa21_csa_component_fa56_and0 | u_CSAwallace_cska32_csa21_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa57_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa57_and0 = u_CSAwallace_cska32_csa16_csa_component_fa57_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa57_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa57_xor0 ^ u_CSAwallace_cska32_and_26_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa57_and1 = u_CSAwallace_cska32_csa21_csa_component_fa57_xor0 & u_CSAwallace_cska32_and_26_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa57_or0 = u_CSAwallace_cska32_csa21_csa_component_fa57_and0 | u_CSAwallace_cska32_csa21_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa58_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa58_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa58_and0 = u_CSAwallace_cska32_csa16_csa_component_fa58_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa58_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa58_xor0 ^ u_CSAwallace_cska32_and_27_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa58_and1 = u_CSAwallace_cska32_csa21_csa_component_fa58_xor0 & u_CSAwallace_cska32_and_27_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa58_or0 = u_CSAwallace_cska32_csa21_csa_component_fa58_and0 | u_CSAwallace_cska32_csa21_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa59_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa59_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa59_and0 = u_CSAwallace_cska32_csa16_csa_component_fa59_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa59_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa59_xor0 ^ u_CSAwallace_cska32_and_28_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa59_and1 = u_CSAwallace_cska32_csa21_csa_component_fa59_xor0 & u_CSAwallace_cska32_and_28_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa59_or0 = u_CSAwallace_cska32_csa21_csa_component_fa59_and0 | u_CSAwallace_cska32_csa21_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa60_xor0 = u_CSAwallace_cska32_csa16_csa_component_fa60_xor1 ^ u_CSAwallace_cska32_csa16_csa_component_fa59_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa60_and0 = u_CSAwallace_cska32_csa16_csa_component_fa60_xor1 & u_CSAwallace_cska32_csa16_csa_component_fa59_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa60_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa60_xor0 ^ u_CSAwallace_cska32_and_29_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa60_and1 = u_CSAwallace_cska32_csa21_csa_component_fa60_xor0 & u_CSAwallace_cska32_and_29_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa60_or0 = u_CSAwallace_cska32_csa21_csa_component_fa60_and0 | u_CSAwallace_cska32_csa21_csa_component_fa60_and1;
  assign u_CSAwallace_cska32_csa21_csa_component_fa61_xor0 = u_CSAwallace_cska32_and_31_30 ^ u_CSAwallace_cska32_csa16_csa_component_fa60_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa61_and0 = u_CSAwallace_cska32_and_31_30 & u_CSAwallace_cska32_csa16_csa_component_fa60_or0;
  assign u_CSAwallace_cska32_csa21_csa_component_fa61_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa61_xor0 ^ u_CSAwallace_cska32_and_30_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa61_and1 = u_CSAwallace_cska32_csa21_csa_component_fa61_xor0 & u_CSAwallace_cska32_and_30_31;
  assign u_CSAwallace_cska32_csa21_csa_component_fa61_or0 = u_CSAwallace_cska32_csa21_csa_component_fa61_and0 | u_CSAwallace_cska32_csa21_csa_component_fa61_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa4_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa4_xor0 ^ u_CSAwallace_cska32_csa17_csa_component_fa3_and0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa4_and0 = u_CSAwallace_cska32_csa17_csa_component_fa4_xor0 & u_CSAwallace_cska32_csa17_csa_component_fa3_and0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa5_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa5_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa4_and0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa5_and0 = u_CSAwallace_cska32_csa17_csa_component_fa5_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa4_and0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa6_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa6_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa5_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa6_and0 = u_CSAwallace_cska32_csa17_csa_component_fa6_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa5_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa7_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa7_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa6_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa7_and0 = u_CSAwallace_cska32_csa17_csa_component_fa7_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa6_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa7_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa7_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa6_and0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa7_and1 = u_CSAwallace_cska32_csa22_csa_component_fa7_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa6_and0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa7_or0 = u_CSAwallace_cska32_csa22_csa_component_fa7_and0 | u_CSAwallace_cska32_csa22_csa_component_fa7_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa8_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa8_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa7_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa8_and0 = u_CSAwallace_cska32_csa17_csa_component_fa8_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa7_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa8_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_csa11_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa8_and1 = u_CSAwallace_cska32_csa22_csa_component_fa8_xor0 & u_CSAwallace_cska32_csa11_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa8_or0 = u_CSAwallace_cska32_csa22_csa_component_fa8_and0 | u_CSAwallace_cska32_csa22_csa_component_fa8_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa9_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa9_and0 = u_CSAwallace_cska32_csa17_csa_component_fa9_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa9_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa9_xor0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa9_and1 = u_CSAwallace_cska32_csa22_csa_component_fa9_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa9_xor0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa9_or0 = u_CSAwallace_cska32_csa22_csa_component_fa9_and0 | u_CSAwallace_cska32_csa22_csa_component_fa9_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa10_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa10_and0 = u_CSAwallace_cska32_csa17_csa_component_fa10_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa10_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa10_xor0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa10_and1 = u_CSAwallace_cska32_csa22_csa_component_fa10_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa10_xor0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa10_or0 = u_CSAwallace_cska32_csa22_csa_component_fa10_and0 | u_CSAwallace_cska32_csa22_csa_component_fa10_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa11_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa11_and0 = u_CSAwallace_cska32_csa17_csa_component_fa11_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa11_xor0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa11_and1 = u_CSAwallace_cska32_csa22_csa_component_fa11_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa11_xor0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa11_or0 = u_CSAwallace_cska32_csa22_csa_component_fa11_and0 | u_CSAwallace_cska32_csa22_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa12_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa12_and0 = u_CSAwallace_cska32_csa17_csa_component_fa12_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa12_and1 = u_CSAwallace_cska32_csa22_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa12_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa12_or0 = u_CSAwallace_cska32_csa22_csa_component_fa12_and0 | u_CSAwallace_cska32_csa22_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa13_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa13_and0 = u_CSAwallace_cska32_csa17_csa_component_fa13_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa13_and1 = u_CSAwallace_cska32_csa22_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa13_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa13_or0 = u_CSAwallace_cska32_csa22_csa_component_fa13_and0 | u_CSAwallace_cska32_csa22_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa14_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa14_and0 = u_CSAwallace_cska32_csa17_csa_component_fa14_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa14_and1 = u_CSAwallace_cska32_csa22_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa14_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa14_or0 = u_CSAwallace_cska32_csa22_csa_component_fa14_and0 | u_CSAwallace_cska32_csa22_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa15_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa15_and0 = u_CSAwallace_cska32_csa17_csa_component_fa15_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa15_and1 = u_CSAwallace_cska32_csa22_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa15_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa15_or0 = u_CSAwallace_cska32_csa22_csa_component_fa15_and0 | u_CSAwallace_cska32_csa22_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa16_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa16_and0 = u_CSAwallace_cska32_csa17_csa_component_fa16_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa16_and1 = u_CSAwallace_cska32_csa22_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa16_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa16_or0 = u_CSAwallace_cska32_csa22_csa_component_fa16_and0 | u_CSAwallace_cska32_csa22_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa17_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa17_and0 = u_CSAwallace_cska32_csa17_csa_component_fa17_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa17_and1 = u_CSAwallace_cska32_csa22_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa17_or0 = u_CSAwallace_cska32_csa22_csa_component_fa17_and0 | u_CSAwallace_cska32_csa22_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa18_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa18_and0 = u_CSAwallace_cska32_csa17_csa_component_fa18_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa18_and1 = u_CSAwallace_cska32_csa22_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa18_or0 = u_CSAwallace_cska32_csa22_csa_component_fa18_and0 | u_CSAwallace_cska32_csa22_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa19_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa19_and0 = u_CSAwallace_cska32_csa17_csa_component_fa19_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa19_and1 = u_CSAwallace_cska32_csa22_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa19_or0 = u_CSAwallace_cska32_csa22_csa_component_fa19_and0 | u_CSAwallace_cska32_csa22_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa20_and0 = u_CSAwallace_cska32_csa17_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa20_and1 = u_CSAwallace_cska32_csa22_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa20_or0 = u_CSAwallace_cska32_csa22_csa_component_fa20_and0 | u_CSAwallace_cska32_csa22_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa21_and0 = u_CSAwallace_cska32_csa17_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa21_and1 = u_CSAwallace_cska32_csa22_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa21_or0 = u_CSAwallace_cska32_csa22_csa_component_fa21_and0 | u_CSAwallace_cska32_csa22_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa22_and0 = u_CSAwallace_cska32_csa17_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa22_and1 = u_CSAwallace_cska32_csa22_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa22_or0 = u_CSAwallace_cska32_csa22_csa_component_fa22_and0 | u_CSAwallace_cska32_csa22_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa23_and0 = u_CSAwallace_cska32_csa17_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa23_and1 = u_CSAwallace_cska32_csa22_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa23_or0 = u_CSAwallace_cska32_csa22_csa_component_fa23_and0 | u_CSAwallace_cska32_csa22_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa24_and0 = u_CSAwallace_cska32_csa17_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa24_and1 = u_CSAwallace_cska32_csa22_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa24_or0 = u_CSAwallace_cska32_csa22_csa_component_fa24_and0 | u_CSAwallace_cska32_csa22_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa25_and0 = u_CSAwallace_cska32_csa17_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa25_and1 = u_CSAwallace_cska32_csa22_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa25_or0 = u_CSAwallace_cska32_csa22_csa_component_fa25_and0 | u_CSAwallace_cska32_csa22_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa26_and0 = u_CSAwallace_cska32_csa17_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa26_and1 = u_CSAwallace_cska32_csa22_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa26_or0 = u_CSAwallace_cska32_csa22_csa_component_fa26_and0 | u_CSAwallace_cska32_csa22_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa27_and0 = u_CSAwallace_cska32_csa17_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa27_and1 = u_CSAwallace_cska32_csa22_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa27_or0 = u_CSAwallace_cska32_csa22_csa_component_fa27_and0 | u_CSAwallace_cska32_csa22_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa28_and0 = u_CSAwallace_cska32_csa17_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa28_and1 = u_CSAwallace_cska32_csa22_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa28_or0 = u_CSAwallace_cska32_csa22_csa_component_fa28_and0 | u_CSAwallace_cska32_csa22_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa29_and0 = u_CSAwallace_cska32_csa17_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa29_and1 = u_CSAwallace_cska32_csa22_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa29_or0 = u_CSAwallace_cska32_csa22_csa_component_fa29_and0 | u_CSAwallace_cska32_csa22_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa30_and0 = u_CSAwallace_cska32_csa17_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa30_and1 = u_CSAwallace_cska32_csa22_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa30_or0 = u_CSAwallace_cska32_csa22_csa_component_fa30_and0 | u_CSAwallace_cska32_csa22_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa31_and0 = u_CSAwallace_cska32_csa17_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa31_and1 = u_CSAwallace_cska32_csa22_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa31_or0 = u_CSAwallace_cska32_csa22_csa_component_fa31_and0 | u_CSAwallace_cska32_csa22_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa32_and0 = u_CSAwallace_cska32_csa17_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa32_and1 = u_CSAwallace_cska32_csa22_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa32_or0 = u_CSAwallace_cska32_csa22_csa_component_fa32_and0 | u_CSAwallace_cska32_csa22_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa33_and0 = u_CSAwallace_cska32_csa17_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa33_and1 = u_CSAwallace_cska32_csa22_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa33_or0 = u_CSAwallace_cska32_csa22_csa_component_fa33_and0 | u_CSAwallace_cska32_csa22_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa34_and0 = u_CSAwallace_cska32_csa17_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa34_and1 = u_CSAwallace_cska32_csa22_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa34_or0 = u_CSAwallace_cska32_csa22_csa_component_fa34_and0 | u_CSAwallace_cska32_csa22_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa35_and0 = u_CSAwallace_cska32_csa17_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa22_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa35_and1 = u_CSAwallace_cska32_csa22_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa35_or0 = u_CSAwallace_cska32_csa22_csa_component_fa35_and0 | u_CSAwallace_cska32_csa22_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa17_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa36_and0 = u_CSAwallace_cska32_csa17_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa36_and1 = u_CSAwallace_cska32_csa22_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa36_or0 = u_CSAwallace_cska32_csa22_csa_component_fa36_and0 | u_CSAwallace_cska32_csa22_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa11_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa17_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa37_and0 = u_CSAwallace_cska32_csa11_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa17_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa22_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa37_and1 = u_CSAwallace_cska32_csa22_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa37_or0 = u_CSAwallace_cska32_csa22_csa_component_fa37_and0 | u_CSAwallace_cska32_csa22_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa18_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa38_and1 = u_CSAwallace_cska32_csa11_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa18_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa11_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa18_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa22_csa_component_fa39_and1 = u_CSAwallace_cska32_csa11_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa18_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa13_or0 ^ u_CSAwallace_cska32_csa4_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa14_and0 = u_CSAwallace_cska32_csa18_csa_component_fa13_or0 & u_CSAwallace_cska32_csa4_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa14_or0 ^ u_CSAwallace_cska32_csa13_csa_component_fa15_xor0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa15_and0 = u_CSAwallace_cska32_csa18_csa_component_fa14_or0 & u_CSAwallace_cska32_csa13_csa_component_fa15_xor0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa15_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa16_xor0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa16_and0 = u_CSAwallace_cska32_csa18_csa_component_fa15_or0 & u_CSAwallace_cska32_csa19_csa_component_fa16_xor0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa16_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa17_xor0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa17_and0 = u_CSAwallace_cska32_csa18_csa_component_fa16_or0 & u_CSAwallace_cska32_csa19_csa_component_fa17_xor0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa17_and1 = u_CSAwallace_cska32_csa23_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa17_or0 = u_CSAwallace_cska32_csa23_csa_component_fa17_and0 | u_CSAwallace_cska32_csa23_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa17_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa18_and0 = u_CSAwallace_cska32_csa18_csa_component_fa17_or0 & u_CSAwallace_cska32_csa19_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa17_and0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa18_and1 = u_CSAwallace_cska32_csa23_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa17_and0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa18_or0 = u_CSAwallace_cska32_csa23_csa_component_fa18_and0 | u_CSAwallace_cska32_csa23_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa18_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa19_and0 = u_CSAwallace_cska32_csa18_csa_component_fa18_or0 & u_CSAwallace_cska32_csa19_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa19_and1 = u_CSAwallace_cska32_csa23_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa19_or0 = u_CSAwallace_cska32_csa23_csa_component_fa19_and0 | u_CSAwallace_cska32_csa23_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa19_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa20_and0 = u_CSAwallace_cska32_csa18_csa_component_fa19_or0 & u_CSAwallace_cska32_csa19_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa20_and1 = u_CSAwallace_cska32_csa23_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa20_or0 = u_CSAwallace_cska32_csa23_csa_component_fa20_and0 | u_CSAwallace_cska32_csa23_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa20_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa21_and0 = u_CSAwallace_cska32_csa18_csa_component_fa20_or0 & u_CSAwallace_cska32_csa19_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa21_and1 = u_CSAwallace_cska32_csa23_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa21_or0 = u_CSAwallace_cska32_csa23_csa_component_fa21_and0 | u_CSAwallace_cska32_csa23_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa21_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa22_and0 = u_CSAwallace_cska32_csa18_csa_component_fa21_or0 & u_CSAwallace_cska32_csa19_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa22_and1 = u_CSAwallace_cska32_csa23_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa22_or0 = u_CSAwallace_cska32_csa23_csa_component_fa22_and0 | u_CSAwallace_cska32_csa23_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa22_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa23_and0 = u_CSAwallace_cska32_csa18_csa_component_fa22_or0 & u_CSAwallace_cska32_csa19_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa23_and1 = u_CSAwallace_cska32_csa23_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa23_or0 = u_CSAwallace_cska32_csa23_csa_component_fa23_and0 | u_CSAwallace_cska32_csa23_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa23_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa24_and0 = u_CSAwallace_cska32_csa18_csa_component_fa23_or0 & u_CSAwallace_cska32_csa19_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa24_and1 = u_CSAwallace_cska32_csa23_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa24_or0 = u_CSAwallace_cska32_csa23_csa_component_fa24_and0 | u_CSAwallace_cska32_csa23_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa24_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa25_and0 = u_CSAwallace_cska32_csa18_csa_component_fa24_or0 & u_CSAwallace_cska32_csa19_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa25_and1 = u_CSAwallace_cska32_csa23_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa25_or0 = u_CSAwallace_cska32_csa23_csa_component_fa25_and0 | u_CSAwallace_cska32_csa23_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa25_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa26_and0 = u_CSAwallace_cska32_csa18_csa_component_fa25_or0 & u_CSAwallace_cska32_csa19_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa26_and1 = u_CSAwallace_cska32_csa23_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa26_or0 = u_CSAwallace_cska32_csa23_csa_component_fa26_and0 | u_CSAwallace_cska32_csa23_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa26_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa27_and0 = u_CSAwallace_cska32_csa18_csa_component_fa26_or0 & u_CSAwallace_cska32_csa19_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa27_and1 = u_CSAwallace_cska32_csa23_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa27_or0 = u_CSAwallace_cska32_csa23_csa_component_fa27_and0 | u_CSAwallace_cska32_csa23_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa27_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa28_and0 = u_CSAwallace_cska32_csa18_csa_component_fa27_or0 & u_CSAwallace_cska32_csa19_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa28_and1 = u_CSAwallace_cska32_csa23_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa28_or0 = u_CSAwallace_cska32_csa23_csa_component_fa28_and0 | u_CSAwallace_cska32_csa23_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa28_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa29_and0 = u_CSAwallace_cska32_csa18_csa_component_fa28_or0 & u_CSAwallace_cska32_csa19_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa29_and1 = u_CSAwallace_cska32_csa23_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa29_or0 = u_CSAwallace_cska32_csa23_csa_component_fa29_and0 | u_CSAwallace_cska32_csa23_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa29_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa30_and0 = u_CSAwallace_cska32_csa18_csa_component_fa29_or0 & u_CSAwallace_cska32_csa19_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa30_and1 = u_CSAwallace_cska32_csa23_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa30_or0 = u_CSAwallace_cska32_csa23_csa_component_fa30_and0 | u_CSAwallace_cska32_csa23_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa30_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa31_and0 = u_CSAwallace_cska32_csa18_csa_component_fa30_or0 & u_CSAwallace_cska32_csa19_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa31_and1 = u_CSAwallace_cska32_csa23_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa31_or0 = u_CSAwallace_cska32_csa23_csa_component_fa31_and0 | u_CSAwallace_cska32_csa23_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa31_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa32_and0 = u_CSAwallace_cska32_csa18_csa_component_fa31_or0 & u_CSAwallace_cska32_csa19_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa32_and1 = u_CSAwallace_cska32_csa23_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa32_or0 = u_CSAwallace_cska32_csa23_csa_component_fa32_and0 | u_CSAwallace_cska32_csa23_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa32_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa33_and0 = u_CSAwallace_cska32_csa18_csa_component_fa32_or0 & u_CSAwallace_cska32_csa19_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa33_and1 = u_CSAwallace_cska32_csa23_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa33_or0 = u_CSAwallace_cska32_csa23_csa_component_fa33_and0 | u_CSAwallace_cska32_csa23_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa33_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa34_and0 = u_CSAwallace_cska32_csa18_csa_component_fa33_or0 & u_CSAwallace_cska32_csa19_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa34_and1 = u_CSAwallace_cska32_csa23_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa34_or0 = u_CSAwallace_cska32_csa23_csa_component_fa34_and0 | u_CSAwallace_cska32_csa23_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa34_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa35_and0 = u_CSAwallace_cska32_csa18_csa_component_fa34_or0 & u_CSAwallace_cska32_csa19_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa35_and1 = u_CSAwallace_cska32_csa23_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa35_or0 = u_CSAwallace_cska32_csa23_csa_component_fa35_and0 | u_CSAwallace_cska32_csa23_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa35_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa36_and0 = u_CSAwallace_cska32_csa18_csa_component_fa35_or0 & u_CSAwallace_cska32_csa19_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa36_and1 = u_CSAwallace_cska32_csa23_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa36_or0 = u_CSAwallace_cska32_csa23_csa_component_fa36_and0 | u_CSAwallace_cska32_csa23_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa36_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa37_and0 = u_CSAwallace_cska32_csa18_csa_component_fa36_or0 & u_CSAwallace_cska32_csa19_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa37_and1 = u_CSAwallace_cska32_csa23_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa37_or0 = u_CSAwallace_cska32_csa23_csa_component_fa37_and0 | u_CSAwallace_cska32_csa23_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa37_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa38_and0 = u_CSAwallace_cska32_csa18_csa_component_fa37_or0 & u_CSAwallace_cska32_csa19_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa38_and1 = u_CSAwallace_cska32_csa23_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa38_or0 = u_CSAwallace_cska32_csa23_csa_component_fa38_and0 | u_CSAwallace_cska32_csa23_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa38_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa39_and0 = u_CSAwallace_cska32_csa18_csa_component_fa38_or0 & u_CSAwallace_cska32_csa19_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa39_and1 = u_CSAwallace_cska32_csa23_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa39_or0 = u_CSAwallace_cska32_csa23_csa_component_fa39_and0 | u_CSAwallace_cska32_csa23_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa39_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa40_and0 = u_CSAwallace_cska32_csa18_csa_component_fa39_or0 & u_CSAwallace_cska32_csa19_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa40_and1 = u_CSAwallace_cska32_csa23_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa40_or0 = u_CSAwallace_cska32_csa23_csa_component_fa40_and0 | u_CSAwallace_cska32_csa23_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa40_or0 ^ u_CSAwallace_cska32_csa19_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa41_and0 = u_CSAwallace_cska32_csa18_csa_component_fa40_or0 & u_CSAwallace_cska32_csa19_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa41_and1 = u_CSAwallace_cska32_csa23_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa41_or0 = u_CSAwallace_cska32_csa23_csa_component_fa41_and0 | u_CSAwallace_cska32_csa23_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa41_and1 ^ u_CSAwallace_cska32_csa19_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa42_and0 = u_CSAwallace_cska32_csa18_csa_component_fa41_and1 & u_CSAwallace_cska32_csa19_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa42_and1 = u_CSAwallace_cska32_csa23_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa42_or0 = u_CSAwallace_cska32_csa23_csa_component_fa42_and0 | u_CSAwallace_cska32_csa23_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa42_and1 ^ u_CSAwallace_cska32_csa19_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa43_and0 = u_CSAwallace_cska32_csa18_csa_component_fa42_and1 & u_CSAwallace_cska32_csa19_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa43_and1 = u_CSAwallace_cska32_csa23_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa43_or0 = u_CSAwallace_cska32_csa23_csa_component_fa43_and0 | u_CSAwallace_cska32_csa23_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa43_and1 ^ u_CSAwallace_cska32_csa19_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa44_and0 = u_CSAwallace_cska32_csa18_csa_component_fa43_and1 & u_CSAwallace_cska32_csa19_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa19_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa44_and1 = u_CSAwallace_cska32_csa23_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa19_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa44_or0 = u_CSAwallace_cska32_csa23_csa_component_fa44_and0 | u_CSAwallace_cska32_csa23_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa19_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa45_and1 = u_CSAwallace_cska32_csa19_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa19_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa19_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa46_and1 = u_CSAwallace_cska32_csa19_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa19_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa19_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa47_and1 = u_CSAwallace_cska32_csa19_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa19_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa19_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa48_and1 = u_CSAwallace_cska32_csa19_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa19_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa19_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa19_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa49_and1 = u_CSAwallace_cska32_csa19_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa19_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa23_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa19_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa23_csa_component_fa50_and1 = u_CSAwallace_cska32_csa14_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa19_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa20_csa_component_fa23_and0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa24_and0 = u_CSAwallace_cska32_csa20_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa20_csa_component_fa23_and0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa25_and0 = u_CSAwallace_cska32_csa20_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa26_and0 = u_CSAwallace_cska32_csa20_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa27_and0 = u_CSAwallace_cska32_csa20_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_and_0_27;
  assign u_CSAwallace_cska32_csa24_csa_component_fa27_and1 = u_CSAwallace_cska32_csa24_csa_component_fa27_xor0 & u_CSAwallace_cska32_and_0_27;
  assign u_CSAwallace_cska32_csa24_csa_component_fa27_or0 = u_CSAwallace_cska32_csa24_csa_component_fa27_and0 | u_CSAwallace_cska32_csa24_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa28_and0 = u_CSAwallace_cska32_csa20_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa9_csa_component_fa28_xor0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa28_and1 = u_CSAwallace_cska32_csa24_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa9_csa_component_fa28_xor0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa28_or0 = u_CSAwallace_cska32_csa24_csa_component_fa28_and0 | u_CSAwallace_cska32_csa24_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa29_and0 = u_CSAwallace_cska32_csa20_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa16_csa_component_fa29_xor0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa29_and1 = u_CSAwallace_cska32_csa24_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa16_csa_component_fa29_xor0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa29_or0 = u_CSAwallace_cska32_csa24_csa_component_fa29_and0 | u_CSAwallace_cska32_csa24_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa30_and0 = u_CSAwallace_cska32_csa20_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa30_xor0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa30_and1 = u_CSAwallace_cska32_csa24_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa30_xor0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa30_or0 = u_CSAwallace_cska32_csa24_csa_component_fa30_and0 | u_CSAwallace_cska32_csa24_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa31_and0 = u_CSAwallace_cska32_csa20_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa31_and1 = u_CSAwallace_cska32_csa24_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa31_or0 = u_CSAwallace_cska32_csa24_csa_component_fa31_and0 | u_CSAwallace_cska32_csa24_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa32_and0 = u_CSAwallace_cska32_csa20_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa32_and1 = u_CSAwallace_cska32_csa24_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa32_or0 = u_CSAwallace_cska32_csa24_csa_component_fa32_and0 | u_CSAwallace_cska32_csa24_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa33_and0 = u_CSAwallace_cska32_csa20_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa33_and1 = u_CSAwallace_cska32_csa24_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa33_or0 = u_CSAwallace_cska32_csa24_csa_component_fa33_and0 | u_CSAwallace_cska32_csa24_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa34_and0 = u_CSAwallace_cska32_csa20_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa34_and1 = u_CSAwallace_cska32_csa24_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa34_or0 = u_CSAwallace_cska32_csa24_csa_component_fa34_and0 | u_CSAwallace_cska32_csa24_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa35_and0 = u_CSAwallace_cska32_csa20_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa35_and1 = u_CSAwallace_cska32_csa24_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa35_or0 = u_CSAwallace_cska32_csa24_csa_component_fa35_and0 | u_CSAwallace_cska32_csa24_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa36_and0 = u_CSAwallace_cska32_csa20_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa36_and1 = u_CSAwallace_cska32_csa24_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa36_or0 = u_CSAwallace_cska32_csa24_csa_component_fa36_and0 | u_CSAwallace_cska32_csa24_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa37_and0 = u_CSAwallace_cska32_csa20_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa37_and1 = u_CSAwallace_cska32_csa24_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa37_or0 = u_CSAwallace_cska32_csa24_csa_component_fa37_and0 | u_CSAwallace_cska32_csa24_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa38_and0 = u_CSAwallace_cska32_csa20_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa38_and1 = u_CSAwallace_cska32_csa24_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa38_or0 = u_CSAwallace_cska32_csa24_csa_component_fa38_and0 | u_CSAwallace_cska32_csa24_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa39_and0 = u_CSAwallace_cska32_csa20_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa39_and1 = u_CSAwallace_cska32_csa24_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa39_or0 = u_CSAwallace_cska32_csa24_csa_component_fa39_and0 | u_CSAwallace_cska32_csa24_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa40_and0 = u_CSAwallace_cska32_csa20_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa40_and1 = u_CSAwallace_cska32_csa24_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa40_or0 = u_CSAwallace_cska32_csa24_csa_component_fa40_and0 | u_CSAwallace_cska32_csa24_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa41_and0 = u_CSAwallace_cska32_csa20_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa41_and1 = u_CSAwallace_cska32_csa24_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa41_or0 = u_CSAwallace_cska32_csa24_csa_component_fa41_and0 | u_CSAwallace_cska32_csa24_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa42_and0 = u_CSAwallace_cska32_csa20_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa42_and1 = u_CSAwallace_cska32_csa24_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa42_or0 = u_CSAwallace_cska32_csa24_csa_component_fa42_and0 | u_CSAwallace_cska32_csa24_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa43_and0 = u_CSAwallace_cska32_csa20_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa43_and1 = u_CSAwallace_cska32_csa24_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa43_or0 = u_CSAwallace_cska32_csa24_csa_component_fa43_and0 | u_CSAwallace_cska32_csa24_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa44_and0 = u_CSAwallace_cska32_csa20_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa44_and1 = u_CSAwallace_cska32_csa24_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa44_or0 = u_CSAwallace_cska32_csa24_csa_component_fa44_and0 | u_CSAwallace_cska32_csa24_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa45_and0 = u_CSAwallace_cska32_csa20_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa45_and1 = u_CSAwallace_cska32_csa24_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa45_or0 = u_CSAwallace_cska32_csa24_csa_component_fa45_and0 | u_CSAwallace_cska32_csa24_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa46_and0 = u_CSAwallace_cska32_csa20_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa46_and1 = u_CSAwallace_cska32_csa24_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa46_or0 = u_CSAwallace_cska32_csa24_csa_component_fa46_and0 | u_CSAwallace_cska32_csa24_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa47_and0 = u_CSAwallace_cska32_csa20_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa47_and1 = u_CSAwallace_cska32_csa24_csa_component_fa47_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa47_or0 = u_CSAwallace_cska32_csa24_csa_component_fa47_and0 | u_CSAwallace_cska32_csa24_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa48_and0 = u_CSAwallace_cska32_csa20_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa48_and1 = u_CSAwallace_cska32_csa24_csa_component_fa48_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa48_or0 = u_CSAwallace_cska32_csa24_csa_component_fa48_and0 | u_CSAwallace_cska32_csa24_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa49_and0 = u_CSAwallace_cska32_csa20_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa49_and1 = u_CSAwallace_cska32_csa24_csa_component_fa49_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa49_or0 = u_CSAwallace_cska32_csa24_csa_component_fa49_and0 | u_CSAwallace_cska32_csa24_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa50_and0 = u_CSAwallace_cska32_csa20_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa50_and1 = u_CSAwallace_cska32_csa24_csa_component_fa50_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa50_or0 = u_CSAwallace_cska32_csa24_csa_component_fa50_and0 | u_CSAwallace_cska32_csa24_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa51_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa51_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa51_and0 = u_CSAwallace_cska32_csa20_csa_component_fa51_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa51_and1 = u_CSAwallace_cska32_csa24_csa_component_fa51_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa51_or0 = u_CSAwallace_cska32_csa24_csa_component_fa51_and0 | u_CSAwallace_cska32_csa24_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa52_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa52_and0 = u_CSAwallace_cska32_csa20_csa_component_fa52_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa52_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa52_and1 = u_CSAwallace_cska32_csa24_csa_component_fa52_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa52_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa52_or0 = u_CSAwallace_cska32_csa24_csa_component_fa52_and0 | u_CSAwallace_cska32_csa24_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa53_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa53_and0 = u_CSAwallace_cska32_csa20_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa24_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa53_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa53_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa53_and1 = u_CSAwallace_cska32_csa24_csa_component_fa53_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa53_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa53_or0 = u_CSAwallace_cska32_csa24_csa_component_fa53_and0 | u_CSAwallace_cska32_csa24_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa54_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa54_and0 = u_CSAwallace_cska32_csa20_csa_component_fa54_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa54_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa54_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa54_and1 = u_CSAwallace_cska32_csa24_csa_component_fa54_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa54_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa54_or0 = u_CSAwallace_cska32_csa24_csa_component_fa54_and0 | u_CSAwallace_cska32_csa24_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa55_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa55_and0 = u_CSAwallace_cska32_csa20_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa55_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa55_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa55_and1 = u_CSAwallace_cska32_csa24_csa_component_fa55_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa55_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa55_or0 = u_CSAwallace_cska32_csa24_csa_component_fa55_and0 | u_CSAwallace_cska32_csa24_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa56_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa56_and0 = u_CSAwallace_cska32_csa20_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa56_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa56_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa56_and1 = u_CSAwallace_cska32_csa24_csa_component_fa56_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa56_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa56_or0 = u_CSAwallace_cska32_csa24_csa_component_fa56_and0 | u_CSAwallace_cska32_csa24_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa57_xor0 = u_CSAwallace_cska32_csa20_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa20_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa57_and0 = u_CSAwallace_cska32_csa20_csa_component_fa57_xor1 & u_CSAwallace_cska32_csa20_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa57_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa57_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa57_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa57_and1 = u_CSAwallace_cska32_csa24_csa_component_fa57_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa57_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa57_or0 = u_CSAwallace_cska32_csa24_csa_component_fa57_and0 | u_CSAwallace_cska32_csa24_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa58_xor0 = u_CSAwallace_cska32_csa15_csa_component_fa57_and1 ^ u_CSAwallace_cska32_csa20_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa58_and0 = u_CSAwallace_cska32_csa15_csa_component_fa57_and1 & u_CSAwallace_cska32_csa20_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa58_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa58_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa58_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa58_and1 = u_CSAwallace_cska32_csa24_csa_component_fa58_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa58_xor1;
  assign u_CSAwallace_cska32_csa24_csa_component_fa58_or0 = u_CSAwallace_cska32_csa24_csa_component_fa58_and0 | u_CSAwallace_cska32_csa24_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa5_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa5_xor0 ^ u_CSAwallace_cska32_csa22_csa_component_fa4_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa5_and0 = u_CSAwallace_cska32_csa22_csa_component_fa5_xor0 & u_CSAwallace_cska32_csa22_csa_component_fa4_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa6_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa6_xor0 ^ u_CSAwallace_cska32_csa22_csa_component_fa5_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa6_and0 = u_CSAwallace_cska32_csa22_csa_component_fa6_xor0 & u_CSAwallace_cska32_csa22_csa_component_fa5_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa7_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa7_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa6_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa7_and0 = u_CSAwallace_cska32_csa22_csa_component_fa7_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa6_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa8_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa8_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa7_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa8_and0 = u_CSAwallace_cska32_csa22_csa_component_fa8_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa7_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa9_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa9_and0 = u_CSAwallace_cska32_csa22_csa_component_fa9_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa8_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa10_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa10_and0 = u_CSAwallace_cska32_csa22_csa_component_fa10_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa9_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa10_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa10_and1 = u_CSAwallace_cska32_csa25_csa_component_fa10_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa10_or0 = u_CSAwallace_cska32_csa25_csa_component_fa10_and0 | u_CSAwallace_cska32_csa25_csa_component_fa10_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa11_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa11_and0 = u_CSAwallace_cska32_csa22_csa_component_fa11_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa11_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa11_and1 = u_CSAwallace_cska32_csa25_csa_component_fa11_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa11_or0 = u_CSAwallace_cska32_csa25_csa_component_fa11_and0 | u_CSAwallace_cska32_csa25_csa_component_fa11_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa12_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa12_and0 = u_CSAwallace_cska32_csa22_csa_component_fa12_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa12_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa12_and1 = u_CSAwallace_cska32_csa25_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa12_or0 = u_CSAwallace_cska32_csa25_csa_component_fa12_and0 | u_CSAwallace_cska32_csa25_csa_component_fa12_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa13_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa13_and0 = u_CSAwallace_cska32_csa22_csa_component_fa13_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa13_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa18_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa13_and1 = u_CSAwallace_cska32_csa25_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa18_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa13_or0 = u_CSAwallace_cska32_csa25_csa_component_fa13_and0 | u_CSAwallace_cska32_csa25_csa_component_fa13_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa14_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa14_and0 = u_CSAwallace_cska32_csa22_csa_component_fa14_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa14_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa14_xor0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa14_and1 = u_CSAwallace_cska32_csa25_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa14_xor0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa14_or0 = u_CSAwallace_cska32_csa25_csa_component_fa14_and0 | u_CSAwallace_cska32_csa25_csa_component_fa14_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa15_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa15_and0 = u_CSAwallace_cska32_csa22_csa_component_fa15_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa15_xor0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa15_and1 = u_CSAwallace_cska32_csa25_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa15_xor0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa15_or0 = u_CSAwallace_cska32_csa25_csa_component_fa15_and0 | u_CSAwallace_cska32_csa25_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa16_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa16_and0 = u_CSAwallace_cska32_csa22_csa_component_fa16_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa16_xor0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa16_and1 = u_CSAwallace_cska32_csa25_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa16_xor0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa16_or0 = u_CSAwallace_cska32_csa25_csa_component_fa16_and0 | u_CSAwallace_cska32_csa25_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa17_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa17_and0 = u_CSAwallace_cska32_csa22_csa_component_fa17_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa17_and1 = u_CSAwallace_cska32_csa25_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa17_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa17_or0 = u_CSAwallace_cska32_csa25_csa_component_fa17_and0 | u_CSAwallace_cska32_csa25_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa18_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa18_and0 = u_CSAwallace_cska32_csa22_csa_component_fa18_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa18_and1 = u_CSAwallace_cska32_csa25_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa18_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa18_or0 = u_CSAwallace_cska32_csa25_csa_component_fa18_and0 | u_CSAwallace_cska32_csa25_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa19_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa19_and0 = u_CSAwallace_cska32_csa22_csa_component_fa19_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa19_and1 = u_CSAwallace_cska32_csa25_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa19_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa19_or0 = u_CSAwallace_cska32_csa25_csa_component_fa19_and0 | u_CSAwallace_cska32_csa25_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa20_and0 = u_CSAwallace_cska32_csa22_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa20_and1 = u_CSAwallace_cska32_csa25_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa20_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa20_or0 = u_CSAwallace_cska32_csa25_csa_component_fa20_and0 | u_CSAwallace_cska32_csa25_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa21_and0 = u_CSAwallace_cska32_csa22_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa21_and1 = u_CSAwallace_cska32_csa25_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa21_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa21_or0 = u_CSAwallace_cska32_csa25_csa_component_fa21_and0 | u_CSAwallace_cska32_csa25_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa22_and0 = u_CSAwallace_cska32_csa22_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa22_and1 = u_CSAwallace_cska32_csa25_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa22_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa22_or0 = u_CSAwallace_cska32_csa25_csa_component_fa22_and0 | u_CSAwallace_cska32_csa25_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa23_and0 = u_CSAwallace_cska32_csa22_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa23_and1 = u_CSAwallace_cska32_csa25_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa23_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa23_or0 = u_CSAwallace_cska32_csa25_csa_component_fa23_and0 | u_CSAwallace_cska32_csa25_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa24_and0 = u_CSAwallace_cska32_csa22_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa24_and1 = u_CSAwallace_cska32_csa25_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa24_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa24_or0 = u_CSAwallace_cska32_csa25_csa_component_fa24_and0 | u_CSAwallace_cska32_csa25_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa25_and0 = u_CSAwallace_cska32_csa22_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa25_and1 = u_CSAwallace_cska32_csa25_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa25_or0 = u_CSAwallace_cska32_csa25_csa_component_fa25_and0 | u_CSAwallace_cska32_csa25_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa26_and0 = u_CSAwallace_cska32_csa22_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa26_and1 = u_CSAwallace_cska32_csa25_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa26_or0 = u_CSAwallace_cska32_csa25_csa_component_fa26_and0 | u_CSAwallace_cska32_csa25_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa27_and0 = u_CSAwallace_cska32_csa22_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa27_and1 = u_CSAwallace_cska32_csa25_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa27_or0 = u_CSAwallace_cska32_csa25_csa_component_fa27_and0 | u_CSAwallace_cska32_csa25_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa28_and0 = u_CSAwallace_cska32_csa22_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa28_and1 = u_CSAwallace_cska32_csa25_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa28_or0 = u_CSAwallace_cska32_csa25_csa_component_fa28_and0 | u_CSAwallace_cska32_csa25_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa29_and0 = u_CSAwallace_cska32_csa22_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa29_and1 = u_CSAwallace_cska32_csa25_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa29_or0 = u_CSAwallace_cska32_csa25_csa_component_fa29_and0 | u_CSAwallace_cska32_csa25_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa30_and0 = u_CSAwallace_cska32_csa22_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa30_and1 = u_CSAwallace_cska32_csa25_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa30_or0 = u_CSAwallace_cska32_csa25_csa_component_fa30_and0 | u_CSAwallace_cska32_csa25_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa31_and0 = u_CSAwallace_cska32_csa22_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa31_and1 = u_CSAwallace_cska32_csa25_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa31_or0 = u_CSAwallace_cska32_csa25_csa_component_fa31_and0 | u_CSAwallace_cska32_csa25_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa32_and0 = u_CSAwallace_cska32_csa22_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa32_and1 = u_CSAwallace_cska32_csa25_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa32_or0 = u_CSAwallace_cska32_csa25_csa_component_fa32_and0 | u_CSAwallace_cska32_csa25_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa33_and0 = u_CSAwallace_cska32_csa22_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa33_and1 = u_CSAwallace_cska32_csa25_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa33_or0 = u_CSAwallace_cska32_csa25_csa_component_fa33_and0 | u_CSAwallace_cska32_csa25_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa34_and0 = u_CSAwallace_cska32_csa22_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa34_and1 = u_CSAwallace_cska32_csa25_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa34_or0 = u_CSAwallace_cska32_csa25_csa_component_fa34_and0 | u_CSAwallace_cska32_csa25_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa35_and0 = u_CSAwallace_cska32_csa22_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa35_and1 = u_CSAwallace_cska32_csa25_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa35_or0 = u_CSAwallace_cska32_csa25_csa_component_fa35_and0 | u_CSAwallace_cska32_csa25_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa36_and0 = u_CSAwallace_cska32_csa22_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa36_and1 = u_CSAwallace_cska32_csa25_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa36_or0 = u_CSAwallace_cska32_csa25_csa_component_fa36_and0 | u_CSAwallace_cska32_csa25_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa37_and0 = u_CSAwallace_cska32_csa22_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa37_and1 = u_CSAwallace_cska32_csa25_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa37_or0 = u_CSAwallace_cska32_csa25_csa_component_fa37_and0 | u_CSAwallace_cska32_csa25_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa38_and0 = u_CSAwallace_cska32_csa22_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa25_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa38_and1 = u_CSAwallace_cska32_csa25_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa38_or0 = u_CSAwallace_cska32_csa25_csa_component_fa38_and0 | u_CSAwallace_cska32_csa25_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa22_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa39_and0 = u_CSAwallace_cska32_csa22_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa39_and1 = u_CSAwallace_cska32_csa25_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa39_or0 = u_CSAwallace_cska32_csa25_csa_component_fa39_and0 | u_CSAwallace_cska32_csa25_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa18_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa22_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa40_and0 = u_CSAwallace_cska32_csa18_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa22_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa25_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa40_and1 = u_CSAwallace_cska32_csa25_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa40_or0 = u_CSAwallace_cska32_csa25_csa_component_fa40_and0 | u_CSAwallace_cska32_csa25_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa23_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa41_and1 = u_CSAwallace_cska32_csa18_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa23_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa23_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa42_and1 = u_CSAwallace_cska32_csa18_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa23_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa18_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa23_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa43_and1 = u_CSAwallace_cska32_csa18_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa23_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa4_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa23_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa44_and1 = u_CSAwallace_cska32_csa4_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa23_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa45_xor1 = u_CSAwallace_cska32_and_31_14 ^ u_CSAwallace_cska32_csa23_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa25_csa_component_fa45_and1 = u_CSAwallace_cska32_and_31_14 & u_CSAwallace_cska32_csa23_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa20_or0 ^ u_CSAwallace_cska32_csa14_csa_component_fa20_and0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa21_and0 = u_CSAwallace_cska32_csa23_csa_component_fa20_or0 & u_CSAwallace_cska32_csa14_csa_component_fa20_and0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa21_or0 ^ u_CSAwallace_cska32_csa14_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa22_and0 = u_CSAwallace_cska32_csa23_csa_component_fa21_or0 & u_CSAwallace_cska32_csa14_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa22_or0 ^ u_CSAwallace_cska32_csa20_csa_component_fa23_xor0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa23_and0 = u_CSAwallace_cska32_csa23_csa_component_fa22_or0 & u_CSAwallace_cska32_csa20_csa_component_fa23_xor0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa23_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa24_xor0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa24_and0 = u_CSAwallace_cska32_csa23_csa_component_fa23_or0 & u_CSAwallace_cska32_csa24_csa_component_fa24_xor0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa24_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa25_xor0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa25_and0 = u_CSAwallace_cska32_csa23_csa_component_fa24_or0 & u_CSAwallace_cska32_csa24_csa_component_fa25_xor0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa25_and1 = u_CSAwallace_cska32_csa26_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa25_or0 = u_CSAwallace_cska32_csa26_csa_component_fa25_and0 | u_CSAwallace_cska32_csa26_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa25_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa26_xor0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa26_and0 = u_CSAwallace_cska32_csa23_csa_component_fa25_or0 & u_CSAwallace_cska32_csa24_csa_component_fa26_xor0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa26_and1 = u_CSAwallace_cska32_csa26_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa26_or0 = u_CSAwallace_cska32_csa26_csa_component_fa26_and0 | u_CSAwallace_cska32_csa26_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa26_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa27_and0 = u_CSAwallace_cska32_csa23_csa_component_fa26_or0 & u_CSAwallace_cska32_csa24_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa26_and0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa27_and1 = u_CSAwallace_cska32_csa26_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa26_and0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa27_or0 = u_CSAwallace_cska32_csa26_csa_component_fa27_and0 | u_CSAwallace_cska32_csa26_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa27_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa28_and0 = u_CSAwallace_cska32_csa23_csa_component_fa27_or0 & u_CSAwallace_cska32_csa24_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa28_and1 = u_CSAwallace_cska32_csa26_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa28_or0 = u_CSAwallace_cska32_csa26_csa_component_fa28_and0 | u_CSAwallace_cska32_csa26_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa28_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa29_and0 = u_CSAwallace_cska32_csa23_csa_component_fa28_or0 & u_CSAwallace_cska32_csa24_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa29_and1 = u_CSAwallace_cska32_csa26_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa29_or0 = u_CSAwallace_cska32_csa26_csa_component_fa29_and0 | u_CSAwallace_cska32_csa26_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa29_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa30_and0 = u_CSAwallace_cska32_csa23_csa_component_fa29_or0 & u_CSAwallace_cska32_csa24_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa30_and1 = u_CSAwallace_cska32_csa26_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa30_or0 = u_CSAwallace_cska32_csa26_csa_component_fa30_and0 | u_CSAwallace_cska32_csa26_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa30_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa31_and0 = u_CSAwallace_cska32_csa23_csa_component_fa30_or0 & u_CSAwallace_cska32_csa24_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa31_and1 = u_CSAwallace_cska32_csa26_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa31_or0 = u_CSAwallace_cska32_csa26_csa_component_fa31_and0 | u_CSAwallace_cska32_csa26_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa31_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa32_and0 = u_CSAwallace_cska32_csa23_csa_component_fa31_or0 & u_CSAwallace_cska32_csa24_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa32_and1 = u_CSAwallace_cska32_csa26_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa32_or0 = u_CSAwallace_cska32_csa26_csa_component_fa32_and0 | u_CSAwallace_cska32_csa26_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa32_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa33_and0 = u_CSAwallace_cska32_csa23_csa_component_fa32_or0 & u_CSAwallace_cska32_csa24_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa33_and1 = u_CSAwallace_cska32_csa26_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa33_or0 = u_CSAwallace_cska32_csa26_csa_component_fa33_and0 | u_CSAwallace_cska32_csa26_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa33_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa34_and0 = u_CSAwallace_cska32_csa23_csa_component_fa33_or0 & u_CSAwallace_cska32_csa24_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa34_and1 = u_CSAwallace_cska32_csa26_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa34_or0 = u_CSAwallace_cska32_csa26_csa_component_fa34_and0 | u_CSAwallace_cska32_csa26_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa34_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa35_and0 = u_CSAwallace_cska32_csa23_csa_component_fa34_or0 & u_CSAwallace_cska32_csa24_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa35_and1 = u_CSAwallace_cska32_csa26_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa35_or0 = u_CSAwallace_cska32_csa26_csa_component_fa35_and0 | u_CSAwallace_cska32_csa26_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa35_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa36_and0 = u_CSAwallace_cska32_csa23_csa_component_fa35_or0 & u_CSAwallace_cska32_csa24_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa36_and1 = u_CSAwallace_cska32_csa26_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa36_or0 = u_CSAwallace_cska32_csa26_csa_component_fa36_and0 | u_CSAwallace_cska32_csa26_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa36_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa37_and0 = u_CSAwallace_cska32_csa23_csa_component_fa36_or0 & u_CSAwallace_cska32_csa24_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa37_and1 = u_CSAwallace_cska32_csa26_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa37_or0 = u_CSAwallace_cska32_csa26_csa_component_fa37_and0 | u_CSAwallace_cska32_csa26_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa37_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa38_and0 = u_CSAwallace_cska32_csa23_csa_component_fa37_or0 & u_CSAwallace_cska32_csa24_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa38_and1 = u_CSAwallace_cska32_csa26_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa38_or0 = u_CSAwallace_cska32_csa26_csa_component_fa38_and0 | u_CSAwallace_cska32_csa26_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa38_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa39_and0 = u_CSAwallace_cska32_csa23_csa_component_fa38_or0 & u_CSAwallace_cska32_csa24_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa39_and1 = u_CSAwallace_cska32_csa26_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa39_or0 = u_CSAwallace_cska32_csa26_csa_component_fa39_and0 | u_CSAwallace_cska32_csa26_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa39_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa40_and0 = u_CSAwallace_cska32_csa23_csa_component_fa39_or0 & u_CSAwallace_cska32_csa24_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa40_and1 = u_CSAwallace_cska32_csa26_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa40_or0 = u_CSAwallace_cska32_csa26_csa_component_fa40_and0 | u_CSAwallace_cska32_csa26_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa40_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa41_and0 = u_CSAwallace_cska32_csa23_csa_component_fa40_or0 & u_CSAwallace_cska32_csa24_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa41_and1 = u_CSAwallace_cska32_csa26_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa41_or0 = u_CSAwallace_cska32_csa26_csa_component_fa41_and0 | u_CSAwallace_cska32_csa26_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa41_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa42_and0 = u_CSAwallace_cska32_csa23_csa_component_fa41_or0 & u_CSAwallace_cska32_csa24_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa42_and1 = u_CSAwallace_cska32_csa26_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa42_or0 = u_CSAwallace_cska32_csa26_csa_component_fa42_and0 | u_CSAwallace_cska32_csa26_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa42_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa43_and0 = u_CSAwallace_cska32_csa23_csa_component_fa42_or0 & u_CSAwallace_cska32_csa24_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa43_and1 = u_CSAwallace_cska32_csa26_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa43_or0 = u_CSAwallace_cska32_csa26_csa_component_fa43_and0 | u_CSAwallace_cska32_csa26_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa43_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa44_and0 = u_CSAwallace_cska32_csa23_csa_component_fa43_or0 & u_CSAwallace_cska32_csa24_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa44_and1 = u_CSAwallace_cska32_csa26_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa44_or0 = u_CSAwallace_cska32_csa26_csa_component_fa44_and0 | u_CSAwallace_cska32_csa26_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa44_or0 ^ u_CSAwallace_cska32_csa24_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa45_and0 = u_CSAwallace_cska32_csa23_csa_component_fa44_or0 & u_CSAwallace_cska32_csa24_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa45_and1 = u_CSAwallace_cska32_csa26_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa45_or0 = u_CSAwallace_cska32_csa26_csa_component_fa45_and0 | u_CSAwallace_cska32_csa26_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa45_and1 ^ u_CSAwallace_cska32_csa24_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa46_and0 = u_CSAwallace_cska32_csa23_csa_component_fa45_and1 & u_CSAwallace_cska32_csa24_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa46_and1 = u_CSAwallace_cska32_csa26_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa46_or0 = u_CSAwallace_cska32_csa26_csa_component_fa46_and0 | u_CSAwallace_cska32_csa26_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa46_and1 ^ u_CSAwallace_cska32_csa24_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa47_and0 = u_CSAwallace_cska32_csa23_csa_component_fa46_and1 & u_CSAwallace_cska32_csa24_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa47_and1 = u_CSAwallace_cska32_csa26_csa_component_fa47_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa47_or0 = u_CSAwallace_cska32_csa26_csa_component_fa47_and0 | u_CSAwallace_cska32_csa26_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa47_and1 ^ u_CSAwallace_cska32_csa24_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa48_and0 = u_CSAwallace_cska32_csa23_csa_component_fa47_and1 & u_CSAwallace_cska32_csa24_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa48_and1 = u_CSAwallace_cska32_csa26_csa_component_fa48_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa48_or0 = u_CSAwallace_cska32_csa26_csa_component_fa48_and0 | u_CSAwallace_cska32_csa26_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa48_and1 ^ u_CSAwallace_cska32_csa24_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa49_and0 = u_CSAwallace_cska32_csa23_csa_component_fa48_and1 & u_CSAwallace_cska32_csa24_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa49_and1 = u_CSAwallace_cska32_csa26_csa_component_fa49_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa49_or0 = u_CSAwallace_cska32_csa26_csa_component_fa49_and0 | u_CSAwallace_cska32_csa26_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa49_and1 ^ u_CSAwallace_cska32_csa24_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa50_and0 = u_CSAwallace_cska32_csa23_csa_component_fa49_and1 & u_CSAwallace_cska32_csa24_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa50_and1 = u_CSAwallace_cska32_csa26_csa_component_fa50_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa50_or0 = u_CSAwallace_cska32_csa26_csa_component_fa50_and0 | u_CSAwallace_cska32_csa26_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa51_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa50_and1 ^ u_CSAwallace_cska32_csa24_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa51_and0 = u_CSAwallace_cska32_csa23_csa_component_fa50_and1 & u_CSAwallace_cska32_csa24_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_csa24_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa51_and1 = u_CSAwallace_cska32_csa26_csa_component_fa51_xor0 & u_CSAwallace_cska32_csa24_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa51_or0 = u_CSAwallace_cska32_csa26_csa_component_fa51_and0 | u_CSAwallace_cska32_csa26_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa26_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa24_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa52_and1 = u_CSAwallace_cska32_csa24_csa_component_fa52_xor1 & u_CSAwallace_cska32_csa24_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa24_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa53_and1 = u_CSAwallace_cska32_csa24_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa24_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa24_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa54_and1 = u_CSAwallace_cska32_csa24_csa_component_fa54_xor1 & u_CSAwallace_cska32_csa24_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa24_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa55_and1 = u_CSAwallace_cska32_csa24_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa24_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa24_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa56_and1 = u_CSAwallace_cska32_csa24_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa24_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa57_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa24_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa57_and1 = u_CSAwallace_cska32_csa24_csa_component_fa57_xor1 & u_CSAwallace_cska32_csa24_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa58_xor1 = u_CSAwallace_cska32_csa24_csa_component_fa58_xor1 ^ u_CSAwallace_cska32_csa24_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa58_and1 = u_CSAwallace_cska32_csa24_csa_component_fa58_xor1 & u_CSAwallace_cska32_csa24_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa59_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa59_xor1 ^ u_CSAwallace_cska32_csa24_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_csa26_csa_component_fa59_and1 = u_CSAwallace_cska32_csa21_csa_component_fa59_xor1 & u_CSAwallace_cska32_csa24_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa6_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa6_xor0 ^ u_CSAwallace_cska32_csa25_csa_component_fa5_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa6_and0 = u_CSAwallace_cska32_csa25_csa_component_fa6_xor0 & u_CSAwallace_cska32_csa25_csa_component_fa5_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa7_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa7_xor0 ^ u_CSAwallace_cska32_csa25_csa_component_fa6_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa7_and0 = u_CSAwallace_cska32_csa25_csa_component_fa7_xor0 & u_CSAwallace_cska32_csa25_csa_component_fa6_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa8_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_csa25_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa8_and0 = u_CSAwallace_cska32_csa25_csa_component_fa8_xor0 & u_CSAwallace_cska32_csa25_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa25_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa9_and0 = u_CSAwallace_cska32_csa25_csa_component_fa9_xor0 & u_CSAwallace_cska32_csa25_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa10_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa10_and0 = u_CSAwallace_cska32_csa25_csa_component_fa10_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa11_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa11_and0 = u_CSAwallace_cska32_csa25_csa_component_fa11_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa10_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa12_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa12_and0 = u_CSAwallace_cska32_csa25_csa_component_fa12_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa11_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa13_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa13_and0 = u_CSAwallace_cska32_csa25_csa_component_fa13_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa12_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa14_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa14_and0 = u_CSAwallace_cska32_csa25_csa_component_fa14_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa13_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa15_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa15_and0 = u_CSAwallace_cska32_csa25_csa_component_fa15_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa14_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa15_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa15_and1 = u_CSAwallace_cska32_csa27_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa15_or0 = u_CSAwallace_cska32_csa27_csa_component_fa15_and0 | u_CSAwallace_cska32_csa27_csa_component_fa15_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa16_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa16_and0 = u_CSAwallace_cska32_csa25_csa_component_fa16_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa16_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa16_and1 = u_CSAwallace_cska32_csa27_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa16_or0 = u_CSAwallace_cska32_csa27_csa_component_fa16_and0 | u_CSAwallace_cska32_csa27_csa_component_fa16_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa17_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa17_and0 = u_CSAwallace_cska32_csa25_csa_component_fa17_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa17_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa17_and1 = u_CSAwallace_cska32_csa27_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa17_or0 = u_CSAwallace_cska32_csa27_csa_component_fa17_and0 | u_CSAwallace_cska32_csa27_csa_component_fa17_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa18_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa18_and0 = u_CSAwallace_cska32_csa25_csa_component_fa18_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa18_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa18_and1 = u_CSAwallace_cska32_csa27_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa18_or0 = u_CSAwallace_cska32_csa27_csa_component_fa18_and0 | u_CSAwallace_cska32_csa27_csa_component_fa18_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa19_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa19_and0 = u_CSAwallace_cska32_csa25_csa_component_fa19_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa19_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa19_and1 = u_CSAwallace_cska32_csa27_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa19_or0 = u_CSAwallace_cska32_csa27_csa_component_fa19_and0 | u_CSAwallace_cska32_csa27_csa_component_fa19_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa20_and0 = u_CSAwallace_cska32_csa25_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa20_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa23_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa20_and1 = u_CSAwallace_cska32_csa27_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa23_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa20_or0 = u_CSAwallace_cska32_csa27_csa_component_fa20_and0 | u_CSAwallace_cska32_csa27_csa_component_fa20_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa21_and0 = u_CSAwallace_cska32_csa25_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa21_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa21_xor0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa21_and1 = u_CSAwallace_cska32_csa27_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa21_xor0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa21_or0 = u_CSAwallace_cska32_csa27_csa_component_fa21_and0 | u_CSAwallace_cska32_csa27_csa_component_fa21_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa22_and0 = u_CSAwallace_cska32_csa25_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa22_xor0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa22_and1 = u_CSAwallace_cska32_csa27_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa22_xor0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa22_or0 = u_CSAwallace_cska32_csa27_csa_component_fa22_and0 | u_CSAwallace_cska32_csa27_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa23_and0 = u_CSAwallace_cska32_csa25_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa23_xor0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa23_and1 = u_CSAwallace_cska32_csa27_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa23_xor0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa23_or0 = u_CSAwallace_cska32_csa27_csa_component_fa23_and0 | u_CSAwallace_cska32_csa27_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa24_and0 = u_CSAwallace_cska32_csa25_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa24_xor0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa24_and1 = u_CSAwallace_cska32_csa27_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa24_xor0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa24_or0 = u_CSAwallace_cska32_csa27_csa_component_fa24_and0 | u_CSAwallace_cska32_csa27_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa25_and0 = u_CSAwallace_cska32_csa25_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa25_and1 = u_CSAwallace_cska32_csa27_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa25_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa25_or0 = u_CSAwallace_cska32_csa27_csa_component_fa25_and0 | u_CSAwallace_cska32_csa27_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa26_and0 = u_CSAwallace_cska32_csa25_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa26_and1 = u_CSAwallace_cska32_csa27_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa26_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa26_or0 = u_CSAwallace_cska32_csa27_csa_component_fa26_and0 | u_CSAwallace_cska32_csa27_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa27_and0 = u_CSAwallace_cska32_csa25_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa27_and1 = u_CSAwallace_cska32_csa27_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa27_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa27_or0 = u_CSAwallace_cska32_csa27_csa_component_fa27_and0 | u_CSAwallace_cska32_csa27_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa28_and0 = u_CSAwallace_cska32_csa25_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa28_and1 = u_CSAwallace_cska32_csa27_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa28_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa28_or0 = u_CSAwallace_cska32_csa27_csa_component_fa28_and0 | u_CSAwallace_cska32_csa27_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa29_and0 = u_CSAwallace_cska32_csa25_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa29_and1 = u_CSAwallace_cska32_csa27_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa29_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa29_or0 = u_CSAwallace_cska32_csa27_csa_component_fa29_and0 | u_CSAwallace_cska32_csa27_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa30_and0 = u_CSAwallace_cska32_csa25_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa30_and1 = u_CSAwallace_cska32_csa27_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa30_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa30_or0 = u_CSAwallace_cska32_csa27_csa_component_fa30_and0 | u_CSAwallace_cska32_csa27_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa31_and0 = u_CSAwallace_cska32_csa25_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa31_and1 = u_CSAwallace_cska32_csa27_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa31_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa31_or0 = u_CSAwallace_cska32_csa27_csa_component_fa31_and0 | u_CSAwallace_cska32_csa27_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa32_and0 = u_CSAwallace_cska32_csa25_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa32_and1 = u_CSAwallace_cska32_csa27_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa32_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa32_or0 = u_CSAwallace_cska32_csa27_csa_component_fa32_and0 | u_CSAwallace_cska32_csa27_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa33_and0 = u_CSAwallace_cska32_csa25_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa33_and1 = u_CSAwallace_cska32_csa27_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa33_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa33_or0 = u_CSAwallace_cska32_csa27_csa_component_fa33_and0 | u_CSAwallace_cska32_csa27_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa34_and0 = u_CSAwallace_cska32_csa25_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa34_and1 = u_CSAwallace_cska32_csa27_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa34_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa34_or0 = u_CSAwallace_cska32_csa27_csa_component_fa34_and0 | u_CSAwallace_cska32_csa27_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa35_and0 = u_CSAwallace_cska32_csa25_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa35_and1 = u_CSAwallace_cska32_csa27_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa35_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa35_or0 = u_CSAwallace_cska32_csa27_csa_component_fa35_and0 | u_CSAwallace_cska32_csa27_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa36_and0 = u_CSAwallace_cska32_csa25_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa36_and1 = u_CSAwallace_cska32_csa27_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa36_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa36_or0 = u_CSAwallace_cska32_csa27_csa_component_fa36_and0 | u_CSAwallace_cska32_csa27_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa37_and0 = u_CSAwallace_cska32_csa25_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa37_and1 = u_CSAwallace_cska32_csa27_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa37_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa37_or0 = u_CSAwallace_cska32_csa27_csa_component_fa37_and0 | u_CSAwallace_cska32_csa27_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa38_and0 = u_CSAwallace_cska32_csa25_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa38_and1 = u_CSAwallace_cska32_csa27_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa38_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa38_or0 = u_CSAwallace_cska32_csa27_csa_component_fa38_and0 | u_CSAwallace_cska32_csa27_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa39_and0 = u_CSAwallace_cska32_csa25_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa39_and1 = u_CSAwallace_cska32_csa27_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa39_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa39_or0 = u_CSAwallace_cska32_csa27_csa_component_fa39_and0 | u_CSAwallace_cska32_csa27_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa40_and0 = u_CSAwallace_cska32_csa25_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa40_and1 = u_CSAwallace_cska32_csa27_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa40_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa40_or0 = u_CSAwallace_cska32_csa27_csa_component_fa40_and0 | u_CSAwallace_cska32_csa27_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa41_and0 = u_CSAwallace_cska32_csa25_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa27_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa41_and1 = u_CSAwallace_cska32_csa27_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa41_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa41_or0 = u_CSAwallace_cska32_csa27_csa_component_fa41_and0 | u_CSAwallace_cska32_csa27_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa42_and0 = u_CSAwallace_cska32_csa25_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa42_and1 = u_CSAwallace_cska32_csa27_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa42_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa42_or0 = u_CSAwallace_cska32_csa27_csa_component_fa42_and0 | u_CSAwallace_cska32_csa27_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa43_and0 = u_CSAwallace_cska32_csa25_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa43_and1 = u_CSAwallace_cska32_csa27_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa43_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa43_or0 = u_CSAwallace_cska32_csa27_csa_component_fa43_and0 | u_CSAwallace_cska32_csa27_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa44_and0 = u_CSAwallace_cska32_csa25_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa44_and1 = u_CSAwallace_cska32_csa27_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa44_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa44_or0 = u_CSAwallace_cska32_csa27_csa_component_fa44_and0 | u_CSAwallace_cska32_csa27_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa25_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa45_and0 = u_CSAwallace_cska32_csa25_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa45_and1 = u_CSAwallace_cska32_csa27_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa45_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa45_or0 = u_CSAwallace_cska32_csa27_csa_component_fa45_and0 | u_CSAwallace_cska32_csa27_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa23_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa25_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa46_and0 = u_CSAwallace_cska32_csa23_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa25_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa27_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa46_and1 = u_CSAwallace_cska32_csa27_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa46_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa46_or0 = u_CSAwallace_cska32_csa27_csa_component_fa46_and0 | u_CSAwallace_cska32_csa27_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa47_and1 = u_CSAwallace_cska32_csa23_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa47_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa48_and1 = u_CSAwallace_cska32_csa23_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa48_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa49_and1 = u_CSAwallace_cska32_csa23_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa49_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa23_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa50_and1 = u_CSAwallace_cska32_csa23_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa50_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa14_csa_component_fa51_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa51_and1 = u_CSAwallace_cska32_csa14_csa_component_fa51_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa51_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa52_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa52_and1 = u_CSAwallace_cska32_csa7_csa_component_fa52_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa52_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa7_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa53_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa53_and1 = u_CSAwallace_cska32_csa7_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa53_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa54_xor1 = u_CSAwallace_cska32_and_31_23 ^ u_CSAwallace_cska32_csa26_csa_component_fa54_xor1;
  assign u_CSAwallace_cska32_csa27_csa_component_fa54_and1 = u_CSAwallace_cska32_and_31_23 & u_CSAwallace_cska32_csa26_csa_component_fa54_xor1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa7_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa7_xor0 ^ u_CSAwallace_cska32_csa27_csa_component_fa6_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa7_and0 = u_CSAwallace_cska32_csa27_csa_component_fa7_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa6_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa8_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_csa27_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa8_and0 = u_CSAwallace_cska32_csa27_csa_component_fa8_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa27_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa9_and0 = u_CSAwallace_cska32_csa27_csa_component_fa9_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa27_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa10_and0 = u_CSAwallace_cska32_csa27_csa_component_fa10_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa27_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa11_and0 = u_CSAwallace_cska32_csa27_csa_component_fa11_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa27_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa12_and0 = u_CSAwallace_cska32_csa27_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa27_csa_component_fa12_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa13_and0 = u_CSAwallace_cska32_csa27_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa12_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa27_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa14_and0 = u_CSAwallace_cska32_csa27_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa15_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa15_and0 = u_CSAwallace_cska32_csa27_csa_component_fa15_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa16_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa16_and0 = u_CSAwallace_cska32_csa27_csa_component_fa16_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa15_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa17_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa17_and0 = u_CSAwallace_cska32_csa27_csa_component_fa17_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa16_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa18_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa18_and0 = u_CSAwallace_cska32_csa27_csa_component_fa18_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa17_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa19_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa19_and0 = u_CSAwallace_cska32_csa27_csa_component_fa19_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa18_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa20_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa20_and0 = u_CSAwallace_cska32_csa27_csa_component_fa20_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa19_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa21_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa21_and0 = u_CSAwallace_cska32_csa27_csa_component_fa21_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa20_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa22_and0 = u_CSAwallace_cska32_csa27_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa21_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa22_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa21_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa22_and1 = u_CSAwallace_cska32_csa28_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa21_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa22_or0 = u_CSAwallace_cska32_csa28_csa_component_fa22_and0 | u_CSAwallace_cska32_csa28_csa_component_fa22_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa23_and0 = u_CSAwallace_cska32_csa27_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa23_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa22_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa23_and1 = u_CSAwallace_cska32_csa28_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa22_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa23_or0 = u_CSAwallace_cska32_csa28_csa_component_fa23_and0 | u_CSAwallace_cska32_csa28_csa_component_fa23_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa24_and0 = u_CSAwallace_cska32_csa27_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa24_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa23_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa24_and1 = u_CSAwallace_cska32_csa28_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa23_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa24_or0 = u_CSAwallace_cska32_csa28_csa_component_fa24_and0 | u_CSAwallace_cska32_csa28_csa_component_fa24_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa25_and0 = u_CSAwallace_cska32_csa27_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa25_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa25_and1 = u_CSAwallace_cska32_csa28_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa25_or0 = u_CSAwallace_cska32_csa28_csa_component_fa25_and0 | u_CSAwallace_cska32_csa28_csa_component_fa25_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa26_and0 = u_CSAwallace_cska32_csa27_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa26_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa26_and1 = u_CSAwallace_cska32_csa28_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa26_or0 = u_CSAwallace_cska32_csa28_csa_component_fa26_and0 | u_CSAwallace_cska32_csa28_csa_component_fa26_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa27_and0 = u_CSAwallace_cska32_csa27_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa27_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa27_and1 = u_CSAwallace_cska32_csa28_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa27_or0 = u_CSAwallace_cska32_csa28_csa_component_fa27_and0 | u_CSAwallace_cska32_csa28_csa_component_fa27_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa28_and0 = u_CSAwallace_cska32_csa27_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa28_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa28_and1 = u_CSAwallace_cska32_csa28_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa28_or0 = u_CSAwallace_cska32_csa28_csa_component_fa28_and0 | u_CSAwallace_cska32_csa28_csa_component_fa28_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa29_and0 = u_CSAwallace_cska32_csa27_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa29_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa29_and1 = u_CSAwallace_cska32_csa28_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa29_or0 = u_CSAwallace_cska32_csa28_csa_component_fa29_and0 | u_CSAwallace_cska32_csa28_csa_component_fa29_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa30_and0 = u_CSAwallace_cska32_csa27_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa30_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa30_and1 = u_CSAwallace_cska32_csa28_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa30_or0 = u_CSAwallace_cska32_csa28_csa_component_fa30_and0 | u_CSAwallace_cska32_csa28_csa_component_fa30_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa31_and0 = u_CSAwallace_cska32_csa27_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa31_and1 = u_CSAwallace_cska32_csa28_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa31_or0 = u_CSAwallace_cska32_csa28_csa_component_fa31_and0 | u_CSAwallace_cska32_csa28_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa32_and0 = u_CSAwallace_cska32_csa27_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa32_and1 = u_CSAwallace_cska32_csa28_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa32_or0 = u_CSAwallace_cska32_csa28_csa_component_fa32_and0 | u_CSAwallace_cska32_csa28_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa33_and0 = u_CSAwallace_cska32_csa27_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa33_and1 = u_CSAwallace_cska32_csa28_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa33_or0 = u_CSAwallace_cska32_csa28_csa_component_fa33_and0 | u_CSAwallace_cska32_csa28_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa34_and0 = u_CSAwallace_cska32_csa27_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa34_and1 = u_CSAwallace_cska32_csa28_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa34_or0 = u_CSAwallace_cska32_csa28_csa_component_fa34_and0 | u_CSAwallace_cska32_csa28_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa35_and0 = u_CSAwallace_cska32_csa27_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa35_and1 = u_CSAwallace_cska32_csa28_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa35_or0 = u_CSAwallace_cska32_csa28_csa_component_fa35_and0 | u_CSAwallace_cska32_csa28_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa36_and0 = u_CSAwallace_cska32_csa27_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa36_and1 = u_CSAwallace_cska32_csa28_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa36_or0 = u_CSAwallace_cska32_csa28_csa_component_fa36_and0 | u_CSAwallace_cska32_csa28_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa37_and0 = u_CSAwallace_cska32_csa27_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa37_and1 = u_CSAwallace_cska32_csa28_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa37_or0 = u_CSAwallace_cska32_csa28_csa_component_fa37_and0 | u_CSAwallace_cska32_csa28_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa38_and0 = u_CSAwallace_cska32_csa27_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa38_and1 = u_CSAwallace_cska32_csa28_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa38_or0 = u_CSAwallace_cska32_csa28_csa_component_fa38_and0 | u_CSAwallace_cska32_csa28_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa39_and0 = u_CSAwallace_cska32_csa27_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa39_and1 = u_CSAwallace_cska32_csa28_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa39_or0 = u_CSAwallace_cska32_csa28_csa_component_fa39_and0 | u_CSAwallace_cska32_csa28_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa40_and0 = u_CSAwallace_cska32_csa27_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa40_and1 = u_CSAwallace_cska32_csa28_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa40_or0 = u_CSAwallace_cska32_csa28_csa_component_fa40_and0 | u_CSAwallace_cska32_csa28_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa41_and0 = u_CSAwallace_cska32_csa27_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa41_and1 = u_CSAwallace_cska32_csa28_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa41_or0 = u_CSAwallace_cska32_csa28_csa_component_fa41_and0 | u_CSAwallace_cska32_csa28_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa42_and0 = u_CSAwallace_cska32_csa27_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa42_and1 = u_CSAwallace_cska32_csa28_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa42_or0 = u_CSAwallace_cska32_csa28_csa_component_fa42_and0 | u_CSAwallace_cska32_csa28_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa43_and0 = u_CSAwallace_cska32_csa27_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa43_and1 = u_CSAwallace_cska32_csa28_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa43_or0 = u_CSAwallace_cska32_csa28_csa_component_fa43_and0 | u_CSAwallace_cska32_csa28_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa44_and0 = u_CSAwallace_cska32_csa27_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa44_and1 = u_CSAwallace_cska32_csa28_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa44_or0 = u_CSAwallace_cska32_csa28_csa_component_fa44_and0 | u_CSAwallace_cska32_csa28_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa45_and0 = u_CSAwallace_cska32_csa27_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa45_and1 = u_CSAwallace_cska32_csa28_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa45_or0 = u_CSAwallace_cska32_csa28_csa_component_fa45_and0 | u_CSAwallace_cska32_csa28_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa46_and0 = u_CSAwallace_cska32_csa27_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa46_and1 = u_CSAwallace_cska32_csa28_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa46_or0 = u_CSAwallace_cska32_csa28_csa_component_fa46_and0 | u_CSAwallace_cska32_csa28_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa47_and0 = u_CSAwallace_cska32_csa27_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa47_and1 = u_CSAwallace_cska32_csa28_csa_component_fa47_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa47_or0 = u_CSAwallace_cska32_csa28_csa_component_fa47_and0 | u_CSAwallace_cska32_csa28_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa48_and0 = u_CSAwallace_cska32_csa27_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa48_and1 = u_CSAwallace_cska32_csa28_csa_component_fa48_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa48_or0 = u_CSAwallace_cska32_csa28_csa_component_fa48_and0 | u_CSAwallace_cska32_csa28_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa49_and0 = u_CSAwallace_cska32_csa27_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa49_and1 = u_CSAwallace_cska32_csa28_csa_component_fa49_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa49_or0 = u_CSAwallace_cska32_csa28_csa_component_fa49_and0 | u_CSAwallace_cska32_csa28_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa50_and0 = u_CSAwallace_cska32_csa27_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa50_and1 = u_CSAwallace_cska32_csa28_csa_component_fa50_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa50_or0 = u_CSAwallace_cska32_csa28_csa_component_fa50_and0 | u_CSAwallace_cska32_csa28_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa51_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa51_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa51_and0 = u_CSAwallace_cska32_csa27_csa_component_fa51_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa51_and1 = u_CSAwallace_cska32_csa28_csa_component_fa51_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa51_or0 = u_CSAwallace_cska32_csa28_csa_component_fa51_and0 | u_CSAwallace_cska32_csa28_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa52_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa52_and0 = u_CSAwallace_cska32_csa27_csa_component_fa52_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa52_and1 = u_CSAwallace_cska32_csa28_csa_component_fa52_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa28_csa_component_fa52_or0 = u_CSAwallace_cska32_csa28_csa_component_fa52_and0 | u_CSAwallace_cska32_csa28_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa53_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa53_and0 = u_CSAwallace_cska32_csa27_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa53_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa53_and1 = u_CSAwallace_cska32_csa28_csa_component_fa53_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa53_or0 = u_CSAwallace_cska32_csa28_csa_component_fa53_and0 | u_CSAwallace_cska32_csa28_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa54_xor0 = u_CSAwallace_cska32_csa27_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa54_and0 = u_CSAwallace_cska32_csa27_csa_component_fa54_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa54_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa54_and1 = u_CSAwallace_cska32_csa28_csa_component_fa54_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa54_or0 = u_CSAwallace_cska32_csa28_csa_component_fa54_and0 | u_CSAwallace_cska32_csa28_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa55_xor0 = u_CSAwallace_cska32_csa26_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa27_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa55_and0 = u_CSAwallace_cska32_csa26_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa27_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa28_csa_component_fa55_xor0 ^ u_CSAwallace_cska32_csa26_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa55_and1 = u_CSAwallace_cska32_csa28_csa_component_fa55_xor0 & u_CSAwallace_cska32_csa26_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa55_or0 = u_CSAwallace_cska32_csa28_csa_component_fa55_and0 | u_CSAwallace_cska32_csa28_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa56_and1 = u_CSAwallace_cska32_csa26_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa57_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa57_and1 = u_CSAwallace_cska32_csa26_csa_component_fa57_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa58_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa58_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa58_and1 = u_CSAwallace_cska32_csa26_csa_component_fa58_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa59_xor1 = u_CSAwallace_cska32_csa26_csa_component_fa59_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa59_and1 = u_CSAwallace_cska32_csa26_csa_component_fa59_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa60_xor1 = u_CSAwallace_cska32_csa21_csa_component_fa60_xor1 ^ u_CSAwallace_cska32_csa26_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa28_csa_component_fa60_and1 = u_CSAwallace_cska32_csa21_csa_component_fa60_xor1 & u_CSAwallace_cska32_csa26_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa8_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa8_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa8_and0 = u_CSAwallace_cska32_csa28_csa_component_fa8_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa7_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa9_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa9_and0 = u_CSAwallace_cska32_csa28_csa_component_fa9_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa10_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa10_and0 = u_CSAwallace_cska32_csa28_csa_component_fa10_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa11_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa11_and0 = u_CSAwallace_cska32_csa28_csa_component_fa11_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa12_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa12_and0 = u_CSAwallace_cska32_csa28_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa13_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa12_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa13_and0 = u_CSAwallace_cska32_csa28_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa12_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa14_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa14_and0 = u_CSAwallace_cska32_csa28_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa15_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa15_and0 = u_CSAwallace_cska32_csa28_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa16_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa16_and0 = u_CSAwallace_cska32_csa28_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa17_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa17_and0 = u_CSAwallace_cska32_csa28_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa18_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa17_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa18_and0 = u_CSAwallace_cska32_csa28_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa17_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa19_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa18_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa19_and0 = u_CSAwallace_cska32_csa28_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa18_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa20_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa19_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa20_and0 = u_CSAwallace_cska32_csa28_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa19_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa21_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa28_csa_component_fa20_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa21_and0 = u_CSAwallace_cska32_csa28_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa20_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa22_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa22_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa21_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa22_and0 = u_CSAwallace_cska32_csa28_csa_component_fa22_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa21_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa23_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa23_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa23_and0 = u_CSAwallace_cska32_csa28_csa_component_fa23_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa22_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa24_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa24_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa24_and0 = u_CSAwallace_cska32_csa28_csa_component_fa24_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa23_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa25_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa25_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa25_and0 = u_CSAwallace_cska32_csa28_csa_component_fa25_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa24_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa26_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa26_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa26_and0 = u_CSAwallace_cska32_csa28_csa_component_fa26_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa25_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa27_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa27_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa27_and0 = u_CSAwallace_cska32_csa28_csa_component_fa27_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa26_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa28_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa28_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa28_and0 = u_CSAwallace_cska32_csa28_csa_component_fa28_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa27_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa29_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa29_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa29_and0 = u_CSAwallace_cska32_csa28_csa_component_fa29_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa28_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa30_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa30_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa30_and0 = u_CSAwallace_cska32_csa28_csa_component_fa30_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa29_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa31_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa31_and0 = u_CSAwallace_cska32_csa28_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa30_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa31_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa31_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa30_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa31_and1 = u_CSAwallace_cska32_csa29_csa_component_fa31_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa30_and0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa31_or0 = u_CSAwallace_cska32_csa29_csa_component_fa31_and0 | u_CSAwallace_cska32_csa29_csa_component_fa31_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa32_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa32_and0 = u_CSAwallace_cska32_csa28_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa32_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa32_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa32_and1 = u_CSAwallace_cska32_csa29_csa_component_fa32_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa32_or0 = u_CSAwallace_cska32_csa29_csa_component_fa32_and0 | u_CSAwallace_cska32_csa29_csa_component_fa32_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa33_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa33_and0 = u_CSAwallace_cska32_csa28_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa33_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa33_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa33_and1 = u_CSAwallace_cska32_csa29_csa_component_fa33_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa33_or0 = u_CSAwallace_cska32_csa29_csa_component_fa33_and0 | u_CSAwallace_cska32_csa29_csa_component_fa33_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa34_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa34_and0 = u_CSAwallace_cska32_csa28_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa34_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa34_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa34_and1 = u_CSAwallace_cska32_csa29_csa_component_fa34_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa34_or0 = u_CSAwallace_cska32_csa29_csa_component_fa34_and0 | u_CSAwallace_cska32_csa29_csa_component_fa34_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa35_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa35_and0 = u_CSAwallace_cska32_csa28_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa35_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa35_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa35_and1 = u_CSAwallace_cska32_csa29_csa_component_fa35_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa35_or0 = u_CSAwallace_cska32_csa29_csa_component_fa35_and0 | u_CSAwallace_cska32_csa29_csa_component_fa35_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa36_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa36_and0 = u_CSAwallace_cska32_csa28_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa36_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa36_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa36_and1 = u_CSAwallace_cska32_csa29_csa_component_fa36_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa36_or0 = u_CSAwallace_cska32_csa29_csa_component_fa36_and0 | u_CSAwallace_cska32_csa29_csa_component_fa36_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa37_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa37_and0 = u_CSAwallace_cska32_csa28_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa37_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa37_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa37_and1 = u_CSAwallace_cska32_csa29_csa_component_fa37_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa37_or0 = u_CSAwallace_cska32_csa29_csa_component_fa37_and0 | u_CSAwallace_cska32_csa29_csa_component_fa37_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa38_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa38_and0 = u_CSAwallace_cska32_csa28_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa38_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa38_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa38_and1 = u_CSAwallace_cska32_csa29_csa_component_fa38_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa38_or0 = u_CSAwallace_cska32_csa29_csa_component_fa38_and0 | u_CSAwallace_cska32_csa29_csa_component_fa38_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa39_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa39_and0 = u_CSAwallace_cska32_csa28_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa39_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa39_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa39_and1 = u_CSAwallace_cska32_csa29_csa_component_fa39_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa39_or0 = u_CSAwallace_cska32_csa29_csa_component_fa39_and0 | u_CSAwallace_cska32_csa29_csa_component_fa39_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa40_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa40_and0 = u_CSAwallace_cska32_csa28_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa40_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa40_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa40_and1 = u_CSAwallace_cska32_csa29_csa_component_fa40_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa40_or0 = u_CSAwallace_cska32_csa29_csa_component_fa40_and0 | u_CSAwallace_cska32_csa29_csa_component_fa40_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa41_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa41_and0 = u_CSAwallace_cska32_csa28_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa41_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa41_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa41_and1 = u_CSAwallace_cska32_csa29_csa_component_fa41_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa41_or0 = u_CSAwallace_cska32_csa29_csa_component_fa41_and0 | u_CSAwallace_cska32_csa29_csa_component_fa41_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa42_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa42_and0 = u_CSAwallace_cska32_csa28_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa42_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa42_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa42_and1 = u_CSAwallace_cska32_csa29_csa_component_fa42_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa42_or0 = u_CSAwallace_cska32_csa29_csa_component_fa42_and0 | u_CSAwallace_cska32_csa29_csa_component_fa42_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa43_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa43_and0 = u_CSAwallace_cska32_csa28_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa43_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa43_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa43_and1 = u_CSAwallace_cska32_csa29_csa_component_fa43_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa43_or0 = u_CSAwallace_cska32_csa29_csa_component_fa43_and0 | u_CSAwallace_cska32_csa29_csa_component_fa43_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa44_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa44_and0 = u_CSAwallace_cska32_csa28_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa44_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa44_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa44_and1 = u_CSAwallace_cska32_csa29_csa_component_fa44_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa44_or0 = u_CSAwallace_cska32_csa29_csa_component_fa44_and0 | u_CSAwallace_cska32_csa29_csa_component_fa44_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa45_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa45_and0 = u_CSAwallace_cska32_csa28_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa45_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa45_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa45_and1 = u_CSAwallace_cska32_csa29_csa_component_fa45_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa45_or0 = u_CSAwallace_cska32_csa29_csa_component_fa45_and0 | u_CSAwallace_cska32_csa29_csa_component_fa45_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa46_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa46_and0 = u_CSAwallace_cska32_csa28_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa46_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa46_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa46_and1 = u_CSAwallace_cska32_csa29_csa_component_fa46_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa46_or0 = u_CSAwallace_cska32_csa29_csa_component_fa46_and0 | u_CSAwallace_cska32_csa29_csa_component_fa46_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa47_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa47_and0 = u_CSAwallace_cska32_csa28_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa47_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa47_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa47_and1 = u_CSAwallace_cska32_csa29_csa_component_fa47_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa47_or0 = u_CSAwallace_cska32_csa29_csa_component_fa47_and0 | u_CSAwallace_cska32_csa29_csa_component_fa47_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa48_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa48_and0 = u_CSAwallace_cska32_csa28_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa48_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa48_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa48_and1 = u_CSAwallace_cska32_csa29_csa_component_fa48_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa48_or0 = u_CSAwallace_cska32_csa29_csa_component_fa48_and0 | u_CSAwallace_cska32_csa29_csa_component_fa48_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa49_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa49_and0 = u_CSAwallace_cska32_csa28_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa49_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa49_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa49_and1 = u_CSAwallace_cska32_csa29_csa_component_fa49_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa49_or0 = u_CSAwallace_cska32_csa29_csa_component_fa49_and0 | u_CSAwallace_cska32_csa29_csa_component_fa49_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa50_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa50_and0 = u_CSAwallace_cska32_csa28_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa50_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa50_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa50_and1 = u_CSAwallace_cska32_csa29_csa_component_fa50_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa50_or0 = u_CSAwallace_cska32_csa29_csa_component_fa50_and0 | u_CSAwallace_cska32_csa29_csa_component_fa50_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa51_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa51_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa51_and0 = u_CSAwallace_cska32_csa28_csa_component_fa51_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa51_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa51_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa51_and1 = u_CSAwallace_cska32_csa29_csa_component_fa51_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa51_or0 = u_CSAwallace_cska32_csa29_csa_component_fa51_and0 | u_CSAwallace_cska32_csa29_csa_component_fa51_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa52_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa52_and0 = u_CSAwallace_cska32_csa28_csa_component_fa52_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa52_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa52_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa52_and1 = u_CSAwallace_cska32_csa29_csa_component_fa52_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa52_or0 = u_CSAwallace_cska32_csa29_csa_component_fa52_and0 | u_CSAwallace_cska32_csa29_csa_component_fa52_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa53_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa53_and0 = u_CSAwallace_cska32_csa28_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa53_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa53_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa53_and1 = u_CSAwallace_cska32_csa29_csa_component_fa53_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa53_or0 = u_CSAwallace_cska32_csa29_csa_component_fa53_and0 | u_CSAwallace_cska32_csa29_csa_component_fa53_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa54_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa54_and0 = u_CSAwallace_cska32_csa28_csa_component_fa54_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa54_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa54_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa54_and1 = u_CSAwallace_cska32_csa29_csa_component_fa54_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa54_or0 = u_CSAwallace_cska32_csa29_csa_component_fa54_and0 | u_CSAwallace_cska32_csa29_csa_component_fa54_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa55_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa55_and0 = u_CSAwallace_cska32_csa28_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa55_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa55_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa55_and1 = u_CSAwallace_cska32_csa29_csa_component_fa55_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa55_or0 = u_CSAwallace_cska32_csa29_csa_component_fa55_and0 | u_CSAwallace_cska32_csa29_csa_component_fa55_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa56_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa56_and0 = u_CSAwallace_cska32_csa28_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa56_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa56_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa56_and1 = u_CSAwallace_cska32_csa29_csa_component_fa56_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa56_or0 = u_CSAwallace_cska32_csa29_csa_component_fa56_and0 | u_CSAwallace_cska32_csa29_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa57_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa57_and0 = u_CSAwallace_cska32_csa28_csa_component_fa57_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa56_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa57_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa57_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa57_and1 = u_CSAwallace_cska32_csa29_csa_component_fa57_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa57_or0 = u_CSAwallace_cska32_csa29_csa_component_fa57_and0 | u_CSAwallace_cska32_csa29_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa58_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa58_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa58_and0 = u_CSAwallace_cska32_csa28_csa_component_fa58_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa57_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa58_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa58_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa58_and1 = u_CSAwallace_cska32_csa29_csa_component_fa58_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa58_or0 = u_CSAwallace_cska32_csa29_csa_component_fa58_and0 | u_CSAwallace_cska32_csa29_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa59_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa59_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa59_and0 = u_CSAwallace_cska32_csa28_csa_component_fa59_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa58_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa59_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa59_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa59_and1 = u_CSAwallace_cska32_csa29_csa_component_fa59_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa59_or0 = u_CSAwallace_cska32_csa29_csa_component_fa59_and0 | u_CSAwallace_cska32_csa29_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa60_xor0 = u_CSAwallace_cska32_csa28_csa_component_fa60_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa60_and0 = u_CSAwallace_cska32_csa28_csa_component_fa60_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa59_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa60_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa60_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa59_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa60_and1 = u_CSAwallace_cska32_csa29_csa_component_fa60_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa59_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa60_or0 = u_CSAwallace_cska32_csa29_csa_component_fa60_and0 | u_CSAwallace_cska32_csa29_csa_component_fa60_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa61_xor0 = u_CSAwallace_cska32_csa21_csa_component_fa61_xor1 ^ u_CSAwallace_cska32_csa28_csa_component_fa60_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa61_and0 = u_CSAwallace_cska32_csa21_csa_component_fa61_xor1 & u_CSAwallace_cska32_csa28_csa_component_fa60_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa61_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa61_xor0 ^ u_CSAwallace_cska32_csa21_csa_component_fa60_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa61_and1 = u_CSAwallace_cska32_csa29_csa_component_fa61_xor0 & u_CSAwallace_cska32_csa21_csa_component_fa60_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa61_or0 = u_CSAwallace_cska32_csa29_csa_component_fa61_and0 | u_CSAwallace_cska32_csa29_csa_component_fa61_and1;
  assign u_CSAwallace_cska32_csa29_csa_component_fa62_xor1 = u_CSAwallace_cska32_and_31_31 ^ u_CSAwallace_cska32_csa21_csa_component_fa61_or0;
  assign u_CSAwallace_cska32_csa29_csa_component_fa62_and1 = u_CSAwallace_cska32_and_31_31 & u_CSAwallace_cska32_csa21_csa_component_fa61_or0;
  assign u_CSAwallace_cska32_u_cska64_and_propagate00 = u_CSAwallace_cska32_and_0_0 & u_CSAwallace_cska32_csa10_csa_component_fa2_xor0;
  assign u_CSAwallace_cska32_u_cska64_and_propagate01 = u_CSAwallace_cska32_csa0_csa_component_fa1_xor0 & u_CSAwallace_cska32_csa17_csa_component_fa3_xor0;
  assign u_CSAwallace_cska32_u_cska64_and_propagate02 = u_CSAwallace_cska32_u_cska64_and_propagate00 & u_CSAwallace_cska32_u_cska64_and_propagate01;
  assign u_CSAwallace_cska32_u_cska64_mux2to10_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate02;
  assign u_CSAwallace_cska32_u_cska64_and_propagate13 = u_CSAwallace_cska32_csa22_csa_component_fa4_xor0 & u_CSAwallace_cska32_csa27_csa_component_fa6_xor0;
  assign u_CSAwallace_cska32_u_cska64_and_propagate14 = u_CSAwallace_cska32_csa25_csa_component_fa5_xor0 & u_CSAwallace_cska32_csa28_csa_component_fa7_xor0;
  assign u_CSAwallace_cska32_u_cska64_and_propagate15 = u_CSAwallace_cska32_u_cska64_and_propagate13 & u_CSAwallace_cska32_u_cska64_and_propagate14;
  assign u_CSAwallace_cska32_u_cska64_mux2to11_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate15;
  assign u_CSAwallace_cska32_u_cska64_xor9 = u_CSAwallace_cska32_csa29_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_u_cska64_fa8_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa9_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_u_cska64_fa8_and0 = u_CSAwallace_cska32_csa29_csa_component_fa9_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa8_and0;
  assign u_CSAwallace_cska32_u_cska64_xor10 = u_CSAwallace_cska32_csa29_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_u_cska64_fa9_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa10_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_u_cska64_fa9_and0 = u_CSAwallace_cska32_csa29_csa_component_fa10_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa9_and0;
  assign u_CSAwallace_cska32_u_cska64_fa9_xor1 = u_CSAwallace_cska32_u_cska64_fa9_xor0 ^ u_CSAwallace_cska32_u_cska64_fa8_and0;
  assign u_CSAwallace_cska32_u_cska64_fa9_and1 = u_CSAwallace_cska32_u_cska64_fa9_xor0 & u_CSAwallace_cska32_u_cska64_fa8_and0;
  assign u_CSAwallace_cska32_u_cska64_fa9_or0 = u_CSAwallace_cska32_u_cska64_fa9_and0 | u_CSAwallace_cska32_u_cska64_fa9_and1;
  assign u_CSAwallace_cska32_u_cska64_xor11 = u_CSAwallace_cska32_csa29_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_u_cska64_fa10_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa11_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_u_cska64_fa10_and0 = u_CSAwallace_cska32_csa29_csa_component_fa11_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa10_and0;
  assign u_CSAwallace_cska32_u_cska64_fa10_xor1 = u_CSAwallace_cska32_u_cska64_fa10_xor0 ^ u_CSAwallace_cska32_u_cska64_fa9_or0;
  assign u_CSAwallace_cska32_u_cska64_fa10_and1 = u_CSAwallace_cska32_u_cska64_fa10_xor0 & u_CSAwallace_cska32_u_cska64_fa9_or0;
  assign u_CSAwallace_cska32_u_cska64_fa10_or0 = u_CSAwallace_cska32_u_cska64_fa10_and0 | u_CSAwallace_cska32_u_cska64_fa10_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate26 = u_CSAwallace_cska32_csa29_csa_component_fa8_xor0 & u_CSAwallace_cska32_u_cska64_xor10;
  assign u_CSAwallace_cska32_u_cska64_and_propagate27 = u_CSAwallace_cska32_u_cska64_xor9 & u_CSAwallace_cska32_u_cska64_xor11;
  assign u_CSAwallace_cska32_u_cska64_and_propagate28 = u_CSAwallace_cska32_u_cska64_and_propagate26 & u_CSAwallace_cska32_u_cska64_and_propagate27;
  assign u_CSAwallace_cska32_u_cska64_mux2to12_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate28;
  assign u_CSAwallace_cska32_u_cska64_mux2to12_and1 = u_CSAwallace_cska32_u_cska64_fa10_or0 & u_CSAwallace_cska32_u_cska64_mux2to12_not0;
  assign u_CSAwallace_cska32_u_cska64_xor12 = u_CSAwallace_cska32_csa29_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_u_cska64_fa11_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa12_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_u_cska64_fa11_and0 = u_CSAwallace_cska32_csa29_csa_component_fa12_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa11_and0;
  assign u_CSAwallace_cska32_u_cska64_fa11_xor1 = u_CSAwallace_cska32_u_cska64_fa11_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to12_and1;
  assign u_CSAwallace_cska32_u_cska64_fa11_and1 = u_CSAwallace_cska32_u_cska64_fa11_xor0 & u_CSAwallace_cska32_u_cska64_mux2to12_and1;
  assign u_CSAwallace_cska32_u_cska64_fa11_or0 = u_CSAwallace_cska32_u_cska64_fa11_and0 | u_CSAwallace_cska32_u_cska64_fa11_and1;
  assign u_CSAwallace_cska32_u_cska64_xor13 = u_CSAwallace_cska32_csa29_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa12_and0;
  assign u_CSAwallace_cska32_u_cska64_fa12_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa13_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa12_and0;
  assign u_CSAwallace_cska32_u_cska64_fa12_and0 = u_CSAwallace_cska32_csa29_csa_component_fa13_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa12_and0;
  assign u_CSAwallace_cska32_u_cska64_fa12_xor1 = u_CSAwallace_cska32_u_cska64_fa12_xor0 ^ u_CSAwallace_cska32_u_cska64_fa11_or0;
  assign u_CSAwallace_cska32_u_cska64_fa12_and1 = u_CSAwallace_cska32_u_cska64_fa12_xor0 & u_CSAwallace_cska32_u_cska64_fa11_or0;
  assign u_CSAwallace_cska32_u_cska64_fa12_or0 = u_CSAwallace_cska32_u_cska64_fa12_and0 | u_CSAwallace_cska32_u_cska64_fa12_and1;
  assign u_CSAwallace_cska32_u_cska64_xor14 = u_CSAwallace_cska32_csa29_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_u_cska64_fa13_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa14_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_u_cska64_fa13_and0 = u_CSAwallace_cska32_csa29_csa_component_fa14_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa13_and0;
  assign u_CSAwallace_cska32_u_cska64_fa13_xor1 = u_CSAwallace_cska32_u_cska64_fa13_xor0 ^ u_CSAwallace_cska32_u_cska64_fa12_or0;
  assign u_CSAwallace_cska32_u_cska64_fa13_and1 = u_CSAwallace_cska32_u_cska64_fa13_xor0 & u_CSAwallace_cska32_u_cska64_fa12_or0;
  assign u_CSAwallace_cska32_u_cska64_fa13_or0 = u_CSAwallace_cska32_u_cska64_fa13_and0 | u_CSAwallace_cska32_u_cska64_fa13_and1;
  assign u_CSAwallace_cska32_u_cska64_xor15 = u_CSAwallace_cska32_csa29_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_u_cska64_fa14_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa15_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_u_cska64_fa14_and0 = u_CSAwallace_cska32_csa29_csa_component_fa15_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa14_and0;
  assign u_CSAwallace_cska32_u_cska64_fa14_xor1 = u_CSAwallace_cska32_u_cska64_fa14_xor0 ^ u_CSAwallace_cska32_u_cska64_fa13_or0;
  assign u_CSAwallace_cska32_u_cska64_fa14_and1 = u_CSAwallace_cska32_u_cska64_fa14_xor0 & u_CSAwallace_cska32_u_cska64_fa13_or0;
  assign u_CSAwallace_cska32_u_cska64_fa14_or0 = u_CSAwallace_cska32_u_cska64_fa14_and0 | u_CSAwallace_cska32_u_cska64_fa14_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate39 = u_CSAwallace_cska32_u_cska64_xor12 & u_CSAwallace_cska32_u_cska64_xor14;
  assign u_CSAwallace_cska32_u_cska64_and_propagate310 = u_CSAwallace_cska32_u_cska64_xor13 & u_CSAwallace_cska32_u_cska64_xor15;
  assign u_CSAwallace_cska32_u_cska64_and_propagate311 = u_CSAwallace_cska32_u_cska64_and_propagate39 & u_CSAwallace_cska32_u_cska64_and_propagate310;
  assign u_CSAwallace_cska32_u_cska64_mux2to13_and0 = u_CSAwallace_cska32_u_cska64_mux2to12_and1 & u_CSAwallace_cska32_u_cska64_and_propagate311;
  assign u_CSAwallace_cska32_u_cska64_mux2to13_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate311;
  assign u_CSAwallace_cska32_u_cska64_mux2to13_and1 = u_CSAwallace_cska32_u_cska64_fa14_or0 & u_CSAwallace_cska32_u_cska64_mux2to13_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to13_xor0 = u_CSAwallace_cska32_u_cska64_mux2to13_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to13_and1;
  assign u_CSAwallace_cska32_u_cska64_xor16 = u_CSAwallace_cska32_csa29_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_u_cska64_fa15_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa16_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_u_cska64_fa15_and0 = u_CSAwallace_cska32_csa29_csa_component_fa16_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa15_and0;
  assign u_CSAwallace_cska32_u_cska64_fa15_xor1 = u_CSAwallace_cska32_u_cska64_fa15_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to13_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa15_and1 = u_CSAwallace_cska32_u_cska64_fa15_xor0 & u_CSAwallace_cska32_u_cska64_mux2to13_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa15_or0 = u_CSAwallace_cska32_u_cska64_fa15_and0 | u_CSAwallace_cska32_u_cska64_fa15_and1;
  assign u_CSAwallace_cska32_u_cska64_xor17 = u_CSAwallace_cska32_csa29_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_u_cska64_fa16_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa17_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_u_cska64_fa16_and0 = u_CSAwallace_cska32_csa29_csa_component_fa17_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa16_and0;
  assign u_CSAwallace_cska32_u_cska64_fa16_xor1 = u_CSAwallace_cska32_u_cska64_fa16_xor0 ^ u_CSAwallace_cska32_u_cska64_fa15_or0;
  assign u_CSAwallace_cska32_u_cska64_fa16_and1 = u_CSAwallace_cska32_u_cska64_fa16_xor0 & u_CSAwallace_cska32_u_cska64_fa15_or0;
  assign u_CSAwallace_cska32_u_cska64_fa16_or0 = u_CSAwallace_cska32_u_cska64_fa16_and0 | u_CSAwallace_cska32_u_cska64_fa16_and1;
  assign u_CSAwallace_cska32_u_cska64_xor18 = u_CSAwallace_cska32_csa29_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa17_and0;
  assign u_CSAwallace_cska32_u_cska64_fa17_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa18_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa17_and0;
  assign u_CSAwallace_cska32_u_cska64_fa17_and0 = u_CSAwallace_cska32_csa29_csa_component_fa18_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa17_and0;
  assign u_CSAwallace_cska32_u_cska64_fa17_xor1 = u_CSAwallace_cska32_u_cska64_fa17_xor0 ^ u_CSAwallace_cska32_u_cska64_fa16_or0;
  assign u_CSAwallace_cska32_u_cska64_fa17_and1 = u_CSAwallace_cska32_u_cska64_fa17_xor0 & u_CSAwallace_cska32_u_cska64_fa16_or0;
  assign u_CSAwallace_cska32_u_cska64_fa17_or0 = u_CSAwallace_cska32_u_cska64_fa17_and0 | u_CSAwallace_cska32_u_cska64_fa17_and1;
  assign u_CSAwallace_cska32_u_cska64_xor19 = u_CSAwallace_cska32_csa29_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa18_and0;
  assign u_CSAwallace_cska32_u_cska64_fa18_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa19_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa18_and0;
  assign u_CSAwallace_cska32_u_cska64_fa18_and0 = u_CSAwallace_cska32_csa29_csa_component_fa19_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa18_and0;
  assign u_CSAwallace_cska32_u_cska64_fa18_xor1 = u_CSAwallace_cska32_u_cska64_fa18_xor0 ^ u_CSAwallace_cska32_u_cska64_fa17_or0;
  assign u_CSAwallace_cska32_u_cska64_fa18_and1 = u_CSAwallace_cska32_u_cska64_fa18_xor0 & u_CSAwallace_cska32_u_cska64_fa17_or0;
  assign u_CSAwallace_cska32_u_cska64_fa18_or0 = u_CSAwallace_cska32_u_cska64_fa18_and0 | u_CSAwallace_cska32_u_cska64_fa18_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate412 = u_CSAwallace_cska32_u_cska64_xor16 & u_CSAwallace_cska32_u_cska64_xor18;
  assign u_CSAwallace_cska32_u_cska64_and_propagate413 = u_CSAwallace_cska32_u_cska64_xor17 & u_CSAwallace_cska32_u_cska64_xor19;
  assign u_CSAwallace_cska32_u_cska64_and_propagate414 = u_CSAwallace_cska32_u_cska64_and_propagate412 & u_CSAwallace_cska32_u_cska64_and_propagate413;
  assign u_CSAwallace_cska32_u_cska64_mux2to14_and0 = u_CSAwallace_cska32_u_cska64_mux2to13_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate414;
  assign u_CSAwallace_cska32_u_cska64_mux2to14_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate414;
  assign u_CSAwallace_cska32_u_cska64_mux2to14_and1 = u_CSAwallace_cska32_u_cska64_fa18_or0 & u_CSAwallace_cska32_u_cska64_mux2to14_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to14_xor0 = u_CSAwallace_cska32_u_cska64_mux2to14_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to14_and1;
  assign u_CSAwallace_cska32_u_cska64_xor20 = u_CSAwallace_cska32_csa29_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa19_and0;
  assign u_CSAwallace_cska32_u_cska64_fa19_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa20_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa19_and0;
  assign u_CSAwallace_cska32_u_cska64_fa19_and0 = u_CSAwallace_cska32_csa29_csa_component_fa20_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa19_and0;
  assign u_CSAwallace_cska32_u_cska64_fa19_xor1 = u_CSAwallace_cska32_u_cska64_fa19_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to14_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa19_and1 = u_CSAwallace_cska32_u_cska64_fa19_xor0 & u_CSAwallace_cska32_u_cska64_mux2to14_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa19_or0 = u_CSAwallace_cska32_u_cska64_fa19_and0 | u_CSAwallace_cska32_u_cska64_fa19_and1;
  assign u_CSAwallace_cska32_u_cska64_xor21 = u_CSAwallace_cska32_csa29_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa20_and0;
  assign u_CSAwallace_cska32_u_cska64_fa20_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa21_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa20_and0;
  assign u_CSAwallace_cska32_u_cska64_fa20_and0 = u_CSAwallace_cska32_csa29_csa_component_fa21_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa20_and0;
  assign u_CSAwallace_cska32_u_cska64_fa20_xor1 = u_CSAwallace_cska32_u_cska64_fa20_xor0 ^ u_CSAwallace_cska32_u_cska64_fa19_or0;
  assign u_CSAwallace_cska32_u_cska64_fa20_and1 = u_CSAwallace_cska32_u_cska64_fa20_xor0 & u_CSAwallace_cska32_u_cska64_fa19_or0;
  assign u_CSAwallace_cska32_u_cska64_fa20_or0 = u_CSAwallace_cska32_u_cska64_fa20_and0 | u_CSAwallace_cska32_u_cska64_fa20_and1;
  assign u_CSAwallace_cska32_u_cska64_xor22 = u_CSAwallace_cska32_csa29_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa21_and0;
  assign u_CSAwallace_cska32_u_cska64_fa21_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa22_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa21_and0;
  assign u_CSAwallace_cska32_u_cska64_fa21_and0 = u_CSAwallace_cska32_csa29_csa_component_fa22_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa21_and0;
  assign u_CSAwallace_cska32_u_cska64_fa21_xor1 = u_CSAwallace_cska32_u_cska64_fa21_xor0 ^ u_CSAwallace_cska32_u_cska64_fa20_or0;
  assign u_CSAwallace_cska32_u_cska64_fa21_and1 = u_CSAwallace_cska32_u_cska64_fa21_xor0 & u_CSAwallace_cska32_u_cska64_fa20_or0;
  assign u_CSAwallace_cska32_u_cska64_fa21_or0 = u_CSAwallace_cska32_u_cska64_fa21_and0 | u_CSAwallace_cska32_u_cska64_fa21_and1;
  assign u_CSAwallace_cska32_u_cska64_xor23 = u_CSAwallace_cska32_csa29_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa22_and0;
  assign u_CSAwallace_cska32_u_cska64_fa22_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa23_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa22_and0;
  assign u_CSAwallace_cska32_u_cska64_fa22_and0 = u_CSAwallace_cska32_csa29_csa_component_fa23_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa22_and0;
  assign u_CSAwallace_cska32_u_cska64_fa22_xor1 = u_CSAwallace_cska32_u_cska64_fa22_xor0 ^ u_CSAwallace_cska32_u_cska64_fa21_or0;
  assign u_CSAwallace_cska32_u_cska64_fa22_and1 = u_CSAwallace_cska32_u_cska64_fa22_xor0 & u_CSAwallace_cska32_u_cska64_fa21_or0;
  assign u_CSAwallace_cska32_u_cska64_fa22_or0 = u_CSAwallace_cska32_u_cska64_fa22_and0 | u_CSAwallace_cska32_u_cska64_fa22_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate515 = u_CSAwallace_cska32_u_cska64_xor20 & u_CSAwallace_cska32_u_cska64_xor22;
  assign u_CSAwallace_cska32_u_cska64_and_propagate516 = u_CSAwallace_cska32_u_cska64_xor21 & u_CSAwallace_cska32_u_cska64_xor23;
  assign u_CSAwallace_cska32_u_cska64_and_propagate517 = u_CSAwallace_cska32_u_cska64_and_propagate515 & u_CSAwallace_cska32_u_cska64_and_propagate516;
  assign u_CSAwallace_cska32_u_cska64_mux2to15_and0 = u_CSAwallace_cska32_u_cska64_mux2to14_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate517;
  assign u_CSAwallace_cska32_u_cska64_mux2to15_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate517;
  assign u_CSAwallace_cska32_u_cska64_mux2to15_and1 = u_CSAwallace_cska32_u_cska64_fa22_or0 & u_CSAwallace_cska32_u_cska64_mux2to15_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to15_xor0 = u_CSAwallace_cska32_u_cska64_mux2to15_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to15_and1;
  assign u_CSAwallace_cska32_u_cska64_xor24 = u_CSAwallace_cska32_csa29_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa23_and0;
  assign u_CSAwallace_cska32_u_cska64_fa23_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa24_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa23_and0;
  assign u_CSAwallace_cska32_u_cska64_fa23_and0 = u_CSAwallace_cska32_csa29_csa_component_fa24_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa23_and0;
  assign u_CSAwallace_cska32_u_cska64_fa23_xor1 = u_CSAwallace_cska32_u_cska64_fa23_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to15_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa23_and1 = u_CSAwallace_cska32_u_cska64_fa23_xor0 & u_CSAwallace_cska32_u_cska64_mux2to15_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa23_or0 = u_CSAwallace_cska32_u_cska64_fa23_and0 | u_CSAwallace_cska32_u_cska64_fa23_and1;
  assign u_CSAwallace_cska32_u_cska64_xor25 = u_CSAwallace_cska32_csa29_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_u_cska64_fa24_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa25_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_u_cska64_fa24_and0 = u_CSAwallace_cska32_csa29_csa_component_fa25_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa24_and0;
  assign u_CSAwallace_cska32_u_cska64_fa24_xor1 = u_CSAwallace_cska32_u_cska64_fa24_xor0 ^ u_CSAwallace_cska32_u_cska64_fa23_or0;
  assign u_CSAwallace_cska32_u_cska64_fa24_and1 = u_CSAwallace_cska32_u_cska64_fa24_xor0 & u_CSAwallace_cska32_u_cska64_fa23_or0;
  assign u_CSAwallace_cska32_u_cska64_fa24_or0 = u_CSAwallace_cska32_u_cska64_fa24_and0 | u_CSAwallace_cska32_u_cska64_fa24_and1;
  assign u_CSAwallace_cska32_u_cska64_xor26 = u_CSAwallace_cska32_csa29_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_u_cska64_fa25_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa26_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_u_cska64_fa25_and0 = u_CSAwallace_cska32_csa29_csa_component_fa26_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa25_and0;
  assign u_CSAwallace_cska32_u_cska64_fa25_xor1 = u_CSAwallace_cska32_u_cska64_fa25_xor0 ^ u_CSAwallace_cska32_u_cska64_fa24_or0;
  assign u_CSAwallace_cska32_u_cska64_fa25_and1 = u_CSAwallace_cska32_u_cska64_fa25_xor0 & u_CSAwallace_cska32_u_cska64_fa24_or0;
  assign u_CSAwallace_cska32_u_cska64_fa25_or0 = u_CSAwallace_cska32_u_cska64_fa25_and0 | u_CSAwallace_cska32_u_cska64_fa25_and1;
  assign u_CSAwallace_cska32_u_cska64_xor27 = u_CSAwallace_cska32_csa29_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa26_and0;
  assign u_CSAwallace_cska32_u_cska64_fa26_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa27_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa26_and0;
  assign u_CSAwallace_cska32_u_cska64_fa26_and0 = u_CSAwallace_cska32_csa29_csa_component_fa27_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa26_and0;
  assign u_CSAwallace_cska32_u_cska64_fa26_xor1 = u_CSAwallace_cska32_u_cska64_fa26_xor0 ^ u_CSAwallace_cska32_u_cska64_fa25_or0;
  assign u_CSAwallace_cska32_u_cska64_fa26_and1 = u_CSAwallace_cska32_u_cska64_fa26_xor0 & u_CSAwallace_cska32_u_cska64_fa25_or0;
  assign u_CSAwallace_cska32_u_cska64_fa26_or0 = u_CSAwallace_cska32_u_cska64_fa26_and0 | u_CSAwallace_cska32_u_cska64_fa26_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate618 = u_CSAwallace_cska32_u_cska64_xor24 & u_CSAwallace_cska32_u_cska64_xor26;
  assign u_CSAwallace_cska32_u_cska64_and_propagate619 = u_CSAwallace_cska32_u_cska64_xor25 & u_CSAwallace_cska32_u_cska64_xor27;
  assign u_CSAwallace_cska32_u_cska64_and_propagate620 = u_CSAwallace_cska32_u_cska64_and_propagate618 & u_CSAwallace_cska32_u_cska64_and_propagate619;
  assign u_CSAwallace_cska32_u_cska64_mux2to16_and0 = u_CSAwallace_cska32_u_cska64_mux2to15_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate620;
  assign u_CSAwallace_cska32_u_cska64_mux2to16_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate620;
  assign u_CSAwallace_cska32_u_cska64_mux2to16_and1 = u_CSAwallace_cska32_u_cska64_fa26_or0 & u_CSAwallace_cska32_u_cska64_mux2to16_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to16_xor0 = u_CSAwallace_cska32_u_cska64_mux2to16_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to16_and1;
  assign u_CSAwallace_cska32_u_cska64_xor28 = u_CSAwallace_cska32_csa29_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa27_and0;
  assign u_CSAwallace_cska32_u_cska64_fa27_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa28_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa27_and0;
  assign u_CSAwallace_cska32_u_cska64_fa27_and0 = u_CSAwallace_cska32_csa29_csa_component_fa28_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa27_and0;
  assign u_CSAwallace_cska32_u_cska64_fa27_xor1 = u_CSAwallace_cska32_u_cska64_fa27_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to16_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa27_and1 = u_CSAwallace_cska32_u_cska64_fa27_xor0 & u_CSAwallace_cska32_u_cska64_mux2to16_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa27_or0 = u_CSAwallace_cska32_u_cska64_fa27_and0 | u_CSAwallace_cska32_u_cska64_fa27_and1;
  assign u_CSAwallace_cska32_u_cska64_xor29 = u_CSAwallace_cska32_csa29_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa28_and0;
  assign u_CSAwallace_cska32_u_cska64_fa28_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa29_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa28_and0;
  assign u_CSAwallace_cska32_u_cska64_fa28_and0 = u_CSAwallace_cska32_csa29_csa_component_fa29_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa28_and0;
  assign u_CSAwallace_cska32_u_cska64_fa28_xor1 = u_CSAwallace_cska32_u_cska64_fa28_xor0 ^ u_CSAwallace_cska32_u_cska64_fa27_or0;
  assign u_CSAwallace_cska32_u_cska64_fa28_and1 = u_CSAwallace_cska32_u_cska64_fa28_xor0 & u_CSAwallace_cska32_u_cska64_fa27_or0;
  assign u_CSAwallace_cska32_u_cska64_fa28_or0 = u_CSAwallace_cska32_u_cska64_fa28_and0 | u_CSAwallace_cska32_u_cska64_fa28_and1;
  assign u_CSAwallace_cska32_u_cska64_xor30 = u_CSAwallace_cska32_csa29_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa29_and0;
  assign u_CSAwallace_cska32_u_cska64_fa29_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa30_xor0 ^ u_CSAwallace_cska32_csa29_csa_component_fa29_and0;
  assign u_CSAwallace_cska32_u_cska64_fa29_and0 = u_CSAwallace_cska32_csa29_csa_component_fa30_xor0 & u_CSAwallace_cska32_csa29_csa_component_fa29_and0;
  assign u_CSAwallace_cska32_u_cska64_fa29_xor1 = u_CSAwallace_cska32_u_cska64_fa29_xor0 ^ u_CSAwallace_cska32_u_cska64_fa28_or0;
  assign u_CSAwallace_cska32_u_cska64_fa29_and1 = u_CSAwallace_cska32_u_cska64_fa29_xor0 & u_CSAwallace_cska32_u_cska64_fa28_or0;
  assign u_CSAwallace_cska32_u_cska64_fa29_or0 = u_CSAwallace_cska32_u_cska64_fa29_and0 | u_CSAwallace_cska32_u_cska64_fa29_and1;
  assign u_CSAwallace_cska32_u_cska64_xor31 = u_CSAwallace_cska32_csa29_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa30_and0;
  assign u_CSAwallace_cska32_u_cska64_fa30_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa31_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa30_and0;
  assign u_CSAwallace_cska32_u_cska64_fa30_and0 = u_CSAwallace_cska32_csa29_csa_component_fa31_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa30_and0;
  assign u_CSAwallace_cska32_u_cska64_fa30_xor1 = u_CSAwallace_cska32_u_cska64_fa30_xor0 ^ u_CSAwallace_cska32_u_cska64_fa29_or0;
  assign u_CSAwallace_cska32_u_cska64_fa30_and1 = u_CSAwallace_cska32_u_cska64_fa30_xor0 & u_CSAwallace_cska32_u_cska64_fa29_or0;
  assign u_CSAwallace_cska32_u_cska64_fa30_or0 = u_CSAwallace_cska32_u_cska64_fa30_and0 | u_CSAwallace_cska32_u_cska64_fa30_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate721 = u_CSAwallace_cska32_u_cska64_xor28 & u_CSAwallace_cska32_u_cska64_xor30;
  assign u_CSAwallace_cska32_u_cska64_and_propagate722 = u_CSAwallace_cska32_u_cska64_xor29 & u_CSAwallace_cska32_u_cska64_xor31;
  assign u_CSAwallace_cska32_u_cska64_and_propagate723 = u_CSAwallace_cska32_u_cska64_and_propagate721 & u_CSAwallace_cska32_u_cska64_and_propagate722;
  assign u_CSAwallace_cska32_u_cska64_mux2to17_and0 = u_CSAwallace_cska32_u_cska64_mux2to16_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate723;
  assign u_CSAwallace_cska32_u_cska64_mux2to17_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate723;
  assign u_CSAwallace_cska32_u_cska64_mux2to17_and1 = u_CSAwallace_cska32_u_cska64_fa30_or0 & u_CSAwallace_cska32_u_cska64_mux2to17_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to17_xor0 = u_CSAwallace_cska32_u_cska64_mux2to17_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to17_and1;
  assign u_CSAwallace_cska32_u_cska64_xor32 = u_CSAwallace_cska32_csa29_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_u_cska64_fa31_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa32_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_u_cska64_fa31_and0 = u_CSAwallace_cska32_csa29_csa_component_fa32_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa31_or0;
  assign u_CSAwallace_cska32_u_cska64_fa31_xor1 = u_CSAwallace_cska32_u_cska64_fa31_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to17_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa31_and1 = u_CSAwallace_cska32_u_cska64_fa31_xor0 & u_CSAwallace_cska32_u_cska64_mux2to17_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa31_or0 = u_CSAwallace_cska32_u_cska64_fa31_and0 | u_CSAwallace_cska32_u_cska64_fa31_and1;
  assign u_CSAwallace_cska32_u_cska64_xor33 = u_CSAwallace_cska32_csa29_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_u_cska64_fa32_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa33_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_u_cska64_fa32_and0 = u_CSAwallace_cska32_csa29_csa_component_fa33_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa32_or0;
  assign u_CSAwallace_cska32_u_cska64_fa32_xor1 = u_CSAwallace_cska32_u_cska64_fa32_xor0 ^ u_CSAwallace_cska32_u_cska64_fa31_or0;
  assign u_CSAwallace_cska32_u_cska64_fa32_and1 = u_CSAwallace_cska32_u_cska64_fa32_xor0 & u_CSAwallace_cska32_u_cska64_fa31_or0;
  assign u_CSAwallace_cska32_u_cska64_fa32_or0 = u_CSAwallace_cska32_u_cska64_fa32_and0 | u_CSAwallace_cska32_u_cska64_fa32_and1;
  assign u_CSAwallace_cska32_u_cska64_xor34 = u_CSAwallace_cska32_csa29_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_u_cska64_fa33_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa34_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_u_cska64_fa33_and0 = u_CSAwallace_cska32_csa29_csa_component_fa34_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa33_or0;
  assign u_CSAwallace_cska32_u_cska64_fa33_xor1 = u_CSAwallace_cska32_u_cska64_fa33_xor0 ^ u_CSAwallace_cska32_u_cska64_fa32_or0;
  assign u_CSAwallace_cska32_u_cska64_fa33_and1 = u_CSAwallace_cska32_u_cska64_fa33_xor0 & u_CSAwallace_cska32_u_cska64_fa32_or0;
  assign u_CSAwallace_cska32_u_cska64_fa33_or0 = u_CSAwallace_cska32_u_cska64_fa33_and0 | u_CSAwallace_cska32_u_cska64_fa33_and1;
  assign u_CSAwallace_cska32_u_cska64_xor35 = u_CSAwallace_cska32_csa29_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_u_cska64_fa34_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa35_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_u_cska64_fa34_and0 = u_CSAwallace_cska32_csa29_csa_component_fa35_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa34_or0;
  assign u_CSAwallace_cska32_u_cska64_fa34_xor1 = u_CSAwallace_cska32_u_cska64_fa34_xor0 ^ u_CSAwallace_cska32_u_cska64_fa33_or0;
  assign u_CSAwallace_cska32_u_cska64_fa34_and1 = u_CSAwallace_cska32_u_cska64_fa34_xor0 & u_CSAwallace_cska32_u_cska64_fa33_or0;
  assign u_CSAwallace_cska32_u_cska64_fa34_or0 = u_CSAwallace_cska32_u_cska64_fa34_and0 | u_CSAwallace_cska32_u_cska64_fa34_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate824 = u_CSAwallace_cska32_u_cska64_xor32 & u_CSAwallace_cska32_u_cska64_xor34;
  assign u_CSAwallace_cska32_u_cska64_and_propagate825 = u_CSAwallace_cska32_u_cska64_xor33 & u_CSAwallace_cska32_u_cska64_xor35;
  assign u_CSAwallace_cska32_u_cska64_and_propagate826 = u_CSAwallace_cska32_u_cska64_and_propagate824 & u_CSAwallace_cska32_u_cska64_and_propagate825;
  assign u_CSAwallace_cska32_u_cska64_mux2to18_and0 = u_CSAwallace_cska32_u_cska64_mux2to17_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate826;
  assign u_CSAwallace_cska32_u_cska64_mux2to18_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate826;
  assign u_CSAwallace_cska32_u_cska64_mux2to18_and1 = u_CSAwallace_cska32_u_cska64_fa34_or0 & u_CSAwallace_cska32_u_cska64_mux2to18_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to18_xor0 = u_CSAwallace_cska32_u_cska64_mux2to18_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to18_and1;
  assign u_CSAwallace_cska32_u_cska64_xor36 = u_CSAwallace_cska32_csa29_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_u_cska64_fa35_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa36_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_u_cska64_fa35_and0 = u_CSAwallace_cska32_csa29_csa_component_fa36_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa35_or0;
  assign u_CSAwallace_cska32_u_cska64_fa35_xor1 = u_CSAwallace_cska32_u_cska64_fa35_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to18_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa35_and1 = u_CSAwallace_cska32_u_cska64_fa35_xor0 & u_CSAwallace_cska32_u_cska64_mux2to18_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa35_or0 = u_CSAwallace_cska32_u_cska64_fa35_and0 | u_CSAwallace_cska32_u_cska64_fa35_and1;
  assign u_CSAwallace_cska32_u_cska64_xor37 = u_CSAwallace_cska32_csa29_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_u_cska64_fa36_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa37_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_u_cska64_fa36_and0 = u_CSAwallace_cska32_csa29_csa_component_fa37_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa36_or0;
  assign u_CSAwallace_cska32_u_cska64_fa36_xor1 = u_CSAwallace_cska32_u_cska64_fa36_xor0 ^ u_CSAwallace_cska32_u_cska64_fa35_or0;
  assign u_CSAwallace_cska32_u_cska64_fa36_and1 = u_CSAwallace_cska32_u_cska64_fa36_xor0 & u_CSAwallace_cska32_u_cska64_fa35_or0;
  assign u_CSAwallace_cska32_u_cska64_fa36_or0 = u_CSAwallace_cska32_u_cska64_fa36_and0 | u_CSAwallace_cska32_u_cska64_fa36_and1;
  assign u_CSAwallace_cska32_u_cska64_xor38 = u_CSAwallace_cska32_csa29_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_u_cska64_fa37_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa38_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_u_cska64_fa37_and0 = u_CSAwallace_cska32_csa29_csa_component_fa38_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa37_or0;
  assign u_CSAwallace_cska32_u_cska64_fa37_xor1 = u_CSAwallace_cska32_u_cska64_fa37_xor0 ^ u_CSAwallace_cska32_u_cska64_fa36_or0;
  assign u_CSAwallace_cska32_u_cska64_fa37_and1 = u_CSAwallace_cska32_u_cska64_fa37_xor0 & u_CSAwallace_cska32_u_cska64_fa36_or0;
  assign u_CSAwallace_cska32_u_cska64_fa37_or0 = u_CSAwallace_cska32_u_cska64_fa37_and0 | u_CSAwallace_cska32_u_cska64_fa37_and1;
  assign u_CSAwallace_cska32_u_cska64_xor39 = u_CSAwallace_cska32_csa29_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_u_cska64_fa38_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa39_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_u_cska64_fa38_and0 = u_CSAwallace_cska32_csa29_csa_component_fa39_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa38_or0;
  assign u_CSAwallace_cska32_u_cska64_fa38_xor1 = u_CSAwallace_cska32_u_cska64_fa38_xor0 ^ u_CSAwallace_cska32_u_cska64_fa37_or0;
  assign u_CSAwallace_cska32_u_cska64_fa38_and1 = u_CSAwallace_cska32_u_cska64_fa38_xor0 & u_CSAwallace_cska32_u_cska64_fa37_or0;
  assign u_CSAwallace_cska32_u_cska64_fa38_or0 = u_CSAwallace_cska32_u_cska64_fa38_and0 | u_CSAwallace_cska32_u_cska64_fa38_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate927 = u_CSAwallace_cska32_u_cska64_xor36 & u_CSAwallace_cska32_u_cska64_xor38;
  assign u_CSAwallace_cska32_u_cska64_and_propagate928 = u_CSAwallace_cska32_u_cska64_xor37 & u_CSAwallace_cska32_u_cska64_xor39;
  assign u_CSAwallace_cska32_u_cska64_and_propagate929 = u_CSAwallace_cska32_u_cska64_and_propagate927 & u_CSAwallace_cska32_u_cska64_and_propagate928;
  assign u_CSAwallace_cska32_u_cska64_mux2to19_and0 = u_CSAwallace_cska32_u_cska64_mux2to18_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate929;
  assign u_CSAwallace_cska32_u_cska64_mux2to19_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate929;
  assign u_CSAwallace_cska32_u_cska64_mux2to19_and1 = u_CSAwallace_cska32_u_cska64_fa38_or0 & u_CSAwallace_cska32_u_cska64_mux2to19_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to19_xor0 = u_CSAwallace_cska32_u_cska64_mux2to19_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to19_and1;
  assign u_CSAwallace_cska32_u_cska64_xor40 = u_CSAwallace_cska32_csa29_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_u_cska64_fa39_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa40_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_u_cska64_fa39_and0 = u_CSAwallace_cska32_csa29_csa_component_fa40_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa39_or0;
  assign u_CSAwallace_cska32_u_cska64_fa39_xor1 = u_CSAwallace_cska32_u_cska64_fa39_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to19_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa39_and1 = u_CSAwallace_cska32_u_cska64_fa39_xor0 & u_CSAwallace_cska32_u_cska64_mux2to19_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa39_or0 = u_CSAwallace_cska32_u_cska64_fa39_and0 | u_CSAwallace_cska32_u_cska64_fa39_and1;
  assign u_CSAwallace_cska32_u_cska64_xor41 = u_CSAwallace_cska32_csa29_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_u_cska64_fa40_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa41_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_u_cska64_fa40_and0 = u_CSAwallace_cska32_csa29_csa_component_fa41_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa40_or0;
  assign u_CSAwallace_cska32_u_cska64_fa40_xor1 = u_CSAwallace_cska32_u_cska64_fa40_xor0 ^ u_CSAwallace_cska32_u_cska64_fa39_or0;
  assign u_CSAwallace_cska32_u_cska64_fa40_and1 = u_CSAwallace_cska32_u_cska64_fa40_xor0 & u_CSAwallace_cska32_u_cska64_fa39_or0;
  assign u_CSAwallace_cska32_u_cska64_fa40_or0 = u_CSAwallace_cska32_u_cska64_fa40_and0 | u_CSAwallace_cska32_u_cska64_fa40_and1;
  assign u_CSAwallace_cska32_u_cska64_xor42 = u_CSAwallace_cska32_csa29_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_u_cska64_fa41_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa42_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_u_cska64_fa41_and0 = u_CSAwallace_cska32_csa29_csa_component_fa42_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa41_or0;
  assign u_CSAwallace_cska32_u_cska64_fa41_xor1 = u_CSAwallace_cska32_u_cska64_fa41_xor0 ^ u_CSAwallace_cska32_u_cska64_fa40_or0;
  assign u_CSAwallace_cska32_u_cska64_fa41_and1 = u_CSAwallace_cska32_u_cska64_fa41_xor0 & u_CSAwallace_cska32_u_cska64_fa40_or0;
  assign u_CSAwallace_cska32_u_cska64_fa41_or0 = u_CSAwallace_cska32_u_cska64_fa41_and0 | u_CSAwallace_cska32_u_cska64_fa41_and1;
  assign u_CSAwallace_cska32_u_cska64_xor43 = u_CSAwallace_cska32_csa29_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_u_cska64_fa42_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa43_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_u_cska64_fa42_and0 = u_CSAwallace_cska32_csa29_csa_component_fa43_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa42_or0;
  assign u_CSAwallace_cska32_u_cska64_fa42_xor1 = u_CSAwallace_cska32_u_cska64_fa42_xor0 ^ u_CSAwallace_cska32_u_cska64_fa41_or0;
  assign u_CSAwallace_cska32_u_cska64_fa42_and1 = u_CSAwallace_cska32_u_cska64_fa42_xor0 & u_CSAwallace_cska32_u_cska64_fa41_or0;
  assign u_CSAwallace_cska32_u_cska64_fa42_or0 = u_CSAwallace_cska32_u_cska64_fa42_and0 | u_CSAwallace_cska32_u_cska64_fa42_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1030 = u_CSAwallace_cska32_u_cska64_xor40 & u_CSAwallace_cska32_u_cska64_xor42;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1031 = u_CSAwallace_cska32_u_cska64_xor41 & u_CSAwallace_cska32_u_cska64_xor43;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1032 = u_CSAwallace_cska32_u_cska64_and_propagate1030 & u_CSAwallace_cska32_u_cska64_and_propagate1031;
  assign u_CSAwallace_cska32_u_cska64_mux2to110_and0 = u_CSAwallace_cska32_u_cska64_mux2to19_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate1032;
  assign u_CSAwallace_cska32_u_cska64_mux2to110_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate1032;
  assign u_CSAwallace_cska32_u_cska64_mux2to110_and1 = u_CSAwallace_cska32_u_cska64_fa42_or0 & u_CSAwallace_cska32_u_cska64_mux2to110_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to110_xor0 = u_CSAwallace_cska32_u_cska64_mux2to110_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to110_and1;
  assign u_CSAwallace_cska32_u_cska64_xor44 = u_CSAwallace_cska32_csa29_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_u_cska64_fa43_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa44_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_u_cska64_fa43_and0 = u_CSAwallace_cska32_csa29_csa_component_fa44_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa43_or0;
  assign u_CSAwallace_cska32_u_cska64_fa43_xor1 = u_CSAwallace_cska32_u_cska64_fa43_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to110_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa43_and1 = u_CSAwallace_cska32_u_cska64_fa43_xor0 & u_CSAwallace_cska32_u_cska64_mux2to110_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa43_or0 = u_CSAwallace_cska32_u_cska64_fa43_and0 | u_CSAwallace_cska32_u_cska64_fa43_and1;
  assign u_CSAwallace_cska32_u_cska64_xor45 = u_CSAwallace_cska32_csa29_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_u_cska64_fa44_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa45_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_u_cska64_fa44_and0 = u_CSAwallace_cska32_csa29_csa_component_fa45_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa44_or0;
  assign u_CSAwallace_cska32_u_cska64_fa44_xor1 = u_CSAwallace_cska32_u_cska64_fa44_xor0 ^ u_CSAwallace_cska32_u_cska64_fa43_or0;
  assign u_CSAwallace_cska32_u_cska64_fa44_and1 = u_CSAwallace_cska32_u_cska64_fa44_xor0 & u_CSAwallace_cska32_u_cska64_fa43_or0;
  assign u_CSAwallace_cska32_u_cska64_fa44_or0 = u_CSAwallace_cska32_u_cska64_fa44_and0 | u_CSAwallace_cska32_u_cska64_fa44_and1;
  assign u_CSAwallace_cska32_u_cska64_xor46 = u_CSAwallace_cska32_csa29_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_u_cska64_fa45_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa46_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_u_cska64_fa45_and0 = u_CSAwallace_cska32_csa29_csa_component_fa46_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa45_or0;
  assign u_CSAwallace_cska32_u_cska64_fa45_xor1 = u_CSAwallace_cska32_u_cska64_fa45_xor0 ^ u_CSAwallace_cska32_u_cska64_fa44_or0;
  assign u_CSAwallace_cska32_u_cska64_fa45_and1 = u_CSAwallace_cska32_u_cska64_fa45_xor0 & u_CSAwallace_cska32_u_cska64_fa44_or0;
  assign u_CSAwallace_cska32_u_cska64_fa45_or0 = u_CSAwallace_cska32_u_cska64_fa45_and0 | u_CSAwallace_cska32_u_cska64_fa45_and1;
  assign u_CSAwallace_cska32_u_cska64_xor47 = u_CSAwallace_cska32_csa29_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_u_cska64_fa46_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa47_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_u_cska64_fa46_and0 = u_CSAwallace_cska32_csa29_csa_component_fa47_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa46_or0;
  assign u_CSAwallace_cska32_u_cska64_fa46_xor1 = u_CSAwallace_cska32_u_cska64_fa46_xor0 ^ u_CSAwallace_cska32_u_cska64_fa45_or0;
  assign u_CSAwallace_cska32_u_cska64_fa46_and1 = u_CSAwallace_cska32_u_cska64_fa46_xor0 & u_CSAwallace_cska32_u_cska64_fa45_or0;
  assign u_CSAwallace_cska32_u_cska64_fa46_or0 = u_CSAwallace_cska32_u_cska64_fa46_and0 | u_CSAwallace_cska32_u_cska64_fa46_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1133 = u_CSAwallace_cska32_u_cska64_xor44 & u_CSAwallace_cska32_u_cska64_xor46;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1134 = u_CSAwallace_cska32_u_cska64_xor45 & u_CSAwallace_cska32_u_cska64_xor47;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1135 = u_CSAwallace_cska32_u_cska64_and_propagate1133 & u_CSAwallace_cska32_u_cska64_and_propagate1134;
  assign u_CSAwallace_cska32_u_cska64_mux2to111_and0 = u_CSAwallace_cska32_u_cska64_mux2to110_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate1135;
  assign u_CSAwallace_cska32_u_cska64_mux2to111_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate1135;
  assign u_CSAwallace_cska32_u_cska64_mux2to111_and1 = u_CSAwallace_cska32_u_cska64_fa46_or0 & u_CSAwallace_cska32_u_cska64_mux2to111_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to111_xor0 = u_CSAwallace_cska32_u_cska64_mux2to111_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to111_and1;
  assign u_CSAwallace_cska32_u_cska64_xor48 = u_CSAwallace_cska32_csa29_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_u_cska64_fa47_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa48_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_u_cska64_fa47_and0 = u_CSAwallace_cska32_csa29_csa_component_fa48_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa47_or0;
  assign u_CSAwallace_cska32_u_cska64_fa47_xor1 = u_CSAwallace_cska32_u_cska64_fa47_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to111_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa47_and1 = u_CSAwallace_cska32_u_cska64_fa47_xor0 & u_CSAwallace_cska32_u_cska64_mux2to111_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa47_or0 = u_CSAwallace_cska32_u_cska64_fa47_and0 | u_CSAwallace_cska32_u_cska64_fa47_and1;
  assign u_CSAwallace_cska32_u_cska64_xor49 = u_CSAwallace_cska32_csa29_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_u_cska64_fa48_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa49_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_u_cska64_fa48_and0 = u_CSAwallace_cska32_csa29_csa_component_fa49_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa48_or0;
  assign u_CSAwallace_cska32_u_cska64_fa48_xor1 = u_CSAwallace_cska32_u_cska64_fa48_xor0 ^ u_CSAwallace_cska32_u_cska64_fa47_or0;
  assign u_CSAwallace_cska32_u_cska64_fa48_and1 = u_CSAwallace_cska32_u_cska64_fa48_xor0 & u_CSAwallace_cska32_u_cska64_fa47_or0;
  assign u_CSAwallace_cska32_u_cska64_fa48_or0 = u_CSAwallace_cska32_u_cska64_fa48_and0 | u_CSAwallace_cska32_u_cska64_fa48_and1;
  assign u_CSAwallace_cska32_u_cska64_xor50 = u_CSAwallace_cska32_csa29_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_u_cska64_fa49_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa50_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_u_cska64_fa49_and0 = u_CSAwallace_cska32_csa29_csa_component_fa50_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa49_or0;
  assign u_CSAwallace_cska32_u_cska64_fa49_xor1 = u_CSAwallace_cska32_u_cska64_fa49_xor0 ^ u_CSAwallace_cska32_u_cska64_fa48_or0;
  assign u_CSAwallace_cska32_u_cska64_fa49_and1 = u_CSAwallace_cska32_u_cska64_fa49_xor0 & u_CSAwallace_cska32_u_cska64_fa48_or0;
  assign u_CSAwallace_cska32_u_cska64_fa49_or0 = u_CSAwallace_cska32_u_cska64_fa49_and0 | u_CSAwallace_cska32_u_cska64_fa49_and1;
  assign u_CSAwallace_cska32_u_cska64_xor51 = u_CSAwallace_cska32_csa29_csa_component_fa51_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_u_cska64_fa50_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa51_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_u_cska64_fa50_and0 = u_CSAwallace_cska32_csa29_csa_component_fa51_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa50_or0;
  assign u_CSAwallace_cska32_u_cska64_fa50_xor1 = u_CSAwallace_cska32_u_cska64_fa50_xor0 ^ u_CSAwallace_cska32_u_cska64_fa49_or0;
  assign u_CSAwallace_cska32_u_cska64_fa50_and1 = u_CSAwallace_cska32_u_cska64_fa50_xor0 & u_CSAwallace_cska32_u_cska64_fa49_or0;
  assign u_CSAwallace_cska32_u_cska64_fa50_or0 = u_CSAwallace_cska32_u_cska64_fa50_and0 | u_CSAwallace_cska32_u_cska64_fa50_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1236 = u_CSAwallace_cska32_u_cska64_xor48 & u_CSAwallace_cska32_u_cska64_xor50;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1237 = u_CSAwallace_cska32_u_cska64_xor49 & u_CSAwallace_cska32_u_cska64_xor51;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1238 = u_CSAwallace_cska32_u_cska64_and_propagate1236 & u_CSAwallace_cska32_u_cska64_and_propagate1237;
  assign u_CSAwallace_cska32_u_cska64_mux2to112_and0 = u_CSAwallace_cska32_u_cska64_mux2to111_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate1238;
  assign u_CSAwallace_cska32_u_cska64_mux2to112_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate1238;
  assign u_CSAwallace_cska32_u_cska64_mux2to112_and1 = u_CSAwallace_cska32_u_cska64_fa50_or0 & u_CSAwallace_cska32_u_cska64_mux2to112_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to112_xor0 = u_CSAwallace_cska32_u_cska64_mux2to112_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to112_and1;
  assign u_CSAwallace_cska32_u_cska64_xor52 = u_CSAwallace_cska32_csa29_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_u_cska64_fa51_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa52_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_u_cska64_fa51_and0 = u_CSAwallace_cska32_csa29_csa_component_fa52_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa51_or0;
  assign u_CSAwallace_cska32_u_cska64_fa51_xor1 = u_CSAwallace_cska32_u_cska64_fa51_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to112_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa51_and1 = u_CSAwallace_cska32_u_cska64_fa51_xor0 & u_CSAwallace_cska32_u_cska64_mux2to112_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa51_or0 = u_CSAwallace_cska32_u_cska64_fa51_and0 | u_CSAwallace_cska32_u_cska64_fa51_and1;
  assign u_CSAwallace_cska32_u_cska64_xor53 = u_CSAwallace_cska32_csa29_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_u_cska64_fa52_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa53_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_u_cska64_fa52_and0 = u_CSAwallace_cska32_csa29_csa_component_fa53_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa52_or0;
  assign u_CSAwallace_cska32_u_cska64_fa52_xor1 = u_CSAwallace_cska32_u_cska64_fa52_xor0 ^ u_CSAwallace_cska32_u_cska64_fa51_or0;
  assign u_CSAwallace_cska32_u_cska64_fa52_and1 = u_CSAwallace_cska32_u_cska64_fa52_xor0 & u_CSAwallace_cska32_u_cska64_fa51_or0;
  assign u_CSAwallace_cska32_u_cska64_fa52_or0 = u_CSAwallace_cska32_u_cska64_fa52_and0 | u_CSAwallace_cska32_u_cska64_fa52_and1;
  assign u_CSAwallace_cska32_u_cska64_xor54 = u_CSAwallace_cska32_csa29_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_u_cska64_fa53_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa54_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_u_cska64_fa53_and0 = u_CSAwallace_cska32_csa29_csa_component_fa54_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa53_or0;
  assign u_CSAwallace_cska32_u_cska64_fa53_xor1 = u_CSAwallace_cska32_u_cska64_fa53_xor0 ^ u_CSAwallace_cska32_u_cska64_fa52_or0;
  assign u_CSAwallace_cska32_u_cska64_fa53_and1 = u_CSAwallace_cska32_u_cska64_fa53_xor0 & u_CSAwallace_cska32_u_cska64_fa52_or0;
  assign u_CSAwallace_cska32_u_cska64_fa53_or0 = u_CSAwallace_cska32_u_cska64_fa53_and0 | u_CSAwallace_cska32_u_cska64_fa53_and1;
  assign u_CSAwallace_cska32_u_cska64_xor55 = u_CSAwallace_cska32_csa29_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_u_cska64_fa54_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa55_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_u_cska64_fa54_and0 = u_CSAwallace_cska32_csa29_csa_component_fa55_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa54_or0;
  assign u_CSAwallace_cska32_u_cska64_fa54_xor1 = u_CSAwallace_cska32_u_cska64_fa54_xor0 ^ u_CSAwallace_cska32_u_cska64_fa53_or0;
  assign u_CSAwallace_cska32_u_cska64_fa54_and1 = u_CSAwallace_cska32_u_cska64_fa54_xor0 & u_CSAwallace_cska32_u_cska64_fa53_or0;
  assign u_CSAwallace_cska32_u_cska64_fa54_or0 = u_CSAwallace_cska32_u_cska64_fa54_and0 | u_CSAwallace_cska32_u_cska64_fa54_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1339 = u_CSAwallace_cska32_u_cska64_xor52 & u_CSAwallace_cska32_u_cska64_xor54;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1340 = u_CSAwallace_cska32_u_cska64_xor53 & u_CSAwallace_cska32_u_cska64_xor55;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1341 = u_CSAwallace_cska32_u_cska64_and_propagate1339 & u_CSAwallace_cska32_u_cska64_and_propagate1340;
  assign u_CSAwallace_cska32_u_cska64_mux2to113_and0 = u_CSAwallace_cska32_u_cska64_mux2to112_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate1341;
  assign u_CSAwallace_cska32_u_cska64_mux2to113_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate1341;
  assign u_CSAwallace_cska32_u_cska64_mux2to113_and1 = u_CSAwallace_cska32_u_cska64_fa54_or0 & u_CSAwallace_cska32_u_cska64_mux2to113_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to113_xor0 = u_CSAwallace_cska32_u_cska64_mux2to113_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to113_and1;
  assign u_CSAwallace_cska32_u_cska64_xor56 = u_CSAwallace_cska32_csa29_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_u_cska64_fa55_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa56_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_u_cska64_fa55_and0 = u_CSAwallace_cska32_csa29_csa_component_fa56_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa55_or0;
  assign u_CSAwallace_cska32_u_cska64_fa55_xor1 = u_CSAwallace_cska32_u_cska64_fa55_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to113_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa55_and1 = u_CSAwallace_cska32_u_cska64_fa55_xor0 & u_CSAwallace_cska32_u_cska64_mux2to113_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa55_or0 = u_CSAwallace_cska32_u_cska64_fa55_and0 | u_CSAwallace_cska32_u_cska64_fa55_and1;
  assign u_CSAwallace_cska32_u_cska64_xor57 = u_CSAwallace_cska32_csa29_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_u_cska64_fa56_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa57_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_u_cska64_fa56_and0 = u_CSAwallace_cska32_csa29_csa_component_fa57_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa56_or0;
  assign u_CSAwallace_cska32_u_cska64_fa56_xor1 = u_CSAwallace_cska32_u_cska64_fa56_xor0 ^ u_CSAwallace_cska32_u_cska64_fa55_or0;
  assign u_CSAwallace_cska32_u_cska64_fa56_and1 = u_CSAwallace_cska32_u_cska64_fa56_xor0 & u_CSAwallace_cska32_u_cska64_fa55_or0;
  assign u_CSAwallace_cska32_u_cska64_fa56_or0 = u_CSAwallace_cska32_u_cska64_fa56_and0 | u_CSAwallace_cska32_u_cska64_fa56_and1;
  assign u_CSAwallace_cska32_u_cska64_xor58 = u_CSAwallace_cska32_csa29_csa_component_fa58_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_u_cska64_fa57_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa58_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_u_cska64_fa57_and0 = u_CSAwallace_cska32_csa29_csa_component_fa58_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa57_or0;
  assign u_CSAwallace_cska32_u_cska64_fa57_xor1 = u_CSAwallace_cska32_u_cska64_fa57_xor0 ^ u_CSAwallace_cska32_u_cska64_fa56_or0;
  assign u_CSAwallace_cska32_u_cska64_fa57_and1 = u_CSAwallace_cska32_u_cska64_fa57_xor0 & u_CSAwallace_cska32_u_cska64_fa56_or0;
  assign u_CSAwallace_cska32_u_cska64_fa57_or0 = u_CSAwallace_cska32_u_cska64_fa57_and0 | u_CSAwallace_cska32_u_cska64_fa57_and1;
  assign u_CSAwallace_cska32_u_cska64_xor59 = u_CSAwallace_cska32_csa29_csa_component_fa59_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_u_cska64_fa58_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa59_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_u_cska64_fa58_and0 = u_CSAwallace_cska32_csa29_csa_component_fa59_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa58_or0;
  assign u_CSAwallace_cska32_u_cska64_fa58_xor1 = u_CSAwallace_cska32_u_cska64_fa58_xor0 ^ u_CSAwallace_cska32_u_cska64_fa57_or0;
  assign u_CSAwallace_cska32_u_cska64_fa58_and1 = u_CSAwallace_cska32_u_cska64_fa58_xor0 & u_CSAwallace_cska32_u_cska64_fa57_or0;
  assign u_CSAwallace_cska32_u_cska64_fa58_or0 = u_CSAwallace_cska32_u_cska64_fa58_and0 | u_CSAwallace_cska32_u_cska64_fa58_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1442 = u_CSAwallace_cska32_u_cska64_xor56 & u_CSAwallace_cska32_u_cska64_xor58;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1443 = u_CSAwallace_cska32_u_cska64_xor57 & u_CSAwallace_cska32_u_cska64_xor59;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1444 = u_CSAwallace_cska32_u_cska64_and_propagate1442 & u_CSAwallace_cska32_u_cska64_and_propagate1443;
  assign u_CSAwallace_cska32_u_cska64_mux2to114_and0 = u_CSAwallace_cska32_u_cska64_mux2to113_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate1444;
  assign u_CSAwallace_cska32_u_cska64_mux2to114_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate1444;
  assign u_CSAwallace_cska32_u_cska64_mux2to114_and1 = u_CSAwallace_cska32_u_cska64_fa58_or0 & u_CSAwallace_cska32_u_cska64_mux2to114_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to114_xor0 = u_CSAwallace_cska32_u_cska64_mux2to114_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to114_and1;
  assign u_CSAwallace_cska32_u_cska64_xor60 = u_CSAwallace_cska32_csa29_csa_component_fa60_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa59_or0;
  assign u_CSAwallace_cska32_u_cska64_fa59_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa60_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa59_or0;
  assign u_CSAwallace_cska32_u_cska64_fa59_and0 = u_CSAwallace_cska32_csa29_csa_component_fa60_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa59_or0;
  assign u_CSAwallace_cska32_u_cska64_fa59_xor1 = u_CSAwallace_cska32_u_cska64_fa59_xor0 ^ u_CSAwallace_cska32_u_cska64_mux2to114_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa59_and1 = u_CSAwallace_cska32_u_cska64_fa59_xor0 & u_CSAwallace_cska32_u_cska64_mux2to114_xor0;
  assign u_CSAwallace_cska32_u_cska64_fa59_or0 = u_CSAwallace_cska32_u_cska64_fa59_and0 | u_CSAwallace_cska32_u_cska64_fa59_and1;
  assign u_CSAwallace_cska32_u_cska64_xor61 = u_CSAwallace_cska32_csa29_csa_component_fa61_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa60_or0;
  assign u_CSAwallace_cska32_u_cska64_fa60_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa61_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa60_or0;
  assign u_CSAwallace_cska32_u_cska64_fa60_and0 = u_CSAwallace_cska32_csa29_csa_component_fa61_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa60_or0;
  assign u_CSAwallace_cska32_u_cska64_fa60_xor1 = u_CSAwallace_cska32_u_cska64_fa60_xor0 ^ u_CSAwallace_cska32_u_cska64_fa59_or0;
  assign u_CSAwallace_cska32_u_cska64_fa60_and1 = u_CSAwallace_cska32_u_cska64_fa60_xor0 & u_CSAwallace_cska32_u_cska64_fa59_or0;
  assign u_CSAwallace_cska32_u_cska64_fa60_or0 = u_CSAwallace_cska32_u_cska64_fa60_and0 | u_CSAwallace_cska32_u_cska64_fa60_and1;
  assign u_CSAwallace_cska32_u_cska64_xor62 = u_CSAwallace_cska32_csa29_csa_component_fa62_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa61_or0;
  assign u_CSAwallace_cska32_u_cska64_fa61_xor0 = u_CSAwallace_cska32_csa29_csa_component_fa62_xor1 ^ u_CSAwallace_cska32_csa29_csa_component_fa61_or0;
  assign u_CSAwallace_cska32_u_cska64_fa61_and0 = u_CSAwallace_cska32_csa29_csa_component_fa62_xor1 & u_CSAwallace_cska32_csa29_csa_component_fa61_or0;
  assign u_CSAwallace_cska32_u_cska64_fa61_xor1 = u_CSAwallace_cska32_u_cska64_fa61_xor0 ^ u_CSAwallace_cska32_u_cska64_fa60_or0;
  assign u_CSAwallace_cska32_u_cska64_fa61_and1 = u_CSAwallace_cska32_u_cska64_fa61_xor0 & u_CSAwallace_cska32_u_cska64_fa60_or0;
  assign u_CSAwallace_cska32_u_cska64_fa61_or0 = u_CSAwallace_cska32_u_cska64_fa61_and0 | u_CSAwallace_cska32_u_cska64_fa61_and1;
  assign u_CSAwallace_cska32_u_cska64_fa62_xor1 = u_CSAwallace_cska32_csa29_csa_component_fa62_and1 ^ u_CSAwallace_cska32_u_cska64_fa61_or0;
  assign u_CSAwallace_cska32_u_cska64_fa62_and1 = u_CSAwallace_cska32_csa29_csa_component_fa62_and1 & u_CSAwallace_cska32_u_cska64_fa61_or0;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1545 = u_CSAwallace_cska32_u_cska64_xor60 & u_CSAwallace_cska32_u_cska64_xor62;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1546 = u_CSAwallace_cska32_u_cska64_xor61 & u_CSAwallace_cska32_csa29_csa_component_fa62_and1;
  assign u_CSAwallace_cska32_u_cska64_and_propagate1547 = u_CSAwallace_cska32_u_cska64_and_propagate1545 & u_CSAwallace_cska32_u_cska64_and_propagate1546;
  assign u_CSAwallace_cska32_u_cska64_mux2to115_and0 = u_CSAwallace_cska32_u_cska64_mux2to114_xor0 & u_CSAwallace_cska32_u_cska64_and_propagate1547;
  assign u_CSAwallace_cska32_u_cska64_mux2to115_not0 = ~u_CSAwallace_cska32_u_cska64_and_propagate1547;
  assign u_CSAwallace_cska32_u_cska64_mux2to115_and1 = u_CSAwallace_cska32_u_cska64_fa62_and1 & u_CSAwallace_cska32_u_cska64_mux2to115_not0;
  assign u_CSAwallace_cska32_u_cska64_mux2to115_xor0 = u_CSAwallace_cska32_u_cska64_mux2to115_and0 ^ u_CSAwallace_cska32_u_cska64_mux2to115_and1;

  assign u_CSAwallace_cska32_out[0] = u_CSAwallace_cska32_and_0_0;
  assign u_CSAwallace_cska32_out[1] = u_CSAwallace_cska32_csa0_csa_component_fa1_xor0;
  assign u_CSAwallace_cska32_out[2] = u_CSAwallace_cska32_csa10_csa_component_fa2_xor0;
  assign u_CSAwallace_cska32_out[3] = u_CSAwallace_cska32_csa17_csa_component_fa3_xor0;
  assign u_CSAwallace_cska32_out[4] = u_CSAwallace_cska32_csa22_csa_component_fa4_xor0;
  assign u_CSAwallace_cska32_out[5] = u_CSAwallace_cska32_csa25_csa_component_fa5_xor0;
  assign u_CSAwallace_cska32_out[6] = u_CSAwallace_cska32_csa27_csa_component_fa6_xor0;
  assign u_CSAwallace_cska32_out[7] = u_CSAwallace_cska32_csa28_csa_component_fa7_xor0;
  assign u_CSAwallace_cska32_out[8] = u_CSAwallace_cska32_csa29_csa_component_fa8_xor0;
  assign u_CSAwallace_cska32_out[9] = u_CSAwallace_cska32_u_cska64_fa8_xor0;
  assign u_CSAwallace_cska32_out[10] = u_CSAwallace_cska32_u_cska64_fa9_xor1;
  assign u_CSAwallace_cska32_out[11] = u_CSAwallace_cska32_u_cska64_fa10_xor1;
  assign u_CSAwallace_cska32_out[12] = u_CSAwallace_cska32_u_cska64_fa11_xor1;
  assign u_CSAwallace_cska32_out[13] = u_CSAwallace_cska32_u_cska64_fa12_xor1;
  assign u_CSAwallace_cska32_out[14] = u_CSAwallace_cska32_u_cska64_fa13_xor1;
  assign u_CSAwallace_cska32_out[15] = u_CSAwallace_cska32_u_cska64_fa14_xor1;
  assign u_CSAwallace_cska32_out[16] = u_CSAwallace_cska32_u_cska64_fa15_xor1;
  assign u_CSAwallace_cska32_out[17] = u_CSAwallace_cska32_u_cska64_fa16_xor1;
  assign u_CSAwallace_cska32_out[18] = u_CSAwallace_cska32_u_cska64_fa17_xor1;
  assign u_CSAwallace_cska32_out[19] = u_CSAwallace_cska32_u_cska64_fa18_xor1;
  assign u_CSAwallace_cska32_out[20] = u_CSAwallace_cska32_u_cska64_fa19_xor1;
  assign u_CSAwallace_cska32_out[21] = u_CSAwallace_cska32_u_cska64_fa20_xor1;
  assign u_CSAwallace_cska32_out[22] = u_CSAwallace_cska32_u_cska64_fa21_xor1;
  assign u_CSAwallace_cska32_out[23] = u_CSAwallace_cska32_u_cska64_fa22_xor1;
  assign u_CSAwallace_cska32_out[24] = u_CSAwallace_cska32_u_cska64_fa23_xor1;
  assign u_CSAwallace_cska32_out[25] = u_CSAwallace_cska32_u_cska64_fa24_xor1;
  assign u_CSAwallace_cska32_out[26] = u_CSAwallace_cska32_u_cska64_fa25_xor1;
  assign u_CSAwallace_cska32_out[27] = u_CSAwallace_cska32_u_cska64_fa26_xor1;
  assign u_CSAwallace_cska32_out[28] = u_CSAwallace_cska32_u_cska64_fa27_xor1;
  assign u_CSAwallace_cska32_out[29] = u_CSAwallace_cska32_u_cska64_fa28_xor1;
  assign u_CSAwallace_cska32_out[30] = u_CSAwallace_cska32_u_cska64_fa29_xor1;
  assign u_CSAwallace_cska32_out[31] = u_CSAwallace_cska32_u_cska64_fa30_xor1;
  assign u_CSAwallace_cska32_out[32] = u_CSAwallace_cska32_u_cska64_fa31_xor1;
  assign u_CSAwallace_cska32_out[33] = u_CSAwallace_cska32_u_cska64_fa32_xor1;
  assign u_CSAwallace_cska32_out[34] = u_CSAwallace_cska32_u_cska64_fa33_xor1;
  assign u_CSAwallace_cska32_out[35] = u_CSAwallace_cska32_u_cska64_fa34_xor1;
  assign u_CSAwallace_cska32_out[36] = u_CSAwallace_cska32_u_cska64_fa35_xor1;
  assign u_CSAwallace_cska32_out[37] = u_CSAwallace_cska32_u_cska64_fa36_xor1;
  assign u_CSAwallace_cska32_out[38] = u_CSAwallace_cska32_u_cska64_fa37_xor1;
  assign u_CSAwallace_cska32_out[39] = u_CSAwallace_cska32_u_cska64_fa38_xor1;
  assign u_CSAwallace_cska32_out[40] = u_CSAwallace_cska32_u_cska64_fa39_xor1;
  assign u_CSAwallace_cska32_out[41] = u_CSAwallace_cska32_u_cska64_fa40_xor1;
  assign u_CSAwallace_cska32_out[42] = u_CSAwallace_cska32_u_cska64_fa41_xor1;
  assign u_CSAwallace_cska32_out[43] = u_CSAwallace_cska32_u_cska64_fa42_xor1;
  assign u_CSAwallace_cska32_out[44] = u_CSAwallace_cska32_u_cska64_fa43_xor1;
  assign u_CSAwallace_cska32_out[45] = u_CSAwallace_cska32_u_cska64_fa44_xor1;
  assign u_CSAwallace_cska32_out[46] = u_CSAwallace_cska32_u_cska64_fa45_xor1;
  assign u_CSAwallace_cska32_out[47] = u_CSAwallace_cska32_u_cska64_fa46_xor1;
  assign u_CSAwallace_cska32_out[48] = u_CSAwallace_cska32_u_cska64_fa47_xor1;
  assign u_CSAwallace_cska32_out[49] = u_CSAwallace_cska32_u_cska64_fa48_xor1;
  assign u_CSAwallace_cska32_out[50] = u_CSAwallace_cska32_u_cska64_fa49_xor1;
  assign u_CSAwallace_cska32_out[51] = u_CSAwallace_cska32_u_cska64_fa50_xor1;
  assign u_CSAwallace_cska32_out[52] = u_CSAwallace_cska32_u_cska64_fa51_xor1;
  assign u_CSAwallace_cska32_out[53] = u_CSAwallace_cska32_u_cska64_fa52_xor1;
  assign u_CSAwallace_cska32_out[54] = u_CSAwallace_cska32_u_cska64_fa53_xor1;
  assign u_CSAwallace_cska32_out[55] = u_CSAwallace_cska32_u_cska64_fa54_xor1;
  assign u_CSAwallace_cska32_out[56] = u_CSAwallace_cska32_u_cska64_fa55_xor1;
  assign u_CSAwallace_cska32_out[57] = u_CSAwallace_cska32_u_cska64_fa56_xor1;
  assign u_CSAwallace_cska32_out[58] = u_CSAwallace_cska32_u_cska64_fa57_xor1;
  assign u_CSAwallace_cska32_out[59] = u_CSAwallace_cska32_u_cska64_fa58_xor1;
  assign u_CSAwallace_cska32_out[60] = u_CSAwallace_cska32_u_cska64_fa59_xor1;
  assign u_CSAwallace_cska32_out[61] = u_CSAwallace_cska32_u_cska64_fa60_xor1;
  assign u_CSAwallace_cska32_out[62] = u_CSAwallace_cska32_u_cska64_fa61_xor1;
  assign u_CSAwallace_cska32_out[63] = u_CSAwallace_cska32_u_cska64_fa62_xor1;
endmodule