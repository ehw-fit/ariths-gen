module f_u_arrmul24(input [23:0] a, input [23:0] b, output [47:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire f_u_arrmul24_and0_0_a_0;
  wire f_u_arrmul24_and0_0_b_0;
  wire f_u_arrmul24_and0_0_y0;
  wire f_u_arrmul24_and1_0_a_1;
  wire f_u_arrmul24_and1_0_b_0;
  wire f_u_arrmul24_and1_0_y0;
  wire f_u_arrmul24_and2_0_a_2;
  wire f_u_arrmul24_and2_0_b_0;
  wire f_u_arrmul24_and2_0_y0;
  wire f_u_arrmul24_and3_0_a_3;
  wire f_u_arrmul24_and3_0_b_0;
  wire f_u_arrmul24_and3_0_y0;
  wire f_u_arrmul24_and4_0_a_4;
  wire f_u_arrmul24_and4_0_b_0;
  wire f_u_arrmul24_and4_0_y0;
  wire f_u_arrmul24_and5_0_a_5;
  wire f_u_arrmul24_and5_0_b_0;
  wire f_u_arrmul24_and5_0_y0;
  wire f_u_arrmul24_and6_0_a_6;
  wire f_u_arrmul24_and6_0_b_0;
  wire f_u_arrmul24_and6_0_y0;
  wire f_u_arrmul24_and7_0_a_7;
  wire f_u_arrmul24_and7_0_b_0;
  wire f_u_arrmul24_and7_0_y0;
  wire f_u_arrmul24_and8_0_a_8;
  wire f_u_arrmul24_and8_0_b_0;
  wire f_u_arrmul24_and8_0_y0;
  wire f_u_arrmul24_and9_0_a_9;
  wire f_u_arrmul24_and9_0_b_0;
  wire f_u_arrmul24_and9_0_y0;
  wire f_u_arrmul24_and10_0_a_10;
  wire f_u_arrmul24_and10_0_b_0;
  wire f_u_arrmul24_and10_0_y0;
  wire f_u_arrmul24_and11_0_a_11;
  wire f_u_arrmul24_and11_0_b_0;
  wire f_u_arrmul24_and11_0_y0;
  wire f_u_arrmul24_and12_0_a_12;
  wire f_u_arrmul24_and12_0_b_0;
  wire f_u_arrmul24_and12_0_y0;
  wire f_u_arrmul24_and13_0_a_13;
  wire f_u_arrmul24_and13_0_b_0;
  wire f_u_arrmul24_and13_0_y0;
  wire f_u_arrmul24_and14_0_a_14;
  wire f_u_arrmul24_and14_0_b_0;
  wire f_u_arrmul24_and14_0_y0;
  wire f_u_arrmul24_and15_0_a_15;
  wire f_u_arrmul24_and15_0_b_0;
  wire f_u_arrmul24_and15_0_y0;
  wire f_u_arrmul24_and16_0_a_16;
  wire f_u_arrmul24_and16_0_b_0;
  wire f_u_arrmul24_and16_0_y0;
  wire f_u_arrmul24_and17_0_a_17;
  wire f_u_arrmul24_and17_0_b_0;
  wire f_u_arrmul24_and17_0_y0;
  wire f_u_arrmul24_and18_0_a_18;
  wire f_u_arrmul24_and18_0_b_0;
  wire f_u_arrmul24_and18_0_y0;
  wire f_u_arrmul24_and19_0_a_19;
  wire f_u_arrmul24_and19_0_b_0;
  wire f_u_arrmul24_and19_0_y0;
  wire f_u_arrmul24_and20_0_a_20;
  wire f_u_arrmul24_and20_0_b_0;
  wire f_u_arrmul24_and20_0_y0;
  wire f_u_arrmul24_and21_0_a_21;
  wire f_u_arrmul24_and21_0_b_0;
  wire f_u_arrmul24_and21_0_y0;
  wire f_u_arrmul24_and22_0_a_22;
  wire f_u_arrmul24_and22_0_b_0;
  wire f_u_arrmul24_and22_0_y0;
  wire f_u_arrmul24_and23_0_a_23;
  wire f_u_arrmul24_and23_0_b_0;
  wire f_u_arrmul24_and23_0_y0;
  wire f_u_arrmul24_and0_1_a_0;
  wire f_u_arrmul24_and0_1_b_1;
  wire f_u_arrmul24_and0_1_y0;
  wire f_u_arrmul24_ha0_1_f_u_arrmul24_and0_1_y0;
  wire f_u_arrmul24_ha0_1_f_u_arrmul24_and1_0_y0;
  wire f_u_arrmul24_ha0_1_y0;
  wire f_u_arrmul24_ha0_1_y1;
  wire f_u_arrmul24_and1_1_a_1;
  wire f_u_arrmul24_and1_1_b_1;
  wire f_u_arrmul24_and1_1_y0;
  wire f_u_arrmul24_fa1_1_f_u_arrmul24_and1_1_y0;
  wire f_u_arrmul24_fa1_1_f_u_arrmul24_and2_0_y0;
  wire f_u_arrmul24_fa1_1_y0;
  wire f_u_arrmul24_fa1_1_y1;
  wire f_u_arrmul24_fa1_1_f_u_arrmul24_ha0_1_y1;
  wire f_u_arrmul24_fa1_1_y2;
  wire f_u_arrmul24_fa1_1_y3;
  wire f_u_arrmul24_fa1_1_y4;
  wire f_u_arrmul24_and2_1_a_2;
  wire f_u_arrmul24_and2_1_b_1;
  wire f_u_arrmul24_and2_1_y0;
  wire f_u_arrmul24_fa2_1_f_u_arrmul24_and2_1_y0;
  wire f_u_arrmul24_fa2_1_f_u_arrmul24_and3_0_y0;
  wire f_u_arrmul24_fa2_1_y0;
  wire f_u_arrmul24_fa2_1_y1;
  wire f_u_arrmul24_fa2_1_f_u_arrmul24_fa1_1_y4;
  wire f_u_arrmul24_fa2_1_y2;
  wire f_u_arrmul24_fa2_1_y3;
  wire f_u_arrmul24_fa2_1_y4;
  wire f_u_arrmul24_and3_1_a_3;
  wire f_u_arrmul24_and3_1_b_1;
  wire f_u_arrmul24_and3_1_y0;
  wire f_u_arrmul24_fa3_1_f_u_arrmul24_and3_1_y0;
  wire f_u_arrmul24_fa3_1_f_u_arrmul24_and4_0_y0;
  wire f_u_arrmul24_fa3_1_y0;
  wire f_u_arrmul24_fa3_1_y1;
  wire f_u_arrmul24_fa3_1_f_u_arrmul24_fa2_1_y4;
  wire f_u_arrmul24_fa3_1_y2;
  wire f_u_arrmul24_fa3_1_y3;
  wire f_u_arrmul24_fa3_1_y4;
  wire f_u_arrmul24_and4_1_a_4;
  wire f_u_arrmul24_and4_1_b_1;
  wire f_u_arrmul24_and4_1_y0;
  wire f_u_arrmul24_fa4_1_f_u_arrmul24_and4_1_y0;
  wire f_u_arrmul24_fa4_1_f_u_arrmul24_and5_0_y0;
  wire f_u_arrmul24_fa4_1_y0;
  wire f_u_arrmul24_fa4_1_y1;
  wire f_u_arrmul24_fa4_1_f_u_arrmul24_fa3_1_y4;
  wire f_u_arrmul24_fa4_1_y2;
  wire f_u_arrmul24_fa4_1_y3;
  wire f_u_arrmul24_fa4_1_y4;
  wire f_u_arrmul24_and5_1_a_5;
  wire f_u_arrmul24_and5_1_b_1;
  wire f_u_arrmul24_and5_1_y0;
  wire f_u_arrmul24_fa5_1_f_u_arrmul24_and5_1_y0;
  wire f_u_arrmul24_fa5_1_f_u_arrmul24_and6_0_y0;
  wire f_u_arrmul24_fa5_1_y0;
  wire f_u_arrmul24_fa5_1_y1;
  wire f_u_arrmul24_fa5_1_f_u_arrmul24_fa4_1_y4;
  wire f_u_arrmul24_fa5_1_y2;
  wire f_u_arrmul24_fa5_1_y3;
  wire f_u_arrmul24_fa5_1_y4;
  wire f_u_arrmul24_and6_1_a_6;
  wire f_u_arrmul24_and6_1_b_1;
  wire f_u_arrmul24_and6_1_y0;
  wire f_u_arrmul24_fa6_1_f_u_arrmul24_and6_1_y0;
  wire f_u_arrmul24_fa6_1_f_u_arrmul24_and7_0_y0;
  wire f_u_arrmul24_fa6_1_y0;
  wire f_u_arrmul24_fa6_1_y1;
  wire f_u_arrmul24_fa6_1_f_u_arrmul24_fa5_1_y4;
  wire f_u_arrmul24_fa6_1_y2;
  wire f_u_arrmul24_fa6_1_y3;
  wire f_u_arrmul24_fa6_1_y4;
  wire f_u_arrmul24_and7_1_a_7;
  wire f_u_arrmul24_and7_1_b_1;
  wire f_u_arrmul24_and7_1_y0;
  wire f_u_arrmul24_fa7_1_f_u_arrmul24_and7_1_y0;
  wire f_u_arrmul24_fa7_1_f_u_arrmul24_and8_0_y0;
  wire f_u_arrmul24_fa7_1_y0;
  wire f_u_arrmul24_fa7_1_y1;
  wire f_u_arrmul24_fa7_1_f_u_arrmul24_fa6_1_y4;
  wire f_u_arrmul24_fa7_1_y2;
  wire f_u_arrmul24_fa7_1_y3;
  wire f_u_arrmul24_fa7_1_y4;
  wire f_u_arrmul24_and8_1_a_8;
  wire f_u_arrmul24_and8_1_b_1;
  wire f_u_arrmul24_and8_1_y0;
  wire f_u_arrmul24_fa8_1_f_u_arrmul24_and8_1_y0;
  wire f_u_arrmul24_fa8_1_f_u_arrmul24_and9_0_y0;
  wire f_u_arrmul24_fa8_1_y0;
  wire f_u_arrmul24_fa8_1_y1;
  wire f_u_arrmul24_fa8_1_f_u_arrmul24_fa7_1_y4;
  wire f_u_arrmul24_fa8_1_y2;
  wire f_u_arrmul24_fa8_1_y3;
  wire f_u_arrmul24_fa8_1_y4;
  wire f_u_arrmul24_and9_1_a_9;
  wire f_u_arrmul24_and9_1_b_1;
  wire f_u_arrmul24_and9_1_y0;
  wire f_u_arrmul24_fa9_1_f_u_arrmul24_and9_1_y0;
  wire f_u_arrmul24_fa9_1_f_u_arrmul24_and10_0_y0;
  wire f_u_arrmul24_fa9_1_y0;
  wire f_u_arrmul24_fa9_1_y1;
  wire f_u_arrmul24_fa9_1_f_u_arrmul24_fa8_1_y4;
  wire f_u_arrmul24_fa9_1_y2;
  wire f_u_arrmul24_fa9_1_y3;
  wire f_u_arrmul24_fa9_1_y4;
  wire f_u_arrmul24_and10_1_a_10;
  wire f_u_arrmul24_and10_1_b_1;
  wire f_u_arrmul24_and10_1_y0;
  wire f_u_arrmul24_fa10_1_f_u_arrmul24_and10_1_y0;
  wire f_u_arrmul24_fa10_1_f_u_arrmul24_and11_0_y0;
  wire f_u_arrmul24_fa10_1_y0;
  wire f_u_arrmul24_fa10_1_y1;
  wire f_u_arrmul24_fa10_1_f_u_arrmul24_fa9_1_y4;
  wire f_u_arrmul24_fa10_1_y2;
  wire f_u_arrmul24_fa10_1_y3;
  wire f_u_arrmul24_fa10_1_y4;
  wire f_u_arrmul24_and11_1_a_11;
  wire f_u_arrmul24_and11_1_b_1;
  wire f_u_arrmul24_and11_1_y0;
  wire f_u_arrmul24_fa11_1_f_u_arrmul24_and11_1_y0;
  wire f_u_arrmul24_fa11_1_f_u_arrmul24_and12_0_y0;
  wire f_u_arrmul24_fa11_1_y0;
  wire f_u_arrmul24_fa11_1_y1;
  wire f_u_arrmul24_fa11_1_f_u_arrmul24_fa10_1_y4;
  wire f_u_arrmul24_fa11_1_y2;
  wire f_u_arrmul24_fa11_1_y3;
  wire f_u_arrmul24_fa11_1_y4;
  wire f_u_arrmul24_and12_1_a_12;
  wire f_u_arrmul24_and12_1_b_1;
  wire f_u_arrmul24_and12_1_y0;
  wire f_u_arrmul24_fa12_1_f_u_arrmul24_and12_1_y0;
  wire f_u_arrmul24_fa12_1_f_u_arrmul24_and13_0_y0;
  wire f_u_arrmul24_fa12_1_y0;
  wire f_u_arrmul24_fa12_1_y1;
  wire f_u_arrmul24_fa12_1_f_u_arrmul24_fa11_1_y4;
  wire f_u_arrmul24_fa12_1_y2;
  wire f_u_arrmul24_fa12_1_y3;
  wire f_u_arrmul24_fa12_1_y4;
  wire f_u_arrmul24_and13_1_a_13;
  wire f_u_arrmul24_and13_1_b_1;
  wire f_u_arrmul24_and13_1_y0;
  wire f_u_arrmul24_fa13_1_f_u_arrmul24_and13_1_y0;
  wire f_u_arrmul24_fa13_1_f_u_arrmul24_and14_0_y0;
  wire f_u_arrmul24_fa13_1_y0;
  wire f_u_arrmul24_fa13_1_y1;
  wire f_u_arrmul24_fa13_1_f_u_arrmul24_fa12_1_y4;
  wire f_u_arrmul24_fa13_1_y2;
  wire f_u_arrmul24_fa13_1_y3;
  wire f_u_arrmul24_fa13_1_y4;
  wire f_u_arrmul24_and14_1_a_14;
  wire f_u_arrmul24_and14_1_b_1;
  wire f_u_arrmul24_and14_1_y0;
  wire f_u_arrmul24_fa14_1_f_u_arrmul24_and14_1_y0;
  wire f_u_arrmul24_fa14_1_f_u_arrmul24_and15_0_y0;
  wire f_u_arrmul24_fa14_1_y0;
  wire f_u_arrmul24_fa14_1_y1;
  wire f_u_arrmul24_fa14_1_f_u_arrmul24_fa13_1_y4;
  wire f_u_arrmul24_fa14_1_y2;
  wire f_u_arrmul24_fa14_1_y3;
  wire f_u_arrmul24_fa14_1_y4;
  wire f_u_arrmul24_and15_1_a_15;
  wire f_u_arrmul24_and15_1_b_1;
  wire f_u_arrmul24_and15_1_y0;
  wire f_u_arrmul24_fa15_1_f_u_arrmul24_and15_1_y0;
  wire f_u_arrmul24_fa15_1_f_u_arrmul24_and16_0_y0;
  wire f_u_arrmul24_fa15_1_y0;
  wire f_u_arrmul24_fa15_1_y1;
  wire f_u_arrmul24_fa15_1_f_u_arrmul24_fa14_1_y4;
  wire f_u_arrmul24_fa15_1_y2;
  wire f_u_arrmul24_fa15_1_y3;
  wire f_u_arrmul24_fa15_1_y4;
  wire f_u_arrmul24_and16_1_a_16;
  wire f_u_arrmul24_and16_1_b_1;
  wire f_u_arrmul24_and16_1_y0;
  wire f_u_arrmul24_fa16_1_f_u_arrmul24_and16_1_y0;
  wire f_u_arrmul24_fa16_1_f_u_arrmul24_and17_0_y0;
  wire f_u_arrmul24_fa16_1_y0;
  wire f_u_arrmul24_fa16_1_y1;
  wire f_u_arrmul24_fa16_1_f_u_arrmul24_fa15_1_y4;
  wire f_u_arrmul24_fa16_1_y2;
  wire f_u_arrmul24_fa16_1_y3;
  wire f_u_arrmul24_fa16_1_y4;
  wire f_u_arrmul24_and17_1_a_17;
  wire f_u_arrmul24_and17_1_b_1;
  wire f_u_arrmul24_and17_1_y0;
  wire f_u_arrmul24_fa17_1_f_u_arrmul24_and17_1_y0;
  wire f_u_arrmul24_fa17_1_f_u_arrmul24_and18_0_y0;
  wire f_u_arrmul24_fa17_1_y0;
  wire f_u_arrmul24_fa17_1_y1;
  wire f_u_arrmul24_fa17_1_f_u_arrmul24_fa16_1_y4;
  wire f_u_arrmul24_fa17_1_y2;
  wire f_u_arrmul24_fa17_1_y3;
  wire f_u_arrmul24_fa17_1_y4;
  wire f_u_arrmul24_and18_1_a_18;
  wire f_u_arrmul24_and18_1_b_1;
  wire f_u_arrmul24_and18_1_y0;
  wire f_u_arrmul24_fa18_1_f_u_arrmul24_and18_1_y0;
  wire f_u_arrmul24_fa18_1_f_u_arrmul24_and19_0_y0;
  wire f_u_arrmul24_fa18_1_y0;
  wire f_u_arrmul24_fa18_1_y1;
  wire f_u_arrmul24_fa18_1_f_u_arrmul24_fa17_1_y4;
  wire f_u_arrmul24_fa18_1_y2;
  wire f_u_arrmul24_fa18_1_y3;
  wire f_u_arrmul24_fa18_1_y4;
  wire f_u_arrmul24_and19_1_a_19;
  wire f_u_arrmul24_and19_1_b_1;
  wire f_u_arrmul24_and19_1_y0;
  wire f_u_arrmul24_fa19_1_f_u_arrmul24_and19_1_y0;
  wire f_u_arrmul24_fa19_1_f_u_arrmul24_and20_0_y0;
  wire f_u_arrmul24_fa19_1_y0;
  wire f_u_arrmul24_fa19_1_y1;
  wire f_u_arrmul24_fa19_1_f_u_arrmul24_fa18_1_y4;
  wire f_u_arrmul24_fa19_1_y2;
  wire f_u_arrmul24_fa19_1_y3;
  wire f_u_arrmul24_fa19_1_y4;
  wire f_u_arrmul24_and20_1_a_20;
  wire f_u_arrmul24_and20_1_b_1;
  wire f_u_arrmul24_and20_1_y0;
  wire f_u_arrmul24_fa20_1_f_u_arrmul24_and20_1_y0;
  wire f_u_arrmul24_fa20_1_f_u_arrmul24_and21_0_y0;
  wire f_u_arrmul24_fa20_1_y0;
  wire f_u_arrmul24_fa20_1_y1;
  wire f_u_arrmul24_fa20_1_f_u_arrmul24_fa19_1_y4;
  wire f_u_arrmul24_fa20_1_y2;
  wire f_u_arrmul24_fa20_1_y3;
  wire f_u_arrmul24_fa20_1_y4;
  wire f_u_arrmul24_and21_1_a_21;
  wire f_u_arrmul24_and21_1_b_1;
  wire f_u_arrmul24_and21_1_y0;
  wire f_u_arrmul24_fa21_1_f_u_arrmul24_and21_1_y0;
  wire f_u_arrmul24_fa21_1_f_u_arrmul24_and22_0_y0;
  wire f_u_arrmul24_fa21_1_y0;
  wire f_u_arrmul24_fa21_1_y1;
  wire f_u_arrmul24_fa21_1_f_u_arrmul24_fa20_1_y4;
  wire f_u_arrmul24_fa21_1_y2;
  wire f_u_arrmul24_fa21_1_y3;
  wire f_u_arrmul24_fa21_1_y4;
  wire f_u_arrmul24_and22_1_a_22;
  wire f_u_arrmul24_and22_1_b_1;
  wire f_u_arrmul24_and22_1_y0;
  wire f_u_arrmul24_fa22_1_f_u_arrmul24_and22_1_y0;
  wire f_u_arrmul24_fa22_1_f_u_arrmul24_and23_0_y0;
  wire f_u_arrmul24_fa22_1_y0;
  wire f_u_arrmul24_fa22_1_y1;
  wire f_u_arrmul24_fa22_1_f_u_arrmul24_fa21_1_y4;
  wire f_u_arrmul24_fa22_1_y2;
  wire f_u_arrmul24_fa22_1_y3;
  wire f_u_arrmul24_fa22_1_y4;
  wire f_u_arrmul24_and23_1_a_23;
  wire f_u_arrmul24_and23_1_b_1;
  wire f_u_arrmul24_and23_1_y0;
  wire f_u_arrmul24_ha23_1_f_u_arrmul24_and23_1_y0;
  wire f_u_arrmul24_ha23_1_f_u_arrmul24_fa22_1_y4;
  wire f_u_arrmul24_ha23_1_y0;
  wire f_u_arrmul24_ha23_1_y1;
  wire f_u_arrmul24_and0_2_a_0;
  wire f_u_arrmul24_and0_2_b_2;
  wire f_u_arrmul24_and0_2_y0;
  wire f_u_arrmul24_ha0_2_f_u_arrmul24_and0_2_y0;
  wire f_u_arrmul24_ha0_2_f_u_arrmul24_fa1_1_y2;
  wire f_u_arrmul24_ha0_2_y0;
  wire f_u_arrmul24_ha0_2_y1;
  wire f_u_arrmul24_and1_2_a_1;
  wire f_u_arrmul24_and1_2_b_2;
  wire f_u_arrmul24_and1_2_y0;
  wire f_u_arrmul24_fa1_2_f_u_arrmul24_and1_2_y0;
  wire f_u_arrmul24_fa1_2_f_u_arrmul24_fa2_1_y2;
  wire f_u_arrmul24_fa1_2_y0;
  wire f_u_arrmul24_fa1_2_y1;
  wire f_u_arrmul24_fa1_2_f_u_arrmul24_ha0_2_y1;
  wire f_u_arrmul24_fa1_2_y2;
  wire f_u_arrmul24_fa1_2_y3;
  wire f_u_arrmul24_fa1_2_y4;
  wire f_u_arrmul24_and2_2_a_2;
  wire f_u_arrmul24_and2_2_b_2;
  wire f_u_arrmul24_and2_2_y0;
  wire f_u_arrmul24_fa2_2_f_u_arrmul24_and2_2_y0;
  wire f_u_arrmul24_fa2_2_f_u_arrmul24_fa3_1_y2;
  wire f_u_arrmul24_fa2_2_y0;
  wire f_u_arrmul24_fa2_2_y1;
  wire f_u_arrmul24_fa2_2_f_u_arrmul24_fa1_2_y4;
  wire f_u_arrmul24_fa2_2_y2;
  wire f_u_arrmul24_fa2_2_y3;
  wire f_u_arrmul24_fa2_2_y4;
  wire f_u_arrmul24_and3_2_a_3;
  wire f_u_arrmul24_and3_2_b_2;
  wire f_u_arrmul24_and3_2_y0;
  wire f_u_arrmul24_fa3_2_f_u_arrmul24_and3_2_y0;
  wire f_u_arrmul24_fa3_2_f_u_arrmul24_fa4_1_y2;
  wire f_u_arrmul24_fa3_2_y0;
  wire f_u_arrmul24_fa3_2_y1;
  wire f_u_arrmul24_fa3_2_f_u_arrmul24_fa2_2_y4;
  wire f_u_arrmul24_fa3_2_y2;
  wire f_u_arrmul24_fa3_2_y3;
  wire f_u_arrmul24_fa3_2_y4;
  wire f_u_arrmul24_and4_2_a_4;
  wire f_u_arrmul24_and4_2_b_2;
  wire f_u_arrmul24_and4_2_y0;
  wire f_u_arrmul24_fa4_2_f_u_arrmul24_and4_2_y0;
  wire f_u_arrmul24_fa4_2_f_u_arrmul24_fa5_1_y2;
  wire f_u_arrmul24_fa4_2_y0;
  wire f_u_arrmul24_fa4_2_y1;
  wire f_u_arrmul24_fa4_2_f_u_arrmul24_fa3_2_y4;
  wire f_u_arrmul24_fa4_2_y2;
  wire f_u_arrmul24_fa4_2_y3;
  wire f_u_arrmul24_fa4_2_y4;
  wire f_u_arrmul24_and5_2_a_5;
  wire f_u_arrmul24_and5_2_b_2;
  wire f_u_arrmul24_and5_2_y0;
  wire f_u_arrmul24_fa5_2_f_u_arrmul24_and5_2_y0;
  wire f_u_arrmul24_fa5_2_f_u_arrmul24_fa6_1_y2;
  wire f_u_arrmul24_fa5_2_y0;
  wire f_u_arrmul24_fa5_2_y1;
  wire f_u_arrmul24_fa5_2_f_u_arrmul24_fa4_2_y4;
  wire f_u_arrmul24_fa5_2_y2;
  wire f_u_arrmul24_fa5_2_y3;
  wire f_u_arrmul24_fa5_2_y4;
  wire f_u_arrmul24_and6_2_a_6;
  wire f_u_arrmul24_and6_2_b_2;
  wire f_u_arrmul24_and6_2_y0;
  wire f_u_arrmul24_fa6_2_f_u_arrmul24_and6_2_y0;
  wire f_u_arrmul24_fa6_2_f_u_arrmul24_fa7_1_y2;
  wire f_u_arrmul24_fa6_2_y0;
  wire f_u_arrmul24_fa6_2_y1;
  wire f_u_arrmul24_fa6_2_f_u_arrmul24_fa5_2_y4;
  wire f_u_arrmul24_fa6_2_y2;
  wire f_u_arrmul24_fa6_2_y3;
  wire f_u_arrmul24_fa6_2_y4;
  wire f_u_arrmul24_and7_2_a_7;
  wire f_u_arrmul24_and7_2_b_2;
  wire f_u_arrmul24_and7_2_y0;
  wire f_u_arrmul24_fa7_2_f_u_arrmul24_and7_2_y0;
  wire f_u_arrmul24_fa7_2_f_u_arrmul24_fa8_1_y2;
  wire f_u_arrmul24_fa7_2_y0;
  wire f_u_arrmul24_fa7_2_y1;
  wire f_u_arrmul24_fa7_2_f_u_arrmul24_fa6_2_y4;
  wire f_u_arrmul24_fa7_2_y2;
  wire f_u_arrmul24_fa7_2_y3;
  wire f_u_arrmul24_fa7_2_y4;
  wire f_u_arrmul24_and8_2_a_8;
  wire f_u_arrmul24_and8_2_b_2;
  wire f_u_arrmul24_and8_2_y0;
  wire f_u_arrmul24_fa8_2_f_u_arrmul24_and8_2_y0;
  wire f_u_arrmul24_fa8_2_f_u_arrmul24_fa9_1_y2;
  wire f_u_arrmul24_fa8_2_y0;
  wire f_u_arrmul24_fa8_2_y1;
  wire f_u_arrmul24_fa8_2_f_u_arrmul24_fa7_2_y4;
  wire f_u_arrmul24_fa8_2_y2;
  wire f_u_arrmul24_fa8_2_y3;
  wire f_u_arrmul24_fa8_2_y4;
  wire f_u_arrmul24_and9_2_a_9;
  wire f_u_arrmul24_and9_2_b_2;
  wire f_u_arrmul24_and9_2_y0;
  wire f_u_arrmul24_fa9_2_f_u_arrmul24_and9_2_y0;
  wire f_u_arrmul24_fa9_2_f_u_arrmul24_fa10_1_y2;
  wire f_u_arrmul24_fa9_2_y0;
  wire f_u_arrmul24_fa9_2_y1;
  wire f_u_arrmul24_fa9_2_f_u_arrmul24_fa8_2_y4;
  wire f_u_arrmul24_fa9_2_y2;
  wire f_u_arrmul24_fa9_2_y3;
  wire f_u_arrmul24_fa9_2_y4;
  wire f_u_arrmul24_and10_2_a_10;
  wire f_u_arrmul24_and10_2_b_2;
  wire f_u_arrmul24_and10_2_y0;
  wire f_u_arrmul24_fa10_2_f_u_arrmul24_and10_2_y0;
  wire f_u_arrmul24_fa10_2_f_u_arrmul24_fa11_1_y2;
  wire f_u_arrmul24_fa10_2_y0;
  wire f_u_arrmul24_fa10_2_y1;
  wire f_u_arrmul24_fa10_2_f_u_arrmul24_fa9_2_y4;
  wire f_u_arrmul24_fa10_2_y2;
  wire f_u_arrmul24_fa10_2_y3;
  wire f_u_arrmul24_fa10_2_y4;
  wire f_u_arrmul24_and11_2_a_11;
  wire f_u_arrmul24_and11_2_b_2;
  wire f_u_arrmul24_and11_2_y0;
  wire f_u_arrmul24_fa11_2_f_u_arrmul24_and11_2_y0;
  wire f_u_arrmul24_fa11_2_f_u_arrmul24_fa12_1_y2;
  wire f_u_arrmul24_fa11_2_y0;
  wire f_u_arrmul24_fa11_2_y1;
  wire f_u_arrmul24_fa11_2_f_u_arrmul24_fa10_2_y4;
  wire f_u_arrmul24_fa11_2_y2;
  wire f_u_arrmul24_fa11_2_y3;
  wire f_u_arrmul24_fa11_2_y4;
  wire f_u_arrmul24_and12_2_a_12;
  wire f_u_arrmul24_and12_2_b_2;
  wire f_u_arrmul24_and12_2_y0;
  wire f_u_arrmul24_fa12_2_f_u_arrmul24_and12_2_y0;
  wire f_u_arrmul24_fa12_2_f_u_arrmul24_fa13_1_y2;
  wire f_u_arrmul24_fa12_2_y0;
  wire f_u_arrmul24_fa12_2_y1;
  wire f_u_arrmul24_fa12_2_f_u_arrmul24_fa11_2_y4;
  wire f_u_arrmul24_fa12_2_y2;
  wire f_u_arrmul24_fa12_2_y3;
  wire f_u_arrmul24_fa12_2_y4;
  wire f_u_arrmul24_and13_2_a_13;
  wire f_u_arrmul24_and13_2_b_2;
  wire f_u_arrmul24_and13_2_y0;
  wire f_u_arrmul24_fa13_2_f_u_arrmul24_and13_2_y0;
  wire f_u_arrmul24_fa13_2_f_u_arrmul24_fa14_1_y2;
  wire f_u_arrmul24_fa13_2_y0;
  wire f_u_arrmul24_fa13_2_y1;
  wire f_u_arrmul24_fa13_2_f_u_arrmul24_fa12_2_y4;
  wire f_u_arrmul24_fa13_2_y2;
  wire f_u_arrmul24_fa13_2_y3;
  wire f_u_arrmul24_fa13_2_y4;
  wire f_u_arrmul24_and14_2_a_14;
  wire f_u_arrmul24_and14_2_b_2;
  wire f_u_arrmul24_and14_2_y0;
  wire f_u_arrmul24_fa14_2_f_u_arrmul24_and14_2_y0;
  wire f_u_arrmul24_fa14_2_f_u_arrmul24_fa15_1_y2;
  wire f_u_arrmul24_fa14_2_y0;
  wire f_u_arrmul24_fa14_2_y1;
  wire f_u_arrmul24_fa14_2_f_u_arrmul24_fa13_2_y4;
  wire f_u_arrmul24_fa14_2_y2;
  wire f_u_arrmul24_fa14_2_y3;
  wire f_u_arrmul24_fa14_2_y4;
  wire f_u_arrmul24_and15_2_a_15;
  wire f_u_arrmul24_and15_2_b_2;
  wire f_u_arrmul24_and15_2_y0;
  wire f_u_arrmul24_fa15_2_f_u_arrmul24_and15_2_y0;
  wire f_u_arrmul24_fa15_2_f_u_arrmul24_fa16_1_y2;
  wire f_u_arrmul24_fa15_2_y0;
  wire f_u_arrmul24_fa15_2_y1;
  wire f_u_arrmul24_fa15_2_f_u_arrmul24_fa14_2_y4;
  wire f_u_arrmul24_fa15_2_y2;
  wire f_u_arrmul24_fa15_2_y3;
  wire f_u_arrmul24_fa15_2_y4;
  wire f_u_arrmul24_and16_2_a_16;
  wire f_u_arrmul24_and16_2_b_2;
  wire f_u_arrmul24_and16_2_y0;
  wire f_u_arrmul24_fa16_2_f_u_arrmul24_and16_2_y0;
  wire f_u_arrmul24_fa16_2_f_u_arrmul24_fa17_1_y2;
  wire f_u_arrmul24_fa16_2_y0;
  wire f_u_arrmul24_fa16_2_y1;
  wire f_u_arrmul24_fa16_2_f_u_arrmul24_fa15_2_y4;
  wire f_u_arrmul24_fa16_2_y2;
  wire f_u_arrmul24_fa16_2_y3;
  wire f_u_arrmul24_fa16_2_y4;
  wire f_u_arrmul24_and17_2_a_17;
  wire f_u_arrmul24_and17_2_b_2;
  wire f_u_arrmul24_and17_2_y0;
  wire f_u_arrmul24_fa17_2_f_u_arrmul24_and17_2_y0;
  wire f_u_arrmul24_fa17_2_f_u_arrmul24_fa18_1_y2;
  wire f_u_arrmul24_fa17_2_y0;
  wire f_u_arrmul24_fa17_2_y1;
  wire f_u_arrmul24_fa17_2_f_u_arrmul24_fa16_2_y4;
  wire f_u_arrmul24_fa17_2_y2;
  wire f_u_arrmul24_fa17_2_y3;
  wire f_u_arrmul24_fa17_2_y4;
  wire f_u_arrmul24_and18_2_a_18;
  wire f_u_arrmul24_and18_2_b_2;
  wire f_u_arrmul24_and18_2_y0;
  wire f_u_arrmul24_fa18_2_f_u_arrmul24_and18_2_y0;
  wire f_u_arrmul24_fa18_2_f_u_arrmul24_fa19_1_y2;
  wire f_u_arrmul24_fa18_2_y0;
  wire f_u_arrmul24_fa18_2_y1;
  wire f_u_arrmul24_fa18_2_f_u_arrmul24_fa17_2_y4;
  wire f_u_arrmul24_fa18_2_y2;
  wire f_u_arrmul24_fa18_2_y3;
  wire f_u_arrmul24_fa18_2_y4;
  wire f_u_arrmul24_and19_2_a_19;
  wire f_u_arrmul24_and19_2_b_2;
  wire f_u_arrmul24_and19_2_y0;
  wire f_u_arrmul24_fa19_2_f_u_arrmul24_and19_2_y0;
  wire f_u_arrmul24_fa19_2_f_u_arrmul24_fa20_1_y2;
  wire f_u_arrmul24_fa19_2_y0;
  wire f_u_arrmul24_fa19_2_y1;
  wire f_u_arrmul24_fa19_2_f_u_arrmul24_fa18_2_y4;
  wire f_u_arrmul24_fa19_2_y2;
  wire f_u_arrmul24_fa19_2_y3;
  wire f_u_arrmul24_fa19_2_y4;
  wire f_u_arrmul24_and20_2_a_20;
  wire f_u_arrmul24_and20_2_b_2;
  wire f_u_arrmul24_and20_2_y0;
  wire f_u_arrmul24_fa20_2_f_u_arrmul24_and20_2_y0;
  wire f_u_arrmul24_fa20_2_f_u_arrmul24_fa21_1_y2;
  wire f_u_arrmul24_fa20_2_y0;
  wire f_u_arrmul24_fa20_2_y1;
  wire f_u_arrmul24_fa20_2_f_u_arrmul24_fa19_2_y4;
  wire f_u_arrmul24_fa20_2_y2;
  wire f_u_arrmul24_fa20_2_y3;
  wire f_u_arrmul24_fa20_2_y4;
  wire f_u_arrmul24_and21_2_a_21;
  wire f_u_arrmul24_and21_2_b_2;
  wire f_u_arrmul24_and21_2_y0;
  wire f_u_arrmul24_fa21_2_f_u_arrmul24_and21_2_y0;
  wire f_u_arrmul24_fa21_2_f_u_arrmul24_fa22_1_y2;
  wire f_u_arrmul24_fa21_2_y0;
  wire f_u_arrmul24_fa21_2_y1;
  wire f_u_arrmul24_fa21_2_f_u_arrmul24_fa20_2_y4;
  wire f_u_arrmul24_fa21_2_y2;
  wire f_u_arrmul24_fa21_2_y3;
  wire f_u_arrmul24_fa21_2_y4;
  wire f_u_arrmul24_and22_2_a_22;
  wire f_u_arrmul24_and22_2_b_2;
  wire f_u_arrmul24_and22_2_y0;
  wire f_u_arrmul24_fa22_2_f_u_arrmul24_and22_2_y0;
  wire f_u_arrmul24_fa22_2_f_u_arrmul24_ha23_1_y0;
  wire f_u_arrmul24_fa22_2_y0;
  wire f_u_arrmul24_fa22_2_y1;
  wire f_u_arrmul24_fa22_2_f_u_arrmul24_fa21_2_y4;
  wire f_u_arrmul24_fa22_2_y2;
  wire f_u_arrmul24_fa22_2_y3;
  wire f_u_arrmul24_fa22_2_y4;
  wire f_u_arrmul24_and23_2_a_23;
  wire f_u_arrmul24_and23_2_b_2;
  wire f_u_arrmul24_and23_2_y0;
  wire f_u_arrmul24_fa23_2_f_u_arrmul24_and23_2_y0;
  wire f_u_arrmul24_fa23_2_f_u_arrmul24_ha23_1_y1;
  wire f_u_arrmul24_fa23_2_y0;
  wire f_u_arrmul24_fa23_2_y1;
  wire f_u_arrmul24_fa23_2_f_u_arrmul24_fa22_2_y4;
  wire f_u_arrmul24_fa23_2_y2;
  wire f_u_arrmul24_fa23_2_y3;
  wire f_u_arrmul24_fa23_2_y4;
  wire f_u_arrmul24_and0_3_a_0;
  wire f_u_arrmul24_and0_3_b_3;
  wire f_u_arrmul24_and0_3_y0;
  wire f_u_arrmul24_ha0_3_f_u_arrmul24_and0_3_y0;
  wire f_u_arrmul24_ha0_3_f_u_arrmul24_fa1_2_y2;
  wire f_u_arrmul24_ha0_3_y0;
  wire f_u_arrmul24_ha0_3_y1;
  wire f_u_arrmul24_and1_3_a_1;
  wire f_u_arrmul24_and1_3_b_3;
  wire f_u_arrmul24_and1_3_y0;
  wire f_u_arrmul24_fa1_3_f_u_arrmul24_and1_3_y0;
  wire f_u_arrmul24_fa1_3_f_u_arrmul24_fa2_2_y2;
  wire f_u_arrmul24_fa1_3_y0;
  wire f_u_arrmul24_fa1_3_y1;
  wire f_u_arrmul24_fa1_3_f_u_arrmul24_ha0_3_y1;
  wire f_u_arrmul24_fa1_3_y2;
  wire f_u_arrmul24_fa1_3_y3;
  wire f_u_arrmul24_fa1_3_y4;
  wire f_u_arrmul24_and2_3_a_2;
  wire f_u_arrmul24_and2_3_b_3;
  wire f_u_arrmul24_and2_3_y0;
  wire f_u_arrmul24_fa2_3_f_u_arrmul24_and2_3_y0;
  wire f_u_arrmul24_fa2_3_f_u_arrmul24_fa3_2_y2;
  wire f_u_arrmul24_fa2_3_y0;
  wire f_u_arrmul24_fa2_3_y1;
  wire f_u_arrmul24_fa2_3_f_u_arrmul24_fa1_3_y4;
  wire f_u_arrmul24_fa2_3_y2;
  wire f_u_arrmul24_fa2_3_y3;
  wire f_u_arrmul24_fa2_3_y4;
  wire f_u_arrmul24_and3_3_a_3;
  wire f_u_arrmul24_and3_3_b_3;
  wire f_u_arrmul24_and3_3_y0;
  wire f_u_arrmul24_fa3_3_f_u_arrmul24_and3_3_y0;
  wire f_u_arrmul24_fa3_3_f_u_arrmul24_fa4_2_y2;
  wire f_u_arrmul24_fa3_3_y0;
  wire f_u_arrmul24_fa3_3_y1;
  wire f_u_arrmul24_fa3_3_f_u_arrmul24_fa2_3_y4;
  wire f_u_arrmul24_fa3_3_y2;
  wire f_u_arrmul24_fa3_3_y3;
  wire f_u_arrmul24_fa3_3_y4;
  wire f_u_arrmul24_and4_3_a_4;
  wire f_u_arrmul24_and4_3_b_3;
  wire f_u_arrmul24_and4_3_y0;
  wire f_u_arrmul24_fa4_3_f_u_arrmul24_and4_3_y0;
  wire f_u_arrmul24_fa4_3_f_u_arrmul24_fa5_2_y2;
  wire f_u_arrmul24_fa4_3_y0;
  wire f_u_arrmul24_fa4_3_y1;
  wire f_u_arrmul24_fa4_3_f_u_arrmul24_fa3_3_y4;
  wire f_u_arrmul24_fa4_3_y2;
  wire f_u_arrmul24_fa4_3_y3;
  wire f_u_arrmul24_fa4_3_y4;
  wire f_u_arrmul24_and5_3_a_5;
  wire f_u_arrmul24_and5_3_b_3;
  wire f_u_arrmul24_and5_3_y0;
  wire f_u_arrmul24_fa5_3_f_u_arrmul24_and5_3_y0;
  wire f_u_arrmul24_fa5_3_f_u_arrmul24_fa6_2_y2;
  wire f_u_arrmul24_fa5_3_y0;
  wire f_u_arrmul24_fa5_3_y1;
  wire f_u_arrmul24_fa5_3_f_u_arrmul24_fa4_3_y4;
  wire f_u_arrmul24_fa5_3_y2;
  wire f_u_arrmul24_fa5_3_y3;
  wire f_u_arrmul24_fa5_3_y4;
  wire f_u_arrmul24_and6_3_a_6;
  wire f_u_arrmul24_and6_3_b_3;
  wire f_u_arrmul24_and6_3_y0;
  wire f_u_arrmul24_fa6_3_f_u_arrmul24_and6_3_y0;
  wire f_u_arrmul24_fa6_3_f_u_arrmul24_fa7_2_y2;
  wire f_u_arrmul24_fa6_3_y0;
  wire f_u_arrmul24_fa6_3_y1;
  wire f_u_arrmul24_fa6_3_f_u_arrmul24_fa5_3_y4;
  wire f_u_arrmul24_fa6_3_y2;
  wire f_u_arrmul24_fa6_3_y3;
  wire f_u_arrmul24_fa6_3_y4;
  wire f_u_arrmul24_and7_3_a_7;
  wire f_u_arrmul24_and7_3_b_3;
  wire f_u_arrmul24_and7_3_y0;
  wire f_u_arrmul24_fa7_3_f_u_arrmul24_and7_3_y0;
  wire f_u_arrmul24_fa7_3_f_u_arrmul24_fa8_2_y2;
  wire f_u_arrmul24_fa7_3_y0;
  wire f_u_arrmul24_fa7_3_y1;
  wire f_u_arrmul24_fa7_3_f_u_arrmul24_fa6_3_y4;
  wire f_u_arrmul24_fa7_3_y2;
  wire f_u_arrmul24_fa7_3_y3;
  wire f_u_arrmul24_fa7_3_y4;
  wire f_u_arrmul24_and8_3_a_8;
  wire f_u_arrmul24_and8_3_b_3;
  wire f_u_arrmul24_and8_3_y0;
  wire f_u_arrmul24_fa8_3_f_u_arrmul24_and8_3_y0;
  wire f_u_arrmul24_fa8_3_f_u_arrmul24_fa9_2_y2;
  wire f_u_arrmul24_fa8_3_y0;
  wire f_u_arrmul24_fa8_3_y1;
  wire f_u_arrmul24_fa8_3_f_u_arrmul24_fa7_3_y4;
  wire f_u_arrmul24_fa8_3_y2;
  wire f_u_arrmul24_fa8_3_y3;
  wire f_u_arrmul24_fa8_3_y4;
  wire f_u_arrmul24_and9_3_a_9;
  wire f_u_arrmul24_and9_3_b_3;
  wire f_u_arrmul24_and9_3_y0;
  wire f_u_arrmul24_fa9_3_f_u_arrmul24_and9_3_y0;
  wire f_u_arrmul24_fa9_3_f_u_arrmul24_fa10_2_y2;
  wire f_u_arrmul24_fa9_3_y0;
  wire f_u_arrmul24_fa9_3_y1;
  wire f_u_arrmul24_fa9_3_f_u_arrmul24_fa8_3_y4;
  wire f_u_arrmul24_fa9_3_y2;
  wire f_u_arrmul24_fa9_3_y3;
  wire f_u_arrmul24_fa9_3_y4;
  wire f_u_arrmul24_and10_3_a_10;
  wire f_u_arrmul24_and10_3_b_3;
  wire f_u_arrmul24_and10_3_y0;
  wire f_u_arrmul24_fa10_3_f_u_arrmul24_and10_3_y0;
  wire f_u_arrmul24_fa10_3_f_u_arrmul24_fa11_2_y2;
  wire f_u_arrmul24_fa10_3_y0;
  wire f_u_arrmul24_fa10_3_y1;
  wire f_u_arrmul24_fa10_3_f_u_arrmul24_fa9_3_y4;
  wire f_u_arrmul24_fa10_3_y2;
  wire f_u_arrmul24_fa10_3_y3;
  wire f_u_arrmul24_fa10_3_y4;
  wire f_u_arrmul24_and11_3_a_11;
  wire f_u_arrmul24_and11_3_b_3;
  wire f_u_arrmul24_and11_3_y0;
  wire f_u_arrmul24_fa11_3_f_u_arrmul24_and11_3_y0;
  wire f_u_arrmul24_fa11_3_f_u_arrmul24_fa12_2_y2;
  wire f_u_arrmul24_fa11_3_y0;
  wire f_u_arrmul24_fa11_3_y1;
  wire f_u_arrmul24_fa11_3_f_u_arrmul24_fa10_3_y4;
  wire f_u_arrmul24_fa11_3_y2;
  wire f_u_arrmul24_fa11_3_y3;
  wire f_u_arrmul24_fa11_3_y4;
  wire f_u_arrmul24_and12_3_a_12;
  wire f_u_arrmul24_and12_3_b_3;
  wire f_u_arrmul24_and12_3_y0;
  wire f_u_arrmul24_fa12_3_f_u_arrmul24_and12_3_y0;
  wire f_u_arrmul24_fa12_3_f_u_arrmul24_fa13_2_y2;
  wire f_u_arrmul24_fa12_3_y0;
  wire f_u_arrmul24_fa12_3_y1;
  wire f_u_arrmul24_fa12_3_f_u_arrmul24_fa11_3_y4;
  wire f_u_arrmul24_fa12_3_y2;
  wire f_u_arrmul24_fa12_3_y3;
  wire f_u_arrmul24_fa12_3_y4;
  wire f_u_arrmul24_and13_3_a_13;
  wire f_u_arrmul24_and13_3_b_3;
  wire f_u_arrmul24_and13_3_y0;
  wire f_u_arrmul24_fa13_3_f_u_arrmul24_and13_3_y0;
  wire f_u_arrmul24_fa13_3_f_u_arrmul24_fa14_2_y2;
  wire f_u_arrmul24_fa13_3_y0;
  wire f_u_arrmul24_fa13_3_y1;
  wire f_u_arrmul24_fa13_3_f_u_arrmul24_fa12_3_y4;
  wire f_u_arrmul24_fa13_3_y2;
  wire f_u_arrmul24_fa13_3_y3;
  wire f_u_arrmul24_fa13_3_y4;
  wire f_u_arrmul24_and14_3_a_14;
  wire f_u_arrmul24_and14_3_b_3;
  wire f_u_arrmul24_and14_3_y0;
  wire f_u_arrmul24_fa14_3_f_u_arrmul24_and14_3_y0;
  wire f_u_arrmul24_fa14_3_f_u_arrmul24_fa15_2_y2;
  wire f_u_arrmul24_fa14_3_y0;
  wire f_u_arrmul24_fa14_3_y1;
  wire f_u_arrmul24_fa14_3_f_u_arrmul24_fa13_3_y4;
  wire f_u_arrmul24_fa14_3_y2;
  wire f_u_arrmul24_fa14_3_y3;
  wire f_u_arrmul24_fa14_3_y4;
  wire f_u_arrmul24_and15_3_a_15;
  wire f_u_arrmul24_and15_3_b_3;
  wire f_u_arrmul24_and15_3_y0;
  wire f_u_arrmul24_fa15_3_f_u_arrmul24_and15_3_y0;
  wire f_u_arrmul24_fa15_3_f_u_arrmul24_fa16_2_y2;
  wire f_u_arrmul24_fa15_3_y0;
  wire f_u_arrmul24_fa15_3_y1;
  wire f_u_arrmul24_fa15_3_f_u_arrmul24_fa14_3_y4;
  wire f_u_arrmul24_fa15_3_y2;
  wire f_u_arrmul24_fa15_3_y3;
  wire f_u_arrmul24_fa15_3_y4;
  wire f_u_arrmul24_and16_3_a_16;
  wire f_u_arrmul24_and16_3_b_3;
  wire f_u_arrmul24_and16_3_y0;
  wire f_u_arrmul24_fa16_3_f_u_arrmul24_and16_3_y0;
  wire f_u_arrmul24_fa16_3_f_u_arrmul24_fa17_2_y2;
  wire f_u_arrmul24_fa16_3_y0;
  wire f_u_arrmul24_fa16_3_y1;
  wire f_u_arrmul24_fa16_3_f_u_arrmul24_fa15_3_y4;
  wire f_u_arrmul24_fa16_3_y2;
  wire f_u_arrmul24_fa16_3_y3;
  wire f_u_arrmul24_fa16_3_y4;
  wire f_u_arrmul24_and17_3_a_17;
  wire f_u_arrmul24_and17_3_b_3;
  wire f_u_arrmul24_and17_3_y0;
  wire f_u_arrmul24_fa17_3_f_u_arrmul24_and17_3_y0;
  wire f_u_arrmul24_fa17_3_f_u_arrmul24_fa18_2_y2;
  wire f_u_arrmul24_fa17_3_y0;
  wire f_u_arrmul24_fa17_3_y1;
  wire f_u_arrmul24_fa17_3_f_u_arrmul24_fa16_3_y4;
  wire f_u_arrmul24_fa17_3_y2;
  wire f_u_arrmul24_fa17_3_y3;
  wire f_u_arrmul24_fa17_3_y4;
  wire f_u_arrmul24_and18_3_a_18;
  wire f_u_arrmul24_and18_3_b_3;
  wire f_u_arrmul24_and18_3_y0;
  wire f_u_arrmul24_fa18_3_f_u_arrmul24_and18_3_y0;
  wire f_u_arrmul24_fa18_3_f_u_arrmul24_fa19_2_y2;
  wire f_u_arrmul24_fa18_3_y0;
  wire f_u_arrmul24_fa18_3_y1;
  wire f_u_arrmul24_fa18_3_f_u_arrmul24_fa17_3_y4;
  wire f_u_arrmul24_fa18_3_y2;
  wire f_u_arrmul24_fa18_3_y3;
  wire f_u_arrmul24_fa18_3_y4;
  wire f_u_arrmul24_and19_3_a_19;
  wire f_u_arrmul24_and19_3_b_3;
  wire f_u_arrmul24_and19_3_y0;
  wire f_u_arrmul24_fa19_3_f_u_arrmul24_and19_3_y0;
  wire f_u_arrmul24_fa19_3_f_u_arrmul24_fa20_2_y2;
  wire f_u_arrmul24_fa19_3_y0;
  wire f_u_arrmul24_fa19_3_y1;
  wire f_u_arrmul24_fa19_3_f_u_arrmul24_fa18_3_y4;
  wire f_u_arrmul24_fa19_3_y2;
  wire f_u_arrmul24_fa19_3_y3;
  wire f_u_arrmul24_fa19_3_y4;
  wire f_u_arrmul24_and20_3_a_20;
  wire f_u_arrmul24_and20_3_b_3;
  wire f_u_arrmul24_and20_3_y0;
  wire f_u_arrmul24_fa20_3_f_u_arrmul24_and20_3_y0;
  wire f_u_arrmul24_fa20_3_f_u_arrmul24_fa21_2_y2;
  wire f_u_arrmul24_fa20_3_y0;
  wire f_u_arrmul24_fa20_3_y1;
  wire f_u_arrmul24_fa20_3_f_u_arrmul24_fa19_3_y4;
  wire f_u_arrmul24_fa20_3_y2;
  wire f_u_arrmul24_fa20_3_y3;
  wire f_u_arrmul24_fa20_3_y4;
  wire f_u_arrmul24_and21_3_a_21;
  wire f_u_arrmul24_and21_3_b_3;
  wire f_u_arrmul24_and21_3_y0;
  wire f_u_arrmul24_fa21_3_f_u_arrmul24_and21_3_y0;
  wire f_u_arrmul24_fa21_3_f_u_arrmul24_fa22_2_y2;
  wire f_u_arrmul24_fa21_3_y0;
  wire f_u_arrmul24_fa21_3_y1;
  wire f_u_arrmul24_fa21_3_f_u_arrmul24_fa20_3_y4;
  wire f_u_arrmul24_fa21_3_y2;
  wire f_u_arrmul24_fa21_3_y3;
  wire f_u_arrmul24_fa21_3_y4;
  wire f_u_arrmul24_and22_3_a_22;
  wire f_u_arrmul24_and22_3_b_3;
  wire f_u_arrmul24_and22_3_y0;
  wire f_u_arrmul24_fa22_3_f_u_arrmul24_and22_3_y0;
  wire f_u_arrmul24_fa22_3_f_u_arrmul24_fa23_2_y2;
  wire f_u_arrmul24_fa22_3_y0;
  wire f_u_arrmul24_fa22_3_y1;
  wire f_u_arrmul24_fa22_3_f_u_arrmul24_fa21_3_y4;
  wire f_u_arrmul24_fa22_3_y2;
  wire f_u_arrmul24_fa22_3_y3;
  wire f_u_arrmul24_fa22_3_y4;
  wire f_u_arrmul24_and23_3_a_23;
  wire f_u_arrmul24_and23_3_b_3;
  wire f_u_arrmul24_and23_3_y0;
  wire f_u_arrmul24_fa23_3_f_u_arrmul24_and23_3_y0;
  wire f_u_arrmul24_fa23_3_f_u_arrmul24_fa23_2_y4;
  wire f_u_arrmul24_fa23_3_y0;
  wire f_u_arrmul24_fa23_3_y1;
  wire f_u_arrmul24_fa23_3_f_u_arrmul24_fa22_3_y4;
  wire f_u_arrmul24_fa23_3_y2;
  wire f_u_arrmul24_fa23_3_y3;
  wire f_u_arrmul24_fa23_3_y4;
  wire f_u_arrmul24_and0_4_a_0;
  wire f_u_arrmul24_and0_4_b_4;
  wire f_u_arrmul24_and0_4_y0;
  wire f_u_arrmul24_ha0_4_f_u_arrmul24_and0_4_y0;
  wire f_u_arrmul24_ha0_4_f_u_arrmul24_fa1_3_y2;
  wire f_u_arrmul24_ha0_4_y0;
  wire f_u_arrmul24_ha0_4_y1;
  wire f_u_arrmul24_and1_4_a_1;
  wire f_u_arrmul24_and1_4_b_4;
  wire f_u_arrmul24_and1_4_y0;
  wire f_u_arrmul24_fa1_4_f_u_arrmul24_and1_4_y0;
  wire f_u_arrmul24_fa1_4_f_u_arrmul24_fa2_3_y2;
  wire f_u_arrmul24_fa1_4_y0;
  wire f_u_arrmul24_fa1_4_y1;
  wire f_u_arrmul24_fa1_4_f_u_arrmul24_ha0_4_y1;
  wire f_u_arrmul24_fa1_4_y2;
  wire f_u_arrmul24_fa1_4_y3;
  wire f_u_arrmul24_fa1_4_y4;
  wire f_u_arrmul24_and2_4_a_2;
  wire f_u_arrmul24_and2_4_b_4;
  wire f_u_arrmul24_and2_4_y0;
  wire f_u_arrmul24_fa2_4_f_u_arrmul24_and2_4_y0;
  wire f_u_arrmul24_fa2_4_f_u_arrmul24_fa3_3_y2;
  wire f_u_arrmul24_fa2_4_y0;
  wire f_u_arrmul24_fa2_4_y1;
  wire f_u_arrmul24_fa2_4_f_u_arrmul24_fa1_4_y4;
  wire f_u_arrmul24_fa2_4_y2;
  wire f_u_arrmul24_fa2_4_y3;
  wire f_u_arrmul24_fa2_4_y4;
  wire f_u_arrmul24_and3_4_a_3;
  wire f_u_arrmul24_and3_4_b_4;
  wire f_u_arrmul24_and3_4_y0;
  wire f_u_arrmul24_fa3_4_f_u_arrmul24_and3_4_y0;
  wire f_u_arrmul24_fa3_4_f_u_arrmul24_fa4_3_y2;
  wire f_u_arrmul24_fa3_4_y0;
  wire f_u_arrmul24_fa3_4_y1;
  wire f_u_arrmul24_fa3_4_f_u_arrmul24_fa2_4_y4;
  wire f_u_arrmul24_fa3_4_y2;
  wire f_u_arrmul24_fa3_4_y3;
  wire f_u_arrmul24_fa3_4_y4;
  wire f_u_arrmul24_and4_4_a_4;
  wire f_u_arrmul24_and4_4_b_4;
  wire f_u_arrmul24_and4_4_y0;
  wire f_u_arrmul24_fa4_4_f_u_arrmul24_and4_4_y0;
  wire f_u_arrmul24_fa4_4_f_u_arrmul24_fa5_3_y2;
  wire f_u_arrmul24_fa4_4_y0;
  wire f_u_arrmul24_fa4_4_y1;
  wire f_u_arrmul24_fa4_4_f_u_arrmul24_fa3_4_y4;
  wire f_u_arrmul24_fa4_4_y2;
  wire f_u_arrmul24_fa4_4_y3;
  wire f_u_arrmul24_fa4_4_y4;
  wire f_u_arrmul24_and5_4_a_5;
  wire f_u_arrmul24_and5_4_b_4;
  wire f_u_arrmul24_and5_4_y0;
  wire f_u_arrmul24_fa5_4_f_u_arrmul24_and5_4_y0;
  wire f_u_arrmul24_fa5_4_f_u_arrmul24_fa6_3_y2;
  wire f_u_arrmul24_fa5_4_y0;
  wire f_u_arrmul24_fa5_4_y1;
  wire f_u_arrmul24_fa5_4_f_u_arrmul24_fa4_4_y4;
  wire f_u_arrmul24_fa5_4_y2;
  wire f_u_arrmul24_fa5_4_y3;
  wire f_u_arrmul24_fa5_4_y4;
  wire f_u_arrmul24_and6_4_a_6;
  wire f_u_arrmul24_and6_4_b_4;
  wire f_u_arrmul24_and6_4_y0;
  wire f_u_arrmul24_fa6_4_f_u_arrmul24_and6_4_y0;
  wire f_u_arrmul24_fa6_4_f_u_arrmul24_fa7_3_y2;
  wire f_u_arrmul24_fa6_4_y0;
  wire f_u_arrmul24_fa6_4_y1;
  wire f_u_arrmul24_fa6_4_f_u_arrmul24_fa5_4_y4;
  wire f_u_arrmul24_fa6_4_y2;
  wire f_u_arrmul24_fa6_4_y3;
  wire f_u_arrmul24_fa6_4_y4;
  wire f_u_arrmul24_and7_4_a_7;
  wire f_u_arrmul24_and7_4_b_4;
  wire f_u_arrmul24_and7_4_y0;
  wire f_u_arrmul24_fa7_4_f_u_arrmul24_and7_4_y0;
  wire f_u_arrmul24_fa7_4_f_u_arrmul24_fa8_3_y2;
  wire f_u_arrmul24_fa7_4_y0;
  wire f_u_arrmul24_fa7_4_y1;
  wire f_u_arrmul24_fa7_4_f_u_arrmul24_fa6_4_y4;
  wire f_u_arrmul24_fa7_4_y2;
  wire f_u_arrmul24_fa7_4_y3;
  wire f_u_arrmul24_fa7_4_y4;
  wire f_u_arrmul24_and8_4_a_8;
  wire f_u_arrmul24_and8_4_b_4;
  wire f_u_arrmul24_and8_4_y0;
  wire f_u_arrmul24_fa8_4_f_u_arrmul24_and8_4_y0;
  wire f_u_arrmul24_fa8_4_f_u_arrmul24_fa9_3_y2;
  wire f_u_arrmul24_fa8_4_y0;
  wire f_u_arrmul24_fa8_4_y1;
  wire f_u_arrmul24_fa8_4_f_u_arrmul24_fa7_4_y4;
  wire f_u_arrmul24_fa8_4_y2;
  wire f_u_arrmul24_fa8_4_y3;
  wire f_u_arrmul24_fa8_4_y4;
  wire f_u_arrmul24_and9_4_a_9;
  wire f_u_arrmul24_and9_4_b_4;
  wire f_u_arrmul24_and9_4_y0;
  wire f_u_arrmul24_fa9_4_f_u_arrmul24_and9_4_y0;
  wire f_u_arrmul24_fa9_4_f_u_arrmul24_fa10_3_y2;
  wire f_u_arrmul24_fa9_4_y0;
  wire f_u_arrmul24_fa9_4_y1;
  wire f_u_arrmul24_fa9_4_f_u_arrmul24_fa8_4_y4;
  wire f_u_arrmul24_fa9_4_y2;
  wire f_u_arrmul24_fa9_4_y3;
  wire f_u_arrmul24_fa9_4_y4;
  wire f_u_arrmul24_and10_4_a_10;
  wire f_u_arrmul24_and10_4_b_4;
  wire f_u_arrmul24_and10_4_y0;
  wire f_u_arrmul24_fa10_4_f_u_arrmul24_and10_4_y0;
  wire f_u_arrmul24_fa10_4_f_u_arrmul24_fa11_3_y2;
  wire f_u_arrmul24_fa10_4_y0;
  wire f_u_arrmul24_fa10_4_y1;
  wire f_u_arrmul24_fa10_4_f_u_arrmul24_fa9_4_y4;
  wire f_u_arrmul24_fa10_4_y2;
  wire f_u_arrmul24_fa10_4_y3;
  wire f_u_arrmul24_fa10_4_y4;
  wire f_u_arrmul24_and11_4_a_11;
  wire f_u_arrmul24_and11_4_b_4;
  wire f_u_arrmul24_and11_4_y0;
  wire f_u_arrmul24_fa11_4_f_u_arrmul24_and11_4_y0;
  wire f_u_arrmul24_fa11_4_f_u_arrmul24_fa12_3_y2;
  wire f_u_arrmul24_fa11_4_y0;
  wire f_u_arrmul24_fa11_4_y1;
  wire f_u_arrmul24_fa11_4_f_u_arrmul24_fa10_4_y4;
  wire f_u_arrmul24_fa11_4_y2;
  wire f_u_arrmul24_fa11_4_y3;
  wire f_u_arrmul24_fa11_4_y4;
  wire f_u_arrmul24_and12_4_a_12;
  wire f_u_arrmul24_and12_4_b_4;
  wire f_u_arrmul24_and12_4_y0;
  wire f_u_arrmul24_fa12_4_f_u_arrmul24_and12_4_y0;
  wire f_u_arrmul24_fa12_4_f_u_arrmul24_fa13_3_y2;
  wire f_u_arrmul24_fa12_4_y0;
  wire f_u_arrmul24_fa12_4_y1;
  wire f_u_arrmul24_fa12_4_f_u_arrmul24_fa11_4_y4;
  wire f_u_arrmul24_fa12_4_y2;
  wire f_u_arrmul24_fa12_4_y3;
  wire f_u_arrmul24_fa12_4_y4;
  wire f_u_arrmul24_and13_4_a_13;
  wire f_u_arrmul24_and13_4_b_4;
  wire f_u_arrmul24_and13_4_y0;
  wire f_u_arrmul24_fa13_4_f_u_arrmul24_and13_4_y0;
  wire f_u_arrmul24_fa13_4_f_u_arrmul24_fa14_3_y2;
  wire f_u_arrmul24_fa13_4_y0;
  wire f_u_arrmul24_fa13_4_y1;
  wire f_u_arrmul24_fa13_4_f_u_arrmul24_fa12_4_y4;
  wire f_u_arrmul24_fa13_4_y2;
  wire f_u_arrmul24_fa13_4_y3;
  wire f_u_arrmul24_fa13_4_y4;
  wire f_u_arrmul24_and14_4_a_14;
  wire f_u_arrmul24_and14_4_b_4;
  wire f_u_arrmul24_and14_4_y0;
  wire f_u_arrmul24_fa14_4_f_u_arrmul24_and14_4_y0;
  wire f_u_arrmul24_fa14_4_f_u_arrmul24_fa15_3_y2;
  wire f_u_arrmul24_fa14_4_y0;
  wire f_u_arrmul24_fa14_4_y1;
  wire f_u_arrmul24_fa14_4_f_u_arrmul24_fa13_4_y4;
  wire f_u_arrmul24_fa14_4_y2;
  wire f_u_arrmul24_fa14_4_y3;
  wire f_u_arrmul24_fa14_4_y4;
  wire f_u_arrmul24_and15_4_a_15;
  wire f_u_arrmul24_and15_4_b_4;
  wire f_u_arrmul24_and15_4_y0;
  wire f_u_arrmul24_fa15_4_f_u_arrmul24_and15_4_y0;
  wire f_u_arrmul24_fa15_4_f_u_arrmul24_fa16_3_y2;
  wire f_u_arrmul24_fa15_4_y0;
  wire f_u_arrmul24_fa15_4_y1;
  wire f_u_arrmul24_fa15_4_f_u_arrmul24_fa14_4_y4;
  wire f_u_arrmul24_fa15_4_y2;
  wire f_u_arrmul24_fa15_4_y3;
  wire f_u_arrmul24_fa15_4_y4;
  wire f_u_arrmul24_and16_4_a_16;
  wire f_u_arrmul24_and16_4_b_4;
  wire f_u_arrmul24_and16_4_y0;
  wire f_u_arrmul24_fa16_4_f_u_arrmul24_and16_4_y0;
  wire f_u_arrmul24_fa16_4_f_u_arrmul24_fa17_3_y2;
  wire f_u_arrmul24_fa16_4_y0;
  wire f_u_arrmul24_fa16_4_y1;
  wire f_u_arrmul24_fa16_4_f_u_arrmul24_fa15_4_y4;
  wire f_u_arrmul24_fa16_4_y2;
  wire f_u_arrmul24_fa16_4_y3;
  wire f_u_arrmul24_fa16_4_y4;
  wire f_u_arrmul24_and17_4_a_17;
  wire f_u_arrmul24_and17_4_b_4;
  wire f_u_arrmul24_and17_4_y0;
  wire f_u_arrmul24_fa17_4_f_u_arrmul24_and17_4_y0;
  wire f_u_arrmul24_fa17_4_f_u_arrmul24_fa18_3_y2;
  wire f_u_arrmul24_fa17_4_y0;
  wire f_u_arrmul24_fa17_4_y1;
  wire f_u_arrmul24_fa17_4_f_u_arrmul24_fa16_4_y4;
  wire f_u_arrmul24_fa17_4_y2;
  wire f_u_arrmul24_fa17_4_y3;
  wire f_u_arrmul24_fa17_4_y4;
  wire f_u_arrmul24_and18_4_a_18;
  wire f_u_arrmul24_and18_4_b_4;
  wire f_u_arrmul24_and18_4_y0;
  wire f_u_arrmul24_fa18_4_f_u_arrmul24_and18_4_y0;
  wire f_u_arrmul24_fa18_4_f_u_arrmul24_fa19_3_y2;
  wire f_u_arrmul24_fa18_4_y0;
  wire f_u_arrmul24_fa18_4_y1;
  wire f_u_arrmul24_fa18_4_f_u_arrmul24_fa17_4_y4;
  wire f_u_arrmul24_fa18_4_y2;
  wire f_u_arrmul24_fa18_4_y3;
  wire f_u_arrmul24_fa18_4_y4;
  wire f_u_arrmul24_and19_4_a_19;
  wire f_u_arrmul24_and19_4_b_4;
  wire f_u_arrmul24_and19_4_y0;
  wire f_u_arrmul24_fa19_4_f_u_arrmul24_and19_4_y0;
  wire f_u_arrmul24_fa19_4_f_u_arrmul24_fa20_3_y2;
  wire f_u_arrmul24_fa19_4_y0;
  wire f_u_arrmul24_fa19_4_y1;
  wire f_u_arrmul24_fa19_4_f_u_arrmul24_fa18_4_y4;
  wire f_u_arrmul24_fa19_4_y2;
  wire f_u_arrmul24_fa19_4_y3;
  wire f_u_arrmul24_fa19_4_y4;
  wire f_u_arrmul24_and20_4_a_20;
  wire f_u_arrmul24_and20_4_b_4;
  wire f_u_arrmul24_and20_4_y0;
  wire f_u_arrmul24_fa20_4_f_u_arrmul24_and20_4_y0;
  wire f_u_arrmul24_fa20_4_f_u_arrmul24_fa21_3_y2;
  wire f_u_arrmul24_fa20_4_y0;
  wire f_u_arrmul24_fa20_4_y1;
  wire f_u_arrmul24_fa20_4_f_u_arrmul24_fa19_4_y4;
  wire f_u_arrmul24_fa20_4_y2;
  wire f_u_arrmul24_fa20_4_y3;
  wire f_u_arrmul24_fa20_4_y4;
  wire f_u_arrmul24_and21_4_a_21;
  wire f_u_arrmul24_and21_4_b_4;
  wire f_u_arrmul24_and21_4_y0;
  wire f_u_arrmul24_fa21_4_f_u_arrmul24_and21_4_y0;
  wire f_u_arrmul24_fa21_4_f_u_arrmul24_fa22_3_y2;
  wire f_u_arrmul24_fa21_4_y0;
  wire f_u_arrmul24_fa21_4_y1;
  wire f_u_arrmul24_fa21_4_f_u_arrmul24_fa20_4_y4;
  wire f_u_arrmul24_fa21_4_y2;
  wire f_u_arrmul24_fa21_4_y3;
  wire f_u_arrmul24_fa21_4_y4;
  wire f_u_arrmul24_and22_4_a_22;
  wire f_u_arrmul24_and22_4_b_4;
  wire f_u_arrmul24_and22_4_y0;
  wire f_u_arrmul24_fa22_4_f_u_arrmul24_and22_4_y0;
  wire f_u_arrmul24_fa22_4_f_u_arrmul24_fa23_3_y2;
  wire f_u_arrmul24_fa22_4_y0;
  wire f_u_arrmul24_fa22_4_y1;
  wire f_u_arrmul24_fa22_4_f_u_arrmul24_fa21_4_y4;
  wire f_u_arrmul24_fa22_4_y2;
  wire f_u_arrmul24_fa22_4_y3;
  wire f_u_arrmul24_fa22_4_y4;
  wire f_u_arrmul24_and23_4_a_23;
  wire f_u_arrmul24_and23_4_b_4;
  wire f_u_arrmul24_and23_4_y0;
  wire f_u_arrmul24_fa23_4_f_u_arrmul24_and23_4_y0;
  wire f_u_arrmul24_fa23_4_f_u_arrmul24_fa23_3_y4;
  wire f_u_arrmul24_fa23_4_y0;
  wire f_u_arrmul24_fa23_4_y1;
  wire f_u_arrmul24_fa23_4_f_u_arrmul24_fa22_4_y4;
  wire f_u_arrmul24_fa23_4_y2;
  wire f_u_arrmul24_fa23_4_y3;
  wire f_u_arrmul24_fa23_4_y4;
  wire f_u_arrmul24_and0_5_a_0;
  wire f_u_arrmul24_and0_5_b_5;
  wire f_u_arrmul24_and0_5_y0;
  wire f_u_arrmul24_ha0_5_f_u_arrmul24_and0_5_y0;
  wire f_u_arrmul24_ha0_5_f_u_arrmul24_fa1_4_y2;
  wire f_u_arrmul24_ha0_5_y0;
  wire f_u_arrmul24_ha0_5_y1;
  wire f_u_arrmul24_and1_5_a_1;
  wire f_u_arrmul24_and1_5_b_5;
  wire f_u_arrmul24_and1_5_y0;
  wire f_u_arrmul24_fa1_5_f_u_arrmul24_and1_5_y0;
  wire f_u_arrmul24_fa1_5_f_u_arrmul24_fa2_4_y2;
  wire f_u_arrmul24_fa1_5_y0;
  wire f_u_arrmul24_fa1_5_y1;
  wire f_u_arrmul24_fa1_5_f_u_arrmul24_ha0_5_y1;
  wire f_u_arrmul24_fa1_5_y2;
  wire f_u_arrmul24_fa1_5_y3;
  wire f_u_arrmul24_fa1_5_y4;
  wire f_u_arrmul24_and2_5_a_2;
  wire f_u_arrmul24_and2_5_b_5;
  wire f_u_arrmul24_and2_5_y0;
  wire f_u_arrmul24_fa2_5_f_u_arrmul24_and2_5_y0;
  wire f_u_arrmul24_fa2_5_f_u_arrmul24_fa3_4_y2;
  wire f_u_arrmul24_fa2_5_y0;
  wire f_u_arrmul24_fa2_5_y1;
  wire f_u_arrmul24_fa2_5_f_u_arrmul24_fa1_5_y4;
  wire f_u_arrmul24_fa2_5_y2;
  wire f_u_arrmul24_fa2_5_y3;
  wire f_u_arrmul24_fa2_5_y4;
  wire f_u_arrmul24_and3_5_a_3;
  wire f_u_arrmul24_and3_5_b_5;
  wire f_u_arrmul24_and3_5_y0;
  wire f_u_arrmul24_fa3_5_f_u_arrmul24_and3_5_y0;
  wire f_u_arrmul24_fa3_5_f_u_arrmul24_fa4_4_y2;
  wire f_u_arrmul24_fa3_5_y0;
  wire f_u_arrmul24_fa3_5_y1;
  wire f_u_arrmul24_fa3_5_f_u_arrmul24_fa2_5_y4;
  wire f_u_arrmul24_fa3_5_y2;
  wire f_u_arrmul24_fa3_5_y3;
  wire f_u_arrmul24_fa3_5_y4;
  wire f_u_arrmul24_and4_5_a_4;
  wire f_u_arrmul24_and4_5_b_5;
  wire f_u_arrmul24_and4_5_y0;
  wire f_u_arrmul24_fa4_5_f_u_arrmul24_and4_5_y0;
  wire f_u_arrmul24_fa4_5_f_u_arrmul24_fa5_4_y2;
  wire f_u_arrmul24_fa4_5_y0;
  wire f_u_arrmul24_fa4_5_y1;
  wire f_u_arrmul24_fa4_5_f_u_arrmul24_fa3_5_y4;
  wire f_u_arrmul24_fa4_5_y2;
  wire f_u_arrmul24_fa4_5_y3;
  wire f_u_arrmul24_fa4_5_y4;
  wire f_u_arrmul24_and5_5_a_5;
  wire f_u_arrmul24_and5_5_b_5;
  wire f_u_arrmul24_and5_5_y0;
  wire f_u_arrmul24_fa5_5_f_u_arrmul24_and5_5_y0;
  wire f_u_arrmul24_fa5_5_f_u_arrmul24_fa6_4_y2;
  wire f_u_arrmul24_fa5_5_y0;
  wire f_u_arrmul24_fa5_5_y1;
  wire f_u_arrmul24_fa5_5_f_u_arrmul24_fa4_5_y4;
  wire f_u_arrmul24_fa5_5_y2;
  wire f_u_arrmul24_fa5_5_y3;
  wire f_u_arrmul24_fa5_5_y4;
  wire f_u_arrmul24_and6_5_a_6;
  wire f_u_arrmul24_and6_5_b_5;
  wire f_u_arrmul24_and6_5_y0;
  wire f_u_arrmul24_fa6_5_f_u_arrmul24_and6_5_y0;
  wire f_u_arrmul24_fa6_5_f_u_arrmul24_fa7_4_y2;
  wire f_u_arrmul24_fa6_5_y0;
  wire f_u_arrmul24_fa6_5_y1;
  wire f_u_arrmul24_fa6_5_f_u_arrmul24_fa5_5_y4;
  wire f_u_arrmul24_fa6_5_y2;
  wire f_u_arrmul24_fa6_5_y3;
  wire f_u_arrmul24_fa6_5_y4;
  wire f_u_arrmul24_and7_5_a_7;
  wire f_u_arrmul24_and7_5_b_5;
  wire f_u_arrmul24_and7_5_y0;
  wire f_u_arrmul24_fa7_5_f_u_arrmul24_and7_5_y0;
  wire f_u_arrmul24_fa7_5_f_u_arrmul24_fa8_4_y2;
  wire f_u_arrmul24_fa7_5_y0;
  wire f_u_arrmul24_fa7_5_y1;
  wire f_u_arrmul24_fa7_5_f_u_arrmul24_fa6_5_y4;
  wire f_u_arrmul24_fa7_5_y2;
  wire f_u_arrmul24_fa7_5_y3;
  wire f_u_arrmul24_fa7_5_y4;
  wire f_u_arrmul24_and8_5_a_8;
  wire f_u_arrmul24_and8_5_b_5;
  wire f_u_arrmul24_and8_5_y0;
  wire f_u_arrmul24_fa8_5_f_u_arrmul24_and8_5_y0;
  wire f_u_arrmul24_fa8_5_f_u_arrmul24_fa9_4_y2;
  wire f_u_arrmul24_fa8_5_y0;
  wire f_u_arrmul24_fa8_5_y1;
  wire f_u_arrmul24_fa8_5_f_u_arrmul24_fa7_5_y4;
  wire f_u_arrmul24_fa8_5_y2;
  wire f_u_arrmul24_fa8_5_y3;
  wire f_u_arrmul24_fa8_5_y4;
  wire f_u_arrmul24_and9_5_a_9;
  wire f_u_arrmul24_and9_5_b_5;
  wire f_u_arrmul24_and9_5_y0;
  wire f_u_arrmul24_fa9_5_f_u_arrmul24_and9_5_y0;
  wire f_u_arrmul24_fa9_5_f_u_arrmul24_fa10_4_y2;
  wire f_u_arrmul24_fa9_5_y0;
  wire f_u_arrmul24_fa9_5_y1;
  wire f_u_arrmul24_fa9_5_f_u_arrmul24_fa8_5_y4;
  wire f_u_arrmul24_fa9_5_y2;
  wire f_u_arrmul24_fa9_5_y3;
  wire f_u_arrmul24_fa9_5_y4;
  wire f_u_arrmul24_and10_5_a_10;
  wire f_u_arrmul24_and10_5_b_5;
  wire f_u_arrmul24_and10_5_y0;
  wire f_u_arrmul24_fa10_5_f_u_arrmul24_and10_5_y0;
  wire f_u_arrmul24_fa10_5_f_u_arrmul24_fa11_4_y2;
  wire f_u_arrmul24_fa10_5_y0;
  wire f_u_arrmul24_fa10_5_y1;
  wire f_u_arrmul24_fa10_5_f_u_arrmul24_fa9_5_y4;
  wire f_u_arrmul24_fa10_5_y2;
  wire f_u_arrmul24_fa10_5_y3;
  wire f_u_arrmul24_fa10_5_y4;
  wire f_u_arrmul24_and11_5_a_11;
  wire f_u_arrmul24_and11_5_b_5;
  wire f_u_arrmul24_and11_5_y0;
  wire f_u_arrmul24_fa11_5_f_u_arrmul24_and11_5_y0;
  wire f_u_arrmul24_fa11_5_f_u_arrmul24_fa12_4_y2;
  wire f_u_arrmul24_fa11_5_y0;
  wire f_u_arrmul24_fa11_5_y1;
  wire f_u_arrmul24_fa11_5_f_u_arrmul24_fa10_5_y4;
  wire f_u_arrmul24_fa11_5_y2;
  wire f_u_arrmul24_fa11_5_y3;
  wire f_u_arrmul24_fa11_5_y4;
  wire f_u_arrmul24_and12_5_a_12;
  wire f_u_arrmul24_and12_5_b_5;
  wire f_u_arrmul24_and12_5_y0;
  wire f_u_arrmul24_fa12_5_f_u_arrmul24_and12_5_y0;
  wire f_u_arrmul24_fa12_5_f_u_arrmul24_fa13_4_y2;
  wire f_u_arrmul24_fa12_5_y0;
  wire f_u_arrmul24_fa12_5_y1;
  wire f_u_arrmul24_fa12_5_f_u_arrmul24_fa11_5_y4;
  wire f_u_arrmul24_fa12_5_y2;
  wire f_u_arrmul24_fa12_5_y3;
  wire f_u_arrmul24_fa12_5_y4;
  wire f_u_arrmul24_and13_5_a_13;
  wire f_u_arrmul24_and13_5_b_5;
  wire f_u_arrmul24_and13_5_y0;
  wire f_u_arrmul24_fa13_5_f_u_arrmul24_and13_5_y0;
  wire f_u_arrmul24_fa13_5_f_u_arrmul24_fa14_4_y2;
  wire f_u_arrmul24_fa13_5_y0;
  wire f_u_arrmul24_fa13_5_y1;
  wire f_u_arrmul24_fa13_5_f_u_arrmul24_fa12_5_y4;
  wire f_u_arrmul24_fa13_5_y2;
  wire f_u_arrmul24_fa13_5_y3;
  wire f_u_arrmul24_fa13_5_y4;
  wire f_u_arrmul24_and14_5_a_14;
  wire f_u_arrmul24_and14_5_b_5;
  wire f_u_arrmul24_and14_5_y0;
  wire f_u_arrmul24_fa14_5_f_u_arrmul24_and14_5_y0;
  wire f_u_arrmul24_fa14_5_f_u_arrmul24_fa15_4_y2;
  wire f_u_arrmul24_fa14_5_y0;
  wire f_u_arrmul24_fa14_5_y1;
  wire f_u_arrmul24_fa14_5_f_u_arrmul24_fa13_5_y4;
  wire f_u_arrmul24_fa14_5_y2;
  wire f_u_arrmul24_fa14_5_y3;
  wire f_u_arrmul24_fa14_5_y4;
  wire f_u_arrmul24_and15_5_a_15;
  wire f_u_arrmul24_and15_5_b_5;
  wire f_u_arrmul24_and15_5_y0;
  wire f_u_arrmul24_fa15_5_f_u_arrmul24_and15_5_y0;
  wire f_u_arrmul24_fa15_5_f_u_arrmul24_fa16_4_y2;
  wire f_u_arrmul24_fa15_5_y0;
  wire f_u_arrmul24_fa15_5_y1;
  wire f_u_arrmul24_fa15_5_f_u_arrmul24_fa14_5_y4;
  wire f_u_arrmul24_fa15_5_y2;
  wire f_u_arrmul24_fa15_5_y3;
  wire f_u_arrmul24_fa15_5_y4;
  wire f_u_arrmul24_and16_5_a_16;
  wire f_u_arrmul24_and16_5_b_5;
  wire f_u_arrmul24_and16_5_y0;
  wire f_u_arrmul24_fa16_5_f_u_arrmul24_and16_5_y0;
  wire f_u_arrmul24_fa16_5_f_u_arrmul24_fa17_4_y2;
  wire f_u_arrmul24_fa16_5_y0;
  wire f_u_arrmul24_fa16_5_y1;
  wire f_u_arrmul24_fa16_5_f_u_arrmul24_fa15_5_y4;
  wire f_u_arrmul24_fa16_5_y2;
  wire f_u_arrmul24_fa16_5_y3;
  wire f_u_arrmul24_fa16_5_y4;
  wire f_u_arrmul24_and17_5_a_17;
  wire f_u_arrmul24_and17_5_b_5;
  wire f_u_arrmul24_and17_5_y0;
  wire f_u_arrmul24_fa17_5_f_u_arrmul24_and17_5_y0;
  wire f_u_arrmul24_fa17_5_f_u_arrmul24_fa18_4_y2;
  wire f_u_arrmul24_fa17_5_y0;
  wire f_u_arrmul24_fa17_5_y1;
  wire f_u_arrmul24_fa17_5_f_u_arrmul24_fa16_5_y4;
  wire f_u_arrmul24_fa17_5_y2;
  wire f_u_arrmul24_fa17_5_y3;
  wire f_u_arrmul24_fa17_5_y4;
  wire f_u_arrmul24_and18_5_a_18;
  wire f_u_arrmul24_and18_5_b_5;
  wire f_u_arrmul24_and18_5_y0;
  wire f_u_arrmul24_fa18_5_f_u_arrmul24_and18_5_y0;
  wire f_u_arrmul24_fa18_5_f_u_arrmul24_fa19_4_y2;
  wire f_u_arrmul24_fa18_5_y0;
  wire f_u_arrmul24_fa18_5_y1;
  wire f_u_arrmul24_fa18_5_f_u_arrmul24_fa17_5_y4;
  wire f_u_arrmul24_fa18_5_y2;
  wire f_u_arrmul24_fa18_5_y3;
  wire f_u_arrmul24_fa18_5_y4;
  wire f_u_arrmul24_and19_5_a_19;
  wire f_u_arrmul24_and19_5_b_5;
  wire f_u_arrmul24_and19_5_y0;
  wire f_u_arrmul24_fa19_5_f_u_arrmul24_and19_5_y0;
  wire f_u_arrmul24_fa19_5_f_u_arrmul24_fa20_4_y2;
  wire f_u_arrmul24_fa19_5_y0;
  wire f_u_arrmul24_fa19_5_y1;
  wire f_u_arrmul24_fa19_5_f_u_arrmul24_fa18_5_y4;
  wire f_u_arrmul24_fa19_5_y2;
  wire f_u_arrmul24_fa19_5_y3;
  wire f_u_arrmul24_fa19_5_y4;
  wire f_u_arrmul24_and20_5_a_20;
  wire f_u_arrmul24_and20_5_b_5;
  wire f_u_arrmul24_and20_5_y0;
  wire f_u_arrmul24_fa20_5_f_u_arrmul24_and20_5_y0;
  wire f_u_arrmul24_fa20_5_f_u_arrmul24_fa21_4_y2;
  wire f_u_arrmul24_fa20_5_y0;
  wire f_u_arrmul24_fa20_5_y1;
  wire f_u_arrmul24_fa20_5_f_u_arrmul24_fa19_5_y4;
  wire f_u_arrmul24_fa20_5_y2;
  wire f_u_arrmul24_fa20_5_y3;
  wire f_u_arrmul24_fa20_5_y4;
  wire f_u_arrmul24_and21_5_a_21;
  wire f_u_arrmul24_and21_5_b_5;
  wire f_u_arrmul24_and21_5_y0;
  wire f_u_arrmul24_fa21_5_f_u_arrmul24_and21_5_y0;
  wire f_u_arrmul24_fa21_5_f_u_arrmul24_fa22_4_y2;
  wire f_u_arrmul24_fa21_5_y0;
  wire f_u_arrmul24_fa21_5_y1;
  wire f_u_arrmul24_fa21_5_f_u_arrmul24_fa20_5_y4;
  wire f_u_arrmul24_fa21_5_y2;
  wire f_u_arrmul24_fa21_5_y3;
  wire f_u_arrmul24_fa21_5_y4;
  wire f_u_arrmul24_and22_5_a_22;
  wire f_u_arrmul24_and22_5_b_5;
  wire f_u_arrmul24_and22_5_y0;
  wire f_u_arrmul24_fa22_5_f_u_arrmul24_and22_5_y0;
  wire f_u_arrmul24_fa22_5_f_u_arrmul24_fa23_4_y2;
  wire f_u_arrmul24_fa22_5_y0;
  wire f_u_arrmul24_fa22_5_y1;
  wire f_u_arrmul24_fa22_5_f_u_arrmul24_fa21_5_y4;
  wire f_u_arrmul24_fa22_5_y2;
  wire f_u_arrmul24_fa22_5_y3;
  wire f_u_arrmul24_fa22_5_y4;
  wire f_u_arrmul24_and23_5_a_23;
  wire f_u_arrmul24_and23_5_b_5;
  wire f_u_arrmul24_and23_5_y0;
  wire f_u_arrmul24_fa23_5_f_u_arrmul24_and23_5_y0;
  wire f_u_arrmul24_fa23_5_f_u_arrmul24_fa23_4_y4;
  wire f_u_arrmul24_fa23_5_y0;
  wire f_u_arrmul24_fa23_5_y1;
  wire f_u_arrmul24_fa23_5_f_u_arrmul24_fa22_5_y4;
  wire f_u_arrmul24_fa23_5_y2;
  wire f_u_arrmul24_fa23_5_y3;
  wire f_u_arrmul24_fa23_5_y4;
  wire f_u_arrmul24_and0_6_a_0;
  wire f_u_arrmul24_and0_6_b_6;
  wire f_u_arrmul24_and0_6_y0;
  wire f_u_arrmul24_ha0_6_f_u_arrmul24_and0_6_y0;
  wire f_u_arrmul24_ha0_6_f_u_arrmul24_fa1_5_y2;
  wire f_u_arrmul24_ha0_6_y0;
  wire f_u_arrmul24_ha0_6_y1;
  wire f_u_arrmul24_and1_6_a_1;
  wire f_u_arrmul24_and1_6_b_6;
  wire f_u_arrmul24_and1_6_y0;
  wire f_u_arrmul24_fa1_6_f_u_arrmul24_and1_6_y0;
  wire f_u_arrmul24_fa1_6_f_u_arrmul24_fa2_5_y2;
  wire f_u_arrmul24_fa1_6_y0;
  wire f_u_arrmul24_fa1_6_y1;
  wire f_u_arrmul24_fa1_6_f_u_arrmul24_ha0_6_y1;
  wire f_u_arrmul24_fa1_6_y2;
  wire f_u_arrmul24_fa1_6_y3;
  wire f_u_arrmul24_fa1_6_y4;
  wire f_u_arrmul24_and2_6_a_2;
  wire f_u_arrmul24_and2_6_b_6;
  wire f_u_arrmul24_and2_6_y0;
  wire f_u_arrmul24_fa2_6_f_u_arrmul24_and2_6_y0;
  wire f_u_arrmul24_fa2_6_f_u_arrmul24_fa3_5_y2;
  wire f_u_arrmul24_fa2_6_y0;
  wire f_u_arrmul24_fa2_6_y1;
  wire f_u_arrmul24_fa2_6_f_u_arrmul24_fa1_6_y4;
  wire f_u_arrmul24_fa2_6_y2;
  wire f_u_arrmul24_fa2_6_y3;
  wire f_u_arrmul24_fa2_6_y4;
  wire f_u_arrmul24_and3_6_a_3;
  wire f_u_arrmul24_and3_6_b_6;
  wire f_u_arrmul24_and3_6_y0;
  wire f_u_arrmul24_fa3_6_f_u_arrmul24_and3_6_y0;
  wire f_u_arrmul24_fa3_6_f_u_arrmul24_fa4_5_y2;
  wire f_u_arrmul24_fa3_6_y0;
  wire f_u_arrmul24_fa3_6_y1;
  wire f_u_arrmul24_fa3_6_f_u_arrmul24_fa2_6_y4;
  wire f_u_arrmul24_fa3_6_y2;
  wire f_u_arrmul24_fa3_6_y3;
  wire f_u_arrmul24_fa3_6_y4;
  wire f_u_arrmul24_and4_6_a_4;
  wire f_u_arrmul24_and4_6_b_6;
  wire f_u_arrmul24_and4_6_y0;
  wire f_u_arrmul24_fa4_6_f_u_arrmul24_and4_6_y0;
  wire f_u_arrmul24_fa4_6_f_u_arrmul24_fa5_5_y2;
  wire f_u_arrmul24_fa4_6_y0;
  wire f_u_arrmul24_fa4_6_y1;
  wire f_u_arrmul24_fa4_6_f_u_arrmul24_fa3_6_y4;
  wire f_u_arrmul24_fa4_6_y2;
  wire f_u_arrmul24_fa4_6_y3;
  wire f_u_arrmul24_fa4_6_y4;
  wire f_u_arrmul24_and5_6_a_5;
  wire f_u_arrmul24_and5_6_b_6;
  wire f_u_arrmul24_and5_6_y0;
  wire f_u_arrmul24_fa5_6_f_u_arrmul24_and5_6_y0;
  wire f_u_arrmul24_fa5_6_f_u_arrmul24_fa6_5_y2;
  wire f_u_arrmul24_fa5_6_y0;
  wire f_u_arrmul24_fa5_6_y1;
  wire f_u_arrmul24_fa5_6_f_u_arrmul24_fa4_6_y4;
  wire f_u_arrmul24_fa5_6_y2;
  wire f_u_arrmul24_fa5_6_y3;
  wire f_u_arrmul24_fa5_6_y4;
  wire f_u_arrmul24_and6_6_a_6;
  wire f_u_arrmul24_and6_6_b_6;
  wire f_u_arrmul24_and6_6_y0;
  wire f_u_arrmul24_fa6_6_f_u_arrmul24_and6_6_y0;
  wire f_u_arrmul24_fa6_6_f_u_arrmul24_fa7_5_y2;
  wire f_u_arrmul24_fa6_6_y0;
  wire f_u_arrmul24_fa6_6_y1;
  wire f_u_arrmul24_fa6_6_f_u_arrmul24_fa5_6_y4;
  wire f_u_arrmul24_fa6_6_y2;
  wire f_u_arrmul24_fa6_6_y3;
  wire f_u_arrmul24_fa6_6_y4;
  wire f_u_arrmul24_and7_6_a_7;
  wire f_u_arrmul24_and7_6_b_6;
  wire f_u_arrmul24_and7_6_y0;
  wire f_u_arrmul24_fa7_6_f_u_arrmul24_and7_6_y0;
  wire f_u_arrmul24_fa7_6_f_u_arrmul24_fa8_5_y2;
  wire f_u_arrmul24_fa7_6_y0;
  wire f_u_arrmul24_fa7_6_y1;
  wire f_u_arrmul24_fa7_6_f_u_arrmul24_fa6_6_y4;
  wire f_u_arrmul24_fa7_6_y2;
  wire f_u_arrmul24_fa7_6_y3;
  wire f_u_arrmul24_fa7_6_y4;
  wire f_u_arrmul24_and8_6_a_8;
  wire f_u_arrmul24_and8_6_b_6;
  wire f_u_arrmul24_and8_6_y0;
  wire f_u_arrmul24_fa8_6_f_u_arrmul24_and8_6_y0;
  wire f_u_arrmul24_fa8_6_f_u_arrmul24_fa9_5_y2;
  wire f_u_arrmul24_fa8_6_y0;
  wire f_u_arrmul24_fa8_6_y1;
  wire f_u_arrmul24_fa8_6_f_u_arrmul24_fa7_6_y4;
  wire f_u_arrmul24_fa8_6_y2;
  wire f_u_arrmul24_fa8_6_y3;
  wire f_u_arrmul24_fa8_6_y4;
  wire f_u_arrmul24_and9_6_a_9;
  wire f_u_arrmul24_and9_6_b_6;
  wire f_u_arrmul24_and9_6_y0;
  wire f_u_arrmul24_fa9_6_f_u_arrmul24_and9_6_y0;
  wire f_u_arrmul24_fa9_6_f_u_arrmul24_fa10_5_y2;
  wire f_u_arrmul24_fa9_6_y0;
  wire f_u_arrmul24_fa9_6_y1;
  wire f_u_arrmul24_fa9_6_f_u_arrmul24_fa8_6_y4;
  wire f_u_arrmul24_fa9_6_y2;
  wire f_u_arrmul24_fa9_6_y3;
  wire f_u_arrmul24_fa9_6_y4;
  wire f_u_arrmul24_and10_6_a_10;
  wire f_u_arrmul24_and10_6_b_6;
  wire f_u_arrmul24_and10_6_y0;
  wire f_u_arrmul24_fa10_6_f_u_arrmul24_and10_6_y0;
  wire f_u_arrmul24_fa10_6_f_u_arrmul24_fa11_5_y2;
  wire f_u_arrmul24_fa10_6_y0;
  wire f_u_arrmul24_fa10_6_y1;
  wire f_u_arrmul24_fa10_6_f_u_arrmul24_fa9_6_y4;
  wire f_u_arrmul24_fa10_6_y2;
  wire f_u_arrmul24_fa10_6_y3;
  wire f_u_arrmul24_fa10_6_y4;
  wire f_u_arrmul24_and11_6_a_11;
  wire f_u_arrmul24_and11_6_b_6;
  wire f_u_arrmul24_and11_6_y0;
  wire f_u_arrmul24_fa11_6_f_u_arrmul24_and11_6_y0;
  wire f_u_arrmul24_fa11_6_f_u_arrmul24_fa12_5_y2;
  wire f_u_arrmul24_fa11_6_y0;
  wire f_u_arrmul24_fa11_6_y1;
  wire f_u_arrmul24_fa11_6_f_u_arrmul24_fa10_6_y4;
  wire f_u_arrmul24_fa11_6_y2;
  wire f_u_arrmul24_fa11_6_y3;
  wire f_u_arrmul24_fa11_6_y4;
  wire f_u_arrmul24_and12_6_a_12;
  wire f_u_arrmul24_and12_6_b_6;
  wire f_u_arrmul24_and12_6_y0;
  wire f_u_arrmul24_fa12_6_f_u_arrmul24_and12_6_y0;
  wire f_u_arrmul24_fa12_6_f_u_arrmul24_fa13_5_y2;
  wire f_u_arrmul24_fa12_6_y0;
  wire f_u_arrmul24_fa12_6_y1;
  wire f_u_arrmul24_fa12_6_f_u_arrmul24_fa11_6_y4;
  wire f_u_arrmul24_fa12_6_y2;
  wire f_u_arrmul24_fa12_6_y3;
  wire f_u_arrmul24_fa12_6_y4;
  wire f_u_arrmul24_and13_6_a_13;
  wire f_u_arrmul24_and13_6_b_6;
  wire f_u_arrmul24_and13_6_y0;
  wire f_u_arrmul24_fa13_6_f_u_arrmul24_and13_6_y0;
  wire f_u_arrmul24_fa13_6_f_u_arrmul24_fa14_5_y2;
  wire f_u_arrmul24_fa13_6_y0;
  wire f_u_arrmul24_fa13_6_y1;
  wire f_u_arrmul24_fa13_6_f_u_arrmul24_fa12_6_y4;
  wire f_u_arrmul24_fa13_6_y2;
  wire f_u_arrmul24_fa13_6_y3;
  wire f_u_arrmul24_fa13_6_y4;
  wire f_u_arrmul24_and14_6_a_14;
  wire f_u_arrmul24_and14_6_b_6;
  wire f_u_arrmul24_and14_6_y0;
  wire f_u_arrmul24_fa14_6_f_u_arrmul24_and14_6_y0;
  wire f_u_arrmul24_fa14_6_f_u_arrmul24_fa15_5_y2;
  wire f_u_arrmul24_fa14_6_y0;
  wire f_u_arrmul24_fa14_6_y1;
  wire f_u_arrmul24_fa14_6_f_u_arrmul24_fa13_6_y4;
  wire f_u_arrmul24_fa14_6_y2;
  wire f_u_arrmul24_fa14_6_y3;
  wire f_u_arrmul24_fa14_6_y4;
  wire f_u_arrmul24_and15_6_a_15;
  wire f_u_arrmul24_and15_6_b_6;
  wire f_u_arrmul24_and15_6_y0;
  wire f_u_arrmul24_fa15_6_f_u_arrmul24_and15_6_y0;
  wire f_u_arrmul24_fa15_6_f_u_arrmul24_fa16_5_y2;
  wire f_u_arrmul24_fa15_6_y0;
  wire f_u_arrmul24_fa15_6_y1;
  wire f_u_arrmul24_fa15_6_f_u_arrmul24_fa14_6_y4;
  wire f_u_arrmul24_fa15_6_y2;
  wire f_u_arrmul24_fa15_6_y3;
  wire f_u_arrmul24_fa15_6_y4;
  wire f_u_arrmul24_and16_6_a_16;
  wire f_u_arrmul24_and16_6_b_6;
  wire f_u_arrmul24_and16_6_y0;
  wire f_u_arrmul24_fa16_6_f_u_arrmul24_and16_6_y0;
  wire f_u_arrmul24_fa16_6_f_u_arrmul24_fa17_5_y2;
  wire f_u_arrmul24_fa16_6_y0;
  wire f_u_arrmul24_fa16_6_y1;
  wire f_u_arrmul24_fa16_6_f_u_arrmul24_fa15_6_y4;
  wire f_u_arrmul24_fa16_6_y2;
  wire f_u_arrmul24_fa16_6_y3;
  wire f_u_arrmul24_fa16_6_y4;
  wire f_u_arrmul24_and17_6_a_17;
  wire f_u_arrmul24_and17_6_b_6;
  wire f_u_arrmul24_and17_6_y0;
  wire f_u_arrmul24_fa17_6_f_u_arrmul24_and17_6_y0;
  wire f_u_arrmul24_fa17_6_f_u_arrmul24_fa18_5_y2;
  wire f_u_arrmul24_fa17_6_y0;
  wire f_u_arrmul24_fa17_6_y1;
  wire f_u_arrmul24_fa17_6_f_u_arrmul24_fa16_6_y4;
  wire f_u_arrmul24_fa17_6_y2;
  wire f_u_arrmul24_fa17_6_y3;
  wire f_u_arrmul24_fa17_6_y4;
  wire f_u_arrmul24_and18_6_a_18;
  wire f_u_arrmul24_and18_6_b_6;
  wire f_u_arrmul24_and18_6_y0;
  wire f_u_arrmul24_fa18_6_f_u_arrmul24_and18_6_y0;
  wire f_u_arrmul24_fa18_6_f_u_arrmul24_fa19_5_y2;
  wire f_u_arrmul24_fa18_6_y0;
  wire f_u_arrmul24_fa18_6_y1;
  wire f_u_arrmul24_fa18_6_f_u_arrmul24_fa17_6_y4;
  wire f_u_arrmul24_fa18_6_y2;
  wire f_u_arrmul24_fa18_6_y3;
  wire f_u_arrmul24_fa18_6_y4;
  wire f_u_arrmul24_and19_6_a_19;
  wire f_u_arrmul24_and19_6_b_6;
  wire f_u_arrmul24_and19_6_y0;
  wire f_u_arrmul24_fa19_6_f_u_arrmul24_and19_6_y0;
  wire f_u_arrmul24_fa19_6_f_u_arrmul24_fa20_5_y2;
  wire f_u_arrmul24_fa19_6_y0;
  wire f_u_arrmul24_fa19_6_y1;
  wire f_u_arrmul24_fa19_6_f_u_arrmul24_fa18_6_y4;
  wire f_u_arrmul24_fa19_6_y2;
  wire f_u_arrmul24_fa19_6_y3;
  wire f_u_arrmul24_fa19_6_y4;
  wire f_u_arrmul24_and20_6_a_20;
  wire f_u_arrmul24_and20_6_b_6;
  wire f_u_arrmul24_and20_6_y0;
  wire f_u_arrmul24_fa20_6_f_u_arrmul24_and20_6_y0;
  wire f_u_arrmul24_fa20_6_f_u_arrmul24_fa21_5_y2;
  wire f_u_arrmul24_fa20_6_y0;
  wire f_u_arrmul24_fa20_6_y1;
  wire f_u_arrmul24_fa20_6_f_u_arrmul24_fa19_6_y4;
  wire f_u_arrmul24_fa20_6_y2;
  wire f_u_arrmul24_fa20_6_y3;
  wire f_u_arrmul24_fa20_6_y4;
  wire f_u_arrmul24_and21_6_a_21;
  wire f_u_arrmul24_and21_6_b_6;
  wire f_u_arrmul24_and21_6_y0;
  wire f_u_arrmul24_fa21_6_f_u_arrmul24_and21_6_y0;
  wire f_u_arrmul24_fa21_6_f_u_arrmul24_fa22_5_y2;
  wire f_u_arrmul24_fa21_6_y0;
  wire f_u_arrmul24_fa21_6_y1;
  wire f_u_arrmul24_fa21_6_f_u_arrmul24_fa20_6_y4;
  wire f_u_arrmul24_fa21_6_y2;
  wire f_u_arrmul24_fa21_6_y3;
  wire f_u_arrmul24_fa21_6_y4;
  wire f_u_arrmul24_and22_6_a_22;
  wire f_u_arrmul24_and22_6_b_6;
  wire f_u_arrmul24_and22_6_y0;
  wire f_u_arrmul24_fa22_6_f_u_arrmul24_and22_6_y0;
  wire f_u_arrmul24_fa22_6_f_u_arrmul24_fa23_5_y2;
  wire f_u_arrmul24_fa22_6_y0;
  wire f_u_arrmul24_fa22_6_y1;
  wire f_u_arrmul24_fa22_6_f_u_arrmul24_fa21_6_y4;
  wire f_u_arrmul24_fa22_6_y2;
  wire f_u_arrmul24_fa22_6_y3;
  wire f_u_arrmul24_fa22_6_y4;
  wire f_u_arrmul24_and23_6_a_23;
  wire f_u_arrmul24_and23_6_b_6;
  wire f_u_arrmul24_and23_6_y0;
  wire f_u_arrmul24_fa23_6_f_u_arrmul24_and23_6_y0;
  wire f_u_arrmul24_fa23_6_f_u_arrmul24_fa23_5_y4;
  wire f_u_arrmul24_fa23_6_y0;
  wire f_u_arrmul24_fa23_6_y1;
  wire f_u_arrmul24_fa23_6_f_u_arrmul24_fa22_6_y4;
  wire f_u_arrmul24_fa23_6_y2;
  wire f_u_arrmul24_fa23_6_y3;
  wire f_u_arrmul24_fa23_6_y4;
  wire f_u_arrmul24_and0_7_a_0;
  wire f_u_arrmul24_and0_7_b_7;
  wire f_u_arrmul24_and0_7_y0;
  wire f_u_arrmul24_ha0_7_f_u_arrmul24_and0_7_y0;
  wire f_u_arrmul24_ha0_7_f_u_arrmul24_fa1_6_y2;
  wire f_u_arrmul24_ha0_7_y0;
  wire f_u_arrmul24_ha0_7_y1;
  wire f_u_arrmul24_and1_7_a_1;
  wire f_u_arrmul24_and1_7_b_7;
  wire f_u_arrmul24_and1_7_y0;
  wire f_u_arrmul24_fa1_7_f_u_arrmul24_and1_7_y0;
  wire f_u_arrmul24_fa1_7_f_u_arrmul24_fa2_6_y2;
  wire f_u_arrmul24_fa1_7_y0;
  wire f_u_arrmul24_fa1_7_y1;
  wire f_u_arrmul24_fa1_7_f_u_arrmul24_ha0_7_y1;
  wire f_u_arrmul24_fa1_7_y2;
  wire f_u_arrmul24_fa1_7_y3;
  wire f_u_arrmul24_fa1_7_y4;
  wire f_u_arrmul24_and2_7_a_2;
  wire f_u_arrmul24_and2_7_b_7;
  wire f_u_arrmul24_and2_7_y0;
  wire f_u_arrmul24_fa2_7_f_u_arrmul24_and2_7_y0;
  wire f_u_arrmul24_fa2_7_f_u_arrmul24_fa3_6_y2;
  wire f_u_arrmul24_fa2_7_y0;
  wire f_u_arrmul24_fa2_7_y1;
  wire f_u_arrmul24_fa2_7_f_u_arrmul24_fa1_7_y4;
  wire f_u_arrmul24_fa2_7_y2;
  wire f_u_arrmul24_fa2_7_y3;
  wire f_u_arrmul24_fa2_7_y4;
  wire f_u_arrmul24_and3_7_a_3;
  wire f_u_arrmul24_and3_7_b_7;
  wire f_u_arrmul24_and3_7_y0;
  wire f_u_arrmul24_fa3_7_f_u_arrmul24_and3_7_y0;
  wire f_u_arrmul24_fa3_7_f_u_arrmul24_fa4_6_y2;
  wire f_u_arrmul24_fa3_7_y0;
  wire f_u_arrmul24_fa3_7_y1;
  wire f_u_arrmul24_fa3_7_f_u_arrmul24_fa2_7_y4;
  wire f_u_arrmul24_fa3_7_y2;
  wire f_u_arrmul24_fa3_7_y3;
  wire f_u_arrmul24_fa3_7_y4;
  wire f_u_arrmul24_and4_7_a_4;
  wire f_u_arrmul24_and4_7_b_7;
  wire f_u_arrmul24_and4_7_y0;
  wire f_u_arrmul24_fa4_7_f_u_arrmul24_and4_7_y0;
  wire f_u_arrmul24_fa4_7_f_u_arrmul24_fa5_6_y2;
  wire f_u_arrmul24_fa4_7_y0;
  wire f_u_arrmul24_fa4_7_y1;
  wire f_u_arrmul24_fa4_7_f_u_arrmul24_fa3_7_y4;
  wire f_u_arrmul24_fa4_7_y2;
  wire f_u_arrmul24_fa4_7_y3;
  wire f_u_arrmul24_fa4_7_y4;
  wire f_u_arrmul24_and5_7_a_5;
  wire f_u_arrmul24_and5_7_b_7;
  wire f_u_arrmul24_and5_7_y0;
  wire f_u_arrmul24_fa5_7_f_u_arrmul24_and5_7_y0;
  wire f_u_arrmul24_fa5_7_f_u_arrmul24_fa6_6_y2;
  wire f_u_arrmul24_fa5_7_y0;
  wire f_u_arrmul24_fa5_7_y1;
  wire f_u_arrmul24_fa5_7_f_u_arrmul24_fa4_7_y4;
  wire f_u_arrmul24_fa5_7_y2;
  wire f_u_arrmul24_fa5_7_y3;
  wire f_u_arrmul24_fa5_7_y4;
  wire f_u_arrmul24_and6_7_a_6;
  wire f_u_arrmul24_and6_7_b_7;
  wire f_u_arrmul24_and6_7_y0;
  wire f_u_arrmul24_fa6_7_f_u_arrmul24_and6_7_y0;
  wire f_u_arrmul24_fa6_7_f_u_arrmul24_fa7_6_y2;
  wire f_u_arrmul24_fa6_7_y0;
  wire f_u_arrmul24_fa6_7_y1;
  wire f_u_arrmul24_fa6_7_f_u_arrmul24_fa5_7_y4;
  wire f_u_arrmul24_fa6_7_y2;
  wire f_u_arrmul24_fa6_7_y3;
  wire f_u_arrmul24_fa6_7_y4;
  wire f_u_arrmul24_and7_7_a_7;
  wire f_u_arrmul24_and7_7_b_7;
  wire f_u_arrmul24_and7_7_y0;
  wire f_u_arrmul24_fa7_7_f_u_arrmul24_and7_7_y0;
  wire f_u_arrmul24_fa7_7_f_u_arrmul24_fa8_6_y2;
  wire f_u_arrmul24_fa7_7_y0;
  wire f_u_arrmul24_fa7_7_y1;
  wire f_u_arrmul24_fa7_7_f_u_arrmul24_fa6_7_y4;
  wire f_u_arrmul24_fa7_7_y2;
  wire f_u_arrmul24_fa7_7_y3;
  wire f_u_arrmul24_fa7_7_y4;
  wire f_u_arrmul24_and8_7_a_8;
  wire f_u_arrmul24_and8_7_b_7;
  wire f_u_arrmul24_and8_7_y0;
  wire f_u_arrmul24_fa8_7_f_u_arrmul24_and8_7_y0;
  wire f_u_arrmul24_fa8_7_f_u_arrmul24_fa9_6_y2;
  wire f_u_arrmul24_fa8_7_y0;
  wire f_u_arrmul24_fa8_7_y1;
  wire f_u_arrmul24_fa8_7_f_u_arrmul24_fa7_7_y4;
  wire f_u_arrmul24_fa8_7_y2;
  wire f_u_arrmul24_fa8_7_y3;
  wire f_u_arrmul24_fa8_7_y4;
  wire f_u_arrmul24_and9_7_a_9;
  wire f_u_arrmul24_and9_7_b_7;
  wire f_u_arrmul24_and9_7_y0;
  wire f_u_arrmul24_fa9_7_f_u_arrmul24_and9_7_y0;
  wire f_u_arrmul24_fa9_7_f_u_arrmul24_fa10_6_y2;
  wire f_u_arrmul24_fa9_7_y0;
  wire f_u_arrmul24_fa9_7_y1;
  wire f_u_arrmul24_fa9_7_f_u_arrmul24_fa8_7_y4;
  wire f_u_arrmul24_fa9_7_y2;
  wire f_u_arrmul24_fa9_7_y3;
  wire f_u_arrmul24_fa9_7_y4;
  wire f_u_arrmul24_and10_7_a_10;
  wire f_u_arrmul24_and10_7_b_7;
  wire f_u_arrmul24_and10_7_y0;
  wire f_u_arrmul24_fa10_7_f_u_arrmul24_and10_7_y0;
  wire f_u_arrmul24_fa10_7_f_u_arrmul24_fa11_6_y2;
  wire f_u_arrmul24_fa10_7_y0;
  wire f_u_arrmul24_fa10_7_y1;
  wire f_u_arrmul24_fa10_7_f_u_arrmul24_fa9_7_y4;
  wire f_u_arrmul24_fa10_7_y2;
  wire f_u_arrmul24_fa10_7_y3;
  wire f_u_arrmul24_fa10_7_y4;
  wire f_u_arrmul24_and11_7_a_11;
  wire f_u_arrmul24_and11_7_b_7;
  wire f_u_arrmul24_and11_7_y0;
  wire f_u_arrmul24_fa11_7_f_u_arrmul24_and11_7_y0;
  wire f_u_arrmul24_fa11_7_f_u_arrmul24_fa12_6_y2;
  wire f_u_arrmul24_fa11_7_y0;
  wire f_u_arrmul24_fa11_7_y1;
  wire f_u_arrmul24_fa11_7_f_u_arrmul24_fa10_7_y4;
  wire f_u_arrmul24_fa11_7_y2;
  wire f_u_arrmul24_fa11_7_y3;
  wire f_u_arrmul24_fa11_7_y4;
  wire f_u_arrmul24_and12_7_a_12;
  wire f_u_arrmul24_and12_7_b_7;
  wire f_u_arrmul24_and12_7_y0;
  wire f_u_arrmul24_fa12_7_f_u_arrmul24_and12_7_y0;
  wire f_u_arrmul24_fa12_7_f_u_arrmul24_fa13_6_y2;
  wire f_u_arrmul24_fa12_7_y0;
  wire f_u_arrmul24_fa12_7_y1;
  wire f_u_arrmul24_fa12_7_f_u_arrmul24_fa11_7_y4;
  wire f_u_arrmul24_fa12_7_y2;
  wire f_u_arrmul24_fa12_7_y3;
  wire f_u_arrmul24_fa12_7_y4;
  wire f_u_arrmul24_and13_7_a_13;
  wire f_u_arrmul24_and13_7_b_7;
  wire f_u_arrmul24_and13_7_y0;
  wire f_u_arrmul24_fa13_7_f_u_arrmul24_and13_7_y0;
  wire f_u_arrmul24_fa13_7_f_u_arrmul24_fa14_6_y2;
  wire f_u_arrmul24_fa13_7_y0;
  wire f_u_arrmul24_fa13_7_y1;
  wire f_u_arrmul24_fa13_7_f_u_arrmul24_fa12_7_y4;
  wire f_u_arrmul24_fa13_7_y2;
  wire f_u_arrmul24_fa13_7_y3;
  wire f_u_arrmul24_fa13_7_y4;
  wire f_u_arrmul24_and14_7_a_14;
  wire f_u_arrmul24_and14_7_b_7;
  wire f_u_arrmul24_and14_7_y0;
  wire f_u_arrmul24_fa14_7_f_u_arrmul24_and14_7_y0;
  wire f_u_arrmul24_fa14_7_f_u_arrmul24_fa15_6_y2;
  wire f_u_arrmul24_fa14_7_y0;
  wire f_u_arrmul24_fa14_7_y1;
  wire f_u_arrmul24_fa14_7_f_u_arrmul24_fa13_7_y4;
  wire f_u_arrmul24_fa14_7_y2;
  wire f_u_arrmul24_fa14_7_y3;
  wire f_u_arrmul24_fa14_7_y4;
  wire f_u_arrmul24_and15_7_a_15;
  wire f_u_arrmul24_and15_7_b_7;
  wire f_u_arrmul24_and15_7_y0;
  wire f_u_arrmul24_fa15_7_f_u_arrmul24_and15_7_y0;
  wire f_u_arrmul24_fa15_7_f_u_arrmul24_fa16_6_y2;
  wire f_u_arrmul24_fa15_7_y0;
  wire f_u_arrmul24_fa15_7_y1;
  wire f_u_arrmul24_fa15_7_f_u_arrmul24_fa14_7_y4;
  wire f_u_arrmul24_fa15_7_y2;
  wire f_u_arrmul24_fa15_7_y3;
  wire f_u_arrmul24_fa15_7_y4;
  wire f_u_arrmul24_and16_7_a_16;
  wire f_u_arrmul24_and16_7_b_7;
  wire f_u_arrmul24_and16_7_y0;
  wire f_u_arrmul24_fa16_7_f_u_arrmul24_and16_7_y0;
  wire f_u_arrmul24_fa16_7_f_u_arrmul24_fa17_6_y2;
  wire f_u_arrmul24_fa16_7_y0;
  wire f_u_arrmul24_fa16_7_y1;
  wire f_u_arrmul24_fa16_7_f_u_arrmul24_fa15_7_y4;
  wire f_u_arrmul24_fa16_7_y2;
  wire f_u_arrmul24_fa16_7_y3;
  wire f_u_arrmul24_fa16_7_y4;
  wire f_u_arrmul24_and17_7_a_17;
  wire f_u_arrmul24_and17_7_b_7;
  wire f_u_arrmul24_and17_7_y0;
  wire f_u_arrmul24_fa17_7_f_u_arrmul24_and17_7_y0;
  wire f_u_arrmul24_fa17_7_f_u_arrmul24_fa18_6_y2;
  wire f_u_arrmul24_fa17_7_y0;
  wire f_u_arrmul24_fa17_7_y1;
  wire f_u_arrmul24_fa17_7_f_u_arrmul24_fa16_7_y4;
  wire f_u_arrmul24_fa17_7_y2;
  wire f_u_arrmul24_fa17_7_y3;
  wire f_u_arrmul24_fa17_7_y4;
  wire f_u_arrmul24_and18_7_a_18;
  wire f_u_arrmul24_and18_7_b_7;
  wire f_u_arrmul24_and18_7_y0;
  wire f_u_arrmul24_fa18_7_f_u_arrmul24_and18_7_y0;
  wire f_u_arrmul24_fa18_7_f_u_arrmul24_fa19_6_y2;
  wire f_u_arrmul24_fa18_7_y0;
  wire f_u_arrmul24_fa18_7_y1;
  wire f_u_arrmul24_fa18_7_f_u_arrmul24_fa17_7_y4;
  wire f_u_arrmul24_fa18_7_y2;
  wire f_u_arrmul24_fa18_7_y3;
  wire f_u_arrmul24_fa18_7_y4;
  wire f_u_arrmul24_and19_7_a_19;
  wire f_u_arrmul24_and19_7_b_7;
  wire f_u_arrmul24_and19_7_y0;
  wire f_u_arrmul24_fa19_7_f_u_arrmul24_and19_7_y0;
  wire f_u_arrmul24_fa19_7_f_u_arrmul24_fa20_6_y2;
  wire f_u_arrmul24_fa19_7_y0;
  wire f_u_arrmul24_fa19_7_y1;
  wire f_u_arrmul24_fa19_7_f_u_arrmul24_fa18_7_y4;
  wire f_u_arrmul24_fa19_7_y2;
  wire f_u_arrmul24_fa19_7_y3;
  wire f_u_arrmul24_fa19_7_y4;
  wire f_u_arrmul24_and20_7_a_20;
  wire f_u_arrmul24_and20_7_b_7;
  wire f_u_arrmul24_and20_7_y0;
  wire f_u_arrmul24_fa20_7_f_u_arrmul24_and20_7_y0;
  wire f_u_arrmul24_fa20_7_f_u_arrmul24_fa21_6_y2;
  wire f_u_arrmul24_fa20_7_y0;
  wire f_u_arrmul24_fa20_7_y1;
  wire f_u_arrmul24_fa20_7_f_u_arrmul24_fa19_7_y4;
  wire f_u_arrmul24_fa20_7_y2;
  wire f_u_arrmul24_fa20_7_y3;
  wire f_u_arrmul24_fa20_7_y4;
  wire f_u_arrmul24_and21_7_a_21;
  wire f_u_arrmul24_and21_7_b_7;
  wire f_u_arrmul24_and21_7_y0;
  wire f_u_arrmul24_fa21_7_f_u_arrmul24_and21_7_y0;
  wire f_u_arrmul24_fa21_7_f_u_arrmul24_fa22_6_y2;
  wire f_u_arrmul24_fa21_7_y0;
  wire f_u_arrmul24_fa21_7_y1;
  wire f_u_arrmul24_fa21_7_f_u_arrmul24_fa20_7_y4;
  wire f_u_arrmul24_fa21_7_y2;
  wire f_u_arrmul24_fa21_7_y3;
  wire f_u_arrmul24_fa21_7_y4;
  wire f_u_arrmul24_and22_7_a_22;
  wire f_u_arrmul24_and22_7_b_7;
  wire f_u_arrmul24_and22_7_y0;
  wire f_u_arrmul24_fa22_7_f_u_arrmul24_and22_7_y0;
  wire f_u_arrmul24_fa22_7_f_u_arrmul24_fa23_6_y2;
  wire f_u_arrmul24_fa22_7_y0;
  wire f_u_arrmul24_fa22_7_y1;
  wire f_u_arrmul24_fa22_7_f_u_arrmul24_fa21_7_y4;
  wire f_u_arrmul24_fa22_7_y2;
  wire f_u_arrmul24_fa22_7_y3;
  wire f_u_arrmul24_fa22_7_y4;
  wire f_u_arrmul24_and23_7_a_23;
  wire f_u_arrmul24_and23_7_b_7;
  wire f_u_arrmul24_and23_7_y0;
  wire f_u_arrmul24_fa23_7_f_u_arrmul24_and23_7_y0;
  wire f_u_arrmul24_fa23_7_f_u_arrmul24_fa23_6_y4;
  wire f_u_arrmul24_fa23_7_y0;
  wire f_u_arrmul24_fa23_7_y1;
  wire f_u_arrmul24_fa23_7_f_u_arrmul24_fa22_7_y4;
  wire f_u_arrmul24_fa23_7_y2;
  wire f_u_arrmul24_fa23_7_y3;
  wire f_u_arrmul24_fa23_7_y4;
  wire f_u_arrmul24_and0_8_a_0;
  wire f_u_arrmul24_and0_8_b_8;
  wire f_u_arrmul24_and0_8_y0;
  wire f_u_arrmul24_ha0_8_f_u_arrmul24_and0_8_y0;
  wire f_u_arrmul24_ha0_8_f_u_arrmul24_fa1_7_y2;
  wire f_u_arrmul24_ha0_8_y0;
  wire f_u_arrmul24_ha0_8_y1;
  wire f_u_arrmul24_and1_8_a_1;
  wire f_u_arrmul24_and1_8_b_8;
  wire f_u_arrmul24_and1_8_y0;
  wire f_u_arrmul24_fa1_8_f_u_arrmul24_and1_8_y0;
  wire f_u_arrmul24_fa1_8_f_u_arrmul24_fa2_7_y2;
  wire f_u_arrmul24_fa1_8_y0;
  wire f_u_arrmul24_fa1_8_y1;
  wire f_u_arrmul24_fa1_8_f_u_arrmul24_ha0_8_y1;
  wire f_u_arrmul24_fa1_8_y2;
  wire f_u_arrmul24_fa1_8_y3;
  wire f_u_arrmul24_fa1_8_y4;
  wire f_u_arrmul24_and2_8_a_2;
  wire f_u_arrmul24_and2_8_b_8;
  wire f_u_arrmul24_and2_8_y0;
  wire f_u_arrmul24_fa2_8_f_u_arrmul24_and2_8_y0;
  wire f_u_arrmul24_fa2_8_f_u_arrmul24_fa3_7_y2;
  wire f_u_arrmul24_fa2_8_y0;
  wire f_u_arrmul24_fa2_8_y1;
  wire f_u_arrmul24_fa2_8_f_u_arrmul24_fa1_8_y4;
  wire f_u_arrmul24_fa2_8_y2;
  wire f_u_arrmul24_fa2_8_y3;
  wire f_u_arrmul24_fa2_8_y4;
  wire f_u_arrmul24_and3_8_a_3;
  wire f_u_arrmul24_and3_8_b_8;
  wire f_u_arrmul24_and3_8_y0;
  wire f_u_arrmul24_fa3_8_f_u_arrmul24_and3_8_y0;
  wire f_u_arrmul24_fa3_8_f_u_arrmul24_fa4_7_y2;
  wire f_u_arrmul24_fa3_8_y0;
  wire f_u_arrmul24_fa3_8_y1;
  wire f_u_arrmul24_fa3_8_f_u_arrmul24_fa2_8_y4;
  wire f_u_arrmul24_fa3_8_y2;
  wire f_u_arrmul24_fa3_8_y3;
  wire f_u_arrmul24_fa3_8_y4;
  wire f_u_arrmul24_and4_8_a_4;
  wire f_u_arrmul24_and4_8_b_8;
  wire f_u_arrmul24_and4_8_y0;
  wire f_u_arrmul24_fa4_8_f_u_arrmul24_and4_8_y0;
  wire f_u_arrmul24_fa4_8_f_u_arrmul24_fa5_7_y2;
  wire f_u_arrmul24_fa4_8_y0;
  wire f_u_arrmul24_fa4_8_y1;
  wire f_u_arrmul24_fa4_8_f_u_arrmul24_fa3_8_y4;
  wire f_u_arrmul24_fa4_8_y2;
  wire f_u_arrmul24_fa4_8_y3;
  wire f_u_arrmul24_fa4_8_y4;
  wire f_u_arrmul24_and5_8_a_5;
  wire f_u_arrmul24_and5_8_b_8;
  wire f_u_arrmul24_and5_8_y0;
  wire f_u_arrmul24_fa5_8_f_u_arrmul24_and5_8_y0;
  wire f_u_arrmul24_fa5_8_f_u_arrmul24_fa6_7_y2;
  wire f_u_arrmul24_fa5_8_y0;
  wire f_u_arrmul24_fa5_8_y1;
  wire f_u_arrmul24_fa5_8_f_u_arrmul24_fa4_8_y4;
  wire f_u_arrmul24_fa5_8_y2;
  wire f_u_arrmul24_fa5_8_y3;
  wire f_u_arrmul24_fa5_8_y4;
  wire f_u_arrmul24_and6_8_a_6;
  wire f_u_arrmul24_and6_8_b_8;
  wire f_u_arrmul24_and6_8_y0;
  wire f_u_arrmul24_fa6_8_f_u_arrmul24_and6_8_y0;
  wire f_u_arrmul24_fa6_8_f_u_arrmul24_fa7_7_y2;
  wire f_u_arrmul24_fa6_8_y0;
  wire f_u_arrmul24_fa6_8_y1;
  wire f_u_arrmul24_fa6_8_f_u_arrmul24_fa5_8_y4;
  wire f_u_arrmul24_fa6_8_y2;
  wire f_u_arrmul24_fa6_8_y3;
  wire f_u_arrmul24_fa6_8_y4;
  wire f_u_arrmul24_and7_8_a_7;
  wire f_u_arrmul24_and7_8_b_8;
  wire f_u_arrmul24_and7_8_y0;
  wire f_u_arrmul24_fa7_8_f_u_arrmul24_and7_8_y0;
  wire f_u_arrmul24_fa7_8_f_u_arrmul24_fa8_7_y2;
  wire f_u_arrmul24_fa7_8_y0;
  wire f_u_arrmul24_fa7_8_y1;
  wire f_u_arrmul24_fa7_8_f_u_arrmul24_fa6_8_y4;
  wire f_u_arrmul24_fa7_8_y2;
  wire f_u_arrmul24_fa7_8_y3;
  wire f_u_arrmul24_fa7_8_y4;
  wire f_u_arrmul24_and8_8_a_8;
  wire f_u_arrmul24_and8_8_b_8;
  wire f_u_arrmul24_and8_8_y0;
  wire f_u_arrmul24_fa8_8_f_u_arrmul24_and8_8_y0;
  wire f_u_arrmul24_fa8_8_f_u_arrmul24_fa9_7_y2;
  wire f_u_arrmul24_fa8_8_y0;
  wire f_u_arrmul24_fa8_8_y1;
  wire f_u_arrmul24_fa8_8_f_u_arrmul24_fa7_8_y4;
  wire f_u_arrmul24_fa8_8_y2;
  wire f_u_arrmul24_fa8_8_y3;
  wire f_u_arrmul24_fa8_8_y4;
  wire f_u_arrmul24_and9_8_a_9;
  wire f_u_arrmul24_and9_8_b_8;
  wire f_u_arrmul24_and9_8_y0;
  wire f_u_arrmul24_fa9_8_f_u_arrmul24_and9_8_y0;
  wire f_u_arrmul24_fa9_8_f_u_arrmul24_fa10_7_y2;
  wire f_u_arrmul24_fa9_8_y0;
  wire f_u_arrmul24_fa9_8_y1;
  wire f_u_arrmul24_fa9_8_f_u_arrmul24_fa8_8_y4;
  wire f_u_arrmul24_fa9_8_y2;
  wire f_u_arrmul24_fa9_8_y3;
  wire f_u_arrmul24_fa9_8_y4;
  wire f_u_arrmul24_and10_8_a_10;
  wire f_u_arrmul24_and10_8_b_8;
  wire f_u_arrmul24_and10_8_y0;
  wire f_u_arrmul24_fa10_8_f_u_arrmul24_and10_8_y0;
  wire f_u_arrmul24_fa10_8_f_u_arrmul24_fa11_7_y2;
  wire f_u_arrmul24_fa10_8_y0;
  wire f_u_arrmul24_fa10_8_y1;
  wire f_u_arrmul24_fa10_8_f_u_arrmul24_fa9_8_y4;
  wire f_u_arrmul24_fa10_8_y2;
  wire f_u_arrmul24_fa10_8_y3;
  wire f_u_arrmul24_fa10_8_y4;
  wire f_u_arrmul24_and11_8_a_11;
  wire f_u_arrmul24_and11_8_b_8;
  wire f_u_arrmul24_and11_8_y0;
  wire f_u_arrmul24_fa11_8_f_u_arrmul24_and11_8_y0;
  wire f_u_arrmul24_fa11_8_f_u_arrmul24_fa12_7_y2;
  wire f_u_arrmul24_fa11_8_y0;
  wire f_u_arrmul24_fa11_8_y1;
  wire f_u_arrmul24_fa11_8_f_u_arrmul24_fa10_8_y4;
  wire f_u_arrmul24_fa11_8_y2;
  wire f_u_arrmul24_fa11_8_y3;
  wire f_u_arrmul24_fa11_8_y4;
  wire f_u_arrmul24_and12_8_a_12;
  wire f_u_arrmul24_and12_8_b_8;
  wire f_u_arrmul24_and12_8_y0;
  wire f_u_arrmul24_fa12_8_f_u_arrmul24_and12_8_y0;
  wire f_u_arrmul24_fa12_8_f_u_arrmul24_fa13_7_y2;
  wire f_u_arrmul24_fa12_8_y0;
  wire f_u_arrmul24_fa12_8_y1;
  wire f_u_arrmul24_fa12_8_f_u_arrmul24_fa11_8_y4;
  wire f_u_arrmul24_fa12_8_y2;
  wire f_u_arrmul24_fa12_8_y3;
  wire f_u_arrmul24_fa12_8_y4;
  wire f_u_arrmul24_and13_8_a_13;
  wire f_u_arrmul24_and13_8_b_8;
  wire f_u_arrmul24_and13_8_y0;
  wire f_u_arrmul24_fa13_8_f_u_arrmul24_and13_8_y0;
  wire f_u_arrmul24_fa13_8_f_u_arrmul24_fa14_7_y2;
  wire f_u_arrmul24_fa13_8_y0;
  wire f_u_arrmul24_fa13_8_y1;
  wire f_u_arrmul24_fa13_8_f_u_arrmul24_fa12_8_y4;
  wire f_u_arrmul24_fa13_8_y2;
  wire f_u_arrmul24_fa13_8_y3;
  wire f_u_arrmul24_fa13_8_y4;
  wire f_u_arrmul24_and14_8_a_14;
  wire f_u_arrmul24_and14_8_b_8;
  wire f_u_arrmul24_and14_8_y0;
  wire f_u_arrmul24_fa14_8_f_u_arrmul24_and14_8_y0;
  wire f_u_arrmul24_fa14_8_f_u_arrmul24_fa15_7_y2;
  wire f_u_arrmul24_fa14_8_y0;
  wire f_u_arrmul24_fa14_8_y1;
  wire f_u_arrmul24_fa14_8_f_u_arrmul24_fa13_8_y4;
  wire f_u_arrmul24_fa14_8_y2;
  wire f_u_arrmul24_fa14_8_y3;
  wire f_u_arrmul24_fa14_8_y4;
  wire f_u_arrmul24_and15_8_a_15;
  wire f_u_arrmul24_and15_8_b_8;
  wire f_u_arrmul24_and15_8_y0;
  wire f_u_arrmul24_fa15_8_f_u_arrmul24_and15_8_y0;
  wire f_u_arrmul24_fa15_8_f_u_arrmul24_fa16_7_y2;
  wire f_u_arrmul24_fa15_8_y0;
  wire f_u_arrmul24_fa15_8_y1;
  wire f_u_arrmul24_fa15_8_f_u_arrmul24_fa14_8_y4;
  wire f_u_arrmul24_fa15_8_y2;
  wire f_u_arrmul24_fa15_8_y3;
  wire f_u_arrmul24_fa15_8_y4;
  wire f_u_arrmul24_and16_8_a_16;
  wire f_u_arrmul24_and16_8_b_8;
  wire f_u_arrmul24_and16_8_y0;
  wire f_u_arrmul24_fa16_8_f_u_arrmul24_and16_8_y0;
  wire f_u_arrmul24_fa16_8_f_u_arrmul24_fa17_7_y2;
  wire f_u_arrmul24_fa16_8_y0;
  wire f_u_arrmul24_fa16_8_y1;
  wire f_u_arrmul24_fa16_8_f_u_arrmul24_fa15_8_y4;
  wire f_u_arrmul24_fa16_8_y2;
  wire f_u_arrmul24_fa16_8_y3;
  wire f_u_arrmul24_fa16_8_y4;
  wire f_u_arrmul24_and17_8_a_17;
  wire f_u_arrmul24_and17_8_b_8;
  wire f_u_arrmul24_and17_8_y0;
  wire f_u_arrmul24_fa17_8_f_u_arrmul24_and17_8_y0;
  wire f_u_arrmul24_fa17_8_f_u_arrmul24_fa18_7_y2;
  wire f_u_arrmul24_fa17_8_y0;
  wire f_u_arrmul24_fa17_8_y1;
  wire f_u_arrmul24_fa17_8_f_u_arrmul24_fa16_8_y4;
  wire f_u_arrmul24_fa17_8_y2;
  wire f_u_arrmul24_fa17_8_y3;
  wire f_u_arrmul24_fa17_8_y4;
  wire f_u_arrmul24_and18_8_a_18;
  wire f_u_arrmul24_and18_8_b_8;
  wire f_u_arrmul24_and18_8_y0;
  wire f_u_arrmul24_fa18_8_f_u_arrmul24_and18_8_y0;
  wire f_u_arrmul24_fa18_8_f_u_arrmul24_fa19_7_y2;
  wire f_u_arrmul24_fa18_8_y0;
  wire f_u_arrmul24_fa18_8_y1;
  wire f_u_arrmul24_fa18_8_f_u_arrmul24_fa17_8_y4;
  wire f_u_arrmul24_fa18_8_y2;
  wire f_u_arrmul24_fa18_8_y3;
  wire f_u_arrmul24_fa18_8_y4;
  wire f_u_arrmul24_and19_8_a_19;
  wire f_u_arrmul24_and19_8_b_8;
  wire f_u_arrmul24_and19_8_y0;
  wire f_u_arrmul24_fa19_8_f_u_arrmul24_and19_8_y0;
  wire f_u_arrmul24_fa19_8_f_u_arrmul24_fa20_7_y2;
  wire f_u_arrmul24_fa19_8_y0;
  wire f_u_arrmul24_fa19_8_y1;
  wire f_u_arrmul24_fa19_8_f_u_arrmul24_fa18_8_y4;
  wire f_u_arrmul24_fa19_8_y2;
  wire f_u_arrmul24_fa19_8_y3;
  wire f_u_arrmul24_fa19_8_y4;
  wire f_u_arrmul24_and20_8_a_20;
  wire f_u_arrmul24_and20_8_b_8;
  wire f_u_arrmul24_and20_8_y0;
  wire f_u_arrmul24_fa20_8_f_u_arrmul24_and20_8_y0;
  wire f_u_arrmul24_fa20_8_f_u_arrmul24_fa21_7_y2;
  wire f_u_arrmul24_fa20_8_y0;
  wire f_u_arrmul24_fa20_8_y1;
  wire f_u_arrmul24_fa20_8_f_u_arrmul24_fa19_8_y4;
  wire f_u_arrmul24_fa20_8_y2;
  wire f_u_arrmul24_fa20_8_y3;
  wire f_u_arrmul24_fa20_8_y4;
  wire f_u_arrmul24_and21_8_a_21;
  wire f_u_arrmul24_and21_8_b_8;
  wire f_u_arrmul24_and21_8_y0;
  wire f_u_arrmul24_fa21_8_f_u_arrmul24_and21_8_y0;
  wire f_u_arrmul24_fa21_8_f_u_arrmul24_fa22_7_y2;
  wire f_u_arrmul24_fa21_8_y0;
  wire f_u_arrmul24_fa21_8_y1;
  wire f_u_arrmul24_fa21_8_f_u_arrmul24_fa20_8_y4;
  wire f_u_arrmul24_fa21_8_y2;
  wire f_u_arrmul24_fa21_8_y3;
  wire f_u_arrmul24_fa21_8_y4;
  wire f_u_arrmul24_and22_8_a_22;
  wire f_u_arrmul24_and22_8_b_8;
  wire f_u_arrmul24_and22_8_y0;
  wire f_u_arrmul24_fa22_8_f_u_arrmul24_and22_8_y0;
  wire f_u_arrmul24_fa22_8_f_u_arrmul24_fa23_7_y2;
  wire f_u_arrmul24_fa22_8_y0;
  wire f_u_arrmul24_fa22_8_y1;
  wire f_u_arrmul24_fa22_8_f_u_arrmul24_fa21_8_y4;
  wire f_u_arrmul24_fa22_8_y2;
  wire f_u_arrmul24_fa22_8_y3;
  wire f_u_arrmul24_fa22_8_y4;
  wire f_u_arrmul24_and23_8_a_23;
  wire f_u_arrmul24_and23_8_b_8;
  wire f_u_arrmul24_and23_8_y0;
  wire f_u_arrmul24_fa23_8_f_u_arrmul24_and23_8_y0;
  wire f_u_arrmul24_fa23_8_f_u_arrmul24_fa23_7_y4;
  wire f_u_arrmul24_fa23_8_y0;
  wire f_u_arrmul24_fa23_8_y1;
  wire f_u_arrmul24_fa23_8_f_u_arrmul24_fa22_8_y4;
  wire f_u_arrmul24_fa23_8_y2;
  wire f_u_arrmul24_fa23_8_y3;
  wire f_u_arrmul24_fa23_8_y4;
  wire f_u_arrmul24_and0_9_a_0;
  wire f_u_arrmul24_and0_9_b_9;
  wire f_u_arrmul24_and0_9_y0;
  wire f_u_arrmul24_ha0_9_f_u_arrmul24_and0_9_y0;
  wire f_u_arrmul24_ha0_9_f_u_arrmul24_fa1_8_y2;
  wire f_u_arrmul24_ha0_9_y0;
  wire f_u_arrmul24_ha0_9_y1;
  wire f_u_arrmul24_and1_9_a_1;
  wire f_u_arrmul24_and1_9_b_9;
  wire f_u_arrmul24_and1_9_y0;
  wire f_u_arrmul24_fa1_9_f_u_arrmul24_and1_9_y0;
  wire f_u_arrmul24_fa1_9_f_u_arrmul24_fa2_8_y2;
  wire f_u_arrmul24_fa1_9_y0;
  wire f_u_arrmul24_fa1_9_y1;
  wire f_u_arrmul24_fa1_9_f_u_arrmul24_ha0_9_y1;
  wire f_u_arrmul24_fa1_9_y2;
  wire f_u_arrmul24_fa1_9_y3;
  wire f_u_arrmul24_fa1_9_y4;
  wire f_u_arrmul24_and2_9_a_2;
  wire f_u_arrmul24_and2_9_b_9;
  wire f_u_arrmul24_and2_9_y0;
  wire f_u_arrmul24_fa2_9_f_u_arrmul24_and2_9_y0;
  wire f_u_arrmul24_fa2_9_f_u_arrmul24_fa3_8_y2;
  wire f_u_arrmul24_fa2_9_y0;
  wire f_u_arrmul24_fa2_9_y1;
  wire f_u_arrmul24_fa2_9_f_u_arrmul24_fa1_9_y4;
  wire f_u_arrmul24_fa2_9_y2;
  wire f_u_arrmul24_fa2_9_y3;
  wire f_u_arrmul24_fa2_9_y4;
  wire f_u_arrmul24_and3_9_a_3;
  wire f_u_arrmul24_and3_9_b_9;
  wire f_u_arrmul24_and3_9_y0;
  wire f_u_arrmul24_fa3_9_f_u_arrmul24_and3_9_y0;
  wire f_u_arrmul24_fa3_9_f_u_arrmul24_fa4_8_y2;
  wire f_u_arrmul24_fa3_9_y0;
  wire f_u_arrmul24_fa3_9_y1;
  wire f_u_arrmul24_fa3_9_f_u_arrmul24_fa2_9_y4;
  wire f_u_arrmul24_fa3_9_y2;
  wire f_u_arrmul24_fa3_9_y3;
  wire f_u_arrmul24_fa3_9_y4;
  wire f_u_arrmul24_and4_9_a_4;
  wire f_u_arrmul24_and4_9_b_9;
  wire f_u_arrmul24_and4_9_y0;
  wire f_u_arrmul24_fa4_9_f_u_arrmul24_and4_9_y0;
  wire f_u_arrmul24_fa4_9_f_u_arrmul24_fa5_8_y2;
  wire f_u_arrmul24_fa4_9_y0;
  wire f_u_arrmul24_fa4_9_y1;
  wire f_u_arrmul24_fa4_9_f_u_arrmul24_fa3_9_y4;
  wire f_u_arrmul24_fa4_9_y2;
  wire f_u_arrmul24_fa4_9_y3;
  wire f_u_arrmul24_fa4_9_y4;
  wire f_u_arrmul24_and5_9_a_5;
  wire f_u_arrmul24_and5_9_b_9;
  wire f_u_arrmul24_and5_9_y0;
  wire f_u_arrmul24_fa5_9_f_u_arrmul24_and5_9_y0;
  wire f_u_arrmul24_fa5_9_f_u_arrmul24_fa6_8_y2;
  wire f_u_arrmul24_fa5_9_y0;
  wire f_u_arrmul24_fa5_9_y1;
  wire f_u_arrmul24_fa5_9_f_u_arrmul24_fa4_9_y4;
  wire f_u_arrmul24_fa5_9_y2;
  wire f_u_arrmul24_fa5_9_y3;
  wire f_u_arrmul24_fa5_9_y4;
  wire f_u_arrmul24_and6_9_a_6;
  wire f_u_arrmul24_and6_9_b_9;
  wire f_u_arrmul24_and6_9_y0;
  wire f_u_arrmul24_fa6_9_f_u_arrmul24_and6_9_y0;
  wire f_u_arrmul24_fa6_9_f_u_arrmul24_fa7_8_y2;
  wire f_u_arrmul24_fa6_9_y0;
  wire f_u_arrmul24_fa6_9_y1;
  wire f_u_arrmul24_fa6_9_f_u_arrmul24_fa5_9_y4;
  wire f_u_arrmul24_fa6_9_y2;
  wire f_u_arrmul24_fa6_9_y3;
  wire f_u_arrmul24_fa6_9_y4;
  wire f_u_arrmul24_and7_9_a_7;
  wire f_u_arrmul24_and7_9_b_9;
  wire f_u_arrmul24_and7_9_y0;
  wire f_u_arrmul24_fa7_9_f_u_arrmul24_and7_9_y0;
  wire f_u_arrmul24_fa7_9_f_u_arrmul24_fa8_8_y2;
  wire f_u_arrmul24_fa7_9_y0;
  wire f_u_arrmul24_fa7_9_y1;
  wire f_u_arrmul24_fa7_9_f_u_arrmul24_fa6_9_y4;
  wire f_u_arrmul24_fa7_9_y2;
  wire f_u_arrmul24_fa7_9_y3;
  wire f_u_arrmul24_fa7_9_y4;
  wire f_u_arrmul24_and8_9_a_8;
  wire f_u_arrmul24_and8_9_b_9;
  wire f_u_arrmul24_and8_9_y0;
  wire f_u_arrmul24_fa8_9_f_u_arrmul24_and8_9_y0;
  wire f_u_arrmul24_fa8_9_f_u_arrmul24_fa9_8_y2;
  wire f_u_arrmul24_fa8_9_y0;
  wire f_u_arrmul24_fa8_9_y1;
  wire f_u_arrmul24_fa8_9_f_u_arrmul24_fa7_9_y4;
  wire f_u_arrmul24_fa8_9_y2;
  wire f_u_arrmul24_fa8_9_y3;
  wire f_u_arrmul24_fa8_9_y4;
  wire f_u_arrmul24_and9_9_a_9;
  wire f_u_arrmul24_and9_9_b_9;
  wire f_u_arrmul24_and9_9_y0;
  wire f_u_arrmul24_fa9_9_f_u_arrmul24_and9_9_y0;
  wire f_u_arrmul24_fa9_9_f_u_arrmul24_fa10_8_y2;
  wire f_u_arrmul24_fa9_9_y0;
  wire f_u_arrmul24_fa9_9_y1;
  wire f_u_arrmul24_fa9_9_f_u_arrmul24_fa8_9_y4;
  wire f_u_arrmul24_fa9_9_y2;
  wire f_u_arrmul24_fa9_9_y3;
  wire f_u_arrmul24_fa9_9_y4;
  wire f_u_arrmul24_and10_9_a_10;
  wire f_u_arrmul24_and10_9_b_9;
  wire f_u_arrmul24_and10_9_y0;
  wire f_u_arrmul24_fa10_9_f_u_arrmul24_and10_9_y0;
  wire f_u_arrmul24_fa10_9_f_u_arrmul24_fa11_8_y2;
  wire f_u_arrmul24_fa10_9_y0;
  wire f_u_arrmul24_fa10_9_y1;
  wire f_u_arrmul24_fa10_9_f_u_arrmul24_fa9_9_y4;
  wire f_u_arrmul24_fa10_9_y2;
  wire f_u_arrmul24_fa10_9_y3;
  wire f_u_arrmul24_fa10_9_y4;
  wire f_u_arrmul24_and11_9_a_11;
  wire f_u_arrmul24_and11_9_b_9;
  wire f_u_arrmul24_and11_9_y0;
  wire f_u_arrmul24_fa11_9_f_u_arrmul24_and11_9_y0;
  wire f_u_arrmul24_fa11_9_f_u_arrmul24_fa12_8_y2;
  wire f_u_arrmul24_fa11_9_y0;
  wire f_u_arrmul24_fa11_9_y1;
  wire f_u_arrmul24_fa11_9_f_u_arrmul24_fa10_9_y4;
  wire f_u_arrmul24_fa11_9_y2;
  wire f_u_arrmul24_fa11_9_y3;
  wire f_u_arrmul24_fa11_9_y4;
  wire f_u_arrmul24_and12_9_a_12;
  wire f_u_arrmul24_and12_9_b_9;
  wire f_u_arrmul24_and12_9_y0;
  wire f_u_arrmul24_fa12_9_f_u_arrmul24_and12_9_y0;
  wire f_u_arrmul24_fa12_9_f_u_arrmul24_fa13_8_y2;
  wire f_u_arrmul24_fa12_9_y0;
  wire f_u_arrmul24_fa12_9_y1;
  wire f_u_arrmul24_fa12_9_f_u_arrmul24_fa11_9_y4;
  wire f_u_arrmul24_fa12_9_y2;
  wire f_u_arrmul24_fa12_9_y3;
  wire f_u_arrmul24_fa12_9_y4;
  wire f_u_arrmul24_and13_9_a_13;
  wire f_u_arrmul24_and13_9_b_9;
  wire f_u_arrmul24_and13_9_y0;
  wire f_u_arrmul24_fa13_9_f_u_arrmul24_and13_9_y0;
  wire f_u_arrmul24_fa13_9_f_u_arrmul24_fa14_8_y2;
  wire f_u_arrmul24_fa13_9_y0;
  wire f_u_arrmul24_fa13_9_y1;
  wire f_u_arrmul24_fa13_9_f_u_arrmul24_fa12_9_y4;
  wire f_u_arrmul24_fa13_9_y2;
  wire f_u_arrmul24_fa13_9_y3;
  wire f_u_arrmul24_fa13_9_y4;
  wire f_u_arrmul24_and14_9_a_14;
  wire f_u_arrmul24_and14_9_b_9;
  wire f_u_arrmul24_and14_9_y0;
  wire f_u_arrmul24_fa14_9_f_u_arrmul24_and14_9_y0;
  wire f_u_arrmul24_fa14_9_f_u_arrmul24_fa15_8_y2;
  wire f_u_arrmul24_fa14_9_y0;
  wire f_u_arrmul24_fa14_9_y1;
  wire f_u_arrmul24_fa14_9_f_u_arrmul24_fa13_9_y4;
  wire f_u_arrmul24_fa14_9_y2;
  wire f_u_arrmul24_fa14_9_y3;
  wire f_u_arrmul24_fa14_9_y4;
  wire f_u_arrmul24_and15_9_a_15;
  wire f_u_arrmul24_and15_9_b_9;
  wire f_u_arrmul24_and15_9_y0;
  wire f_u_arrmul24_fa15_9_f_u_arrmul24_and15_9_y0;
  wire f_u_arrmul24_fa15_9_f_u_arrmul24_fa16_8_y2;
  wire f_u_arrmul24_fa15_9_y0;
  wire f_u_arrmul24_fa15_9_y1;
  wire f_u_arrmul24_fa15_9_f_u_arrmul24_fa14_9_y4;
  wire f_u_arrmul24_fa15_9_y2;
  wire f_u_arrmul24_fa15_9_y3;
  wire f_u_arrmul24_fa15_9_y4;
  wire f_u_arrmul24_and16_9_a_16;
  wire f_u_arrmul24_and16_9_b_9;
  wire f_u_arrmul24_and16_9_y0;
  wire f_u_arrmul24_fa16_9_f_u_arrmul24_and16_9_y0;
  wire f_u_arrmul24_fa16_9_f_u_arrmul24_fa17_8_y2;
  wire f_u_arrmul24_fa16_9_y0;
  wire f_u_arrmul24_fa16_9_y1;
  wire f_u_arrmul24_fa16_9_f_u_arrmul24_fa15_9_y4;
  wire f_u_arrmul24_fa16_9_y2;
  wire f_u_arrmul24_fa16_9_y3;
  wire f_u_arrmul24_fa16_9_y4;
  wire f_u_arrmul24_and17_9_a_17;
  wire f_u_arrmul24_and17_9_b_9;
  wire f_u_arrmul24_and17_9_y0;
  wire f_u_arrmul24_fa17_9_f_u_arrmul24_and17_9_y0;
  wire f_u_arrmul24_fa17_9_f_u_arrmul24_fa18_8_y2;
  wire f_u_arrmul24_fa17_9_y0;
  wire f_u_arrmul24_fa17_9_y1;
  wire f_u_arrmul24_fa17_9_f_u_arrmul24_fa16_9_y4;
  wire f_u_arrmul24_fa17_9_y2;
  wire f_u_arrmul24_fa17_9_y3;
  wire f_u_arrmul24_fa17_9_y4;
  wire f_u_arrmul24_and18_9_a_18;
  wire f_u_arrmul24_and18_9_b_9;
  wire f_u_arrmul24_and18_9_y0;
  wire f_u_arrmul24_fa18_9_f_u_arrmul24_and18_9_y0;
  wire f_u_arrmul24_fa18_9_f_u_arrmul24_fa19_8_y2;
  wire f_u_arrmul24_fa18_9_y0;
  wire f_u_arrmul24_fa18_9_y1;
  wire f_u_arrmul24_fa18_9_f_u_arrmul24_fa17_9_y4;
  wire f_u_arrmul24_fa18_9_y2;
  wire f_u_arrmul24_fa18_9_y3;
  wire f_u_arrmul24_fa18_9_y4;
  wire f_u_arrmul24_and19_9_a_19;
  wire f_u_arrmul24_and19_9_b_9;
  wire f_u_arrmul24_and19_9_y0;
  wire f_u_arrmul24_fa19_9_f_u_arrmul24_and19_9_y0;
  wire f_u_arrmul24_fa19_9_f_u_arrmul24_fa20_8_y2;
  wire f_u_arrmul24_fa19_9_y0;
  wire f_u_arrmul24_fa19_9_y1;
  wire f_u_arrmul24_fa19_9_f_u_arrmul24_fa18_9_y4;
  wire f_u_arrmul24_fa19_9_y2;
  wire f_u_arrmul24_fa19_9_y3;
  wire f_u_arrmul24_fa19_9_y4;
  wire f_u_arrmul24_and20_9_a_20;
  wire f_u_arrmul24_and20_9_b_9;
  wire f_u_arrmul24_and20_9_y0;
  wire f_u_arrmul24_fa20_9_f_u_arrmul24_and20_9_y0;
  wire f_u_arrmul24_fa20_9_f_u_arrmul24_fa21_8_y2;
  wire f_u_arrmul24_fa20_9_y0;
  wire f_u_arrmul24_fa20_9_y1;
  wire f_u_arrmul24_fa20_9_f_u_arrmul24_fa19_9_y4;
  wire f_u_arrmul24_fa20_9_y2;
  wire f_u_arrmul24_fa20_9_y3;
  wire f_u_arrmul24_fa20_9_y4;
  wire f_u_arrmul24_and21_9_a_21;
  wire f_u_arrmul24_and21_9_b_9;
  wire f_u_arrmul24_and21_9_y0;
  wire f_u_arrmul24_fa21_9_f_u_arrmul24_and21_9_y0;
  wire f_u_arrmul24_fa21_9_f_u_arrmul24_fa22_8_y2;
  wire f_u_arrmul24_fa21_9_y0;
  wire f_u_arrmul24_fa21_9_y1;
  wire f_u_arrmul24_fa21_9_f_u_arrmul24_fa20_9_y4;
  wire f_u_arrmul24_fa21_9_y2;
  wire f_u_arrmul24_fa21_9_y3;
  wire f_u_arrmul24_fa21_9_y4;
  wire f_u_arrmul24_and22_9_a_22;
  wire f_u_arrmul24_and22_9_b_9;
  wire f_u_arrmul24_and22_9_y0;
  wire f_u_arrmul24_fa22_9_f_u_arrmul24_and22_9_y0;
  wire f_u_arrmul24_fa22_9_f_u_arrmul24_fa23_8_y2;
  wire f_u_arrmul24_fa22_9_y0;
  wire f_u_arrmul24_fa22_9_y1;
  wire f_u_arrmul24_fa22_9_f_u_arrmul24_fa21_9_y4;
  wire f_u_arrmul24_fa22_9_y2;
  wire f_u_arrmul24_fa22_9_y3;
  wire f_u_arrmul24_fa22_9_y4;
  wire f_u_arrmul24_and23_9_a_23;
  wire f_u_arrmul24_and23_9_b_9;
  wire f_u_arrmul24_and23_9_y0;
  wire f_u_arrmul24_fa23_9_f_u_arrmul24_and23_9_y0;
  wire f_u_arrmul24_fa23_9_f_u_arrmul24_fa23_8_y4;
  wire f_u_arrmul24_fa23_9_y0;
  wire f_u_arrmul24_fa23_9_y1;
  wire f_u_arrmul24_fa23_9_f_u_arrmul24_fa22_9_y4;
  wire f_u_arrmul24_fa23_9_y2;
  wire f_u_arrmul24_fa23_9_y3;
  wire f_u_arrmul24_fa23_9_y4;
  wire f_u_arrmul24_and0_10_a_0;
  wire f_u_arrmul24_and0_10_b_10;
  wire f_u_arrmul24_and0_10_y0;
  wire f_u_arrmul24_ha0_10_f_u_arrmul24_and0_10_y0;
  wire f_u_arrmul24_ha0_10_f_u_arrmul24_fa1_9_y2;
  wire f_u_arrmul24_ha0_10_y0;
  wire f_u_arrmul24_ha0_10_y1;
  wire f_u_arrmul24_and1_10_a_1;
  wire f_u_arrmul24_and1_10_b_10;
  wire f_u_arrmul24_and1_10_y0;
  wire f_u_arrmul24_fa1_10_f_u_arrmul24_and1_10_y0;
  wire f_u_arrmul24_fa1_10_f_u_arrmul24_fa2_9_y2;
  wire f_u_arrmul24_fa1_10_y0;
  wire f_u_arrmul24_fa1_10_y1;
  wire f_u_arrmul24_fa1_10_f_u_arrmul24_ha0_10_y1;
  wire f_u_arrmul24_fa1_10_y2;
  wire f_u_arrmul24_fa1_10_y3;
  wire f_u_arrmul24_fa1_10_y4;
  wire f_u_arrmul24_and2_10_a_2;
  wire f_u_arrmul24_and2_10_b_10;
  wire f_u_arrmul24_and2_10_y0;
  wire f_u_arrmul24_fa2_10_f_u_arrmul24_and2_10_y0;
  wire f_u_arrmul24_fa2_10_f_u_arrmul24_fa3_9_y2;
  wire f_u_arrmul24_fa2_10_y0;
  wire f_u_arrmul24_fa2_10_y1;
  wire f_u_arrmul24_fa2_10_f_u_arrmul24_fa1_10_y4;
  wire f_u_arrmul24_fa2_10_y2;
  wire f_u_arrmul24_fa2_10_y3;
  wire f_u_arrmul24_fa2_10_y4;
  wire f_u_arrmul24_and3_10_a_3;
  wire f_u_arrmul24_and3_10_b_10;
  wire f_u_arrmul24_and3_10_y0;
  wire f_u_arrmul24_fa3_10_f_u_arrmul24_and3_10_y0;
  wire f_u_arrmul24_fa3_10_f_u_arrmul24_fa4_9_y2;
  wire f_u_arrmul24_fa3_10_y0;
  wire f_u_arrmul24_fa3_10_y1;
  wire f_u_arrmul24_fa3_10_f_u_arrmul24_fa2_10_y4;
  wire f_u_arrmul24_fa3_10_y2;
  wire f_u_arrmul24_fa3_10_y3;
  wire f_u_arrmul24_fa3_10_y4;
  wire f_u_arrmul24_and4_10_a_4;
  wire f_u_arrmul24_and4_10_b_10;
  wire f_u_arrmul24_and4_10_y0;
  wire f_u_arrmul24_fa4_10_f_u_arrmul24_and4_10_y0;
  wire f_u_arrmul24_fa4_10_f_u_arrmul24_fa5_9_y2;
  wire f_u_arrmul24_fa4_10_y0;
  wire f_u_arrmul24_fa4_10_y1;
  wire f_u_arrmul24_fa4_10_f_u_arrmul24_fa3_10_y4;
  wire f_u_arrmul24_fa4_10_y2;
  wire f_u_arrmul24_fa4_10_y3;
  wire f_u_arrmul24_fa4_10_y4;
  wire f_u_arrmul24_and5_10_a_5;
  wire f_u_arrmul24_and5_10_b_10;
  wire f_u_arrmul24_and5_10_y0;
  wire f_u_arrmul24_fa5_10_f_u_arrmul24_and5_10_y0;
  wire f_u_arrmul24_fa5_10_f_u_arrmul24_fa6_9_y2;
  wire f_u_arrmul24_fa5_10_y0;
  wire f_u_arrmul24_fa5_10_y1;
  wire f_u_arrmul24_fa5_10_f_u_arrmul24_fa4_10_y4;
  wire f_u_arrmul24_fa5_10_y2;
  wire f_u_arrmul24_fa5_10_y3;
  wire f_u_arrmul24_fa5_10_y4;
  wire f_u_arrmul24_and6_10_a_6;
  wire f_u_arrmul24_and6_10_b_10;
  wire f_u_arrmul24_and6_10_y0;
  wire f_u_arrmul24_fa6_10_f_u_arrmul24_and6_10_y0;
  wire f_u_arrmul24_fa6_10_f_u_arrmul24_fa7_9_y2;
  wire f_u_arrmul24_fa6_10_y0;
  wire f_u_arrmul24_fa6_10_y1;
  wire f_u_arrmul24_fa6_10_f_u_arrmul24_fa5_10_y4;
  wire f_u_arrmul24_fa6_10_y2;
  wire f_u_arrmul24_fa6_10_y3;
  wire f_u_arrmul24_fa6_10_y4;
  wire f_u_arrmul24_and7_10_a_7;
  wire f_u_arrmul24_and7_10_b_10;
  wire f_u_arrmul24_and7_10_y0;
  wire f_u_arrmul24_fa7_10_f_u_arrmul24_and7_10_y0;
  wire f_u_arrmul24_fa7_10_f_u_arrmul24_fa8_9_y2;
  wire f_u_arrmul24_fa7_10_y0;
  wire f_u_arrmul24_fa7_10_y1;
  wire f_u_arrmul24_fa7_10_f_u_arrmul24_fa6_10_y4;
  wire f_u_arrmul24_fa7_10_y2;
  wire f_u_arrmul24_fa7_10_y3;
  wire f_u_arrmul24_fa7_10_y4;
  wire f_u_arrmul24_and8_10_a_8;
  wire f_u_arrmul24_and8_10_b_10;
  wire f_u_arrmul24_and8_10_y0;
  wire f_u_arrmul24_fa8_10_f_u_arrmul24_and8_10_y0;
  wire f_u_arrmul24_fa8_10_f_u_arrmul24_fa9_9_y2;
  wire f_u_arrmul24_fa8_10_y0;
  wire f_u_arrmul24_fa8_10_y1;
  wire f_u_arrmul24_fa8_10_f_u_arrmul24_fa7_10_y4;
  wire f_u_arrmul24_fa8_10_y2;
  wire f_u_arrmul24_fa8_10_y3;
  wire f_u_arrmul24_fa8_10_y4;
  wire f_u_arrmul24_and9_10_a_9;
  wire f_u_arrmul24_and9_10_b_10;
  wire f_u_arrmul24_and9_10_y0;
  wire f_u_arrmul24_fa9_10_f_u_arrmul24_and9_10_y0;
  wire f_u_arrmul24_fa9_10_f_u_arrmul24_fa10_9_y2;
  wire f_u_arrmul24_fa9_10_y0;
  wire f_u_arrmul24_fa9_10_y1;
  wire f_u_arrmul24_fa9_10_f_u_arrmul24_fa8_10_y4;
  wire f_u_arrmul24_fa9_10_y2;
  wire f_u_arrmul24_fa9_10_y3;
  wire f_u_arrmul24_fa9_10_y4;
  wire f_u_arrmul24_and10_10_a_10;
  wire f_u_arrmul24_and10_10_b_10;
  wire f_u_arrmul24_and10_10_y0;
  wire f_u_arrmul24_fa10_10_f_u_arrmul24_and10_10_y0;
  wire f_u_arrmul24_fa10_10_f_u_arrmul24_fa11_9_y2;
  wire f_u_arrmul24_fa10_10_y0;
  wire f_u_arrmul24_fa10_10_y1;
  wire f_u_arrmul24_fa10_10_f_u_arrmul24_fa9_10_y4;
  wire f_u_arrmul24_fa10_10_y2;
  wire f_u_arrmul24_fa10_10_y3;
  wire f_u_arrmul24_fa10_10_y4;
  wire f_u_arrmul24_and11_10_a_11;
  wire f_u_arrmul24_and11_10_b_10;
  wire f_u_arrmul24_and11_10_y0;
  wire f_u_arrmul24_fa11_10_f_u_arrmul24_and11_10_y0;
  wire f_u_arrmul24_fa11_10_f_u_arrmul24_fa12_9_y2;
  wire f_u_arrmul24_fa11_10_y0;
  wire f_u_arrmul24_fa11_10_y1;
  wire f_u_arrmul24_fa11_10_f_u_arrmul24_fa10_10_y4;
  wire f_u_arrmul24_fa11_10_y2;
  wire f_u_arrmul24_fa11_10_y3;
  wire f_u_arrmul24_fa11_10_y4;
  wire f_u_arrmul24_and12_10_a_12;
  wire f_u_arrmul24_and12_10_b_10;
  wire f_u_arrmul24_and12_10_y0;
  wire f_u_arrmul24_fa12_10_f_u_arrmul24_and12_10_y0;
  wire f_u_arrmul24_fa12_10_f_u_arrmul24_fa13_9_y2;
  wire f_u_arrmul24_fa12_10_y0;
  wire f_u_arrmul24_fa12_10_y1;
  wire f_u_arrmul24_fa12_10_f_u_arrmul24_fa11_10_y4;
  wire f_u_arrmul24_fa12_10_y2;
  wire f_u_arrmul24_fa12_10_y3;
  wire f_u_arrmul24_fa12_10_y4;
  wire f_u_arrmul24_and13_10_a_13;
  wire f_u_arrmul24_and13_10_b_10;
  wire f_u_arrmul24_and13_10_y0;
  wire f_u_arrmul24_fa13_10_f_u_arrmul24_and13_10_y0;
  wire f_u_arrmul24_fa13_10_f_u_arrmul24_fa14_9_y2;
  wire f_u_arrmul24_fa13_10_y0;
  wire f_u_arrmul24_fa13_10_y1;
  wire f_u_arrmul24_fa13_10_f_u_arrmul24_fa12_10_y4;
  wire f_u_arrmul24_fa13_10_y2;
  wire f_u_arrmul24_fa13_10_y3;
  wire f_u_arrmul24_fa13_10_y4;
  wire f_u_arrmul24_and14_10_a_14;
  wire f_u_arrmul24_and14_10_b_10;
  wire f_u_arrmul24_and14_10_y0;
  wire f_u_arrmul24_fa14_10_f_u_arrmul24_and14_10_y0;
  wire f_u_arrmul24_fa14_10_f_u_arrmul24_fa15_9_y2;
  wire f_u_arrmul24_fa14_10_y0;
  wire f_u_arrmul24_fa14_10_y1;
  wire f_u_arrmul24_fa14_10_f_u_arrmul24_fa13_10_y4;
  wire f_u_arrmul24_fa14_10_y2;
  wire f_u_arrmul24_fa14_10_y3;
  wire f_u_arrmul24_fa14_10_y4;
  wire f_u_arrmul24_and15_10_a_15;
  wire f_u_arrmul24_and15_10_b_10;
  wire f_u_arrmul24_and15_10_y0;
  wire f_u_arrmul24_fa15_10_f_u_arrmul24_and15_10_y0;
  wire f_u_arrmul24_fa15_10_f_u_arrmul24_fa16_9_y2;
  wire f_u_arrmul24_fa15_10_y0;
  wire f_u_arrmul24_fa15_10_y1;
  wire f_u_arrmul24_fa15_10_f_u_arrmul24_fa14_10_y4;
  wire f_u_arrmul24_fa15_10_y2;
  wire f_u_arrmul24_fa15_10_y3;
  wire f_u_arrmul24_fa15_10_y4;
  wire f_u_arrmul24_and16_10_a_16;
  wire f_u_arrmul24_and16_10_b_10;
  wire f_u_arrmul24_and16_10_y0;
  wire f_u_arrmul24_fa16_10_f_u_arrmul24_and16_10_y0;
  wire f_u_arrmul24_fa16_10_f_u_arrmul24_fa17_9_y2;
  wire f_u_arrmul24_fa16_10_y0;
  wire f_u_arrmul24_fa16_10_y1;
  wire f_u_arrmul24_fa16_10_f_u_arrmul24_fa15_10_y4;
  wire f_u_arrmul24_fa16_10_y2;
  wire f_u_arrmul24_fa16_10_y3;
  wire f_u_arrmul24_fa16_10_y4;
  wire f_u_arrmul24_and17_10_a_17;
  wire f_u_arrmul24_and17_10_b_10;
  wire f_u_arrmul24_and17_10_y0;
  wire f_u_arrmul24_fa17_10_f_u_arrmul24_and17_10_y0;
  wire f_u_arrmul24_fa17_10_f_u_arrmul24_fa18_9_y2;
  wire f_u_arrmul24_fa17_10_y0;
  wire f_u_arrmul24_fa17_10_y1;
  wire f_u_arrmul24_fa17_10_f_u_arrmul24_fa16_10_y4;
  wire f_u_arrmul24_fa17_10_y2;
  wire f_u_arrmul24_fa17_10_y3;
  wire f_u_arrmul24_fa17_10_y4;
  wire f_u_arrmul24_and18_10_a_18;
  wire f_u_arrmul24_and18_10_b_10;
  wire f_u_arrmul24_and18_10_y0;
  wire f_u_arrmul24_fa18_10_f_u_arrmul24_and18_10_y0;
  wire f_u_arrmul24_fa18_10_f_u_arrmul24_fa19_9_y2;
  wire f_u_arrmul24_fa18_10_y0;
  wire f_u_arrmul24_fa18_10_y1;
  wire f_u_arrmul24_fa18_10_f_u_arrmul24_fa17_10_y4;
  wire f_u_arrmul24_fa18_10_y2;
  wire f_u_arrmul24_fa18_10_y3;
  wire f_u_arrmul24_fa18_10_y4;
  wire f_u_arrmul24_and19_10_a_19;
  wire f_u_arrmul24_and19_10_b_10;
  wire f_u_arrmul24_and19_10_y0;
  wire f_u_arrmul24_fa19_10_f_u_arrmul24_and19_10_y0;
  wire f_u_arrmul24_fa19_10_f_u_arrmul24_fa20_9_y2;
  wire f_u_arrmul24_fa19_10_y0;
  wire f_u_arrmul24_fa19_10_y1;
  wire f_u_arrmul24_fa19_10_f_u_arrmul24_fa18_10_y4;
  wire f_u_arrmul24_fa19_10_y2;
  wire f_u_arrmul24_fa19_10_y3;
  wire f_u_arrmul24_fa19_10_y4;
  wire f_u_arrmul24_and20_10_a_20;
  wire f_u_arrmul24_and20_10_b_10;
  wire f_u_arrmul24_and20_10_y0;
  wire f_u_arrmul24_fa20_10_f_u_arrmul24_and20_10_y0;
  wire f_u_arrmul24_fa20_10_f_u_arrmul24_fa21_9_y2;
  wire f_u_arrmul24_fa20_10_y0;
  wire f_u_arrmul24_fa20_10_y1;
  wire f_u_arrmul24_fa20_10_f_u_arrmul24_fa19_10_y4;
  wire f_u_arrmul24_fa20_10_y2;
  wire f_u_arrmul24_fa20_10_y3;
  wire f_u_arrmul24_fa20_10_y4;
  wire f_u_arrmul24_and21_10_a_21;
  wire f_u_arrmul24_and21_10_b_10;
  wire f_u_arrmul24_and21_10_y0;
  wire f_u_arrmul24_fa21_10_f_u_arrmul24_and21_10_y0;
  wire f_u_arrmul24_fa21_10_f_u_arrmul24_fa22_9_y2;
  wire f_u_arrmul24_fa21_10_y0;
  wire f_u_arrmul24_fa21_10_y1;
  wire f_u_arrmul24_fa21_10_f_u_arrmul24_fa20_10_y4;
  wire f_u_arrmul24_fa21_10_y2;
  wire f_u_arrmul24_fa21_10_y3;
  wire f_u_arrmul24_fa21_10_y4;
  wire f_u_arrmul24_and22_10_a_22;
  wire f_u_arrmul24_and22_10_b_10;
  wire f_u_arrmul24_and22_10_y0;
  wire f_u_arrmul24_fa22_10_f_u_arrmul24_and22_10_y0;
  wire f_u_arrmul24_fa22_10_f_u_arrmul24_fa23_9_y2;
  wire f_u_arrmul24_fa22_10_y0;
  wire f_u_arrmul24_fa22_10_y1;
  wire f_u_arrmul24_fa22_10_f_u_arrmul24_fa21_10_y4;
  wire f_u_arrmul24_fa22_10_y2;
  wire f_u_arrmul24_fa22_10_y3;
  wire f_u_arrmul24_fa22_10_y4;
  wire f_u_arrmul24_and23_10_a_23;
  wire f_u_arrmul24_and23_10_b_10;
  wire f_u_arrmul24_and23_10_y0;
  wire f_u_arrmul24_fa23_10_f_u_arrmul24_and23_10_y0;
  wire f_u_arrmul24_fa23_10_f_u_arrmul24_fa23_9_y4;
  wire f_u_arrmul24_fa23_10_y0;
  wire f_u_arrmul24_fa23_10_y1;
  wire f_u_arrmul24_fa23_10_f_u_arrmul24_fa22_10_y4;
  wire f_u_arrmul24_fa23_10_y2;
  wire f_u_arrmul24_fa23_10_y3;
  wire f_u_arrmul24_fa23_10_y4;
  wire f_u_arrmul24_and0_11_a_0;
  wire f_u_arrmul24_and0_11_b_11;
  wire f_u_arrmul24_and0_11_y0;
  wire f_u_arrmul24_ha0_11_f_u_arrmul24_and0_11_y0;
  wire f_u_arrmul24_ha0_11_f_u_arrmul24_fa1_10_y2;
  wire f_u_arrmul24_ha0_11_y0;
  wire f_u_arrmul24_ha0_11_y1;
  wire f_u_arrmul24_and1_11_a_1;
  wire f_u_arrmul24_and1_11_b_11;
  wire f_u_arrmul24_and1_11_y0;
  wire f_u_arrmul24_fa1_11_f_u_arrmul24_and1_11_y0;
  wire f_u_arrmul24_fa1_11_f_u_arrmul24_fa2_10_y2;
  wire f_u_arrmul24_fa1_11_y0;
  wire f_u_arrmul24_fa1_11_y1;
  wire f_u_arrmul24_fa1_11_f_u_arrmul24_ha0_11_y1;
  wire f_u_arrmul24_fa1_11_y2;
  wire f_u_arrmul24_fa1_11_y3;
  wire f_u_arrmul24_fa1_11_y4;
  wire f_u_arrmul24_and2_11_a_2;
  wire f_u_arrmul24_and2_11_b_11;
  wire f_u_arrmul24_and2_11_y0;
  wire f_u_arrmul24_fa2_11_f_u_arrmul24_and2_11_y0;
  wire f_u_arrmul24_fa2_11_f_u_arrmul24_fa3_10_y2;
  wire f_u_arrmul24_fa2_11_y0;
  wire f_u_arrmul24_fa2_11_y1;
  wire f_u_arrmul24_fa2_11_f_u_arrmul24_fa1_11_y4;
  wire f_u_arrmul24_fa2_11_y2;
  wire f_u_arrmul24_fa2_11_y3;
  wire f_u_arrmul24_fa2_11_y4;
  wire f_u_arrmul24_and3_11_a_3;
  wire f_u_arrmul24_and3_11_b_11;
  wire f_u_arrmul24_and3_11_y0;
  wire f_u_arrmul24_fa3_11_f_u_arrmul24_and3_11_y0;
  wire f_u_arrmul24_fa3_11_f_u_arrmul24_fa4_10_y2;
  wire f_u_arrmul24_fa3_11_y0;
  wire f_u_arrmul24_fa3_11_y1;
  wire f_u_arrmul24_fa3_11_f_u_arrmul24_fa2_11_y4;
  wire f_u_arrmul24_fa3_11_y2;
  wire f_u_arrmul24_fa3_11_y3;
  wire f_u_arrmul24_fa3_11_y4;
  wire f_u_arrmul24_and4_11_a_4;
  wire f_u_arrmul24_and4_11_b_11;
  wire f_u_arrmul24_and4_11_y0;
  wire f_u_arrmul24_fa4_11_f_u_arrmul24_and4_11_y0;
  wire f_u_arrmul24_fa4_11_f_u_arrmul24_fa5_10_y2;
  wire f_u_arrmul24_fa4_11_y0;
  wire f_u_arrmul24_fa4_11_y1;
  wire f_u_arrmul24_fa4_11_f_u_arrmul24_fa3_11_y4;
  wire f_u_arrmul24_fa4_11_y2;
  wire f_u_arrmul24_fa4_11_y3;
  wire f_u_arrmul24_fa4_11_y4;
  wire f_u_arrmul24_and5_11_a_5;
  wire f_u_arrmul24_and5_11_b_11;
  wire f_u_arrmul24_and5_11_y0;
  wire f_u_arrmul24_fa5_11_f_u_arrmul24_and5_11_y0;
  wire f_u_arrmul24_fa5_11_f_u_arrmul24_fa6_10_y2;
  wire f_u_arrmul24_fa5_11_y0;
  wire f_u_arrmul24_fa5_11_y1;
  wire f_u_arrmul24_fa5_11_f_u_arrmul24_fa4_11_y4;
  wire f_u_arrmul24_fa5_11_y2;
  wire f_u_arrmul24_fa5_11_y3;
  wire f_u_arrmul24_fa5_11_y4;
  wire f_u_arrmul24_and6_11_a_6;
  wire f_u_arrmul24_and6_11_b_11;
  wire f_u_arrmul24_and6_11_y0;
  wire f_u_arrmul24_fa6_11_f_u_arrmul24_and6_11_y0;
  wire f_u_arrmul24_fa6_11_f_u_arrmul24_fa7_10_y2;
  wire f_u_arrmul24_fa6_11_y0;
  wire f_u_arrmul24_fa6_11_y1;
  wire f_u_arrmul24_fa6_11_f_u_arrmul24_fa5_11_y4;
  wire f_u_arrmul24_fa6_11_y2;
  wire f_u_arrmul24_fa6_11_y3;
  wire f_u_arrmul24_fa6_11_y4;
  wire f_u_arrmul24_and7_11_a_7;
  wire f_u_arrmul24_and7_11_b_11;
  wire f_u_arrmul24_and7_11_y0;
  wire f_u_arrmul24_fa7_11_f_u_arrmul24_and7_11_y0;
  wire f_u_arrmul24_fa7_11_f_u_arrmul24_fa8_10_y2;
  wire f_u_arrmul24_fa7_11_y0;
  wire f_u_arrmul24_fa7_11_y1;
  wire f_u_arrmul24_fa7_11_f_u_arrmul24_fa6_11_y4;
  wire f_u_arrmul24_fa7_11_y2;
  wire f_u_arrmul24_fa7_11_y3;
  wire f_u_arrmul24_fa7_11_y4;
  wire f_u_arrmul24_and8_11_a_8;
  wire f_u_arrmul24_and8_11_b_11;
  wire f_u_arrmul24_and8_11_y0;
  wire f_u_arrmul24_fa8_11_f_u_arrmul24_and8_11_y0;
  wire f_u_arrmul24_fa8_11_f_u_arrmul24_fa9_10_y2;
  wire f_u_arrmul24_fa8_11_y0;
  wire f_u_arrmul24_fa8_11_y1;
  wire f_u_arrmul24_fa8_11_f_u_arrmul24_fa7_11_y4;
  wire f_u_arrmul24_fa8_11_y2;
  wire f_u_arrmul24_fa8_11_y3;
  wire f_u_arrmul24_fa8_11_y4;
  wire f_u_arrmul24_and9_11_a_9;
  wire f_u_arrmul24_and9_11_b_11;
  wire f_u_arrmul24_and9_11_y0;
  wire f_u_arrmul24_fa9_11_f_u_arrmul24_and9_11_y0;
  wire f_u_arrmul24_fa9_11_f_u_arrmul24_fa10_10_y2;
  wire f_u_arrmul24_fa9_11_y0;
  wire f_u_arrmul24_fa9_11_y1;
  wire f_u_arrmul24_fa9_11_f_u_arrmul24_fa8_11_y4;
  wire f_u_arrmul24_fa9_11_y2;
  wire f_u_arrmul24_fa9_11_y3;
  wire f_u_arrmul24_fa9_11_y4;
  wire f_u_arrmul24_and10_11_a_10;
  wire f_u_arrmul24_and10_11_b_11;
  wire f_u_arrmul24_and10_11_y0;
  wire f_u_arrmul24_fa10_11_f_u_arrmul24_and10_11_y0;
  wire f_u_arrmul24_fa10_11_f_u_arrmul24_fa11_10_y2;
  wire f_u_arrmul24_fa10_11_y0;
  wire f_u_arrmul24_fa10_11_y1;
  wire f_u_arrmul24_fa10_11_f_u_arrmul24_fa9_11_y4;
  wire f_u_arrmul24_fa10_11_y2;
  wire f_u_arrmul24_fa10_11_y3;
  wire f_u_arrmul24_fa10_11_y4;
  wire f_u_arrmul24_and11_11_a_11;
  wire f_u_arrmul24_and11_11_b_11;
  wire f_u_arrmul24_and11_11_y0;
  wire f_u_arrmul24_fa11_11_f_u_arrmul24_and11_11_y0;
  wire f_u_arrmul24_fa11_11_f_u_arrmul24_fa12_10_y2;
  wire f_u_arrmul24_fa11_11_y0;
  wire f_u_arrmul24_fa11_11_y1;
  wire f_u_arrmul24_fa11_11_f_u_arrmul24_fa10_11_y4;
  wire f_u_arrmul24_fa11_11_y2;
  wire f_u_arrmul24_fa11_11_y3;
  wire f_u_arrmul24_fa11_11_y4;
  wire f_u_arrmul24_and12_11_a_12;
  wire f_u_arrmul24_and12_11_b_11;
  wire f_u_arrmul24_and12_11_y0;
  wire f_u_arrmul24_fa12_11_f_u_arrmul24_and12_11_y0;
  wire f_u_arrmul24_fa12_11_f_u_arrmul24_fa13_10_y2;
  wire f_u_arrmul24_fa12_11_y0;
  wire f_u_arrmul24_fa12_11_y1;
  wire f_u_arrmul24_fa12_11_f_u_arrmul24_fa11_11_y4;
  wire f_u_arrmul24_fa12_11_y2;
  wire f_u_arrmul24_fa12_11_y3;
  wire f_u_arrmul24_fa12_11_y4;
  wire f_u_arrmul24_and13_11_a_13;
  wire f_u_arrmul24_and13_11_b_11;
  wire f_u_arrmul24_and13_11_y0;
  wire f_u_arrmul24_fa13_11_f_u_arrmul24_and13_11_y0;
  wire f_u_arrmul24_fa13_11_f_u_arrmul24_fa14_10_y2;
  wire f_u_arrmul24_fa13_11_y0;
  wire f_u_arrmul24_fa13_11_y1;
  wire f_u_arrmul24_fa13_11_f_u_arrmul24_fa12_11_y4;
  wire f_u_arrmul24_fa13_11_y2;
  wire f_u_arrmul24_fa13_11_y3;
  wire f_u_arrmul24_fa13_11_y4;
  wire f_u_arrmul24_and14_11_a_14;
  wire f_u_arrmul24_and14_11_b_11;
  wire f_u_arrmul24_and14_11_y0;
  wire f_u_arrmul24_fa14_11_f_u_arrmul24_and14_11_y0;
  wire f_u_arrmul24_fa14_11_f_u_arrmul24_fa15_10_y2;
  wire f_u_arrmul24_fa14_11_y0;
  wire f_u_arrmul24_fa14_11_y1;
  wire f_u_arrmul24_fa14_11_f_u_arrmul24_fa13_11_y4;
  wire f_u_arrmul24_fa14_11_y2;
  wire f_u_arrmul24_fa14_11_y3;
  wire f_u_arrmul24_fa14_11_y4;
  wire f_u_arrmul24_and15_11_a_15;
  wire f_u_arrmul24_and15_11_b_11;
  wire f_u_arrmul24_and15_11_y0;
  wire f_u_arrmul24_fa15_11_f_u_arrmul24_and15_11_y0;
  wire f_u_arrmul24_fa15_11_f_u_arrmul24_fa16_10_y2;
  wire f_u_arrmul24_fa15_11_y0;
  wire f_u_arrmul24_fa15_11_y1;
  wire f_u_arrmul24_fa15_11_f_u_arrmul24_fa14_11_y4;
  wire f_u_arrmul24_fa15_11_y2;
  wire f_u_arrmul24_fa15_11_y3;
  wire f_u_arrmul24_fa15_11_y4;
  wire f_u_arrmul24_and16_11_a_16;
  wire f_u_arrmul24_and16_11_b_11;
  wire f_u_arrmul24_and16_11_y0;
  wire f_u_arrmul24_fa16_11_f_u_arrmul24_and16_11_y0;
  wire f_u_arrmul24_fa16_11_f_u_arrmul24_fa17_10_y2;
  wire f_u_arrmul24_fa16_11_y0;
  wire f_u_arrmul24_fa16_11_y1;
  wire f_u_arrmul24_fa16_11_f_u_arrmul24_fa15_11_y4;
  wire f_u_arrmul24_fa16_11_y2;
  wire f_u_arrmul24_fa16_11_y3;
  wire f_u_arrmul24_fa16_11_y4;
  wire f_u_arrmul24_and17_11_a_17;
  wire f_u_arrmul24_and17_11_b_11;
  wire f_u_arrmul24_and17_11_y0;
  wire f_u_arrmul24_fa17_11_f_u_arrmul24_and17_11_y0;
  wire f_u_arrmul24_fa17_11_f_u_arrmul24_fa18_10_y2;
  wire f_u_arrmul24_fa17_11_y0;
  wire f_u_arrmul24_fa17_11_y1;
  wire f_u_arrmul24_fa17_11_f_u_arrmul24_fa16_11_y4;
  wire f_u_arrmul24_fa17_11_y2;
  wire f_u_arrmul24_fa17_11_y3;
  wire f_u_arrmul24_fa17_11_y4;
  wire f_u_arrmul24_and18_11_a_18;
  wire f_u_arrmul24_and18_11_b_11;
  wire f_u_arrmul24_and18_11_y0;
  wire f_u_arrmul24_fa18_11_f_u_arrmul24_and18_11_y0;
  wire f_u_arrmul24_fa18_11_f_u_arrmul24_fa19_10_y2;
  wire f_u_arrmul24_fa18_11_y0;
  wire f_u_arrmul24_fa18_11_y1;
  wire f_u_arrmul24_fa18_11_f_u_arrmul24_fa17_11_y4;
  wire f_u_arrmul24_fa18_11_y2;
  wire f_u_arrmul24_fa18_11_y3;
  wire f_u_arrmul24_fa18_11_y4;
  wire f_u_arrmul24_and19_11_a_19;
  wire f_u_arrmul24_and19_11_b_11;
  wire f_u_arrmul24_and19_11_y0;
  wire f_u_arrmul24_fa19_11_f_u_arrmul24_and19_11_y0;
  wire f_u_arrmul24_fa19_11_f_u_arrmul24_fa20_10_y2;
  wire f_u_arrmul24_fa19_11_y0;
  wire f_u_arrmul24_fa19_11_y1;
  wire f_u_arrmul24_fa19_11_f_u_arrmul24_fa18_11_y4;
  wire f_u_arrmul24_fa19_11_y2;
  wire f_u_arrmul24_fa19_11_y3;
  wire f_u_arrmul24_fa19_11_y4;
  wire f_u_arrmul24_and20_11_a_20;
  wire f_u_arrmul24_and20_11_b_11;
  wire f_u_arrmul24_and20_11_y0;
  wire f_u_arrmul24_fa20_11_f_u_arrmul24_and20_11_y0;
  wire f_u_arrmul24_fa20_11_f_u_arrmul24_fa21_10_y2;
  wire f_u_arrmul24_fa20_11_y0;
  wire f_u_arrmul24_fa20_11_y1;
  wire f_u_arrmul24_fa20_11_f_u_arrmul24_fa19_11_y4;
  wire f_u_arrmul24_fa20_11_y2;
  wire f_u_arrmul24_fa20_11_y3;
  wire f_u_arrmul24_fa20_11_y4;
  wire f_u_arrmul24_and21_11_a_21;
  wire f_u_arrmul24_and21_11_b_11;
  wire f_u_arrmul24_and21_11_y0;
  wire f_u_arrmul24_fa21_11_f_u_arrmul24_and21_11_y0;
  wire f_u_arrmul24_fa21_11_f_u_arrmul24_fa22_10_y2;
  wire f_u_arrmul24_fa21_11_y0;
  wire f_u_arrmul24_fa21_11_y1;
  wire f_u_arrmul24_fa21_11_f_u_arrmul24_fa20_11_y4;
  wire f_u_arrmul24_fa21_11_y2;
  wire f_u_arrmul24_fa21_11_y3;
  wire f_u_arrmul24_fa21_11_y4;
  wire f_u_arrmul24_and22_11_a_22;
  wire f_u_arrmul24_and22_11_b_11;
  wire f_u_arrmul24_and22_11_y0;
  wire f_u_arrmul24_fa22_11_f_u_arrmul24_and22_11_y0;
  wire f_u_arrmul24_fa22_11_f_u_arrmul24_fa23_10_y2;
  wire f_u_arrmul24_fa22_11_y0;
  wire f_u_arrmul24_fa22_11_y1;
  wire f_u_arrmul24_fa22_11_f_u_arrmul24_fa21_11_y4;
  wire f_u_arrmul24_fa22_11_y2;
  wire f_u_arrmul24_fa22_11_y3;
  wire f_u_arrmul24_fa22_11_y4;
  wire f_u_arrmul24_and23_11_a_23;
  wire f_u_arrmul24_and23_11_b_11;
  wire f_u_arrmul24_and23_11_y0;
  wire f_u_arrmul24_fa23_11_f_u_arrmul24_and23_11_y0;
  wire f_u_arrmul24_fa23_11_f_u_arrmul24_fa23_10_y4;
  wire f_u_arrmul24_fa23_11_y0;
  wire f_u_arrmul24_fa23_11_y1;
  wire f_u_arrmul24_fa23_11_f_u_arrmul24_fa22_11_y4;
  wire f_u_arrmul24_fa23_11_y2;
  wire f_u_arrmul24_fa23_11_y3;
  wire f_u_arrmul24_fa23_11_y4;
  wire f_u_arrmul24_and0_12_a_0;
  wire f_u_arrmul24_and0_12_b_12;
  wire f_u_arrmul24_and0_12_y0;
  wire f_u_arrmul24_ha0_12_f_u_arrmul24_and0_12_y0;
  wire f_u_arrmul24_ha0_12_f_u_arrmul24_fa1_11_y2;
  wire f_u_arrmul24_ha0_12_y0;
  wire f_u_arrmul24_ha0_12_y1;
  wire f_u_arrmul24_and1_12_a_1;
  wire f_u_arrmul24_and1_12_b_12;
  wire f_u_arrmul24_and1_12_y0;
  wire f_u_arrmul24_fa1_12_f_u_arrmul24_and1_12_y0;
  wire f_u_arrmul24_fa1_12_f_u_arrmul24_fa2_11_y2;
  wire f_u_arrmul24_fa1_12_y0;
  wire f_u_arrmul24_fa1_12_y1;
  wire f_u_arrmul24_fa1_12_f_u_arrmul24_ha0_12_y1;
  wire f_u_arrmul24_fa1_12_y2;
  wire f_u_arrmul24_fa1_12_y3;
  wire f_u_arrmul24_fa1_12_y4;
  wire f_u_arrmul24_and2_12_a_2;
  wire f_u_arrmul24_and2_12_b_12;
  wire f_u_arrmul24_and2_12_y0;
  wire f_u_arrmul24_fa2_12_f_u_arrmul24_and2_12_y0;
  wire f_u_arrmul24_fa2_12_f_u_arrmul24_fa3_11_y2;
  wire f_u_arrmul24_fa2_12_y0;
  wire f_u_arrmul24_fa2_12_y1;
  wire f_u_arrmul24_fa2_12_f_u_arrmul24_fa1_12_y4;
  wire f_u_arrmul24_fa2_12_y2;
  wire f_u_arrmul24_fa2_12_y3;
  wire f_u_arrmul24_fa2_12_y4;
  wire f_u_arrmul24_and3_12_a_3;
  wire f_u_arrmul24_and3_12_b_12;
  wire f_u_arrmul24_and3_12_y0;
  wire f_u_arrmul24_fa3_12_f_u_arrmul24_and3_12_y0;
  wire f_u_arrmul24_fa3_12_f_u_arrmul24_fa4_11_y2;
  wire f_u_arrmul24_fa3_12_y0;
  wire f_u_arrmul24_fa3_12_y1;
  wire f_u_arrmul24_fa3_12_f_u_arrmul24_fa2_12_y4;
  wire f_u_arrmul24_fa3_12_y2;
  wire f_u_arrmul24_fa3_12_y3;
  wire f_u_arrmul24_fa3_12_y4;
  wire f_u_arrmul24_and4_12_a_4;
  wire f_u_arrmul24_and4_12_b_12;
  wire f_u_arrmul24_and4_12_y0;
  wire f_u_arrmul24_fa4_12_f_u_arrmul24_and4_12_y0;
  wire f_u_arrmul24_fa4_12_f_u_arrmul24_fa5_11_y2;
  wire f_u_arrmul24_fa4_12_y0;
  wire f_u_arrmul24_fa4_12_y1;
  wire f_u_arrmul24_fa4_12_f_u_arrmul24_fa3_12_y4;
  wire f_u_arrmul24_fa4_12_y2;
  wire f_u_arrmul24_fa4_12_y3;
  wire f_u_arrmul24_fa4_12_y4;
  wire f_u_arrmul24_and5_12_a_5;
  wire f_u_arrmul24_and5_12_b_12;
  wire f_u_arrmul24_and5_12_y0;
  wire f_u_arrmul24_fa5_12_f_u_arrmul24_and5_12_y0;
  wire f_u_arrmul24_fa5_12_f_u_arrmul24_fa6_11_y2;
  wire f_u_arrmul24_fa5_12_y0;
  wire f_u_arrmul24_fa5_12_y1;
  wire f_u_arrmul24_fa5_12_f_u_arrmul24_fa4_12_y4;
  wire f_u_arrmul24_fa5_12_y2;
  wire f_u_arrmul24_fa5_12_y3;
  wire f_u_arrmul24_fa5_12_y4;
  wire f_u_arrmul24_and6_12_a_6;
  wire f_u_arrmul24_and6_12_b_12;
  wire f_u_arrmul24_and6_12_y0;
  wire f_u_arrmul24_fa6_12_f_u_arrmul24_and6_12_y0;
  wire f_u_arrmul24_fa6_12_f_u_arrmul24_fa7_11_y2;
  wire f_u_arrmul24_fa6_12_y0;
  wire f_u_arrmul24_fa6_12_y1;
  wire f_u_arrmul24_fa6_12_f_u_arrmul24_fa5_12_y4;
  wire f_u_arrmul24_fa6_12_y2;
  wire f_u_arrmul24_fa6_12_y3;
  wire f_u_arrmul24_fa6_12_y4;
  wire f_u_arrmul24_and7_12_a_7;
  wire f_u_arrmul24_and7_12_b_12;
  wire f_u_arrmul24_and7_12_y0;
  wire f_u_arrmul24_fa7_12_f_u_arrmul24_and7_12_y0;
  wire f_u_arrmul24_fa7_12_f_u_arrmul24_fa8_11_y2;
  wire f_u_arrmul24_fa7_12_y0;
  wire f_u_arrmul24_fa7_12_y1;
  wire f_u_arrmul24_fa7_12_f_u_arrmul24_fa6_12_y4;
  wire f_u_arrmul24_fa7_12_y2;
  wire f_u_arrmul24_fa7_12_y3;
  wire f_u_arrmul24_fa7_12_y4;
  wire f_u_arrmul24_and8_12_a_8;
  wire f_u_arrmul24_and8_12_b_12;
  wire f_u_arrmul24_and8_12_y0;
  wire f_u_arrmul24_fa8_12_f_u_arrmul24_and8_12_y0;
  wire f_u_arrmul24_fa8_12_f_u_arrmul24_fa9_11_y2;
  wire f_u_arrmul24_fa8_12_y0;
  wire f_u_arrmul24_fa8_12_y1;
  wire f_u_arrmul24_fa8_12_f_u_arrmul24_fa7_12_y4;
  wire f_u_arrmul24_fa8_12_y2;
  wire f_u_arrmul24_fa8_12_y3;
  wire f_u_arrmul24_fa8_12_y4;
  wire f_u_arrmul24_and9_12_a_9;
  wire f_u_arrmul24_and9_12_b_12;
  wire f_u_arrmul24_and9_12_y0;
  wire f_u_arrmul24_fa9_12_f_u_arrmul24_and9_12_y0;
  wire f_u_arrmul24_fa9_12_f_u_arrmul24_fa10_11_y2;
  wire f_u_arrmul24_fa9_12_y0;
  wire f_u_arrmul24_fa9_12_y1;
  wire f_u_arrmul24_fa9_12_f_u_arrmul24_fa8_12_y4;
  wire f_u_arrmul24_fa9_12_y2;
  wire f_u_arrmul24_fa9_12_y3;
  wire f_u_arrmul24_fa9_12_y4;
  wire f_u_arrmul24_and10_12_a_10;
  wire f_u_arrmul24_and10_12_b_12;
  wire f_u_arrmul24_and10_12_y0;
  wire f_u_arrmul24_fa10_12_f_u_arrmul24_and10_12_y0;
  wire f_u_arrmul24_fa10_12_f_u_arrmul24_fa11_11_y2;
  wire f_u_arrmul24_fa10_12_y0;
  wire f_u_arrmul24_fa10_12_y1;
  wire f_u_arrmul24_fa10_12_f_u_arrmul24_fa9_12_y4;
  wire f_u_arrmul24_fa10_12_y2;
  wire f_u_arrmul24_fa10_12_y3;
  wire f_u_arrmul24_fa10_12_y4;
  wire f_u_arrmul24_and11_12_a_11;
  wire f_u_arrmul24_and11_12_b_12;
  wire f_u_arrmul24_and11_12_y0;
  wire f_u_arrmul24_fa11_12_f_u_arrmul24_and11_12_y0;
  wire f_u_arrmul24_fa11_12_f_u_arrmul24_fa12_11_y2;
  wire f_u_arrmul24_fa11_12_y0;
  wire f_u_arrmul24_fa11_12_y1;
  wire f_u_arrmul24_fa11_12_f_u_arrmul24_fa10_12_y4;
  wire f_u_arrmul24_fa11_12_y2;
  wire f_u_arrmul24_fa11_12_y3;
  wire f_u_arrmul24_fa11_12_y4;
  wire f_u_arrmul24_and12_12_a_12;
  wire f_u_arrmul24_and12_12_b_12;
  wire f_u_arrmul24_and12_12_y0;
  wire f_u_arrmul24_fa12_12_f_u_arrmul24_and12_12_y0;
  wire f_u_arrmul24_fa12_12_f_u_arrmul24_fa13_11_y2;
  wire f_u_arrmul24_fa12_12_y0;
  wire f_u_arrmul24_fa12_12_y1;
  wire f_u_arrmul24_fa12_12_f_u_arrmul24_fa11_12_y4;
  wire f_u_arrmul24_fa12_12_y2;
  wire f_u_arrmul24_fa12_12_y3;
  wire f_u_arrmul24_fa12_12_y4;
  wire f_u_arrmul24_and13_12_a_13;
  wire f_u_arrmul24_and13_12_b_12;
  wire f_u_arrmul24_and13_12_y0;
  wire f_u_arrmul24_fa13_12_f_u_arrmul24_and13_12_y0;
  wire f_u_arrmul24_fa13_12_f_u_arrmul24_fa14_11_y2;
  wire f_u_arrmul24_fa13_12_y0;
  wire f_u_arrmul24_fa13_12_y1;
  wire f_u_arrmul24_fa13_12_f_u_arrmul24_fa12_12_y4;
  wire f_u_arrmul24_fa13_12_y2;
  wire f_u_arrmul24_fa13_12_y3;
  wire f_u_arrmul24_fa13_12_y4;
  wire f_u_arrmul24_and14_12_a_14;
  wire f_u_arrmul24_and14_12_b_12;
  wire f_u_arrmul24_and14_12_y0;
  wire f_u_arrmul24_fa14_12_f_u_arrmul24_and14_12_y0;
  wire f_u_arrmul24_fa14_12_f_u_arrmul24_fa15_11_y2;
  wire f_u_arrmul24_fa14_12_y0;
  wire f_u_arrmul24_fa14_12_y1;
  wire f_u_arrmul24_fa14_12_f_u_arrmul24_fa13_12_y4;
  wire f_u_arrmul24_fa14_12_y2;
  wire f_u_arrmul24_fa14_12_y3;
  wire f_u_arrmul24_fa14_12_y4;
  wire f_u_arrmul24_and15_12_a_15;
  wire f_u_arrmul24_and15_12_b_12;
  wire f_u_arrmul24_and15_12_y0;
  wire f_u_arrmul24_fa15_12_f_u_arrmul24_and15_12_y0;
  wire f_u_arrmul24_fa15_12_f_u_arrmul24_fa16_11_y2;
  wire f_u_arrmul24_fa15_12_y0;
  wire f_u_arrmul24_fa15_12_y1;
  wire f_u_arrmul24_fa15_12_f_u_arrmul24_fa14_12_y4;
  wire f_u_arrmul24_fa15_12_y2;
  wire f_u_arrmul24_fa15_12_y3;
  wire f_u_arrmul24_fa15_12_y4;
  wire f_u_arrmul24_and16_12_a_16;
  wire f_u_arrmul24_and16_12_b_12;
  wire f_u_arrmul24_and16_12_y0;
  wire f_u_arrmul24_fa16_12_f_u_arrmul24_and16_12_y0;
  wire f_u_arrmul24_fa16_12_f_u_arrmul24_fa17_11_y2;
  wire f_u_arrmul24_fa16_12_y0;
  wire f_u_arrmul24_fa16_12_y1;
  wire f_u_arrmul24_fa16_12_f_u_arrmul24_fa15_12_y4;
  wire f_u_arrmul24_fa16_12_y2;
  wire f_u_arrmul24_fa16_12_y3;
  wire f_u_arrmul24_fa16_12_y4;
  wire f_u_arrmul24_and17_12_a_17;
  wire f_u_arrmul24_and17_12_b_12;
  wire f_u_arrmul24_and17_12_y0;
  wire f_u_arrmul24_fa17_12_f_u_arrmul24_and17_12_y0;
  wire f_u_arrmul24_fa17_12_f_u_arrmul24_fa18_11_y2;
  wire f_u_arrmul24_fa17_12_y0;
  wire f_u_arrmul24_fa17_12_y1;
  wire f_u_arrmul24_fa17_12_f_u_arrmul24_fa16_12_y4;
  wire f_u_arrmul24_fa17_12_y2;
  wire f_u_arrmul24_fa17_12_y3;
  wire f_u_arrmul24_fa17_12_y4;
  wire f_u_arrmul24_and18_12_a_18;
  wire f_u_arrmul24_and18_12_b_12;
  wire f_u_arrmul24_and18_12_y0;
  wire f_u_arrmul24_fa18_12_f_u_arrmul24_and18_12_y0;
  wire f_u_arrmul24_fa18_12_f_u_arrmul24_fa19_11_y2;
  wire f_u_arrmul24_fa18_12_y0;
  wire f_u_arrmul24_fa18_12_y1;
  wire f_u_arrmul24_fa18_12_f_u_arrmul24_fa17_12_y4;
  wire f_u_arrmul24_fa18_12_y2;
  wire f_u_arrmul24_fa18_12_y3;
  wire f_u_arrmul24_fa18_12_y4;
  wire f_u_arrmul24_and19_12_a_19;
  wire f_u_arrmul24_and19_12_b_12;
  wire f_u_arrmul24_and19_12_y0;
  wire f_u_arrmul24_fa19_12_f_u_arrmul24_and19_12_y0;
  wire f_u_arrmul24_fa19_12_f_u_arrmul24_fa20_11_y2;
  wire f_u_arrmul24_fa19_12_y0;
  wire f_u_arrmul24_fa19_12_y1;
  wire f_u_arrmul24_fa19_12_f_u_arrmul24_fa18_12_y4;
  wire f_u_arrmul24_fa19_12_y2;
  wire f_u_arrmul24_fa19_12_y3;
  wire f_u_arrmul24_fa19_12_y4;
  wire f_u_arrmul24_and20_12_a_20;
  wire f_u_arrmul24_and20_12_b_12;
  wire f_u_arrmul24_and20_12_y0;
  wire f_u_arrmul24_fa20_12_f_u_arrmul24_and20_12_y0;
  wire f_u_arrmul24_fa20_12_f_u_arrmul24_fa21_11_y2;
  wire f_u_arrmul24_fa20_12_y0;
  wire f_u_arrmul24_fa20_12_y1;
  wire f_u_arrmul24_fa20_12_f_u_arrmul24_fa19_12_y4;
  wire f_u_arrmul24_fa20_12_y2;
  wire f_u_arrmul24_fa20_12_y3;
  wire f_u_arrmul24_fa20_12_y4;
  wire f_u_arrmul24_and21_12_a_21;
  wire f_u_arrmul24_and21_12_b_12;
  wire f_u_arrmul24_and21_12_y0;
  wire f_u_arrmul24_fa21_12_f_u_arrmul24_and21_12_y0;
  wire f_u_arrmul24_fa21_12_f_u_arrmul24_fa22_11_y2;
  wire f_u_arrmul24_fa21_12_y0;
  wire f_u_arrmul24_fa21_12_y1;
  wire f_u_arrmul24_fa21_12_f_u_arrmul24_fa20_12_y4;
  wire f_u_arrmul24_fa21_12_y2;
  wire f_u_arrmul24_fa21_12_y3;
  wire f_u_arrmul24_fa21_12_y4;
  wire f_u_arrmul24_and22_12_a_22;
  wire f_u_arrmul24_and22_12_b_12;
  wire f_u_arrmul24_and22_12_y0;
  wire f_u_arrmul24_fa22_12_f_u_arrmul24_and22_12_y0;
  wire f_u_arrmul24_fa22_12_f_u_arrmul24_fa23_11_y2;
  wire f_u_arrmul24_fa22_12_y0;
  wire f_u_arrmul24_fa22_12_y1;
  wire f_u_arrmul24_fa22_12_f_u_arrmul24_fa21_12_y4;
  wire f_u_arrmul24_fa22_12_y2;
  wire f_u_arrmul24_fa22_12_y3;
  wire f_u_arrmul24_fa22_12_y4;
  wire f_u_arrmul24_and23_12_a_23;
  wire f_u_arrmul24_and23_12_b_12;
  wire f_u_arrmul24_and23_12_y0;
  wire f_u_arrmul24_fa23_12_f_u_arrmul24_and23_12_y0;
  wire f_u_arrmul24_fa23_12_f_u_arrmul24_fa23_11_y4;
  wire f_u_arrmul24_fa23_12_y0;
  wire f_u_arrmul24_fa23_12_y1;
  wire f_u_arrmul24_fa23_12_f_u_arrmul24_fa22_12_y4;
  wire f_u_arrmul24_fa23_12_y2;
  wire f_u_arrmul24_fa23_12_y3;
  wire f_u_arrmul24_fa23_12_y4;
  wire f_u_arrmul24_and0_13_a_0;
  wire f_u_arrmul24_and0_13_b_13;
  wire f_u_arrmul24_and0_13_y0;
  wire f_u_arrmul24_ha0_13_f_u_arrmul24_and0_13_y0;
  wire f_u_arrmul24_ha0_13_f_u_arrmul24_fa1_12_y2;
  wire f_u_arrmul24_ha0_13_y0;
  wire f_u_arrmul24_ha0_13_y1;
  wire f_u_arrmul24_and1_13_a_1;
  wire f_u_arrmul24_and1_13_b_13;
  wire f_u_arrmul24_and1_13_y0;
  wire f_u_arrmul24_fa1_13_f_u_arrmul24_and1_13_y0;
  wire f_u_arrmul24_fa1_13_f_u_arrmul24_fa2_12_y2;
  wire f_u_arrmul24_fa1_13_y0;
  wire f_u_arrmul24_fa1_13_y1;
  wire f_u_arrmul24_fa1_13_f_u_arrmul24_ha0_13_y1;
  wire f_u_arrmul24_fa1_13_y2;
  wire f_u_arrmul24_fa1_13_y3;
  wire f_u_arrmul24_fa1_13_y4;
  wire f_u_arrmul24_and2_13_a_2;
  wire f_u_arrmul24_and2_13_b_13;
  wire f_u_arrmul24_and2_13_y0;
  wire f_u_arrmul24_fa2_13_f_u_arrmul24_and2_13_y0;
  wire f_u_arrmul24_fa2_13_f_u_arrmul24_fa3_12_y2;
  wire f_u_arrmul24_fa2_13_y0;
  wire f_u_arrmul24_fa2_13_y1;
  wire f_u_arrmul24_fa2_13_f_u_arrmul24_fa1_13_y4;
  wire f_u_arrmul24_fa2_13_y2;
  wire f_u_arrmul24_fa2_13_y3;
  wire f_u_arrmul24_fa2_13_y4;
  wire f_u_arrmul24_and3_13_a_3;
  wire f_u_arrmul24_and3_13_b_13;
  wire f_u_arrmul24_and3_13_y0;
  wire f_u_arrmul24_fa3_13_f_u_arrmul24_and3_13_y0;
  wire f_u_arrmul24_fa3_13_f_u_arrmul24_fa4_12_y2;
  wire f_u_arrmul24_fa3_13_y0;
  wire f_u_arrmul24_fa3_13_y1;
  wire f_u_arrmul24_fa3_13_f_u_arrmul24_fa2_13_y4;
  wire f_u_arrmul24_fa3_13_y2;
  wire f_u_arrmul24_fa3_13_y3;
  wire f_u_arrmul24_fa3_13_y4;
  wire f_u_arrmul24_and4_13_a_4;
  wire f_u_arrmul24_and4_13_b_13;
  wire f_u_arrmul24_and4_13_y0;
  wire f_u_arrmul24_fa4_13_f_u_arrmul24_and4_13_y0;
  wire f_u_arrmul24_fa4_13_f_u_arrmul24_fa5_12_y2;
  wire f_u_arrmul24_fa4_13_y0;
  wire f_u_arrmul24_fa4_13_y1;
  wire f_u_arrmul24_fa4_13_f_u_arrmul24_fa3_13_y4;
  wire f_u_arrmul24_fa4_13_y2;
  wire f_u_arrmul24_fa4_13_y3;
  wire f_u_arrmul24_fa4_13_y4;
  wire f_u_arrmul24_and5_13_a_5;
  wire f_u_arrmul24_and5_13_b_13;
  wire f_u_arrmul24_and5_13_y0;
  wire f_u_arrmul24_fa5_13_f_u_arrmul24_and5_13_y0;
  wire f_u_arrmul24_fa5_13_f_u_arrmul24_fa6_12_y2;
  wire f_u_arrmul24_fa5_13_y0;
  wire f_u_arrmul24_fa5_13_y1;
  wire f_u_arrmul24_fa5_13_f_u_arrmul24_fa4_13_y4;
  wire f_u_arrmul24_fa5_13_y2;
  wire f_u_arrmul24_fa5_13_y3;
  wire f_u_arrmul24_fa5_13_y4;
  wire f_u_arrmul24_and6_13_a_6;
  wire f_u_arrmul24_and6_13_b_13;
  wire f_u_arrmul24_and6_13_y0;
  wire f_u_arrmul24_fa6_13_f_u_arrmul24_and6_13_y0;
  wire f_u_arrmul24_fa6_13_f_u_arrmul24_fa7_12_y2;
  wire f_u_arrmul24_fa6_13_y0;
  wire f_u_arrmul24_fa6_13_y1;
  wire f_u_arrmul24_fa6_13_f_u_arrmul24_fa5_13_y4;
  wire f_u_arrmul24_fa6_13_y2;
  wire f_u_arrmul24_fa6_13_y3;
  wire f_u_arrmul24_fa6_13_y4;
  wire f_u_arrmul24_and7_13_a_7;
  wire f_u_arrmul24_and7_13_b_13;
  wire f_u_arrmul24_and7_13_y0;
  wire f_u_arrmul24_fa7_13_f_u_arrmul24_and7_13_y0;
  wire f_u_arrmul24_fa7_13_f_u_arrmul24_fa8_12_y2;
  wire f_u_arrmul24_fa7_13_y0;
  wire f_u_arrmul24_fa7_13_y1;
  wire f_u_arrmul24_fa7_13_f_u_arrmul24_fa6_13_y4;
  wire f_u_arrmul24_fa7_13_y2;
  wire f_u_arrmul24_fa7_13_y3;
  wire f_u_arrmul24_fa7_13_y4;
  wire f_u_arrmul24_and8_13_a_8;
  wire f_u_arrmul24_and8_13_b_13;
  wire f_u_arrmul24_and8_13_y0;
  wire f_u_arrmul24_fa8_13_f_u_arrmul24_and8_13_y0;
  wire f_u_arrmul24_fa8_13_f_u_arrmul24_fa9_12_y2;
  wire f_u_arrmul24_fa8_13_y0;
  wire f_u_arrmul24_fa8_13_y1;
  wire f_u_arrmul24_fa8_13_f_u_arrmul24_fa7_13_y4;
  wire f_u_arrmul24_fa8_13_y2;
  wire f_u_arrmul24_fa8_13_y3;
  wire f_u_arrmul24_fa8_13_y4;
  wire f_u_arrmul24_and9_13_a_9;
  wire f_u_arrmul24_and9_13_b_13;
  wire f_u_arrmul24_and9_13_y0;
  wire f_u_arrmul24_fa9_13_f_u_arrmul24_and9_13_y0;
  wire f_u_arrmul24_fa9_13_f_u_arrmul24_fa10_12_y2;
  wire f_u_arrmul24_fa9_13_y0;
  wire f_u_arrmul24_fa9_13_y1;
  wire f_u_arrmul24_fa9_13_f_u_arrmul24_fa8_13_y4;
  wire f_u_arrmul24_fa9_13_y2;
  wire f_u_arrmul24_fa9_13_y3;
  wire f_u_arrmul24_fa9_13_y4;
  wire f_u_arrmul24_and10_13_a_10;
  wire f_u_arrmul24_and10_13_b_13;
  wire f_u_arrmul24_and10_13_y0;
  wire f_u_arrmul24_fa10_13_f_u_arrmul24_and10_13_y0;
  wire f_u_arrmul24_fa10_13_f_u_arrmul24_fa11_12_y2;
  wire f_u_arrmul24_fa10_13_y0;
  wire f_u_arrmul24_fa10_13_y1;
  wire f_u_arrmul24_fa10_13_f_u_arrmul24_fa9_13_y4;
  wire f_u_arrmul24_fa10_13_y2;
  wire f_u_arrmul24_fa10_13_y3;
  wire f_u_arrmul24_fa10_13_y4;
  wire f_u_arrmul24_and11_13_a_11;
  wire f_u_arrmul24_and11_13_b_13;
  wire f_u_arrmul24_and11_13_y0;
  wire f_u_arrmul24_fa11_13_f_u_arrmul24_and11_13_y0;
  wire f_u_arrmul24_fa11_13_f_u_arrmul24_fa12_12_y2;
  wire f_u_arrmul24_fa11_13_y0;
  wire f_u_arrmul24_fa11_13_y1;
  wire f_u_arrmul24_fa11_13_f_u_arrmul24_fa10_13_y4;
  wire f_u_arrmul24_fa11_13_y2;
  wire f_u_arrmul24_fa11_13_y3;
  wire f_u_arrmul24_fa11_13_y4;
  wire f_u_arrmul24_and12_13_a_12;
  wire f_u_arrmul24_and12_13_b_13;
  wire f_u_arrmul24_and12_13_y0;
  wire f_u_arrmul24_fa12_13_f_u_arrmul24_and12_13_y0;
  wire f_u_arrmul24_fa12_13_f_u_arrmul24_fa13_12_y2;
  wire f_u_arrmul24_fa12_13_y0;
  wire f_u_arrmul24_fa12_13_y1;
  wire f_u_arrmul24_fa12_13_f_u_arrmul24_fa11_13_y4;
  wire f_u_arrmul24_fa12_13_y2;
  wire f_u_arrmul24_fa12_13_y3;
  wire f_u_arrmul24_fa12_13_y4;
  wire f_u_arrmul24_and13_13_a_13;
  wire f_u_arrmul24_and13_13_b_13;
  wire f_u_arrmul24_and13_13_y0;
  wire f_u_arrmul24_fa13_13_f_u_arrmul24_and13_13_y0;
  wire f_u_arrmul24_fa13_13_f_u_arrmul24_fa14_12_y2;
  wire f_u_arrmul24_fa13_13_y0;
  wire f_u_arrmul24_fa13_13_y1;
  wire f_u_arrmul24_fa13_13_f_u_arrmul24_fa12_13_y4;
  wire f_u_arrmul24_fa13_13_y2;
  wire f_u_arrmul24_fa13_13_y3;
  wire f_u_arrmul24_fa13_13_y4;
  wire f_u_arrmul24_and14_13_a_14;
  wire f_u_arrmul24_and14_13_b_13;
  wire f_u_arrmul24_and14_13_y0;
  wire f_u_arrmul24_fa14_13_f_u_arrmul24_and14_13_y0;
  wire f_u_arrmul24_fa14_13_f_u_arrmul24_fa15_12_y2;
  wire f_u_arrmul24_fa14_13_y0;
  wire f_u_arrmul24_fa14_13_y1;
  wire f_u_arrmul24_fa14_13_f_u_arrmul24_fa13_13_y4;
  wire f_u_arrmul24_fa14_13_y2;
  wire f_u_arrmul24_fa14_13_y3;
  wire f_u_arrmul24_fa14_13_y4;
  wire f_u_arrmul24_and15_13_a_15;
  wire f_u_arrmul24_and15_13_b_13;
  wire f_u_arrmul24_and15_13_y0;
  wire f_u_arrmul24_fa15_13_f_u_arrmul24_and15_13_y0;
  wire f_u_arrmul24_fa15_13_f_u_arrmul24_fa16_12_y2;
  wire f_u_arrmul24_fa15_13_y0;
  wire f_u_arrmul24_fa15_13_y1;
  wire f_u_arrmul24_fa15_13_f_u_arrmul24_fa14_13_y4;
  wire f_u_arrmul24_fa15_13_y2;
  wire f_u_arrmul24_fa15_13_y3;
  wire f_u_arrmul24_fa15_13_y4;
  wire f_u_arrmul24_and16_13_a_16;
  wire f_u_arrmul24_and16_13_b_13;
  wire f_u_arrmul24_and16_13_y0;
  wire f_u_arrmul24_fa16_13_f_u_arrmul24_and16_13_y0;
  wire f_u_arrmul24_fa16_13_f_u_arrmul24_fa17_12_y2;
  wire f_u_arrmul24_fa16_13_y0;
  wire f_u_arrmul24_fa16_13_y1;
  wire f_u_arrmul24_fa16_13_f_u_arrmul24_fa15_13_y4;
  wire f_u_arrmul24_fa16_13_y2;
  wire f_u_arrmul24_fa16_13_y3;
  wire f_u_arrmul24_fa16_13_y4;
  wire f_u_arrmul24_and17_13_a_17;
  wire f_u_arrmul24_and17_13_b_13;
  wire f_u_arrmul24_and17_13_y0;
  wire f_u_arrmul24_fa17_13_f_u_arrmul24_and17_13_y0;
  wire f_u_arrmul24_fa17_13_f_u_arrmul24_fa18_12_y2;
  wire f_u_arrmul24_fa17_13_y0;
  wire f_u_arrmul24_fa17_13_y1;
  wire f_u_arrmul24_fa17_13_f_u_arrmul24_fa16_13_y4;
  wire f_u_arrmul24_fa17_13_y2;
  wire f_u_arrmul24_fa17_13_y3;
  wire f_u_arrmul24_fa17_13_y4;
  wire f_u_arrmul24_and18_13_a_18;
  wire f_u_arrmul24_and18_13_b_13;
  wire f_u_arrmul24_and18_13_y0;
  wire f_u_arrmul24_fa18_13_f_u_arrmul24_and18_13_y0;
  wire f_u_arrmul24_fa18_13_f_u_arrmul24_fa19_12_y2;
  wire f_u_arrmul24_fa18_13_y0;
  wire f_u_arrmul24_fa18_13_y1;
  wire f_u_arrmul24_fa18_13_f_u_arrmul24_fa17_13_y4;
  wire f_u_arrmul24_fa18_13_y2;
  wire f_u_arrmul24_fa18_13_y3;
  wire f_u_arrmul24_fa18_13_y4;
  wire f_u_arrmul24_and19_13_a_19;
  wire f_u_arrmul24_and19_13_b_13;
  wire f_u_arrmul24_and19_13_y0;
  wire f_u_arrmul24_fa19_13_f_u_arrmul24_and19_13_y0;
  wire f_u_arrmul24_fa19_13_f_u_arrmul24_fa20_12_y2;
  wire f_u_arrmul24_fa19_13_y0;
  wire f_u_arrmul24_fa19_13_y1;
  wire f_u_arrmul24_fa19_13_f_u_arrmul24_fa18_13_y4;
  wire f_u_arrmul24_fa19_13_y2;
  wire f_u_arrmul24_fa19_13_y3;
  wire f_u_arrmul24_fa19_13_y4;
  wire f_u_arrmul24_and20_13_a_20;
  wire f_u_arrmul24_and20_13_b_13;
  wire f_u_arrmul24_and20_13_y0;
  wire f_u_arrmul24_fa20_13_f_u_arrmul24_and20_13_y0;
  wire f_u_arrmul24_fa20_13_f_u_arrmul24_fa21_12_y2;
  wire f_u_arrmul24_fa20_13_y0;
  wire f_u_arrmul24_fa20_13_y1;
  wire f_u_arrmul24_fa20_13_f_u_arrmul24_fa19_13_y4;
  wire f_u_arrmul24_fa20_13_y2;
  wire f_u_arrmul24_fa20_13_y3;
  wire f_u_arrmul24_fa20_13_y4;
  wire f_u_arrmul24_and21_13_a_21;
  wire f_u_arrmul24_and21_13_b_13;
  wire f_u_arrmul24_and21_13_y0;
  wire f_u_arrmul24_fa21_13_f_u_arrmul24_and21_13_y0;
  wire f_u_arrmul24_fa21_13_f_u_arrmul24_fa22_12_y2;
  wire f_u_arrmul24_fa21_13_y0;
  wire f_u_arrmul24_fa21_13_y1;
  wire f_u_arrmul24_fa21_13_f_u_arrmul24_fa20_13_y4;
  wire f_u_arrmul24_fa21_13_y2;
  wire f_u_arrmul24_fa21_13_y3;
  wire f_u_arrmul24_fa21_13_y4;
  wire f_u_arrmul24_and22_13_a_22;
  wire f_u_arrmul24_and22_13_b_13;
  wire f_u_arrmul24_and22_13_y0;
  wire f_u_arrmul24_fa22_13_f_u_arrmul24_and22_13_y0;
  wire f_u_arrmul24_fa22_13_f_u_arrmul24_fa23_12_y2;
  wire f_u_arrmul24_fa22_13_y0;
  wire f_u_arrmul24_fa22_13_y1;
  wire f_u_arrmul24_fa22_13_f_u_arrmul24_fa21_13_y4;
  wire f_u_arrmul24_fa22_13_y2;
  wire f_u_arrmul24_fa22_13_y3;
  wire f_u_arrmul24_fa22_13_y4;
  wire f_u_arrmul24_and23_13_a_23;
  wire f_u_arrmul24_and23_13_b_13;
  wire f_u_arrmul24_and23_13_y0;
  wire f_u_arrmul24_fa23_13_f_u_arrmul24_and23_13_y0;
  wire f_u_arrmul24_fa23_13_f_u_arrmul24_fa23_12_y4;
  wire f_u_arrmul24_fa23_13_y0;
  wire f_u_arrmul24_fa23_13_y1;
  wire f_u_arrmul24_fa23_13_f_u_arrmul24_fa22_13_y4;
  wire f_u_arrmul24_fa23_13_y2;
  wire f_u_arrmul24_fa23_13_y3;
  wire f_u_arrmul24_fa23_13_y4;
  wire f_u_arrmul24_and0_14_a_0;
  wire f_u_arrmul24_and0_14_b_14;
  wire f_u_arrmul24_and0_14_y0;
  wire f_u_arrmul24_ha0_14_f_u_arrmul24_and0_14_y0;
  wire f_u_arrmul24_ha0_14_f_u_arrmul24_fa1_13_y2;
  wire f_u_arrmul24_ha0_14_y0;
  wire f_u_arrmul24_ha0_14_y1;
  wire f_u_arrmul24_and1_14_a_1;
  wire f_u_arrmul24_and1_14_b_14;
  wire f_u_arrmul24_and1_14_y0;
  wire f_u_arrmul24_fa1_14_f_u_arrmul24_and1_14_y0;
  wire f_u_arrmul24_fa1_14_f_u_arrmul24_fa2_13_y2;
  wire f_u_arrmul24_fa1_14_y0;
  wire f_u_arrmul24_fa1_14_y1;
  wire f_u_arrmul24_fa1_14_f_u_arrmul24_ha0_14_y1;
  wire f_u_arrmul24_fa1_14_y2;
  wire f_u_arrmul24_fa1_14_y3;
  wire f_u_arrmul24_fa1_14_y4;
  wire f_u_arrmul24_and2_14_a_2;
  wire f_u_arrmul24_and2_14_b_14;
  wire f_u_arrmul24_and2_14_y0;
  wire f_u_arrmul24_fa2_14_f_u_arrmul24_and2_14_y0;
  wire f_u_arrmul24_fa2_14_f_u_arrmul24_fa3_13_y2;
  wire f_u_arrmul24_fa2_14_y0;
  wire f_u_arrmul24_fa2_14_y1;
  wire f_u_arrmul24_fa2_14_f_u_arrmul24_fa1_14_y4;
  wire f_u_arrmul24_fa2_14_y2;
  wire f_u_arrmul24_fa2_14_y3;
  wire f_u_arrmul24_fa2_14_y4;
  wire f_u_arrmul24_and3_14_a_3;
  wire f_u_arrmul24_and3_14_b_14;
  wire f_u_arrmul24_and3_14_y0;
  wire f_u_arrmul24_fa3_14_f_u_arrmul24_and3_14_y0;
  wire f_u_arrmul24_fa3_14_f_u_arrmul24_fa4_13_y2;
  wire f_u_arrmul24_fa3_14_y0;
  wire f_u_arrmul24_fa3_14_y1;
  wire f_u_arrmul24_fa3_14_f_u_arrmul24_fa2_14_y4;
  wire f_u_arrmul24_fa3_14_y2;
  wire f_u_arrmul24_fa3_14_y3;
  wire f_u_arrmul24_fa3_14_y4;
  wire f_u_arrmul24_and4_14_a_4;
  wire f_u_arrmul24_and4_14_b_14;
  wire f_u_arrmul24_and4_14_y0;
  wire f_u_arrmul24_fa4_14_f_u_arrmul24_and4_14_y0;
  wire f_u_arrmul24_fa4_14_f_u_arrmul24_fa5_13_y2;
  wire f_u_arrmul24_fa4_14_y0;
  wire f_u_arrmul24_fa4_14_y1;
  wire f_u_arrmul24_fa4_14_f_u_arrmul24_fa3_14_y4;
  wire f_u_arrmul24_fa4_14_y2;
  wire f_u_arrmul24_fa4_14_y3;
  wire f_u_arrmul24_fa4_14_y4;
  wire f_u_arrmul24_and5_14_a_5;
  wire f_u_arrmul24_and5_14_b_14;
  wire f_u_arrmul24_and5_14_y0;
  wire f_u_arrmul24_fa5_14_f_u_arrmul24_and5_14_y0;
  wire f_u_arrmul24_fa5_14_f_u_arrmul24_fa6_13_y2;
  wire f_u_arrmul24_fa5_14_y0;
  wire f_u_arrmul24_fa5_14_y1;
  wire f_u_arrmul24_fa5_14_f_u_arrmul24_fa4_14_y4;
  wire f_u_arrmul24_fa5_14_y2;
  wire f_u_arrmul24_fa5_14_y3;
  wire f_u_arrmul24_fa5_14_y4;
  wire f_u_arrmul24_and6_14_a_6;
  wire f_u_arrmul24_and6_14_b_14;
  wire f_u_arrmul24_and6_14_y0;
  wire f_u_arrmul24_fa6_14_f_u_arrmul24_and6_14_y0;
  wire f_u_arrmul24_fa6_14_f_u_arrmul24_fa7_13_y2;
  wire f_u_arrmul24_fa6_14_y0;
  wire f_u_arrmul24_fa6_14_y1;
  wire f_u_arrmul24_fa6_14_f_u_arrmul24_fa5_14_y4;
  wire f_u_arrmul24_fa6_14_y2;
  wire f_u_arrmul24_fa6_14_y3;
  wire f_u_arrmul24_fa6_14_y4;
  wire f_u_arrmul24_and7_14_a_7;
  wire f_u_arrmul24_and7_14_b_14;
  wire f_u_arrmul24_and7_14_y0;
  wire f_u_arrmul24_fa7_14_f_u_arrmul24_and7_14_y0;
  wire f_u_arrmul24_fa7_14_f_u_arrmul24_fa8_13_y2;
  wire f_u_arrmul24_fa7_14_y0;
  wire f_u_arrmul24_fa7_14_y1;
  wire f_u_arrmul24_fa7_14_f_u_arrmul24_fa6_14_y4;
  wire f_u_arrmul24_fa7_14_y2;
  wire f_u_arrmul24_fa7_14_y3;
  wire f_u_arrmul24_fa7_14_y4;
  wire f_u_arrmul24_and8_14_a_8;
  wire f_u_arrmul24_and8_14_b_14;
  wire f_u_arrmul24_and8_14_y0;
  wire f_u_arrmul24_fa8_14_f_u_arrmul24_and8_14_y0;
  wire f_u_arrmul24_fa8_14_f_u_arrmul24_fa9_13_y2;
  wire f_u_arrmul24_fa8_14_y0;
  wire f_u_arrmul24_fa8_14_y1;
  wire f_u_arrmul24_fa8_14_f_u_arrmul24_fa7_14_y4;
  wire f_u_arrmul24_fa8_14_y2;
  wire f_u_arrmul24_fa8_14_y3;
  wire f_u_arrmul24_fa8_14_y4;
  wire f_u_arrmul24_and9_14_a_9;
  wire f_u_arrmul24_and9_14_b_14;
  wire f_u_arrmul24_and9_14_y0;
  wire f_u_arrmul24_fa9_14_f_u_arrmul24_and9_14_y0;
  wire f_u_arrmul24_fa9_14_f_u_arrmul24_fa10_13_y2;
  wire f_u_arrmul24_fa9_14_y0;
  wire f_u_arrmul24_fa9_14_y1;
  wire f_u_arrmul24_fa9_14_f_u_arrmul24_fa8_14_y4;
  wire f_u_arrmul24_fa9_14_y2;
  wire f_u_arrmul24_fa9_14_y3;
  wire f_u_arrmul24_fa9_14_y4;
  wire f_u_arrmul24_and10_14_a_10;
  wire f_u_arrmul24_and10_14_b_14;
  wire f_u_arrmul24_and10_14_y0;
  wire f_u_arrmul24_fa10_14_f_u_arrmul24_and10_14_y0;
  wire f_u_arrmul24_fa10_14_f_u_arrmul24_fa11_13_y2;
  wire f_u_arrmul24_fa10_14_y0;
  wire f_u_arrmul24_fa10_14_y1;
  wire f_u_arrmul24_fa10_14_f_u_arrmul24_fa9_14_y4;
  wire f_u_arrmul24_fa10_14_y2;
  wire f_u_arrmul24_fa10_14_y3;
  wire f_u_arrmul24_fa10_14_y4;
  wire f_u_arrmul24_and11_14_a_11;
  wire f_u_arrmul24_and11_14_b_14;
  wire f_u_arrmul24_and11_14_y0;
  wire f_u_arrmul24_fa11_14_f_u_arrmul24_and11_14_y0;
  wire f_u_arrmul24_fa11_14_f_u_arrmul24_fa12_13_y2;
  wire f_u_arrmul24_fa11_14_y0;
  wire f_u_arrmul24_fa11_14_y1;
  wire f_u_arrmul24_fa11_14_f_u_arrmul24_fa10_14_y4;
  wire f_u_arrmul24_fa11_14_y2;
  wire f_u_arrmul24_fa11_14_y3;
  wire f_u_arrmul24_fa11_14_y4;
  wire f_u_arrmul24_and12_14_a_12;
  wire f_u_arrmul24_and12_14_b_14;
  wire f_u_arrmul24_and12_14_y0;
  wire f_u_arrmul24_fa12_14_f_u_arrmul24_and12_14_y0;
  wire f_u_arrmul24_fa12_14_f_u_arrmul24_fa13_13_y2;
  wire f_u_arrmul24_fa12_14_y0;
  wire f_u_arrmul24_fa12_14_y1;
  wire f_u_arrmul24_fa12_14_f_u_arrmul24_fa11_14_y4;
  wire f_u_arrmul24_fa12_14_y2;
  wire f_u_arrmul24_fa12_14_y3;
  wire f_u_arrmul24_fa12_14_y4;
  wire f_u_arrmul24_and13_14_a_13;
  wire f_u_arrmul24_and13_14_b_14;
  wire f_u_arrmul24_and13_14_y0;
  wire f_u_arrmul24_fa13_14_f_u_arrmul24_and13_14_y0;
  wire f_u_arrmul24_fa13_14_f_u_arrmul24_fa14_13_y2;
  wire f_u_arrmul24_fa13_14_y0;
  wire f_u_arrmul24_fa13_14_y1;
  wire f_u_arrmul24_fa13_14_f_u_arrmul24_fa12_14_y4;
  wire f_u_arrmul24_fa13_14_y2;
  wire f_u_arrmul24_fa13_14_y3;
  wire f_u_arrmul24_fa13_14_y4;
  wire f_u_arrmul24_and14_14_a_14;
  wire f_u_arrmul24_and14_14_b_14;
  wire f_u_arrmul24_and14_14_y0;
  wire f_u_arrmul24_fa14_14_f_u_arrmul24_and14_14_y0;
  wire f_u_arrmul24_fa14_14_f_u_arrmul24_fa15_13_y2;
  wire f_u_arrmul24_fa14_14_y0;
  wire f_u_arrmul24_fa14_14_y1;
  wire f_u_arrmul24_fa14_14_f_u_arrmul24_fa13_14_y4;
  wire f_u_arrmul24_fa14_14_y2;
  wire f_u_arrmul24_fa14_14_y3;
  wire f_u_arrmul24_fa14_14_y4;
  wire f_u_arrmul24_and15_14_a_15;
  wire f_u_arrmul24_and15_14_b_14;
  wire f_u_arrmul24_and15_14_y0;
  wire f_u_arrmul24_fa15_14_f_u_arrmul24_and15_14_y0;
  wire f_u_arrmul24_fa15_14_f_u_arrmul24_fa16_13_y2;
  wire f_u_arrmul24_fa15_14_y0;
  wire f_u_arrmul24_fa15_14_y1;
  wire f_u_arrmul24_fa15_14_f_u_arrmul24_fa14_14_y4;
  wire f_u_arrmul24_fa15_14_y2;
  wire f_u_arrmul24_fa15_14_y3;
  wire f_u_arrmul24_fa15_14_y4;
  wire f_u_arrmul24_and16_14_a_16;
  wire f_u_arrmul24_and16_14_b_14;
  wire f_u_arrmul24_and16_14_y0;
  wire f_u_arrmul24_fa16_14_f_u_arrmul24_and16_14_y0;
  wire f_u_arrmul24_fa16_14_f_u_arrmul24_fa17_13_y2;
  wire f_u_arrmul24_fa16_14_y0;
  wire f_u_arrmul24_fa16_14_y1;
  wire f_u_arrmul24_fa16_14_f_u_arrmul24_fa15_14_y4;
  wire f_u_arrmul24_fa16_14_y2;
  wire f_u_arrmul24_fa16_14_y3;
  wire f_u_arrmul24_fa16_14_y4;
  wire f_u_arrmul24_and17_14_a_17;
  wire f_u_arrmul24_and17_14_b_14;
  wire f_u_arrmul24_and17_14_y0;
  wire f_u_arrmul24_fa17_14_f_u_arrmul24_and17_14_y0;
  wire f_u_arrmul24_fa17_14_f_u_arrmul24_fa18_13_y2;
  wire f_u_arrmul24_fa17_14_y0;
  wire f_u_arrmul24_fa17_14_y1;
  wire f_u_arrmul24_fa17_14_f_u_arrmul24_fa16_14_y4;
  wire f_u_arrmul24_fa17_14_y2;
  wire f_u_arrmul24_fa17_14_y3;
  wire f_u_arrmul24_fa17_14_y4;
  wire f_u_arrmul24_and18_14_a_18;
  wire f_u_arrmul24_and18_14_b_14;
  wire f_u_arrmul24_and18_14_y0;
  wire f_u_arrmul24_fa18_14_f_u_arrmul24_and18_14_y0;
  wire f_u_arrmul24_fa18_14_f_u_arrmul24_fa19_13_y2;
  wire f_u_arrmul24_fa18_14_y0;
  wire f_u_arrmul24_fa18_14_y1;
  wire f_u_arrmul24_fa18_14_f_u_arrmul24_fa17_14_y4;
  wire f_u_arrmul24_fa18_14_y2;
  wire f_u_arrmul24_fa18_14_y3;
  wire f_u_arrmul24_fa18_14_y4;
  wire f_u_arrmul24_and19_14_a_19;
  wire f_u_arrmul24_and19_14_b_14;
  wire f_u_arrmul24_and19_14_y0;
  wire f_u_arrmul24_fa19_14_f_u_arrmul24_and19_14_y0;
  wire f_u_arrmul24_fa19_14_f_u_arrmul24_fa20_13_y2;
  wire f_u_arrmul24_fa19_14_y0;
  wire f_u_arrmul24_fa19_14_y1;
  wire f_u_arrmul24_fa19_14_f_u_arrmul24_fa18_14_y4;
  wire f_u_arrmul24_fa19_14_y2;
  wire f_u_arrmul24_fa19_14_y3;
  wire f_u_arrmul24_fa19_14_y4;
  wire f_u_arrmul24_and20_14_a_20;
  wire f_u_arrmul24_and20_14_b_14;
  wire f_u_arrmul24_and20_14_y0;
  wire f_u_arrmul24_fa20_14_f_u_arrmul24_and20_14_y0;
  wire f_u_arrmul24_fa20_14_f_u_arrmul24_fa21_13_y2;
  wire f_u_arrmul24_fa20_14_y0;
  wire f_u_arrmul24_fa20_14_y1;
  wire f_u_arrmul24_fa20_14_f_u_arrmul24_fa19_14_y4;
  wire f_u_arrmul24_fa20_14_y2;
  wire f_u_arrmul24_fa20_14_y3;
  wire f_u_arrmul24_fa20_14_y4;
  wire f_u_arrmul24_and21_14_a_21;
  wire f_u_arrmul24_and21_14_b_14;
  wire f_u_arrmul24_and21_14_y0;
  wire f_u_arrmul24_fa21_14_f_u_arrmul24_and21_14_y0;
  wire f_u_arrmul24_fa21_14_f_u_arrmul24_fa22_13_y2;
  wire f_u_arrmul24_fa21_14_y0;
  wire f_u_arrmul24_fa21_14_y1;
  wire f_u_arrmul24_fa21_14_f_u_arrmul24_fa20_14_y4;
  wire f_u_arrmul24_fa21_14_y2;
  wire f_u_arrmul24_fa21_14_y3;
  wire f_u_arrmul24_fa21_14_y4;
  wire f_u_arrmul24_and22_14_a_22;
  wire f_u_arrmul24_and22_14_b_14;
  wire f_u_arrmul24_and22_14_y0;
  wire f_u_arrmul24_fa22_14_f_u_arrmul24_and22_14_y0;
  wire f_u_arrmul24_fa22_14_f_u_arrmul24_fa23_13_y2;
  wire f_u_arrmul24_fa22_14_y0;
  wire f_u_arrmul24_fa22_14_y1;
  wire f_u_arrmul24_fa22_14_f_u_arrmul24_fa21_14_y4;
  wire f_u_arrmul24_fa22_14_y2;
  wire f_u_arrmul24_fa22_14_y3;
  wire f_u_arrmul24_fa22_14_y4;
  wire f_u_arrmul24_and23_14_a_23;
  wire f_u_arrmul24_and23_14_b_14;
  wire f_u_arrmul24_and23_14_y0;
  wire f_u_arrmul24_fa23_14_f_u_arrmul24_and23_14_y0;
  wire f_u_arrmul24_fa23_14_f_u_arrmul24_fa23_13_y4;
  wire f_u_arrmul24_fa23_14_y0;
  wire f_u_arrmul24_fa23_14_y1;
  wire f_u_arrmul24_fa23_14_f_u_arrmul24_fa22_14_y4;
  wire f_u_arrmul24_fa23_14_y2;
  wire f_u_arrmul24_fa23_14_y3;
  wire f_u_arrmul24_fa23_14_y4;
  wire f_u_arrmul24_and0_15_a_0;
  wire f_u_arrmul24_and0_15_b_15;
  wire f_u_arrmul24_and0_15_y0;
  wire f_u_arrmul24_ha0_15_f_u_arrmul24_and0_15_y0;
  wire f_u_arrmul24_ha0_15_f_u_arrmul24_fa1_14_y2;
  wire f_u_arrmul24_ha0_15_y0;
  wire f_u_arrmul24_ha0_15_y1;
  wire f_u_arrmul24_and1_15_a_1;
  wire f_u_arrmul24_and1_15_b_15;
  wire f_u_arrmul24_and1_15_y0;
  wire f_u_arrmul24_fa1_15_f_u_arrmul24_and1_15_y0;
  wire f_u_arrmul24_fa1_15_f_u_arrmul24_fa2_14_y2;
  wire f_u_arrmul24_fa1_15_y0;
  wire f_u_arrmul24_fa1_15_y1;
  wire f_u_arrmul24_fa1_15_f_u_arrmul24_ha0_15_y1;
  wire f_u_arrmul24_fa1_15_y2;
  wire f_u_arrmul24_fa1_15_y3;
  wire f_u_arrmul24_fa1_15_y4;
  wire f_u_arrmul24_and2_15_a_2;
  wire f_u_arrmul24_and2_15_b_15;
  wire f_u_arrmul24_and2_15_y0;
  wire f_u_arrmul24_fa2_15_f_u_arrmul24_and2_15_y0;
  wire f_u_arrmul24_fa2_15_f_u_arrmul24_fa3_14_y2;
  wire f_u_arrmul24_fa2_15_y0;
  wire f_u_arrmul24_fa2_15_y1;
  wire f_u_arrmul24_fa2_15_f_u_arrmul24_fa1_15_y4;
  wire f_u_arrmul24_fa2_15_y2;
  wire f_u_arrmul24_fa2_15_y3;
  wire f_u_arrmul24_fa2_15_y4;
  wire f_u_arrmul24_and3_15_a_3;
  wire f_u_arrmul24_and3_15_b_15;
  wire f_u_arrmul24_and3_15_y0;
  wire f_u_arrmul24_fa3_15_f_u_arrmul24_and3_15_y0;
  wire f_u_arrmul24_fa3_15_f_u_arrmul24_fa4_14_y2;
  wire f_u_arrmul24_fa3_15_y0;
  wire f_u_arrmul24_fa3_15_y1;
  wire f_u_arrmul24_fa3_15_f_u_arrmul24_fa2_15_y4;
  wire f_u_arrmul24_fa3_15_y2;
  wire f_u_arrmul24_fa3_15_y3;
  wire f_u_arrmul24_fa3_15_y4;
  wire f_u_arrmul24_and4_15_a_4;
  wire f_u_arrmul24_and4_15_b_15;
  wire f_u_arrmul24_and4_15_y0;
  wire f_u_arrmul24_fa4_15_f_u_arrmul24_and4_15_y0;
  wire f_u_arrmul24_fa4_15_f_u_arrmul24_fa5_14_y2;
  wire f_u_arrmul24_fa4_15_y0;
  wire f_u_arrmul24_fa4_15_y1;
  wire f_u_arrmul24_fa4_15_f_u_arrmul24_fa3_15_y4;
  wire f_u_arrmul24_fa4_15_y2;
  wire f_u_arrmul24_fa4_15_y3;
  wire f_u_arrmul24_fa4_15_y4;
  wire f_u_arrmul24_and5_15_a_5;
  wire f_u_arrmul24_and5_15_b_15;
  wire f_u_arrmul24_and5_15_y0;
  wire f_u_arrmul24_fa5_15_f_u_arrmul24_and5_15_y0;
  wire f_u_arrmul24_fa5_15_f_u_arrmul24_fa6_14_y2;
  wire f_u_arrmul24_fa5_15_y0;
  wire f_u_arrmul24_fa5_15_y1;
  wire f_u_arrmul24_fa5_15_f_u_arrmul24_fa4_15_y4;
  wire f_u_arrmul24_fa5_15_y2;
  wire f_u_arrmul24_fa5_15_y3;
  wire f_u_arrmul24_fa5_15_y4;
  wire f_u_arrmul24_and6_15_a_6;
  wire f_u_arrmul24_and6_15_b_15;
  wire f_u_arrmul24_and6_15_y0;
  wire f_u_arrmul24_fa6_15_f_u_arrmul24_and6_15_y0;
  wire f_u_arrmul24_fa6_15_f_u_arrmul24_fa7_14_y2;
  wire f_u_arrmul24_fa6_15_y0;
  wire f_u_arrmul24_fa6_15_y1;
  wire f_u_arrmul24_fa6_15_f_u_arrmul24_fa5_15_y4;
  wire f_u_arrmul24_fa6_15_y2;
  wire f_u_arrmul24_fa6_15_y3;
  wire f_u_arrmul24_fa6_15_y4;
  wire f_u_arrmul24_and7_15_a_7;
  wire f_u_arrmul24_and7_15_b_15;
  wire f_u_arrmul24_and7_15_y0;
  wire f_u_arrmul24_fa7_15_f_u_arrmul24_and7_15_y0;
  wire f_u_arrmul24_fa7_15_f_u_arrmul24_fa8_14_y2;
  wire f_u_arrmul24_fa7_15_y0;
  wire f_u_arrmul24_fa7_15_y1;
  wire f_u_arrmul24_fa7_15_f_u_arrmul24_fa6_15_y4;
  wire f_u_arrmul24_fa7_15_y2;
  wire f_u_arrmul24_fa7_15_y3;
  wire f_u_arrmul24_fa7_15_y4;
  wire f_u_arrmul24_and8_15_a_8;
  wire f_u_arrmul24_and8_15_b_15;
  wire f_u_arrmul24_and8_15_y0;
  wire f_u_arrmul24_fa8_15_f_u_arrmul24_and8_15_y0;
  wire f_u_arrmul24_fa8_15_f_u_arrmul24_fa9_14_y2;
  wire f_u_arrmul24_fa8_15_y0;
  wire f_u_arrmul24_fa8_15_y1;
  wire f_u_arrmul24_fa8_15_f_u_arrmul24_fa7_15_y4;
  wire f_u_arrmul24_fa8_15_y2;
  wire f_u_arrmul24_fa8_15_y3;
  wire f_u_arrmul24_fa8_15_y4;
  wire f_u_arrmul24_and9_15_a_9;
  wire f_u_arrmul24_and9_15_b_15;
  wire f_u_arrmul24_and9_15_y0;
  wire f_u_arrmul24_fa9_15_f_u_arrmul24_and9_15_y0;
  wire f_u_arrmul24_fa9_15_f_u_arrmul24_fa10_14_y2;
  wire f_u_arrmul24_fa9_15_y0;
  wire f_u_arrmul24_fa9_15_y1;
  wire f_u_arrmul24_fa9_15_f_u_arrmul24_fa8_15_y4;
  wire f_u_arrmul24_fa9_15_y2;
  wire f_u_arrmul24_fa9_15_y3;
  wire f_u_arrmul24_fa9_15_y4;
  wire f_u_arrmul24_and10_15_a_10;
  wire f_u_arrmul24_and10_15_b_15;
  wire f_u_arrmul24_and10_15_y0;
  wire f_u_arrmul24_fa10_15_f_u_arrmul24_and10_15_y0;
  wire f_u_arrmul24_fa10_15_f_u_arrmul24_fa11_14_y2;
  wire f_u_arrmul24_fa10_15_y0;
  wire f_u_arrmul24_fa10_15_y1;
  wire f_u_arrmul24_fa10_15_f_u_arrmul24_fa9_15_y4;
  wire f_u_arrmul24_fa10_15_y2;
  wire f_u_arrmul24_fa10_15_y3;
  wire f_u_arrmul24_fa10_15_y4;
  wire f_u_arrmul24_and11_15_a_11;
  wire f_u_arrmul24_and11_15_b_15;
  wire f_u_arrmul24_and11_15_y0;
  wire f_u_arrmul24_fa11_15_f_u_arrmul24_and11_15_y0;
  wire f_u_arrmul24_fa11_15_f_u_arrmul24_fa12_14_y2;
  wire f_u_arrmul24_fa11_15_y0;
  wire f_u_arrmul24_fa11_15_y1;
  wire f_u_arrmul24_fa11_15_f_u_arrmul24_fa10_15_y4;
  wire f_u_arrmul24_fa11_15_y2;
  wire f_u_arrmul24_fa11_15_y3;
  wire f_u_arrmul24_fa11_15_y4;
  wire f_u_arrmul24_and12_15_a_12;
  wire f_u_arrmul24_and12_15_b_15;
  wire f_u_arrmul24_and12_15_y0;
  wire f_u_arrmul24_fa12_15_f_u_arrmul24_and12_15_y0;
  wire f_u_arrmul24_fa12_15_f_u_arrmul24_fa13_14_y2;
  wire f_u_arrmul24_fa12_15_y0;
  wire f_u_arrmul24_fa12_15_y1;
  wire f_u_arrmul24_fa12_15_f_u_arrmul24_fa11_15_y4;
  wire f_u_arrmul24_fa12_15_y2;
  wire f_u_arrmul24_fa12_15_y3;
  wire f_u_arrmul24_fa12_15_y4;
  wire f_u_arrmul24_and13_15_a_13;
  wire f_u_arrmul24_and13_15_b_15;
  wire f_u_arrmul24_and13_15_y0;
  wire f_u_arrmul24_fa13_15_f_u_arrmul24_and13_15_y0;
  wire f_u_arrmul24_fa13_15_f_u_arrmul24_fa14_14_y2;
  wire f_u_arrmul24_fa13_15_y0;
  wire f_u_arrmul24_fa13_15_y1;
  wire f_u_arrmul24_fa13_15_f_u_arrmul24_fa12_15_y4;
  wire f_u_arrmul24_fa13_15_y2;
  wire f_u_arrmul24_fa13_15_y3;
  wire f_u_arrmul24_fa13_15_y4;
  wire f_u_arrmul24_and14_15_a_14;
  wire f_u_arrmul24_and14_15_b_15;
  wire f_u_arrmul24_and14_15_y0;
  wire f_u_arrmul24_fa14_15_f_u_arrmul24_and14_15_y0;
  wire f_u_arrmul24_fa14_15_f_u_arrmul24_fa15_14_y2;
  wire f_u_arrmul24_fa14_15_y0;
  wire f_u_arrmul24_fa14_15_y1;
  wire f_u_arrmul24_fa14_15_f_u_arrmul24_fa13_15_y4;
  wire f_u_arrmul24_fa14_15_y2;
  wire f_u_arrmul24_fa14_15_y3;
  wire f_u_arrmul24_fa14_15_y4;
  wire f_u_arrmul24_and15_15_a_15;
  wire f_u_arrmul24_and15_15_b_15;
  wire f_u_arrmul24_and15_15_y0;
  wire f_u_arrmul24_fa15_15_f_u_arrmul24_and15_15_y0;
  wire f_u_arrmul24_fa15_15_f_u_arrmul24_fa16_14_y2;
  wire f_u_arrmul24_fa15_15_y0;
  wire f_u_arrmul24_fa15_15_y1;
  wire f_u_arrmul24_fa15_15_f_u_arrmul24_fa14_15_y4;
  wire f_u_arrmul24_fa15_15_y2;
  wire f_u_arrmul24_fa15_15_y3;
  wire f_u_arrmul24_fa15_15_y4;
  wire f_u_arrmul24_and16_15_a_16;
  wire f_u_arrmul24_and16_15_b_15;
  wire f_u_arrmul24_and16_15_y0;
  wire f_u_arrmul24_fa16_15_f_u_arrmul24_and16_15_y0;
  wire f_u_arrmul24_fa16_15_f_u_arrmul24_fa17_14_y2;
  wire f_u_arrmul24_fa16_15_y0;
  wire f_u_arrmul24_fa16_15_y1;
  wire f_u_arrmul24_fa16_15_f_u_arrmul24_fa15_15_y4;
  wire f_u_arrmul24_fa16_15_y2;
  wire f_u_arrmul24_fa16_15_y3;
  wire f_u_arrmul24_fa16_15_y4;
  wire f_u_arrmul24_and17_15_a_17;
  wire f_u_arrmul24_and17_15_b_15;
  wire f_u_arrmul24_and17_15_y0;
  wire f_u_arrmul24_fa17_15_f_u_arrmul24_and17_15_y0;
  wire f_u_arrmul24_fa17_15_f_u_arrmul24_fa18_14_y2;
  wire f_u_arrmul24_fa17_15_y0;
  wire f_u_arrmul24_fa17_15_y1;
  wire f_u_arrmul24_fa17_15_f_u_arrmul24_fa16_15_y4;
  wire f_u_arrmul24_fa17_15_y2;
  wire f_u_arrmul24_fa17_15_y3;
  wire f_u_arrmul24_fa17_15_y4;
  wire f_u_arrmul24_and18_15_a_18;
  wire f_u_arrmul24_and18_15_b_15;
  wire f_u_arrmul24_and18_15_y0;
  wire f_u_arrmul24_fa18_15_f_u_arrmul24_and18_15_y0;
  wire f_u_arrmul24_fa18_15_f_u_arrmul24_fa19_14_y2;
  wire f_u_arrmul24_fa18_15_y0;
  wire f_u_arrmul24_fa18_15_y1;
  wire f_u_arrmul24_fa18_15_f_u_arrmul24_fa17_15_y4;
  wire f_u_arrmul24_fa18_15_y2;
  wire f_u_arrmul24_fa18_15_y3;
  wire f_u_arrmul24_fa18_15_y4;
  wire f_u_arrmul24_and19_15_a_19;
  wire f_u_arrmul24_and19_15_b_15;
  wire f_u_arrmul24_and19_15_y0;
  wire f_u_arrmul24_fa19_15_f_u_arrmul24_and19_15_y0;
  wire f_u_arrmul24_fa19_15_f_u_arrmul24_fa20_14_y2;
  wire f_u_arrmul24_fa19_15_y0;
  wire f_u_arrmul24_fa19_15_y1;
  wire f_u_arrmul24_fa19_15_f_u_arrmul24_fa18_15_y4;
  wire f_u_arrmul24_fa19_15_y2;
  wire f_u_arrmul24_fa19_15_y3;
  wire f_u_arrmul24_fa19_15_y4;
  wire f_u_arrmul24_and20_15_a_20;
  wire f_u_arrmul24_and20_15_b_15;
  wire f_u_arrmul24_and20_15_y0;
  wire f_u_arrmul24_fa20_15_f_u_arrmul24_and20_15_y0;
  wire f_u_arrmul24_fa20_15_f_u_arrmul24_fa21_14_y2;
  wire f_u_arrmul24_fa20_15_y0;
  wire f_u_arrmul24_fa20_15_y1;
  wire f_u_arrmul24_fa20_15_f_u_arrmul24_fa19_15_y4;
  wire f_u_arrmul24_fa20_15_y2;
  wire f_u_arrmul24_fa20_15_y3;
  wire f_u_arrmul24_fa20_15_y4;
  wire f_u_arrmul24_and21_15_a_21;
  wire f_u_arrmul24_and21_15_b_15;
  wire f_u_arrmul24_and21_15_y0;
  wire f_u_arrmul24_fa21_15_f_u_arrmul24_and21_15_y0;
  wire f_u_arrmul24_fa21_15_f_u_arrmul24_fa22_14_y2;
  wire f_u_arrmul24_fa21_15_y0;
  wire f_u_arrmul24_fa21_15_y1;
  wire f_u_arrmul24_fa21_15_f_u_arrmul24_fa20_15_y4;
  wire f_u_arrmul24_fa21_15_y2;
  wire f_u_arrmul24_fa21_15_y3;
  wire f_u_arrmul24_fa21_15_y4;
  wire f_u_arrmul24_and22_15_a_22;
  wire f_u_arrmul24_and22_15_b_15;
  wire f_u_arrmul24_and22_15_y0;
  wire f_u_arrmul24_fa22_15_f_u_arrmul24_and22_15_y0;
  wire f_u_arrmul24_fa22_15_f_u_arrmul24_fa23_14_y2;
  wire f_u_arrmul24_fa22_15_y0;
  wire f_u_arrmul24_fa22_15_y1;
  wire f_u_arrmul24_fa22_15_f_u_arrmul24_fa21_15_y4;
  wire f_u_arrmul24_fa22_15_y2;
  wire f_u_arrmul24_fa22_15_y3;
  wire f_u_arrmul24_fa22_15_y4;
  wire f_u_arrmul24_and23_15_a_23;
  wire f_u_arrmul24_and23_15_b_15;
  wire f_u_arrmul24_and23_15_y0;
  wire f_u_arrmul24_fa23_15_f_u_arrmul24_and23_15_y0;
  wire f_u_arrmul24_fa23_15_f_u_arrmul24_fa23_14_y4;
  wire f_u_arrmul24_fa23_15_y0;
  wire f_u_arrmul24_fa23_15_y1;
  wire f_u_arrmul24_fa23_15_f_u_arrmul24_fa22_15_y4;
  wire f_u_arrmul24_fa23_15_y2;
  wire f_u_arrmul24_fa23_15_y3;
  wire f_u_arrmul24_fa23_15_y4;
  wire f_u_arrmul24_and0_16_a_0;
  wire f_u_arrmul24_and0_16_b_16;
  wire f_u_arrmul24_and0_16_y0;
  wire f_u_arrmul24_ha0_16_f_u_arrmul24_and0_16_y0;
  wire f_u_arrmul24_ha0_16_f_u_arrmul24_fa1_15_y2;
  wire f_u_arrmul24_ha0_16_y0;
  wire f_u_arrmul24_ha0_16_y1;
  wire f_u_arrmul24_and1_16_a_1;
  wire f_u_arrmul24_and1_16_b_16;
  wire f_u_arrmul24_and1_16_y0;
  wire f_u_arrmul24_fa1_16_f_u_arrmul24_and1_16_y0;
  wire f_u_arrmul24_fa1_16_f_u_arrmul24_fa2_15_y2;
  wire f_u_arrmul24_fa1_16_y0;
  wire f_u_arrmul24_fa1_16_y1;
  wire f_u_arrmul24_fa1_16_f_u_arrmul24_ha0_16_y1;
  wire f_u_arrmul24_fa1_16_y2;
  wire f_u_arrmul24_fa1_16_y3;
  wire f_u_arrmul24_fa1_16_y4;
  wire f_u_arrmul24_and2_16_a_2;
  wire f_u_arrmul24_and2_16_b_16;
  wire f_u_arrmul24_and2_16_y0;
  wire f_u_arrmul24_fa2_16_f_u_arrmul24_and2_16_y0;
  wire f_u_arrmul24_fa2_16_f_u_arrmul24_fa3_15_y2;
  wire f_u_arrmul24_fa2_16_y0;
  wire f_u_arrmul24_fa2_16_y1;
  wire f_u_arrmul24_fa2_16_f_u_arrmul24_fa1_16_y4;
  wire f_u_arrmul24_fa2_16_y2;
  wire f_u_arrmul24_fa2_16_y3;
  wire f_u_arrmul24_fa2_16_y4;
  wire f_u_arrmul24_and3_16_a_3;
  wire f_u_arrmul24_and3_16_b_16;
  wire f_u_arrmul24_and3_16_y0;
  wire f_u_arrmul24_fa3_16_f_u_arrmul24_and3_16_y0;
  wire f_u_arrmul24_fa3_16_f_u_arrmul24_fa4_15_y2;
  wire f_u_arrmul24_fa3_16_y0;
  wire f_u_arrmul24_fa3_16_y1;
  wire f_u_arrmul24_fa3_16_f_u_arrmul24_fa2_16_y4;
  wire f_u_arrmul24_fa3_16_y2;
  wire f_u_arrmul24_fa3_16_y3;
  wire f_u_arrmul24_fa3_16_y4;
  wire f_u_arrmul24_and4_16_a_4;
  wire f_u_arrmul24_and4_16_b_16;
  wire f_u_arrmul24_and4_16_y0;
  wire f_u_arrmul24_fa4_16_f_u_arrmul24_and4_16_y0;
  wire f_u_arrmul24_fa4_16_f_u_arrmul24_fa5_15_y2;
  wire f_u_arrmul24_fa4_16_y0;
  wire f_u_arrmul24_fa4_16_y1;
  wire f_u_arrmul24_fa4_16_f_u_arrmul24_fa3_16_y4;
  wire f_u_arrmul24_fa4_16_y2;
  wire f_u_arrmul24_fa4_16_y3;
  wire f_u_arrmul24_fa4_16_y4;
  wire f_u_arrmul24_and5_16_a_5;
  wire f_u_arrmul24_and5_16_b_16;
  wire f_u_arrmul24_and5_16_y0;
  wire f_u_arrmul24_fa5_16_f_u_arrmul24_and5_16_y0;
  wire f_u_arrmul24_fa5_16_f_u_arrmul24_fa6_15_y2;
  wire f_u_arrmul24_fa5_16_y0;
  wire f_u_arrmul24_fa5_16_y1;
  wire f_u_arrmul24_fa5_16_f_u_arrmul24_fa4_16_y4;
  wire f_u_arrmul24_fa5_16_y2;
  wire f_u_arrmul24_fa5_16_y3;
  wire f_u_arrmul24_fa5_16_y4;
  wire f_u_arrmul24_and6_16_a_6;
  wire f_u_arrmul24_and6_16_b_16;
  wire f_u_arrmul24_and6_16_y0;
  wire f_u_arrmul24_fa6_16_f_u_arrmul24_and6_16_y0;
  wire f_u_arrmul24_fa6_16_f_u_arrmul24_fa7_15_y2;
  wire f_u_arrmul24_fa6_16_y0;
  wire f_u_arrmul24_fa6_16_y1;
  wire f_u_arrmul24_fa6_16_f_u_arrmul24_fa5_16_y4;
  wire f_u_arrmul24_fa6_16_y2;
  wire f_u_arrmul24_fa6_16_y3;
  wire f_u_arrmul24_fa6_16_y4;
  wire f_u_arrmul24_and7_16_a_7;
  wire f_u_arrmul24_and7_16_b_16;
  wire f_u_arrmul24_and7_16_y0;
  wire f_u_arrmul24_fa7_16_f_u_arrmul24_and7_16_y0;
  wire f_u_arrmul24_fa7_16_f_u_arrmul24_fa8_15_y2;
  wire f_u_arrmul24_fa7_16_y0;
  wire f_u_arrmul24_fa7_16_y1;
  wire f_u_arrmul24_fa7_16_f_u_arrmul24_fa6_16_y4;
  wire f_u_arrmul24_fa7_16_y2;
  wire f_u_arrmul24_fa7_16_y3;
  wire f_u_arrmul24_fa7_16_y4;
  wire f_u_arrmul24_and8_16_a_8;
  wire f_u_arrmul24_and8_16_b_16;
  wire f_u_arrmul24_and8_16_y0;
  wire f_u_arrmul24_fa8_16_f_u_arrmul24_and8_16_y0;
  wire f_u_arrmul24_fa8_16_f_u_arrmul24_fa9_15_y2;
  wire f_u_arrmul24_fa8_16_y0;
  wire f_u_arrmul24_fa8_16_y1;
  wire f_u_arrmul24_fa8_16_f_u_arrmul24_fa7_16_y4;
  wire f_u_arrmul24_fa8_16_y2;
  wire f_u_arrmul24_fa8_16_y3;
  wire f_u_arrmul24_fa8_16_y4;
  wire f_u_arrmul24_and9_16_a_9;
  wire f_u_arrmul24_and9_16_b_16;
  wire f_u_arrmul24_and9_16_y0;
  wire f_u_arrmul24_fa9_16_f_u_arrmul24_and9_16_y0;
  wire f_u_arrmul24_fa9_16_f_u_arrmul24_fa10_15_y2;
  wire f_u_arrmul24_fa9_16_y0;
  wire f_u_arrmul24_fa9_16_y1;
  wire f_u_arrmul24_fa9_16_f_u_arrmul24_fa8_16_y4;
  wire f_u_arrmul24_fa9_16_y2;
  wire f_u_arrmul24_fa9_16_y3;
  wire f_u_arrmul24_fa9_16_y4;
  wire f_u_arrmul24_and10_16_a_10;
  wire f_u_arrmul24_and10_16_b_16;
  wire f_u_arrmul24_and10_16_y0;
  wire f_u_arrmul24_fa10_16_f_u_arrmul24_and10_16_y0;
  wire f_u_arrmul24_fa10_16_f_u_arrmul24_fa11_15_y2;
  wire f_u_arrmul24_fa10_16_y0;
  wire f_u_arrmul24_fa10_16_y1;
  wire f_u_arrmul24_fa10_16_f_u_arrmul24_fa9_16_y4;
  wire f_u_arrmul24_fa10_16_y2;
  wire f_u_arrmul24_fa10_16_y3;
  wire f_u_arrmul24_fa10_16_y4;
  wire f_u_arrmul24_and11_16_a_11;
  wire f_u_arrmul24_and11_16_b_16;
  wire f_u_arrmul24_and11_16_y0;
  wire f_u_arrmul24_fa11_16_f_u_arrmul24_and11_16_y0;
  wire f_u_arrmul24_fa11_16_f_u_arrmul24_fa12_15_y2;
  wire f_u_arrmul24_fa11_16_y0;
  wire f_u_arrmul24_fa11_16_y1;
  wire f_u_arrmul24_fa11_16_f_u_arrmul24_fa10_16_y4;
  wire f_u_arrmul24_fa11_16_y2;
  wire f_u_arrmul24_fa11_16_y3;
  wire f_u_arrmul24_fa11_16_y4;
  wire f_u_arrmul24_and12_16_a_12;
  wire f_u_arrmul24_and12_16_b_16;
  wire f_u_arrmul24_and12_16_y0;
  wire f_u_arrmul24_fa12_16_f_u_arrmul24_and12_16_y0;
  wire f_u_arrmul24_fa12_16_f_u_arrmul24_fa13_15_y2;
  wire f_u_arrmul24_fa12_16_y0;
  wire f_u_arrmul24_fa12_16_y1;
  wire f_u_arrmul24_fa12_16_f_u_arrmul24_fa11_16_y4;
  wire f_u_arrmul24_fa12_16_y2;
  wire f_u_arrmul24_fa12_16_y3;
  wire f_u_arrmul24_fa12_16_y4;
  wire f_u_arrmul24_and13_16_a_13;
  wire f_u_arrmul24_and13_16_b_16;
  wire f_u_arrmul24_and13_16_y0;
  wire f_u_arrmul24_fa13_16_f_u_arrmul24_and13_16_y0;
  wire f_u_arrmul24_fa13_16_f_u_arrmul24_fa14_15_y2;
  wire f_u_arrmul24_fa13_16_y0;
  wire f_u_arrmul24_fa13_16_y1;
  wire f_u_arrmul24_fa13_16_f_u_arrmul24_fa12_16_y4;
  wire f_u_arrmul24_fa13_16_y2;
  wire f_u_arrmul24_fa13_16_y3;
  wire f_u_arrmul24_fa13_16_y4;
  wire f_u_arrmul24_and14_16_a_14;
  wire f_u_arrmul24_and14_16_b_16;
  wire f_u_arrmul24_and14_16_y0;
  wire f_u_arrmul24_fa14_16_f_u_arrmul24_and14_16_y0;
  wire f_u_arrmul24_fa14_16_f_u_arrmul24_fa15_15_y2;
  wire f_u_arrmul24_fa14_16_y0;
  wire f_u_arrmul24_fa14_16_y1;
  wire f_u_arrmul24_fa14_16_f_u_arrmul24_fa13_16_y4;
  wire f_u_arrmul24_fa14_16_y2;
  wire f_u_arrmul24_fa14_16_y3;
  wire f_u_arrmul24_fa14_16_y4;
  wire f_u_arrmul24_and15_16_a_15;
  wire f_u_arrmul24_and15_16_b_16;
  wire f_u_arrmul24_and15_16_y0;
  wire f_u_arrmul24_fa15_16_f_u_arrmul24_and15_16_y0;
  wire f_u_arrmul24_fa15_16_f_u_arrmul24_fa16_15_y2;
  wire f_u_arrmul24_fa15_16_y0;
  wire f_u_arrmul24_fa15_16_y1;
  wire f_u_arrmul24_fa15_16_f_u_arrmul24_fa14_16_y4;
  wire f_u_arrmul24_fa15_16_y2;
  wire f_u_arrmul24_fa15_16_y3;
  wire f_u_arrmul24_fa15_16_y4;
  wire f_u_arrmul24_and16_16_a_16;
  wire f_u_arrmul24_and16_16_b_16;
  wire f_u_arrmul24_and16_16_y0;
  wire f_u_arrmul24_fa16_16_f_u_arrmul24_and16_16_y0;
  wire f_u_arrmul24_fa16_16_f_u_arrmul24_fa17_15_y2;
  wire f_u_arrmul24_fa16_16_y0;
  wire f_u_arrmul24_fa16_16_y1;
  wire f_u_arrmul24_fa16_16_f_u_arrmul24_fa15_16_y4;
  wire f_u_arrmul24_fa16_16_y2;
  wire f_u_arrmul24_fa16_16_y3;
  wire f_u_arrmul24_fa16_16_y4;
  wire f_u_arrmul24_and17_16_a_17;
  wire f_u_arrmul24_and17_16_b_16;
  wire f_u_arrmul24_and17_16_y0;
  wire f_u_arrmul24_fa17_16_f_u_arrmul24_and17_16_y0;
  wire f_u_arrmul24_fa17_16_f_u_arrmul24_fa18_15_y2;
  wire f_u_arrmul24_fa17_16_y0;
  wire f_u_arrmul24_fa17_16_y1;
  wire f_u_arrmul24_fa17_16_f_u_arrmul24_fa16_16_y4;
  wire f_u_arrmul24_fa17_16_y2;
  wire f_u_arrmul24_fa17_16_y3;
  wire f_u_arrmul24_fa17_16_y4;
  wire f_u_arrmul24_and18_16_a_18;
  wire f_u_arrmul24_and18_16_b_16;
  wire f_u_arrmul24_and18_16_y0;
  wire f_u_arrmul24_fa18_16_f_u_arrmul24_and18_16_y0;
  wire f_u_arrmul24_fa18_16_f_u_arrmul24_fa19_15_y2;
  wire f_u_arrmul24_fa18_16_y0;
  wire f_u_arrmul24_fa18_16_y1;
  wire f_u_arrmul24_fa18_16_f_u_arrmul24_fa17_16_y4;
  wire f_u_arrmul24_fa18_16_y2;
  wire f_u_arrmul24_fa18_16_y3;
  wire f_u_arrmul24_fa18_16_y4;
  wire f_u_arrmul24_and19_16_a_19;
  wire f_u_arrmul24_and19_16_b_16;
  wire f_u_arrmul24_and19_16_y0;
  wire f_u_arrmul24_fa19_16_f_u_arrmul24_and19_16_y0;
  wire f_u_arrmul24_fa19_16_f_u_arrmul24_fa20_15_y2;
  wire f_u_arrmul24_fa19_16_y0;
  wire f_u_arrmul24_fa19_16_y1;
  wire f_u_arrmul24_fa19_16_f_u_arrmul24_fa18_16_y4;
  wire f_u_arrmul24_fa19_16_y2;
  wire f_u_arrmul24_fa19_16_y3;
  wire f_u_arrmul24_fa19_16_y4;
  wire f_u_arrmul24_and20_16_a_20;
  wire f_u_arrmul24_and20_16_b_16;
  wire f_u_arrmul24_and20_16_y0;
  wire f_u_arrmul24_fa20_16_f_u_arrmul24_and20_16_y0;
  wire f_u_arrmul24_fa20_16_f_u_arrmul24_fa21_15_y2;
  wire f_u_arrmul24_fa20_16_y0;
  wire f_u_arrmul24_fa20_16_y1;
  wire f_u_arrmul24_fa20_16_f_u_arrmul24_fa19_16_y4;
  wire f_u_arrmul24_fa20_16_y2;
  wire f_u_arrmul24_fa20_16_y3;
  wire f_u_arrmul24_fa20_16_y4;
  wire f_u_arrmul24_and21_16_a_21;
  wire f_u_arrmul24_and21_16_b_16;
  wire f_u_arrmul24_and21_16_y0;
  wire f_u_arrmul24_fa21_16_f_u_arrmul24_and21_16_y0;
  wire f_u_arrmul24_fa21_16_f_u_arrmul24_fa22_15_y2;
  wire f_u_arrmul24_fa21_16_y0;
  wire f_u_arrmul24_fa21_16_y1;
  wire f_u_arrmul24_fa21_16_f_u_arrmul24_fa20_16_y4;
  wire f_u_arrmul24_fa21_16_y2;
  wire f_u_arrmul24_fa21_16_y3;
  wire f_u_arrmul24_fa21_16_y4;
  wire f_u_arrmul24_and22_16_a_22;
  wire f_u_arrmul24_and22_16_b_16;
  wire f_u_arrmul24_and22_16_y0;
  wire f_u_arrmul24_fa22_16_f_u_arrmul24_and22_16_y0;
  wire f_u_arrmul24_fa22_16_f_u_arrmul24_fa23_15_y2;
  wire f_u_arrmul24_fa22_16_y0;
  wire f_u_arrmul24_fa22_16_y1;
  wire f_u_arrmul24_fa22_16_f_u_arrmul24_fa21_16_y4;
  wire f_u_arrmul24_fa22_16_y2;
  wire f_u_arrmul24_fa22_16_y3;
  wire f_u_arrmul24_fa22_16_y4;
  wire f_u_arrmul24_and23_16_a_23;
  wire f_u_arrmul24_and23_16_b_16;
  wire f_u_arrmul24_and23_16_y0;
  wire f_u_arrmul24_fa23_16_f_u_arrmul24_and23_16_y0;
  wire f_u_arrmul24_fa23_16_f_u_arrmul24_fa23_15_y4;
  wire f_u_arrmul24_fa23_16_y0;
  wire f_u_arrmul24_fa23_16_y1;
  wire f_u_arrmul24_fa23_16_f_u_arrmul24_fa22_16_y4;
  wire f_u_arrmul24_fa23_16_y2;
  wire f_u_arrmul24_fa23_16_y3;
  wire f_u_arrmul24_fa23_16_y4;
  wire f_u_arrmul24_and0_17_a_0;
  wire f_u_arrmul24_and0_17_b_17;
  wire f_u_arrmul24_and0_17_y0;
  wire f_u_arrmul24_ha0_17_f_u_arrmul24_and0_17_y0;
  wire f_u_arrmul24_ha0_17_f_u_arrmul24_fa1_16_y2;
  wire f_u_arrmul24_ha0_17_y0;
  wire f_u_arrmul24_ha0_17_y1;
  wire f_u_arrmul24_and1_17_a_1;
  wire f_u_arrmul24_and1_17_b_17;
  wire f_u_arrmul24_and1_17_y0;
  wire f_u_arrmul24_fa1_17_f_u_arrmul24_and1_17_y0;
  wire f_u_arrmul24_fa1_17_f_u_arrmul24_fa2_16_y2;
  wire f_u_arrmul24_fa1_17_y0;
  wire f_u_arrmul24_fa1_17_y1;
  wire f_u_arrmul24_fa1_17_f_u_arrmul24_ha0_17_y1;
  wire f_u_arrmul24_fa1_17_y2;
  wire f_u_arrmul24_fa1_17_y3;
  wire f_u_arrmul24_fa1_17_y4;
  wire f_u_arrmul24_and2_17_a_2;
  wire f_u_arrmul24_and2_17_b_17;
  wire f_u_arrmul24_and2_17_y0;
  wire f_u_arrmul24_fa2_17_f_u_arrmul24_and2_17_y0;
  wire f_u_arrmul24_fa2_17_f_u_arrmul24_fa3_16_y2;
  wire f_u_arrmul24_fa2_17_y0;
  wire f_u_arrmul24_fa2_17_y1;
  wire f_u_arrmul24_fa2_17_f_u_arrmul24_fa1_17_y4;
  wire f_u_arrmul24_fa2_17_y2;
  wire f_u_arrmul24_fa2_17_y3;
  wire f_u_arrmul24_fa2_17_y4;
  wire f_u_arrmul24_and3_17_a_3;
  wire f_u_arrmul24_and3_17_b_17;
  wire f_u_arrmul24_and3_17_y0;
  wire f_u_arrmul24_fa3_17_f_u_arrmul24_and3_17_y0;
  wire f_u_arrmul24_fa3_17_f_u_arrmul24_fa4_16_y2;
  wire f_u_arrmul24_fa3_17_y0;
  wire f_u_arrmul24_fa3_17_y1;
  wire f_u_arrmul24_fa3_17_f_u_arrmul24_fa2_17_y4;
  wire f_u_arrmul24_fa3_17_y2;
  wire f_u_arrmul24_fa3_17_y3;
  wire f_u_arrmul24_fa3_17_y4;
  wire f_u_arrmul24_and4_17_a_4;
  wire f_u_arrmul24_and4_17_b_17;
  wire f_u_arrmul24_and4_17_y0;
  wire f_u_arrmul24_fa4_17_f_u_arrmul24_and4_17_y0;
  wire f_u_arrmul24_fa4_17_f_u_arrmul24_fa5_16_y2;
  wire f_u_arrmul24_fa4_17_y0;
  wire f_u_arrmul24_fa4_17_y1;
  wire f_u_arrmul24_fa4_17_f_u_arrmul24_fa3_17_y4;
  wire f_u_arrmul24_fa4_17_y2;
  wire f_u_arrmul24_fa4_17_y3;
  wire f_u_arrmul24_fa4_17_y4;
  wire f_u_arrmul24_and5_17_a_5;
  wire f_u_arrmul24_and5_17_b_17;
  wire f_u_arrmul24_and5_17_y0;
  wire f_u_arrmul24_fa5_17_f_u_arrmul24_and5_17_y0;
  wire f_u_arrmul24_fa5_17_f_u_arrmul24_fa6_16_y2;
  wire f_u_arrmul24_fa5_17_y0;
  wire f_u_arrmul24_fa5_17_y1;
  wire f_u_arrmul24_fa5_17_f_u_arrmul24_fa4_17_y4;
  wire f_u_arrmul24_fa5_17_y2;
  wire f_u_arrmul24_fa5_17_y3;
  wire f_u_arrmul24_fa5_17_y4;
  wire f_u_arrmul24_and6_17_a_6;
  wire f_u_arrmul24_and6_17_b_17;
  wire f_u_arrmul24_and6_17_y0;
  wire f_u_arrmul24_fa6_17_f_u_arrmul24_and6_17_y0;
  wire f_u_arrmul24_fa6_17_f_u_arrmul24_fa7_16_y2;
  wire f_u_arrmul24_fa6_17_y0;
  wire f_u_arrmul24_fa6_17_y1;
  wire f_u_arrmul24_fa6_17_f_u_arrmul24_fa5_17_y4;
  wire f_u_arrmul24_fa6_17_y2;
  wire f_u_arrmul24_fa6_17_y3;
  wire f_u_arrmul24_fa6_17_y4;
  wire f_u_arrmul24_and7_17_a_7;
  wire f_u_arrmul24_and7_17_b_17;
  wire f_u_arrmul24_and7_17_y0;
  wire f_u_arrmul24_fa7_17_f_u_arrmul24_and7_17_y0;
  wire f_u_arrmul24_fa7_17_f_u_arrmul24_fa8_16_y2;
  wire f_u_arrmul24_fa7_17_y0;
  wire f_u_arrmul24_fa7_17_y1;
  wire f_u_arrmul24_fa7_17_f_u_arrmul24_fa6_17_y4;
  wire f_u_arrmul24_fa7_17_y2;
  wire f_u_arrmul24_fa7_17_y3;
  wire f_u_arrmul24_fa7_17_y4;
  wire f_u_arrmul24_and8_17_a_8;
  wire f_u_arrmul24_and8_17_b_17;
  wire f_u_arrmul24_and8_17_y0;
  wire f_u_arrmul24_fa8_17_f_u_arrmul24_and8_17_y0;
  wire f_u_arrmul24_fa8_17_f_u_arrmul24_fa9_16_y2;
  wire f_u_arrmul24_fa8_17_y0;
  wire f_u_arrmul24_fa8_17_y1;
  wire f_u_arrmul24_fa8_17_f_u_arrmul24_fa7_17_y4;
  wire f_u_arrmul24_fa8_17_y2;
  wire f_u_arrmul24_fa8_17_y3;
  wire f_u_arrmul24_fa8_17_y4;
  wire f_u_arrmul24_and9_17_a_9;
  wire f_u_arrmul24_and9_17_b_17;
  wire f_u_arrmul24_and9_17_y0;
  wire f_u_arrmul24_fa9_17_f_u_arrmul24_and9_17_y0;
  wire f_u_arrmul24_fa9_17_f_u_arrmul24_fa10_16_y2;
  wire f_u_arrmul24_fa9_17_y0;
  wire f_u_arrmul24_fa9_17_y1;
  wire f_u_arrmul24_fa9_17_f_u_arrmul24_fa8_17_y4;
  wire f_u_arrmul24_fa9_17_y2;
  wire f_u_arrmul24_fa9_17_y3;
  wire f_u_arrmul24_fa9_17_y4;
  wire f_u_arrmul24_and10_17_a_10;
  wire f_u_arrmul24_and10_17_b_17;
  wire f_u_arrmul24_and10_17_y0;
  wire f_u_arrmul24_fa10_17_f_u_arrmul24_and10_17_y0;
  wire f_u_arrmul24_fa10_17_f_u_arrmul24_fa11_16_y2;
  wire f_u_arrmul24_fa10_17_y0;
  wire f_u_arrmul24_fa10_17_y1;
  wire f_u_arrmul24_fa10_17_f_u_arrmul24_fa9_17_y4;
  wire f_u_arrmul24_fa10_17_y2;
  wire f_u_arrmul24_fa10_17_y3;
  wire f_u_arrmul24_fa10_17_y4;
  wire f_u_arrmul24_and11_17_a_11;
  wire f_u_arrmul24_and11_17_b_17;
  wire f_u_arrmul24_and11_17_y0;
  wire f_u_arrmul24_fa11_17_f_u_arrmul24_and11_17_y0;
  wire f_u_arrmul24_fa11_17_f_u_arrmul24_fa12_16_y2;
  wire f_u_arrmul24_fa11_17_y0;
  wire f_u_arrmul24_fa11_17_y1;
  wire f_u_arrmul24_fa11_17_f_u_arrmul24_fa10_17_y4;
  wire f_u_arrmul24_fa11_17_y2;
  wire f_u_arrmul24_fa11_17_y3;
  wire f_u_arrmul24_fa11_17_y4;
  wire f_u_arrmul24_and12_17_a_12;
  wire f_u_arrmul24_and12_17_b_17;
  wire f_u_arrmul24_and12_17_y0;
  wire f_u_arrmul24_fa12_17_f_u_arrmul24_and12_17_y0;
  wire f_u_arrmul24_fa12_17_f_u_arrmul24_fa13_16_y2;
  wire f_u_arrmul24_fa12_17_y0;
  wire f_u_arrmul24_fa12_17_y1;
  wire f_u_arrmul24_fa12_17_f_u_arrmul24_fa11_17_y4;
  wire f_u_arrmul24_fa12_17_y2;
  wire f_u_arrmul24_fa12_17_y3;
  wire f_u_arrmul24_fa12_17_y4;
  wire f_u_arrmul24_and13_17_a_13;
  wire f_u_arrmul24_and13_17_b_17;
  wire f_u_arrmul24_and13_17_y0;
  wire f_u_arrmul24_fa13_17_f_u_arrmul24_and13_17_y0;
  wire f_u_arrmul24_fa13_17_f_u_arrmul24_fa14_16_y2;
  wire f_u_arrmul24_fa13_17_y0;
  wire f_u_arrmul24_fa13_17_y1;
  wire f_u_arrmul24_fa13_17_f_u_arrmul24_fa12_17_y4;
  wire f_u_arrmul24_fa13_17_y2;
  wire f_u_arrmul24_fa13_17_y3;
  wire f_u_arrmul24_fa13_17_y4;
  wire f_u_arrmul24_and14_17_a_14;
  wire f_u_arrmul24_and14_17_b_17;
  wire f_u_arrmul24_and14_17_y0;
  wire f_u_arrmul24_fa14_17_f_u_arrmul24_and14_17_y0;
  wire f_u_arrmul24_fa14_17_f_u_arrmul24_fa15_16_y2;
  wire f_u_arrmul24_fa14_17_y0;
  wire f_u_arrmul24_fa14_17_y1;
  wire f_u_arrmul24_fa14_17_f_u_arrmul24_fa13_17_y4;
  wire f_u_arrmul24_fa14_17_y2;
  wire f_u_arrmul24_fa14_17_y3;
  wire f_u_arrmul24_fa14_17_y4;
  wire f_u_arrmul24_and15_17_a_15;
  wire f_u_arrmul24_and15_17_b_17;
  wire f_u_arrmul24_and15_17_y0;
  wire f_u_arrmul24_fa15_17_f_u_arrmul24_and15_17_y0;
  wire f_u_arrmul24_fa15_17_f_u_arrmul24_fa16_16_y2;
  wire f_u_arrmul24_fa15_17_y0;
  wire f_u_arrmul24_fa15_17_y1;
  wire f_u_arrmul24_fa15_17_f_u_arrmul24_fa14_17_y4;
  wire f_u_arrmul24_fa15_17_y2;
  wire f_u_arrmul24_fa15_17_y3;
  wire f_u_arrmul24_fa15_17_y4;
  wire f_u_arrmul24_and16_17_a_16;
  wire f_u_arrmul24_and16_17_b_17;
  wire f_u_arrmul24_and16_17_y0;
  wire f_u_arrmul24_fa16_17_f_u_arrmul24_and16_17_y0;
  wire f_u_arrmul24_fa16_17_f_u_arrmul24_fa17_16_y2;
  wire f_u_arrmul24_fa16_17_y0;
  wire f_u_arrmul24_fa16_17_y1;
  wire f_u_arrmul24_fa16_17_f_u_arrmul24_fa15_17_y4;
  wire f_u_arrmul24_fa16_17_y2;
  wire f_u_arrmul24_fa16_17_y3;
  wire f_u_arrmul24_fa16_17_y4;
  wire f_u_arrmul24_and17_17_a_17;
  wire f_u_arrmul24_and17_17_b_17;
  wire f_u_arrmul24_and17_17_y0;
  wire f_u_arrmul24_fa17_17_f_u_arrmul24_and17_17_y0;
  wire f_u_arrmul24_fa17_17_f_u_arrmul24_fa18_16_y2;
  wire f_u_arrmul24_fa17_17_y0;
  wire f_u_arrmul24_fa17_17_y1;
  wire f_u_arrmul24_fa17_17_f_u_arrmul24_fa16_17_y4;
  wire f_u_arrmul24_fa17_17_y2;
  wire f_u_arrmul24_fa17_17_y3;
  wire f_u_arrmul24_fa17_17_y4;
  wire f_u_arrmul24_and18_17_a_18;
  wire f_u_arrmul24_and18_17_b_17;
  wire f_u_arrmul24_and18_17_y0;
  wire f_u_arrmul24_fa18_17_f_u_arrmul24_and18_17_y0;
  wire f_u_arrmul24_fa18_17_f_u_arrmul24_fa19_16_y2;
  wire f_u_arrmul24_fa18_17_y0;
  wire f_u_arrmul24_fa18_17_y1;
  wire f_u_arrmul24_fa18_17_f_u_arrmul24_fa17_17_y4;
  wire f_u_arrmul24_fa18_17_y2;
  wire f_u_arrmul24_fa18_17_y3;
  wire f_u_arrmul24_fa18_17_y4;
  wire f_u_arrmul24_and19_17_a_19;
  wire f_u_arrmul24_and19_17_b_17;
  wire f_u_arrmul24_and19_17_y0;
  wire f_u_arrmul24_fa19_17_f_u_arrmul24_and19_17_y0;
  wire f_u_arrmul24_fa19_17_f_u_arrmul24_fa20_16_y2;
  wire f_u_arrmul24_fa19_17_y0;
  wire f_u_arrmul24_fa19_17_y1;
  wire f_u_arrmul24_fa19_17_f_u_arrmul24_fa18_17_y4;
  wire f_u_arrmul24_fa19_17_y2;
  wire f_u_arrmul24_fa19_17_y3;
  wire f_u_arrmul24_fa19_17_y4;
  wire f_u_arrmul24_and20_17_a_20;
  wire f_u_arrmul24_and20_17_b_17;
  wire f_u_arrmul24_and20_17_y0;
  wire f_u_arrmul24_fa20_17_f_u_arrmul24_and20_17_y0;
  wire f_u_arrmul24_fa20_17_f_u_arrmul24_fa21_16_y2;
  wire f_u_arrmul24_fa20_17_y0;
  wire f_u_arrmul24_fa20_17_y1;
  wire f_u_arrmul24_fa20_17_f_u_arrmul24_fa19_17_y4;
  wire f_u_arrmul24_fa20_17_y2;
  wire f_u_arrmul24_fa20_17_y3;
  wire f_u_arrmul24_fa20_17_y4;
  wire f_u_arrmul24_and21_17_a_21;
  wire f_u_arrmul24_and21_17_b_17;
  wire f_u_arrmul24_and21_17_y0;
  wire f_u_arrmul24_fa21_17_f_u_arrmul24_and21_17_y0;
  wire f_u_arrmul24_fa21_17_f_u_arrmul24_fa22_16_y2;
  wire f_u_arrmul24_fa21_17_y0;
  wire f_u_arrmul24_fa21_17_y1;
  wire f_u_arrmul24_fa21_17_f_u_arrmul24_fa20_17_y4;
  wire f_u_arrmul24_fa21_17_y2;
  wire f_u_arrmul24_fa21_17_y3;
  wire f_u_arrmul24_fa21_17_y4;
  wire f_u_arrmul24_and22_17_a_22;
  wire f_u_arrmul24_and22_17_b_17;
  wire f_u_arrmul24_and22_17_y0;
  wire f_u_arrmul24_fa22_17_f_u_arrmul24_and22_17_y0;
  wire f_u_arrmul24_fa22_17_f_u_arrmul24_fa23_16_y2;
  wire f_u_arrmul24_fa22_17_y0;
  wire f_u_arrmul24_fa22_17_y1;
  wire f_u_arrmul24_fa22_17_f_u_arrmul24_fa21_17_y4;
  wire f_u_arrmul24_fa22_17_y2;
  wire f_u_arrmul24_fa22_17_y3;
  wire f_u_arrmul24_fa22_17_y4;
  wire f_u_arrmul24_and23_17_a_23;
  wire f_u_arrmul24_and23_17_b_17;
  wire f_u_arrmul24_and23_17_y0;
  wire f_u_arrmul24_fa23_17_f_u_arrmul24_and23_17_y0;
  wire f_u_arrmul24_fa23_17_f_u_arrmul24_fa23_16_y4;
  wire f_u_arrmul24_fa23_17_y0;
  wire f_u_arrmul24_fa23_17_y1;
  wire f_u_arrmul24_fa23_17_f_u_arrmul24_fa22_17_y4;
  wire f_u_arrmul24_fa23_17_y2;
  wire f_u_arrmul24_fa23_17_y3;
  wire f_u_arrmul24_fa23_17_y4;
  wire f_u_arrmul24_and0_18_a_0;
  wire f_u_arrmul24_and0_18_b_18;
  wire f_u_arrmul24_and0_18_y0;
  wire f_u_arrmul24_ha0_18_f_u_arrmul24_and0_18_y0;
  wire f_u_arrmul24_ha0_18_f_u_arrmul24_fa1_17_y2;
  wire f_u_arrmul24_ha0_18_y0;
  wire f_u_arrmul24_ha0_18_y1;
  wire f_u_arrmul24_and1_18_a_1;
  wire f_u_arrmul24_and1_18_b_18;
  wire f_u_arrmul24_and1_18_y0;
  wire f_u_arrmul24_fa1_18_f_u_arrmul24_and1_18_y0;
  wire f_u_arrmul24_fa1_18_f_u_arrmul24_fa2_17_y2;
  wire f_u_arrmul24_fa1_18_y0;
  wire f_u_arrmul24_fa1_18_y1;
  wire f_u_arrmul24_fa1_18_f_u_arrmul24_ha0_18_y1;
  wire f_u_arrmul24_fa1_18_y2;
  wire f_u_arrmul24_fa1_18_y3;
  wire f_u_arrmul24_fa1_18_y4;
  wire f_u_arrmul24_and2_18_a_2;
  wire f_u_arrmul24_and2_18_b_18;
  wire f_u_arrmul24_and2_18_y0;
  wire f_u_arrmul24_fa2_18_f_u_arrmul24_and2_18_y0;
  wire f_u_arrmul24_fa2_18_f_u_arrmul24_fa3_17_y2;
  wire f_u_arrmul24_fa2_18_y0;
  wire f_u_arrmul24_fa2_18_y1;
  wire f_u_arrmul24_fa2_18_f_u_arrmul24_fa1_18_y4;
  wire f_u_arrmul24_fa2_18_y2;
  wire f_u_arrmul24_fa2_18_y3;
  wire f_u_arrmul24_fa2_18_y4;
  wire f_u_arrmul24_and3_18_a_3;
  wire f_u_arrmul24_and3_18_b_18;
  wire f_u_arrmul24_and3_18_y0;
  wire f_u_arrmul24_fa3_18_f_u_arrmul24_and3_18_y0;
  wire f_u_arrmul24_fa3_18_f_u_arrmul24_fa4_17_y2;
  wire f_u_arrmul24_fa3_18_y0;
  wire f_u_arrmul24_fa3_18_y1;
  wire f_u_arrmul24_fa3_18_f_u_arrmul24_fa2_18_y4;
  wire f_u_arrmul24_fa3_18_y2;
  wire f_u_arrmul24_fa3_18_y3;
  wire f_u_arrmul24_fa3_18_y4;
  wire f_u_arrmul24_and4_18_a_4;
  wire f_u_arrmul24_and4_18_b_18;
  wire f_u_arrmul24_and4_18_y0;
  wire f_u_arrmul24_fa4_18_f_u_arrmul24_and4_18_y0;
  wire f_u_arrmul24_fa4_18_f_u_arrmul24_fa5_17_y2;
  wire f_u_arrmul24_fa4_18_y0;
  wire f_u_arrmul24_fa4_18_y1;
  wire f_u_arrmul24_fa4_18_f_u_arrmul24_fa3_18_y4;
  wire f_u_arrmul24_fa4_18_y2;
  wire f_u_arrmul24_fa4_18_y3;
  wire f_u_arrmul24_fa4_18_y4;
  wire f_u_arrmul24_and5_18_a_5;
  wire f_u_arrmul24_and5_18_b_18;
  wire f_u_arrmul24_and5_18_y0;
  wire f_u_arrmul24_fa5_18_f_u_arrmul24_and5_18_y0;
  wire f_u_arrmul24_fa5_18_f_u_arrmul24_fa6_17_y2;
  wire f_u_arrmul24_fa5_18_y0;
  wire f_u_arrmul24_fa5_18_y1;
  wire f_u_arrmul24_fa5_18_f_u_arrmul24_fa4_18_y4;
  wire f_u_arrmul24_fa5_18_y2;
  wire f_u_arrmul24_fa5_18_y3;
  wire f_u_arrmul24_fa5_18_y4;
  wire f_u_arrmul24_and6_18_a_6;
  wire f_u_arrmul24_and6_18_b_18;
  wire f_u_arrmul24_and6_18_y0;
  wire f_u_arrmul24_fa6_18_f_u_arrmul24_and6_18_y0;
  wire f_u_arrmul24_fa6_18_f_u_arrmul24_fa7_17_y2;
  wire f_u_arrmul24_fa6_18_y0;
  wire f_u_arrmul24_fa6_18_y1;
  wire f_u_arrmul24_fa6_18_f_u_arrmul24_fa5_18_y4;
  wire f_u_arrmul24_fa6_18_y2;
  wire f_u_arrmul24_fa6_18_y3;
  wire f_u_arrmul24_fa6_18_y4;
  wire f_u_arrmul24_and7_18_a_7;
  wire f_u_arrmul24_and7_18_b_18;
  wire f_u_arrmul24_and7_18_y0;
  wire f_u_arrmul24_fa7_18_f_u_arrmul24_and7_18_y0;
  wire f_u_arrmul24_fa7_18_f_u_arrmul24_fa8_17_y2;
  wire f_u_arrmul24_fa7_18_y0;
  wire f_u_arrmul24_fa7_18_y1;
  wire f_u_arrmul24_fa7_18_f_u_arrmul24_fa6_18_y4;
  wire f_u_arrmul24_fa7_18_y2;
  wire f_u_arrmul24_fa7_18_y3;
  wire f_u_arrmul24_fa7_18_y4;
  wire f_u_arrmul24_and8_18_a_8;
  wire f_u_arrmul24_and8_18_b_18;
  wire f_u_arrmul24_and8_18_y0;
  wire f_u_arrmul24_fa8_18_f_u_arrmul24_and8_18_y0;
  wire f_u_arrmul24_fa8_18_f_u_arrmul24_fa9_17_y2;
  wire f_u_arrmul24_fa8_18_y0;
  wire f_u_arrmul24_fa8_18_y1;
  wire f_u_arrmul24_fa8_18_f_u_arrmul24_fa7_18_y4;
  wire f_u_arrmul24_fa8_18_y2;
  wire f_u_arrmul24_fa8_18_y3;
  wire f_u_arrmul24_fa8_18_y4;
  wire f_u_arrmul24_and9_18_a_9;
  wire f_u_arrmul24_and9_18_b_18;
  wire f_u_arrmul24_and9_18_y0;
  wire f_u_arrmul24_fa9_18_f_u_arrmul24_and9_18_y0;
  wire f_u_arrmul24_fa9_18_f_u_arrmul24_fa10_17_y2;
  wire f_u_arrmul24_fa9_18_y0;
  wire f_u_arrmul24_fa9_18_y1;
  wire f_u_arrmul24_fa9_18_f_u_arrmul24_fa8_18_y4;
  wire f_u_arrmul24_fa9_18_y2;
  wire f_u_arrmul24_fa9_18_y3;
  wire f_u_arrmul24_fa9_18_y4;
  wire f_u_arrmul24_and10_18_a_10;
  wire f_u_arrmul24_and10_18_b_18;
  wire f_u_arrmul24_and10_18_y0;
  wire f_u_arrmul24_fa10_18_f_u_arrmul24_and10_18_y0;
  wire f_u_arrmul24_fa10_18_f_u_arrmul24_fa11_17_y2;
  wire f_u_arrmul24_fa10_18_y0;
  wire f_u_arrmul24_fa10_18_y1;
  wire f_u_arrmul24_fa10_18_f_u_arrmul24_fa9_18_y4;
  wire f_u_arrmul24_fa10_18_y2;
  wire f_u_arrmul24_fa10_18_y3;
  wire f_u_arrmul24_fa10_18_y4;
  wire f_u_arrmul24_and11_18_a_11;
  wire f_u_arrmul24_and11_18_b_18;
  wire f_u_arrmul24_and11_18_y0;
  wire f_u_arrmul24_fa11_18_f_u_arrmul24_and11_18_y0;
  wire f_u_arrmul24_fa11_18_f_u_arrmul24_fa12_17_y2;
  wire f_u_arrmul24_fa11_18_y0;
  wire f_u_arrmul24_fa11_18_y1;
  wire f_u_arrmul24_fa11_18_f_u_arrmul24_fa10_18_y4;
  wire f_u_arrmul24_fa11_18_y2;
  wire f_u_arrmul24_fa11_18_y3;
  wire f_u_arrmul24_fa11_18_y4;
  wire f_u_arrmul24_and12_18_a_12;
  wire f_u_arrmul24_and12_18_b_18;
  wire f_u_arrmul24_and12_18_y0;
  wire f_u_arrmul24_fa12_18_f_u_arrmul24_and12_18_y0;
  wire f_u_arrmul24_fa12_18_f_u_arrmul24_fa13_17_y2;
  wire f_u_arrmul24_fa12_18_y0;
  wire f_u_arrmul24_fa12_18_y1;
  wire f_u_arrmul24_fa12_18_f_u_arrmul24_fa11_18_y4;
  wire f_u_arrmul24_fa12_18_y2;
  wire f_u_arrmul24_fa12_18_y3;
  wire f_u_arrmul24_fa12_18_y4;
  wire f_u_arrmul24_and13_18_a_13;
  wire f_u_arrmul24_and13_18_b_18;
  wire f_u_arrmul24_and13_18_y0;
  wire f_u_arrmul24_fa13_18_f_u_arrmul24_and13_18_y0;
  wire f_u_arrmul24_fa13_18_f_u_arrmul24_fa14_17_y2;
  wire f_u_arrmul24_fa13_18_y0;
  wire f_u_arrmul24_fa13_18_y1;
  wire f_u_arrmul24_fa13_18_f_u_arrmul24_fa12_18_y4;
  wire f_u_arrmul24_fa13_18_y2;
  wire f_u_arrmul24_fa13_18_y3;
  wire f_u_arrmul24_fa13_18_y4;
  wire f_u_arrmul24_and14_18_a_14;
  wire f_u_arrmul24_and14_18_b_18;
  wire f_u_arrmul24_and14_18_y0;
  wire f_u_arrmul24_fa14_18_f_u_arrmul24_and14_18_y0;
  wire f_u_arrmul24_fa14_18_f_u_arrmul24_fa15_17_y2;
  wire f_u_arrmul24_fa14_18_y0;
  wire f_u_arrmul24_fa14_18_y1;
  wire f_u_arrmul24_fa14_18_f_u_arrmul24_fa13_18_y4;
  wire f_u_arrmul24_fa14_18_y2;
  wire f_u_arrmul24_fa14_18_y3;
  wire f_u_arrmul24_fa14_18_y4;
  wire f_u_arrmul24_and15_18_a_15;
  wire f_u_arrmul24_and15_18_b_18;
  wire f_u_arrmul24_and15_18_y0;
  wire f_u_arrmul24_fa15_18_f_u_arrmul24_and15_18_y0;
  wire f_u_arrmul24_fa15_18_f_u_arrmul24_fa16_17_y2;
  wire f_u_arrmul24_fa15_18_y0;
  wire f_u_arrmul24_fa15_18_y1;
  wire f_u_arrmul24_fa15_18_f_u_arrmul24_fa14_18_y4;
  wire f_u_arrmul24_fa15_18_y2;
  wire f_u_arrmul24_fa15_18_y3;
  wire f_u_arrmul24_fa15_18_y4;
  wire f_u_arrmul24_and16_18_a_16;
  wire f_u_arrmul24_and16_18_b_18;
  wire f_u_arrmul24_and16_18_y0;
  wire f_u_arrmul24_fa16_18_f_u_arrmul24_and16_18_y0;
  wire f_u_arrmul24_fa16_18_f_u_arrmul24_fa17_17_y2;
  wire f_u_arrmul24_fa16_18_y0;
  wire f_u_arrmul24_fa16_18_y1;
  wire f_u_arrmul24_fa16_18_f_u_arrmul24_fa15_18_y4;
  wire f_u_arrmul24_fa16_18_y2;
  wire f_u_arrmul24_fa16_18_y3;
  wire f_u_arrmul24_fa16_18_y4;
  wire f_u_arrmul24_and17_18_a_17;
  wire f_u_arrmul24_and17_18_b_18;
  wire f_u_arrmul24_and17_18_y0;
  wire f_u_arrmul24_fa17_18_f_u_arrmul24_and17_18_y0;
  wire f_u_arrmul24_fa17_18_f_u_arrmul24_fa18_17_y2;
  wire f_u_arrmul24_fa17_18_y0;
  wire f_u_arrmul24_fa17_18_y1;
  wire f_u_arrmul24_fa17_18_f_u_arrmul24_fa16_18_y4;
  wire f_u_arrmul24_fa17_18_y2;
  wire f_u_arrmul24_fa17_18_y3;
  wire f_u_arrmul24_fa17_18_y4;
  wire f_u_arrmul24_and18_18_a_18;
  wire f_u_arrmul24_and18_18_b_18;
  wire f_u_arrmul24_and18_18_y0;
  wire f_u_arrmul24_fa18_18_f_u_arrmul24_and18_18_y0;
  wire f_u_arrmul24_fa18_18_f_u_arrmul24_fa19_17_y2;
  wire f_u_arrmul24_fa18_18_y0;
  wire f_u_arrmul24_fa18_18_y1;
  wire f_u_arrmul24_fa18_18_f_u_arrmul24_fa17_18_y4;
  wire f_u_arrmul24_fa18_18_y2;
  wire f_u_arrmul24_fa18_18_y3;
  wire f_u_arrmul24_fa18_18_y4;
  wire f_u_arrmul24_and19_18_a_19;
  wire f_u_arrmul24_and19_18_b_18;
  wire f_u_arrmul24_and19_18_y0;
  wire f_u_arrmul24_fa19_18_f_u_arrmul24_and19_18_y0;
  wire f_u_arrmul24_fa19_18_f_u_arrmul24_fa20_17_y2;
  wire f_u_arrmul24_fa19_18_y0;
  wire f_u_arrmul24_fa19_18_y1;
  wire f_u_arrmul24_fa19_18_f_u_arrmul24_fa18_18_y4;
  wire f_u_arrmul24_fa19_18_y2;
  wire f_u_arrmul24_fa19_18_y3;
  wire f_u_arrmul24_fa19_18_y4;
  wire f_u_arrmul24_and20_18_a_20;
  wire f_u_arrmul24_and20_18_b_18;
  wire f_u_arrmul24_and20_18_y0;
  wire f_u_arrmul24_fa20_18_f_u_arrmul24_and20_18_y0;
  wire f_u_arrmul24_fa20_18_f_u_arrmul24_fa21_17_y2;
  wire f_u_arrmul24_fa20_18_y0;
  wire f_u_arrmul24_fa20_18_y1;
  wire f_u_arrmul24_fa20_18_f_u_arrmul24_fa19_18_y4;
  wire f_u_arrmul24_fa20_18_y2;
  wire f_u_arrmul24_fa20_18_y3;
  wire f_u_arrmul24_fa20_18_y4;
  wire f_u_arrmul24_and21_18_a_21;
  wire f_u_arrmul24_and21_18_b_18;
  wire f_u_arrmul24_and21_18_y0;
  wire f_u_arrmul24_fa21_18_f_u_arrmul24_and21_18_y0;
  wire f_u_arrmul24_fa21_18_f_u_arrmul24_fa22_17_y2;
  wire f_u_arrmul24_fa21_18_y0;
  wire f_u_arrmul24_fa21_18_y1;
  wire f_u_arrmul24_fa21_18_f_u_arrmul24_fa20_18_y4;
  wire f_u_arrmul24_fa21_18_y2;
  wire f_u_arrmul24_fa21_18_y3;
  wire f_u_arrmul24_fa21_18_y4;
  wire f_u_arrmul24_and22_18_a_22;
  wire f_u_arrmul24_and22_18_b_18;
  wire f_u_arrmul24_and22_18_y0;
  wire f_u_arrmul24_fa22_18_f_u_arrmul24_and22_18_y0;
  wire f_u_arrmul24_fa22_18_f_u_arrmul24_fa23_17_y2;
  wire f_u_arrmul24_fa22_18_y0;
  wire f_u_arrmul24_fa22_18_y1;
  wire f_u_arrmul24_fa22_18_f_u_arrmul24_fa21_18_y4;
  wire f_u_arrmul24_fa22_18_y2;
  wire f_u_arrmul24_fa22_18_y3;
  wire f_u_arrmul24_fa22_18_y4;
  wire f_u_arrmul24_and23_18_a_23;
  wire f_u_arrmul24_and23_18_b_18;
  wire f_u_arrmul24_and23_18_y0;
  wire f_u_arrmul24_fa23_18_f_u_arrmul24_and23_18_y0;
  wire f_u_arrmul24_fa23_18_f_u_arrmul24_fa23_17_y4;
  wire f_u_arrmul24_fa23_18_y0;
  wire f_u_arrmul24_fa23_18_y1;
  wire f_u_arrmul24_fa23_18_f_u_arrmul24_fa22_18_y4;
  wire f_u_arrmul24_fa23_18_y2;
  wire f_u_arrmul24_fa23_18_y3;
  wire f_u_arrmul24_fa23_18_y4;
  wire f_u_arrmul24_and0_19_a_0;
  wire f_u_arrmul24_and0_19_b_19;
  wire f_u_arrmul24_and0_19_y0;
  wire f_u_arrmul24_ha0_19_f_u_arrmul24_and0_19_y0;
  wire f_u_arrmul24_ha0_19_f_u_arrmul24_fa1_18_y2;
  wire f_u_arrmul24_ha0_19_y0;
  wire f_u_arrmul24_ha0_19_y1;
  wire f_u_arrmul24_and1_19_a_1;
  wire f_u_arrmul24_and1_19_b_19;
  wire f_u_arrmul24_and1_19_y0;
  wire f_u_arrmul24_fa1_19_f_u_arrmul24_and1_19_y0;
  wire f_u_arrmul24_fa1_19_f_u_arrmul24_fa2_18_y2;
  wire f_u_arrmul24_fa1_19_y0;
  wire f_u_arrmul24_fa1_19_y1;
  wire f_u_arrmul24_fa1_19_f_u_arrmul24_ha0_19_y1;
  wire f_u_arrmul24_fa1_19_y2;
  wire f_u_arrmul24_fa1_19_y3;
  wire f_u_arrmul24_fa1_19_y4;
  wire f_u_arrmul24_and2_19_a_2;
  wire f_u_arrmul24_and2_19_b_19;
  wire f_u_arrmul24_and2_19_y0;
  wire f_u_arrmul24_fa2_19_f_u_arrmul24_and2_19_y0;
  wire f_u_arrmul24_fa2_19_f_u_arrmul24_fa3_18_y2;
  wire f_u_arrmul24_fa2_19_y0;
  wire f_u_arrmul24_fa2_19_y1;
  wire f_u_arrmul24_fa2_19_f_u_arrmul24_fa1_19_y4;
  wire f_u_arrmul24_fa2_19_y2;
  wire f_u_arrmul24_fa2_19_y3;
  wire f_u_arrmul24_fa2_19_y4;
  wire f_u_arrmul24_and3_19_a_3;
  wire f_u_arrmul24_and3_19_b_19;
  wire f_u_arrmul24_and3_19_y0;
  wire f_u_arrmul24_fa3_19_f_u_arrmul24_and3_19_y0;
  wire f_u_arrmul24_fa3_19_f_u_arrmul24_fa4_18_y2;
  wire f_u_arrmul24_fa3_19_y0;
  wire f_u_arrmul24_fa3_19_y1;
  wire f_u_arrmul24_fa3_19_f_u_arrmul24_fa2_19_y4;
  wire f_u_arrmul24_fa3_19_y2;
  wire f_u_arrmul24_fa3_19_y3;
  wire f_u_arrmul24_fa3_19_y4;
  wire f_u_arrmul24_and4_19_a_4;
  wire f_u_arrmul24_and4_19_b_19;
  wire f_u_arrmul24_and4_19_y0;
  wire f_u_arrmul24_fa4_19_f_u_arrmul24_and4_19_y0;
  wire f_u_arrmul24_fa4_19_f_u_arrmul24_fa5_18_y2;
  wire f_u_arrmul24_fa4_19_y0;
  wire f_u_arrmul24_fa4_19_y1;
  wire f_u_arrmul24_fa4_19_f_u_arrmul24_fa3_19_y4;
  wire f_u_arrmul24_fa4_19_y2;
  wire f_u_arrmul24_fa4_19_y3;
  wire f_u_arrmul24_fa4_19_y4;
  wire f_u_arrmul24_and5_19_a_5;
  wire f_u_arrmul24_and5_19_b_19;
  wire f_u_arrmul24_and5_19_y0;
  wire f_u_arrmul24_fa5_19_f_u_arrmul24_and5_19_y0;
  wire f_u_arrmul24_fa5_19_f_u_arrmul24_fa6_18_y2;
  wire f_u_arrmul24_fa5_19_y0;
  wire f_u_arrmul24_fa5_19_y1;
  wire f_u_arrmul24_fa5_19_f_u_arrmul24_fa4_19_y4;
  wire f_u_arrmul24_fa5_19_y2;
  wire f_u_arrmul24_fa5_19_y3;
  wire f_u_arrmul24_fa5_19_y4;
  wire f_u_arrmul24_and6_19_a_6;
  wire f_u_arrmul24_and6_19_b_19;
  wire f_u_arrmul24_and6_19_y0;
  wire f_u_arrmul24_fa6_19_f_u_arrmul24_and6_19_y0;
  wire f_u_arrmul24_fa6_19_f_u_arrmul24_fa7_18_y2;
  wire f_u_arrmul24_fa6_19_y0;
  wire f_u_arrmul24_fa6_19_y1;
  wire f_u_arrmul24_fa6_19_f_u_arrmul24_fa5_19_y4;
  wire f_u_arrmul24_fa6_19_y2;
  wire f_u_arrmul24_fa6_19_y3;
  wire f_u_arrmul24_fa6_19_y4;
  wire f_u_arrmul24_and7_19_a_7;
  wire f_u_arrmul24_and7_19_b_19;
  wire f_u_arrmul24_and7_19_y0;
  wire f_u_arrmul24_fa7_19_f_u_arrmul24_and7_19_y0;
  wire f_u_arrmul24_fa7_19_f_u_arrmul24_fa8_18_y2;
  wire f_u_arrmul24_fa7_19_y0;
  wire f_u_arrmul24_fa7_19_y1;
  wire f_u_arrmul24_fa7_19_f_u_arrmul24_fa6_19_y4;
  wire f_u_arrmul24_fa7_19_y2;
  wire f_u_arrmul24_fa7_19_y3;
  wire f_u_arrmul24_fa7_19_y4;
  wire f_u_arrmul24_and8_19_a_8;
  wire f_u_arrmul24_and8_19_b_19;
  wire f_u_arrmul24_and8_19_y0;
  wire f_u_arrmul24_fa8_19_f_u_arrmul24_and8_19_y0;
  wire f_u_arrmul24_fa8_19_f_u_arrmul24_fa9_18_y2;
  wire f_u_arrmul24_fa8_19_y0;
  wire f_u_arrmul24_fa8_19_y1;
  wire f_u_arrmul24_fa8_19_f_u_arrmul24_fa7_19_y4;
  wire f_u_arrmul24_fa8_19_y2;
  wire f_u_arrmul24_fa8_19_y3;
  wire f_u_arrmul24_fa8_19_y4;
  wire f_u_arrmul24_and9_19_a_9;
  wire f_u_arrmul24_and9_19_b_19;
  wire f_u_arrmul24_and9_19_y0;
  wire f_u_arrmul24_fa9_19_f_u_arrmul24_and9_19_y0;
  wire f_u_arrmul24_fa9_19_f_u_arrmul24_fa10_18_y2;
  wire f_u_arrmul24_fa9_19_y0;
  wire f_u_arrmul24_fa9_19_y1;
  wire f_u_arrmul24_fa9_19_f_u_arrmul24_fa8_19_y4;
  wire f_u_arrmul24_fa9_19_y2;
  wire f_u_arrmul24_fa9_19_y3;
  wire f_u_arrmul24_fa9_19_y4;
  wire f_u_arrmul24_and10_19_a_10;
  wire f_u_arrmul24_and10_19_b_19;
  wire f_u_arrmul24_and10_19_y0;
  wire f_u_arrmul24_fa10_19_f_u_arrmul24_and10_19_y0;
  wire f_u_arrmul24_fa10_19_f_u_arrmul24_fa11_18_y2;
  wire f_u_arrmul24_fa10_19_y0;
  wire f_u_arrmul24_fa10_19_y1;
  wire f_u_arrmul24_fa10_19_f_u_arrmul24_fa9_19_y4;
  wire f_u_arrmul24_fa10_19_y2;
  wire f_u_arrmul24_fa10_19_y3;
  wire f_u_arrmul24_fa10_19_y4;
  wire f_u_arrmul24_and11_19_a_11;
  wire f_u_arrmul24_and11_19_b_19;
  wire f_u_arrmul24_and11_19_y0;
  wire f_u_arrmul24_fa11_19_f_u_arrmul24_and11_19_y0;
  wire f_u_arrmul24_fa11_19_f_u_arrmul24_fa12_18_y2;
  wire f_u_arrmul24_fa11_19_y0;
  wire f_u_arrmul24_fa11_19_y1;
  wire f_u_arrmul24_fa11_19_f_u_arrmul24_fa10_19_y4;
  wire f_u_arrmul24_fa11_19_y2;
  wire f_u_arrmul24_fa11_19_y3;
  wire f_u_arrmul24_fa11_19_y4;
  wire f_u_arrmul24_and12_19_a_12;
  wire f_u_arrmul24_and12_19_b_19;
  wire f_u_arrmul24_and12_19_y0;
  wire f_u_arrmul24_fa12_19_f_u_arrmul24_and12_19_y0;
  wire f_u_arrmul24_fa12_19_f_u_arrmul24_fa13_18_y2;
  wire f_u_arrmul24_fa12_19_y0;
  wire f_u_arrmul24_fa12_19_y1;
  wire f_u_arrmul24_fa12_19_f_u_arrmul24_fa11_19_y4;
  wire f_u_arrmul24_fa12_19_y2;
  wire f_u_arrmul24_fa12_19_y3;
  wire f_u_arrmul24_fa12_19_y4;
  wire f_u_arrmul24_and13_19_a_13;
  wire f_u_arrmul24_and13_19_b_19;
  wire f_u_arrmul24_and13_19_y0;
  wire f_u_arrmul24_fa13_19_f_u_arrmul24_and13_19_y0;
  wire f_u_arrmul24_fa13_19_f_u_arrmul24_fa14_18_y2;
  wire f_u_arrmul24_fa13_19_y0;
  wire f_u_arrmul24_fa13_19_y1;
  wire f_u_arrmul24_fa13_19_f_u_arrmul24_fa12_19_y4;
  wire f_u_arrmul24_fa13_19_y2;
  wire f_u_arrmul24_fa13_19_y3;
  wire f_u_arrmul24_fa13_19_y4;
  wire f_u_arrmul24_and14_19_a_14;
  wire f_u_arrmul24_and14_19_b_19;
  wire f_u_arrmul24_and14_19_y0;
  wire f_u_arrmul24_fa14_19_f_u_arrmul24_and14_19_y0;
  wire f_u_arrmul24_fa14_19_f_u_arrmul24_fa15_18_y2;
  wire f_u_arrmul24_fa14_19_y0;
  wire f_u_arrmul24_fa14_19_y1;
  wire f_u_arrmul24_fa14_19_f_u_arrmul24_fa13_19_y4;
  wire f_u_arrmul24_fa14_19_y2;
  wire f_u_arrmul24_fa14_19_y3;
  wire f_u_arrmul24_fa14_19_y4;
  wire f_u_arrmul24_and15_19_a_15;
  wire f_u_arrmul24_and15_19_b_19;
  wire f_u_arrmul24_and15_19_y0;
  wire f_u_arrmul24_fa15_19_f_u_arrmul24_and15_19_y0;
  wire f_u_arrmul24_fa15_19_f_u_arrmul24_fa16_18_y2;
  wire f_u_arrmul24_fa15_19_y0;
  wire f_u_arrmul24_fa15_19_y1;
  wire f_u_arrmul24_fa15_19_f_u_arrmul24_fa14_19_y4;
  wire f_u_arrmul24_fa15_19_y2;
  wire f_u_arrmul24_fa15_19_y3;
  wire f_u_arrmul24_fa15_19_y4;
  wire f_u_arrmul24_and16_19_a_16;
  wire f_u_arrmul24_and16_19_b_19;
  wire f_u_arrmul24_and16_19_y0;
  wire f_u_arrmul24_fa16_19_f_u_arrmul24_and16_19_y0;
  wire f_u_arrmul24_fa16_19_f_u_arrmul24_fa17_18_y2;
  wire f_u_arrmul24_fa16_19_y0;
  wire f_u_arrmul24_fa16_19_y1;
  wire f_u_arrmul24_fa16_19_f_u_arrmul24_fa15_19_y4;
  wire f_u_arrmul24_fa16_19_y2;
  wire f_u_arrmul24_fa16_19_y3;
  wire f_u_arrmul24_fa16_19_y4;
  wire f_u_arrmul24_and17_19_a_17;
  wire f_u_arrmul24_and17_19_b_19;
  wire f_u_arrmul24_and17_19_y0;
  wire f_u_arrmul24_fa17_19_f_u_arrmul24_and17_19_y0;
  wire f_u_arrmul24_fa17_19_f_u_arrmul24_fa18_18_y2;
  wire f_u_arrmul24_fa17_19_y0;
  wire f_u_arrmul24_fa17_19_y1;
  wire f_u_arrmul24_fa17_19_f_u_arrmul24_fa16_19_y4;
  wire f_u_arrmul24_fa17_19_y2;
  wire f_u_arrmul24_fa17_19_y3;
  wire f_u_arrmul24_fa17_19_y4;
  wire f_u_arrmul24_and18_19_a_18;
  wire f_u_arrmul24_and18_19_b_19;
  wire f_u_arrmul24_and18_19_y0;
  wire f_u_arrmul24_fa18_19_f_u_arrmul24_and18_19_y0;
  wire f_u_arrmul24_fa18_19_f_u_arrmul24_fa19_18_y2;
  wire f_u_arrmul24_fa18_19_y0;
  wire f_u_arrmul24_fa18_19_y1;
  wire f_u_arrmul24_fa18_19_f_u_arrmul24_fa17_19_y4;
  wire f_u_arrmul24_fa18_19_y2;
  wire f_u_arrmul24_fa18_19_y3;
  wire f_u_arrmul24_fa18_19_y4;
  wire f_u_arrmul24_and19_19_a_19;
  wire f_u_arrmul24_and19_19_b_19;
  wire f_u_arrmul24_and19_19_y0;
  wire f_u_arrmul24_fa19_19_f_u_arrmul24_and19_19_y0;
  wire f_u_arrmul24_fa19_19_f_u_arrmul24_fa20_18_y2;
  wire f_u_arrmul24_fa19_19_y0;
  wire f_u_arrmul24_fa19_19_y1;
  wire f_u_arrmul24_fa19_19_f_u_arrmul24_fa18_19_y4;
  wire f_u_arrmul24_fa19_19_y2;
  wire f_u_arrmul24_fa19_19_y3;
  wire f_u_arrmul24_fa19_19_y4;
  wire f_u_arrmul24_and20_19_a_20;
  wire f_u_arrmul24_and20_19_b_19;
  wire f_u_arrmul24_and20_19_y0;
  wire f_u_arrmul24_fa20_19_f_u_arrmul24_and20_19_y0;
  wire f_u_arrmul24_fa20_19_f_u_arrmul24_fa21_18_y2;
  wire f_u_arrmul24_fa20_19_y0;
  wire f_u_arrmul24_fa20_19_y1;
  wire f_u_arrmul24_fa20_19_f_u_arrmul24_fa19_19_y4;
  wire f_u_arrmul24_fa20_19_y2;
  wire f_u_arrmul24_fa20_19_y3;
  wire f_u_arrmul24_fa20_19_y4;
  wire f_u_arrmul24_and21_19_a_21;
  wire f_u_arrmul24_and21_19_b_19;
  wire f_u_arrmul24_and21_19_y0;
  wire f_u_arrmul24_fa21_19_f_u_arrmul24_and21_19_y0;
  wire f_u_arrmul24_fa21_19_f_u_arrmul24_fa22_18_y2;
  wire f_u_arrmul24_fa21_19_y0;
  wire f_u_arrmul24_fa21_19_y1;
  wire f_u_arrmul24_fa21_19_f_u_arrmul24_fa20_19_y4;
  wire f_u_arrmul24_fa21_19_y2;
  wire f_u_arrmul24_fa21_19_y3;
  wire f_u_arrmul24_fa21_19_y4;
  wire f_u_arrmul24_and22_19_a_22;
  wire f_u_arrmul24_and22_19_b_19;
  wire f_u_arrmul24_and22_19_y0;
  wire f_u_arrmul24_fa22_19_f_u_arrmul24_and22_19_y0;
  wire f_u_arrmul24_fa22_19_f_u_arrmul24_fa23_18_y2;
  wire f_u_arrmul24_fa22_19_y0;
  wire f_u_arrmul24_fa22_19_y1;
  wire f_u_arrmul24_fa22_19_f_u_arrmul24_fa21_19_y4;
  wire f_u_arrmul24_fa22_19_y2;
  wire f_u_arrmul24_fa22_19_y3;
  wire f_u_arrmul24_fa22_19_y4;
  wire f_u_arrmul24_and23_19_a_23;
  wire f_u_arrmul24_and23_19_b_19;
  wire f_u_arrmul24_and23_19_y0;
  wire f_u_arrmul24_fa23_19_f_u_arrmul24_and23_19_y0;
  wire f_u_arrmul24_fa23_19_f_u_arrmul24_fa23_18_y4;
  wire f_u_arrmul24_fa23_19_y0;
  wire f_u_arrmul24_fa23_19_y1;
  wire f_u_arrmul24_fa23_19_f_u_arrmul24_fa22_19_y4;
  wire f_u_arrmul24_fa23_19_y2;
  wire f_u_arrmul24_fa23_19_y3;
  wire f_u_arrmul24_fa23_19_y4;
  wire f_u_arrmul24_and0_20_a_0;
  wire f_u_arrmul24_and0_20_b_20;
  wire f_u_arrmul24_and0_20_y0;
  wire f_u_arrmul24_ha0_20_f_u_arrmul24_and0_20_y0;
  wire f_u_arrmul24_ha0_20_f_u_arrmul24_fa1_19_y2;
  wire f_u_arrmul24_ha0_20_y0;
  wire f_u_arrmul24_ha0_20_y1;
  wire f_u_arrmul24_and1_20_a_1;
  wire f_u_arrmul24_and1_20_b_20;
  wire f_u_arrmul24_and1_20_y0;
  wire f_u_arrmul24_fa1_20_f_u_arrmul24_and1_20_y0;
  wire f_u_arrmul24_fa1_20_f_u_arrmul24_fa2_19_y2;
  wire f_u_arrmul24_fa1_20_y0;
  wire f_u_arrmul24_fa1_20_y1;
  wire f_u_arrmul24_fa1_20_f_u_arrmul24_ha0_20_y1;
  wire f_u_arrmul24_fa1_20_y2;
  wire f_u_arrmul24_fa1_20_y3;
  wire f_u_arrmul24_fa1_20_y4;
  wire f_u_arrmul24_and2_20_a_2;
  wire f_u_arrmul24_and2_20_b_20;
  wire f_u_arrmul24_and2_20_y0;
  wire f_u_arrmul24_fa2_20_f_u_arrmul24_and2_20_y0;
  wire f_u_arrmul24_fa2_20_f_u_arrmul24_fa3_19_y2;
  wire f_u_arrmul24_fa2_20_y0;
  wire f_u_arrmul24_fa2_20_y1;
  wire f_u_arrmul24_fa2_20_f_u_arrmul24_fa1_20_y4;
  wire f_u_arrmul24_fa2_20_y2;
  wire f_u_arrmul24_fa2_20_y3;
  wire f_u_arrmul24_fa2_20_y4;
  wire f_u_arrmul24_and3_20_a_3;
  wire f_u_arrmul24_and3_20_b_20;
  wire f_u_arrmul24_and3_20_y0;
  wire f_u_arrmul24_fa3_20_f_u_arrmul24_and3_20_y0;
  wire f_u_arrmul24_fa3_20_f_u_arrmul24_fa4_19_y2;
  wire f_u_arrmul24_fa3_20_y0;
  wire f_u_arrmul24_fa3_20_y1;
  wire f_u_arrmul24_fa3_20_f_u_arrmul24_fa2_20_y4;
  wire f_u_arrmul24_fa3_20_y2;
  wire f_u_arrmul24_fa3_20_y3;
  wire f_u_arrmul24_fa3_20_y4;
  wire f_u_arrmul24_and4_20_a_4;
  wire f_u_arrmul24_and4_20_b_20;
  wire f_u_arrmul24_and4_20_y0;
  wire f_u_arrmul24_fa4_20_f_u_arrmul24_and4_20_y0;
  wire f_u_arrmul24_fa4_20_f_u_arrmul24_fa5_19_y2;
  wire f_u_arrmul24_fa4_20_y0;
  wire f_u_arrmul24_fa4_20_y1;
  wire f_u_arrmul24_fa4_20_f_u_arrmul24_fa3_20_y4;
  wire f_u_arrmul24_fa4_20_y2;
  wire f_u_arrmul24_fa4_20_y3;
  wire f_u_arrmul24_fa4_20_y4;
  wire f_u_arrmul24_and5_20_a_5;
  wire f_u_arrmul24_and5_20_b_20;
  wire f_u_arrmul24_and5_20_y0;
  wire f_u_arrmul24_fa5_20_f_u_arrmul24_and5_20_y0;
  wire f_u_arrmul24_fa5_20_f_u_arrmul24_fa6_19_y2;
  wire f_u_arrmul24_fa5_20_y0;
  wire f_u_arrmul24_fa5_20_y1;
  wire f_u_arrmul24_fa5_20_f_u_arrmul24_fa4_20_y4;
  wire f_u_arrmul24_fa5_20_y2;
  wire f_u_arrmul24_fa5_20_y3;
  wire f_u_arrmul24_fa5_20_y4;
  wire f_u_arrmul24_and6_20_a_6;
  wire f_u_arrmul24_and6_20_b_20;
  wire f_u_arrmul24_and6_20_y0;
  wire f_u_arrmul24_fa6_20_f_u_arrmul24_and6_20_y0;
  wire f_u_arrmul24_fa6_20_f_u_arrmul24_fa7_19_y2;
  wire f_u_arrmul24_fa6_20_y0;
  wire f_u_arrmul24_fa6_20_y1;
  wire f_u_arrmul24_fa6_20_f_u_arrmul24_fa5_20_y4;
  wire f_u_arrmul24_fa6_20_y2;
  wire f_u_arrmul24_fa6_20_y3;
  wire f_u_arrmul24_fa6_20_y4;
  wire f_u_arrmul24_and7_20_a_7;
  wire f_u_arrmul24_and7_20_b_20;
  wire f_u_arrmul24_and7_20_y0;
  wire f_u_arrmul24_fa7_20_f_u_arrmul24_and7_20_y0;
  wire f_u_arrmul24_fa7_20_f_u_arrmul24_fa8_19_y2;
  wire f_u_arrmul24_fa7_20_y0;
  wire f_u_arrmul24_fa7_20_y1;
  wire f_u_arrmul24_fa7_20_f_u_arrmul24_fa6_20_y4;
  wire f_u_arrmul24_fa7_20_y2;
  wire f_u_arrmul24_fa7_20_y3;
  wire f_u_arrmul24_fa7_20_y4;
  wire f_u_arrmul24_and8_20_a_8;
  wire f_u_arrmul24_and8_20_b_20;
  wire f_u_arrmul24_and8_20_y0;
  wire f_u_arrmul24_fa8_20_f_u_arrmul24_and8_20_y0;
  wire f_u_arrmul24_fa8_20_f_u_arrmul24_fa9_19_y2;
  wire f_u_arrmul24_fa8_20_y0;
  wire f_u_arrmul24_fa8_20_y1;
  wire f_u_arrmul24_fa8_20_f_u_arrmul24_fa7_20_y4;
  wire f_u_arrmul24_fa8_20_y2;
  wire f_u_arrmul24_fa8_20_y3;
  wire f_u_arrmul24_fa8_20_y4;
  wire f_u_arrmul24_and9_20_a_9;
  wire f_u_arrmul24_and9_20_b_20;
  wire f_u_arrmul24_and9_20_y0;
  wire f_u_arrmul24_fa9_20_f_u_arrmul24_and9_20_y0;
  wire f_u_arrmul24_fa9_20_f_u_arrmul24_fa10_19_y2;
  wire f_u_arrmul24_fa9_20_y0;
  wire f_u_arrmul24_fa9_20_y1;
  wire f_u_arrmul24_fa9_20_f_u_arrmul24_fa8_20_y4;
  wire f_u_arrmul24_fa9_20_y2;
  wire f_u_arrmul24_fa9_20_y3;
  wire f_u_arrmul24_fa9_20_y4;
  wire f_u_arrmul24_and10_20_a_10;
  wire f_u_arrmul24_and10_20_b_20;
  wire f_u_arrmul24_and10_20_y0;
  wire f_u_arrmul24_fa10_20_f_u_arrmul24_and10_20_y0;
  wire f_u_arrmul24_fa10_20_f_u_arrmul24_fa11_19_y2;
  wire f_u_arrmul24_fa10_20_y0;
  wire f_u_arrmul24_fa10_20_y1;
  wire f_u_arrmul24_fa10_20_f_u_arrmul24_fa9_20_y4;
  wire f_u_arrmul24_fa10_20_y2;
  wire f_u_arrmul24_fa10_20_y3;
  wire f_u_arrmul24_fa10_20_y4;
  wire f_u_arrmul24_and11_20_a_11;
  wire f_u_arrmul24_and11_20_b_20;
  wire f_u_arrmul24_and11_20_y0;
  wire f_u_arrmul24_fa11_20_f_u_arrmul24_and11_20_y0;
  wire f_u_arrmul24_fa11_20_f_u_arrmul24_fa12_19_y2;
  wire f_u_arrmul24_fa11_20_y0;
  wire f_u_arrmul24_fa11_20_y1;
  wire f_u_arrmul24_fa11_20_f_u_arrmul24_fa10_20_y4;
  wire f_u_arrmul24_fa11_20_y2;
  wire f_u_arrmul24_fa11_20_y3;
  wire f_u_arrmul24_fa11_20_y4;
  wire f_u_arrmul24_and12_20_a_12;
  wire f_u_arrmul24_and12_20_b_20;
  wire f_u_arrmul24_and12_20_y0;
  wire f_u_arrmul24_fa12_20_f_u_arrmul24_and12_20_y0;
  wire f_u_arrmul24_fa12_20_f_u_arrmul24_fa13_19_y2;
  wire f_u_arrmul24_fa12_20_y0;
  wire f_u_arrmul24_fa12_20_y1;
  wire f_u_arrmul24_fa12_20_f_u_arrmul24_fa11_20_y4;
  wire f_u_arrmul24_fa12_20_y2;
  wire f_u_arrmul24_fa12_20_y3;
  wire f_u_arrmul24_fa12_20_y4;
  wire f_u_arrmul24_and13_20_a_13;
  wire f_u_arrmul24_and13_20_b_20;
  wire f_u_arrmul24_and13_20_y0;
  wire f_u_arrmul24_fa13_20_f_u_arrmul24_and13_20_y0;
  wire f_u_arrmul24_fa13_20_f_u_arrmul24_fa14_19_y2;
  wire f_u_arrmul24_fa13_20_y0;
  wire f_u_arrmul24_fa13_20_y1;
  wire f_u_arrmul24_fa13_20_f_u_arrmul24_fa12_20_y4;
  wire f_u_arrmul24_fa13_20_y2;
  wire f_u_arrmul24_fa13_20_y3;
  wire f_u_arrmul24_fa13_20_y4;
  wire f_u_arrmul24_and14_20_a_14;
  wire f_u_arrmul24_and14_20_b_20;
  wire f_u_arrmul24_and14_20_y0;
  wire f_u_arrmul24_fa14_20_f_u_arrmul24_and14_20_y0;
  wire f_u_arrmul24_fa14_20_f_u_arrmul24_fa15_19_y2;
  wire f_u_arrmul24_fa14_20_y0;
  wire f_u_arrmul24_fa14_20_y1;
  wire f_u_arrmul24_fa14_20_f_u_arrmul24_fa13_20_y4;
  wire f_u_arrmul24_fa14_20_y2;
  wire f_u_arrmul24_fa14_20_y3;
  wire f_u_arrmul24_fa14_20_y4;
  wire f_u_arrmul24_and15_20_a_15;
  wire f_u_arrmul24_and15_20_b_20;
  wire f_u_arrmul24_and15_20_y0;
  wire f_u_arrmul24_fa15_20_f_u_arrmul24_and15_20_y0;
  wire f_u_arrmul24_fa15_20_f_u_arrmul24_fa16_19_y2;
  wire f_u_arrmul24_fa15_20_y0;
  wire f_u_arrmul24_fa15_20_y1;
  wire f_u_arrmul24_fa15_20_f_u_arrmul24_fa14_20_y4;
  wire f_u_arrmul24_fa15_20_y2;
  wire f_u_arrmul24_fa15_20_y3;
  wire f_u_arrmul24_fa15_20_y4;
  wire f_u_arrmul24_and16_20_a_16;
  wire f_u_arrmul24_and16_20_b_20;
  wire f_u_arrmul24_and16_20_y0;
  wire f_u_arrmul24_fa16_20_f_u_arrmul24_and16_20_y0;
  wire f_u_arrmul24_fa16_20_f_u_arrmul24_fa17_19_y2;
  wire f_u_arrmul24_fa16_20_y0;
  wire f_u_arrmul24_fa16_20_y1;
  wire f_u_arrmul24_fa16_20_f_u_arrmul24_fa15_20_y4;
  wire f_u_arrmul24_fa16_20_y2;
  wire f_u_arrmul24_fa16_20_y3;
  wire f_u_arrmul24_fa16_20_y4;
  wire f_u_arrmul24_and17_20_a_17;
  wire f_u_arrmul24_and17_20_b_20;
  wire f_u_arrmul24_and17_20_y0;
  wire f_u_arrmul24_fa17_20_f_u_arrmul24_and17_20_y0;
  wire f_u_arrmul24_fa17_20_f_u_arrmul24_fa18_19_y2;
  wire f_u_arrmul24_fa17_20_y0;
  wire f_u_arrmul24_fa17_20_y1;
  wire f_u_arrmul24_fa17_20_f_u_arrmul24_fa16_20_y4;
  wire f_u_arrmul24_fa17_20_y2;
  wire f_u_arrmul24_fa17_20_y3;
  wire f_u_arrmul24_fa17_20_y4;
  wire f_u_arrmul24_and18_20_a_18;
  wire f_u_arrmul24_and18_20_b_20;
  wire f_u_arrmul24_and18_20_y0;
  wire f_u_arrmul24_fa18_20_f_u_arrmul24_and18_20_y0;
  wire f_u_arrmul24_fa18_20_f_u_arrmul24_fa19_19_y2;
  wire f_u_arrmul24_fa18_20_y0;
  wire f_u_arrmul24_fa18_20_y1;
  wire f_u_arrmul24_fa18_20_f_u_arrmul24_fa17_20_y4;
  wire f_u_arrmul24_fa18_20_y2;
  wire f_u_arrmul24_fa18_20_y3;
  wire f_u_arrmul24_fa18_20_y4;
  wire f_u_arrmul24_and19_20_a_19;
  wire f_u_arrmul24_and19_20_b_20;
  wire f_u_arrmul24_and19_20_y0;
  wire f_u_arrmul24_fa19_20_f_u_arrmul24_and19_20_y0;
  wire f_u_arrmul24_fa19_20_f_u_arrmul24_fa20_19_y2;
  wire f_u_arrmul24_fa19_20_y0;
  wire f_u_arrmul24_fa19_20_y1;
  wire f_u_arrmul24_fa19_20_f_u_arrmul24_fa18_20_y4;
  wire f_u_arrmul24_fa19_20_y2;
  wire f_u_arrmul24_fa19_20_y3;
  wire f_u_arrmul24_fa19_20_y4;
  wire f_u_arrmul24_and20_20_a_20;
  wire f_u_arrmul24_and20_20_b_20;
  wire f_u_arrmul24_and20_20_y0;
  wire f_u_arrmul24_fa20_20_f_u_arrmul24_and20_20_y0;
  wire f_u_arrmul24_fa20_20_f_u_arrmul24_fa21_19_y2;
  wire f_u_arrmul24_fa20_20_y0;
  wire f_u_arrmul24_fa20_20_y1;
  wire f_u_arrmul24_fa20_20_f_u_arrmul24_fa19_20_y4;
  wire f_u_arrmul24_fa20_20_y2;
  wire f_u_arrmul24_fa20_20_y3;
  wire f_u_arrmul24_fa20_20_y4;
  wire f_u_arrmul24_and21_20_a_21;
  wire f_u_arrmul24_and21_20_b_20;
  wire f_u_arrmul24_and21_20_y0;
  wire f_u_arrmul24_fa21_20_f_u_arrmul24_and21_20_y0;
  wire f_u_arrmul24_fa21_20_f_u_arrmul24_fa22_19_y2;
  wire f_u_arrmul24_fa21_20_y0;
  wire f_u_arrmul24_fa21_20_y1;
  wire f_u_arrmul24_fa21_20_f_u_arrmul24_fa20_20_y4;
  wire f_u_arrmul24_fa21_20_y2;
  wire f_u_arrmul24_fa21_20_y3;
  wire f_u_arrmul24_fa21_20_y4;
  wire f_u_arrmul24_and22_20_a_22;
  wire f_u_arrmul24_and22_20_b_20;
  wire f_u_arrmul24_and22_20_y0;
  wire f_u_arrmul24_fa22_20_f_u_arrmul24_and22_20_y0;
  wire f_u_arrmul24_fa22_20_f_u_arrmul24_fa23_19_y2;
  wire f_u_arrmul24_fa22_20_y0;
  wire f_u_arrmul24_fa22_20_y1;
  wire f_u_arrmul24_fa22_20_f_u_arrmul24_fa21_20_y4;
  wire f_u_arrmul24_fa22_20_y2;
  wire f_u_arrmul24_fa22_20_y3;
  wire f_u_arrmul24_fa22_20_y4;
  wire f_u_arrmul24_and23_20_a_23;
  wire f_u_arrmul24_and23_20_b_20;
  wire f_u_arrmul24_and23_20_y0;
  wire f_u_arrmul24_fa23_20_f_u_arrmul24_and23_20_y0;
  wire f_u_arrmul24_fa23_20_f_u_arrmul24_fa23_19_y4;
  wire f_u_arrmul24_fa23_20_y0;
  wire f_u_arrmul24_fa23_20_y1;
  wire f_u_arrmul24_fa23_20_f_u_arrmul24_fa22_20_y4;
  wire f_u_arrmul24_fa23_20_y2;
  wire f_u_arrmul24_fa23_20_y3;
  wire f_u_arrmul24_fa23_20_y4;
  wire f_u_arrmul24_and0_21_a_0;
  wire f_u_arrmul24_and0_21_b_21;
  wire f_u_arrmul24_and0_21_y0;
  wire f_u_arrmul24_ha0_21_f_u_arrmul24_and0_21_y0;
  wire f_u_arrmul24_ha0_21_f_u_arrmul24_fa1_20_y2;
  wire f_u_arrmul24_ha0_21_y0;
  wire f_u_arrmul24_ha0_21_y1;
  wire f_u_arrmul24_and1_21_a_1;
  wire f_u_arrmul24_and1_21_b_21;
  wire f_u_arrmul24_and1_21_y0;
  wire f_u_arrmul24_fa1_21_f_u_arrmul24_and1_21_y0;
  wire f_u_arrmul24_fa1_21_f_u_arrmul24_fa2_20_y2;
  wire f_u_arrmul24_fa1_21_y0;
  wire f_u_arrmul24_fa1_21_y1;
  wire f_u_arrmul24_fa1_21_f_u_arrmul24_ha0_21_y1;
  wire f_u_arrmul24_fa1_21_y2;
  wire f_u_arrmul24_fa1_21_y3;
  wire f_u_arrmul24_fa1_21_y4;
  wire f_u_arrmul24_and2_21_a_2;
  wire f_u_arrmul24_and2_21_b_21;
  wire f_u_arrmul24_and2_21_y0;
  wire f_u_arrmul24_fa2_21_f_u_arrmul24_and2_21_y0;
  wire f_u_arrmul24_fa2_21_f_u_arrmul24_fa3_20_y2;
  wire f_u_arrmul24_fa2_21_y0;
  wire f_u_arrmul24_fa2_21_y1;
  wire f_u_arrmul24_fa2_21_f_u_arrmul24_fa1_21_y4;
  wire f_u_arrmul24_fa2_21_y2;
  wire f_u_arrmul24_fa2_21_y3;
  wire f_u_arrmul24_fa2_21_y4;
  wire f_u_arrmul24_and3_21_a_3;
  wire f_u_arrmul24_and3_21_b_21;
  wire f_u_arrmul24_and3_21_y0;
  wire f_u_arrmul24_fa3_21_f_u_arrmul24_and3_21_y0;
  wire f_u_arrmul24_fa3_21_f_u_arrmul24_fa4_20_y2;
  wire f_u_arrmul24_fa3_21_y0;
  wire f_u_arrmul24_fa3_21_y1;
  wire f_u_arrmul24_fa3_21_f_u_arrmul24_fa2_21_y4;
  wire f_u_arrmul24_fa3_21_y2;
  wire f_u_arrmul24_fa3_21_y3;
  wire f_u_arrmul24_fa3_21_y4;
  wire f_u_arrmul24_and4_21_a_4;
  wire f_u_arrmul24_and4_21_b_21;
  wire f_u_arrmul24_and4_21_y0;
  wire f_u_arrmul24_fa4_21_f_u_arrmul24_and4_21_y0;
  wire f_u_arrmul24_fa4_21_f_u_arrmul24_fa5_20_y2;
  wire f_u_arrmul24_fa4_21_y0;
  wire f_u_arrmul24_fa4_21_y1;
  wire f_u_arrmul24_fa4_21_f_u_arrmul24_fa3_21_y4;
  wire f_u_arrmul24_fa4_21_y2;
  wire f_u_arrmul24_fa4_21_y3;
  wire f_u_arrmul24_fa4_21_y4;
  wire f_u_arrmul24_and5_21_a_5;
  wire f_u_arrmul24_and5_21_b_21;
  wire f_u_arrmul24_and5_21_y0;
  wire f_u_arrmul24_fa5_21_f_u_arrmul24_and5_21_y0;
  wire f_u_arrmul24_fa5_21_f_u_arrmul24_fa6_20_y2;
  wire f_u_arrmul24_fa5_21_y0;
  wire f_u_arrmul24_fa5_21_y1;
  wire f_u_arrmul24_fa5_21_f_u_arrmul24_fa4_21_y4;
  wire f_u_arrmul24_fa5_21_y2;
  wire f_u_arrmul24_fa5_21_y3;
  wire f_u_arrmul24_fa5_21_y4;
  wire f_u_arrmul24_and6_21_a_6;
  wire f_u_arrmul24_and6_21_b_21;
  wire f_u_arrmul24_and6_21_y0;
  wire f_u_arrmul24_fa6_21_f_u_arrmul24_and6_21_y0;
  wire f_u_arrmul24_fa6_21_f_u_arrmul24_fa7_20_y2;
  wire f_u_arrmul24_fa6_21_y0;
  wire f_u_arrmul24_fa6_21_y1;
  wire f_u_arrmul24_fa6_21_f_u_arrmul24_fa5_21_y4;
  wire f_u_arrmul24_fa6_21_y2;
  wire f_u_arrmul24_fa6_21_y3;
  wire f_u_arrmul24_fa6_21_y4;
  wire f_u_arrmul24_and7_21_a_7;
  wire f_u_arrmul24_and7_21_b_21;
  wire f_u_arrmul24_and7_21_y0;
  wire f_u_arrmul24_fa7_21_f_u_arrmul24_and7_21_y0;
  wire f_u_arrmul24_fa7_21_f_u_arrmul24_fa8_20_y2;
  wire f_u_arrmul24_fa7_21_y0;
  wire f_u_arrmul24_fa7_21_y1;
  wire f_u_arrmul24_fa7_21_f_u_arrmul24_fa6_21_y4;
  wire f_u_arrmul24_fa7_21_y2;
  wire f_u_arrmul24_fa7_21_y3;
  wire f_u_arrmul24_fa7_21_y4;
  wire f_u_arrmul24_and8_21_a_8;
  wire f_u_arrmul24_and8_21_b_21;
  wire f_u_arrmul24_and8_21_y0;
  wire f_u_arrmul24_fa8_21_f_u_arrmul24_and8_21_y0;
  wire f_u_arrmul24_fa8_21_f_u_arrmul24_fa9_20_y2;
  wire f_u_arrmul24_fa8_21_y0;
  wire f_u_arrmul24_fa8_21_y1;
  wire f_u_arrmul24_fa8_21_f_u_arrmul24_fa7_21_y4;
  wire f_u_arrmul24_fa8_21_y2;
  wire f_u_arrmul24_fa8_21_y3;
  wire f_u_arrmul24_fa8_21_y4;
  wire f_u_arrmul24_and9_21_a_9;
  wire f_u_arrmul24_and9_21_b_21;
  wire f_u_arrmul24_and9_21_y0;
  wire f_u_arrmul24_fa9_21_f_u_arrmul24_and9_21_y0;
  wire f_u_arrmul24_fa9_21_f_u_arrmul24_fa10_20_y2;
  wire f_u_arrmul24_fa9_21_y0;
  wire f_u_arrmul24_fa9_21_y1;
  wire f_u_arrmul24_fa9_21_f_u_arrmul24_fa8_21_y4;
  wire f_u_arrmul24_fa9_21_y2;
  wire f_u_arrmul24_fa9_21_y3;
  wire f_u_arrmul24_fa9_21_y4;
  wire f_u_arrmul24_and10_21_a_10;
  wire f_u_arrmul24_and10_21_b_21;
  wire f_u_arrmul24_and10_21_y0;
  wire f_u_arrmul24_fa10_21_f_u_arrmul24_and10_21_y0;
  wire f_u_arrmul24_fa10_21_f_u_arrmul24_fa11_20_y2;
  wire f_u_arrmul24_fa10_21_y0;
  wire f_u_arrmul24_fa10_21_y1;
  wire f_u_arrmul24_fa10_21_f_u_arrmul24_fa9_21_y4;
  wire f_u_arrmul24_fa10_21_y2;
  wire f_u_arrmul24_fa10_21_y3;
  wire f_u_arrmul24_fa10_21_y4;
  wire f_u_arrmul24_and11_21_a_11;
  wire f_u_arrmul24_and11_21_b_21;
  wire f_u_arrmul24_and11_21_y0;
  wire f_u_arrmul24_fa11_21_f_u_arrmul24_and11_21_y0;
  wire f_u_arrmul24_fa11_21_f_u_arrmul24_fa12_20_y2;
  wire f_u_arrmul24_fa11_21_y0;
  wire f_u_arrmul24_fa11_21_y1;
  wire f_u_arrmul24_fa11_21_f_u_arrmul24_fa10_21_y4;
  wire f_u_arrmul24_fa11_21_y2;
  wire f_u_arrmul24_fa11_21_y3;
  wire f_u_arrmul24_fa11_21_y4;
  wire f_u_arrmul24_and12_21_a_12;
  wire f_u_arrmul24_and12_21_b_21;
  wire f_u_arrmul24_and12_21_y0;
  wire f_u_arrmul24_fa12_21_f_u_arrmul24_and12_21_y0;
  wire f_u_arrmul24_fa12_21_f_u_arrmul24_fa13_20_y2;
  wire f_u_arrmul24_fa12_21_y0;
  wire f_u_arrmul24_fa12_21_y1;
  wire f_u_arrmul24_fa12_21_f_u_arrmul24_fa11_21_y4;
  wire f_u_arrmul24_fa12_21_y2;
  wire f_u_arrmul24_fa12_21_y3;
  wire f_u_arrmul24_fa12_21_y4;
  wire f_u_arrmul24_and13_21_a_13;
  wire f_u_arrmul24_and13_21_b_21;
  wire f_u_arrmul24_and13_21_y0;
  wire f_u_arrmul24_fa13_21_f_u_arrmul24_and13_21_y0;
  wire f_u_arrmul24_fa13_21_f_u_arrmul24_fa14_20_y2;
  wire f_u_arrmul24_fa13_21_y0;
  wire f_u_arrmul24_fa13_21_y1;
  wire f_u_arrmul24_fa13_21_f_u_arrmul24_fa12_21_y4;
  wire f_u_arrmul24_fa13_21_y2;
  wire f_u_arrmul24_fa13_21_y3;
  wire f_u_arrmul24_fa13_21_y4;
  wire f_u_arrmul24_and14_21_a_14;
  wire f_u_arrmul24_and14_21_b_21;
  wire f_u_arrmul24_and14_21_y0;
  wire f_u_arrmul24_fa14_21_f_u_arrmul24_and14_21_y0;
  wire f_u_arrmul24_fa14_21_f_u_arrmul24_fa15_20_y2;
  wire f_u_arrmul24_fa14_21_y0;
  wire f_u_arrmul24_fa14_21_y1;
  wire f_u_arrmul24_fa14_21_f_u_arrmul24_fa13_21_y4;
  wire f_u_arrmul24_fa14_21_y2;
  wire f_u_arrmul24_fa14_21_y3;
  wire f_u_arrmul24_fa14_21_y4;
  wire f_u_arrmul24_and15_21_a_15;
  wire f_u_arrmul24_and15_21_b_21;
  wire f_u_arrmul24_and15_21_y0;
  wire f_u_arrmul24_fa15_21_f_u_arrmul24_and15_21_y0;
  wire f_u_arrmul24_fa15_21_f_u_arrmul24_fa16_20_y2;
  wire f_u_arrmul24_fa15_21_y0;
  wire f_u_arrmul24_fa15_21_y1;
  wire f_u_arrmul24_fa15_21_f_u_arrmul24_fa14_21_y4;
  wire f_u_arrmul24_fa15_21_y2;
  wire f_u_arrmul24_fa15_21_y3;
  wire f_u_arrmul24_fa15_21_y4;
  wire f_u_arrmul24_and16_21_a_16;
  wire f_u_arrmul24_and16_21_b_21;
  wire f_u_arrmul24_and16_21_y0;
  wire f_u_arrmul24_fa16_21_f_u_arrmul24_and16_21_y0;
  wire f_u_arrmul24_fa16_21_f_u_arrmul24_fa17_20_y2;
  wire f_u_arrmul24_fa16_21_y0;
  wire f_u_arrmul24_fa16_21_y1;
  wire f_u_arrmul24_fa16_21_f_u_arrmul24_fa15_21_y4;
  wire f_u_arrmul24_fa16_21_y2;
  wire f_u_arrmul24_fa16_21_y3;
  wire f_u_arrmul24_fa16_21_y4;
  wire f_u_arrmul24_and17_21_a_17;
  wire f_u_arrmul24_and17_21_b_21;
  wire f_u_arrmul24_and17_21_y0;
  wire f_u_arrmul24_fa17_21_f_u_arrmul24_and17_21_y0;
  wire f_u_arrmul24_fa17_21_f_u_arrmul24_fa18_20_y2;
  wire f_u_arrmul24_fa17_21_y0;
  wire f_u_arrmul24_fa17_21_y1;
  wire f_u_arrmul24_fa17_21_f_u_arrmul24_fa16_21_y4;
  wire f_u_arrmul24_fa17_21_y2;
  wire f_u_arrmul24_fa17_21_y3;
  wire f_u_arrmul24_fa17_21_y4;
  wire f_u_arrmul24_and18_21_a_18;
  wire f_u_arrmul24_and18_21_b_21;
  wire f_u_arrmul24_and18_21_y0;
  wire f_u_arrmul24_fa18_21_f_u_arrmul24_and18_21_y0;
  wire f_u_arrmul24_fa18_21_f_u_arrmul24_fa19_20_y2;
  wire f_u_arrmul24_fa18_21_y0;
  wire f_u_arrmul24_fa18_21_y1;
  wire f_u_arrmul24_fa18_21_f_u_arrmul24_fa17_21_y4;
  wire f_u_arrmul24_fa18_21_y2;
  wire f_u_arrmul24_fa18_21_y3;
  wire f_u_arrmul24_fa18_21_y4;
  wire f_u_arrmul24_and19_21_a_19;
  wire f_u_arrmul24_and19_21_b_21;
  wire f_u_arrmul24_and19_21_y0;
  wire f_u_arrmul24_fa19_21_f_u_arrmul24_and19_21_y0;
  wire f_u_arrmul24_fa19_21_f_u_arrmul24_fa20_20_y2;
  wire f_u_arrmul24_fa19_21_y0;
  wire f_u_arrmul24_fa19_21_y1;
  wire f_u_arrmul24_fa19_21_f_u_arrmul24_fa18_21_y4;
  wire f_u_arrmul24_fa19_21_y2;
  wire f_u_arrmul24_fa19_21_y3;
  wire f_u_arrmul24_fa19_21_y4;
  wire f_u_arrmul24_and20_21_a_20;
  wire f_u_arrmul24_and20_21_b_21;
  wire f_u_arrmul24_and20_21_y0;
  wire f_u_arrmul24_fa20_21_f_u_arrmul24_and20_21_y0;
  wire f_u_arrmul24_fa20_21_f_u_arrmul24_fa21_20_y2;
  wire f_u_arrmul24_fa20_21_y0;
  wire f_u_arrmul24_fa20_21_y1;
  wire f_u_arrmul24_fa20_21_f_u_arrmul24_fa19_21_y4;
  wire f_u_arrmul24_fa20_21_y2;
  wire f_u_arrmul24_fa20_21_y3;
  wire f_u_arrmul24_fa20_21_y4;
  wire f_u_arrmul24_and21_21_a_21;
  wire f_u_arrmul24_and21_21_b_21;
  wire f_u_arrmul24_and21_21_y0;
  wire f_u_arrmul24_fa21_21_f_u_arrmul24_and21_21_y0;
  wire f_u_arrmul24_fa21_21_f_u_arrmul24_fa22_20_y2;
  wire f_u_arrmul24_fa21_21_y0;
  wire f_u_arrmul24_fa21_21_y1;
  wire f_u_arrmul24_fa21_21_f_u_arrmul24_fa20_21_y4;
  wire f_u_arrmul24_fa21_21_y2;
  wire f_u_arrmul24_fa21_21_y3;
  wire f_u_arrmul24_fa21_21_y4;
  wire f_u_arrmul24_and22_21_a_22;
  wire f_u_arrmul24_and22_21_b_21;
  wire f_u_arrmul24_and22_21_y0;
  wire f_u_arrmul24_fa22_21_f_u_arrmul24_and22_21_y0;
  wire f_u_arrmul24_fa22_21_f_u_arrmul24_fa23_20_y2;
  wire f_u_arrmul24_fa22_21_y0;
  wire f_u_arrmul24_fa22_21_y1;
  wire f_u_arrmul24_fa22_21_f_u_arrmul24_fa21_21_y4;
  wire f_u_arrmul24_fa22_21_y2;
  wire f_u_arrmul24_fa22_21_y3;
  wire f_u_arrmul24_fa22_21_y4;
  wire f_u_arrmul24_and23_21_a_23;
  wire f_u_arrmul24_and23_21_b_21;
  wire f_u_arrmul24_and23_21_y0;
  wire f_u_arrmul24_fa23_21_f_u_arrmul24_and23_21_y0;
  wire f_u_arrmul24_fa23_21_f_u_arrmul24_fa23_20_y4;
  wire f_u_arrmul24_fa23_21_y0;
  wire f_u_arrmul24_fa23_21_y1;
  wire f_u_arrmul24_fa23_21_f_u_arrmul24_fa22_21_y4;
  wire f_u_arrmul24_fa23_21_y2;
  wire f_u_arrmul24_fa23_21_y3;
  wire f_u_arrmul24_fa23_21_y4;
  wire f_u_arrmul24_and0_22_a_0;
  wire f_u_arrmul24_and0_22_b_22;
  wire f_u_arrmul24_and0_22_y0;
  wire f_u_arrmul24_ha0_22_f_u_arrmul24_and0_22_y0;
  wire f_u_arrmul24_ha0_22_f_u_arrmul24_fa1_21_y2;
  wire f_u_arrmul24_ha0_22_y0;
  wire f_u_arrmul24_ha0_22_y1;
  wire f_u_arrmul24_and1_22_a_1;
  wire f_u_arrmul24_and1_22_b_22;
  wire f_u_arrmul24_and1_22_y0;
  wire f_u_arrmul24_fa1_22_f_u_arrmul24_and1_22_y0;
  wire f_u_arrmul24_fa1_22_f_u_arrmul24_fa2_21_y2;
  wire f_u_arrmul24_fa1_22_y0;
  wire f_u_arrmul24_fa1_22_y1;
  wire f_u_arrmul24_fa1_22_f_u_arrmul24_ha0_22_y1;
  wire f_u_arrmul24_fa1_22_y2;
  wire f_u_arrmul24_fa1_22_y3;
  wire f_u_arrmul24_fa1_22_y4;
  wire f_u_arrmul24_and2_22_a_2;
  wire f_u_arrmul24_and2_22_b_22;
  wire f_u_arrmul24_and2_22_y0;
  wire f_u_arrmul24_fa2_22_f_u_arrmul24_and2_22_y0;
  wire f_u_arrmul24_fa2_22_f_u_arrmul24_fa3_21_y2;
  wire f_u_arrmul24_fa2_22_y0;
  wire f_u_arrmul24_fa2_22_y1;
  wire f_u_arrmul24_fa2_22_f_u_arrmul24_fa1_22_y4;
  wire f_u_arrmul24_fa2_22_y2;
  wire f_u_arrmul24_fa2_22_y3;
  wire f_u_arrmul24_fa2_22_y4;
  wire f_u_arrmul24_and3_22_a_3;
  wire f_u_arrmul24_and3_22_b_22;
  wire f_u_arrmul24_and3_22_y0;
  wire f_u_arrmul24_fa3_22_f_u_arrmul24_and3_22_y0;
  wire f_u_arrmul24_fa3_22_f_u_arrmul24_fa4_21_y2;
  wire f_u_arrmul24_fa3_22_y0;
  wire f_u_arrmul24_fa3_22_y1;
  wire f_u_arrmul24_fa3_22_f_u_arrmul24_fa2_22_y4;
  wire f_u_arrmul24_fa3_22_y2;
  wire f_u_arrmul24_fa3_22_y3;
  wire f_u_arrmul24_fa3_22_y4;
  wire f_u_arrmul24_and4_22_a_4;
  wire f_u_arrmul24_and4_22_b_22;
  wire f_u_arrmul24_and4_22_y0;
  wire f_u_arrmul24_fa4_22_f_u_arrmul24_and4_22_y0;
  wire f_u_arrmul24_fa4_22_f_u_arrmul24_fa5_21_y2;
  wire f_u_arrmul24_fa4_22_y0;
  wire f_u_arrmul24_fa4_22_y1;
  wire f_u_arrmul24_fa4_22_f_u_arrmul24_fa3_22_y4;
  wire f_u_arrmul24_fa4_22_y2;
  wire f_u_arrmul24_fa4_22_y3;
  wire f_u_arrmul24_fa4_22_y4;
  wire f_u_arrmul24_and5_22_a_5;
  wire f_u_arrmul24_and5_22_b_22;
  wire f_u_arrmul24_and5_22_y0;
  wire f_u_arrmul24_fa5_22_f_u_arrmul24_and5_22_y0;
  wire f_u_arrmul24_fa5_22_f_u_arrmul24_fa6_21_y2;
  wire f_u_arrmul24_fa5_22_y0;
  wire f_u_arrmul24_fa5_22_y1;
  wire f_u_arrmul24_fa5_22_f_u_arrmul24_fa4_22_y4;
  wire f_u_arrmul24_fa5_22_y2;
  wire f_u_arrmul24_fa5_22_y3;
  wire f_u_arrmul24_fa5_22_y4;
  wire f_u_arrmul24_and6_22_a_6;
  wire f_u_arrmul24_and6_22_b_22;
  wire f_u_arrmul24_and6_22_y0;
  wire f_u_arrmul24_fa6_22_f_u_arrmul24_and6_22_y0;
  wire f_u_arrmul24_fa6_22_f_u_arrmul24_fa7_21_y2;
  wire f_u_arrmul24_fa6_22_y0;
  wire f_u_arrmul24_fa6_22_y1;
  wire f_u_arrmul24_fa6_22_f_u_arrmul24_fa5_22_y4;
  wire f_u_arrmul24_fa6_22_y2;
  wire f_u_arrmul24_fa6_22_y3;
  wire f_u_arrmul24_fa6_22_y4;
  wire f_u_arrmul24_and7_22_a_7;
  wire f_u_arrmul24_and7_22_b_22;
  wire f_u_arrmul24_and7_22_y0;
  wire f_u_arrmul24_fa7_22_f_u_arrmul24_and7_22_y0;
  wire f_u_arrmul24_fa7_22_f_u_arrmul24_fa8_21_y2;
  wire f_u_arrmul24_fa7_22_y0;
  wire f_u_arrmul24_fa7_22_y1;
  wire f_u_arrmul24_fa7_22_f_u_arrmul24_fa6_22_y4;
  wire f_u_arrmul24_fa7_22_y2;
  wire f_u_arrmul24_fa7_22_y3;
  wire f_u_arrmul24_fa7_22_y4;
  wire f_u_arrmul24_and8_22_a_8;
  wire f_u_arrmul24_and8_22_b_22;
  wire f_u_arrmul24_and8_22_y0;
  wire f_u_arrmul24_fa8_22_f_u_arrmul24_and8_22_y0;
  wire f_u_arrmul24_fa8_22_f_u_arrmul24_fa9_21_y2;
  wire f_u_arrmul24_fa8_22_y0;
  wire f_u_arrmul24_fa8_22_y1;
  wire f_u_arrmul24_fa8_22_f_u_arrmul24_fa7_22_y4;
  wire f_u_arrmul24_fa8_22_y2;
  wire f_u_arrmul24_fa8_22_y3;
  wire f_u_arrmul24_fa8_22_y4;
  wire f_u_arrmul24_and9_22_a_9;
  wire f_u_arrmul24_and9_22_b_22;
  wire f_u_arrmul24_and9_22_y0;
  wire f_u_arrmul24_fa9_22_f_u_arrmul24_and9_22_y0;
  wire f_u_arrmul24_fa9_22_f_u_arrmul24_fa10_21_y2;
  wire f_u_arrmul24_fa9_22_y0;
  wire f_u_arrmul24_fa9_22_y1;
  wire f_u_arrmul24_fa9_22_f_u_arrmul24_fa8_22_y4;
  wire f_u_arrmul24_fa9_22_y2;
  wire f_u_arrmul24_fa9_22_y3;
  wire f_u_arrmul24_fa9_22_y4;
  wire f_u_arrmul24_and10_22_a_10;
  wire f_u_arrmul24_and10_22_b_22;
  wire f_u_arrmul24_and10_22_y0;
  wire f_u_arrmul24_fa10_22_f_u_arrmul24_and10_22_y0;
  wire f_u_arrmul24_fa10_22_f_u_arrmul24_fa11_21_y2;
  wire f_u_arrmul24_fa10_22_y0;
  wire f_u_arrmul24_fa10_22_y1;
  wire f_u_arrmul24_fa10_22_f_u_arrmul24_fa9_22_y4;
  wire f_u_arrmul24_fa10_22_y2;
  wire f_u_arrmul24_fa10_22_y3;
  wire f_u_arrmul24_fa10_22_y4;
  wire f_u_arrmul24_and11_22_a_11;
  wire f_u_arrmul24_and11_22_b_22;
  wire f_u_arrmul24_and11_22_y0;
  wire f_u_arrmul24_fa11_22_f_u_arrmul24_and11_22_y0;
  wire f_u_arrmul24_fa11_22_f_u_arrmul24_fa12_21_y2;
  wire f_u_arrmul24_fa11_22_y0;
  wire f_u_arrmul24_fa11_22_y1;
  wire f_u_arrmul24_fa11_22_f_u_arrmul24_fa10_22_y4;
  wire f_u_arrmul24_fa11_22_y2;
  wire f_u_arrmul24_fa11_22_y3;
  wire f_u_arrmul24_fa11_22_y4;
  wire f_u_arrmul24_and12_22_a_12;
  wire f_u_arrmul24_and12_22_b_22;
  wire f_u_arrmul24_and12_22_y0;
  wire f_u_arrmul24_fa12_22_f_u_arrmul24_and12_22_y0;
  wire f_u_arrmul24_fa12_22_f_u_arrmul24_fa13_21_y2;
  wire f_u_arrmul24_fa12_22_y0;
  wire f_u_arrmul24_fa12_22_y1;
  wire f_u_arrmul24_fa12_22_f_u_arrmul24_fa11_22_y4;
  wire f_u_arrmul24_fa12_22_y2;
  wire f_u_arrmul24_fa12_22_y3;
  wire f_u_arrmul24_fa12_22_y4;
  wire f_u_arrmul24_and13_22_a_13;
  wire f_u_arrmul24_and13_22_b_22;
  wire f_u_arrmul24_and13_22_y0;
  wire f_u_arrmul24_fa13_22_f_u_arrmul24_and13_22_y0;
  wire f_u_arrmul24_fa13_22_f_u_arrmul24_fa14_21_y2;
  wire f_u_arrmul24_fa13_22_y0;
  wire f_u_arrmul24_fa13_22_y1;
  wire f_u_arrmul24_fa13_22_f_u_arrmul24_fa12_22_y4;
  wire f_u_arrmul24_fa13_22_y2;
  wire f_u_arrmul24_fa13_22_y3;
  wire f_u_arrmul24_fa13_22_y4;
  wire f_u_arrmul24_and14_22_a_14;
  wire f_u_arrmul24_and14_22_b_22;
  wire f_u_arrmul24_and14_22_y0;
  wire f_u_arrmul24_fa14_22_f_u_arrmul24_and14_22_y0;
  wire f_u_arrmul24_fa14_22_f_u_arrmul24_fa15_21_y2;
  wire f_u_arrmul24_fa14_22_y0;
  wire f_u_arrmul24_fa14_22_y1;
  wire f_u_arrmul24_fa14_22_f_u_arrmul24_fa13_22_y4;
  wire f_u_arrmul24_fa14_22_y2;
  wire f_u_arrmul24_fa14_22_y3;
  wire f_u_arrmul24_fa14_22_y4;
  wire f_u_arrmul24_and15_22_a_15;
  wire f_u_arrmul24_and15_22_b_22;
  wire f_u_arrmul24_and15_22_y0;
  wire f_u_arrmul24_fa15_22_f_u_arrmul24_and15_22_y0;
  wire f_u_arrmul24_fa15_22_f_u_arrmul24_fa16_21_y2;
  wire f_u_arrmul24_fa15_22_y0;
  wire f_u_arrmul24_fa15_22_y1;
  wire f_u_arrmul24_fa15_22_f_u_arrmul24_fa14_22_y4;
  wire f_u_arrmul24_fa15_22_y2;
  wire f_u_arrmul24_fa15_22_y3;
  wire f_u_arrmul24_fa15_22_y4;
  wire f_u_arrmul24_and16_22_a_16;
  wire f_u_arrmul24_and16_22_b_22;
  wire f_u_arrmul24_and16_22_y0;
  wire f_u_arrmul24_fa16_22_f_u_arrmul24_and16_22_y0;
  wire f_u_arrmul24_fa16_22_f_u_arrmul24_fa17_21_y2;
  wire f_u_arrmul24_fa16_22_y0;
  wire f_u_arrmul24_fa16_22_y1;
  wire f_u_arrmul24_fa16_22_f_u_arrmul24_fa15_22_y4;
  wire f_u_arrmul24_fa16_22_y2;
  wire f_u_arrmul24_fa16_22_y3;
  wire f_u_arrmul24_fa16_22_y4;
  wire f_u_arrmul24_and17_22_a_17;
  wire f_u_arrmul24_and17_22_b_22;
  wire f_u_arrmul24_and17_22_y0;
  wire f_u_arrmul24_fa17_22_f_u_arrmul24_and17_22_y0;
  wire f_u_arrmul24_fa17_22_f_u_arrmul24_fa18_21_y2;
  wire f_u_arrmul24_fa17_22_y0;
  wire f_u_arrmul24_fa17_22_y1;
  wire f_u_arrmul24_fa17_22_f_u_arrmul24_fa16_22_y4;
  wire f_u_arrmul24_fa17_22_y2;
  wire f_u_arrmul24_fa17_22_y3;
  wire f_u_arrmul24_fa17_22_y4;
  wire f_u_arrmul24_and18_22_a_18;
  wire f_u_arrmul24_and18_22_b_22;
  wire f_u_arrmul24_and18_22_y0;
  wire f_u_arrmul24_fa18_22_f_u_arrmul24_and18_22_y0;
  wire f_u_arrmul24_fa18_22_f_u_arrmul24_fa19_21_y2;
  wire f_u_arrmul24_fa18_22_y0;
  wire f_u_arrmul24_fa18_22_y1;
  wire f_u_arrmul24_fa18_22_f_u_arrmul24_fa17_22_y4;
  wire f_u_arrmul24_fa18_22_y2;
  wire f_u_arrmul24_fa18_22_y3;
  wire f_u_arrmul24_fa18_22_y4;
  wire f_u_arrmul24_and19_22_a_19;
  wire f_u_arrmul24_and19_22_b_22;
  wire f_u_arrmul24_and19_22_y0;
  wire f_u_arrmul24_fa19_22_f_u_arrmul24_and19_22_y0;
  wire f_u_arrmul24_fa19_22_f_u_arrmul24_fa20_21_y2;
  wire f_u_arrmul24_fa19_22_y0;
  wire f_u_arrmul24_fa19_22_y1;
  wire f_u_arrmul24_fa19_22_f_u_arrmul24_fa18_22_y4;
  wire f_u_arrmul24_fa19_22_y2;
  wire f_u_arrmul24_fa19_22_y3;
  wire f_u_arrmul24_fa19_22_y4;
  wire f_u_arrmul24_and20_22_a_20;
  wire f_u_arrmul24_and20_22_b_22;
  wire f_u_arrmul24_and20_22_y0;
  wire f_u_arrmul24_fa20_22_f_u_arrmul24_and20_22_y0;
  wire f_u_arrmul24_fa20_22_f_u_arrmul24_fa21_21_y2;
  wire f_u_arrmul24_fa20_22_y0;
  wire f_u_arrmul24_fa20_22_y1;
  wire f_u_arrmul24_fa20_22_f_u_arrmul24_fa19_22_y4;
  wire f_u_arrmul24_fa20_22_y2;
  wire f_u_arrmul24_fa20_22_y3;
  wire f_u_arrmul24_fa20_22_y4;
  wire f_u_arrmul24_and21_22_a_21;
  wire f_u_arrmul24_and21_22_b_22;
  wire f_u_arrmul24_and21_22_y0;
  wire f_u_arrmul24_fa21_22_f_u_arrmul24_and21_22_y0;
  wire f_u_arrmul24_fa21_22_f_u_arrmul24_fa22_21_y2;
  wire f_u_arrmul24_fa21_22_y0;
  wire f_u_arrmul24_fa21_22_y1;
  wire f_u_arrmul24_fa21_22_f_u_arrmul24_fa20_22_y4;
  wire f_u_arrmul24_fa21_22_y2;
  wire f_u_arrmul24_fa21_22_y3;
  wire f_u_arrmul24_fa21_22_y4;
  wire f_u_arrmul24_and22_22_a_22;
  wire f_u_arrmul24_and22_22_b_22;
  wire f_u_arrmul24_and22_22_y0;
  wire f_u_arrmul24_fa22_22_f_u_arrmul24_and22_22_y0;
  wire f_u_arrmul24_fa22_22_f_u_arrmul24_fa23_21_y2;
  wire f_u_arrmul24_fa22_22_y0;
  wire f_u_arrmul24_fa22_22_y1;
  wire f_u_arrmul24_fa22_22_f_u_arrmul24_fa21_22_y4;
  wire f_u_arrmul24_fa22_22_y2;
  wire f_u_arrmul24_fa22_22_y3;
  wire f_u_arrmul24_fa22_22_y4;
  wire f_u_arrmul24_and23_22_a_23;
  wire f_u_arrmul24_and23_22_b_22;
  wire f_u_arrmul24_and23_22_y0;
  wire f_u_arrmul24_fa23_22_f_u_arrmul24_and23_22_y0;
  wire f_u_arrmul24_fa23_22_f_u_arrmul24_fa23_21_y4;
  wire f_u_arrmul24_fa23_22_y0;
  wire f_u_arrmul24_fa23_22_y1;
  wire f_u_arrmul24_fa23_22_f_u_arrmul24_fa22_22_y4;
  wire f_u_arrmul24_fa23_22_y2;
  wire f_u_arrmul24_fa23_22_y3;
  wire f_u_arrmul24_fa23_22_y4;
  wire f_u_arrmul24_and0_23_a_0;
  wire f_u_arrmul24_and0_23_b_23;
  wire f_u_arrmul24_and0_23_y0;
  wire f_u_arrmul24_ha0_23_f_u_arrmul24_and0_23_y0;
  wire f_u_arrmul24_ha0_23_f_u_arrmul24_fa1_22_y2;
  wire f_u_arrmul24_ha0_23_y0;
  wire f_u_arrmul24_ha0_23_y1;
  wire f_u_arrmul24_and1_23_a_1;
  wire f_u_arrmul24_and1_23_b_23;
  wire f_u_arrmul24_and1_23_y0;
  wire f_u_arrmul24_fa1_23_f_u_arrmul24_and1_23_y0;
  wire f_u_arrmul24_fa1_23_f_u_arrmul24_fa2_22_y2;
  wire f_u_arrmul24_fa1_23_y0;
  wire f_u_arrmul24_fa1_23_y1;
  wire f_u_arrmul24_fa1_23_f_u_arrmul24_ha0_23_y1;
  wire f_u_arrmul24_fa1_23_y2;
  wire f_u_arrmul24_fa1_23_y3;
  wire f_u_arrmul24_fa1_23_y4;
  wire f_u_arrmul24_and2_23_a_2;
  wire f_u_arrmul24_and2_23_b_23;
  wire f_u_arrmul24_and2_23_y0;
  wire f_u_arrmul24_fa2_23_f_u_arrmul24_and2_23_y0;
  wire f_u_arrmul24_fa2_23_f_u_arrmul24_fa3_22_y2;
  wire f_u_arrmul24_fa2_23_y0;
  wire f_u_arrmul24_fa2_23_y1;
  wire f_u_arrmul24_fa2_23_f_u_arrmul24_fa1_23_y4;
  wire f_u_arrmul24_fa2_23_y2;
  wire f_u_arrmul24_fa2_23_y3;
  wire f_u_arrmul24_fa2_23_y4;
  wire f_u_arrmul24_and3_23_a_3;
  wire f_u_arrmul24_and3_23_b_23;
  wire f_u_arrmul24_and3_23_y0;
  wire f_u_arrmul24_fa3_23_f_u_arrmul24_and3_23_y0;
  wire f_u_arrmul24_fa3_23_f_u_arrmul24_fa4_22_y2;
  wire f_u_arrmul24_fa3_23_y0;
  wire f_u_arrmul24_fa3_23_y1;
  wire f_u_arrmul24_fa3_23_f_u_arrmul24_fa2_23_y4;
  wire f_u_arrmul24_fa3_23_y2;
  wire f_u_arrmul24_fa3_23_y3;
  wire f_u_arrmul24_fa3_23_y4;
  wire f_u_arrmul24_and4_23_a_4;
  wire f_u_arrmul24_and4_23_b_23;
  wire f_u_arrmul24_and4_23_y0;
  wire f_u_arrmul24_fa4_23_f_u_arrmul24_and4_23_y0;
  wire f_u_arrmul24_fa4_23_f_u_arrmul24_fa5_22_y2;
  wire f_u_arrmul24_fa4_23_y0;
  wire f_u_arrmul24_fa4_23_y1;
  wire f_u_arrmul24_fa4_23_f_u_arrmul24_fa3_23_y4;
  wire f_u_arrmul24_fa4_23_y2;
  wire f_u_arrmul24_fa4_23_y3;
  wire f_u_arrmul24_fa4_23_y4;
  wire f_u_arrmul24_and5_23_a_5;
  wire f_u_arrmul24_and5_23_b_23;
  wire f_u_arrmul24_and5_23_y0;
  wire f_u_arrmul24_fa5_23_f_u_arrmul24_and5_23_y0;
  wire f_u_arrmul24_fa5_23_f_u_arrmul24_fa6_22_y2;
  wire f_u_arrmul24_fa5_23_y0;
  wire f_u_arrmul24_fa5_23_y1;
  wire f_u_arrmul24_fa5_23_f_u_arrmul24_fa4_23_y4;
  wire f_u_arrmul24_fa5_23_y2;
  wire f_u_arrmul24_fa5_23_y3;
  wire f_u_arrmul24_fa5_23_y4;
  wire f_u_arrmul24_and6_23_a_6;
  wire f_u_arrmul24_and6_23_b_23;
  wire f_u_arrmul24_and6_23_y0;
  wire f_u_arrmul24_fa6_23_f_u_arrmul24_and6_23_y0;
  wire f_u_arrmul24_fa6_23_f_u_arrmul24_fa7_22_y2;
  wire f_u_arrmul24_fa6_23_y0;
  wire f_u_arrmul24_fa6_23_y1;
  wire f_u_arrmul24_fa6_23_f_u_arrmul24_fa5_23_y4;
  wire f_u_arrmul24_fa6_23_y2;
  wire f_u_arrmul24_fa6_23_y3;
  wire f_u_arrmul24_fa6_23_y4;
  wire f_u_arrmul24_and7_23_a_7;
  wire f_u_arrmul24_and7_23_b_23;
  wire f_u_arrmul24_and7_23_y0;
  wire f_u_arrmul24_fa7_23_f_u_arrmul24_and7_23_y0;
  wire f_u_arrmul24_fa7_23_f_u_arrmul24_fa8_22_y2;
  wire f_u_arrmul24_fa7_23_y0;
  wire f_u_arrmul24_fa7_23_y1;
  wire f_u_arrmul24_fa7_23_f_u_arrmul24_fa6_23_y4;
  wire f_u_arrmul24_fa7_23_y2;
  wire f_u_arrmul24_fa7_23_y3;
  wire f_u_arrmul24_fa7_23_y4;
  wire f_u_arrmul24_and8_23_a_8;
  wire f_u_arrmul24_and8_23_b_23;
  wire f_u_arrmul24_and8_23_y0;
  wire f_u_arrmul24_fa8_23_f_u_arrmul24_and8_23_y0;
  wire f_u_arrmul24_fa8_23_f_u_arrmul24_fa9_22_y2;
  wire f_u_arrmul24_fa8_23_y0;
  wire f_u_arrmul24_fa8_23_y1;
  wire f_u_arrmul24_fa8_23_f_u_arrmul24_fa7_23_y4;
  wire f_u_arrmul24_fa8_23_y2;
  wire f_u_arrmul24_fa8_23_y3;
  wire f_u_arrmul24_fa8_23_y4;
  wire f_u_arrmul24_and9_23_a_9;
  wire f_u_arrmul24_and9_23_b_23;
  wire f_u_arrmul24_and9_23_y0;
  wire f_u_arrmul24_fa9_23_f_u_arrmul24_and9_23_y0;
  wire f_u_arrmul24_fa9_23_f_u_arrmul24_fa10_22_y2;
  wire f_u_arrmul24_fa9_23_y0;
  wire f_u_arrmul24_fa9_23_y1;
  wire f_u_arrmul24_fa9_23_f_u_arrmul24_fa8_23_y4;
  wire f_u_arrmul24_fa9_23_y2;
  wire f_u_arrmul24_fa9_23_y3;
  wire f_u_arrmul24_fa9_23_y4;
  wire f_u_arrmul24_and10_23_a_10;
  wire f_u_arrmul24_and10_23_b_23;
  wire f_u_arrmul24_and10_23_y0;
  wire f_u_arrmul24_fa10_23_f_u_arrmul24_and10_23_y0;
  wire f_u_arrmul24_fa10_23_f_u_arrmul24_fa11_22_y2;
  wire f_u_arrmul24_fa10_23_y0;
  wire f_u_arrmul24_fa10_23_y1;
  wire f_u_arrmul24_fa10_23_f_u_arrmul24_fa9_23_y4;
  wire f_u_arrmul24_fa10_23_y2;
  wire f_u_arrmul24_fa10_23_y3;
  wire f_u_arrmul24_fa10_23_y4;
  wire f_u_arrmul24_and11_23_a_11;
  wire f_u_arrmul24_and11_23_b_23;
  wire f_u_arrmul24_and11_23_y0;
  wire f_u_arrmul24_fa11_23_f_u_arrmul24_and11_23_y0;
  wire f_u_arrmul24_fa11_23_f_u_arrmul24_fa12_22_y2;
  wire f_u_arrmul24_fa11_23_y0;
  wire f_u_arrmul24_fa11_23_y1;
  wire f_u_arrmul24_fa11_23_f_u_arrmul24_fa10_23_y4;
  wire f_u_arrmul24_fa11_23_y2;
  wire f_u_arrmul24_fa11_23_y3;
  wire f_u_arrmul24_fa11_23_y4;
  wire f_u_arrmul24_and12_23_a_12;
  wire f_u_arrmul24_and12_23_b_23;
  wire f_u_arrmul24_and12_23_y0;
  wire f_u_arrmul24_fa12_23_f_u_arrmul24_and12_23_y0;
  wire f_u_arrmul24_fa12_23_f_u_arrmul24_fa13_22_y2;
  wire f_u_arrmul24_fa12_23_y0;
  wire f_u_arrmul24_fa12_23_y1;
  wire f_u_arrmul24_fa12_23_f_u_arrmul24_fa11_23_y4;
  wire f_u_arrmul24_fa12_23_y2;
  wire f_u_arrmul24_fa12_23_y3;
  wire f_u_arrmul24_fa12_23_y4;
  wire f_u_arrmul24_and13_23_a_13;
  wire f_u_arrmul24_and13_23_b_23;
  wire f_u_arrmul24_and13_23_y0;
  wire f_u_arrmul24_fa13_23_f_u_arrmul24_and13_23_y0;
  wire f_u_arrmul24_fa13_23_f_u_arrmul24_fa14_22_y2;
  wire f_u_arrmul24_fa13_23_y0;
  wire f_u_arrmul24_fa13_23_y1;
  wire f_u_arrmul24_fa13_23_f_u_arrmul24_fa12_23_y4;
  wire f_u_arrmul24_fa13_23_y2;
  wire f_u_arrmul24_fa13_23_y3;
  wire f_u_arrmul24_fa13_23_y4;
  wire f_u_arrmul24_and14_23_a_14;
  wire f_u_arrmul24_and14_23_b_23;
  wire f_u_arrmul24_and14_23_y0;
  wire f_u_arrmul24_fa14_23_f_u_arrmul24_and14_23_y0;
  wire f_u_arrmul24_fa14_23_f_u_arrmul24_fa15_22_y2;
  wire f_u_arrmul24_fa14_23_y0;
  wire f_u_arrmul24_fa14_23_y1;
  wire f_u_arrmul24_fa14_23_f_u_arrmul24_fa13_23_y4;
  wire f_u_arrmul24_fa14_23_y2;
  wire f_u_arrmul24_fa14_23_y3;
  wire f_u_arrmul24_fa14_23_y4;
  wire f_u_arrmul24_and15_23_a_15;
  wire f_u_arrmul24_and15_23_b_23;
  wire f_u_arrmul24_and15_23_y0;
  wire f_u_arrmul24_fa15_23_f_u_arrmul24_and15_23_y0;
  wire f_u_arrmul24_fa15_23_f_u_arrmul24_fa16_22_y2;
  wire f_u_arrmul24_fa15_23_y0;
  wire f_u_arrmul24_fa15_23_y1;
  wire f_u_arrmul24_fa15_23_f_u_arrmul24_fa14_23_y4;
  wire f_u_arrmul24_fa15_23_y2;
  wire f_u_arrmul24_fa15_23_y3;
  wire f_u_arrmul24_fa15_23_y4;
  wire f_u_arrmul24_and16_23_a_16;
  wire f_u_arrmul24_and16_23_b_23;
  wire f_u_arrmul24_and16_23_y0;
  wire f_u_arrmul24_fa16_23_f_u_arrmul24_and16_23_y0;
  wire f_u_arrmul24_fa16_23_f_u_arrmul24_fa17_22_y2;
  wire f_u_arrmul24_fa16_23_y0;
  wire f_u_arrmul24_fa16_23_y1;
  wire f_u_arrmul24_fa16_23_f_u_arrmul24_fa15_23_y4;
  wire f_u_arrmul24_fa16_23_y2;
  wire f_u_arrmul24_fa16_23_y3;
  wire f_u_arrmul24_fa16_23_y4;
  wire f_u_arrmul24_and17_23_a_17;
  wire f_u_arrmul24_and17_23_b_23;
  wire f_u_arrmul24_and17_23_y0;
  wire f_u_arrmul24_fa17_23_f_u_arrmul24_and17_23_y0;
  wire f_u_arrmul24_fa17_23_f_u_arrmul24_fa18_22_y2;
  wire f_u_arrmul24_fa17_23_y0;
  wire f_u_arrmul24_fa17_23_y1;
  wire f_u_arrmul24_fa17_23_f_u_arrmul24_fa16_23_y4;
  wire f_u_arrmul24_fa17_23_y2;
  wire f_u_arrmul24_fa17_23_y3;
  wire f_u_arrmul24_fa17_23_y4;
  wire f_u_arrmul24_and18_23_a_18;
  wire f_u_arrmul24_and18_23_b_23;
  wire f_u_arrmul24_and18_23_y0;
  wire f_u_arrmul24_fa18_23_f_u_arrmul24_and18_23_y0;
  wire f_u_arrmul24_fa18_23_f_u_arrmul24_fa19_22_y2;
  wire f_u_arrmul24_fa18_23_y0;
  wire f_u_arrmul24_fa18_23_y1;
  wire f_u_arrmul24_fa18_23_f_u_arrmul24_fa17_23_y4;
  wire f_u_arrmul24_fa18_23_y2;
  wire f_u_arrmul24_fa18_23_y3;
  wire f_u_arrmul24_fa18_23_y4;
  wire f_u_arrmul24_and19_23_a_19;
  wire f_u_arrmul24_and19_23_b_23;
  wire f_u_arrmul24_and19_23_y0;
  wire f_u_arrmul24_fa19_23_f_u_arrmul24_and19_23_y0;
  wire f_u_arrmul24_fa19_23_f_u_arrmul24_fa20_22_y2;
  wire f_u_arrmul24_fa19_23_y0;
  wire f_u_arrmul24_fa19_23_y1;
  wire f_u_arrmul24_fa19_23_f_u_arrmul24_fa18_23_y4;
  wire f_u_arrmul24_fa19_23_y2;
  wire f_u_arrmul24_fa19_23_y3;
  wire f_u_arrmul24_fa19_23_y4;
  wire f_u_arrmul24_and20_23_a_20;
  wire f_u_arrmul24_and20_23_b_23;
  wire f_u_arrmul24_and20_23_y0;
  wire f_u_arrmul24_fa20_23_f_u_arrmul24_and20_23_y0;
  wire f_u_arrmul24_fa20_23_f_u_arrmul24_fa21_22_y2;
  wire f_u_arrmul24_fa20_23_y0;
  wire f_u_arrmul24_fa20_23_y1;
  wire f_u_arrmul24_fa20_23_f_u_arrmul24_fa19_23_y4;
  wire f_u_arrmul24_fa20_23_y2;
  wire f_u_arrmul24_fa20_23_y3;
  wire f_u_arrmul24_fa20_23_y4;
  wire f_u_arrmul24_and21_23_a_21;
  wire f_u_arrmul24_and21_23_b_23;
  wire f_u_arrmul24_and21_23_y0;
  wire f_u_arrmul24_fa21_23_f_u_arrmul24_and21_23_y0;
  wire f_u_arrmul24_fa21_23_f_u_arrmul24_fa22_22_y2;
  wire f_u_arrmul24_fa21_23_y0;
  wire f_u_arrmul24_fa21_23_y1;
  wire f_u_arrmul24_fa21_23_f_u_arrmul24_fa20_23_y4;
  wire f_u_arrmul24_fa21_23_y2;
  wire f_u_arrmul24_fa21_23_y3;
  wire f_u_arrmul24_fa21_23_y4;
  wire f_u_arrmul24_and22_23_a_22;
  wire f_u_arrmul24_and22_23_b_23;
  wire f_u_arrmul24_and22_23_y0;
  wire f_u_arrmul24_fa22_23_f_u_arrmul24_and22_23_y0;
  wire f_u_arrmul24_fa22_23_f_u_arrmul24_fa23_22_y2;
  wire f_u_arrmul24_fa22_23_y0;
  wire f_u_arrmul24_fa22_23_y1;
  wire f_u_arrmul24_fa22_23_f_u_arrmul24_fa21_23_y4;
  wire f_u_arrmul24_fa22_23_y2;
  wire f_u_arrmul24_fa22_23_y3;
  wire f_u_arrmul24_fa22_23_y4;
  wire f_u_arrmul24_and23_23_a_23;
  wire f_u_arrmul24_and23_23_b_23;
  wire f_u_arrmul24_and23_23_y0;
  wire f_u_arrmul24_fa23_23_f_u_arrmul24_and23_23_y0;
  wire f_u_arrmul24_fa23_23_f_u_arrmul24_fa23_22_y4;
  wire f_u_arrmul24_fa23_23_y0;
  wire f_u_arrmul24_fa23_23_y1;
  wire f_u_arrmul24_fa23_23_f_u_arrmul24_fa22_23_y4;
  wire f_u_arrmul24_fa23_23_y2;
  wire f_u_arrmul24_fa23_23_y3;
  wire f_u_arrmul24_fa23_23_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign f_u_arrmul24_and0_0_a_0 = a_0;
  assign f_u_arrmul24_and0_0_b_0 = b_0;
  assign f_u_arrmul24_and0_0_y0 = f_u_arrmul24_and0_0_a_0 & f_u_arrmul24_and0_0_b_0;
  assign f_u_arrmul24_and1_0_a_1 = a_1;
  assign f_u_arrmul24_and1_0_b_0 = b_0;
  assign f_u_arrmul24_and1_0_y0 = f_u_arrmul24_and1_0_a_1 & f_u_arrmul24_and1_0_b_0;
  assign f_u_arrmul24_and2_0_a_2 = a_2;
  assign f_u_arrmul24_and2_0_b_0 = b_0;
  assign f_u_arrmul24_and2_0_y0 = f_u_arrmul24_and2_0_a_2 & f_u_arrmul24_and2_0_b_0;
  assign f_u_arrmul24_and3_0_a_3 = a_3;
  assign f_u_arrmul24_and3_0_b_0 = b_0;
  assign f_u_arrmul24_and3_0_y0 = f_u_arrmul24_and3_0_a_3 & f_u_arrmul24_and3_0_b_0;
  assign f_u_arrmul24_and4_0_a_4 = a_4;
  assign f_u_arrmul24_and4_0_b_0 = b_0;
  assign f_u_arrmul24_and4_0_y0 = f_u_arrmul24_and4_0_a_4 & f_u_arrmul24_and4_0_b_0;
  assign f_u_arrmul24_and5_0_a_5 = a_5;
  assign f_u_arrmul24_and5_0_b_0 = b_0;
  assign f_u_arrmul24_and5_0_y0 = f_u_arrmul24_and5_0_a_5 & f_u_arrmul24_and5_0_b_0;
  assign f_u_arrmul24_and6_0_a_6 = a_6;
  assign f_u_arrmul24_and6_0_b_0 = b_0;
  assign f_u_arrmul24_and6_0_y0 = f_u_arrmul24_and6_0_a_6 & f_u_arrmul24_and6_0_b_0;
  assign f_u_arrmul24_and7_0_a_7 = a_7;
  assign f_u_arrmul24_and7_0_b_0 = b_0;
  assign f_u_arrmul24_and7_0_y0 = f_u_arrmul24_and7_0_a_7 & f_u_arrmul24_and7_0_b_0;
  assign f_u_arrmul24_and8_0_a_8 = a_8;
  assign f_u_arrmul24_and8_0_b_0 = b_0;
  assign f_u_arrmul24_and8_0_y0 = f_u_arrmul24_and8_0_a_8 & f_u_arrmul24_and8_0_b_0;
  assign f_u_arrmul24_and9_0_a_9 = a_9;
  assign f_u_arrmul24_and9_0_b_0 = b_0;
  assign f_u_arrmul24_and9_0_y0 = f_u_arrmul24_and9_0_a_9 & f_u_arrmul24_and9_0_b_0;
  assign f_u_arrmul24_and10_0_a_10 = a_10;
  assign f_u_arrmul24_and10_0_b_0 = b_0;
  assign f_u_arrmul24_and10_0_y0 = f_u_arrmul24_and10_0_a_10 & f_u_arrmul24_and10_0_b_0;
  assign f_u_arrmul24_and11_0_a_11 = a_11;
  assign f_u_arrmul24_and11_0_b_0 = b_0;
  assign f_u_arrmul24_and11_0_y0 = f_u_arrmul24_and11_0_a_11 & f_u_arrmul24_and11_0_b_0;
  assign f_u_arrmul24_and12_0_a_12 = a_12;
  assign f_u_arrmul24_and12_0_b_0 = b_0;
  assign f_u_arrmul24_and12_0_y0 = f_u_arrmul24_and12_0_a_12 & f_u_arrmul24_and12_0_b_0;
  assign f_u_arrmul24_and13_0_a_13 = a_13;
  assign f_u_arrmul24_and13_0_b_0 = b_0;
  assign f_u_arrmul24_and13_0_y0 = f_u_arrmul24_and13_0_a_13 & f_u_arrmul24_and13_0_b_0;
  assign f_u_arrmul24_and14_0_a_14 = a_14;
  assign f_u_arrmul24_and14_0_b_0 = b_0;
  assign f_u_arrmul24_and14_0_y0 = f_u_arrmul24_and14_0_a_14 & f_u_arrmul24_and14_0_b_0;
  assign f_u_arrmul24_and15_0_a_15 = a_15;
  assign f_u_arrmul24_and15_0_b_0 = b_0;
  assign f_u_arrmul24_and15_0_y0 = f_u_arrmul24_and15_0_a_15 & f_u_arrmul24_and15_0_b_0;
  assign f_u_arrmul24_and16_0_a_16 = a_16;
  assign f_u_arrmul24_and16_0_b_0 = b_0;
  assign f_u_arrmul24_and16_0_y0 = f_u_arrmul24_and16_0_a_16 & f_u_arrmul24_and16_0_b_0;
  assign f_u_arrmul24_and17_0_a_17 = a_17;
  assign f_u_arrmul24_and17_0_b_0 = b_0;
  assign f_u_arrmul24_and17_0_y0 = f_u_arrmul24_and17_0_a_17 & f_u_arrmul24_and17_0_b_0;
  assign f_u_arrmul24_and18_0_a_18 = a_18;
  assign f_u_arrmul24_and18_0_b_0 = b_0;
  assign f_u_arrmul24_and18_0_y0 = f_u_arrmul24_and18_0_a_18 & f_u_arrmul24_and18_0_b_0;
  assign f_u_arrmul24_and19_0_a_19 = a_19;
  assign f_u_arrmul24_and19_0_b_0 = b_0;
  assign f_u_arrmul24_and19_0_y0 = f_u_arrmul24_and19_0_a_19 & f_u_arrmul24_and19_0_b_0;
  assign f_u_arrmul24_and20_0_a_20 = a_20;
  assign f_u_arrmul24_and20_0_b_0 = b_0;
  assign f_u_arrmul24_and20_0_y0 = f_u_arrmul24_and20_0_a_20 & f_u_arrmul24_and20_0_b_0;
  assign f_u_arrmul24_and21_0_a_21 = a_21;
  assign f_u_arrmul24_and21_0_b_0 = b_0;
  assign f_u_arrmul24_and21_0_y0 = f_u_arrmul24_and21_0_a_21 & f_u_arrmul24_and21_0_b_0;
  assign f_u_arrmul24_and22_0_a_22 = a_22;
  assign f_u_arrmul24_and22_0_b_0 = b_0;
  assign f_u_arrmul24_and22_0_y0 = f_u_arrmul24_and22_0_a_22 & f_u_arrmul24_and22_0_b_0;
  assign f_u_arrmul24_and23_0_a_23 = a_23;
  assign f_u_arrmul24_and23_0_b_0 = b_0;
  assign f_u_arrmul24_and23_0_y0 = f_u_arrmul24_and23_0_a_23 & f_u_arrmul24_and23_0_b_0;
  assign f_u_arrmul24_and0_1_a_0 = a_0;
  assign f_u_arrmul24_and0_1_b_1 = b_1;
  assign f_u_arrmul24_and0_1_y0 = f_u_arrmul24_and0_1_a_0 & f_u_arrmul24_and0_1_b_1;
  assign f_u_arrmul24_ha0_1_f_u_arrmul24_and0_1_y0 = f_u_arrmul24_and0_1_y0;
  assign f_u_arrmul24_ha0_1_f_u_arrmul24_and1_0_y0 = f_u_arrmul24_and1_0_y0;
  assign f_u_arrmul24_ha0_1_y0 = f_u_arrmul24_ha0_1_f_u_arrmul24_and0_1_y0 ^ f_u_arrmul24_ha0_1_f_u_arrmul24_and1_0_y0;
  assign f_u_arrmul24_ha0_1_y1 = f_u_arrmul24_ha0_1_f_u_arrmul24_and0_1_y0 & f_u_arrmul24_ha0_1_f_u_arrmul24_and1_0_y0;
  assign f_u_arrmul24_and1_1_a_1 = a_1;
  assign f_u_arrmul24_and1_1_b_1 = b_1;
  assign f_u_arrmul24_and1_1_y0 = f_u_arrmul24_and1_1_a_1 & f_u_arrmul24_and1_1_b_1;
  assign f_u_arrmul24_fa1_1_f_u_arrmul24_and1_1_y0 = f_u_arrmul24_and1_1_y0;
  assign f_u_arrmul24_fa1_1_f_u_arrmul24_and2_0_y0 = f_u_arrmul24_and2_0_y0;
  assign f_u_arrmul24_fa1_1_f_u_arrmul24_ha0_1_y1 = f_u_arrmul24_ha0_1_y1;
  assign f_u_arrmul24_fa1_1_y0 = f_u_arrmul24_fa1_1_f_u_arrmul24_and1_1_y0 ^ f_u_arrmul24_fa1_1_f_u_arrmul24_and2_0_y0;
  assign f_u_arrmul24_fa1_1_y1 = f_u_arrmul24_fa1_1_f_u_arrmul24_and1_1_y0 & f_u_arrmul24_fa1_1_f_u_arrmul24_and2_0_y0;
  assign f_u_arrmul24_fa1_1_y2 = f_u_arrmul24_fa1_1_y0 ^ f_u_arrmul24_fa1_1_f_u_arrmul24_ha0_1_y1;
  assign f_u_arrmul24_fa1_1_y3 = f_u_arrmul24_fa1_1_y0 & f_u_arrmul24_fa1_1_f_u_arrmul24_ha0_1_y1;
  assign f_u_arrmul24_fa1_1_y4 = f_u_arrmul24_fa1_1_y1 | f_u_arrmul24_fa1_1_y3;
  assign f_u_arrmul24_and2_1_a_2 = a_2;
  assign f_u_arrmul24_and2_1_b_1 = b_1;
  assign f_u_arrmul24_and2_1_y0 = f_u_arrmul24_and2_1_a_2 & f_u_arrmul24_and2_1_b_1;
  assign f_u_arrmul24_fa2_1_f_u_arrmul24_and2_1_y0 = f_u_arrmul24_and2_1_y0;
  assign f_u_arrmul24_fa2_1_f_u_arrmul24_and3_0_y0 = f_u_arrmul24_and3_0_y0;
  assign f_u_arrmul24_fa2_1_f_u_arrmul24_fa1_1_y4 = f_u_arrmul24_fa1_1_y4;
  assign f_u_arrmul24_fa2_1_y0 = f_u_arrmul24_fa2_1_f_u_arrmul24_and2_1_y0 ^ f_u_arrmul24_fa2_1_f_u_arrmul24_and3_0_y0;
  assign f_u_arrmul24_fa2_1_y1 = f_u_arrmul24_fa2_1_f_u_arrmul24_and2_1_y0 & f_u_arrmul24_fa2_1_f_u_arrmul24_and3_0_y0;
  assign f_u_arrmul24_fa2_1_y2 = f_u_arrmul24_fa2_1_y0 ^ f_u_arrmul24_fa2_1_f_u_arrmul24_fa1_1_y4;
  assign f_u_arrmul24_fa2_1_y3 = f_u_arrmul24_fa2_1_y0 & f_u_arrmul24_fa2_1_f_u_arrmul24_fa1_1_y4;
  assign f_u_arrmul24_fa2_1_y4 = f_u_arrmul24_fa2_1_y1 | f_u_arrmul24_fa2_1_y3;
  assign f_u_arrmul24_and3_1_a_3 = a_3;
  assign f_u_arrmul24_and3_1_b_1 = b_1;
  assign f_u_arrmul24_and3_1_y0 = f_u_arrmul24_and3_1_a_3 & f_u_arrmul24_and3_1_b_1;
  assign f_u_arrmul24_fa3_1_f_u_arrmul24_and3_1_y0 = f_u_arrmul24_and3_1_y0;
  assign f_u_arrmul24_fa3_1_f_u_arrmul24_and4_0_y0 = f_u_arrmul24_and4_0_y0;
  assign f_u_arrmul24_fa3_1_f_u_arrmul24_fa2_1_y4 = f_u_arrmul24_fa2_1_y4;
  assign f_u_arrmul24_fa3_1_y0 = f_u_arrmul24_fa3_1_f_u_arrmul24_and3_1_y0 ^ f_u_arrmul24_fa3_1_f_u_arrmul24_and4_0_y0;
  assign f_u_arrmul24_fa3_1_y1 = f_u_arrmul24_fa3_1_f_u_arrmul24_and3_1_y0 & f_u_arrmul24_fa3_1_f_u_arrmul24_and4_0_y0;
  assign f_u_arrmul24_fa3_1_y2 = f_u_arrmul24_fa3_1_y0 ^ f_u_arrmul24_fa3_1_f_u_arrmul24_fa2_1_y4;
  assign f_u_arrmul24_fa3_1_y3 = f_u_arrmul24_fa3_1_y0 & f_u_arrmul24_fa3_1_f_u_arrmul24_fa2_1_y4;
  assign f_u_arrmul24_fa3_1_y4 = f_u_arrmul24_fa3_1_y1 | f_u_arrmul24_fa3_1_y3;
  assign f_u_arrmul24_and4_1_a_4 = a_4;
  assign f_u_arrmul24_and4_1_b_1 = b_1;
  assign f_u_arrmul24_and4_1_y0 = f_u_arrmul24_and4_1_a_4 & f_u_arrmul24_and4_1_b_1;
  assign f_u_arrmul24_fa4_1_f_u_arrmul24_and4_1_y0 = f_u_arrmul24_and4_1_y0;
  assign f_u_arrmul24_fa4_1_f_u_arrmul24_and5_0_y0 = f_u_arrmul24_and5_0_y0;
  assign f_u_arrmul24_fa4_1_f_u_arrmul24_fa3_1_y4 = f_u_arrmul24_fa3_1_y4;
  assign f_u_arrmul24_fa4_1_y0 = f_u_arrmul24_fa4_1_f_u_arrmul24_and4_1_y0 ^ f_u_arrmul24_fa4_1_f_u_arrmul24_and5_0_y0;
  assign f_u_arrmul24_fa4_1_y1 = f_u_arrmul24_fa4_1_f_u_arrmul24_and4_1_y0 & f_u_arrmul24_fa4_1_f_u_arrmul24_and5_0_y0;
  assign f_u_arrmul24_fa4_1_y2 = f_u_arrmul24_fa4_1_y0 ^ f_u_arrmul24_fa4_1_f_u_arrmul24_fa3_1_y4;
  assign f_u_arrmul24_fa4_1_y3 = f_u_arrmul24_fa4_1_y0 & f_u_arrmul24_fa4_1_f_u_arrmul24_fa3_1_y4;
  assign f_u_arrmul24_fa4_1_y4 = f_u_arrmul24_fa4_1_y1 | f_u_arrmul24_fa4_1_y3;
  assign f_u_arrmul24_and5_1_a_5 = a_5;
  assign f_u_arrmul24_and5_1_b_1 = b_1;
  assign f_u_arrmul24_and5_1_y0 = f_u_arrmul24_and5_1_a_5 & f_u_arrmul24_and5_1_b_1;
  assign f_u_arrmul24_fa5_1_f_u_arrmul24_and5_1_y0 = f_u_arrmul24_and5_1_y0;
  assign f_u_arrmul24_fa5_1_f_u_arrmul24_and6_0_y0 = f_u_arrmul24_and6_0_y0;
  assign f_u_arrmul24_fa5_1_f_u_arrmul24_fa4_1_y4 = f_u_arrmul24_fa4_1_y4;
  assign f_u_arrmul24_fa5_1_y0 = f_u_arrmul24_fa5_1_f_u_arrmul24_and5_1_y0 ^ f_u_arrmul24_fa5_1_f_u_arrmul24_and6_0_y0;
  assign f_u_arrmul24_fa5_1_y1 = f_u_arrmul24_fa5_1_f_u_arrmul24_and5_1_y0 & f_u_arrmul24_fa5_1_f_u_arrmul24_and6_0_y0;
  assign f_u_arrmul24_fa5_1_y2 = f_u_arrmul24_fa5_1_y0 ^ f_u_arrmul24_fa5_1_f_u_arrmul24_fa4_1_y4;
  assign f_u_arrmul24_fa5_1_y3 = f_u_arrmul24_fa5_1_y0 & f_u_arrmul24_fa5_1_f_u_arrmul24_fa4_1_y4;
  assign f_u_arrmul24_fa5_1_y4 = f_u_arrmul24_fa5_1_y1 | f_u_arrmul24_fa5_1_y3;
  assign f_u_arrmul24_and6_1_a_6 = a_6;
  assign f_u_arrmul24_and6_1_b_1 = b_1;
  assign f_u_arrmul24_and6_1_y0 = f_u_arrmul24_and6_1_a_6 & f_u_arrmul24_and6_1_b_1;
  assign f_u_arrmul24_fa6_1_f_u_arrmul24_and6_1_y0 = f_u_arrmul24_and6_1_y0;
  assign f_u_arrmul24_fa6_1_f_u_arrmul24_and7_0_y0 = f_u_arrmul24_and7_0_y0;
  assign f_u_arrmul24_fa6_1_f_u_arrmul24_fa5_1_y4 = f_u_arrmul24_fa5_1_y4;
  assign f_u_arrmul24_fa6_1_y0 = f_u_arrmul24_fa6_1_f_u_arrmul24_and6_1_y0 ^ f_u_arrmul24_fa6_1_f_u_arrmul24_and7_0_y0;
  assign f_u_arrmul24_fa6_1_y1 = f_u_arrmul24_fa6_1_f_u_arrmul24_and6_1_y0 & f_u_arrmul24_fa6_1_f_u_arrmul24_and7_0_y0;
  assign f_u_arrmul24_fa6_1_y2 = f_u_arrmul24_fa6_1_y0 ^ f_u_arrmul24_fa6_1_f_u_arrmul24_fa5_1_y4;
  assign f_u_arrmul24_fa6_1_y3 = f_u_arrmul24_fa6_1_y0 & f_u_arrmul24_fa6_1_f_u_arrmul24_fa5_1_y4;
  assign f_u_arrmul24_fa6_1_y4 = f_u_arrmul24_fa6_1_y1 | f_u_arrmul24_fa6_1_y3;
  assign f_u_arrmul24_and7_1_a_7 = a_7;
  assign f_u_arrmul24_and7_1_b_1 = b_1;
  assign f_u_arrmul24_and7_1_y0 = f_u_arrmul24_and7_1_a_7 & f_u_arrmul24_and7_1_b_1;
  assign f_u_arrmul24_fa7_1_f_u_arrmul24_and7_1_y0 = f_u_arrmul24_and7_1_y0;
  assign f_u_arrmul24_fa7_1_f_u_arrmul24_and8_0_y0 = f_u_arrmul24_and8_0_y0;
  assign f_u_arrmul24_fa7_1_f_u_arrmul24_fa6_1_y4 = f_u_arrmul24_fa6_1_y4;
  assign f_u_arrmul24_fa7_1_y0 = f_u_arrmul24_fa7_1_f_u_arrmul24_and7_1_y0 ^ f_u_arrmul24_fa7_1_f_u_arrmul24_and8_0_y0;
  assign f_u_arrmul24_fa7_1_y1 = f_u_arrmul24_fa7_1_f_u_arrmul24_and7_1_y0 & f_u_arrmul24_fa7_1_f_u_arrmul24_and8_0_y0;
  assign f_u_arrmul24_fa7_1_y2 = f_u_arrmul24_fa7_1_y0 ^ f_u_arrmul24_fa7_1_f_u_arrmul24_fa6_1_y4;
  assign f_u_arrmul24_fa7_1_y3 = f_u_arrmul24_fa7_1_y0 & f_u_arrmul24_fa7_1_f_u_arrmul24_fa6_1_y4;
  assign f_u_arrmul24_fa7_1_y4 = f_u_arrmul24_fa7_1_y1 | f_u_arrmul24_fa7_1_y3;
  assign f_u_arrmul24_and8_1_a_8 = a_8;
  assign f_u_arrmul24_and8_1_b_1 = b_1;
  assign f_u_arrmul24_and8_1_y0 = f_u_arrmul24_and8_1_a_8 & f_u_arrmul24_and8_1_b_1;
  assign f_u_arrmul24_fa8_1_f_u_arrmul24_and8_1_y0 = f_u_arrmul24_and8_1_y0;
  assign f_u_arrmul24_fa8_1_f_u_arrmul24_and9_0_y0 = f_u_arrmul24_and9_0_y0;
  assign f_u_arrmul24_fa8_1_f_u_arrmul24_fa7_1_y4 = f_u_arrmul24_fa7_1_y4;
  assign f_u_arrmul24_fa8_1_y0 = f_u_arrmul24_fa8_1_f_u_arrmul24_and8_1_y0 ^ f_u_arrmul24_fa8_1_f_u_arrmul24_and9_0_y0;
  assign f_u_arrmul24_fa8_1_y1 = f_u_arrmul24_fa8_1_f_u_arrmul24_and8_1_y0 & f_u_arrmul24_fa8_1_f_u_arrmul24_and9_0_y0;
  assign f_u_arrmul24_fa8_1_y2 = f_u_arrmul24_fa8_1_y0 ^ f_u_arrmul24_fa8_1_f_u_arrmul24_fa7_1_y4;
  assign f_u_arrmul24_fa8_1_y3 = f_u_arrmul24_fa8_1_y0 & f_u_arrmul24_fa8_1_f_u_arrmul24_fa7_1_y4;
  assign f_u_arrmul24_fa8_1_y4 = f_u_arrmul24_fa8_1_y1 | f_u_arrmul24_fa8_1_y3;
  assign f_u_arrmul24_and9_1_a_9 = a_9;
  assign f_u_arrmul24_and9_1_b_1 = b_1;
  assign f_u_arrmul24_and9_1_y0 = f_u_arrmul24_and9_1_a_9 & f_u_arrmul24_and9_1_b_1;
  assign f_u_arrmul24_fa9_1_f_u_arrmul24_and9_1_y0 = f_u_arrmul24_and9_1_y0;
  assign f_u_arrmul24_fa9_1_f_u_arrmul24_and10_0_y0 = f_u_arrmul24_and10_0_y0;
  assign f_u_arrmul24_fa9_1_f_u_arrmul24_fa8_1_y4 = f_u_arrmul24_fa8_1_y4;
  assign f_u_arrmul24_fa9_1_y0 = f_u_arrmul24_fa9_1_f_u_arrmul24_and9_1_y0 ^ f_u_arrmul24_fa9_1_f_u_arrmul24_and10_0_y0;
  assign f_u_arrmul24_fa9_1_y1 = f_u_arrmul24_fa9_1_f_u_arrmul24_and9_1_y0 & f_u_arrmul24_fa9_1_f_u_arrmul24_and10_0_y0;
  assign f_u_arrmul24_fa9_1_y2 = f_u_arrmul24_fa9_1_y0 ^ f_u_arrmul24_fa9_1_f_u_arrmul24_fa8_1_y4;
  assign f_u_arrmul24_fa9_1_y3 = f_u_arrmul24_fa9_1_y0 & f_u_arrmul24_fa9_1_f_u_arrmul24_fa8_1_y4;
  assign f_u_arrmul24_fa9_1_y4 = f_u_arrmul24_fa9_1_y1 | f_u_arrmul24_fa9_1_y3;
  assign f_u_arrmul24_and10_1_a_10 = a_10;
  assign f_u_arrmul24_and10_1_b_1 = b_1;
  assign f_u_arrmul24_and10_1_y0 = f_u_arrmul24_and10_1_a_10 & f_u_arrmul24_and10_1_b_1;
  assign f_u_arrmul24_fa10_1_f_u_arrmul24_and10_1_y0 = f_u_arrmul24_and10_1_y0;
  assign f_u_arrmul24_fa10_1_f_u_arrmul24_and11_0_y0 = f_u_arrmul24_and11_0_y0;
  assign f_u_arrmul24_fa10_1_f_u_arrmul24_fa9_1_y4 = f_u_arrmul24_fa9_1_y4;
  assign f_u_arrmul24_fa10_1_y0 = f_u_arrmul24_fa10_1_f_u_arrmul24_and10_1_y0 ^ f_u_arrmul24_fa10_1_f_u_arrmul24_and11_0_y0;
  assign f_u_arrmul24_fa10_1_y1 = f_u_arrmul24_fa10_1_f_u_arrmul24_and10_1_y0 & f_u_arrmul24_fa10_1_f_u_arrmul24_and11_0_y0;
  assign f_u_arrmul24_fa10_1_y2 = f_u_arrmul24_fa10_1_y0 ^ f_u_arrmul24_fa10_1_f_u_arrmul24_fa9_1_y4;
  assign f_u_arrmul24_fa10_1_y3 = f_u_arrmul24_fa10_1_y0 & f_u_arrmul24_fa10_1_f_u_arrmul24_fa9_1_y4;
  assign f_u_arrmul24_fa10_1_y4 = f_u_arrmul24_fa10_1_y1 | f_u_arrmul24_fa10_1_y3;
  assign f_u_arrmul24_and11_1_a_11 = a_11;
  assign f_u_arrmul24_and11_1_b_1 = b_1;
  assign f_u_arrmul24_and11_1_y0 = f_u_arrmul24_and11_1_a_11 & f_u_arrmul24_and11_1_b_1;
  assign f_u_arrmul24_fa11_1_f_u_arrmul24_and11_1_y0 = f_u_arrmul24_and11_1_y0;
  assign f_u_arrmul24_fa11_1_f_u_arrmul24_and12_0_y0 = f_u_arrmul24_and12_0_y0;
  assign f_u_arrmul24_fa11_1_f_u_arrmul24_fa10_1_y4 = f_u_arrmul24_fa10_1_y4;
  assign f_u_arrmul24_fa11_1_y0 = f_u_arrmul24_fa11_1_f_u_arrmul24_and11_1_y0 ^ f_u_arrmul24_fa11_1_f_u_arrmul24_and12_0_y0;
  assign f_u_arrmul24_fa11_1_y1 = f_u_arrmul24_fa11_1_f_u_arrmul24_and11_1_y0 & f_u_arrmul24_fa11_1_f_u_arrmul24_and12_0_y0;
  assign f_u_arrmul24_fa11_1_y2 = f_u_arrmul24_fa11_1_y0 ^ f_u_arrmul24_fa11_1_f_u_arrmul24_fa10_1_y4;
  assign f_u_arrmul24_fa11_1_y3 = f_u_arrmul24_fa11_1_y0 & f_u_arrmul24_fa11_1_f_u_arrmul24_fa10_1_y4;
  assign f_u_arrmul24_fa11_1_y4 = f_u_arrmul24_fa11_1_y1 | f_u_arrmul24_fa11_1_y3;
  assign f_u_arrmul24_and12_1_a_12 = a_12;
  assign f_u_arrmul24_and12_1_b_1 = b_1;
  assign f_u_arrmul24_and12_1_y0 = f_u_arrmul24_and12_1_a_12 & f_u_arrmul24_and12_1_b_1;
  assign f_u_arrmul24_fa12_1_f_u_arrmul24_and12_1_y0 = f_u_arrmul24_and12_1_y0;
  assign f_u_arrmul24_fa12_1_f_u_arrmul24_and13_0_y0 = f_u_arrmul24_and13_0_y0;
  assign f_u_arrmul24_fa12_1_f_u_arrmul24_fa11_1_y4 = f_u_arrmul24_fa11_1_y4;
  assign f_u_arrmul24_fa12_1_y0 = f_u_arrmul24_fa12_1_f_u_arrmul24_and12_1_y0 ^ f_u_arrmul24_fa12_1_f_u_arrmul24_and13_0_y0;
  assign f_u_arrmul24_fa12_1_y1 = f_u_arrmul24_fa12_1_f_u_arrmul24_and12_1_y0 & f_u_arrmul24_fa12_1_f_u_arrmul24_and13_0_y0;
  assign f_u_arrmul24_fa12_1_y2 = f_u_arrmul24_fa12_1_y0 ^ f_u_arrmul24_fa12_1_f_u_arrmul24_fa11_1_y4;
  assign f_u_arrmul24_fa12_1_y3 = f_u_arrmul24_fa12_1_y0 & f_u_arrmul24_fa12_1_f_u_arrmul24_fa11_1_y4;
  assign f_u_arrmul24_fa12_1_y4 = f_u_arrmul24_fa12_1_y1 | f_u_arrmul24_fa12_1_y3;
  assign f_u_arrmul24_and13_1_a_13 = a_13;
  assign f_u_arrmul24_and13_1_b_1 = b_1;
  assign f_u_arrmul24_and13_1_y0 = f_u_arrmul24_and13_1_a_13 & f_u_arrmul24_and13_1_b_1;
  assign f_u_arrmul24_fa13_1_f_u_arrmul24_and13_1_y0 = f_u_arrmul24_and13_1_y0;
  assign f_u_arrmul24_fa13_1_f_u_arrmul24_and14_0_y0 = f_u_arrmul24_and14_0_y0;
  assign f_u_arrmul24_fa13_1_f_u_arrmul24_fa12_1_y4 = f_u_arrmul24_fa12_1_y4;
  assign f_u_arrmul24_fa13_1_y0 = f_u_arrmul24_fa13_1_f_u_arrmul24_and13_1_y0 ^ f_u_arrmul24_fa13_1_f_u_arrmul24_and14_0_y0;
  assign f_u_arrmul24_fa13_1_y1 = f_u_arrmul24_fa13_1_f_u_arrmul24_and13_1_y0 & f_u_arrmul24_fa13_1_f_u_arrmul24_and14_0_y0;
  assign f_u_arrmul24_fa13_1_y2 = f_u_arrmul24_fa13_1_y0 ^ f_u_arrmul24_fa13_1_f_u_arrmul24_fa12_1_y4;
  assign f_u_arrmul24_fa13_1_y3 = f_u_arrmul24_fa13_1_y0 & f_u_arrmul24_fa13_1_f_u_arrmul24_fa12_1_y4;
  assign f_u_arrmul24_fa13_1_y4 = f_u_arrmul24_fa13_1_y1 | f_u_arrmul24_fa13_1_y3;
  assign f_u_arrmul24_and14_1_a_14 = a_14;
  assign f_u_arrmul24_and14_1_b_1 = b_1;
  assign f_u_arrmul24_and14_1_y0 = f_u_arrmul24_and14_1_a_14 & f_u_arrmul24_and14_1_b_1;
  assign f_u_arrmul24_fa14_1_f_u_arrmul24_and14_1_y0 = f_u_arrmul24_and14_1_y0;
  assign f_u_arrmul24_fa14_1_f_u_arrmul24_and15_0_y0 = f_u_arrmul24_and15_0_y0;
  assign f_u_arrmul24_fa14_1_f_u_arrmul24_fa13_1_y4 = f_u_arrmul24_fa13_1_y4;
  assign f_u_arrmul24_fa14_1_y0 = f_u_arrmul24_fa14_1_f_u_arrmul24_and14_1_y0 ^ f_u_arrmul24_fa14_1_f_u_arrmul24_and15_0_y0;
  assign f_u_arrmul24_fa14_1_y1 = f_u_arrmul24_fa14_1_f_u_arrmul24_and14_1_y0 & f_u_arrmul24_fa14_1_f_u_arrmul24_and15_0_y0;
  assign f_u_arrmul24_fa14_1_y2 = f_u_arrmul24_fa14_1_y0 ^ f_u_arrmul24_fa14_1_f_u_arrmul24_fa13_1_y4;
  assign f_u_arrmul24_fa14_1_y3 = f_u_arrmul24_fa14_1_y0 & f_u_arrmul24_fa14_1_f_u_arrmul24_fa13_1_y4;
  assign f_u_arrmul24_fa14_1_y4 = f_u_arrmul24_fa14_1_y1 | f_u_arrmul24_fa14_1_y3;
  assign f_u_arrmul24_and15_1_a_15 = a_15;
  assign f_u_arrmul24_and15_1_b_1 = b_1;
  assign f_u_arrmul24_and15_1_y0 = f_u_arrmul24_and15_1_a_15 & f_u_arrmul24_and15_1_b_1;
  assign f_u_arrmul24_fa15_1_f_u_arrmul24_and15_1_y0 = f_u_arrmul24_and15_1_y0;
  assign f_u_arrmul24_fa15_1_f_u_arrmul24_and16_0_y0 = f_u_arrmul24_and16_0_y0;
  assign f_u_arrmul24_fa15_1_f_u_arrmul24_fa14_1_y4 = f_u_arrmul24_fa14_1_y4;
  assign f_u_arrmul24_fa15_1_y0 = f_u_arrmul24_fa15_1_f_u_arrmul24_and15_1_y0 ^ f_u_arrmul24_fa15_1_f_u_arrmul24_and16_0_y0;
  assign f_u_arrmul24_fa15_1_y1 = f_u_arrmul24_fa15_1_f_u_arrmul24_and15_1_y0 & f_u_arrmul24_fa15_1_f_u_arrmul24_and16_0_y0;
  assign f_u_arrmul24_fa15_1_y2 = f_u_arrmul24_fa15_1_y0 ^ f_u_arrmul24_fa15_1_f_u_arrmul24_fa14_1_y4;
  assign f_u_arrmul24_fa15_1_y3 = f_u_arrmul24_fa15_1_y0 & f_u_arrmul24_fa15_1_f_u_arrmul24_fa14_1_y4;
  assign f_u_arrmul24_fa15_1_y4 = f_u_arrmul24_fa15_1_y1 | f_u_arrmul24_fa15_1_y3;
  assign f_u_arrmul24_and16_1_a_16 = a_16;
  assign f_u_arrmul24_and16_1_b_1 = b_1;
  assign f_u_arrmul24_and16_1_y0 = f_u_arrmul24_and16_1_a_16 & f_u_arrmul24_and16_1_b_1;
  assign f_u_arrmul24_fa16_1_f_u_arrmul24_and16_1_y0 = f_u_arrmul24_and16_1_y0;
  assign f_u_arrmul24_fa16_1_f_u_arrmul24_and17_0_y0 = f_u_arrmul24_and17_0_y0;
  assign f_u_arrmul24_fa16_1_f_u_arrmul24_fa15_1_y4 = f_u_arrmul24_fa15_1_y4;
  assign f_u_arrmul24_fa16_1_y0 = f_u_arrmul24_fa16_1_f_u_arrmul24_and16_1_y0 ^ f_u_arrmul24_fa16_1_f_u_arrmul24_and17_0_y0;
  assign f_u_arrmul24_fa16_1_y1 = f_u_arrmul24_fa16_1_f_u_arrmul24_and16_1_y0 & f_u_arrmul24_fa16_1_f_u_arrmul24_and17_0_y0;
  assign f_u_arrmul24_fa16_1_y2 = f_u_arrmul24_fa16_1_y0 ^ f_u_arrmul24_fa16_1_f_u_arrmul24_fa15_1_y4;
  assign f_u_arrmul24_fa16_1_y3 = f_u_arrmul24_fa16_1_y0 & f_u_arrmul24_fa16_1_f_u_arrmul24_fa15_1_y4;
  assign f_u_arrmul24_fa16_1_y4 = f_u_arrmul24_fa16_1_y1 | f_u_arrmul24_fa16_1_y3;
  assign f_u_arrmul24_and17_1_a_17 = a_17;
  assign f_u_arrmul24_and17_1_b_1 = b_1;
  assign f_u_arrmul24_and17_1_y0 = f_u_arrmul24_and17_1_a_17 & f_u_arrmul24_and17_1_b_1;
  assign f_u_arrmul24_fa17_1_f_u_arrmul24_and17_1_y0 = f_u_arrmul24_and17_1_y0;
  assign f_u_arrmul24_fa17_1_f_u_arrmul24_and18_0_y0 = f_u_arrmul24_and18_0_y0;
  assign f_u_arrmul24_fa17_1_f_u_arrmul24_fa16_1_y4 = f_u_arrmul24_fa16_1_y4;
  assign f_u_arrmul24_fa17_1_y0 = f_u_arrmul24_fa17_1_f_u_arrmul24_and17_1_y0 ^ f_u_arrmul24_fa17_1_f_u_arrmul24_and18_0_y0;
  assign f_u_arrmul24_fa17_1_y1 = f_u_arrmul24_fa17_1_f_u_arrmul24_and17_1_y0 & f_u_arrmul24_fa17_1_f_u_arrmul24_and18_0_y0;
  assign f_u_arrmul24_fa17_1_y2 = f_u_arrmul24_fa17_1_y0 ^ f_u_arrmul24_fa17_1_f_u_arrmul24_fa16_1_y4;
  assign f_u_arrmul24_fa17_1_y3 = f_u_arrmul24_fa17_1_y0 & f_u_arrmul24_fa17_1_f_u_arrmul24_fa16_1_y4;
  assign f_u_arrmul24_fa17_1_y4 = f_u_arrmul24_fa17_1_y1 | f_u_arrmul24_fa17_1_y3;
  assign f_u_arrmul24_and18_1_a_18 = a_18;
  assign f_u_arrmul24_and18_1_b_1 = b_1;
  assign f_u_arrmul24_and18_1_y0 = f_u_arrmul24_and18_1_a_18 & f_u_arrmul24_and18_1_b_1;
  assign f_u_arrmul24_fa18_1_f_u_arrmul24_and18_1_y0 = f_u_arrmul24_and18_1_y0;
  assign f_u_arrmul24_fa18_1_f_u_arrmul24_and19_0_y0 = f_u_arrmul24_and19_0_y0;
  assign f_u_arrmul24_fa18_1_f_u_arrmul24_fa17_1_y4 = f_u_arrmul24_fa17_1_y4;
  assign f_u_arrmul24_fa18_1_y0 = f_u_arrmul24_fa18_1_f_u_arrmul24_and18_1_y0 ^ f_u_arrmul24_fa18_1_f_u_arrmul24_and19_0_y0;
  assign f_u_arrmul24_fa18_1_y1 = f_u_arrmul24_fa18_1_f_u_arrmul24_and18_1_y0 & f_u_arrmul24_fa18_1_f_u_arrmul24_and19_0_y0;
  assign f_u_arrmul24_fa18_1_y2 = f_u_arrmul24_fa18_1_y0 ^ f_u_arrmul24_fa18_1_f_u_arrmul24_fa17_1_y4;
  assign f_u_arrmul24_fa18_1_y3 = f_u_arrmul24_fa18_1_y0 & f_u_arrmul24_fa18_1_f_u_arrmul24_fa17_1_y4;
  assign f_u_arrmul24_fa18_1_y4 = f_u_arrmul24_fa18_1_y1 | f_u_arrmul24_fa18_1_y3;
  assign f_u_arrmul24_and19_1_a_19 = a_19;
  assign f_u_arrmul24_and19_1_b_1 = b_1;
  assign f_u_arrmul24_and19_1_y0 = f_u_arrmul24_and19_1_a_19 & f_u_arrmul24_and19_1_b_1;
  assign f_u_arrmul24_fa19_1_f_u_arrmul24_and19_1_y0 = f_u_arrmul24_and19_1_y0;
  assign f_u_arrmul24_fa19_1_f_u_arrmul24_and20_0_y0 = f_u_arrmul24_and20_0_y0;
  assign f_u_arrmul24_fa19_1_f_u_arrmul24_fa18_1_y4 = f_u_arrmul24_fa18_1_y4;
  assign f_u_arrmul24_fa19_1_y0 = f_u_arrmul24_fa19_1_f_u_arrmul24_and19_1_y0 ^ f_u_arrmul24_fa19_1_f_u_arrmul24_and20_0_y0;
  assign f_u_arrmul24_fa19_1_y1 = f_u_arrmul24_fa19_1_f_u_arrmul24_and19_1_y0 & f_u_arrmul24_fa19_1_f_u_arrmul24_and20_0_y0;
  assign f_u_arrmul24_fa19_1_y2 = f_u_arrmul24_fa19_1_y0 ^ f_u_arrmul24_fa19_1_f_u_arrmul24_fa18_1_y4;
  assign f_u_arrmul24_fa19_1_y3 = f_u_arrmul24_fa19_1_y0 & f_u_arrmul24_fa19_1_f_u_arrmul24_fa18_1_y4;
  assign f_u_arrmul24_fa19_1_y4 = f_u_arrmul24_fa19_1_y1 | f_u_arrmul24_fa19_1_y3;
  assign f_u_arrmul24_and20_1_a_20 = a_20;
  assign f_u_arrmul24_and20_1_b_1 = b_1;
  assign f_u_arrmul24_and20_1_y0 = f_u_arrmul24_and20_1_a_20 & f_u_arrmul24_and20_1_b_1;
  assign f_u_arrmul24_fa20_1_f_u_arrmul24_and20_1_y0 = f_u_arrmul24_and20_1_y0;
  assign f_u_arrmul24_fa20_1_f_u_arrmul24_and21_0_y0 = f_u_arrmul24_and21_0_y0;
  assign f_u_arrmul24_fa20_1_f_u_arrmul24_fa19_1_y4 = f_u_arrmul24_fa19_1_y4;
  assign f_u_arrmul24_fa20_1_y0 = f_u_arrmul24_fa20_1_f_u_arrmul24_and20_1_y0 ^ f_u_arrmul24_fa20_1_f_u_arrmul24_and21_0_y0;
  assign f_u_arrmul24_fa20_1_y1 = f_u_arrmul24_fa20_1_f_u_arrmul24_and20_1_y0 & f_u_arrmul24_fa20_1_f_u_arrmul24_and21_0_y0;
  assign f_u_arrmul24_fa20_1_y2 = f_u_arrmul24_fa20_1_y0 ^ f_u_arrmul24_fa20_1_f_u_arrmul24_fa19_1_y4;
  assign f_u_arrmul24_fa20_1_y3 = f_u_arrmul24_fa20_1_y0 & f_u_arrmul24_fa20_1_f_u_arrmul24_fa19_1_y4;
  assign f_u_arrmul24_fa20_1_y4 = f_u_arrmul24_fa20_1_y1 | f_u_arrmul24_fa20_1_y3;
  assign f_u_arrmul24_and21_1_a_21 = a_21;
  assign f_u_arrmul24_and21_1_b_1 = b_1;
  assign f_u_arrmul24_and21_1_y0 = f_u_arrmul24_and21_1_a_21 & f_u_arrmul24_and21_1_b_1;
  assign f_u_arrmul24_fa21_1_f_u_arrmul24_and21_1_y0 = f_u_arrmul24_and21_1_y0;
  assign f_u_arrmul24_fa21_1_f_u_arrmul24_and22_0_y0 = f_u_arrmul24_and22_0_y0;
  assign f_u_arrmul24_fa21_1_f_u_arrmul24_fa20_1_y4 = f_u_arrmul24_fa20_1_y4;
  assign f_u_arrmul24_fa21_1_y0 = f_u_arrmul24_fa21_1_f_u_arrmul24_and21_1_y0 ^ f_u_arrmul24_fa21_1_f_u_arrmul24_and22_0_y0;
  assign f_u_arrmul24_fa21_1_y1 = f_u_arrmul24_fa21_1_f_u_arrmul24_and21_1_y0 & f_u_arrmul24_fa21_1_f_u_arrmul24_and22_0_y0;
  assign f_u_arrmul24_fa21_1_y2 = f_u_arrmul24_fa21_1_y0 ^ f_u_arrmul24_fa21_1_f_u_arrmul24_fa20_1_y4;
  assign f_u_arrmul24_fa21_1_y3 = f_u_arrmul24_fa21_1_y0 & f_u_arrmul24_fa21_1_f_u_arrmul24_fa20_1_y4;
  assign f_u_arrmul24_fa21_1_y4 = f_u_arrmul24_fa21_1_y1 | f_u_arrmul24_fa21_1_y3;
  assign f_u_arrmul24_and22_1_a_22 = a_22;
  assign f_u_arrmul24_and22_1_b_1 = b_1;
  assign f_u_arrmul24_and22_1_y0 = f_u_arrmul24_and22_1_a_22 & f_u_arrmul24_and22_1_b_1;
  assign f_u_arrmul24_fa22_1_f_u_arrmul24_and22_1_y0 = f_u_arrmul24_and22_1_y0;
  assign f_u_arrmul24_fa22_1_f_u_arrmul24_and23_0_y0 = f_u_arrmul24_and23_0_y0;
  assign f_u_arrmul24_fa22_1_f_u_arrmul24_fa21_1_y4 = f_u_arrmul24_fa21_1_y4;
  assign f_u_arrmul24_fa22_1_y0 = f_u_arrmul24_fa22_1_f_u_arrmul24_and22_1_y0 ^ f_u_arrmul24_fa22_1_f_u_arrmul24_and23_0_y0;
  assign f_u_arrmul24_fa22_1_y1 = f_u_arrmul24_fa22_1_f_u_arrmul24_and22_1_y0 & f_u_arrmul24_fa22_1_f_u_arrmul24_and23_0_y0;
  assign f_u_arrmul24_fa22_1_y2 = f_u_arrmul24_fa22_1_y0 ^ f_u_arrmul24_fa22_1_f_u_arrmul24_fa21_1_y4;
  assign f_u_arrmul24_fa22_1_y3 = f_u_arrmul24_fa22_1_y0 & f_u_arrmul24_fa22_1_f_u_arrmul24_fa21_1_y4;
  assign f_u_arrmul24_fa22_1_y4 = f_u_arrmul24_fa22_1_y1 | f_u_arrmul24_fa22_1_y3;
  assign f_u_arrmul24_and23_1_a_23 = a_23;
  assign f_u_arrmul24_and23_1_b_1 = b_1;
  assign f_u_arrmul24_and23_1_y0 = f_u_arrmul24_and23_1_a_23 & f_u_arrmul24_and23_1_b_1;
  assign f_u_arrmul24_ha23_1_f_u_arrmul24_and23_1_y0 = f_u_arrmul24_and23_1_y0;
  assign f_u_arrmul24_ha23_1_f_u_arrmul24_fa22_1_y4 = f_u_arrmul24_fa22_1_y4;
  assign f_u_arrmul24_ha23_1_y0 = f_u_arrmul24_ha23_1_f_u_arrmul24_and23_1_y0 ^ f_u_arrmul24_ha23_1_f_u_arrmul24_fa22_1_y4;
  assign f_u_arrmul24_ha23_1_y1 = f_u_arrmul24_ha23_1_f_u_arrmul24_and23_1_y0 & f_u_arrmul24_ha23_1_f_u_arrmul24_fa22_1_y4;
  assign f_u_arrmul24_and0_2_a_0 = a_0;
  assign f_u_arrmul24_and0_2_b_2 = b_2;
  assign f_u_arrmul24_and0_2_y0 = f_u_arrmul24_and0_2_a_0 & f_u_arrmul24_and0_2_b_2;
  assign f_u_arrmul24_ha0_2_f_u_arrmul24_and0_2_y0 = f_u_arrmul24_and0_2_y0;
  assign f_u_arrmul24_ha0_2_f_u_arrmul24_fa1_1_y2 = f_u_arrmul24_fa1_1_y2;
  assign f_u_arrmul24_ha0_2_y0 = f_u_arrmul24_ha0_2_f_u_arrmul24_and0_2_y0 ^ f_u_arrmul24_ha0_2_f_u_arrmul24_fa1_1_y2;
  assign f_u_arrmul24_ha0_2_y1 = f_u_arrmul24_ha0_2_f_u_arrmul24_and0_2_y0 & f_u_arrmul24_ha0_2_f_u_arrmul24_fa1_1_y2;
  assign f_u_arrmul24_and1_2_a_1 = a_1;
  assign f_u_arrmul24_and1_2_b_2 = b_2;
  assign f_u_arrmul24_and1_2_y0 = f_u_arrmul24_and1_2_a_1 & f_u_arrmul24_and1_2_b_2;
  assign f_u_arrmul24_fa1_2_f_u_arrmul24_and1_2_y0 = f_u_arrmul24_and1_2_y0;
  assign f_u_arrmul24_fa1_2_f_u_arrmul24_fa2_1_y2 = f_u_arrmul24_fa2_1_y2;
  assign f_u_arrmul24_fa1_2_f_u_arrmul24_ha0_2_y1 = f_u_arrmul24_ha0_2_y1;
  assign f_u_arrmul24_fa1_2_y0 = f_u_arrmul24_fa1_2_f_u_arrmul24_and1_2_y0 ^ f_u_arrmul24_fa1_2_f_u_arrmul24_fa2_1_y2;
  assign f_u_arrmul24_fa1_2_y1 = f_u_arrmul24_fa1_2_f_u_arrmul24_and1_2_y0 & f_u_arrmul24_fa1_2_f_u_arrmul24_fa2_1_y2;
  assign f_u_arrmul24_fa1_2_y2 = f_u_arrmul24_fa1_2_y0 ^ f_u_arrmul24_fa1_2_f_u_arrmul24_ha0_2_y1;
  assign f_u_arrmul24_fa1_2_y3 = f_u_arrmul24_fa1_2_y0 & f_u_arrmul24_fa1_2_f_u_arrmul24_ha0_2_y1;
  assign f_u_arrmul24_fa1_2_y4 = f_u_arrmul24_fa1_2_y1 | f_u_arrmul24_fa1_2_y3;
  assign f_u_arrmul24_and2_2_a_2 = a_2;
  assign f_u_arrmul24_and2_2_b_2 = b_2;
  assign f_u_arrmul24_and2_2_y0 = f_u_arrmul24_and2_2_a_2 & f_u_arrmul24_and2_2_b_2;
  assign f_u_arrmul24_fa2_2_f_u_arrmul24_and2_2_y0 = f_u_arrmul24_and2_2_y0;
  assign f_u_arrmul24_fa2_2_f_u_arrmul24_fa3_1_y2 = f_u_arrmul24_fa3_1_y2;
  assign f_u_arrmul24_fa2_2_f_u_arrmul24_fa1_2_y4 = f_u_arrmul24_fa1_2_y4;
  assign f_u_arrmul24_fa2_2_y0 = f_u_arrmul24_fa2_2_f_u_arrmul24_and2_2_y0 ^ f_u_arrmul24_fa2_2_f_u_arrmul24_fa3_1_y2;
  assign f_u_arrmul24_fa2_2_y1 = f_u_arrmul24_fa2_2_f_u_arrmul24_and2_2_y0 & f_u_arrmul24_fa2_2_f_u_arrmul24_fa3_1_y2;
  assign f_u_arrmul24_fa2_2_y2 = f_u_arrmul24_fa2_2_y0 ^ f_u_arrmul24_fa2_2_f_u_arrmul24_fa1_2_y4;
  assign f_u_arrmul24_fa2_2_y3 = f_u_arrmul24_fa2_2_y0 & f_u_arrmul24_fa2_2_f_u_arrmul24_fa1_2_y4;
  assign f_u_arrmul24_fa2_2_y4 = f_u_arrmul24_fa2_2_y1 | f_u_arrmul24_fa2_2_y3;
  assign f_u_arrmul24_and3_2_a_3 = a_3;
  assign f_u_arrmul24_and3_2_b_2 = b_2;
  assign f_u_arrmul24_and3_2_y0 = f_u_arrmul24_and3_2_a_3 & f_u_arrmul24_and3_2_b_2;
  assign f_u_arrmul24_fa3_2_f_u_arrmul24_and3_2_y0 = f_u_arrmul24_and3_2_y0;
  assign f_u_arrmul24_fa3_2_f_u_arrmul24_fa4_1_y2 = f_u_arrmul24_fa4_1_y2;
  assign f_u_arrmul24_fa3_2_f_u_arrmul24_fa2_2_y4 = f_u_arrmul24_fa2_2_y4;
  assign f_u_arrmul24_fa3_2_y0 = f_u_arrmul24_fa3_2_f_u_arrmul24_and3_2_y0 ^ f_u_arrmul24_fa3_2_f_u_arrmul24_fa4_1_y2;
  assign f_u_arrmul24_fa3_2_y1 = f_u_arrmul24_fa3_2_f_u_arrmul24_and3_2_y0 & f_u_arrmul24_fa3_2_f_u_arrmul24_fa4_1_y2;
  assign f_u_arrmul24_fa3_2_y2 = f_u_arrmul24_fa3_2_y0 ^ f_u_arrmul24_fa3_2_f_u_arrmul24_fa2_2_y4;
  assign f_u_arrmul24_fa3_2_y3 = f_u_arrmul24_fa3_2_y0 & f_u_arrmul24_fa3_2_f_u_arrmul24_fa2_2_y4;
  assign f_u_arrmul24_fa3_2_y4 = f_u_arrmul24_fa3_2_y1 | f_u_arrmul24_fa3_2_y3;
  assign f_u_arrmul24_and4_2_a_4 = a_4;
  assign f_u_arrmul24_and4_2_b_2 = b_2;
  assign f_u_arrmul24_and4_2_y0 = f_u_arrmul24_and4_2_a_4 & f_u_arrmul24_and4_2_b_2;
  assign f_u_arrmul24_fa4_2_f_u_arrmul24_and4_2_y0 = f_u_arrmul24_and4_2_y0;
  assign f_u_arrmul24_fa4_2_f_u_arrmul24_fa5_1_y2 = f_u_arrmul24_fa5_1_y2;
  assign f_u_arrmul24_fa4_2_f_u_arrmul24_fa3_2_y4 = f_u_arrmul24_fa3_2_y4;
  assign f_u_arrmul24_fa4_2_y0 = f_u_arrmul24_fa4_2_f_u_arrmul24_and4_2_y0 ^ f_u_arrmul24_fa4_2_f_u_arrmul24_fa5_1_y2;
  assign f_u_arrmul24_fa4_2_y1 = f_u_arrmul24_fa4_2_f_u_arrmul24_and4_2_y0 & f_u_arrmul24_fa4_2_f_u_arrmul24_fa5_1_y2;
  assign f_u_arrmul24_fa4_2_y2 = f_u_arrmul24_fa4_2_y0 ^ f_u_arrmul24_fa4_2_f_u_arrmul24_fa3_2_y4;
  assign f_u_arrmul24_fa4_2_y3 = f_u_arrmul24_fa4_2_y0 & f_u_arrmul24_fa4_2_f_u_arrmul24_fa3_2_y4;
  assign f_u_arrmul24_fa4_2_y4 = f_u_arrmul24_fa4_2_y1 | f_u_arrmul24_fa4_2_y3;
  assign f_u_arrmul24_and5_2_a_5 = a_5;
  assign f_u_arrmul24_and5_2_b_2 = b_2;
  assign f_u_arrmul24_and5_2_y0 = f_u_arrmul24_and5_2_a_5 & f_u_arrmul24_and5_2_b_2;
  assign f_u_arrmul24_fa5_2_f_u_arrmul24_and5_2_y0 = f_u_arrmul24_and5_2_y0;
  assign f_u_arrmul24_fa5_2_f_u_arrmul24_fa6_1_y2 = f_u_arrmul24_fa6_1_y2;
  assign f_u_arrmul24_fa5_2_f_u_arrmul24_fa4_2_y4 = f_u_arrmul24_fa4_2_y4;
  assign f_u_arrmul24_fa5_2_y0 = f_u_arrmul24_fa5_2_f_u_arrmul24_and5_2_y0 ^ f_u_arrmul24_fa5_2_f_u_arrmul24_fa6_1_y2;
  assign f_u_arrmul24_fa5_2_y1 = f_u_arrmul24_fa5_2_f_u_arrmul24_and5_2_y0 & f_u_arrmul24_fa5_2_f_u_arrmul24_fa6_1_y2;
  assign f_u_arrmul24_fa5_2_y2 = f_u_arrmul24_fa5_2_y0 ^ f_u_arrmul24_fa5_2_f_u_arrmul24_fa4_2_y4;
  assign f_u_arrmul24_fa5_2_y3 = f_u_arrmul24_fa5_2_y0 & f_u_arrmul24_fa5_2_f_u_arrmul24_fa4_2_y4;
  assign f_u_arrmul24_fa5_2_y4 = f_u_arrmul24_fa5_2_y1 | f_u_arrmul24_fa5_2_y3;
  assign f_u_arrmul24_and6_2_a_6 = a_6;
  assign f_u_arrmul24_and6_2_b_2 = b_2;
  assign f_u_arrmul24_and6_2_y0 = f_u_arrmul24_and6_2_a_6 & f_u_arrmul24_and6_2_b_2;
  assign f_u_arrmul24_fa6_2_f_u_arrmul24_and6_2_y0 = f_u_arrmul24_and6_2_y0;
  assign f_u_arrmul24_fa6_2_f_u_arrmul24_fa7_1_y2 = f_u_arrmul24_fa7_1_y2;
  assign f_u_arrmul24_fa6_2_f_u_arrmul24_fa5_2_y4 = f_u_arrmul24_fa5_2_y4;
  assign f_u_arrmul24_fa6_2_y0 = f_u_arrmul24_fa6_2_f_u_arrmul24_and6_2_y0 ^ f_u_arrmul24_fa6_2_f_u_arrmul24_fa7_1_y2;
  assign f_u_arrmul24_fa6_2_y1 = f_u_arrmul24_fa6_2_f_u_arrmul24_and6_2_y0 & f_u_arrmul24_fa6_2_f_u_arrmul24_fa7_1_y2;
  assign f_u_arrmul24_fa6_2_y2 = f_u_arrmul24_fa6_2_y0 ^ f_u_arrmul24_fa6_2_f_u_arrmul24_fa5_2_y4;
  assign f_u_arrmul24_fa6_2_y3 = f_u_arrmul24_fa6_2_y0 & f_u_arrmul24_fa6_2_f_u_arrmul24_fa5_2_y4;
  assign f_u_arrmul24_fa6_2_y4 = f_u_arrmul24_fa6_2_y1 | f_u_arrmul24_fa6_2_y3;
  assign f_u_arrmul24_and7_2_a_7 = a_7;
  assign f_u_arrmul24_and7_2_b_2 = b_2;
  assign f_u_arrmul24_and7_2_y0 = f_u_arrmul24_and7_2_a_7 & f_u_arrmul24_and7_2_b_2;
  assign f_u_arrmul24_fa7_2_f_u_arrmul24_and7_2_y0 = f_u_arrmul24_and7_2_y0;
  assign f_u_arrmul24_fa7_2_f_u_arrmul24_fa8_1_y2 = f_u_arrmul24_fa8_1_y2;
  assign f_u_arrmul24_fa7_2_f_u_arrmul24_fa6_2_y4 = f_u_arrmul24_fa6_2_y4;
  assign f_u_arrmul24_fa7_2_y0 = f_u_arrmul24_fa7_2_f_u_arrmul24_and7_2_y0 ^ f_u_arrmul24_fa7_2_f_u_arrmul24_fa8_1_y2;
  assign f_u_arrmul24_fa7_2_y1 = f_u_arrmul24_fa7_2_f_u_arrmul24_and7_2_y0 & f_u_arrmul24_fa7_2_f_u_arrmul24_fa8_1_y2;
  assign f_u_arrmul24_fa7_2_y2 = f_u_arrmul24_fa7_2_y0 ^ f_u_arrmul24_fa7_2_f_u_arrmul24_fa6_2_y4;
  assign f_u_arrmul24_fa7_2_y3 = f_u_arrmul24_fa7_2_y0 & f_u_arrmul24_fa7_2_f_u_arrmul24_fa6_2_y4;
  assign f_u_arrmul24_fa7_2_y4 = f_u_arrmul24_fa7_2_y1 | f_u_arrmul24_fa7_2_y3;
  assign f_u_arrmul24_and8_2_a_8 = a_8;
  assign f_u_arrmul24_and8_2_b_2 = b_2;
  assign f_u_arrmul24_and8_2_y0 = f_u_arrmul24_and8_2_a_8 & f_u_arrmul24_and8_2_b_2;
  assign f_u_arrmul24_fa8_2_f_u_arrmul24_and8_2_y0 = f_u_arrmul24_and8_2_y0;
  assign f_u_arrmul24_fa8_2_f_u_arrmul24_fa9_1_y2 = f_u_arrmul24_fa9_1_y2;
  assign f_u_arrmul24_fa8_2_f_u_arrmul24_fa7_2_y4 = f_u_arrmul24_fa7_2_y4;
  assign f_u_arrmul24_fa8_2_y0 = f_u_arrmul24_fa8_2_f_u_arrmul24_and8_2_y0 ^ f_u_arrmul24_fa8_2_f_u_arrmul24_fa9_1_y2;
  assign f_u_arrmul24_fa8_2_y1 = f_u_arrmul24_fa8_2_f_u_arrmul24_and8_2_y0 & f_u_arrmul24_fa8_2_f_u_arrmul24_fa9_1_y2;
  assign f_u_arrmul24_fa8_2_y2 = f_u_arrmul24_fa8_2_y0 ^ f_u_arrmul24_fa8_2_f_u_arrmul24_fa7_2_y4;
  assign f_u_arrmul24_fa8_2_y3 = f_u_arrmul24_fa8_2_y0 & f_u_arrmul24_fa8_2_f_u_arrmul24_fa7_2_y4;
  assign f_u_arrmul24_fa8_2_y4 = f_u_arrmul24_fa8_2_y1 | f_u_arrmul24_fa8_2_y3;
  assign f_u_arrmul24_and9_2_a_9 = a_9;
  assign f_u_arrmul24_and9_2_b_2 = b_2;
  assign f_u_arrmul24_and9_2_y0 = f_u_arrmul24_and9_2_a_9 & f_u_arrmul24_and9_2_b_2;
  assign f_u_arrmul24_fa9_2_f_u_arrmul24_and9_2_y0 = f_u_arrmul24_and9_2_y0;
  assign f_u_arrmul24_fa9_2_f_u_arrmul24_fa10_1_y2 = f_u_arrmul24_fa10_1_y2;
  assign f_u_arrmul24_fa9_2_f_u_arrmul24_fa8_2_y4 = f_u_arrmul24_fa8_2_y4;
  assign f_u_arrmul24_fa9_2_y0 = f_u_arrmul24_fa9_2_f_u_arrmul24_and9_2_y0 ^ f_u_arrmul24_fa9_2_f_u_arrmul24_fa10_1_y2;
  assign f_u_arrmul24_fa9_2_y1 = f_u_arrmul24_fa9_2_f_u_arrmul24_and9_2_y0 & f_u_arrmul24_fa9_2_f_u_arrmul24_fa10_1_y2;
  assign f_u_arrmul24_fa9_2_y2 = f_u_arrmul24_fa9_2_y0 ^ f_u_arrmul24_fa9_2_f_u_arrmul24_fa8_2_y4;
  assign f_u_arrmul24_fa9_2_y3 = f_u_arrmul24_fa9_2_y0 & f_u_arrmul24_fa9_2_f_u_arrmul24_fa8_2_y4;
  assign f_u_arrmul24_fa9_2_y4 = f_u_arrmul24_fa9_2_y1 | f_u_arrmul24_fa9_2_y3;
  assign f_u_arrmul24_and10_2_a_10 = a_10;
  assign f_u_arrmul24_and10_2_b_2 = b_2;
  assign f_u_arrmul24_and10_2_y0 = f_u_arrmul24_and10_2_a_10 & f_u_arrmul24_and10_2_b_2;
  assign f_u_arrmul24_fa10_2_f_u_arrmul24_and10_2_y0 = f_u_arrmul24_and10_2_y0;
  assign f_u_arrmul24_fa10_2_f_u_arrmul24_fa11_1_y2 = f_u_arrmul24_fa11_1_y2;
  assign f_u_arrmul24_fa10_2_f_u_arrmul24_fa9_2_y4 = f_u_arrmul24_fa9_2_y4;
  assign f_u_arrmul24_fa10_2_y0 = f_u_arrmul24_fa10_2_f_u_arrmul24_and10_2_y0 ^ f_u_arrmul24_fa10_2_f_u_arrmul24_fa11_1_y2;
  assign f_u_arrmul24_fa10_2_y1 = f_u_arrmul24_fa10_2_f_u_arrmul24_and10_2_y0 & f_u_arrmul24_fa10_2_f_u_arrmul24_fa11_1_y2;
  assign f_u_arrmul24_fa10_2_y2 = f_u_arrmul24_fa10_2_y0 ^ f_u_arrmul24_fa10_2_f_u_arrmul24_fa9_2_y4;
  assign f_u_arrmul24_fa10_2_y3 = f_u_arrmul24_fa10_2_y0 & f_u_arrmul24_fa10_2_f_u_arrmul24_fa9_2_y4;
  assign f_u_arrmul24_fa10_2_y4 = f_u_arrmul24_fa10_2_y1 | f_u_arrmul24_fa10_2_y3;
  assign f_u_arrmul24_and11_2_a_11 = a_11;
  assign f_u_arrmul24_and11_2_b_2 = b_2;
  assign f_u_arrmul24_and11_2_y0 = f_u_arrmul24_and11_2_a_11 & f_u_arrmul24_and11_2_b_2;
  assign f_u_arrmul24_fa11_2_f_u_arrmul24_and11_2_y0 = f_u_arrmul24_and11_2_y0;
  assign f_u_arrmul24_fa11_2_f_u_arrmul24_fa12_1_y2 = f_u_arrmul24_fa12_1_y2;
  assign f_u_arrmul24_fa11_2_f_u_arrmul24_fa10_2_y4 = f_u_arrmul24_fa10_2_y4;
  assign f_u_arrmul24_fa11_2_y0 = f_u_arrmul24_fa11_2_f_u_arrmul24_and11_2_y0 ^ f_u_arrmul24_fa11_2_f_u_arrmul24_fa12_1_y2;
  assign f_u_arrmul24_fa11_2_y1 = f_u_arrmul24_fa11_2_f_u_arrmul24_and11_2_y0 & f_u_arrmul24_fa11_2_f_u_arrmul24_fa12_1_y2;
  assign f_u_arrmul24_fa11_2_y2 = f_u_arrmul24_fa11_2_y0 ^ f_u_arrmul24_fa11_2_f_u_arrmul24_fa10_2_y4;
  assign f_u_arrmul24_fa11_2_y3 = f_u_arrmul24_fa11_2_y0 & f_u_arrmul24_fa11_2_f_u_arrmul24_fa10_2_y4;
  assign f_u_arrmul24_fa11_2_y4 = f_u_arrmul24_fa11_2_y1 | f_u_arrmul24_fa11_2_y3;
  assign f_u_arrmul24_and12_2_a_12 = a_12;
  assign f_u_arrmul24_and12_2_b_2 = b_2;
  assign f_u_arrmul24_and12_2_y0 = f_u_arrmul24_and12_2_a_12 & f_u_arrmul24_and12_2_b_2;
  assign f_u_arrmul24_fa12_2_f_u_arrmul24_and12_2_y0 = f_u_arrmul24_and12_2_y0;
  assign f_u_arrmul24_fa12_2_f_u_arrmul24_fa13_1_y2 = f_u_arrmul24_fa13_1_y2;
  assign f_u_arrmul24_fa12_2_f_u_arrmul24_fa11_2_y4 = f_u_arrmul24_fa11_2_y4;
  assign f_u_arrmul24_fa12_2_y0 = f_u_arrmul24_fa12_2_f_u_arrmul24_and12_2_y0 ^ f_u_arrmul24_fa12_2_f_u_arrmul24_fa13_1_y2;
  assign f_u_arrmul24_fa12_2_y1 = f_u_arrmul24_fa12_2_f_u_arrmul24_and12_2_y0 & f_u_arrmul24_fa12_2_f_u_arrmul24_fa13_1_y2;
  assign f_u_arrmul24_fa12_2_y2 = f_u_arrmul24_fa12_2_y0 ^ f_u_arrmul24_fa12_2_f_u_arrmul24_fa11_2_y4;
  assign f_u_arrmul24_fa12_2_y3 = f_u_arrmul24_fa12_2_y0 & f_u_arrmul24_fa12_2_f_u_arrmul24_fa11_2_y4;
  assign f_u_arrmul24_fa12_2_y4 = f_u_arrmul24_fa12_2_y1 | f_u_arrmul24_fa12_2_y3;
  assign f_u_arrmul24_and13_2_a_13 = a_13;
  assign f_u_arrmul24_and13_2_b_2 = b_2;
  assign f_u_arrmul24_and13_2_y0 = f_u_arrmul24_and13_2_a_13 & f_u_arrmul24_and13_2_b_2;
  assign f_u_arrmul24_fa13_2_f_u_arrmul24_and13_2_y0 = f_u_arrmul24_and13_2_y0;
  assign f_u_arrmul24_fa13_2_f_u_arrmul24_fa14_1_y2 = f_u_arrmul24_fa14_1_y2;
  assign f_u_arrmul24_fa13_2_f_u_arrmul24_fa12_2_y4 = f_u_arrmul24_fa12_2_y4;
  assign f_u_arrmul24_fa13_2_y0 = f_u_arrmul24_fa13_2_f_u_arrmul24_and13_2_y0 ^ f_u_arrmul24_fa13_2_f_u_arrmul24_fa14_1_y2;
  assign f_u_arrmul24_fa13_2_y1 = f_u_arrmul24_fa13_2_f_u_arrmul24_and13_2_y0 & f_u_arrmul24_fa13_2_f_u_arrmul24_fa14_1_y2;
  assign f_u_arrmul24_fa13_2_y2 = f_u_arrmul24_fa13_2_y0 ^ f_u_arrmul24_fa13_2_f_u_arrmul24_fa12_2_y4;
  assign f_u_arrmul24_fa13_2_y3 = f_u_arrmul24_fa13_2_y0 & f_u_arrmul24_fa13_2_f_u_arrmul24_fa12_2_y4;
  assign f_u_arrmul24_fa13_2_y4 = f_u_arrmul24_fa13_2_y1 | f_u_arrmul24_fa13_2_y3;
  assign f_u_arrmul24_and14_2_a_14 = a_14;
  assign f_u_arrmul24_and14_2_b_2 = b_2;
  assign f_u_arrmul24_and14_2_y0 = f_u_arrmul24_and14_2_a_14 & f_u_arrmul24_and14_2_b_2;
  assign f_u_arrmul24_fa14_2_f_u_arrmul24_and14_2_y0 = f_u_arrmul24_and14_2_y0;
  assign f_u_arrmul24_fa14_2_f_u_arrmul24_fa15_1_y2 = f_u_arrmul24_fa15_1_y2;
  assign f_u_arrmul24_fa14_2_f_u_arrmul24_fa13_2_y4 = f_u_arrmul24_fa13_2_y4;
  assign f_u_arrmul24_fa14_2_y0 = f_u_arrmul24_fa14_2_f_u_arrmul24_and14_2_y0 ^ f_u_arrmul24_fa14_2_f_u_arrmul24_fa15_1_y2;
  assign f_u_arrmul24_fa14_2_y1 = f_u_arrmul24_fa14_2_f_u_arrmul24_and14_2_y0 & f_u_arrmul24_fa14_2_f_u_arrmul24_fa15_1_y2;
  assign f_u_arrmul24_fa14_2_y2 = f_u_arrmul24_fa14_2_y0 ^ f_u_arrmul24_fa14_2_f_u_arrmul24_fa13_2_y4;
  assign f_u_arrmul24_fa14_2_y3 = f_u_arrmul24_fa14_2_y0 & f_u_arrmul24_fa14_2_f_u_arrmul24_fa13_2_y4;
  assign f_u_arrmul24_fa14_2_y4 = f_u_arrmul24_fa14_2_y1 | f_u_arrmul24_fa14_2_y3;
  assign f_u_arrmul24_and15_2_a_15 = a_15;
  assign f_u_arrmul24_and15_2_b_2 = b_2;
  assign f_u_arrmul24_and15_2_y0 = f_u_arrmul24_and15_2_a_15 & f_u_arrmul24_and15_2_b_2;
  assign f_u_arrmul24_fa15_2_f_u_arrmul24_and15_2_y0 = f_u_arrmul24_and15_2_y0;
  assign f_u_arrmul24_fa15_2_f_u_arrmul24_fa16_1_y2 = f_u_arrmul24_fa16_1_y2;
  assign f_u_arrmul24_fa15_2_f_u_arrmul24_fa14_2_y4 = f_u_arrmul24_fa14_2_y4;
  assign f_u_arrmul24_fa15_2_y0 = f_u_arrmul24_fa15_2_f_u_arrmul24_and15_2_y0 ^ f_u_arrmul24_fa15_2_f_u_arrmul24_fa16_1_y2;
  assign f_u_arrmul24_fa15_2_y1 = f_u_arrmul24_fa15_2_f_u_arrmul24_and15_2_y0 & f_u_arrmul24_fa15_2_f_u_arrmul24_fa16_1_y2;
  assign f_u_arrmul24_fa15_2_y2 = f_u_arrmul24_fa15_2_y0 ^ f_u_arrmul24_fa15_2_f_u_arrmul24_fa14_2_y4;
  assign f_u_arrmul24_fa15_2_y3 = f_u_arrmul24_fa15_2_y0 & f_u_arrmul24_fa15_2_f_u_arrmul24_fa14_2_y4;
  assign f_u_arrmul24_fa15_2_y4 = f_u_arrmul24_fa15_2_y1 | f_u_arrmul24_fa15_2_y3;
  assign f_u_arrmul24_and16_2_a_16 = a_16;
  assign f_u_arrmul24_and16_2_b_2 = b_2;
  assign f_u_arrmul24_and16_2_y0 = f_u_arrmul24_and16_2_a_16 & f_u_arrmul24_and16_2_b_2;
  assign f_u_arrmul24_fa16_2_f_u_arrmul24_and16_2_y0 = f_u_arrmul24_and16_2_y0;
  assign f_u_arrmul24_fa16_2_f_u_arrmul24_fa17_1_y2 = f_u_arrmul24_fa17_1_y2;
  assign f_u_arrmul24_fa16_2_f_u_arrmul24_fa15_2_y4 = f_u_arrmul24_fa15_2_y4;
  assign f_u_arrmul24_fa16_2_y0 = f_u_arrmul24_fa16_2_f_u_arrmul24_and16_2_y0 ^ f_u_arrmul24_fa16_2_f_u_arrmul24_fa17_1_y2;
  assign f_u_arrmul24_fa16_2_y1 = f_u_arrmul24_fa16_2_f_u_arrmul24_and16_2_y0 & f_u_arrmul24_fa16_2_f_u_arrmul24_fa17_1_y2;
  assign f_u_arrmul24_fa16_2_y2 = f_u_arrmul24_fa16_2_y0 ^ f_u_arrmul24_fa16_2_f_u_arrmul24_fa15_2_y4;
  assign f_u_arrmul24_fa16_2_y3 = f_u_arrmul24_fa16_2_y0 & f_u_arrmul24_fa16_2_f_u_arrmul24_fa15_2_y4;
  assign f_u_arrmul24_fa16_2_y4 = f_u_arrmul24_fa16_2_y1 | f_u_arrmul24_fa16_2_y3;
  assign f_u_arrmul24_and17_2_a_17 = a_17;
  assign f_u_arrmul24_and17_2_b_2 = b_2;
  assign f_u_arrmul24_and17_2_y0 = f_u_arrmul24_and17_2_a_17 & f_u_arrmul24_and17_2_b_2;
  assign f_u_arrmul24_fa17_2_f_u_arrmul24_and17_2_y0 = f_u_arrmul24_and17_2_y0;
  assign f_u_arrmul24_fa17_2_f_u_arrmul24_fa18_1_y2 = f_u_arrmul24_fa18_1_y2;
  assign f_u_arrmul24_fa17_2_f_u_arrmul24_fa16_2_y4 = f_u_arrmul24_fa16_2_y4;
  assign f_u_arrmul24_fa17_2_y0 = f_u_arrmul24_fa17_2_f_u_arrmul24_and17_2_y0 ^ f_u_arrmul24_fa17_2_f_u_arrmul24_fa18_1_y2;
  assign f_u_arrmul24_fa17_2_y1 = f_u_arrmul24_fa17_2_f_u_arrmul24_and17_2_y0 & f_u_arrmul24_fa17_2_f_u_arrmul24_fa18_1_y2;
  assign f_u_arrmul24_fa17_2_y2 = f_u_arrmul24_fa17_2_y0 ^ f_u_arrmul24_fa17_2_f_u_arrmul24_fa16_2_y4;
  assign f_u_arrmul24_fa17_2_y3 = f_u_arrmul24_fa17_2_y0 & f_u_arrmul24_fa17_2_f_u_arrmul24_fa16_2_y4;
  assign f_u_arrmul24_fa17_2_y4 = f_u_arrmul24_fa17_2_y1 | f_u_arrmul24_fa17_2_y3;
  assign f_u_arrmul24_and18_2_a_18 = a_18;
  assign f_u_arrmul24_and18_2_b_2 = b_2;
  assign f_u_arrmul24_and18_2_y0 = f_u_arrmul24_and18_2_a_18 & f_u_arrmul24_and18_2_b_2;
  assign f_u_arrmul24_fa18_2_f_u_arrmul24_and18_2_y0 = f_u_arrmul24_and18_2_y0;
  assign f_u_arrmul24_fa18_2_f_u_arrmul24_fa19_1_y2 = f_u_arrmul24_fa19_1_y2;
  assign f_u_arrmul24_fa18_2_f_u_arrmul24_fa17_2_y4 = f_u_arrmul24_fa17_2_y4;
  assign f_u_arrmul24_fa18_2_y0 = f_u_arrmul24_fa18_2_f_u_arrmul24_and18_2_y0 ^ f_u_arrmul24_fa18_2_f_u_arrmul24_fa19_1_y2;
  assign f_u_arrmul24_fa18_2_y1 = f_u_arrmul24_fa18_2_f_u_arrmul24_and18_2_y0 & f_u_arrmul24_fa18_2_f_u_arrmul24_fa19_1_y2;
  assign f_u_arrmul24_fa18_2_y2 = f_u_arrmul24_fa18_2_y0 ^ f_u_arrmul24_fa18_2_f_u_arrmul24_fa17_2_y4;
  assign f_u_arrmul24_fa18_2_y3 = f_u_arrmul24_fa18_2_y0 & f_u_arrmul24_fa18_2_f_u_arrmul24_fa17_2_y4;
  assign f_u_arrmul24_fa18_2_y4 = f_u_arrmul24_fa18_2_y1 | f_u_arrmul24_fa18_2_y3;
  assign f_u_arrmul24_and19_2_a_19 = a_19;
  assign f_u_arrmul24_and19_2_b_2 = b_2;
  assign f_u_arrmul24_and19_2_y0 = f_u_arrmul24_and19_2_a_19 & f_u_arrmul24_and19_2_b_2;
  assign f_u_arrmul24_fa19_2_f_u_arrmul24_and19_2_y0 = f_u_arrmul24_and19_2_y0;
  assign f_u_arrmul24_fa19_2_f_u_arrmul24_fa20_1_y2 = f_u_arrmul24_fa20_1_y2;
  assign f_u_arrmul24_fa19_2_f_u_arrmul24_fa18_2_y4 = f_u_arrmul24_fa18_2_y4;
  assign f_u_arrmul24_fa19_2_y0 = f_u_arrmul24_fa19_2_f_u_arrmul24_and19_2_y0 ^ f_u_arrmul24_fa19_2_f_u_arrmul24_fa20_1_y2;
  assign f_u_arrmul24_fa19_2_y1 = f_u_arrmul24_fa19_2_f_u_arrmul24_and19_2_y0 & f_u_arrmul24_fa19_2_f_u_arrmul24_fa20_1_y2;
  assign f_u_arrmul24_fa19_2_y2 = f_u_arrmul24_fa19_2_y0 ^ f_u_arrmul24_fa19_2_f_u_arrmul24_fa18_2_y4;
  assign f_u_arrmul24_fa19_2_y3 = f_u_arrmul24_fa19_2_y0 & f_u_arrmul24_fa19_2_f_u_arrmul24_fa18_2_y4;
  assign f_u_arrmul24_fa19_2_y4 = f_u_arrmul24_fa19_2_y1 | f_u_arrmul24_fa19_2_y3;
  assign f_u_arrmul24_and20_2_a_20 = a_20;
  assign f_u_arrmul24_and20_2_b_2 = b_2;
  assign f_u_arrmul24_and20_2_y0 = f_u_arrmul24_and20_2_a_20 & f_u_arrmul24_and20_2_b_2;
  assign f_u_arrmul24_fa20_2_f_u_arrmul24_and20_2_y0 = f_u_arrmul24_and20_2_y0;
  assign f_u_arrmul24_fa20_2_f_u_arrmul24_fa21_1_y2 = f_u_arrmul24_fa21_1_y2;
  assign f_u_arrmul24_fa20_2_f_u_arrmul24_fa19_2_y4 = f_u_arrmul24_fa19_2_y4;
  assign f_u_arrmul24_fa20_2_y0 = f_u_arrmul24_fa20_2_f_u_arrmul24_and20_2_y0 ^ f_u_arrmul24_fa20_2_f_u_arrmul24_fa21_1_y2;
  assign f_u_arrmul24_fa20_2_y1 = f_u_arrmul24_fa20_2_f_u_arrmul24_and20_2_y0 & f_u_arrmul24_fa20_2_f_u_arrmul24_fa21_1_y2;
  assign f_u_arrmul24_fa20_2_y2 = f_u_arrmul24_fa20_2_y0 ^ f_u_arrmul24_fa20_2_f_u_arrmul24_fa19_2_y4;
  assign f_u_arrmul24_fa20_2_y3 = f_u_arrmul24_fa20_2_y0 & f_u_arrmul24_fa20_2_f_u_arrmul24_fa19_2_y4;
  assign f_u_arrmul24_fa20_2_y4 = f_u_arrmul24_fa20_2_y1 | f_u_arrmul24_fa20_2_y3;
  assign f_u_arrmul24_and21_2_a_21 = a_21;
  assign f_u_arrmul24_and21_2_b_2 = b_2;
  assign f_u_arrmul24_and21_2_y0 = f_u_arrmul24_and21_2_a_21 & f_u_arrmul24_and21_2_b_2;
  assign f_u_arrmul24_fa21_2_f_u_arrmul24_and21_2_y0 = f_u_arrmul24_and21_2_y0;
  assign f_u_arrmul24_fa21_2_f_u_arrmul24_fa22_1_y2 = f_u_arrmul24_fa22_1_y2;
  assign f_u_arrmul24_fa21_2_f_u_arrmul24_fa20_2_y4 = f_u_arrmul24_fa20_2_y4;
  assign f_u_arrmul24_fa21_2_y0 = f_u_arrmul24_fa21_2_f_u_arrmul24_and21_2_y0 ^ f_u_arrmul24_fa21_2_f_u_arrmul24_fa22_1_y2;
  assign f_u_arrmul24_fa21_2_y1 = f_u_arrmul24_fa21_2_f_u_arrmul24_and21_2_y0 & f_u_arrmul24_fa21_2_f_u_arrmul24_fa22_1_y2;
  assign f_u_arrmul24_fa21_2_y2 = f_u_arrmul24_fa21_2_y0 ^ f_u_arrmul24_fa21_2_f_u_arrmul24_fa20_2_y4;
  assign f_u_arrmul24_fa21_2_y3 = f_u_arrmul24_fa21_2_y0 & f_u_arrmul24_fa21_2_f_u_arrmul24_fa20_2_y4;
  assign f_u_arrmul24_fa21_2_y4 = f_u_arrmul24_fa21_2_y1 | f_u_arrmul24_fa21_2_y3;
  assign f_u_arrmul24_and22_2_a_22 = a_22;
  assign f_u_arrmul24_and22_2_b_2 = b_2;
  assign f_u_arrmul24_and22_2_y0 = f_u_arrmul24_and22_2_a_22 & f_u_arrmul24_and22_2_b_2;
  assign f_u_arrmul24_fa22_2_f_u_arrmul24_and22_2_y0 = f_u_arrmul24_and22_2_y0;
  assign f_u_arrmul24_fa22_2_f_u_arrmul24_ha23_1_y0 = f_u_arrmul24_ha23_1_y0;
  assign f_u_arrmul24_fa22_2_f_u_arrmul24_fa21_2_y4 = f_u_arrmul24_fa21_2_y4;
  assign f_u_arrmul24_fa22_2_y0 = f_u_arrmul24_fa22_2_f_u_arrmul24_and22_2_y0 ^ f_u_arrmul24_fa22_2_f_u_arrmul24_ha23_1_y0;
  assign f_u_arrmul24_fa22_2_y1 = f_u_arrmul24_fa22_2_f_u_arrmul24_and22_2_y0 & f_u_arrmul24_fa22_2_f_u_arrmul24_ha23_1_y0;
  assign f_u_arrmul24_fa22_2_y2 = f_u_arrmul24_fa22_2_y0 ^ f_u_arrmul24_fa22_2_f_u_arrmul24_fa21_2_y4;
  assign f_u_arrmul24_fa22_2_y3 = f_u_arrmul24_fa22_2_y0 & f_u_arrmul24_fa22_2_f_u_arrmul24_fa21_2_y4;
  assign f_u_arrmul24_fa22_2_y4 = f_u_arrmul24_fa22_2_y1 | f_u_arrmul24_fa22_2_y3;
  assign f_u_arrmul24_and23_2_a_23 = a_23;
  assign f_u_arrmul24_and23_2_b_2 = b_2;
  assign f_u_arrmul24_and23_2_y0 = f_u_arrmul24_and23_2_a_23 & f_u_arrmul24_and23_2_b_2;
  assign f_u_arrmul24_fa23_2_f_u_arrmul24_and23_2_y0 = f_u_arrmul24_and23_2_y0;
  assign f_u_arrmul24_fa23_2_f_u_arrmul24_ha23_1_y1 = f_u_arrmul24_ha23_1_y1;
  assign f_u_arrmul24_fa23_2_f_u_arrmul24_fa22_2_y4 = f_u_arrmul24_fa22_2_y4;
  assign f_u_arrmul24_fa23_2_y0 = f_u_arrmul24_fa23_2_f_u_arrmul24_and23_2_y0 ^ f_u_arrmul24_fa23_2_f_u_arrmul24_ha23_1_y1;
  assign f_u_arrmul24_fa23_2_y1 = f_u_arrmul24_fa23_2_f_u_arrmul24_and23_2_y0 & f_u_arrmul24_fa23_2_f_u_arrmul24_ha23_1_y1;
  assign f_u_arrmul24_fa23_2_y2 = f_u_arrmul24_fa23_2_y0 ^ f_u_arrmul24_fa23_2_f_u_arrmul24_fa22_2_y4;
  assign f_u_arrmul24_fa23_2_y3 = f_u_arrmul24_fa23_2_y0 & f_u_arrmul24_fa23_2_f_u_arrmul24_fa22_2_y4;
  assign f_u_arrmul24_fa23_2_y4 = f_u_arrmul24_fa23_2_y1 | f_u_arrmul24_fa23_2_y3;
  assign f_u_arrmul24_and0_3_a_0 = a_0;
  assign f_u_arrmul24_and0_3_b_3 = b_3;
  assign f_u_arrmul24_and0_3_y0 = f_u_arrmul24_and0_3_a_0 & f_u_arrmul24_and0_3_b_3;
  assign f_u_arrmul24_ha0_3_f_u_arrmul24_and0_3_y0 = f_u_arrmul24_and0_3_y0;
  assign f_u_arrmul24_ha0_3_f_u_arrmul24_fa1_2_y2 = f_u_arrmul24_fa1_2_y2;
  assign f_u_arrmul24_ha0_3_y0 = f_u_arrmul24_ha0_3_f_u_arrmul24_and0_3_y0 ^ f_u_arrmul24_ha0_3_f_u_arrmul24_fa1_2_y2;
  assign f_u_arrmul24_ha0_3_y1 = f_u_arrmul24_ha0_3_f_u_arrmul24_and0_3_y0 & f_u_arrmul24_ha0_3_f_u_arrmul24_fa1_2_y2;
  assign f_u_arrmul24_and1_3_a_1 = a_1;
  assign f_u_arrmul24_and1_3_b_3 = b_3;
  assign f_u_arrmul24_and1_3_y0 = f_u_arrmul24_and1_3_a_1 & f_u_arrmul24_and1_3_b_3;
  assign f_u_arrmul24_fa1_3_f_u_arrmul24_and1_3_y0 = f_u_arrmul24_and1_3_y0;
  assign f_u_arrmul24_fa1_3_f_u_arrmul24_fa2_2_y2 = f_u_arrmul24_fa2_2_y2;
  assign f_u_arrmul24_fa1_3_f_u_arrmul24_ha0_3_y1 = f_u_arrmul24_ha0_3_y1;
  assign f_u_arrmul24_fa1_3_y0 = f_u_arrmul24_fa1_3_f_u_arrmul24_and1_3_y0 ^ f_u_arrmul24_fa1_3_f_u_arrmul24_fa2_2_y2;
  assign f_u_arrmul24_fa1_3_y1 = f_u_arrmul24_fa1_3_f_u_arrmul24_and1_3_y0 & f_u_arrmul24_fa1_3_f_u_arrmul24_fa2_2_y2;
  assign f_u_arrmul24_fa1_3_y2 = f_u_arrmul24_fa1_3_y0 ^ f_u_arrmul24_fa1_3_f_u_arrmul24_ha0_3_y1;
  assign f_u_arrmul24_fa1_3_y3 = f_u_arrmul24_fa1_3_y0 & f_u_arrmul24_fa1_3_f_u_arrmul24_ha0_3_y1;
  assign f_u_arrmul24_fa1_3_y4 = f_u_arrmul24_fa1_3_y1 | f_u_arrmul24_fa1_3_y3;
  assign f_u_arrmul24_and2_3_a_2 = a_2;
  assign f_u_arrmul24_and2_3_b_3 = b_3;
  assign f_u_arrmul24_and2_3_y0 = f_u_arrmul24_and2_3_a_2 & f_u_arrmul24_and2_3_b_3;
  assign f_u_arrmul24_fa2_3_f_u_arrmul24_and2_3_y0 = f_u_arrmul24_and2_3_y0;
  assign f_u_arrmul24_fa2_3_f_u_arrmul24_fa3_2_y2 = f_u_arrmul24_fa3_2_y2;
  assign f_u_arrmul24_fa2_3_f_u_arrmul24_fa1_3_y4 = f_u_arrmul24_fa1_3_y4;
  assign f_u_arrmul24_fa2_3_y0 = f_u_arrmul24_fa2_3_f_u_arrmul24_and2_3_y0 ^ f_u_arrmul24_fa2_3_f_u_arrmul24_fa3_2_y2;
  assign f_u_arrmul24_fa2_3_y1 = f_u_arrmul24_fa2_3_f_u_arrmul24_and2_3_y0 & f_u_arrmul24_fa2_3_f_u_arrmul24_fa3_2_y2;
  assign f_u_arrmul24_fa2_3_y2 = f_u_arrmul24_fa2_3_y0 ^ f_u_arrmul24_fa2_3_f_u_arrmul24_fa1_3_y4;
  assign f_u_arrmul24_fa2_3_y3 = f_u_arrmul24_fa2_3_y0 & f_u_arrmul24_fa2_3_f_u_arrmul24_fa1_3_y4;
  assign f_u_arrmul24_fa2_3_y4 = f_u_arrmul24_fa2_3_y1 | f_u_arrmul24_fa2_3_y3;
  assign f_u_arrmul24_and3_3_a_3 = a_3;
  assign f_u_arrmul24_and3_3_b_3 = b_3;
  assign f_u_arrmul24_and3_3_y0 = f_u_arrmul24_and3_3_a_3 & f_u_arrmul24_and3_3_b_3;
  assign f_u_arrmul24_fa3_3_f_u_arrmul24_and3_3_y0 = f_u_arrmul24_and3_3_y0;
  assign f_u_arrmul24_fa3_3_f_u_arrmul24_fa4_2_y2 = f_u_arrmul24_fa4_2_y2;
  assign f_u_arrmul24_fa3_3_f_u_arrmul24_fa2_3_y4 = f_u_arrmul24_fa2_3_y4;
  assign f_u_arrmul24_fa3_3_y0 = f_u_arrmul24_fa3_3_f_u_arrmul24_and3_3_y0 ^ f_u_arrmul24_fa3_3_f_u_arrmul24_fa4_2_y2;
  assign f_u_arrmul24_fa3_3_y1 = f_u_arrmul24_fa3_3_f_u_arrmul24_and3_3_y0 & f_u_arrmul24_fa3_3_f_u_arrmul24_fa4_2_y2;
  assign f_u_arrmul24_fa3_3_y2 = f_u_arrmul24_fa3_3_y0 ^ f_u_arrmul24_fa3_3_f_u_arrmul24_fa2_3_y4;
  assign f_u_arrmul24_fa3_3_y3 = f_u_arrmul24_fa3_3_y0 & f_u_arrmul24_fa3_3_f_u_arrmul24_fa2_3_y4;
  assign f_u_arrmul24_fa3_3_y4 = f_u_arrmul24_fa3_3_y1 | f_u_arrmul24_fa3_3_y3;
  assign f_u_arrmul24_and4_3_a_4 = a_4;
  assign f_u_arrmul24_and4_3_b_3 = b_3;
  assign f_u_arrmul24_and4_3_y0 = f_u_arrmul24_and4_3_a_4 & f_u_arrmul24_and4_3_b_3;
  assign f_u_arrmul24_fa4_3_f_u_arrmul24_and4_3_y0 = f_u_arrmul24_and4_3_y0;
  assign f_u_arrmul24_fa4_3_f_u_arrmul24_fa5_2_y2 = f_u_arrmul24_fa5_2_y2;
  assign f_u_arrmul24_fa4_3_f_u_arrmul24_fa3_3_y4 = f_u_arrmul24_fa3_3_y4;
  assign f_u_arrmul24_fa4_3_y0 = f_u_arrmul24_fa4_3_f_u_arrmul24_and4_3_y0 ^ f_u_arrmul24_fa4_3_f_u_arrmul24_fa5_2_y2;
  assign f_u_arrmul24_fa4_3_y1 = f_u_arrmul24_fa4_3_f_u_arrmul24_and4_3_y0 & f_u_arrmul24_fa4_3_f_u_arrmul24_fa5_2_y2;
  assign f_u_arrmul24_fa4_3_y2 = f_u_arrmul24_fa4_3_y0 ^ f_u_arrmul24_fa4_3_f_u_arrmul24_fa3_3_y4;
  assign f_u_arrmul24_fa4_3_y3 = f_u_arrmul24_fa4_3_y0 & f_u_arrmul24_fa4_3_f_u_arrmul24_fa3_3_y4;
  assign f_u_arrmul24_fa4_3_y4 = f_u_arrmul24_fa4_3_y1 | f_u_arrmul24_fa4_3_y3;
  assign f_u_arrmul24_and5_3_a_5 = a_5;
  assign f_u_arrmul24_and5_3_b_3 = b_3;
  assign f_u_arrmul24_and5_3_y0 = f_u_arrmul24_and5_3_a_5 & f_u_arrmul24_and5_3_b_3;
  assign f_u_arrmul24_fa5_3_f_u_arrmul24_and5_3_y0 = f_u_arrmul24_and5_3_y0;
  assign f_u_arrmul24_fa5_3_f_u_arrmul24_fa6_2_y2 = f_u_arrmul24_fa6_2_y2;
  assign f_u_arrmul24_fa5_3_f_u_arrmul24_fa4_3_y4 = f_u_arrmul24_fa4_3_y4;
  assign f_u_arrmul24_fa5_3_y0 = f_u_arrmul24_fa5_3_f_u_arrmul24_and5_3_y0 ^ f_u_arrmul24_fa5_3_f_u_arrmul24_fa6_2_y2;
  assign f_u_arrmul24_fa5_3_y1 = f_u_arrmul24_fa5_3_f_u_arrmul24_and5_3_y0 & f_u_arrmul24_fa5_3_f_u_arrmul24_fa6_2_y2;
  assign f_u_arrmul24_fa5_3_y2 = f_u_arrmul24_fa5_3_y0 ^ f_u_arrmul24_fa5_3_f_u_arrmul24_fa4_3_y4;
  assign f_u_arrmul24_fa5_3_y3 = f_u_arrmul24_fa5_3_y0 & f_u_arrmul24_fa5_3_f_u_arrmul24_fa4_3_y4;
  assign f_u_arrmul24_fa5_3_y4 = f_u_arrmul24_fa5_3_y1 | f_u_arrmul24_fa5_3_y3;
  assign f_u_arrmul24_and6_3_a_6 = a_6;
  assign f_u_arrmul24_and6_3_b_3 = b_3;
  assign f_u_arrmul24_and6_3_y0 = f_u_arrmul24_and6_3_a_6 & f_u_arrmul24_and6_3_b_3;
  assign f_u_arrmul24_fa6_3_f_u_arrmul24_and6_3_y0 = f_u_arrmul24_and6_3_y0;
  assign f_u_arrmul24_fa6_3_f_u_arrmul24_fa7_2_y2 = f_u_arrmul24_fa7_2_y2;
  assign f_u_arrmul24_fa6_3_f_u_arrmul24_fa5_3_y4 = f_u_arrmul24_fa5_3_y4;
  assign f_u_arrmul24_fa6_3_y0 = f_u_arrmul24_fa6_3_f_u_arrmul24_and6_3_y0 ^ f_u_arrmul24_fa6_3_f_u_arrmul24_fa7_2_y2;
  assign f_u_arrmul24_fa6_3_y1 = f_u_arrmul24_fa6_3_f_u_arrmul24_and6_3_y0 & f_u_arrmul24_fa6_3_f_u_arrmul24_fa7_2_y2;
  assign f_u_arrmul24_fa6_3_y2 = f_u_arrmul24_fa6_3_y0 ^ f_u_arrmul24_fa6_3_f_u_arrmul24_fa5_3_y4;
  assign f_u_arrmul24_fa6_3_y3 = f_u_arrmul24_fa6_3_y0 & f_u_arrmul24_fa6_3_f_u_arrmul24_fa5_3_y4;
  assign f_u_arrmul24_fa6_3_y4 = f_u_arrmul24_fa6_3_y1 | f_u_arrmul24_fa6_3_y3;
  assign f_u_arrmul24_and7_3_a_7 = a_7;
  assign f_u_arrmul24_and7_3_b_3 = b_3;
  assign f_u_arrmul24_and7_3_y0 = f_u_arrmul24_and7_3_a_7 & f_u_arrmul24_and7_3_b_3;
  assign f_u_arrmul24_fa7_3_f_u_arrmul24_and7_3_y0 = f_u_arrmul24_and7_3_y0;
  assign f_u_arrmul24_fa7_3_f_u_arrmul24_fa8_2_y2 = f_u_arrmul24_fa8_2_y2;
  assign f_u_arrmul24_fa7_3_f_u_arrmul24_fa6_3_y4 = f_u_arrmul24_fa6_3_y4;
  assign f_u_arrmul24_fa7_3_y0 = f_u_arrmul24_fa7_3_f_u_arrmul24_and7_3_y0 ^ f_u_arrmul24_fa7_3_f_u_arrmul24_fa8_2_y2;
  assign f_u_arrmul24_fa7_3_y1 = f_u_arrmul24_fa7_3_f_u_arrmul24_and7_3_y0 & f_u_arrmul24_fa7_3_f_u_arrmul24_fa8_2_y2;
  assign f_u_arrmul24_fa7_3_y2 = f_u_arrmul24_fa7_3_y0 ^ f_u_arrmul24_fa7_3_f_u_arrmul24_fa6_3_y4;
  assign f_u_arrmul24_fa7_3_y3 = f_u_arrmul24_fa7_3_y0 & f_u_arrmul24_fa7_3_f_u_arrmul24_fa6_3_y4;
  assign f_u_arrmul24_fa7_3_y4 = f_u_arrmul24_fa7_3_y1 | f_u_arrmul24_fa7_3_y3;
  assign f_u_arrmul24_and8_3_a_8 = a_8;
  assign f_u_arrmul24_and8_3_b_3 = b_3;
  assign f_u_arrmul24_and8_3_y0 = f_u_arrmul24_and8_3_a_8 & f_u_arrmul24_and8_3_b_3;
  assign f_u_arrmul24_fa8_3_f_u_arrmul24_and8_3_y0 = f_u_arrmul24_and8_3_y0;
  assign f_u_arrmul24_fa8_3_f_u_arrmul24_fa9_2_y2 = f_u_arrmul24_fa9_2_y2;
  assign f_u_arrmul24_fa8_3_f_u_arrmul24_fa7_3_y4 = f_u_arrmul24_fa7_3_y4;
  assign f_u_arrmul24_fa8_3_y0 = f_u_arrmul24_fa8_3_f_u_arrmul24_and8_3_y0 ^ f_u_arrmul24_fa8_3_f_u_arrmul24_fa9_2_y2;
  assign f_u_arrmul24_fa8_3_y1 = f_u_arrmul24_fa8_3_f_u_arrmul24_and8_3_y0 & f_u_arrmul24_fa8_3_f_u_arrmul24_fa9_2_y2;
  assign f_u_arrmul24_fa8_3_y2 = f_u_arrmul24_fa8_3_y0 ^ f_u_arrmul24_fa8_3_f_u_arrmul24_fa7_3_y4;
  assign f_u_arrmul24_fa8_3_y3 = f_u_arrmul24_fa8_3_y0 & f_u_arrmul24_fa8_3_f_u_arrmul24_fa7_3_y4;
  assign f_u_arrmul24_fa8_3_y4 = f_u_arrmul24_fa8_3_y1 | f_u_arrmul24_fa8_3_y3;
  assign f_u_arrmul24_and9_3_a_9 = a_9;
  assign f_u_arrmul24_and9_3_b_3 = b_3;
  assign f_u_arrmul24_and9_3_y0 = f_u_arrmul24_and9_3_a_9 & f_u_arrmul24_and9_3_b_3;
  assign f_u_arrmul24_fa9_3_f_u_arrmul24_and9_3_y0 = f_u_arrmul24_and9_3_y0;
  assign f_u_arrmul24_fa9_3_f_u_arrmul24_fa10_2_y2 = f_u_arrmul24_fa10_2_y2;
  assign f_u_arrmul24_fa9_3_f_u_arrmul24_fa8_3_y4 = f_u_arrmul24_fa8_3_y4;
  assign f_u_arrmul24_fa9_3_y0 = f_u_arrmul24_fa9_3_f_u_arrmul24_and9_3_y0 ^ f_u_arrmul24_fa9_3_f_u_arrmul24_fa10_2_y2;
  assign f_u_arrmul24_fa9_3_y1 = f_u_arrmul24_fa9_3_f_u_arrmul24_and9_3_y0 & f_u_arrmul24_fa9_3_f_u_arrmul24_fa10_2_y2;
  assign f_u_arrmul24_fa9_3_y2 = f_u_arrmul24_fa9_3_y0 ^ f_u_arrmul24_fa9_3_f_u_arrmul24_fa8_3_y4;
  assign f_u_arrmul24_fa9_3_y3 = f_u_arrmul24_fa9_3_y0 & f_u_arrmul24_fa9_3_f_u_arrmul24_fa8_3_y4;
  assign f_u_arrmul24_fa9_3_y4 = f_u_arrmul24_fa9_3_y1 | f_u_arrmul24_fa9_3_y3;
  assign f_u_arrmul24_and10_3_a_10 = a_10;
  assign f_u_arrmul24_and10_3_b_3 = b_3;
  assign f_u_arrmul24_and10_3_y0 = f_u_arrmul24_and10_3_a_10 & f_u_arrmul24_and10_3_b_3;
  assign f_u_arrmul24_fa10_3_f_u_arrmul24_and10_3_y0 = f_u_arrmul24_and10_3_y0;
  assign f_u_arrmul24_fa10_3_f_u_arrmul24_fa11_2_y2 = f_u_arrmul24_fa11_2_y2;
  assign f_u_arrmul24_fa10_3_f_u_arrmul24_fa9_3_y4 = f_u_arrmul24_fa9_3_y4;
  assign f_u_arrmul24_fa10_3_y0 = f_u_arrmul24_fa10_3_f_u_arrmul24_and10_3_y0 ^ f_u_arrmul24_fa10_3_f_u_arrmul24_fa11_2_y2;
  assign f_u_arrmul24_fa10_3_y1 = f_u_arrmul24_fa10_3_f_u_arrmul24_and10_3_y0 & f_u_arrmul24_fa10_3_f_u_arrmul24_fa11_2_y2;
  assign f_u_arrmul24_fa10_3_y2 = f_u_arrmul24_fa10_3_y0 ^ f_u_arrmul24_fa10_3_f_u_arrmul24_fa9_3_y4;
  assign f_u_arrmul24_fa10_3_y3 = f_u_arrmul24_fa10_3_y0 & f_u_arrmul24_fa10_3_f_u_arrmul24_fa9_3_y4;
  assign f_u_arrmul24_fa10_3_y4 = f_u_arrmul24_fa10_3_y1 | f_u_arrmul24_fa10_3_y3;
  assign f_u_arrmul24_and11_3_a_11 = a_11;
  assign f_u_arrmul24_and11_3_b_3 = b_3;
  assign f_u_arrmul24_and11_3_y0 = f_u_arrmul24_and11_3_a_11 & f_u_arrmul24_and11_3_b_3;
  assign f_u_arrmul24_fa11_3_f_u_arrmul24_and11_3_y0 = f_u_arrmul24_and11_3_y0;
  assign f_u_arrmul24_fa11_3_f_u_arrmul24_fa12_2_y2 = f_u_arrmul24_fa12_2_y2;
  assign f_u_arrmul24_fa11_3_f_u_arrmul24_fa10_3_y4 = f_u_arrmul24_fa10_3_y4;
  assign f_u_arrmul24_fa11_3_y0 = f_u_arrmul24_fa11_3_f_u_arrmul24_and11_3_y0 ^ f_u_arrmul24_fa11_3_f_u_arrmul24_fa12_2_y2;
  assign f_u_arrmul24_fa11_3_y1 = f_u_arrmul24_fa11_3_f_u_arrmul24_and11_3_y0 & f_u_arrmul24_fa11_3_f_u_arrmul24_fa12_2_y2;
  assign f_u_arrmul24_fa11_3_y2 = f_u_arrmul24_fa11_3_y0 ^ f_u_arrmul24_fa11_3_f_u_arrmul24_fa10_3_y4;
  assign f_u_arrmul24_fa11_3_y3 = f_u_arrmul24_fa11_3_y0 & f_u_arrmul24_fa11_3_f_u_arrmul24_fa10_3_y4;
  assign f_u_arrmul24_fa11_3_y4 = f_u_arrmul24_fa11_3_y1 | f_u_arrmul24_fa11_3_y3;
  assign f_u_arrmul24_and12_3_a_12 = a_12;
  assign f_u_arrmul24_and12_3_b_3 = b_3;
  assign f_u_arrmul24_and12_3_y0 = f_u_arrmul24_and12_3_a_12 & f_u_arrmul24_and12_3_b_3;
  assign f_u_arrmul24_fa12_3_f_u_arrmul24_and12_3_y0 = f_u_arrmul24_and12_3_y0;
  assign f_u_arrmul24_fa12_3_f_u_arrmul24_fa13_2_y2 = f_u_arrmul24_fa13_2_y2;
  assign f_u_arrmul24_fa12_3_f_u_arrmul24_fa11_3_y4 = f_u_arrmul24_fa11_3_y4;
  assign f_u_arrmul24_fa12_3_y0 = f_u_arrmul24_fa12_3_f_u_arrmul24_and12_3_y0 ^ f_u_arrmul24_fa12_3_f_u_arrmul24_fa13_2_y2;
  assign f_u_arrmul24_fa12_3_y1 = f_u_arrmul24_fa12_3_f_u_arrmul24_and12_3_y0 & f_u_arrmul24_fa12_3_f_u_arrmul24_fa13_2_y2;
  assign f_u_arrmul24_fa12_3_y2 = f_u_arrmul24_fa12_3_y0 ^ f_u_arrmul24_fa12_3_f_u_arrmul24_fa11_3_y4;
  assign f_u_arrmul24_fa12_3_y3 = f_u_arrmul24_fa12_3_y0 & f_u_arrmul24_fa12_3_f_u_arrmul24_fa11_3_y4;
  assign f_u_arrmul24_fa12_3_y4 = f_u_arrmul24_fa12_3_y1 | f_u_arrmul24_fa12_3_y3;
  assign f_u_arrmul24_and13_3_a_13 = a_13;
  assign f_u_arrmul24_and13_3_b_3 = b_3;
  assign f_u_arrmul24_and13_3_y0 = f_u_arrmul24_and13_3_a_13 & f_u_arrmul24_and13_3_b_3;
  assign f_u_arrmul24_fa13_3_f_u_arrmul24_and13_3_y0 = f_u_arrmul24_and13_3_y0;
  assign f_u_arrmul24_fa13_3_f_u_arrmul24_fa14_2_y2 = f_u_arrmul24_fa14_2_y2;
  assign f_u_arrmul24_fa13_3_f_u_arrmul24_fa12_3_y4 = f_u_arrmul24_fa12_3_y4;
  assign f_u_arrmul24_fa13_3_y0 = f_u_arrmul24_fa13_3_f_u_arrmul24_and13_3_y0 ^ f_u_arrmul24_fa13_3_f_u_arrmul24_fa14_2_y2;
  assign f_u_arrmul24_fa13_3_y1 = f_u_arrmul24_fa13_3_f_u_arrmul24_and13_3_y0 & f_u_arrmul24_fa13_3_f_u_arrmul24_fa14_2_y2;
  assign f_u_arrmul24_fa13_3_y2 = f_u_arrmul24_fa13_3_y0 ^ f_u_arrmul24_fa13_3_f_u_arrmul24_fa12_3_y4;
  assign f_u_arrmul24_fa13_3_y3 = f_u_arrmul24_fa13_3_y0 & f_u_arrmul24_fa13_3_f_u_arrmul24_fa12_3_y4;
  assign f_u_arrmul24_fa13_3_y4 = f_u_arrmul24_fa13_3_y1 | f_u_arrmul24_fa13_3_y3;
  assign f_u_arrmul24_and14_3_a_14 = a_14;
  assign f_u_arrmul24_and14_3_b_3 = b_3;
  assign f_u_arrmul24_and14_3_y0 = f_u_arrmul24_and14_3_a_14 & f_u_arrmul24_and14_3_b_3;
  assign f_u_arrmul24_fa14_3_f_u_arrmul24_and14_3_y0 = f_u_arrmul24_and14_3_y0;
  assign f_u_arrmul24_fa14_3_f_u_arrmul24_fa15_2_y2 = f_u_arrmul24_fa15_2_y2;
  assign f_u_arrmul24_fa14_3_f_u_arrmul24_fa13_3_y4 = f_u_arrmul24_fa13_3_y4;
  assign f_u_arrmul24_fa14_3_y0 = f_u_arrmul24_fa14_3_f_u_arrmul24_and14_3_y0 ^ f_u_arrmul24_fa14_3_f_u_arrmul24_fa15_2_y2;
  assign f_u_arrmul24_fa14_3_y1 = f_u_arrmul24_fa14_3_f_u_arrmul24_and14_3_y0 & f_u_arrmul24_fa14_3_f_u_arrmul24_fa15_2_y2;
  assign f_u_arrmul24_fa14_3_y2 = f_u_arrmul24_fa14_3_y0 ^ f_u_arrmul24_fa14_3_f_u_arrmul24_fa13_3_y4;
  assign f_u_arrmul24_fa14_3_y3 = f_u_arrmul24_fa14_3_y0 & f_u_arrmul24_fa14_3_f_u_arrmul24_fa13_3_y4;
  assign f_u_arrmul24_fa14_3_y4 = f_u_arrmul24_fa14_3_y1 | f_u_arrmul24_fa14_3_y3;
  assign f_u_arrmul24_and15_3_a_15 = a_15;
  assign f_u_arrmul24_and15_3_b_3 = b_3;
  assign f_u_arrmul24_and15_3_y0 = f_u_arrmul24_and15_3_a_15 & f_u_arrmul24_and15_3_b_3;
  assign f_u_arrmul24_fa15_3_f_u_arrmul24_and15_3_y0 = f_u_arrmul24_and15_3_y0;
  assign f_u_arrmul24_fa15_3_f_u_arrmul24_fa16_2_y2 = f_u_arrmul24_fa16_2_y2;
  assign f_u_arrmul24_fa15_3_f_u_arrmul24_fa14_3_y4 = f_u_arrmul24_fa14_3_y4;
  assign f_u_arrmul24_fa15_3_y0 = f_u_arrmul24_fa15_3_f_u_arrmul24_and15_3_y0 ^ f_u_arrmul24_fa15_3_f_u_arrmul24_fa16_2_y2;
  assign f_u_arrmul24_fa15_3_y1 = f_u_arrmul24_fa15_3_f_u_arrmul24_and15_3_y0 & f_u_arrmul24_fa15_3_f_u_arrmul24_fa16_2_y2;
  assign f_u_arrmul24_fa15_3_y2 = f_u_arrmul24_fa15_3_y0 ^ f_u_arrmul24_fa15_3_f_u_arrmul24_fa14_3_y4;
  assign f_u_arrmul24_fa15_3_y3 = f_u_arrmul24_fa15_3_y0 & f_u_arrmul24_fa15_3_f_u_arrmul24_fa14_3_y4;
  assign f_u_arrmul24_fa15_3_y4 = f_u_arrmul24_fa15_3_y1 | f_u_arrmul24_fa15_3_y3;
  assign f_u_arrmul24_and16_3_a_16 = a_16;
  assign f_u_arrmul24_and16_3_b_3 = b_3;
  assign f_u_arrmul24_and16_3_y0 = f_u_arrmul24_and16_3_a_16 & f_u_arrmul24_and16_3_b_3;
  assign f_u_arrmul24_fa16_3_f_u_arrmul24_and16_3_y0 = f_u_arrmul24_and16_3_y0;
  assign f_u_arrmul24_fa16_3_f_u_arrmul24_fa17_2_y2 = f_u_arrmul24_fa17_2_y2;
  assign f_u_arrmul24_fa16_3_f_u_arrmul24_fa15_3_y4 = f_u_arrmul24_fa15_3_y4;
  assign f_u_arrmul24_fa16_3_y0 = f_u_arrmul24_fa16_3_f_u_arrmul24_and16_3_y0 ^ f_u_arrmul24_fa16_3_f_u_arrmul24_fa17_2_y2;
  assign f_u_arrmul24_fa16_3_y1 = f_u_arrmul24_fa16_3_f_u_arrmul24_and16_3_y0 & f_u_arrmul24_fa16_3_f_u_arrmul24_fa17_2_y2;
  assign f_u_arrmul24_fa16_3_y2 = f_u_arrmul24_fa16_3_y0 ^ f_u_arrmul24_fa16_3_f_u_arrmul24_fa15_3_y4;
  assign f_u_arrmul24_fa16_3_y3 = f_u_arrmul24_fa16_3_y0 & f_u_arrmul24_fa16_3_f_u_arrmul24_fa15_3_y4;
  assign f_u_arrmul24_fa16_3_y4 = f_u_arrmul24_fa16_3_y1 | f_u_arrmul24_fa16_3_y3;
  assign f_u_arrmul24_and17_3_a_17 = a_17;
  assign f_u_arrmul24_and17_3_b_3 = b_3;
  assign f_u_arrmul24_and17_3_y0 = f_u_arrmul24_and17_3_a_17 & f_u_arrmul24_and17_3_b_3;
  assign f_u_arrmul24_fa17_3_f_u_arrmul24_and17_3_y0 = f_u_arrmul24_and17_3_y0;
  assign f_u_arrmul24_fa17_3_f_u_arrmul24_fa18_2_y2 = f_u_arrmul24_fa18_2_y2;
  assign f_u_arrmul24_fa17_3_f_u_arrmul24_fa16_3_y4 = f_u_arrmul24_fa16_3_y4;
  assign f_u_arrmul24_fa17_3_y0 = f_u_arrmul24_fa17_3_f_u_arrmul24_and17_3_y0 ^ f_u_arrmul24_fa17_3_f_u_arrmul24_fa18_2_y2;
  assign f_u_arrmul24_fa17_3_y1 = f_u_arrmul24_fa17_3_f_u_arrmul24_and17_3_y0 & f_u_arrmul24_fa17_3_f_u_arrmul24_fa18_2_y2;
  assign f_u_arrmul24_fa17_3_y2 = f_u_arrmul24_fa17_3_y0 ^ f_u_arrmul24_fa17_3_f_u_arrmul24_fa16_3_y4;
  assign f_u_arrmul24_fa17_3_y3 = f_u_arrmul24_fa17_3_y0 & f_u_arrmul24_fa17_3_f_u_arrmul24_fa16_3_y4;
  assign f_u_arrmul24_fa17_3_y4 = f_u_arrmul24_fa17_3_y1 | f_u_arrmul24_fa17_3_y3;
  assign f_u_arrmul24_and18_3_a_18 = a_18;
  assign f_u_arrmul24_and18_3_b_3 = b_3;
  assign f_u_arrmul24_and18_3_y0 = f_u_arrmul24_and18_3_a_18 & f_u_arrmul24_and18_3_b_3;
  assign f_u_arrmul24_fa18_3_f_u_arrmul24_and18_3_y0 = f_u_arrmul24_and18_3_y0;
  assign f_u_arrmul24_fa18_3_f_u_arrmul24_fa19_2_y2 = f_u_arrmul24_fa19_2_y2;
  assign f_u_arrmul24_fa18_3_f_u_arrmul24_fa17_3_y4 = f_u_arrmul24_fa17_3_y4;
  assign f_u_arrmul24_fa18_3_y0 = f_u_arrmul24_fa18_3_f_u_arrmul24_and18_3_y0 ^ f_u_arrmul24_fa18_3_f_u_arrmul24_fa19_2_y2;
  assign f_u_arrmul24_fa18_3_y1 = f_u_arrmul24_fa18_3_f_u_arrmul24_and18_3_y0 & f_u_arrmul24_fa18_3_f_u_arrmul24_fa19_2_y2;
  assign f_u_arrmul24_fa18_3_y2 = f_u_arrmul24_fa18_3_y0 ^ f_u_arrmul24_fa18_3_f_u_arrmul24_fa17_3_y4;
  assign f_u_arrmul24_fa18_3_y3 = f_u_arrmul24_fa18_3_y0 & f_u_arrmul24_fa18_3_f_u_arrmul24_fa17_3_y4;
  assign f_u_arrmul24_fa18_3_y4 = f_u_arrmul24_fa18_3_y1 | f_u_arrmul24_fa18_3_y3;
  assign f_u_arrmul24_and19_3_a_19 = a_19;
  assign f_u_arrmul24_and19_3_b_3 = b_3;
  assign f_u_arrmul24_and19_3_y0 = f_u_arrmul24_and19_3_a_19 & f_u_arrmul24_and19_3_b_3;
  assign f_u_arrmul24_fa19_3_f_u_arrmul24_and19_3_y0 = f_u_arrmul24_and19_3_y0;
  assign f_u_arrmul24_fa19_3_f_u_arrmul24_fa20_2_y2 = f_u_arrmul24_fa20_2_y2;
  assign f_u_arrmul24_fa19_3_f_u_arrmul24_fa18_3_y4 = f_u_arrmul24_fa18_3_y4;
  assign f_u_arrmul24_fa19_3_y0 = f_u_arrmul24_fa19_3_f_u_arrmul24_and19_3_y0 ^ f_u_arrmul24_fa19_3_f_u_arrmul24_fa20_2_y2;
  assign f_u_arrmul24_fa19_3_y1 = f_u_arrmul24_fa19_3_f_u_arrmul24_and19_3_y0 & f_u_arrmul24_fa19_3_f_u_arrmul24_fa20_2_y2;
  assign f_u_arrmul24_fa19_3_y2 = f_u_arrmul24_fa19_3_y0 ^ f_u_arrmul24_fa19_3_f_u_arrmul24_fa18_3_y4;
  assign f_u_arrmul24_fa19_3_y3 = f_u_arrmul24_fa19_3_y0 & f_u_arrmul24_fa19_3_f_u_arrmul24_fa18_3_y4;
  assign f_u_arrmul24_fa19_3_y4 = f_u_arrmul24_fa19_3_y1 | f_u_arrmul24_fa19_3_y3;
  assign f_u_arrmul24_and20_3_a_20 = a_20;
  assign f_u_arrmul24_and20_3_b_3 = b_3;
  assign f_u_arrmul24_and20_3_y0 = f_u_arrmul24_and20_3_a_20 & f_u_arrmul24_and20_3_b_3;
  assign f_u_arrmul24_fa20_3_f_u_arrmul24_and20_3_y0 = f_u_arrmul24_and20_3_y0;
  assign f_u_arrmul24_fa20_3_f_u_arrmul24_fa21_2_y2 = f_u_arrmul24_fa21_2_y2;
  assign f_u_arrmul24_fa20_3_f_u_arrmul24_fa19_3_y4 = f_u_arrmul24_fa19_3_y4;
  assign f_u_arrmul24_fa20_3_y0 = f_u_arrmul24_fa20_3_f_u_arrmul24_and20_3_y0 ^ f_u_arrmul24_fa20_3_f_u_arrmul24_fa21_2_y2;
  assign f_u_arrmul24_fa20_3_y1 = f_u_arrmul24_fa20_3_f_u_arrmul24_and20_3_y0 & f_u_arrmul24_fa20_3_f_u_arrmul24_fa21_2_y2;
  assign f_u_arrmul24_fa20_3_y2 = f_u_arrmul24_fa20_3_y0 ^ f_u_arrmul24_fa20_3_f_u_arrmul24_fa19_3_y4;
  assign f_u_arrmul24_fa20_3_y3 = f_u_arrmul24_fa20_3_y0 & f_u_arrmul24_fa20_3_f_u_arrmul24_fa19_3_y4;
  assign f_u_arrmul24_fa20_3_y4 = f_u_arrmul24_fa20_3_y1 | f_u_arrmul24_fa20_3_y3;
  assign f_u_arrmul24_and21_3_a_21 = a_21;
  assign f_u_arrmul24_and21_3_b_3 = b_3;
  assign f_u_arrmul24_and21_3_y0 = f_u_arrmul24_and21_3_a_21 & f_u_arrmul24_and21_3_b_3;
  assign f_u_arrmul24_fa21_3_f_u_arrmul24_and21_3_y0 = f_u_arrmul24_and21_3_y0;
  assign f_u_arrmul24_fa21_3_f_u_arrmul24_fa22_2_y2 = f_u_arrmul24_fa22_2_y2;
  assign f_u_arrmul24_fa21_3_f_u_arrmul24_fa20_3_y4 = f_u_arrmul24_fa20_3_y4;
  assign f_u_arrmul24_fa21_3_y0 = f_u_arrmul24_fa21_3_f_u_arrmul24_and21_3_y0 ^ f_u_arrmul24_fa21_3_f_u_arrmul24_fa22_2_y2;
  assign f_u_arrmul24_fa21_3_y1 = f_u_arrmul24_fa21_3_f_u_arrmul24_and21_3_y0 & f_u_arrmul24_fa21_3_f_u_arrmul24_fa22_2_y2;
  assign f_u_arrmul24_fa21_3_y2 = f_u_arrmul24_fa21_3_y0 ^ f_u_arrmul24_fa21_3_f_u_arrmul24_fa20_3_y4;
  assign f_u_arrmul24_fa21_3_y3 = f_u_arrmul24_fa21_3_y0 & f_u_arrmul24_fa21_3_f_u_arrmul24_fa20_3_y4;
  assign f_u_arrmul24_fa21_3_y4 = f_u_arrmul24_fa21_3_y1 | f_u_arrmul24_fa21_3_y3;
  assign f_u_arrmul24_and22_3_a_22 = a_22;
  assign f_u_arrmul24_and22_3_b_3 = b_3;
  assign f_u_arrmul24_and22_3_y0 = f_u_arrmul24_and22_3_a_22 & f_u_arrmul24_and22_3_b_3;
  assign f_u_arrmul24_fa22_3_f_u_arrmul24_and22_3_y0 = f_u_arrmul24_and22_3_y0;
  assign f_u_arrmul24_fa22_3_f_u_arrmul24_fa23_2_y2 = f_u_arrmul24_fa23_2_y2;
  assign f_u_arrmul24_fa22_3_f_u_arrmul24_fa21_3_y4 = f_u_arrmul24_fa21_3_y4;
  assign f_u_arrmul24_fa22_3_y0 = f_u_arrmul24_fa22_3_f_u_arrmul24_and22_3_y0 ^ f_u_arrmul24_fa22_3_f_u_arrmul24_fa23_2_y2;
  assign f_u_arrmul24_fa22_3_y1 = f_u_arrmul24_fa22_3_f_u_arrmul24_and22_3_y0 & f_u_arrmul24_fa22_3_f_u_arrmul24_fa23_2_y2;
  assign f_u_arrmul24_fa22_3_y2 = f_u_arrmul24_fa22_3_y0 ^ f_u_arrmul24_fa22_3_f_u_arrmul24_fa21_3_y4;
  assign f_u_arrmul24_fa22_3_y3 = f_u_arrmul24_fa22_3_y0 & f_u_arrmul24_fa22_3_f_u_arrmul24_fa21_3_y4;
  assign f_u_arrmul24_fa22_3_y4 = f_u_arrmul24_fa22_3_y1 | f_u_arrmul24_fa22_3_y3;
  assign f_u_arrmul24_and23_3_a_23 = a_23;
  assign f_u_arrmul24_and23_3_b_3 = b_3;
  assign f_u_arrmul24_and23_3_y0 = f_u_arrmul24_and23_3_a_23 & f_u_arrmul24_and23_3_b_3;
  assign f_u_arrmul24_fa23_3_f_u_arrmul24_and23_3_y0 = f_u_arrmul24_and23_3_y0;
  assign f_u_arrmul24_fa23_3_f_u_arrmul24_fa23_2_y4 = f_u_arrmul24_fa23_2_y4;
  assign f_u_arrmul24_fa23_3_f_u_arrmul24_fa22_3_y4 = f_u_arrmul24_fa22_3_y4;
  assign f_u_arrmul24_fa23_3_y0 = f_u_arrmul24_fa23_3_f_u_arrmul24_and23_3_y0 ^ f_u_arrmul24_fa23_3_f_u_arrmul24_fa23_2_y4;
  assign f_u_arrmul24_fa23_3_y1 = f_u_arrmul24_fa23_3_f_u_arrmul24_and23_3_y0 & f_u_arrmul24_fa23_3_f_u_arrmul24_fa23_2_y4;
  assign f_u_arrmul24_fa23_3_y2 = f_u_arrmul24_fa23_3_y0 ^ f_u_arrmul24_fa23_3_f_u_arrmul24_fa22_3_y4;
  assign f_u_arrmul24_fa23_3_y3 = f_u_arrmul24_fa23_3_y0 & f_u_arrmul24_fa23_3_f_u_arrmul24_fa22_3_y4;
  assign f_u_arrmul24_fa23_3_y4 = f_u_arrmul24_fa23_3_y1 | f_u_arrmul24_fa23_3_y3;
  assign f_u_arrmul24_and0_4_a_0 = a_0;
  assign f_u_arrmul24_and0_4_b_4 = b_4;
  assign f_u_arrmul24_and0_4_y0 = f_u_arrmul24_and0_4_a_0 & f_u_arrmul24_and0_4_b_4;
  assign f_u_arrmul24_ha0_4_f_u_arrmul24_and0_4_y0 = f_u_arrmul24_and0_4_y0;
  assign f_u_arrmul24_ha0_4_f_u_arrmul24_fa1_3_y2 = f_u_arrmul24_fa1_3_y2;
  assign f_u_arrmul24_ha0_4_y0 = f_u_arrmul24_ha0_4_f_u_arrmul24_and0_4_y0 ^ f_u_arrmul24_ha0_4_f_u_arrmul24_fa1_3_y2;
  assign f_u_arrmul24_ha0_4_y1 = f_u_arrmul24_ha0_4_f_u_arrmul24_and0_4_y0 & f_u_arrmul24_ha0_4_f_u_arrmul24_fa1_3_y2;
  assign f_u_arrmul24_and1_4_a_1 = a_1;
  assign f_u_arrmul24_and1_4_b_4 = b_4;
  assign f_u_arrmul24_and1_4_y0 = f_u_arrmul24_and1_4_a_1 & f_u_arrmul24_and1_4_b_4;
  assign f_u_arrmul24_fa1_4_f_u_arrmul24_and1_4_y0 = f_u_arrmul24_and1_4_y0;
  assign f_u_arrmul24_fa1_4_f_u_arrmul24_fa2_3_y2 = f_u_arrmul24_fa2_3_y2;
  assign f_u_arrmul24_fa1_4_f_u_arrmul24_ha0_4_y1 = f_u_arrmul24_ha0_4_y1;
  assign f_u_arrmul24_fa1_4_y0 = f_u_arrmul24_fa1_4_f_u_arrmul24_and1_4_y0 ^ f_u_arrmul24_fa1_4_f_u_arrmul24_fa2_3_y2;
  assign f_u_arrmul24_fa1_4_y1 = f_u_arrmul24_fa1_4_f_u_arrmul24_and1_4_y0 & f_u_arrmul24_fa1_4_f_u_arrmul24_fa2_3_y2;
  assign f_u_arrmul24_fa1_4_y2 = f_u_arrmul24_fa1_4_y0 ^ f_u_arrmul24_fa1_4_f_u_arrmul24_ha0_4_y1;
  assign f_u_arrmul24_fa1_4_y3 = f_u_arrmul24_fa1_4_y0 & f_u_arrmul24_fa1_4_f_u_arrmul24_ha0_4_y1;
  assign f_u_arrmul24_fa1_4_y4 = f_u_arrmul24_fa1_4_y1 | f_u_arrmul24_fa1_4_y3;
  assign f_u_arrmul24_and2_4_a_2 = a_2;
  assign f_u_arrmul24_and2_4_b_4 = b_4;
  assign f_u_arrmul24_and2_4_y0 = f_u_arrmul24_and2_4_a_2 & f_u_arrmul24_and2_4_b_4;
  assign f_u_arrmul24_fa2_4_f_u_arrmul24_and2_4_y0 = f_u_arrmul24_and2_4_y0;
  assign f_u_arrmul24_fa2_4_f_u_arrmul24_fa3_3_y2 = f_u_arrmul24_fa3_3_y2;
  assign f_u_arrmul24_fa2_4_f_u_arrmul24_fa1_4_y4 = f_u_arrmul24_fa1_4_y4;
  assign f_u_arrmul24_fa2_4_y0 = f_u_arrmul24_fa2_4_f_u_arrmul24_and2_4_y0 ^ f_u_arrmul24_fa2_4_f_u_arrmul24_fa3_3_y2;
  assign f_u_arrmul24_fa2_4_y1 = f_u_arrmul24_fa2_4_f_u_arrmul24_and2_4_y0 & f_u_arrmul24_fa2_4_f_u_arrmul24_fa3_3_y2;
  assign f_u_arrmul24_fa2_4_y2 = f_u_arrmul24_fa2_4_y0 ^ f_u_arrmul24_fa2_4_f_u_arrmul24_fa1_4_y4;
  assign f_u_arrmul24_fa2_4_y3 = f_u_arrmul24_fa2_4_y0 & f_u_arrmul24_fa2_4_f_u_arrmul24_fa1_4_y4;
  assign f_u_arrmul24_fa2_4_y4 = f_u_arrmul24_fa2_4_y1 | f_u_arrmul24_fa2_4_y3;
  assign f_u_arrmul24_and3_4_a_3 = a_3;
  assign f_u_arrmul24_and3_4_b_4 = b_4;
  assign f_u_arrmul24_and3_4_y0 = f_u_arrmul24_and3_4_a_3 & f_u_arrmul24_and3_4_b_4;
  assign f_u_arrmul24_fa3_4_f_u_arrmul24_and3_4_y0 = f_u_arrmul24_and3_4_y0;
  assign f_u_arrmul24_fa3_4_f_u_arrmul24_fa4_3_y2 = f_u_arrmul24_fa4_3_y2;
  assign f_u_arrmul24_fa3_4_f_u_arrmul24_fa2_4_y4 = f_u_arrmul24_fa2_4_y4;
  assign f_u_arrmul24_fa3_4_y0 = f_u_arrmul24_fa3_4_f_u_arrmul24_and3_4_y0 ^ f_u_arrmul24_fa3_4_f_u_arrmul24_fa4_3_y2;
  assign f_u_arrmul24_fa3_4_y1 = f_u_arrmul24_fa3_4_f_u_arrmul24_and3_4_y0 & f_u_arrmul24_fa3_4_f_u_arrmul24_fa4_3_y2;
  assign f_u_arrmul24_fa3_4_y2 = f_u_arrmul24_fa3_4_y0 ^ f_u_arrmul24_fa3_4_f_u_arrmul24_fa2_4_y4;
  assign f_u_arrmul24_fa3_4_y3 = f_u_arrmul24_fa3_4_y0 & f_u_arrmul24_fa3_4_f_u_arrmul24_fa2_4_y4;
  assign f_u_arrmul24_fa3_4_y4 = f_u_arrmul24_fa3_4_y1 | f_u_arrmul24_fa3_4_y3;
  assign f_u_arrmul24_and4_4_a_4 = a_4;
  assign f_u_arrmul24_and4_4_b_4 = b_4;
  assign f_u_arrmul24_and4_4_y0 = f_u_arrmul24_and4_4_a_4 & f_u_arrmul24_and4_4_b_4;
  assign f_u_arrmul24_fa4_4_f_u_arrmul24_and4_4_y0 = f_u_arrmul24_and4_4_y0;
  assign f_u_arrmul24_fa4_4_f_u_arrmul24_fa5_3_y2 = f_u_arrmul24_fa5_3_y2;
  assign f_u_arrmul24_fa4_4_f_u_arrmul24_fa3_4_y4 = f_u_arrmul24_fa3_4_y4;
  assign f_u_arrmul24_fa4_4_y0 = f_u_arrmul24_fa4_4_f_u_arrmul24_and4_4_y0 ^ f_u_arrmul24_fa4_4_f_u_arrmul24_fa5_3_y2;
  assign f_u_arrmul24_fa4_4_y1 = f_u_arrmul24_fa4_4_f_u_arrmul24_and4_4_y0 & f_u_arrmul24_fa4_4_f_u_arrmul24_fa5_3_y2;
  assign f_u_arrmul24_fa4_4_y2 = f_u_arrmul24_fa4_4_y0 ^ f_u_arrmul24_fa4_4_f_u_arrmul24_fa3_4_y4;
  assign f_u_arrmul24_fa4_4_y3 = f_u_arrmul24_fa4_4_y0 & f_u_arrmul24_fa4_4_f_u_arrmul24_fa3_4_y4;
  assign f_u_arrmul24_fa4_4_y4 = f_u_arrmul24_fa4_4_y1 | f_u_arrmul24_fa4_4_y3;
  assign f_u_arrmul24_and5_4_a_5 = a_5;
  assign f_u_arrmul24_and5_4_b_4 = b_4;
  assign f_u_arrmul24_and5_4_y0 = f_u_arrmul24_and5_4_a_5 & f_u_arrmul24_and5_4_b_4;
  assign f_u_arrmul24_fa5_4_f_u_arrmul24_and5_4_y0 = f_u_arrmul24_and5_4_y0;
  assign f_u_arrmul24_fa5_4_f_u_arrmul24_fa6_3_y2 = f_u_arrmul24_fa6_3_y2;
  assign f_u_arrmul24_fa5_4_f_u_arrmul24_fa4_4_y4 = f_u_arrmul24_fa4_4_y4;
  assign f_u_arrmul24_fa5_4_y0 = f_u_arrmul24_fa5_4_f_u_arrmul24_and5_4_y0 ^ f_u_arrmul24_fa5_4_f_u_arrmul24_fa6_3_y2;
  assign f_u_arrmul24_fa5_4_y1 = f_u_arrmul24_fa5_4_f_u_arrmul24_and5_4_y0 & f_u_arrmul24_fa5_4_f_u_arrmul24_fa6_3_y2;
  assign f_u_arrmul24_fa5_4_y2 = f_u_arrmul24_fa5_4_y0 ^ f_u_arrmul24_fa5_4_f_u_arrmul24_fa4_4_y4;
  assign f_u_arrmul24_fa5_4_y3 = f_u_arrmul24_fa5_4_y0 & f_u_arrmul24_fa5_4_f_u_arrmul24_fa4_4_y4;
  assign f_u_arrmul24_fa5_4_y4 = f_u_arrmul24_fa5_4_y1 | f_u_arrmul24_fa5_4_y3;
  assign f_u_arrmul24_and6_4_a_6 = a_6;
  assign f_u_arrmul24_and6_4_b_4 = b_4;
  assign f_u_arrmul24_and6_4_y0 = f_u_arrmul24_and6_4_a_6 & f_u_arrmul24_and6_4_b_4;
  assign f_u_arrmul24_fa6_4_f_u_arrmul24_and6_4_y0 = f_u_arrmul24_and6_4_y0;
  assign f_u_arrmul24_fa6_4_f_u_arrmul24_fa7_3_y2 = f_u_arrmul24_fa7_3_y2;
  assign f_u_arrmul24_fa6_4_f_u_arrmul24_fa5_4_y4 = f_u_arrmul24_fa5_4_y4;
  assign f_u_arrmul24_fa6_4_y0 = f_u_arrmul24_fa6_4_f_u_arrmul24_and6_4_y0 ^ f_u_arrmul24_fa6_4_f_u_arrmul24_fa7_3_y2;
  assign f_u_arrmul24_fa6_4_y1 = f_u_arrmul24_fa6_4_f_u_arrmul24_and6_4_y0 & f_u_arrmul24_fa6_4_f_u_arrmul24_fa7_3_y2;
  assign f_u_arrmul24_fa6_4_y2 = f_u_arrmul24_fa6_4_y0 ^ f_u_arrmul24_fa6_4_f_u_arrmul24_fa5_4_y4;
  assign f_u_arrmul24_fa6_4_y3 = f_u_arrmul24_fa6_4_y0 & f_u_arrmul24_fa6_4_f_u_arrmul24_fa5_4_y4;
  assign f_u_arrmul24_fa6_4_y4 = f_u_arrmul24_fa6_4_y1 | f_u_arrmul24_fa6_4_y3;
  assign f_u_arrmul24_and7_4_a_7 = a_7;
  assign f_u_arrmul24_and7_4_b_4 = b_4;
  assign f_u_arrmul24_and7_4_y0 = f_u_arrmul24_and7_4_a_7 & f_u_arrmul24_and7_4_b_4;
  assign f_u_arrmul24_fa7_4_f_u_arrmul24_and7_4_y0 = f_u_arrmul24_and7_4_y0;
  assign f_u_arrmul24_fa7_4_f_u_arrmul24_fa8_3_y2 = f_u_arrmul24_fa8_3_y2;
  assign f_u_arrmul24_fa7_4_f_u_arrmul24_fa6_4_y4 = f_u_arrmul24_fa6_4_y4;
  assign f_u_arrmul24_fa7_4_y0 = f_u_arrmul24_fa7_4_f_u_arrmul24_and7_4_y0 ^ f_u_arrmul24_fa7_4_f_u_arrmul24_fa8_3_y2;
  assign f_u_arrmul24_fa7_4_y1 = f_u_arrmul24_fa7_4_f_u_arrmul24_and7_4_y0 & f_u_arrmul24_fa7_4_f_u_arrmul24_fa8_3_y2;
  assign f_u_arrmul24_fa7_4_y2 = f_u_arrmul24_fa7_4_y0 ^ f_u_arrmul24_fa7_4_f_u_arrmul24_fa6_4_y4;
  assign f_u_arrmul24_fa7_4_y3 = f_u_arrmul24_fa7_4_y0 & f_u_arrmul24_fa7_4_f_u_arrmul24_fa6_4_y4;
  assign f_u_arrmul24_fa7_4_y4 = f_u_arrmul24_fa7_4_y1 | f_u_arrmul24_fa7_4_y3;
  assign f_u_arrmul24_and8_4_a_8 = a_8;
  assign f_u_arrmul24_and8_4_b_4 = b_4;
  assign f_u_arrmul24_and8_4_y0 = f_u_arrmul24_and8_4_a_8 & f_u_arrmul24_and8_4_b_4;
  assign f_u_arrmul24_fa8_4_f_u_arrmul24_and8_4_y0 = f_u_arrmul24_and8_4_y0;
  assign f_u_arrmul24_fa8_4_f_u_arrmul24_fa9_3_y2 = f_u_arrmul24_fa9_3_y2;
  assign f_u_arrmul24_fa8_4_f_u_arrmul24_fa7_4_y4 = f_u_arrmul24_fa7_4_y4;
  assign f_u_arrmul24_fa8_4_y0 = f_u_arrmul24_fa8_4_f_u_arrmul24_and8_4_y0 ^ f_u_arrmul24_fa8_4_f_u_arrmul24_fa9_3_y2;
  assign f_u_arrmul24_fa8_4_y1 = f_u_arrmul24_fa8_4_f_u_arrmul24_and8_4_y0 & f_u_arrmul24_fa8_4_f_u_arrmul24_fa9_3_y2;
  assign f_u_arrmul24_fa8_4_y2 = f_u_arrmul24_fa8_4_y0 ^ f_u_arrmul24_fa8_4_f_u_arrmul24_fa7_4_y4;
  assign f_u_arrmul24_fa8_4_y3 = f_u_arrmul24_fa8_4_y0 & f_u_arrmul24_fa8_4_f_u_arrmul24_fa7_4_y4;
  assign f_u_arrmul24_fa8_4_y4 = f_u_arrmul24_fa8_4_y1 | f_u_arrmul24_fa8_4_y3;
  assign f_u_arrmul24_and9_4_a_9 = a_9;
  assign f_u_arrmul24_and9_4_b_4 = b_4;
  assign f_u_arrmul24_and9_4_y0 = f_u_arrmul24_and9_4_a_9 & f_u_arrmul24_and9_4_b_4;
  assign f_u_arrmul24_fa9_4_f_u_arrmul24_and9_4_y0 = f_u_arrmul24_and9_4_y0;
  assign f_u_arrmul24_fa9_4_f_u_arrmul24_fa10_3_y2 = f_u_arrmul24_fa10_3_y2;
  assign f_u_arrmul24_fa9_4_f_u_arrmul24_fa8_4_y4 = f_u_arrmul24_fa8_4_y4;
  assign f_u_arrmul24_fa9_4_y0 = f_u_arrmul24_fa9_4_f_u_arrmul24_and9_4_y0 ^ f_u_arrmul24_fa9_4_f_u_arrmul24_fa10_3_y2;
  assign f_u_arrmul24_fa9_4_y1 = f_u_arrmul24_fa9_4_f_u_arrmul24_and9_4_y0 & f_u_arrmul24_fa9_4_f_u_arrmul24_fa10_3_y2;
  assign f_u_arrmul24_fa9_4_y2 = f_u_arrmul24_fa9_4_y0 ^ f_u_arrmul24_fa9_4_f_u_arrmul24_fa8_4_y4;
  assign f_u_arrmul24_fa9_4_y3 = f_u_arrmul24_fa9_4_y0 & f_u_arrmul24_fa9_4_f_u_arrmul24_fa8_4_y4;
  assign f_u_arrmul24_fa9_4_y4 = f_u_arrmul24_fa9_4_y1 | f_u_arrmul24_fa9_4_y3;
  assign f_u_arrmul24_and10_4_a_10 = a_10;
  assign f_u_arrmul24_and10_4_b_4 = b_4;
  assign f_u_arrmul24_and10_4_y0 = f_u_arrmul24_and10_4_a_10 & f_u_arrmul24_and10_4_b_4;
  assign f_u_arrmul24_fa10_4_f_u_arrmul24_and10_4_y0 = f_u_arrmul24_and10_4_y0;
  assign f_u_arrmul24_fa10_4_f_u_arrmul24_fa11_3_y2 = f_u_arrmul24_fa11_3_y2;
  assign f_u_arrmul24_fa10_4_f_u_arrmul24_fa9_4_y4 = f_u_arrmul24_fa9_4_y4;
  assign f_u_arrmul24_fa10_4_y0 = f_u_arrmul24_fa10_4_f_u_arrmul24_and10_4_y0 ^ f_u_arrmul24_fa10_4_f_u_arrmul24_fa11_3_y2;
  assign f_u_arrmul24_fa10_4_y1 = f_u_arrmul24_fa10_4_f_u_arrmul24_and10_4_y0 & f_u_arrmul24_fa10_4_f_u_arrmul24_fa11_3_y2;
  assign f_u_arrmul24_fa10_4_y2 = f_u_arrmul24_fa10_4_y0 ^ f_u_arrmul24_fa10_4_f_u_arrmul24_fa9_4_y4;
  assign f_u_arrmul24_fa10_4_y3 = f_u_arrmul24_fa10_4_y0 & f_u_arrmul24_fa10_4_f_u_arrmul24_fa9_4_y4;
  assign f_u_arrmul24_fa10_4_y4 = f_u_arrmul24_fa10_4_y1 | f_u_arrmul24_fa10_4_y3;
  assign f_u_arrmul24_and11_4_a_11 = a_11;
  assign f_u_arrmul24_and11_4_b_4 = b_4;
  assign f_u_arrmul24_and11_4_y0 = f_u_arrmul24_and11_4_a_11 & f_u_arrmul24_and11_4_b_4;
  assign f_u_arrmul24_fa11_4_f_u_arrmul24_and11_4_y0 = f_u_arrmul24_and11_4_y0;
  assign f_u_arrmul24_fa11_4_f_u_arrmul24_fa12_3_y2 = f_u_arrmul24_fa12_3_y2;
  assign f_u_arrmul24_fa11_4_f_u_arrmul24_fa10_4_y4 = f_u_arrmul24_fa10_4_y4;
  assign f_u_arrmul24_fa11_4_y0 = f_u_arrmul24_fa11_4_f_u_arrmul24_and11_4_y0 ^ f_u_arrmul24_fa11_4_f_u_arrmul24_fa12_3_y2;
  assign f_u_arrmul24_fa11_4_y1 = f_u_arrmul24_fa11_4_f_u_arrmul24_and11_4_y0 & f_u_arrmul24_fa11_4_f_u_arrmul24_fa12_3_y2;
  assign f_u_arrmul24_fa11_4_y2 = f_u_arrmul24_fa11_4_y0 ^ f_u_arrmul24_fa11_4_f_u_arrmul24_fa10_4_y4;
  assign f_u_arrmul24_fa11_4_y3 = f_u_arrmul24_fa11_4_y0 & f_u_arrmul24_fa11_4_f_u_arrmul24_fa10_4_y4;
  assign f_u_arrmul24_fa11_4_y4 = f_u_arrmul24_fa11_4_y1 | f_u_arrmul24_fa11_4_y3;
  assign f_u_arrmul24_and12_4_a_12 = a_12;
  assign f_u_arrmul24_and12_4_b_4 = b_4;
  assign f_u_arrmul24_and12_4_y0 = f_u_arrmul24_and12_4_a_12 & f_u_arrmul24_and12_4_b_4;
  assign f_u_arrmul24_fa12_4_f_u_arrmul24_and12_4_y0 = f_u_arrmul24_and12_4_y0;
  assign f_u_arrmul24_fa12_4_f_u_arrmul24_fa13_3_y2 = f_u_arrmul24_fa13_3_y2;
  assign f_u_arrmul24_fa12_4_f_u_arrmul24_fa11_4_y4 = f_u_arrmul24_fa11_4_y4;
  assign f_u_arrmul24_fa12_4_y0 = f_u_arrmul24_fa12_4_f_u_arrmul24_and12_4_y0 ^ f_u_arrmul24_fa12_4_f_u_arrmul24_fa13_3_y2;
  assign f_u_arrmul24_fa12_4_y1 = f_u_arrmul24_fa12_4_f_u_arrmul24_and12_4_y0 & f_u_arrmul24_fa12_4_f_u_arrmul24_fa13_3_y2;
  assign f_u_arrmul24_fa12_4_y2 = f_u_arrmul24_fa12_4_y0 ^ f_u_arrmul24_fa12_4_f_u_arrmul24_fa11_4_y4;
  assign f_u_arrmul24_fa12_4_y3 = f_u_arrmul24_fa12_4_y0 & f_u_arrmul24_fa12_4_f_u_arrmul24_fa11_4_y4;
  assign f_u_arrmul24_fa12_4_y4 = f_u_arrmul24_fa12_4_y1 | f_u_arrmul24_fa12_4_y3;
  assign f_u_arrmul24_and13_4_a_13 = a_13;
  assign f_u_arrmul24_and13_4_b_4 = b_4;
  assign f_u_arrmul24_and13_4_y0 = f_u_arrmul24_and13_4_a_13 & f_u_arrmul24_and13_4_b_4;
  assign f_u_arrmul24_fa13_4_f_u_arrmul24_and13_4_y0 = f_u_arrmul24_and13_4_y0;
  assign f_u_arrmul24_fa13_4_f_u_arrmul24_fa14_3_y2 = f_u_arrmul24_fa14_3_y2;
  assign f_u_arrmul24_fa13_4_f_u_arrmul24_fa12_4_y4 = f_u_arrmul24_fa12_4_y4;
  assign f_u_arrmul24_fa13_4_y0 = f_u_arrmul24_fa13_4_f_u_arrmul24_and13_4_y0 ^ f_u_arrmul24_fa13_4_f_u_arrmul24_fa14_3_y2;
  assign f_u_arrmul24_fa13_4_y1 = f_u_arrmul24_fa13_4_f_u_arrmul24_and13_4_y0 & f_u_arrmul24_fa13_4_f_u_arrmul24_fa14_3_y2;
  assign f_u_arrmul24_fa13_4_y2 = f_u_arrmul24_fa13_4_y0 ^ f_u_arrmul24_fa13_4_f_u_arrmul24_fa12_4_y4;
  assign f_u_arrmul24_fa13_4_y3 = f_u_arrmul24_fa13_4_y0 & f_u_arrmul24_fa13_4_f_u_arrmul24_fa12_4_y4;
  assign f_u_arrmul24_fa13_4_y4 = f_u_arrmul24_fa13_4_y1 | f_u_arrmul24_fa13_4_y3;
  assign f_u_arrmul24_and14_4_a_14 = a_14;
  assign f_u_arrmul24_and14_4_b_4 = b_4;
  assign f_u_arrmul24_and14_4_y0 = f_u_arrmul24_and14_4_a_14 & f_u_arrmul24_and14_4_b_4;
  assign f_u_arrmul24_fa14_4_f_u_arrmul24_and14_4_y0 = f_u_arrmul24_and14_4_y0;
  assign f_u_arrmul24_fa14_4_f_u_arrmul24_fa15_3_y2 = f_u_arrmul24_fa15_3_y2;
  assign f_u_arrmul24_fa14_4_f_u_arrmul24_fa13_4_y4 = f_u_arrmul24_fa13_4_y4;
  assign f_u_arrmul24_fa14_4_y0 = f_u_arrmul24_fa14_4_f_u_arrmul24_and14_4_y0 ^ f_u_arrmul24_fa14_4_f_u_arrmul24_fa15_3_y2;
  assign f_u_arrmul24_fa14_4_y1 = f_u_arrmul24_fa14_4_f_u_arrmul24_and14_4_y0 & f_u_arrmul24_fa14_4_f_u_arrmul24_fa15_3_y2;
  assign f_u_arrmul24_fa14_4_y2 = f_u_arrmul24_fa14_4_y0 ^ f_u_arrmul24_fa14_4_f_u_arrmul24_fa13_4_y4;
  assign f_u_arrmul24_fa14_4_y3 = f_u_arrmul24_fa14_4_y0 & f_u_arrmul24_fa14_4_f_u_arrmul24_fa13_4_y4;
  assign f_u_arrmul24_fa14_4_y4 = f_u_arrmul24_fa14_4_y1 | f_u_arrmul24_fa14_4_y3;
  assign f_u_arrmul24_and15_4_a_15 = a_15;
  assign f_u_arrmul24_and15_4_b_4 = b_4;
  assign f_u_arrmul24_and15_4_y0 = f_u_arrmul24_and15_4_a_15 & f_u_arrmul24_and15_4_b_4;
  assign f_u_arrmul24_fa15_4_f_u_arrmul24_and15_4_y0 = f_u_arrmul24_and15_4_y0;
  assign f_u_arrmul24_fa15_4_f_u_arrmul24_fa16_3_y2 = f_u_arrmul24_fa16_3_y2;
  assign f_u_arrmul24_fa15_4_f_u_arrmul24_fa14_4_y4 = f_u_arrmul24_fa14_4_y4;
  assign f_u_arrmul24_fa15_4_y0 = f_u_arrmul24_fa15_4_f_u_arrmul24_and15_4_y0 ^ f_u_arrmul24_fa15_4_f_u_arrmul24_fa16_3_y2;
  assign f_u_arrmul24_fa15_4_y1 = f_u_arrmul24_fa15_4_f_u_arrmul24_and15_4_y0 & f_u_arrmul24_fa15_4_f_u_arrmul24_fa16_3_y2;
  assign f_u_arrmul24_fa15_4_y2 = f_u_arrmul24_fa15_4_y0 ^ f_u_arrmul24_fa15_4_f_u_arrmul24_fa14_4_y4;
  assign f_u_arrmul24_fa15_4_y3 = f_u_arrmul24_fa15_4_y0 & f_u_arrmul24_fa15_4_f_u_arrmul24_fa14_4_y4;
  assign f_u_arrmul24_fa15_4_y4 = f_u_arrmul24_fa15_4_y1 | f_u_arrmul24_fa15_4_y3;
  assign f_u_arrmul24_and16_4_a_16 = a_16;
  assign f_u_arrmul24_and16_4_b_4 = b_4;
  assign f_u_arrmul24_and16_4_y0 = f_u_arrmul24_and16_4_a_16 & f_u_arrmul24_and16_4_b_4;
  assign f_u_arrmul24_fa16_4_f_u_arrmul24_and16_4_y0 = f_u_arrmul24_and16_4_y0;
  assign f_u_arrmul24_fa16_4_f_u_arrmul24_fa17_3_y2 = f_u_arrmul24_fa17_3_y2;
  assign f_u_arrmul24_fa16_4_f_u_arrmul24_fa15_4_y4 = f_u_arrmul24_fa15_4_y4;
  assign f_u_arrmul24_fa16_4_y0 = f_u_arrmul24_fa16_4_f_u_arrmul24_and16_4_y0 ^ f_u_arrmul24_fa16_4_f_u_arrmul24_fa17_3_y2;
  assign f_u_arrmul24_fa16_4_y1 = f_u_arrmul24_fa16_4_f_u_arrmul24_and16_4_y0 & f_u_arrmul24_fa16_4_f_u_arrmul24_fa17_3_y2;
  assign f_u_arrmul24_fa16_4_y2 = f_u_arrmul24_fa16_4_y0 ^ f_u_arrmul24_fa16_4_f_u_arrmul24_fa15_4_y4;
  assign f_u_arrmul24_fa16_4_y3 = f_u_arrmul24_fa16_4_y0 & f_u_arrmul24_fa16_4_f_u_arrmul24_fa15_4_y4;
  assign f_u_arrmul24_fa16_4_y4 = f_u_arrmul24_fa16_4_y1 | f_u_arrmul24_fa16_4_y3;
  assign f_u_arrmul24_and17_4_a_17 = a_17;
  assign f_u_arrmul24_and17_4_b_4 = b_4;
  assign f_u_arrmul24_and17_4_y0 = f_u_arrmul24_and17_4_a_17 & f_u_arrmul24_and17_4_b_4;
  assign f_u_arrmul24_fa17_4_f_u_arrmul24_and17_4_y0 = f_u_arrmul24_and17_4_y0;
  assign f_u_arrmul24_fa17_4_f_u_arrmul24_fa18_3_y2 = f_u_arrmul24_fa18_3_y2;
  assign f_u_arrmul24_fa17_4_f_u_arrmul24_fa16_4_y4 = f_u_arrmul24_fa16_4_y4;
  assign f_u_arrmul24_fa17_4_y0 = f_u_arrmul24_fa17_4_f_u_arrmul24_and17_4_y0 ^ f_u_arrmul24_fa17_4_f_u_arrmul24_fa18_3_y2;
  assign f_u_arrmul24_fa17_4_y1 = f_u_arrmul24_fa17_4_f_u_arrmul24_and17_4_y0 & f_u_arrmul24_fa17_4_f_u_arrmul24_fa18_3_y2;
  assign f_u_arrmul24_fa17_4_y2 = f_u_arrmul24_fa17_4_y0 ^ f_u_arrmul24_fa17_4_f_u_arrmul24_fa16_4_y4;
  assign f_u_arrmul24_fa17_4_y3 = f_u_arrmul24_fa17_4_y0 & f_u_arrmul24_fa17_4_f_u_arrmul24_fa16_4_y4;
  assign f_u_arrmul24_fa17_4_y4 = f_u_arrmul24_fa17_4_y1 | f_u_arrmul24_fa17_4_y3;
  assign f_u_arrmul24_and18_4_a_18 = a_18;
  assign f_u_arrmul24_and18_4_b_4 = b_4;
  assign f_u_arrmul24_and18_4_y0 = f_u_arrmul24_and18_4_a_18 & f_u_arrmul24_and18_4_b_4;
  assign f_u_arrmul24_fa18_4_f_u_arrmul24_and18_4_y0 = f_u_arrmul24_and18_4_y0;
  assign f_u_arrmul24_fa18_4_f_u_arrmul24_fa19_3_y2 = f_u_arrmul24_fa19_3_y2;
  assign f_u_arrmul24_fa18_4_f_u_arrmul24_fa17_4_y4 = f_u_arrmul24_fa17_4_y4;
  assign f_u_arrmul24_fa18_4_y0 = f_u_arrmul24_fa18_4_f_u_arrmul24_and18_4_y0 ^ f_u_arrmul24_fa18_4_f_u_arrmul24_fa19_3_y2;
  assign f_u_arrmul24_fa18_4_y1 = f_u_arrmul24_fa18_4_f_u_arrmul24_and18_4_y0 & f_u_arrmul24_fa18_4_f_u_arrmul24_fa19_3_y2;
  assign f_u_arrmul24_fa18_4_y2 = f_u_arrmul24_fa18_4_y0 ^ f_u_arrmul24_fa18_4_f_u_arrmul24_fa17_4_y4;
  assign f_u_arrmul24_fa18_4_y3 = f_u_arrmul24_fa18_4_y0 & f_u_arrmul24_fa18_4_f_u_arrmul24_fa17_4_y4;
  assign f_u_arrmul24_fa18_4_y4 = f_u_arrmul24_fa18_4_y1 | f_u_arrmul24_fa18_4_y3;
  assign f_u_arrmul24_and19_4_a_19 = a_19;
  assign f_u_arrmul24_and19_4_b_4 = b_4;
  assign f_u_arrmul24_and19_4_y0 = f_u_arrmul24_and19_4_a_19 & f_u_arrmul24_and19_4_b_4;
  assign f_u_arrmul24_fa19_4_f_u_arrmul24_and19_4_y0 = f_u_arrmul24_and19_4_y0;
  assign f_u_arrmul24_fa19_4_f_u_arrmul24_fa20_3_y2 = f_u_arrmul24_fa20_3_y2;
  assign f_u_arrmul24_fa19_4_f_u_arrmul24_fa18_4_y4 = f_u_arrmul24_fa18_4_y4;
  assign f_u_arrmul24_fa19_4_y0 = f_u_arrmul24_fa19_4_f_u_arrmul24_and19_4_y0 ^ f_u_arrmul24_fa19_4_f_u_arrmul24_fa20_3_y2;
  assign f_u_arrmul24_fa19_4_y1 = f_u_arrmul24_fa19_4_f_u_arrmul24_and19_4_y0 & f_u_arrmul24_fa19_4_f_u_arrmul24_fa20_3_y2;
  assign f_u_arrmul24_fa19_4_y2 = f_u_arrmul24_fa19_4_y0 ^ f_u_arrmul24_fa19_4_f_u_arrmul24_fa18_4_y4;
  assign f_u_arrmul24_fa19_4_y3 = f_u_arrmul24_fa19_4_y0 & f_u_arrmul24_fa19_4_f_u_arrmul24_fa18_4_y4;
  assign f_u_arrmul24_fa19_4_y4 = f_u_arrmul24_fa19_4_y1 | f_u_arrmul24_fa19_4_y3;
  assign f_u_arrmul24_and20_4_a_20 = a_20;
  assign f_u_arrmul24_and20_4_b_4 = b_4;
  assign f_u_arrmul24_and20_4_y0 = f_u_arrmul24_and20_4_a_20 & f_u_arrmul24_and20_4_b_4;
  assign f_u_arrmul24_fa20_4_f_u_arrmul24_and20_4_y0 = f_u_arrmul24_and20_4_y0;
  assign f_u_arrmul24_fa20_4_f_u_arrmul24_fa21_3_y2 = f_u_arrmul24_fa21_3_y2;
  assign f_u_arrmul24_fa20_4_f_u_arrmul24_fa19_4_y4 = f_u_arrmul24_fa19_4_y4;
  assign f_u_arrmul24_fa20_4_y0 = f_u_arrmul24_fa20_4_f_u_arrmul24_and20_4_y0 ^ f_u_arrmul24_fa20_4_f_u_arrmul24_fa21_3_y2;
  assign f_u_arrmul24_fa20_4_y1 = f_u_arrmul24_fa20_4_f_u_arrmul24_and20_4_y0 & f_u_arrmul24_fa20_4_f_u_arrmul24_fa21_3_y2;
  assign f_u_arrmul24_fa20_4_y2 = f_u_arrmul24_fa20_4_y0 ^ f_u_arrmul24_fa20_4_f_u_arrmul24_fa19_4_y4;
  assign f_u_arrmul24_fa20_4_y3 = f_u_arrmul24_fa20_4_y0 & f_u_arrmul24_fa20_4_f_u_arrmul24_fa19_4_y4;
  assign f_u_arrmul24_fa20_4_y4 = f_u_arrmul24_fa20_4_y1 | f_u_arrmul24_fa20_4_y3;
  assign f_u_arrmul24_and21_4_a_21 = a_21;
  assign f_u_arrmul24_and21_4_b_4 = b_4;
  assign f_u_arrmul24_and21_4_y0 = f_u_arrmul24_and21_4_a_21 & f_u_arrmul24_and21_4_b_4;
  assign f_u_arrmul24_fa21_4_f_u_arrmul24_and21_4_y0 = f_u_arrmul24_and21_4_y0;
  assign f_u_arrmul24_fa21_4_f_u_arrmul24_fa22_3_y2 = f_u_arrmul24_fa22_3_y2;
  assign f_u_arrmul24_fa21_4_f_u_arrmul24_fa20_4_y4 = f_u_arrmul24_fa20_4_y4;
  assign f_u_arrmul24_fa21_4_y0 = f_u_arrmul24_fa21_4_f_u_arrmul24_and21_4_y0 ^ f_u_arrmul24_fa21_4_f_u_arrmul24_fa22_3_y2;
  assign f_u_arrmul24_fa21_4_y1 = f_u_arrmul24_fa21_4_f_u_arrmul24_and21_4_y0 & f_u_arrmul24_fa21_4_f_u_arrmul24_fa22_3_y2;
  assign f_u_arrmul24_fa21_4_y2 = f_u_arrmul24_fa21_4_y0 ^ f_u_arrmul24_fa21_4_f_u_arrmul24_fa20_4_y4;
  assign f_u_arrmul24_fa21_4_y3 = f_u_arrmul24_fa21_4_y0 & f_u_arrmul24_fa21_4_f_u_arrmul24_fa20_4_y4;
  assign f_u_arrmul24_fa21_4_y4 = f_u_arrmul24_fa21_4_y1 | f_u_arrmul24_fa21_4_y3;
  assign f_u_arrmul24_and22_4_a_22 = a_22;
  assign f_u_arrmul24_and22_4_b_4 = b_4;
  assign f_u_arrmul24_and22_4_y0 = f_u_arrmul24_and22_4_a_22 & f_u_arrmul24_and22_4_b_4;
  assign f_u_arrmul24_fa22_4_f_u_arrmul24_and22_4_y0 = f_u_arrmul24_and22_4_y0;
  assign f_u_arrmul24_fa22_4_f_u_arrmul24_fa23_3_y2 = f_u_arrmul24_fa23_3_y2;
  assign f_u_arrmul24_fa22_4_f_u_arrmul24_fa21_4_y4 = f_u_arrmul24_fa21_4_y4;
  assign f_u_arrmul24_fa22_4_y0 = f_u_arrmul24_fa22_4_f_u_arrmul24_and22_4_y0 ^ f_u_arrmul24_fa22_4_f_u_arrmul24_fa23_3_y2;
  assign f_u_arrmul24_fa22_4_y1 = f_u_arrmul24_fa22_4_f_u_arrmul24_and22_4_y0 & f_u_arrmul24_fa22_4_f_u_arrmul24_fa23_3_y2;
  assign f_u_arrmul24_fa22_4_y2 = f_u_arrmul24_fa22_4_y0 ^ f_u_arrmul24_fa22_4_f_u_arrmul24_fa21_4_y4;
  assign f_u_arrmul24_fa22_4_y3 = f_u_arrmul24_fa22_4_y0 & f_u_arrmul24_fa22_4_f_u_arrmul24_fa21_4_y4;
  assign f_u_arrmul24_fa22_4_y4 = f_u_arrmul24_fa22_4_y1 | f_u_arrmul24_fa22_4_y3;
  assign f_u_arrmul24_and23_4_a_23 = a_23;
  assign f_u_arrmul24_and23_4_b_4 = b_4;
  assign f_u_arrmul24_and23_4_y0 = f_u_arrmul24_and23_4_a_23 & f_u_arrmul24_and23_4_b_4;
  assign f_u_arrmul24_fa23_4_f_u_arrmul24_and23_4_y0 = f_u_arrmul24_and23_4_y0;
  assign f_u_arrmul24_fa23_4_f_u_arrmul24_fa23_3_y4 = f_u_arrmul24_fa23_3_y4;
  assign f_u_arrmul24_fa23_4_f_u_arrmul24_fa22_4_y4 = f_u_arrmul24_fa22_4_y4;
  assign f_u_arrmul24_fa23_4_y0 = f_u_arrmul24_fa23_4_f_u_arrmul24_and23_4_y0 ^ f_u_arrmul24_fa23_4_f_u_arrmul24_fa23_3_y4;
  assign f_u_arrmul24_fa23_4_y1 = f_u_arrmul24_fa23_4_f_u_arrmul24_and23_4_y0 & f_u_arrmul24_fa23_4_f_u_arrmul24_fa23_3_y4;
  assign f_u_arrmul24_fa23_4_y2 = f_u_arrmul24_fa23_4_y0 ^ f_u_arrmul24_fa23_4_f_u_arrmul24_fa22_4_y4;
  assign f_u_arrmul24_fa23_4_y3 = f_u_arrmul24_fa23_4_y0 & f_u_arrmul24_fa23_4_f_u_arrmul24_fa22_4_y4;
  assign f_u_arrmul24_fa23_4_y4 = f_u_arrmul24_fa23_4_y1 | f_u_arrmul24_fa23_4_y3;
  assign f_u_arrmul24_and0_5_a_0 = a_0;
  assign f_u_arrmul24_and0_5_b_5 = b_5;
  assign f_u_arrmul24_and0_5_y0 = f_u_arrmul24_and0_5_a_0 & f_u_arrmul24_and0_5_b_5;
  assign f_u_arrmul24_ha0_5_f_u_arrmul24_and0_5_y0 = f_u_arrmul24_and0_5_y0;
  assign f_u_arrmul24_ha0_5_f_u_arrmul24_fa1_4_y2 = f_u_arrmul24_fa1_4_y2;
  assign f_u_arrmul24_ha0_5_y0 = f_u_arrmul24_ha0_5_f_u_arrmul24_and0_5_y0 ^ f_u_arrmul24_ha0_5_f_u_arrmul24_fa1_4_y2;
  assign f_u_arrmul24_ha0_5_y1 = f_u_arrmul24_ha0_5_f_u_arrmul24_and0_5_y0 & f_u_arrmul24_ha0_5_f_u_arrmul24_fa1_4_y2;
  assign f_u_arrmul24_and1_5_a_1 = a_1;
  assign f_u_arrmul24_and1_5_b_5 = b_5;
  assign f_u_arrmul24_and1_5_y0 = f_u_arrmul24_and1_5_a_1 & f_u_arrmul24_and1_5_b_5;
  assign f_u_arrmul24_fa1_5_f_u_arrmul24_and1_5_y0 = f_u_arrmul24_and1_5_y0;
  assign f_u_arrmul24_fa1_5_f_u_arrmul24_fa2_4_y2 = f_u_arrmul24_fa2_4_y2;
  assign f_u_arrmul24_fa1_5_f_u_arrmul24_ha0_5_y1 = f_u_arrmul24_ha0_5_y1;
  assign f_u_arrmul24_fa1_5_y0 = f_u_arrmul24_fa1_5_f_u_arrmul24_and1_5_y0 ^ f_u_arrmul24_fa1_5_f_u_arrmul24_fa2_4_y2;
  assign f_u_arrmul24_fa1_5_y1 = f_u_arrmul24_fa1_5_f_u_arrmul24_and1_5_y0 & f_u_arrmul24_fa1_5_f_u_arrmul24_fa2_4_y2;
  assign f_u_arrmul24_fa1_5_y2 = f_u_arrmul24_fa1_5_y0 ^ f_u_arrmul24_fa1_5_f_u_arrmul24_ha0_5_y1;
  assign f_u_arrmul24_fa1_5_y3 = f_u_arrmul24_fa1_5_y0 & f_u_arrmul24_fa1_5_f_u_arrmul24_ha0_5_y1;
  assign f_u_arrmul24_fa1_5_y4 = f_u_arrmul24_fa1_5_y1 | f_u_arrmul24_fa1_5_y3;
  assign f_u_arrmul24_and2_5_a_2 = a_2;
  assign f_u_arrmul24_and2_5_b_5 = b_5;
  assign f_u_arrmul24_and2_5_y0 = f_u_arrmul24_and2_5_a_2 & f_u_arrmul24_and2_5_b_5;
  assign f_u_arrmul24_fa2_5_f_u_arrmul24_and2_5_y0 = f_u_arrmul24_and2_5_y0;
  assign f_u_arrmul24_fa2_5_f_u_arrmul24_fa3_4_y2 = f_u_arrmul24_fa3_4_y2;
  assign f_u_arrmul24_fa2_5_f_u_arrmul24_fa1_5_y4 = f_u_arrmul24_fa1_5_y4;
  assign f_u_arrmul24_fa2_5_y0 = f_u_arrmul24_fa2_5_f_u_arrmul24_and2_5_y0 ^ f_u_arrmul24_fa2_5_f_u_arrmul24_fa3_4_y2;
  assign f_u_arrmul24_fa2_5_y1 = f_u_arrmul24_fa2_5_f_u_arrmul24_and2_5_y0 & f_u_arrmul24_fa2_5_f_u_arrmul24_fa3_4_y2;
  assign f_u_arrmul24_fa2_5_y2 = f_u_arrmul24_fa2_5_y0 ^ f_u_arrmul24_fa2_5_f_u_arrmul24_fa1_5_y4;
  assign f_u_arrmul24_fa2_5_y3 = f_u_arrmul24_fa2_5_y0 & f_u_arrmul24_fa2_5_f_u_arrmul24_fa1_5_y4;
  assign f_u_arrmul24_fa2_5_y4 = f_u_arrmul24_fa2_5_y1 | f_u_arrmul24_fa2_5_y3;
  assign f_u_arrmul24_and3_5_a_3 = a_3;
  assign f_u_arrmul24_and3_5_b_5 = b_5;
  assign f_u_arrmul24_and3_5_y0 = f_u_arrmul24_and3_5_a_3 & f_u_arrmul24_and3_5_b_5;
  assign f_u_arrmul24_fa3_5_f_u_arrmul24_and3_5_y0 = f_u_arrmul24_and3_5_y0;
  assign f_u_arrmul24_fa3_5_f_u_arrmul24_fa4_4_y2 = f_u_arrmul24_fa4_4_y2;
  assign f_u_arrmul24_fa3_5_f_u_arrmul24_fa2_5_y4 = f_u_arrmul24_fa2_5_y4;
  assign f_u_arrmul24_fa3_5_y0 = f_u_arrmul24_fa3_5_f_u_arrmul24_and3_5_y0 ^ f_u_arrmul24_fa3_5_f_u_arrmul24_fa4_4_y2;
  assign f_u_arrmul24_fa3_5_y1 = f_u_arrmul24_fa3_5_f_u_arrmul24_and3_5_y0 & f_u_arrmul24_fa3_5_f_u_arrmul24_fa4_4_y2;
  assign f_u_arrmul24_fa3_5_y2 = f_u_arrmul24_fa3_5_y0 ^ f_u_arrmul24_fa3_5_f_u_arrmul24_fa2_5_y4;
  assign f_u_arrmul24_fa3_5_y3 = f_u_arrmul24_fa3_5_y0 & f_u_arrmul24_fa3_5_f_u_arrmul24_fa2_5_y4;
  assign f_u_arrmul24_fa3_5_y4 = f_u_arrmul24_fa3_5_y1 | f_u_arrmul24_fa3_5_y3;
  assign f_u_arrmul24_and4_5_a_4 = a_4;
  assign f_u_arrmul24_and4_5_b_5 = b_5;
  assign f_u_arrmul24_and4_5_y0 = f_u_arrmul24_and4_5_a_4 & f_u_arrmul24_and4_5_b_5;
  assign f_u_arrmul24_fa4_5_f_u_arrmul24_and4_5_y0 = f_u_arrmul24_and4_5_y0;
  assign f_u_arrmul24_fa4_5_f_u_arrmul24_fa5_4_y2 = f_u_arrmul24_fa5_4_y2;
  assign f_u_arrmul24_fa4_5_f_u_arrmul24_fa3_5_y4 = f_u_arrmul24_fa3_5_y4;
  assign f_u_arrmul24_fa4_5_y0 = f_u_arrmul24_fa4_5_f_u_arrmul24_and4_5_y0 ^ f_u_arrmul24_fa4_5_f_u_arrmul24_fa5_4_y2;
  assign f_u_arrmul24_fa4_5_y1 = f_u_arrmul24_fa4_5_f_u_arrmul24_and4_5_y0 & f_u_arrmul24_fa4_5_f_u_arrmul24_fa5_4_y2;
  assign f_u_arrmul24_fa4_5_y2 = f_u_arrmul24_fa4_5_y0 ^ f_u_arrmul24_fa4_5_f_u_arrmul24_fa3_5_y4;
  assign f_u_arrmul24_fa4_5_y3 = f_u_arrmul24_fa4_5_y0 & f_u_arrmul24_fa4_5_f_u_arrmul24_fa3_5_y4;
  assign f_u_arrmul24_fa4_5_y4 = f_u_arrmul24_fa4_5_y1 | f_u_arrmul24_fa4_5_y3;
  assign f_u_arrmul24_and5_5_a_5 = a_5;
  assign f_u_arrmul24_and5_5_b_5 = b_5;
  assign f_u_arrmul24_and5_5_y0 = f_u_arrmul24_and5_5_a_5 & f_u_arrmul24_and5_5_b_5;
  assign f_u_arrmul24_fa5_5_f_u_arrmul24_and5_5_y0 = f_u_arrmul24_and5_5_y0;
  assign f_u_arrmul24_fa5_5_f_u_arrmul24_fa6_4_y2 = f_u_arrmul24_fa6_4_y2;
  assign f_u_arrmul24_fa5_5_f_u_arrmul24_fa4_5_y4 = f_u_arrmul24_fa4_5_y4;
  assign f_u_arrmul24_fa5_5_y0 = f_u_arrmul24_fa5_5_f_u_arrmul24_and5_5_y0 ^ f_u_arrmul24_fa5_5_f_u_arrmul24_fa6_4_y2;
  assign f_u_arrmul24_fa5_5_y1 = f_u_arrmul24_fa5_5_f_u_arrmul24_and5_5_y0 & f_u_arrmul24_fa5_5_f_u_arrmul24_fa6_4_y2;
  assign f_u_arrmul24_fa5_5_y2 = f_u_arrmul24_fa5_5_y0 ^ f_u_arrmul24_fa5_5_f_u_arrmul24_fa4_5_y4;
  assign f_u_arrmul24_fa5_5_y3 = f_u_arrmul24_fa5_5_y0 & f_u_arrmul24_fa5_5_f_u_arrmul24_fa4_5_y4;
  assign f_u_arrmul24_fa5_5_y4 = f_u_arrmul24_fa5_5_y1 | f_u_arrmul24_fa5_5_y3;
  assign f_u_arrmul24_and6_5_a_6 = a_6;
  assign f_u_arrmul24_and6_5_b_5 = b_5;
  assign f_u_arrmul24_and6_5_y0 = f_u_arrmul24_and6_5_a_6 & f_u_arrmul24_and6_5_b_5;
  assign f_u_arrmul24_fa6_5_f_u_arrmul24_and6_5_y0 = f_u_arrmul24_and6_5_y0;
  assign f_u_arrmul24_fa6_5_f_u_arrmul24_fa7_4_y2 = f_u_arrmul24_fa7_4_y2;
  assign f_u_arrmul24_fa6_5_f_u_arrmul24_fa5_5_y4 = f_u_arrmul24_fa5_5_y4;
  assign f_u_arrmul24_fa6_5_y0 = f_u_arrmul24_fa6_5_f_u_arrmul24_and6_5_y0 ^ f_u_arrmul24_fa6_5_f_u_arrmul24_fa7_4_y2;
  assign f_u_arrmul24_fa6_5_y1 = f_u_arrmul24_fa6_5_f_u_arrmul24_and6_5_y0 & f_u_arrmul24_fa6_5_f_u_arrmul24_fa7_4_y2;
  assign f_u_arrmul24_fa6_5_y2 = f_u_arrmul24_fa6_5_y0 ^ f_u_arrmul24_fa6_5_f_u_arrmul24_fa5_5_y4;
  assign f_u_arrmul24_fa6_5_y3 = f_u_arrmul24_fa6_5_y0 & f_u_arrmul24_fa6_5_f_u_arrmul24_fa5_5_y4;
  assign f_u_arrmul24_fa6_5_y4 = f_u_arrmul24_fa6_5_y1 | f_u_arrmul24_fa6_5_y3;
  assign f_u_arrmul24_and7_5_a_7 = a_7;
  assign f_u_arrmul24_and7_5_b_5 = b_5;
  assign f_u_arrmul24_and7_5_y0 = f_u_arrmul24_and7_5_a_7 & f_u_arrmul24_and7_5_b_5;
  assign f_u_arrmul24_fa7_5_f_u_arrmul24_and7_5_y0 = f_u_arrmul24_and7_5_y0;
  assign f_u_arrmul24_fa7_5_f_u_arrmul24_fa8_4_y2 = f_u_arrmul24_fa8_4_y2;
  assign f_u_arrmul24_fa7_5_f_u_arrmul24_fa6_5_y4 = f_u_arrmul24_fa6_5_y4;
  assign f_u_arrmul24_fa7_5_y0 = f_u_arrmul24_fa7_5_f_u_arrmul24_and7_5_y0 ^ f_u_arrmul24_fa7_5_f_u_arrmul24_fa8_4_y2;
  assign f_u_arrmul24_fa7_5_y1 = f_u_arrmul24_fa7_5_f_u_arrmul24_and7_5_y0 & f_u_arrmul24_fa7_5_f_u_arrmul24_fa8_4_y2;
  assign f_u_arrmul24_fa7_5_y2 = f_u_arrmul24_fa7_5_y0 ^ f_u_arrmul24_fa7_5_f_u_arrmul24_fa6_5_y4;
  assign f_u_arrmul24_fa7_5_y3 = f_u_arrmul24_fa7_5_y0 & f_u_arrmul24_fa7_5_f_u_arrmul24_fa6_5_y4;
  assign f_u_arrmul24_fa7_5_y4 = f_u_arrmul24_fa7_5_y1 | f_u_arrmul24_fa7_5_y3;
  assign f_u_arrmul24_and8_5_a_8 = a_8;
  assign f_u_arrmul24_and8_5_b_5 = b_5;
  assign f_u_arrmul24_and8_5_y0 = f_u_arrmul24_and8_5_a_8 & f_u_arrmul24_and8_5_b_5;
  assign f_u_arrmul24_fa8_5_f_u_arrmul24_and8_5_y0 = f_u_arrmul24_and8_5_y0;
  assign f_u_arrmul24_fa8_5_f_u_arrmul24_fa9_4_y2 = f_u_arrmul24_fa9_4_y2;
  assign f_u_arrmul24_fa8_5_f_u_arrmul24_fa7_5_y4 = f_u_arrmul24_fa7_5_y4;
  assign f_u_arrmul24_fa8_5_y0 = f_u_arrmul24_fa8_5_f_u_arrmul24_and8_5_y0 ^ f_u_arrmul24_fa8_5_f_u_arrmul24_fa9_4_y2;
  assign f_u_arrmul24_fa8_5_y1 = f_u_arrmul24_fa8_5_f_u_arrmul24_and8_5_y0 & f_u_arrmul24_fa8_5_f_u_arrmul24_fa9_4_y2;
  assign f_u_arrmul24_fa8_5_y2 = f_u_arrmul24_fa8_5_y0 ^ f_u_arrmul24_fa8_5_f_u_arrmul24_fa7_5_y4;
  assign f_u_arrmul24_fa8_5_y3 = f_u_arrmul24_fa8_5_y0 & f_u_arrmul24_fa8_5_f_u_arrmul24_fa7_5_y4;
  assign f_u_arrmul24_fa8_5_y4 = f_u_arrmul24_fa8_5_y1 | f_u_arrmul24_fa8_5_y3;
  assign f_u_arrmul24_and9_5_a_9 = a_9;
  assign f_u_arrmul24_and9_5_b_5 = b_5;
  assign f_u_arrmul24_and9_5_y0 = f_u_arrmul24_and9_5_a_9 & f_u_arrmul24_and9_5_b_5;
  assign f_u_arrmul24_fa9_5_f_u_arrmul24_and9_5_y0 = f_u_arrmul24_and9_5_y0;
  assign f_u_arrmul24_fa9_5_f_u_arrmul24_fa10_4_y2 = f_u_arrmul24_fa10_4_y2;
  assign f_u_arrmul24_fa9_5_f_u_arrmul24_fa8_5_y4 = f_u_arrmul24_fa8_5_y4;
  assign f_u_arrmul24_fa9_5_y0 = f_u_arrmul24_fa9_5_f_u_arrmul24_and9_5_y0 ^ f_u_arrmul24_fa9_5_f_u_arrmul24_fa10_4_y2;
  assign f_u_arrmul24_fa9_5_y1 = f_u_arrmul24_fa9_5_f_u_arrmul24_and9_5_y0 & f_u_arrmul24_fa9_5_f_u_arrmul24_fa10_4_y2;
  assign f_u_arrmul24_fa9_5_y2 = f_u_arrmul24_fa9_5_y0 ^ f_u_arrmul24_fa9_5_f_u_arrmul24_fa8_5_y4;
  assign f_u_arrmul24_fa9_5_y3 = f_u_arrmul24_fa9_5_y0 & f_u_arrmul24_fa9_5_f_u_arrmul24_fa8_5_y4;
  assign f_u_arrmul24_fa9_5_y4 = f_u_arrmul24_fa9_5_y1 | f_u_arrmul24_fa9_5_y3;
  assign f_u_arrmul24_and10_5_a_10 = a_10;
  assign f_u_arrmul24_and10_5_b_5 = b_5;
  assign f_u_arrmul24_and10_5_y0 = f_u_arrmul24_and10_5_a_10 & f_u_arrmul24_and10_5_b_5;
  assign f_u_arrmul24_fa10_5_f_u_arrmul24_and10_5_y0 = f_u_arrmul24_and10_5_y0;
  assign f_u_arrmul24_fa10_5_f_u_arrmul24_fa11_4_y2 = f_u_arrmul24_fa11_4_y2;
  assign f_u_arrmul24_fa10_5_f_u_arrmul24_fa9_5_y4 = f_u_arrmul24_fa9_5_y4;
  assign f_u_arrmul24_fa10_5_y0 = f_u_arrmul24_fa10_5_f_u_arrmul24_and10_5_y0 ^ f_u_arrmul24_fa10_5_f_u_arrmul24_fa11_4_y2;
  assign f_u_arrmul24_fa10_5_y1 = f_u_arrmul24_fa10_5_f_u_arrmul24_and10_5_y0 & f_u_arrmul24_fa10_5_f_u_arrmul24_fa11_4_y2;
  assign f_u_arrmul24_fa10_5_y2 = f_u_arrmul24_fa10_5_y0 ^ f_u_arrmul24_fa10_5_f_u_arrmul24_fa9_5_y4;
  assign f_u_arrmul24_fa10_5_y3 = f_u_arrmul24_fa10_5_y0 & f_u_arrmul24_fa10_5_f_u_arrmul24_fa9_5_y4;
  assign f_u_arrmul24_fa10_5_y4 = f_u_arrmul24_fa10_5_y1 | f_u_arrmul24_fa10_5_y3;
  assign f_u_arrmul24_and11_5_a_11 = a_11;
  assign f_u_arrmul24_and11_5_b_5 = b_5;
  assign f_u_arrmul24_and11_5_y0 = f_u_arrmul24_and11_5_a_11 & f_u_arrmul24_and11_5_b_5;
  assign f_u_arrmul24_fa11_5_f_u_arrmul24_and11_5_y0 = f_u_arrmul24_and11_5_y0;
  assign f_u_arrmul24_fa11_5_f_u_arrmul24_fa12_4_y2 = f_u_arrmul24_fa12_4_y2;
  assign f_u_arrmul24_fa11_5_f_u_arrmul24_fa10_5_y4 = f_u_arrmul24_fa10_5_y4;
  assign f_u_arrmul24_fa11_5_y0 = f_u_arrmul24_fa11_5_f_u_arrmul24_and11_5_y0 ^ f_u_arrmul24_fa11_5_f_u_arrmul24_fa12_4_y2;
  assign f_u_arrmul24_fa11_5_y1 = f_u_arrmul24_fa11_5_f_u_arrmul24_and11_5_y0 & f_u_arrmul24_fa11_5_f_u_arrmul24_fa12_4_y2;
  assign f_u_arrmul24_fa11_5_y2 = f_u_arrmul24_fa11_5_y0 ^ f_u_arrmul24_fa11_5_f_u_arrmul24_fa10_5_y4;
  assign f_u_arrmul24_fa11_5_y3 = f_u_arrmul24_fa11_5_y0 & f_u_arrmul24_fa11_5_f_u_arrmul24_fa10_5_y4;
  assign f_u_arrmul24_fa11_5_y4 = f_u_arrmul24_fa11_5_y1 | f_u_arrmul24_fa11_5_y3;
  assign f_u_arrmul24_and12_5_a_12 = a_12;
  assign f_u_arrmul24_and12_5_b_5 = b_5;
  assign f_u_arrmul24_and12_5_y0 = f_u_arrmul24_and12_5_a_12 & f_u_arrmul24_and12_5_b_5;
  assign f_u_arrmul24_fa12_5_f_u_arrmul24_and12_5_y0 = f_u_arrmul24_and12_5_y0;
  assign f_u_arrmul24_fa12_5_f_u_arrmul24_fa13_4_y2 = f_u_arrmul24_fa13_4_y2;
  assign f_u_arrmul24_fa12_5_f_u_arrmul24_fa11_5_y4 = f_u_arrmul24_fa11_5_y4;
  assign f_u_arrmul24_fa12_5_y0 = f_u_arrmul24_fa12_5_f_u_arrmul24_and12_5_y0 ^ f_u_arrmul24_fa12_5_f_u_arrmul24_fa13_4_y2;
  assign f_u_arrmul24_fa12_5_y1 = f_u_arrmul24_fa12_5_f_u_arrmul24_and12_5_y0 & f_u_arrmul24_fa12_5_f_u_arrmul24_fa13_4_y2;
  assign f_u_arrmul24_fa12_5_y2 = f_u_arrmul24_fa12_5_y0 ^ f_u_arrmul24_fa12_5_f_u_arrmul24_fa11_5_y4;
  assign f_u_arrmul24_fa12_5_y3 = f_u_arrmul24_fa12_5_y0 & f_u_arrmul24_fa12_5_f_u_arrmul24_fa11_5_y4;
  assign f_u_arrmul24_fa12_5_y4 = f_u_arrmul24_fa12_5_y1 | f_u_arrmul24_fa12_5_y3;
  assign f_u_arrmul24_and13_5_a_13 = a_13;
  assign f_u_arrmul24_and13_5_b_5 = b_5;
  assign f_u_arrmul24_and13_5_y0 = f_u_arrmul24_and13_5_a_13 & f_u_arrmul24_and13_5_b_5;
  assign f_u_arrmul24_fa13_5_f_u_arrmul24_and13_5_y0 = f_u_arrmul24_and13_5_y0;
  assign f_u_arrmul24_fa13_5_f_u_arrmul24_fa14_4_y2 = f_u_arrmul24_fa14_4_y2;
  assign f_u_arrmul24_fa13_5_f_u_arrmul24_fa12_5_y4 = f_u_arrmul24_fa12_5_y4;
  assign f_u_arrmul24_fa13_5_y0 = f_u_arrmul24_fa13_5_f_u_arrmul24_and13_5_y0 ^ f_u_arrmul24_fa13_5_f_u_arrmul24_fa14_4_y2;
  assign f_u_arrmul24_fa13_5_y1 = f_u_arrmul24_fa13_5_f_u_arrmul24_and13_5_y0 & f_u_arrmul24_fa13_5_f_u_arrmul24_fa14_4_y2;
  assign f_u_arrmul24_fa13_5_y2 = f_u_arrmul24_fa13_5_y0 ^ f_u_arrmul24_fa13_5_f_u_arrmul24_fa12_5_y4;
  assign f_u_arrmul24_fa13_5_y3 = f_u_arrmul24_fa13_5_y0 & f_u_arrmul24_fa13_5_f_u_arrmul24_fa12_5_y4;
  assign f_u_arrmul24_fa13_5_y4 = f_u_arrmul24_fa13_5_y1 | f_u_arrmul24_fa13_5_y3;
  assign f_u_arrmul24_and14_5_a_14 = a_14;
  assign f_u_arrmul24_and14_5_b_5 = b_5;
  assign f_u_arrmul24_and14_5_y0 = f_u_arrmul24_and14_5_a_14 & f_u_arrmul24_and14_5_b_5;
  assign f_u_arrmul24_fa14_5_f_u_arrmul24_and14_5_y0 = f_u_arrmul24_and14_5_y0;
  assign f_u_arrmul24_fa14_5_f_u_arrmul24_fa15_4_y2 = f_u_arrmul24_fa15_4_y2;
  assign f_u_arrmul24_fa14_5_f_u_arrmul24_fa13_5_y4 = f_u_arrmul24_fa13_5_y4;
  assign f_u_arrmul24_fa14_5_y0 = f_u_arrmul24_fa14_5_f_u_arrmul24_and14_5_y0 ^ f_u_arrmul24_fa14_5_f_u_arrmul24_fa15_4_y2;
  assign f_u_arrmul24_fa14_5_y1 = f_u_arrmul24_fa14_5_f_u_arrmul24_and14_5_y0 & f_u_arrmul24_fa14_5_f_u_arrmul24_fa15_4_y2;
  assign f_u_arrmul24_fa14_5_y2 = f_u_arrmul24_fa14_5_y0 ^ f_u_arrmul24_fa14_5_f_u_arrmul24_fa13_5_y4;
  assign f_u_arrmul24_fa14_5_y3 = f_u_arrmul24_fa14_5_y0 & f_u_arrmul24_fa14_5_f_u_arrmul24_fa13_5_y4;
  assign f_u_arrmul24_fa14_5_y4 = f_u_arrmul24_fa14_5_y1 | f_u_arrmul24_fa14_5_y3;
  assign f_u_arrmul24_and15_5_a_15 = a_15;
  assign f_u_arrmul24_and15_5_b_5 = b_5;
  assign f_u_arrmul24_and15_5_y0 = f_u_arrmul24_and15_5_a_15 & f_u_arrmul24_and15_5_b_5;
  assign f_u_arrmul24_fa15_5_f_u_arrmul24_and15_5_y0 = f_u_arrmul24_and15_5_y0;
  assign f_u_arrmul24_fa15_5_f_u_arrmul24_fa16_4_y2 = f_u_arrmul24_fa16_4_y2;
  assign f_u_arrmul24_fa15_5_f_u_arrmul24_fa14_5_y4 = f_u_arrmul24_fa14_5_y4;
  assign f_u_arrmul24_fa15_5_y0 = f_u_arrmul24_fa15_5_f_u_arrmul24_and15_5_y0 ^ f_u_arrmul24_fa15_5_f_u_arrmul24_fa16_4_y2;
  assign f_u_arrmul24_fa15_5_y1 = f_u_arrmul24_fa15_5_f_u_arrmul24_and15_5_y0 & f_u_arrmul24_fa15_5_f_u_arrmul24_fa16_4_y2;
  assign f_u_arrmul24_fa15_5_y2 = f_u_arrmul24_fa15_5_y0 ^ f_u_arrmul24_fa15_5_f_u_arrmul24_fa14_5_y4;
  assign f_u_arrmul24_fa15_5_y3 = f_u_arrmul24_fa15_5_y0 & f_u_arrmul24_fa15_5_f_u_arrmul24_fa14_5_y4;
  assign f_u_arrmul24_fa15_5_y4 = f_u_arrmul24_fa15_5_y1 | f_u_arrmul24_fa15_5_y3;
  assign f_u_arrmul24_and16_5_a_16 = a_16;
  assign f_u_arrmul24_and16_5_b_5 = b_5;
  assign f_u_arrmul24_and16_5_y0 = f_u_arrmul24_and16_5_a_16 & f_u_arrmul24_and16_5_b_5;
  assign f_u_arrmul24_fa16_5_f_u_arrmul24_and16_5_y0 = f_u_arrmul24_and16_5_y0;
  assign f_u_arrmul24_fa16_5_f_u_arrmul24_fa17_4_y2 = f_u_arrmul24_fa17_4_y2;
  assign f_u_arrmul24_fa16_5_f_u_arrmul24_fa15_5_y4 = f_u_arrmul24_fa15_5_y4;
  assign f_u_arrmul24_fa16_5_y0 = f_u_arrmul24_fa16_5_f_u_arrmul24_and16_5_y0 ^ f_u_arrmul24_fa16_5_f_u_arrmul24_fa17_4_y2;
  assign f_u_arrmul24_fa16_5_y1 = f_u_arrmul24_fa16_5_f_u_arrmul24_and16_5_y0 & f_u_arrmul24_fa16_5_f_u_arrmul24_fa17_4_y2;
  assign f_u_arrmul24_fa16_5_y2 = f_u_arrmul24_fa16_5_y0 ^ f_u_arrmul24_fa16_5_f_u_arrmul24_fa15_5_y4;
  assign f_u_arrmul24_fa16_5_y3 = f_u_arrmul24_fa16_5_y0 & f_u_arrmul24_fa16_5_f_u_arrmul24_fa15_5_y4;
  assign f_u_arrmul24_fa16_5_y4 = f_u_arrmul24_fa16_5_y1 | f_u_arrmul24_fa16_5_y3;
  assign f_u_arrmul24_and17_5_a_17 = a_17;
  assign f_u_arrmul24_and17_5_b_5 = b_5;
  assign f_u_arrmul24_and17_5_y0 = f_u_arrmul24_and17_5_a_17 & f_u_arrmul24_and17_5_b_5;
  assign f_u_arrmul24_fa17_5_f_u_arrmul24_and17_5_y0 = f_u_arrmul24_and17_5_y0;
  assign f_u_arrmul24_fa17_5_f_u_arrmul24_fa18_4_y2 = f_u_arrmul24_fa18_4_y2;
  assign f_u_arrmul24_fa17_5_f_u_arrmul24_fa16_5_y4 = f_u_arrmul24_fa16_5_y4;
  assign f_u_arrmul24_fa17_5_y0 = f_u_arrmul24_fa17_5_f_u_arrmul24_and17_5_y0 ^ f_u_arrmul24_fa17_5_f_u_arrmul24_fa18_4_y2;
  assign f_u_arrmul24_fa17_5_y1 = f_u_arrmul24_fa17_5_f_u_arrmul24_and17_5_y0 & f_u_arrmul24_fa17_5_f_u_arrmul24_fa18_4_y2;
  assign f_u_arrmul24_fa17_5_y2 = f_u_arrmul24_fa17_5_y0 ^ f_u_arrmul24_fa17_5_f_u_arrmul24_fa16_5_y4;
  assign f_u_arrmul24_fa17_5_y3 = f_u_arrmul24_fa17_5_y0 & f_u_arrmul24_fa17_5_f_u_arrmul24_fa16_5_y4;
  assign f_u_arrmul24_fa17_5_y4 = f_u_arrmul24_fa17_5_y1 | f_u_arrmul24_fa17_5_y3;
  assign f_u_arrmul24_and18_5_a_18 = a_18;
  assign f_u_arrmul24_and18_5_b_5 = b_5;
  assign f_u_arrmul24_and18_5_y0 = f_u_arrmul24_and18_5_a_18 & f_u_arrmul24_and18_5_b_5;
  assign f_u_arrmul24_fa18_5_f_u_arrmul24_and18_5_y0 = f_u_arrmul24_and18_5_y0;
  assign f_u_arrmul24_fa18_5_f_u_arrmul24_fa19_4_y2 = f_u_arrmul24_fa19_4_y2;
  assign f_u_arrmul24_fa18_5_f_u_arrmul24_fa17_5_y4 = f_u_arrmul24_fa17_5_y4;
  assign f_u_arrmul24_fa18_5_y0 = f_u_arrmul24_fa18_5_f_u_arrmul24_and18_5_y0 ^ f_u_arrmul24_fa18_5_f_u_arrmul24_fa19_4_y2;
  assign f_u_arrmul24_fa18_5_y1 = f_u_arrmul24_fa18_5_f_u_arrmul24_and18_5_y0 & f_u_arrmul24_fa18_5_f_u_arrmul24_fa19_4_y2;
  assign f_u_arrmul24_fa18_5_y2 = f_u_arrmul24_fa18_5_y0 ^ f_u_arrmul24_fa18_5_f_u_arrmul24_fa17_5_y4;
  assign f_u_arrmul24_fa18_5_y3 = f_u_arrmul24_fa18_5_y0 & f_u_arrmul24_fa18_5_f_u_arrmul24_fa17_5_y4;
  assign f_u_arrmul24_fa18_5_y4 = f_u_arrmul24_fa18_5_y1 | f_u_arrmul24_fa18_5_y3;
  assign f_u_arrmul24_and19_5_a_19 = a_19;
  assign f_u_arrmul24_and19_5_b_5 = b_5;
  assign f_u_arrmul24_and19_5_y0 = f_u_arrmul24_and19_5_a_19 & f_u_arrmul24_and19_5_b_5;
  assign f_u_arrmul24_fa19_5_f_u_arrmul24_and19_5_y0 = f_u_arrmul24_and19_5_y0;
  assign f_u_arrmul24_fa19_5_f_u_arrmul24_fa20_4_y2 = f_u_arrmul24_fa20_4_y2;
  assign f_u_arrmul24_fa19_5_f_u_arrmul24_fa18_5_y4 = f_u_arrmul24_fa18_5_y4;
  assign f_u_arrmul24_fa19_5_y0 = f_u_arrmul24_fa19_5_f_u_arrmul24_and19_5_y0 ^ f_u_arrmul24_fa19_5_f_u_arrmul24_fa20_4_y2;
  assign f_u_arrmul24_fa19_5_y1 = f_u_arrmul24_fa19_5_f_u_arrmul24_and19_5_y0 & f_u_arrmul24_fa19_5_f_u_arrmul24_fa20_4_y2;
  assign f_u_arrmul24_fa19_5_y2 = f_u_arrmul24_fa19_5_y0 ^ f_u_arrmul24_fa19_5_f_u_arrmul24_fa18_5_y4;
  assign f_u_arrmul24_fa19_5_y3 = f_u_arrmul24_fa19_5_y0 & f_u_arrmul24_fa19_5_f_u_arrmul24_fa18_5_y4;
  assign f_u_arrmul24_fa19_5_y4 = f_u_arrmul24_fa19_5_y1 | f_u_arrmul24_fa19_5_y3;
  assign f_u_arrmul24_and20_5_a_20 = a_20;
  assign f_u_arrmul24_and20_5_b_5 = b_5;
  assign f_u_arrmul24_and20_5_y0 = f_u_arrmul24_and20_5_a_20 & f_u_arrmul24_and20_5_b_5;
  assign f_u_arrmul24_fa20_5_f_u_arrmul24_and20_5_y0 = f_u_arrmul24_and20_5_y0;
  assign f_u_arrmul24_fa20_5_f_u_arrmul24_fa21_4_y2 = f_u_arrmul24_fa21_4_y2;
  assign f_u_arrmul24_fa20_5_f_u_arrmul24_fa19_5_y4 = f_u_arrmul24_fa19_5_y4;
  assign f_u_arrmul24_fa20_5_y0 = f_u_arrmul24_fa20_5_f_u_arrmul24_and20_5_y0 ^ f_u_arrmul24_fa20_5_f_u_arrmul24_fa21_4_y2;
  assign f_u_arrmul24_fa20_5_y1 = f_u_arrmul24_fa20_5_f_u_arrmul24_and20_5_y0 & f_u_arrmul24_fa20_5_f_u_arrmul24_fa21_4_y2;
  assign f_u_arrmul24_fa20_5_y2 = f_u_arrmul24_fa20_5_y0 ^ f_u_arrmul24_fa20_5_f_u_arrmul24_fa19_5_y4;
  assign f_u_arrmul24_fa20_5_y3 = f_u_arrmul24_fa20_5_y0 & f_u_arrmul24_fa20_5_f_u_arrmul24_fa19_5_y4;
  assign f_u_arrmul24_fa20_5_y4 = f_u_arrmul24_fa20_5_y1 | f_u_arrmul24_fa20_5_y3;
  assign f_u_arrmul24_and21_5_a_21 = a_21;
  assign f_u_arrmul24_and21_5_b_5 = b_5;
  assign f_u_arrmul24_and21_5_y0 = f_u_arrmul24_and21_5_a_21 & f_u_arrmul24_and21_5_b_5;
  assign f_u_arrmul24_fa21_5_f_u_arrmul24_and21_5_y0 = f_u_arrmul24_and21_5_y0;
  assign f_u_arrmul24_fa21_5_f_u_arrmul24_fa22_4_y2 = f_u_arrmul24_fa22_4_y2;
  assign f_u_arrmul24_fa21_5_f_u_arrmul24_fa20_5_y4 = f_u_arrmul24_fa20_5_y4;
  assign f_u_arrmul24_fa21_5_y0 = f_u_arrmul24_fa21_5_f_u_arrmul24_and21_5_y0 ^ f_u_arrmul24_fa21_5_f_u_arrmul24_fa22_4_y2;
  assign f_u_arrmul24_fa21_5_y1 = f_u_arrmul24_fa21_5_f_u_arrmul24_and21_5_y0 & f_u_arrmul24_fa21_5_f_u_arrmul24_fa22_4_y2;
  assign f_u_arrmul24_fa21_5_y2 = f_u_arrmul24_fa21_5_y0 ^ f_u_arrmul24_fa21_5_f_u_arrmul24_fa20_5_y4;
  assign f_u_arrmul24_fa21_5_y3 = f_u_arrmul24_fa21_5_y0 & f_u_arrmul24_fa21_5_f_u_arrmul24_fa20_5_y4;
  assign f_u_arrmul24_fa21_5_y4 = f_u_arrmul24_fa21_5_y1 | f_u_arrmul24_fa21_5_y3;
  assign f_u_arrmul24_and22_5_a_22 = a_22;
  assign f_u_arrmul24_and22_5_b_5 = b_5;
  assign f_u_arrmul24_and22_5_y0 = f_u_arrmul24_and22_5_a_22 & f_u_arrmul24_and22_5_b_5;
  assign f_u_arrmul24_fa22_5_f_u_arrmul24_and22_5_y0 = f_u_arrmul24_and22_5_y0;
  assign f_u_arrmul24_fa22_5_f_u_arrmul24_fa23_4_y2 = f_u_arrmul24_fa23_4_y2;
  assign f_u_arrmul24_fa22_5_f_u_arrmul24_fa21_5_y4 = f_u_arrmul24_fa21_5_y4;
  assign f_u_arrmul24_fa22_5_y0 = f_u_arrmul24_fa22_5_f_u_arrmul24_and22_5_y0 ^ f_u_arrmul24_fa22_5_f_u_arrmul24_fa23_4_y2;
  assign f_u_arrmul24_fa22_5_y1 = f_u_arrmul24_fa22_5_f_u_arrmul24_and22_5_y0 & f_u_arrmul24_fa22_5_f_u_arrmul24_fa23_4_y2;
  assign f_u_arrmul24_fa22_5_y2 = f_u_arrmul24_fa22_5_y0 ^ f_u_arrmul24_fa22_5_f_u_arrmul24_fa21_5_y4;
  assign f_u_arrmul24_fa22_5_y3 = f_u_arrmul24_fa22_5_y0 & f_u_arrmul24_fa22_5_f_u_arrmul24_fa21_5_y4;
  assign f_u_arrmul24_fa22_5_y4 = f_u_arrmul24_fa22_5_y1 | f_u_arrmul24_fa22_5_y3;
  assign f_u_arrmul24_and23_5_a_23 = a_23;
  assign f_u_arrmul24_and23_5_b_5 = b_5;
  assign f_u_arrmul24_and23_5_y0 = f_u_arrmul24_and23_5_a_23 & f_u_arrmul24_and23_5_b_5;
  assign f_u_arrmul24_fa23_5_f_u_arrmul24_and23_5_y0 = f_u_arrmul24_and23_5_y0;
  assign f_u_arrmul24_fa23_5_f_u_arrmul24_fa23_4_y4 = f_u_arrmul24_fa23_4_y4;
  assign f_u_arrmul24_fa23_5_f_u_arrmul24_fa22_5_y4 = f_u_arrmul24_fa22_5_y4;
  assign f_u_arrmul24_fa23_5_y0 = f_u_arrmul24_fa23_5_f_u_arrmul24_and23_5_y0 ^ f_u_arrmul24_fa23_5_f_u_arrmul24_fa23_4_y4;
  assign f_u_arrmul24_fa23_5_y1 = f_u_arrmul24_fa23_5_f_u_arrmul24_and23_5_y0 & f_u_arrmul24_fa23_5_f_u_arrmul24_fa23_4_y4;
  assign f_u_arrmul24_fa23_5_y2 = f_u_arrmul24_fa23_5_y0 ^ f_u_arrmul24_fa23_5_f_u_arrmul24_fa22_5_y4;
  assign f_u_arrmul24_fa23_5_y3 = f_u_arrmul24_fa23_5_y0 & f_u_arrmul24_fa23_5_f_u_arrmul24_fa22_5_y4;
  assign f_u_arrmul24_fa23_5_y4 = f_u_arrmul24_fa23_5_y1 | f_u_arrmul24_fa23_5_y3;
  assign f_u_arrmul24_and0_6_a_0 = a_0;
  assign f_u_arrmul24_and0_6_b_6 = b_6;
  assign f_u_arrmul24_and0_6_y0 = f_u_arrmul24_and0_6_a_0 & f_u_arrmul24_and0_6_b_6;
  assign f_u_arrmul24_ha0_6_f_u_arrmul24_and0_6_y0 = f_u_arrmul24_and0_6_y0;
  assign f_u_arrmul24_ha0_6_f_u_arrmul24_fa1_5_y2 = f_u_arrmul24_fa1_5_y2;
  assign f_u_arrmul24_ha0_6_y0 = f_u_arrmul24_ha0_6_f_u_arrmul24_and0_6_y0 ^ f_u_arrmul24_ha0_6_f_u_arrmul24_fa1_5_y2;
  assign f_u_arrmul24_ha0_6_y1 = f_u_arrmul24_ha0_6_f_u_arrmul24_and0_6_y0 & f_u_arrmul24_ha0_6_f_u_arrmul24_fa1_5_y2;
  assign f_u_arrmul24_and1_6_a_1 = a_1;
  assign f_u_arrmul24_and1_6_b_6 = b_6;
  assign f_u_arrmul24_and1_6_y0 = f_u_arrmul24_and1_6_a_1 & f_u_arrmul24_and1_6_b_6;
  assign f_u_arrmul24_fa1_6_f_u_arrmul24_and1_6_y0 = f_u_arrmul24_and1_6_y0;
  assign f_u_arrmul24_fa1_6_f_u_arrmul24_fa2_5_y2 = f_u_arrmul24_fa2_5_y2;
  assign f_u_arrmul24_fa1_6_f_u_arrmul24_ha0_6_y1 = f_u_arrmul24_ha0_6_y1;
  assign f_u_arrmul24_fa1_6_y0 = f_u_arrmul24_fa1_6_f_u_arrmul24_and1_6_y0 ^ f_u_arrmul24_fa1_6_f_u_arrmul24_fa2_5_y2;
  assign f_u_arrmul24_fa1_6_y1 = f_u_arrmul24_fa1_6_f_u_arrmul24_and1_6_y0 & f_u_arrmul24_fa1_6_f_u_arrmul24_fa2_5_y2;
  assign f_u_arrmul24_fa1_6_y2 = f_u_arrmul24_fa1_6_y0 ^ f_u_arrmul24_fa1_6_f_u_arrmul24_ha0_6_y1;
  assign f_u_arrmul24_fa1_6_y3 = f_u_arrmul24_fa1_6_y0 & f_u_arrmul24_fa1_6_f_u_arrmul24_ha0_6_y1;
  assign f_u_arrmul24_fa1_6_y4 = f_u_arrmul24_fa1_6_y1 | f_u_arrmul24_fa1_6_y3;
  assign f_u_arrmul24_and2_6_a_2 = a_2;
  assign f_u_arrmul24_and2_6_b_6 = b_6;
  assign f_u_arrmul24_and2_6_y0 = f_u_arrmul24_and2_6_a_2 & f_u_arrmul24_and2_6_b_6;
  assign f_u_arrmul24_fa2_6_f_u_arrmul24_and2_6_y0 = f_u_arrmul24_and2_6_y0;
  assign f_u_arrmul24_fa2_6_f_u_arrmul24_fa3_5_y2 = f_u_arrmul24_fa3_5_y2;
  assign f_u_arrmul24_fa2_6_f_u_arrmul24_fa1_6_y4 = f_u_arrmul24_fa1_6_y4;
  assign f_u_arrmul24_fa2_6_y0 = f_u_arrmul24_fa2_6_f_u_arrmul24_and2_6_y0 ^ f_u_arrmul24_fa2_6_f_u_arrmul24_fa3_5_y2;
  assign f_u_arrmul24_fa2_6_y1 = f_u_arrmul24_fa2_6_f_u_arrmul24_and2_6_y0 & f_u_arrmul24_fa2_6_f_u_arrmul24_fa3_5_y2;
  assign f_u_arrmul24_fa2_6_y2 = f_u_arrmul24_fa2_6_y0 ^ f_u_arrmul24_fa2_6_f_u_arrmul24_fa1_6_y4;
  assign f_u_arrmul24_fa2_6_y3 = f_u_arrmul24_fa2_6_y0 & f_u_arrmul24_fa2_6_f_u_arrmul24_fa1_6_y4;
  assign f_u_arrmul24_fa2_6_y4 = f_u_arrmul24_fa2_6_y1 | f_u_arrmul24_fa2_6_y3;
  assign f_u_arrmul24_and3_6_a_3 = a_3;
  assign f_u_arrmul24_and3_6_b_6 = b_6;
  assign f_u_arrmul24_and3_6_y0 = f_u_arrmul24_and3_6_a_3 & f_u_arrmul24_and3_6_b_6;
  assign f_u_arrmul24_fa3_6_f_u_arrmul24_and3_6_y0 = f_u_arrmul24_and3_6_y0;
  assign f_u_arrmul24_fa3_6_f_u_arrmul24_fa4_5_y2 = f_u_arrmul24_fa4_5_y2;
  assign f_u_arrmul24_fa3_6_f_u_arrmul24_fa2_6_y4 = f_u_arrmul24_fa2_6_y4;
  assign f_u_arrmul24_fa3_6_y0 = f_u_arrmul24_fa3_6_f_u_arrmul24_and3_6_y0 ^ f_u_arrmul24_fa3_6_f_u_arrmul24_fa4_5_y2;
  assign f_u_arrmul24_fa3_6_y1 = f_u_arrmul24_fa3_6_f_u_arrmul24_and3_6_y0 & f_u_arrmul24_fa3_6_f_u_arrmul24_fa4_5_y2;
  assign f_u_arrmul24_fa3_6_y2 = f_u_arrmul24_fa3_6_y0 ^ f_u_arrmul24_fa3_6_f_u_arrmul24_fa2_6_y4;
  assign f_u_arrmul24_fa3_6_y3 = f_u_arrmul24_fa3_6_y0 & f_u_arrmul24_fa3_6_f_u_arrmul24_fa2_6_y4;
  assign f_u_arrmul24_fa3_6_y4 = f_u_arrmul24_fa3_6_y1 | f_u_arrmul24_fa3_6_y3;
  assign f_u_arrmul24_and4_6_a_4 = a_4;
  assign f_u_arrmul24_and4_6_b_6 = b_6;
  assign f_u_arrmul24_and4_6_y0 = f_u_arrmul24_and4_6_a_4 & f_u_arrmul24_and4_6_b_6;
  assign f_u_arrmul24_fa4_6_f_u_arrmul24_and4_6_y0 = f_u_arrmul24_and4_6_y0;
  assign f_u_arrmul24_fa4_6_f_u_arrmul24_fa5_5_y2 = f_u_arrmul24_fa5_5_y2;
  assign f_u_arrmul24_fa4_6_f_u_arrmul24_fa3_6_y4 = f_u_arrmul24_fa3_6_y4;
  assign f_u_arrmul24_fa4_6_y0 = f_u_arrmul24_fa4_6_f_u_arrmul24_and4_6_y0 ^ f_u_arrmul24_fa4_6_f_u_arrmul24_fa5_5_y2;
  assign f_u_arrmul24_fa4_6_y1 = f_u_arrmul24_fa4_6_f_u_arrmul24_and4_6_y0 & f_u_arrmul24_fa4_6_f_u_arrmul24_fa5_5_y2;
  assign f_u_arrmul24_fa4_6_y2 = f_u_arrmul24_fa4_6_y0 ^ f_u_arrmul24_fa4_6_f_u_arrmul24_fa3_6_y4;
  assign f_u_arrmul24_fa4_6_y3 = f_u_arrmul24_fa4_6_y0 & f_u_arrmul24_fa4_6_f_u_arrmul24_fa3_6_y4;
  assign f_u_arrmul24_fa4_6_y4 = f_u_arrmul24_fa4_6_y1 | f_u_arrmul24_fa4_6_y3;
  assign f_u_arrmul24_and5_6_a_5 = a_5;
  assign f_u_arrmul24_and5_6_b_6 = b_6;
  assign f_u_arrmul24_and5_6_y0 = f_u_arrmul24_and5_6_a_5 & f_u_arrmul24_and5_6_b_6;
  assign f_u_arrmul24_fa5_6_f_u_arrmul24_and5_6_y0 = f_u_arrmul24_and5_6_y0;
  assign f_u_arrmul24_fa5_6_f_u_arrmul24_fa6_5_y2 = f_u_arrmul24_fa6_5_y2;
  assign f_u_arrmul24_fa5_6_f_u_arrmul24_fa4_6_y4 = f_u_arrmul24_fa4_6_y4;
  assign f_u_arrmul24_fa5_6_y0 = f_u_arrmul24_fa5_6_f_u_arrmul24_and5_6_y0 ^ f_u_arrmul24_fa5_6_f_u_arrmul24_fa6_5_y2;
  assign f_u_arrmul24_fa5_6_y1 = f_u_arrmul24_fa5_6_f_u_arrmul24_and5_6_y0 & f_u_arrmul24_fa5_6_f_u_arrmul24_fa6_5_y2;
  assign f_u_arrmul24_fa5_6_y2 = f_u_arrmul24_fa5_6_y0 ^ f_u_arrmul24_fa5_6_f_u_arrmul24_fa4_6_y4;
  assign f_u_arrmul24_fa5_6_y3 = f_u_arrmul24_fa5_6_y0 & f_u_arrmul24_fa5_6_f_u_arrmul24_fa4_6_y4;
  assign f_u_arrmul24_fa5_6_y4 = f_u_arrmul24_fa5_6_y1 | f_u_arrmul24_fa5_6_y3;
  assign f_u_arrmul24_and6_6_a_6 = a_6;
  assign f_u_arrmul24_and6_6_b_6 = b_6;
  assign f_u_arrmul24_and6_6_y0 = f_u_arrmul24_and6_6_a_6 & f_u_arrmul24_and6_6_b_6;
  assign f_u_arrmul24_fa6_6_f_u_arrmul24_and6_6_y0 = f_u_arrmul24_and6_6_y0;
  assign f_u_arrmul24_fa6_6_f_u_arrmul24_fa7_5_y2 = f_u_arrmul24_fa7_5_y2;
  assign f_u_arrmul24_fa6_6_f_u_arrmul24_fa5_6_y4 = f_u_arrmul24_fa5_6_y4;
  assign f_u_arrmul24_fa6_6_y0 = f_u_arrmul24_fa6_6_f_u_arrmul24_and6_6_y0 ^ f_u_arrmul24_fa6_6_f_u_arrmul24_fa7_5_y2;
  assign f_u_arrmul24_fa6_6_y1 = f_u_arrmul24_fa6_6_f_u_arrmul24_and6_6_y0 & f_u_arrmul24_fa6_6_f_u_arrmul24_fa7_5_y2;
  assign f_u_arrmul24_fa6_6_y2 = f_u_arrmul24_fa6_6_y0 ^ f_u_arrmul24_fa6_6_f_u_arrmul24_fa5_6_y4;
  assign f_u_arrmul24_fa6_6_y3 = f_u_arrmul24_fa6_6_y0 & f_u_arrmul24_fa6_6_f_u_arrmul24_fa5_6_y4;
  assign f_u_arrmul24_fa6_6_y4 = f_u_arrmul24_fa6_6_y1 | f_u_arrmul24_fa6_6_y3;
  assign f_u_arrmul24_and7_6_a_7 = a_7;
  assign f_u_arrmul24_and7_6_b_6 = b_6;
  assign f_u_arrmul24_and7_6_y0 = f_u_arrmul24_and7_6_a_7 & f_u_arrmul24_and7_6_b_6;
  assign f_u_arrmul24_fa7_6_f_u_arrmul24_and7_6_y0 = f_u_arrmul24_and7_6_y0;
  assign f_u_arrmul24_fa7_6_f_u_arrmul24_fa8_5_y2 = f_u_arrmul24_fa8_5_y2;
  assign f_u_arrmul24_fa7_6_f_u_arrmul24_fa6_6_y4 = f_u_arrmul24_fa6_6_y4;
  assign f_u_arrmul24_fa7_6_y0 = f_u_arrmul24_fa7_6_f_u_arrmul24_and7_6_y0 ^ f_u_arrmul24_fa7_6_f_u_arrmul24_fa8_5_y2;
  assign f_u_arrmul24_fa7_6_y1 = f_u_arrmul24_fa7_6_f_u_arrmul24_and7_6_y0 & f_u_arrmul24_fa7_6_f_u_arrmul24_fa8_5_y2;
  assign f_u_arrmul24_fa7_6_y2 = f_u_arrmul24_fa7_6_y0 ^ f_u_arrmul24_fa7_6_f_u_arrmul24_fa6_6_y4;
  assign f_u_arrmul24_fa7_6_y3 = f_u_arrmul24_fa7_6_y0 & f_u_arrmul24_fa7_6_f_u_arrmul24_fa6_6_y4;
  assign f_u_arrmul24_fa7_6_y4 = f_u_arrmul24_fa7_6_y1 | f_u_arrmul24_fa7_6_y3;
  assign f_u_arrmul24_and8_6_a_8 = a_8;
  assign f_u_arrmul24_and8_6_b_6 = b_6;
  assign f_u_arrmul24_and8_6_y0 = f_u_arrmul24_and8_6_a_8 & f_u_arrmul24_and8_6_b_6;
  assign f_u_arrmul24_fa8_6_f_u_arrmul24_and8_6_y0 = f_u_arrmul24_and8_6_y0;
  assign f_u_arrmul24_fa8_6_f_u_arrmul24_fa9_5_y2 = f_u_arrmul24_fa9_5_y2;
  assign f_u_arrmul24_fa8_6_f_u_arrmul24_fa7_6_y4 = f_u_arrmul24_fa7_6_y4;
  assign f_u_arrmul24_fa8_6_y0 = f_u_arrmul24_fa8_6_f_u_arrmul24_and8_6_y0 ^ f_u_arrmul24_fa8_6_f_u_arrmul24_fa9_5_y2;
  assign f_u_arrmul24_fa8_6_y1 = f_u_arrmul24_fa8_6_f_u_arrmul24_and8_6_y0 & f_u_arrmul24_fa8_6_f_u_arrmul24_fa9_5_y2;
  assign f_u_arrmul24_fa8_6_y2 = f_u_arrmul24_fa8_6_y0 ^ f_u_arrmul24_fa8_6_f_u_arrmul24_fa7_6_y4;
  assign f_u_arrmul24_fa8_6_y3 = f_u_arrmul24_fa8_6_y0 & f_u_arrmul24_fa8_6_f_u_arrmul24_fa7_6_y4;
  assign f_u_arrmul24_fa8_6_y4 = f_u_arrmul24_fa8_6_y1 | f_u_arrmul24_fa8_6_y3;
  assign f_u_arrmul24_and9_6_a_9 = a_9;
  assign f_u_arrmul24_and9_6_b_6 = b_6;
  assign f_u_arrmul24_and9_6_y0 = f_u_arrmul24_and9_6_a_9 & f_u_arrmul24_and9_6_b_6;
  assign f_u_arrmul24_fa9_6_f_u_arrmul24_and9_6_y0 = f_u_arrmul24_and9_6_y0;
  assign f_u_arrmul24_fa9_6_f_u_arrmul24_fa10_5_y2 = f_u_arrmul24_fa10_5_y2;
  assign f_u_arrmul24_fa9_6_f_u_arrmul24_fa8_6_y4 = f_u_arrmul24_fa8_6_y4;
  assign f_u_arrmul24_fa9_6_y0 = f_u_arrmul24_fa9_6_f_u_arrmul24_and9_6_y0 ^ f_u_arrmul24_fa9_6_f_u_arrmul24_fa10_5_y2;
  assign f_u_arrmul24_fa9_6_y1 = f_u_arrmul24_fa9_6_f_u_arrmul24_and9_6_y0 & f_u_arrmul24_fa9_6_f_u_arrmul24_fa10_5_y2;
  assign f_u_arrmul24_fa9_6_y2 = f_u_arrmul24_fa9_6_y0 ^ f_u_arrmul24_fa9_6_f_u_arrmul24_fa8_6_y4;
  assign f_u_arrmul24_fa9_6_y3 = f_u_arrmul24_fa9_6_y0 & f_u_arrmul24_fa9_6_f_u_arrmul24_fa8_6_y4;
  assign f_u_arrmul24_fa9_6_y4 = f_u_arrmul24_fa9_6_y1 | f_u_arrmul24_fa9_6_y3;
  assign f_u_arrmul24_and10_6_a_10 = a_10;
  assign f_u_arrmul24_and10_6_b_6 = b_6;
  assign f_u_arrmul24_and10_6_y0 = f_u_arrmul24_and10_6_a_10 & f_u_arrmul24_and10_6_b_6;
  assign f_u_arrmul24_fa10_6_f_u_arrmul24_and10_6_y0 = f_u_arrmul24_and10_6_y0;
  assign f_u_arrmul24_fa10_6_f_u_arrmul24_fa11_5_y2 = f_u_arrmul24_fa11_5_y2;
  assign f_u_arrmul24_fa10_6_f_u_arrmul24_fa9_6_y4 = f_u_arrmul24_fa9_6_y4;
  assign f_u_arrmul24_fa10_6_y0 = f_u_arrmul24_fa10_6_f_u_arrmul24_and10_6_y0 ^ f_u_arrmul24_fa10_6_f_u_arrmul24_fa11_5_y2;
  assign f_u_arrmul24_fa10_6_y1 = f_u_arrmul24_fa10_6_f_u_arrmul24_and10_6_y0 & f_u_arrmul24_fa10_6_f_u_arrmul24_fa11_5_y2;
  assign f_u_arrmul24_fa10_6_y2 = f_u_arrmul24_fa10_6_y0 ^ f_u_arrmul24_fa10_6_f_u_arrmul24_fa9_6_y4;
  assign f_u_arrmul24_fa10_6_y3 = f_u_arrmul24_fa10_6_y0 & f_u_arrmul24_fa10_6_f_u_arrmul24_fa9_6_y4;
  assign f_u_arrmul24_fa10_6_y4 = f_u_arrmul24_fa10_6_y1 | f_u_arrmul24_fa10_6_y3;
  assign f_u_arrmul24_and11_6_a_11 = a_11;
  assign f_u_arrmul24_and11_6_b_6 = b_6;
  assign f_u_arrmul24_and11_6_y0 = f_u_arrmul24_and11_6_a_11 & f_u_arrmul24_and11_6_b_6;
  assign f_u_arrmul24_fa11_6_f_u_arrmul24_and11_6_y0 = f_u_arrmul24_and11_6_y0;
  assign f_u_arrmul24_fa11_6_f_u_arrmul24_fa12_5_y2 = f_u_arrmul24_fa12_5_y2;
  assign f_u_arrmul24_fa11_6_f_u_arrmul24_fa10_6_y4 = f_u_arrmul24_fa10_6_y4;
  assign f_u_arrmul24_fa11_6_y0 = f_u_arrmul24_fa11_6_f_u_arrmul24_and11_6_y0 ^ f_u_arrmul24_fa11_6_f_u_arrmul24_fa12_5_y2;
  assign f_u_arrmul24_fa11_6_y1 = f_u_arrmul24_fa11_6_f_u_arrmul24_and11_6_y0 & f_u_arrmul24_fa11_6_f_u_arrmul24_fa12_5_y2;
  assign f_u_arrmul24_fa11_6_y2 = f_u_arrmul24_fa11_6_y0 ^ f_u_arrmul24_fa11_6_f_u_arrmul24_fa10_6_y4;
  assign f_u_arrmul24_fa11_6_y3 = f_u_arrmul24_fa11_6_y0 & f_u_arrmul24_fa11_6_f_u_arrmul24_fa10_6_y4;
  assign f_u_arrmul24_fa11_6_y4 = f_u_arrmul24_fa11_6_y1 | f_u_arrmul24_fa11_6_y3;
  assign f_u_arrmul24_and12_6_a_12 = a_12;
  assign f_u_arrmul24_and12_6_b_6 = b_6;
  assign f_u_arrmul24_and12_6_y0 = f_u_arrmul24_and12_6_a_12 & f_u_arrmul24_and12_6_b_6;
  assign f_u_arrmul24_fa12_6_f_u_arrmul24_and12_6_y0 = f_u_arrmul24_and12_6_y0;
  assign f_u_arrmul24_fa12_6_f_u_arrmul24_fa13_5_y2 = f_u_arrmul24_fa13_5_y2;
  assign f_u_arrmul24_fa12_6_f_u_arrmul24_fa11_6_y4 = f_u_arrmul24_fa11_6_y4;
  assign f_u_arrmul24_fa12_6_y0 = f_u_arrmul24_fa12_6_f_u_arrmul24_and12_6_y0 ^ f_u_arrmul24_fa12_6_f_u_arrmul24_fa13_5_y2;
  assign f_u_arrmul24_fa12_6_y1 = f_u_arrmul24_fa12_6_f_u_arrmul24_and12_6_y0 & f_u_arrmul24_fa12_6_f_u_arrmul24_fa13_5_y2;
  assign f_u_arrmul24_fa12_6_y2 = f_u_arrmul24_fa12_6_y0 ^ f_u_arrmul24_fa12_6_f_u_arrmul24_fa11_6_y4;
  assign f_u_arrmul24_fa12_6_y3 = f_u_arrmul24_fa12_6_y0 & f_u_arrmul24_fa12_6_f_u_arrmul24_fa11_6_y4;
  assign f_u_arrmul24_fa12_6_y4 = f_u_arrmul24_fa12_6_y1 | f_u_arrmul24_fa12_6_y3;
  assign f_u_arrmul24_and13_6_a_13 = a_13;
  assign f_u_arrmul24_and13_6_b_6 = b_6;
  assign f_u_arrmul24_and13_6_y0 = f_u_arrmul24_and13_6_a_13 & f_u_arrmul24_and13_6_b_6;
  assign f_u_arrmul24_fa13_6_f_u_arrmul24_and13_6_y0 = f_u_arrmul24_and13_6_y0;
  assign f_u_arrmul24_fa13_6_f_u_arrmul24_fa14_5_y2 = f_u_arrmul24_fa14_5_y2;
  assign f_u_arrmul24_fa13_6_f_u_arrmul24_fa12_6_y4 = f_u_arrmul24_fa12_6_y4;
  assign f_u_arrmul24_fa13_6_y0 = f_u_arrmul24_fa13_6_f_u_arrmul24_and13_6_y0 ^ f_u_arrmul24_fa13_6_f_u_arrmul24_fa14_5_y2;
  assign f_u_arrmul24_fa13_6_y1 = f_u_arrmul24_fa13_6_f_u_arrmul24_and13_6_y0 & f_u_arrmul24_fa13_6_f_u_arrmul24_fa14_5_y2;
  assign f_u_arrmul24_fa13_6_y2 = f_u_arrmul24_fa13_6_y0 ^ f_u_arrmul24_fa13_6_f_u_arrmul24_fa12_6_y4;
  assign f_u_arrmul24_fa13_6_y3 = f_u_arrmul24_fa13_6_y0 & f_u_arrmul24_fa13_6_f_u_arrmul24_fa12_6_y4;
  assign f_u_arrmul24_fa13_6_y4 = f_u_arrmul24_fa13_6_y1 | f_u_arrmul24_fa13_6_y3;
  assign f_u_arrmul24_and14_6_a_14 = a_14;
  assign f_u_arrmul24_and14_6_b_6 = b_6;
  assign f_u_arrmul24_and14_6_y0 = f_u_arrmul24_and14_6_a_14 & f_u_arrmul24_and14_6_b_6;
  assign f_u_arrmul24_fa14_6_f_u_arrmul24_and14_6_y0 = f_u_arrmul24_and14_6_y0;
  assign f_u_arrmul24_fa14_6_f_u_arrmul24_fa15_5_y2 = f_u_arrmul24_fa15_5_y2;
  assign f_u_arrmul24_fa14_6_f_u_arrmul24_fa13_6_y4 = f_u_arrmul24_fa13_6_y4;
  assign f_u_arrmul24_fa14_6_y0 = f_u_arrmul24_fa14_6_f_u_arrmul24_and14_6_y0 ^ f_u_arrmul24_fa14_6_f_u_arrmul24_fa15_5_y2;
  assign f_u_arrmul24_fa14_6_y1 = f_u_arrmul24_fa14_6_f_u_arrmul24_and14_6_y0 & f_u_arrmul24_fa14_6_f_u_arrmul24_fa15_5_y2;
  assign f_u_arrmul24_fa14_6_y2 = f_u_arrmul24_fa14_6_y0 ^ f_u_arrmul24_fa14_6_f_u_arrmul24_fa13_6_y4;
  assign f_u_arrmul24_fa14_6_y3 = f_u_arrmul24_fa14_6_y0 & f_u_arrmul24_fa14_6_f_u_arrmul24_fa13_6_y4;
  assign f_u_arrmul24_fa14_6_y4 = f_u_arrmul24_fa14_6_y1 | f_u_arrmul24_fa14_6_y3;
  assign f_u_arrmul24_and15_6_a_15 = a_15;
  assign f_u_arrmul24_and15_6_b_6 = b_6;
  assign f_u_arrmul24_and15_6_y0 = f_u_arrmul24_and15_6_a_15 & f_u_arrmul24_and15_6_b_6;
  assign f_u_arrmul24_fa15_6_f_u_arrmul24_and15_6_y0 = f_u_arrmul24_and15_6_y0;
  assign f_u_arrmul24_fa15_6_f_u_arrmul24_fa16_5_y2 = f_u_arrmul24_fa16_5_y2;
  assign f_u_arrmul24_fa15_6_f_u_arrmul24_fa14_6_y4 = f_u_arrmul24_fa14_6_y4;
  assign f_u_arrmul24_fa15_6_y0 = f_u_arrmul24_fa15_6_f_u_arrmul24_and15_6_y0 ^ f_u_arrmul24_fa15_6_f_u_arrmul24_fa16_5_y2;
  assign f_u_arrmul24_fa15_6_y1 = f_u_arrmul24_fa15_6_f_u_arrmul24_and15_6_y0 & f_u_arrmul24_fa15_6_f_u_arrmul24_fa16_5_y2;
  assign f_u_arrmul24_fa15_6_y2 = f_u_arrmul24_fa15_6_y0 ^ f_u_arrmul24_fa15_6_f_u_arrmul24_fa14_6_y4;
  assign f_u_arrmul24_fa15_6_y3 = f_u_arrmul24_fa15_6_y0 & f_u_arrmul24_fa15_6_f_u_arrmul24_fa14_6_y4;
  assign f_u_arrmul24_fa15_6_y4 = f_u_arrmul24_fa15_6_y1 | f_u_arrmul24_fa15_6_y3;
  assign f_u_arrmul24_and16_6_a_16 = a_16;
  assign f_u_arrmul24_and16_6_b_6 = b_6;
  assign f_u_arrmul24_and16_6_y0 = f_u_arrmul24_and16_6_a_16 & f_u_arrmul24_and16_6_b_6;
  assign f_u_arrmul24_fa16_6_f_u_arrmul24_and16_6_y0 = f_u_arrmul24_and16_6_y0;
  assign f_u_arrmul24_fa16_6_f_u_arrmul24_fa17_5_y2 = f_u_arrmul24_fa17_5_y2;
  assign f_u_arrmul24_fa16_6_f_u_arrmul24_fa15_6_y4 = f_u_arrmul24_fa15_6_y4;
  assign f_u_arrmul24_fa16_6_y0 = f_u_arrmul24_fa16_6_f_u_arrmul24_and16_6_y0 ^ f_u_arrmul24_fa16_6_f_u_arrmul24_fa17_5_y2;
  assign f_u_arrmul24_fa16_6_y1 = f_u_arrmul24_fa16_6_f_u_arrmul24_and16_6_y0 & f_u_arrmul24_fa16_6_f_u_arrmul24_fa17_5_y2;
  assign f_u_arrmul24_fa16_6_y2 = f_u_arrmul24_fa16_6_y0 ^ f_u_arrmul24_fa16_6_f_u_arrmul24_fa15_6_y4;
  assign f_u_arrmul24_fa16_6_y3 = f_u_arrmul24_fa16_6_y0 & f_u_arrmul24_fa16_6_f_u_arrmul24_fa15_6_y4;
  assign f_u_arrmul24_fa16_6_y4 = f_u_arrmul24_fa16_6_y1 | f_u_arrmul24_fa16_6_y3;
  assign f_u_arrmul24_and17_6_a_17 = a_17;
  assign f_u_arrmul24_and17_6_b_6 = b_6;
  assign f_u_arrmul24_and17_6_y0 = f_u_arrmul24_and17_6_a_17 & f_u_arrmul24_and17_6_b_6;
  assign f_u_arrmul24_fa17_6_f_u_arrmul24_and17_6_y0 = f_u_arrmul24_and17_6_y0;
  assign f_u_arrmul24_fa17_6_f_u_arrmul24_fa18_5_y2 = f_u_arrmul24_fa18_5_y2;
  assign f_u_arrmul24_fa17_6_f_u_arrmul24_fa16_6_y4 = f_u_arrmul24_fa16_6_y4;
  assign f_u_arrmul24_fa17_6_y0 = f_u_arrmul24_fa17_6_f_u_arrmul24_and17_6_y0 ^ f_u_arrmul24_fa17_6_f_u_arrmul24_fa18_5_y2;
  assign f_u_arrmul24_fa17_6_y1 = f_u_arrmul24_fa17_6_f_u_arrmul24_and17_6_y0 & f_u_arrmul24_fa17_6_f_u_arrmul24_fa18_5_y2;
  assign f_u_arrmul24_fa17_6_y2 = f_u_arrmul24_fa17_6_y0 ^ f_u_arrmul24_fa17_6_f_u_arrmul24_fa16_6_y4;
  assign f_u_arrmul24_fa17_6_y3 = f_u_arrmul24_fa17_6_y0 & f_u_arrmul24_fa17_6_f_u_arrmul24_fa16_6_y4;
  assign f_u_arrmul24_fa17_6_y4 = f_u_arrmul24_fa17_6_y1 | f_u_arrmul24_fa17_6_y3;
  assign f_u_arrmul24_and18_6_a_18 = a_18;
  assign f_u_arrmul24_and18_6_b_6 = b_6;
  assign f_u_arrmul24_and18_6_y0 = f_u_arrmul24_and18_6_a_18 & f_u_arrmul24_and18_6_b_6;
  assign f_u_arrmul24_fa18_6_f_u_arrmul24_and18_6_y0 = f_u_arrmul24_and18_6_y0;
  assign f_u_arrmul24_fa18_6_f_u_arrmul24_fa19_5_y2 = f_u_arrmul24_fa19_5_y2;
  assign f_u_arrmul24_fa18_6_f_u_arrmul24_fa17_6_y4 = f_u_arrmul24_fa17_6_y4;
  assign f_u_arrmul24_fa18_6_y0 = f_u_arrmul24_fa18_6_f_u_arrmul24_and18_6_y0 ^ f_u_arrmul24_fa18_6_f_u_arrmul24_fa19_5_y2;
  assign f_u_arrmul24_fa18_6_y1 = f_u_arrmul24_fa18_6_f_u_arrmul24_and18_6_y0 & f_u_arrmul24_fa18_6_f_u_arrmul24_fa19_5_y2;
  assign f_u_arrmul24_fa18_6_y2 = f_u_arrmul24_fa18_6_y0 ^ f_u_arrmul24_fa18_6_f_u_arrmul24_fa17_6_y4;
  assign f_u_arrmul24_fa18_6_y3 = f_u_arrmul24_fa18_6_y0 & f_u_arrmul24_fa18_6_f_u_arrmul24_fa17_6_y4;
  assign f_u_arrmul24_fa18_6_y4 = f_u_arrmul24_fa18_6_y1 | f_u_arrmul24_fa18_6_y3;
  assign f_u_arrmul24_and19_6_a_19 = a_19;
  assign f_u_arrmul24_and19_6_b_6 = b_6;
  assign f_u_arrmul24_and19_6_y0 = f_u_arrmul24_and19_6_a_19 & f_u_arrmul24_and19_6_b_6;
  assign f_u_arrmul24_fa19_6_f_u_arrmul24_and19_6_y0 = f_u_arrmul24_and19_6_y0;
  assign f_u_arrmul24_fa19_6_f_u_arrmul24_fa20_5_y2 = f_u_arrmul24_fa20_5_y2;
  assign f_u_arrmul24_fa19_6_f_u_arrmul24_fa18_6_y4 = f_u_arrmul24_fa18_6_y4;
  assign f_u_arrmul24_fa19_6_y0 = f_u_arrmul24_fa19_6_f_u_arrmul24_and19_6_y0 ^ f_u_arrmul24_fa19_6_f_u_arrmul24_fa20_5_y2;
  assign f_u_arrmul24_fa19_6_y1 = f_u_arrmul24_fa19_6_f_u_arrmul24_and19_6_y0 & f_u_arrmul24_fa19_6_f_u_arrmul24_fa20_5_y2;
  assign f_u_arrmul24_fa19_6_y2 = f_u_arrmul24_fa19_6_y0 ^ f_u_arrmul24_fa19_6_f_u_arrmul24_fa18_6_y4;
  assign f_u_arrmul24_fa19_6_y3 = f_u_arrmul24_fa19_6_y0 & f_u_arrmul24_fa19_6_f_u_arrmul24_fa18_6_y4;
  assign f_u_arrmul24_fa19_6_y4 = f_u_arrmul24_fa19_6_y1 | f_u_arrmul24_fa19_6_y3;
  assign f_u_arrmul24_and20_6_a_20 = a_20;
  assign f_u_arrmul24_and20_6_b_6 = b_6;
  assign f_u_arrmul24_and20_6_y0 = f_u_arrmul24_and20_6_a_20 & f_u_arrmul24_and20_6_b_6;
  assign f_u_arrmul24_fa20_6_f_u_arrmul24_and20_6_y0 = f_u_arrmul24_and20_6_y0;
  assign f_u_arrmul24_fa20_6_f_u_arrmul24_fa21_5_y2 = f_u_arrmul24_fa21_5_y2;
  assign f_u_arrmul24_fa20_6_f_u_arrmul24_fa19_6_y4 = f_u_arrmul24_fa19_6_y4;
  assign f_u_arrmul24_fa20_6_y0 = f_u_arrmul24_fa20_6_f_u_arrmul24_and20_6_y0 ^ f_u_arrmul24_fa20_6_f_u_arrmul24_fa21_5_y2;
  assign f_u_arrmul24_fa20_6_y1 = f_u_arrmul24_fa20_6_f_u_arrmul24_and20_6_y0 & f_u_arrmul24_fa20_6_f_u_arrmul24_fa21_5_y2;
  assign f_u_arrmul24_fa20_6_y2 = f_u_arrmul24_fa20_6_y0 ^ f_u_arrmul24_fa20_6_f_u_arrmul24_fa19_6_y4;
  assign f_u_arrmul24_fa20_6_y3 = f_u_arrmul24_fa20_6_y0 & f_u_arrmul24_fa20_6_f_u_arrmul24_fa19_6_y4;
  assign f_u_arrmul24_fa20_6_y4 = f_u_arrmul24_fa20_6_y1 | f_u_arrmul24_fa20_6_y3;
  assign f_u_arrmul24_and21_6_a_21 = a_21;
  assign f_u_arrmul24_and21_6_b_6 = b_6;
  assign f_u_arrmul24_and21_6_y0 = f_u_arrmul24_and21_6_a_21 & f_u_arrmul24_and21_6_b_6;
  assign f_u_arrmul24_fa21_6_f_u_arrmul24_and21_6_y0 = f_u_arrmul24_and21_6_y0;
  assign f_u_arrmul24_fa21_6_f_u_arrmul24_fa22_5_y2 = f_u_arrmul24_fa22_5_y2;
  assign f_u_arrmul24_fa21_6_f_u_arrmul24_fa20_6_y4 = f_u_arrmul24_fa20_6_y4;
  assign f_u_arrmul24_fa21_6_y0 = f_u_arrmul24_fa21_6_f_u_arrmul24_and21_6_y0 ^ f_u_arrmul24_fa21_6_f_u_arrmul24_fa22_5_y2;
  assign f_u_arrmul24_fa21_6_y1 = f_u_arrmul24_fa21_6_f_u_arrmul24_and21_6_y0 & f_u_arrmul24_fa21_6_f_u_arrmul24_fa22_5_y2;
  assign f_u_arrmul24_fa21_6_y2 = f_u_arrmul24_fa21_6_y0 ^ f_u_arrmul24_fa21_6_f_u_arrmul24_fa20_6_y4;
  assign f_u_arrmul24_fa21_6_y3 = f_u_arrmul24_fa21_6_y0 & f_u_arrmul24_fa21_6_f_u_arrmul24_fa20_6_y4;
  assign f_u_arrmul24_fa21_6_y4 = f_u_arrmul24_fa21_6_y1 | f_u_arrmul24_fa21_6_y3;
  assign f_u_arrmul24_and22_6_a_22 = a_22;
  assign f_u_arrmul24_and22_6_b_6 = b_6;
  assign f_u_arrmul24_and22_6_y0 = f_u_arrmul24_and22_6_a_22 & f_u_arrmul24_and22_6_b_6;
  assign f_u_arrmul24_fa22_6_f_u_arrmul24_and22_6_y0 = f_u_arrmul24_and22_6_y0;
  assign f_u_arrmul24_fa22_6_f_u_arrmul24_fa23_5_y2 = f_u_arrmul24_fa23_5_y2;
  assign f_u_arrmul24_fa22_6_f_u_arrmul24_fa21_6_y4 = f_u_arrmul24_fa21_6_y4;
  assign f_u_arrmul24_fa22_6_y0 = f_u_arrmul24_fa22_6_f_u_arrmul24_and22_6_y0 ^ f_u_arrmul24_fa22_6_f_u_arrmul24_fa23_5_y2;
  assign f_u_arrmul24_fa22_6_y1 = f_u_arrmul24_fa22_6_f_u_arrmul24_and22_6_y0 & f_u_arrmul24_fa22_6_f_u_arrmul24_fa23_5_y2;
  assign f_u_arrmul24_fa22_6_y2 = f_u_arrmul24_fa22_6_y0 ^ f_u_arrmul24_fa22_6_f_u_arrmul24_fa21_6_y4;
  assign f_u_arrmul24_fa22_6_y3 = f_u_arrmul24_fa22_6_y0 & f_u_arrmul24_fa22_6_f_u_arrmul24_fa21_6_y4;
  assign f_u_arrmul24_fa22_6_y4 = f_u_arrmul24_fa22_6_y1 | f_u_arrmul24_fa22_6_y3;
  assign f_u_arrmul24_and23_6_a_23 = a_23;
  assign f_u_arrmul24_and23_6_b_6 = b_6;
  assign f_u_arrmul24_and23_6_y0 = f_u_arrmul24_and23_6_a_23 & f_u_arrmul24_and23_6_b_6;
  assign f_u_arrmul24_fa23_6_f_u_arrmul24_and23_6_y0 = f_u_arrmul24_and23_6_y0;
  assign f_u_arrmul24_fa23_6_f_u_arrmul24_fa23_5_y4 = f_u_arrmul24_fa23_5_y4;
  assign f_u_arrmul24_fa23_6_f_u_arrmul24_fa22_6_y4 = f_u_arrmul24_fa22_6_y4;
  assign f_u_arrmul24_fa23_6_y0 = f_u_arrmul24_fa23_6_f_u_arrmul24_and23_6_y0 ^ f_u_arrmul24_fa23_6_f_u_arrmul24_fa23_5_y4;
  assign f_u_arrmul24_fa23_6_y1 = f_u_arrmul24_fa23_6_f_u_arrmul24_and23_6_y0 & f_u_arrmul24_fa23_6_f_u_arrmul24_fa23_5_y4;
  assign f_u_arrmul24_fa23_6_y2 = f_u_arrmul24_fa23_6_y0 ^ f_u_arrmul24_fa23_6_f_u_arrmul24_fa22_6_y4;
  assign f_u_arrmul24_fa23_6_y3 = f_u_arrmul24_fa23_6_y0 & f_u_arrmul24_fa23_6_f_u_arrmul24_fa22_6_y4;
  assign f_u_arrmul24_fa23_6_y4 = f_u_arrmul24_fa23_6_y1 | f_u_arrmul24_fa23_6_y3;
  assign f_u_arrmul24_and0_7_a_0 = a_0;
  assign f_u_arrmul24_and0_7_b_7 = b_7;
  assign f_u_arrmul24_and0_7_y0 = f_u_arrmul24_and0_7_a_0 & f_u_arrmul24_and0_7_b_7;
  assign f_u_arrmul24_ha0_7_f_u_arrmul24_and0_7_y0 = f_u_arrmul24_and0_7_y0;
  assign f_u_arrmul24_ha0_7_f_u_arrmul24_fa1_6_y2 = f_u_arrmul24_fa1_6_y2;
  assign f_u_arrmul24_ha0_7_y0 = f_u_arrmul24_ha0_7_f_u_arrmul24_and0_7_y0 ^ f_u_arrmul24_ha0_7_f_u_arrmul24_fa1_6_y2;
  assign f_u_arrmul24_ha0_7_y1 = f_u_arrmul24_ha0_7_f_u_arrmul24_and0_7_y0 & f_u_arrmul24_ha0_7_f_u_arrmul24_fa1_6_y2;
  assign f_u_arrmul24_and1_7_a_1 = a_1;
  assign f_u_arrmul24_and1_7_b_7 = b_7;
  assign f_u_arrmul24_and1_7_y0 = f_u_arrmul24_and1_7_a_1 & f_u_arrmul24_and1_7_b_7;
  assign f_u_arrmul24_fa1_7_f_u_arrmul24_and1_7_y0 = f_u_arrmul24_and1_7_y0;
  assign f_u_arrmul24_fa1_7_f_u_arrmul24_fa2_6_y2 = f_u_arrmul24_fa2_6_y2;
  assign f_u_arrmul24_fa1_7_f_u_arrmul24_ha0_7_y1 = f_u_arrmul24_ha0_7_y1;
  assign f_u_arrmul24_fa1_7_y0 = f_u_arrmul24_fa1_7_f_u_arrmul24_and1_7_y0 ^ f_u_arrmul24_fa1_7_f_u_arrmul24_fa2_6_y2;
  assign f_u_arrmul24_fa1_7_y1 = f_u_arrmul24_fa1_7_f_u_arrmul24_and1_7_y0 & f_u_arrmul24_fa1_7_f_u_arrmul24_fa2_6_y2;
  assign f_u_arrmul24_fa1_7_y2 = f_u_arrmul24_fa1_7_y0 ^ f_u_arrmul24_fa1_7_f_u_arrmul24_ha0_7_y1;
  assign f_u_arrmul24_fa1_7_y3 = f_u_arrmul24_fa1_7_y0 & f_u_arrmul24_fa1_7_f_u_arrmul24_ha0_7_y1;
  assign f_u_arrmul24_fa1_7_y4 = f_u_arrmul24_fa1_7_y1 | f_u_arrmul24_fa1_7_y3;
  assign f_u_arrmul24_and2_7_a_2 = a_2;
  assign f_u_arrmul24_and2_7_b_7 = b_7;
  assign f_u_arrmul24_and2_7_y0 = f_u_arrmul24_and2_7_a_2 & f_u_arrmul24_and2_7_b_7;
  assign f_u_arrmul24_fa2_7_f_u_arrmul24_and2_7_y0 = f_u_arrmul24_and2_7_y0;
  assign f_u_arrmul24_fa2_7_f_u_arrmul24_fa3_6_y2 = f_u_arrmul24_fa3_6_y2;
  assign f_u_arrmul24_fa2_7_f_u_arrmul24_fa1_7_y4 = f_u_arrmul24_fa1_7_y4;
  assign f_u_arrmul24_fa2_7_y0 = f_u_arrmul24_fa2_7_f_u_arrmul24_and2_7_y0 ^ f_u_arrmul24_fa2_7_f_u_arrmul24_fa3_6_y2;
  assign f_u_arrmul24_fa2_7_y1 = f_u_arrmul24_fa2_7_f_u_arrmul24_and2_7_y0 & f_u_arrmul24_fa2_7_f_u_arrmul24_fa3_6_y2;
  assign f_u_arrmul24_fa2_7_y2 = f_u_arrmul24_fa2_7_y0 ^ f_u_arrmul24_fa2_7_f_u_arrmul24_fa1_7_y4;
  assign f_u_arrmul24_fa2_7_y3 = f_u_arrmul24_fa2_7_y0 & f_u_arrmul24_fa2_7_f_u_arrmul24_fa1_7_y4;
  assign f_u_arrmul24_fa2_7_y4 = f_u_arrmul24_fa2_7_y1 | f_u_arrmul24_fa2_7_y3;
  assign f_u_arrmul24_and3_7_a_3 = a_3;
  assign f_u_arrmul24_and3_7_b_7 = b_7;
  assign f_u_arrmul24_and3_7_y0 = f_u_arrmul24_and3_7_a_3 & f_u_arrmul24_and3_7_b_7;
  assign f_u_arrmul24_fa3_7_f_u_arrmul24_and3_7_y0 = f_u_arrmul24_and3_7_y0;
  assign f_u_arrmul24_fa3_7_f_u_arrmul24_fa4_6_y2 = f_u_arrmul24_fa4_6_y2;
  assign f_u_arrmul24_fa3_7_f_u_arrmul24_fa2_7_y4 = f_u_arrmul24_fa2_7_y4;
  assign f_u_arrmul24_fa3_7_y0 = f_u_arrmul24_fa3_7_f_u_arrmul24_and3_7_y0 ^ f_u_arrmul24_fa3_7_f_u_arrmul24_fa4_6_y2;
  assign f_u_arrmul24_fa3_7_y1 = f_u_arrmul24_fa3_7_f_u_arrmul24_and3_7_y0 & f_u_arrmul24_fa3_7_f_u_arrmul24_fa4_6_y2;
  assign f_u_arrmul24_fa3_7_y2 = f_u_arrmul24_fa3_7_y0 ^ f_u_arrmul24_fa3_7_f_u_arrmul24_fa2_7_y4;
  assign f_u_arrmul24_fa3_7_y3 = f_u_arrmul24_fa3_7_y0 & f_u_arrmul24_fa3_7_f_u_arrmul24_fa2_7_y4;
  assign f_u_arrmul24_fa3_7_y4 = f_u_arrmul24_fa3_7_y1 | f_u_arrmul24_fa3_7_y3;
  assign f_u_arrmul24_and4_7_a_4 = a_4;
  assign f_u_arrmul24_and4_7_b_7 = b_7;
  assign f_u_arrmul24_and4_7_y0 = f_u_arrmul24_and4_7_a_4 & f_u_arrmul24_and4_7_b_7;
  assign f_u_arrmul24_fa4_7_f_u_arrmul24_and4_7_y0 = f_u_arrmul24_and4_7_y0;
  assign f_u_arrmul24_fa4_7_f_u_arrmul24_fa5_6_y2 = f_u_arrmul24_fa5_6_y2;
  assign f_u_arrmul24_fa4_7_f_u_arrmul24_fa3_7_y4 = f_u_arrmul24_fa3_7_y4;
  assign f_u_arrmul24_fa4_7_y0 = f_u_arrmul24_fa4_7_f_u_arrmul24_and4_7_y0 ^ f_u_arrmul24_fa4_7_f_u_arrmul24_fa5_6_y2;
  assign f_u_arrmul24_fa4_7_y1 = f_u_arrmul24_fa4_7_f_u_arrmul24_and4_7_y0 & f_u_arrmul24_fa4_7_f_u_arrmul24_fa5_6_y2;
  assign f_u_arrmul24_fa4_7_y2 = f_u_arrmul24_fa4_7_y0 ^ f_u_arrmul24_fa4_7_f_u_arrmul24_fa3_7_y4;
  assign f_u_arrmul24_fa4_7_y3 = f_u_arrmul24_fa4_7_y0 & f_u_arrmul24_fa4_7_f_u_arrmul24_fa3_7_y4;
  assign f_u_arrmul24_fa4_7_y4 = f_u_arrmul24_fa4_7_y1 | f_u_arrmul24_fa4_7_y3;
  assign f_u_arrmul24_and5_7_a_5 = a_5;
  assign f_u_arrmul24_and5_7_b_7 = b_7;
  assign f_u_arrmul24_and5_7_y0 = f_u_arrmul24_and5_7_a_5 & f_u_arrmul24_and5_7_b_7;
  assign f_u_arrmul24_fa5_7_f_u_arrmul24_and5_7_y0 = f_u_arrmul24_and5_7_y0;
  assign f_u_arrmul24_fa5_7_f_u_arrmul24_fa6_6_y2 = f_u_arrmul24_fa6_6_y2;
  assign f_u_arrmul24_fa5_7_f_u_arrmul24_fa4_7_y4 = f_u_arrmul24_fa4_7_y4;
  assign f_u_arrmul24_fa5_7_y0 = f_u_arrmul24_fa5_7_f_u_arrmul24_and5_7_y0 ^ f_u_arrmul24_fa5_7_f_u_arrmul24_fa6_6_y2;
  assign f_u_arrmul24_fa5_7_y1 = f_u_arrmul24_fa5_7_f_u_arrmul24_and5_7_y0 & f_u_arrmul24_fa5_7_f_u_arrmul24_fa6_6_y2;
  assign f_u_arrmul24_fa5_7_y2 = f_u_arrmul24_fa5_7_y0 ^ f_u_arrmul24_fa5_7_f_u_arrmul24_fa4_7_y4;
  assign f_u_arrmul24_fa5_7_y3 = f_u_arrmul24_fa5_7_y0 & f_u_arrmul24_fa5_7_f_u_arrmul24_fa4_7_y4;
  assign f_u_arrmul24_fa5_7_y4 = f_u_arrmul24_fa5_7_y1 | f_u_arrmul24_fa5_7_y3;
  assign f_u_arrmul24_and6_7_a_6 = a_6;
  assign f_u_arrmul24_and6_7_b_7 = b_7;
  assign f_u_arrmul24_and6_7_y0 = f_u_arrmul24_and6_7_a_6 & f_u_arrmul24_and6_7_b_7;
  assign f_u_arrmul24_fa6_7_f_u_arrmul24_and6_7_y0 = f_u_arrmul24_and6_7_y0;
  assign f_u_arrmul24_fa6_7_f_u_arrmul24_fa7_6_y2 = f_u_arrmul24_fa7_6_y2;
  assign f_u_arrmul24_fa6_7_f_u_arrmul24_fa5_7_y4 = f_u_arrmul24_fa5_7_y4;
  assign f_u_arrmul24_fa6_7_y0 = f_u_arrmul24_fa6_7_f_u_arrmul24_and6_7_y0 ^ f_u_arrmul24_fa6_7_f_u_arrmul24_fa7_6_y2;
  assign f_u_arrmul24_fa6_7_y1 = f_u_arrmul24_fa6_7_f_u_arrmul24_and6_7_y0 & f_u_arrmul24_fa6_7_f_u_arrmul24_fa7_6_y2;
  assign f_u_arrmul24_fa6_7_y2 = f_u_arrmul24_fa6_7_y0 ^ f_u_arrmul24_fa6_7_f_u_arrmul24_fa5_7_y4;
  assign f_u_arrmul24_fa6_7_y3 = f_u_arrmul24_fa6_7_y0 & f_u_arrmul24_fa6_7_f_u_arrmul24_fa5_7_y4;
  assign f_u_arrmul24_fa6_7_y4 = f_u_arrmul24_fa6_7_y1 | f_u_arrmul24_fa6_7_y3;
  assign f_u_arrmul24_and7_7_a_7 = a_7;
  assign f_u_arrmul24_and7_7_b_7 = b_7;
  assign f_u_arrmul24_and7_7_y0 = f_u_arrmul24_and7_7_a_7 & f_u_arrmul24_and7_7_b_7;
  assign f_u_arrmul24_fa7_7_f_u_arrmul24_and7_7_y0 = f_u_arrmul24_and7_7_y0;
  assign f_u_arrmul24_fa7_7_f_u_arrmul24_fa8_6_y2 = f_u_arrmul24_fa8_6_y2;
  assign f_u_arrmul24_fa7_7_f_u_arrmul24_fa6_7_y4 = f_u_arrmul24_fa6_7_y4;
  assign f_u_arrmul24_fa7_7_y0 = f_u_arrmul24_fa7_7_f_u_arrmul24_and7_7_y0 ^ f_u_arrmul24_fa7_7_f_u_arrmul24_fa8_6_y2;
  assign f_u_arrmul24_fa7_7_y1 = f_u_arrmul24_fa7_7_f_u_arrmul24_and7_7_y0 & f_u_arrmul24_fa7_7_f_u_arrmul24_fa8_6_y2;
  assign f_u_arrmul24_fa7_7_y2 = f_u_arrmul24_fa7_7_y0 ^ f_u_arrmul24_fa7_7_f_u_arrmul24_fa6_7_y4;
  assign f_u_arrmul24_fa7_7_y3 = f_u_arrmul24_fa7_7_y0 & f_u_arrmul24_fa7_7_f_u_arrmul24_fa6_7_y4;
  assign f_u_arrmul24_fa7_7_y4 = f_u_arrmul24_fa7_7_y1 | f_u_arrmul24_fa7_7_y3;
  assign f_u_arrmul24_and8_7_a_8 = a_8;
  assign f_u_arrmul24_and8_7_b_7 = b_7;
  assign f_u_arrmul24_and8_7_y0 = f_u_arrmul24_and8_7_a_8 & f_u_arrmul24_and8_7_b_7;
  assign f_u_arrmul24_fa8_7_f_u_arrmul24_and8_7_y0 = f_u_arrmul24_and8_7_y0;
  assign f_u_arrmul24_fa8_7_f_u_arrmul24_fa9_6_y2 = f_u_arrmul24_fa9_6_y2;
  assign f_u_arrmul24_fa8_7_f_u_arrmul24_fa7_7_y4 = f_u_arrmul24_fa7_7_y4;
  assign f_u_arrmul24_fa8_7_y0 = f_u_arrmul24_fa8_7_f_u_arrmul24_and8_7_y0 ^ f_u_arrmul24_fa8_7_f_u_arrmul24_fa9_6_y2;
  assign f_u_arrmul24_fa8_7_y1 = f_u_arrmul24_fa8_7_f_u_arrmul24_and8_7_y0 & f_u_arrmul24_fa8_7_f_u_arrmul24_fa9_6_y2;
  assign f_u_arrmul24_fa8_7_y2 = f_u_arrmul24_fa8_7_y0 ^ f_u_arrmul24_fa8_7_f_u_arrmul24_fa7_7_y4;
  assign f_u_arrmul24_fa8_7_y3 = f_u_arrmul24_fa8_7_y0 & f_u_arrmul24_fa8_7_f_u_arrmul24_fa7_7_y4;
  assign f_u_arrmul24_fa8_7_y4 = f_u_arrmul24_fa8_7_y1 | f_u_arrmul24_fa8_7_y3;
  assign f_u_arrmul24_and9_7_a_9 = a_9;
  assign f_u_arrmul24_and9_7_b_7 = b_7;
  assign f_u_arrmul24_and9_7_y0 = f_u_arrmul24_and9_7_a_9 & f_u_arrmul24_and9_7_b_7;
  assign f_u_arrmul24_fa9_7_f_u_arrmul24_and9_7_y0 = f_u_arrmul24_and9_7_y0;
  assign f_u_arrmul24_fa9_7_f_u_arrmul24_fa10_6_y2 = f_u_arrmul24_fa10_6_y2;
  assign f_u_arrmul24_fa9_7_f_u_arrmul24_fa8_7_y4 = f_u_arrmul24_fa8_7_y4;
  assign f_u_arrmul24_fa9_7_y0 = f_u_arrmul24_fa9_7_f_u_arrmul24_and9_7_y0 ^ f_u_arrmul24_fa9_7_f_u_arrmul24_fa10_6_y2;
  assign f_u_arrmul24_fa9_7_y1 = f_u_arrmul24_fa9_7_f_u_arrmul24_and9_7_y0 & f_u_arrmul24_fa9_7_f_u_arrmul24_fa10_6_y2;
  assign f_u_arrmul24_fa9_7_y2 = f_u_arrmul24_fa9_7_y0 ^ f_u_arrmul24_fa9_7_f_u_arrmul24_fa8_7_y4;
  assign f_u_arrmul24_fa9_7_y3 = f_u_arrmul24_fa9_7_y0 & f_u_arrmul24_fa9_7_f_u_arrmul24_fa8_7_y4;
  assign f_u_arrmul24_fa9_7_y4 = f_u_arrmul24_fa9_7_y1 | f_u_arrmul24_fa9_7_y3;
  assign f_u_arrmul24_and10_7_a_10 = a_10;
  assign f_u_arrmul24_and10_7_b_7 = b_7;
  assign f_u_arrmul24_and10_7_y0 = f_u_arrmul24_and10_7_a_10 & f_u_arrmul24_and10_7_b_7;
  assign f_u_arrmul24_fa10_7_f_u_arrmul24_and10_7_y0 = f_u_arrmul24_and10_7_y0;
  assign f_u_arrmul24_fa10_7_f_u_arrmul24_fa11_6_y2 = f_u_arrmul24_fa11_6_y2;
  assign f_u_arrmul24_fa10_7_f_u_arrmul24_fa9_7_y4 = f_u_arrmul24_fa9_7_y4;
  assign f_u_arrmul24_fa10_7_y0 = f_u_arrmul24_fa10_7_f_u_arrmul24_and10_7_y0 ^ f_u_arrmul24_fa10_7_f_u_arrmul24_fa11_6_y2;
  assign f_u_arrmul24_fa10_7_y1 = f_u_arrmul24_fa10_7_f_u_arrmul24_and10_7_y0 & f_u_arrmul24_fa10_7_f_u_arrmul24_fa11_6_y2;
  assign f_u_arrmul24_fa10_7_y2 = f_u_arrmul24_fa10_7_y0 ^ f_u_arrmul24_fa10_7_f_u_arrmul24_fa9_7_y4;
  assign f_u_arrmul24_fa10_7_y3 = f_u_arrmul24_fa10_7_y0 & f_u_arrmul24_fa10_7_f_u_arrmul24_fa9_7_y4;
  assign f_u_arrmul24_fa10_7_y4 = f_u_arrmul24_fa10_7_y1 | f_u_arrmul24_fa10_7_y3;
  assign f_u_arrmul24_and11_7_a_11 = a_11;
  assign f_u_arrmul24_and11_7_b_7 = b_7;
  assign f_u_arrmul24_and11_7_y0 = f_u_arrmul24_and11_7_a_11 & f_u_arrmul24_and11_7_b_7;
  assign f_u_arrmul24_fa11_7_f_u_arrmul24_and11_7_y0 = f_u_arrmul24_and11_7_y0;
  assign f_u_arrmul24_fa11_7_f_u_arrmul24_fa12_6_y2 = f_u_arrmul24_fa12_6_y2;
  assign f_u_arrmul24_fa11_7_f_u_arrmul24_fa10_7_y4 = f_u_arrmul24_fa10_7_y4;
  assign f_u_arrmul24_fa11_7_y0 = f_u_arrmul24_fa11_7_f_u_arrmul24_and11_7_y0 ^ f_u_arrmul24_fa11_7_f_u_arrmul24_fa12_6_y2;
  assign f_u_arrmul24_fa11_7_y1 = f_u_arrmul24_fa11_7_f_u_arrmul24_and11_7_y0 & f_u_arrmul24_fa11_7_f_u_arrmul24_fa12_6_y2;
  assign f_u_arrmul24_fa11_7_y2 = f_u_arrmul24_fa11_7_y0 ^ f_u_arrmul24_fa11_7_f_u_arrmul24_fa10_7_y4;
  assign f_u_arrmul24_fa11_7_y3 = f_u_arrmul24_fa11_7_y0 & f_u_arrmul24_fa11_7_f_u_arrmul24_fa10_7_y4;
  assign f_u_arrmul24_fa11_7_y4 = f_u_arrmul24_fa11_7_y1 | f_u_arrmul24_fa11_7_y3;
  assign f_u_arrmul24_and12_7_a_12 = a_12;
  assign f_u_arrmul24_and12_7_b_7 = b_7;
  assign f_u_arrmul24_and12_7_y0 = f_u_arrmul24_and12_7_a_12 & f_u_arrmul24_and12_7_b_7;
  assign f_u_arrmul24_fa12_7_f_u_arrmul24_and12_7_y0 = f_u_arrmul24_and12_7_y0;
  assign f_u_arrmul24_fa12_7_f_u_arrmul24_fa13_6_y2 = f_u_arrmul24_fa13_6_y2;
  assign f_u_arrmul24_fa12_7_f_u_arrmul24_fa11_7_y4 = f_u_arrmul24_fa11_7_y4;
  assign f_u_arrmul24_fa12_7_y0 = f_u_arrmul24_fa12_7_f_u_arrmul24_and12_7_y0 ^ f_u_arrmul24_fa12_7_f_u_arrmul24_fa13_6_y2;
  assign f_u_arrmul24_fa12_7_y1 = f_u_arrmul24_fa12_7_f_u_arrmul24_and12_7_y0 & f_u_arrmul24_fa12_7_f_u_arrmul24_fa13_6_y2;
  assign f_u_arrmul24_fa12_7_y2 = f_u_arrmul24_fa12_7_y0 ^ f_u_arrmul24_fa12_7_f_u_arrmul24_fa11_7_y4;
  assign f_u_arrmul24_fa12_7_y3 = f_u_arrmul24_fa12_7_y0 & f_u_arrmul24_fa12_7_f_u_arrmul24_fa11_7_y4;
  assign f_u_arrmul24_fa12_7_y4 = f_u_arrmul24_fa12_7_y1 | f_u_arrmul24_fa12_7_y3;
  assign f_u_arrmul24_and13_7_a_13 = a_13;
  assign f_u_arrmul24_and13_7_b_7 = b_7;
  assign f_u_arrmul24_and13_7_y0 = f_u_arrmul24_and13_7_a_13 & f_u_arrmul24_and13_7_b_7;
  assign f_u_arrmul24_fa13_7_f_u_arrmul24_and13_7_y0 = f_u_arrmul24_and13_7_y0;
  assign f_u_arrmul24_fa13_7_f_u_arrmul24_fa14_6_y2 = f_u_arrmul24_fa14_6_y2;
  assign f_u_arrmul24_fa13_7_f_u_arrmul24_fa12_7_y4 = f_u_arrmul24_fa12_7_y4;
  assign f_u_arrmul24_fa13_7_y0 = f_u_arrmul24_fa13_7_f_u_arrmul24_and13_7_y0 ^ f_u_arrmul24_fa13_7_f_u_arrmul24_fa14_6_y2;
  assign f_u_arrmul24_fa13_7_y1 = f_u_arrmul24_fa13_7_f_u_arrmul24_and13_7_y0 & f_u_arrmul24_fa13_7_f_u_arrmul24_fa14_6_y2;
  assign f_u_arrmul24_fa13_7_y2 = f_u_arrmul24_fa13_7_y0 ^ f_u_arrmul24_fa13_7_f_u_arrmul24_fa12_7_y4;
  assign f_u_arrmul24_fa13_7_y3 = f_u_arrmul24_fa13_7_y0 & f_u_arrmul24_fa13_7_f_u_arrmul24_fa12_7_y4;
  assign f_u_arrmul24_fa13_7_y4 = f_u_arrmul24_fa13_7_y1 | f_u_arrmul24_fa13_7_y3;
  assign f_u_arrmul24_and14_7_a_14 = a_14;
  assign f_u_arrmul24_and14_7_b_7 = b_7;
  assign f_u_arrmul24_and14_7_y0 = f_u_arrmul24_and14_7_a_14 & f_u_arrmul24_and14_7_b_7;
  assign f_u_arrmul24_fa14_7_f_u_arrmul24_and14_7_y0 = f_u_arrmul24_and14_7_y0;
  assign f_u_arrmul24_fa14_7_f_u_arrmul24_fa15_6_y2 = f_u_arrmul24_fa15_6_y2;
  assign f_u_arrmul24_fa14_7_f_u_arrmul24_fa13_7_y4 = f_u_arrmul24_fa13_7_y4;
  assign f_u_arrmul24_fa14_7_y0 = f_u_arrmul24_fa14_7_f_u_arrmul24_and14_7_y0 ^ f_u_arrmul24_fa14_7_f_u_arrmul24_fa15_6_y2;
  assign f_u_arrmul24_fa14_7_y1 = f_u_arrmul24_fa14_7_f_u_arrmul24_and14_7_y0 & f_u_arrmul24_fa14_7_f_u_arrmul24_fa15_6_y2;
  assign f_u_arrmul24_fa14_7_y2 = f_u_arrmul24_fa14_7_y0 ^ f_u_arrmul24_fa14_7_f_u_arrmul24_fa13_7_y4;
  assign f_u_arrmul24_fa14_7_y3 = f_u_arrmul24_fa14_7_y0 & f_u_arrmul24_fa14_7_f_u_arrmul24_fa13_7_y4;
  assign f_u_arrmul24_fa14_7_y4 = f_u_arrmul24_fa14_7_y1 | f_u_arrmul24_fa14_7_y3;
  assign f_u_arrmul24_and15_7_a_15 = a_15;
  assign f_u_arrmul24_and15_7_b_7 = b_7;
  assign f_u_arrmul24_and15_7_y0 = f_u_arrmul24_and15_7_a_15 & f_u_arrmul24_and15_7_b_7;
  assign f_u_arrmul24_fa15_7_f_u_arrmul24_and15_7_y0 = f_u_arrmul24_and15_7_y0;
  assign f_u_arrmul24_fa15_7_f_u_arrmul24_fa16_6_y2 = f_u_arrmul24_fa16_6_y2;
  assign f_u_arrmul24_fa15_7_f_u_arrmul24_fa14_7_y4 = f_u_arrmul24_fa14_7_y4;
  assign f_u_arrmul24_fa15_7_y0 = f_u_arrmul24_fa15_7_f_u_arrmul24_and15_7_y0 ^ f_u_arrmul24_fa15_7_f_u_arrmul24_fa16_6_y2;
  assign f_u_arrmul24_fa15_7_y1 = f_u_arrmul24_fa15_7_f_u_arrmul24_and15_7_y0 & f_u_arrmul24_fa15_7_f_u_arrmul24_fa16_6_y2;
  assign f_u_arrmul24_fa15_7_y2 = f_u_arrmul24_fa15_7_y0 ^ f_u_arrmul24_fa15_7_f_u_arrmul24_fa14_7_y4;
  assign f_u_arrmul24_fa15_7_y3 = f_u_arrmul24_fa15_7_y0 & f_u_arrmul24_fa15_7_f_u_arrmul24_fa14_7_y4;
  assign f_u_arrmul24_fa15_7_y4 = f_u_arrmul24_fa15_7_y1 | f_u_arrmul24_fa15_7_y3;
  assign f_u_arrmul24_and16_7_a_16 = a_16;
  assign f_u_arrmul24_and16_7_b_7 = b_7;
  assign f_u_arrmul24_and16_7_y0 = f_u_arrmul24_and16_7_a_16 & f_u_arrmul24_and16_7_b_7;
  assign f_u_arrmul24_fa16_7_f_u_arrmul24_and16_7_y0 = f_u_arrmul24_and16_7_y0;
  assign f_u_arrmul24_fa16_7_f_u_arrmul24_fa17_6_y2 = f_u_arrmul24_fa17_6_y2;
  assign f_u_arrmul24_fa16_7_f_u_arrmul24_fa15_7_y4 = f_u_arrmul24_fa15_7_y4;
  assign f_u_arrmul24_fa16_7_y0 = f_u_arrmul24_fa16_7_f_u_arrmul24_and16_7_y0 ^ f_u_arrmul24_fa16_7_f_u_arrmul24_fa17_6_y2;
  assign f_u_arrmul24_fa16_7_y1 = f_u_arrmul24_fa16_7_f_u_arrmul24_and16_7_y0 & f_u_arrmul24_fa16_7_f_u_arrmul24_fa17_6_y2;
  assign f_u_arrmul24_fa16_7_y2 = f_u_arrmul24_fa16_7_y0 ^ f_u_arrmul24_fa16_7_f_u_arrmul24_fa15_7_y4;
  assign f_u_arrmul24_fa16_7_y3 = f_u_arrmul24_fa16_7_y0 & f_u_arrmul24_fa16_7_f_u_arrmul24_fa15_7_y4;
  assign f_u_arrmul24_fa16_7_y4 = f_u_arrmul24_fa16_7_y1 | f_u_arrmul24_fa16_7_y3;
  assign f_u_arrmul24_and17_7_a_17 = a_17;
  assign f_u_arrmul24_and17_7_b_7 = b_7;
  assign f_u_arrmul24_and17_7_y0 = f_u_arrmul24_and17_7_a_17 & f_u_arrmul24_and17_7_b_7;
  assign f_u_arrmul24_fa17_7_f_u_arrmul24_and17_7_y0 = f_u_arrmul24_and17_7_y0;
  assign f_u_arrmul24_fa17_7_f_u_arrmul24_fa18_6_y2 = f_u_arrmul24_fa18_6_y2;
  assign f_u_arrmul24_fa17_7_f_u_arrmul24_fa16_7_y4 = f_u_arrmul24_fa16_7_y4;
  assign f_u_arrmul24_fa17_7_y0 = f_u_arrmul24_fa17_7_f_u_arrmul24_and17_7_y0 ^ f_u_arrmul24_fa17_7_f_u_arrmul24_fa18_6_y2;
  assign f_u_arrmul24_fa17_7_y1 = f_u_arrmul24_fa17_7_f_u_arrmul24_and17_7_y0 & f_u_arrmul24_fa17_7_f_u_arrmul24_fa18_6_y2;
  assign f_u_arrmul24_fa17_7_y2 = f_u_arrmul24_fa17_7_y0 ^ f_u_arrmul24_fa17_7_f_u_arrmul24_fa16_7_y4;
  assign f_u_arrmul24_fa17_7_y3 = f_u_arrmul24_fa17_7_y0 & f_u_arrmul24_fa17_7_f_u_arrmul24_fa16_7_y4;
  assign f_u_arrmul24_fa17_7_y4 = f_u_arrmul24_fa17_7_y1 | f_u_arrmul24_fa17_7_y3;
  assign f_u_arrmul24_and18_7_a_18 = a_18;
  assign f_u_arrmul24_and18_7_b_7 = b_7;
  assign f_u_arrmul24_and18_7_y0 = f_u_arrmul24_and18_7_a_18 & f_u_arrmul24_and18_7_b_7;
  assign f_u_arrmul24_fa18_7_f_u_arrmul24_and18_7_y0 = f_u_arrmul24_and18_7_y0;
  assign f_u_arrmul24_fa18_7_f_u_arrmul24_fa19_6_y2 = f_u_arrmul24_fa19_6_y2;
  assign f_u_arrmul24_fa18_7_f_u_arrmul24_fa17_7_y4 = f_u_arrmul24_fa17_7_y4;
  assign f_u_arrmul24_fa18_7_y0 = f_u_arrmul24_fa18_7_f_u_arrmul24_and18_7_y0 ^ f_u_arrmul24_fa18_7_f_u_arrmul24_fa19_6_y2;
  assign f_u_arrmul24_fa18_7_y1 = f_u_arrmul24_fa18_7_f_u_arrmul24_and18_7_y0 & f_u_arrmul24_fa18_7_f_u_arrmul24_fa19_6_y2;
  assign f_u_arrmul24_fa18_7_y2 = f_u_arrmul24_fa18_7_y0 ^ f_u_arrmul24_fa18_7_f_u_arrmul24_fa17_7_y4;
  assign f_u_arrmul24_fa18_7_y3 = f_u_arrmul24_fa18_7_y0 & f_u_arrmul24_fa18_7_f_u_arrmul24_fa17_7_y4;
  assign f_u_arrmul24_fa18_7_y4 = f_u_arrmul24_fa18_7_y1 | f_u_arrmul24_fa18_7_y3;
  assign f_u_arrmul24_and19_7_a_19 = a_19;
  assign f_u_arrmul24_and19_7_b_7 = b_7;
  assign f_u_arrmul24_and19_7_y0 = f_u_arrmul24_and19_7_a_19 & f_u_arrmul24_and19_7_b_7;
  assign f_u_arrmul24_fa19_7_f_u_arrmul24_and19_7_y0 = f_u_arrmul24_and19_7_y0;
  assign f_u_arrmul24_fa19_7_f_u_arrmul24_fa20_6_y2 = f_u_arrmul24_fa20_6_y2;
  assign f_u_arrmul24_fa19_7_f_u_arrmul24_fa18_7_y4 = f_u_arrmul24_fa18_7_y4;
  assign f_u_arrmul24_fa19_7_y0 = f_u_arrmul24_fa19_7_f_u_arrmul24_and19_7_y0 ^ f_u_arrmul24_fa19_7_f_u_arrmul24_fa20_6_y2;
  assign f_u_arrmul24_fa19_7_y1 = f_u_arrmul24_fa19_7_f_u_arrmul24_and19_7_y0 & f_u_arrmul24_fa19_7_f_u_arrmul24_fa20_6_y2;
  assign f_u_arrmul24_fa19_7_y2 = f_u_arrmul24_fa19_7_y0 ^ f_u_arrmul24_fa19_7_f_u_arrmul24_fa18_7_y4;
  assign f_u_arrmul24_fa19_7_y3 = f_u_arrmul24_fa19_7_y0 & f_u_arrmul24_fa19_7_f_u_arrmul24_fa18_7_y4;
  assign f_u_arrmul24_fa19_7_y4 = f_u_arrmul24_fa19_7_y1 | f_u_arrmul24_fa19_7_y3;
  assign f_u_arrmul24_and20_7_a_20 = a_20;
  assign f_u_arrmul24_and20_7_b_7 = b_7;
  assign f_u_arrmul24_and20_7_y0 = f_u_arrmul24_and20_7_a_20 & f_u_arrmul24_and20_7_b_7;
  assign f_u_arrmul24_fa20_7_f_u_arrmul24_and20_7_y0 = f_u_arrmul24_and20_7_y0;
  assign f_u_arrmul24_fa20_7_f_u_arrmul24_fa21_6_y2 = f_u_arrmul24_fa21_6_y2;
  assign f_u_arrmul24_fa20_7_f_u_arrmul24_fa19_7_y4 = f_u_arrmul24_fa19_7_y4;
  assign f_u_arrmul24_fa20_7_y0 = f_u_arrmul24_fa20_7_f_u_arrmul24_and20_7_y0 ^ f_u_arrmul24_fa20_7_f_u_arrmul24_fa21_6_y2;
  assign f_u_arrmul24_fa20_7_y1 = f_u_arrmul24_fa20_7_f_u_arrmul24_and20_7_y0 & f_u_arrmul24_fa20_7_f_u_arrmul24_fa21_6_y2;
  assign f_u_arrmul24_fa20_7_y2 = f_u_arrmul24_fa20_7_y0 ^ f_u_arrmul24_fa20_7_f_u_arrmul24_fa19_7_y4;
  assign f_u_arrmul24_fa20_7_y3 = f_u_arrmul24_fa20_7_y0 & f_u_arrmul24_fa20_7_f_u_arrmul24_fa19_7_y4;
  assign f_u_arrmul24_fa20_7_y4 = f_u_arrmul24_fa20_7_y1 | f_u_arrmul24_fa20_7_y3;
  assign f_u_arrmul24_and21_7_a_21 = a_21;
  assign f_u_arrmul24_and21_7_b_7 = b_7;
  assign f_u_arrmul24_and21_7_y0 = f_u_arrmul24_and21_7_a_21 & f_u_arrmul24_and21_7_b_7;
  assign f_u_arrmul24_fa21_7_f_u_arrmul24_and21_7_y0 = f_u_arrmul24_and21_7_y0;
  assign f_u_arrmul24_fa21_7_f_u_arrmul24_fa22_6_y2 = f_u_arrmul24_fa22_6_y2;
  assign f_u_arrmul24_fa21_7_f_u_arrmul24_fa20_7_y4 = f_u_arrmul24_fa20_7_y4;
  assign f_u_arrmul24_fa21_7_y0 = f_u_arrmul24_fa21_7_f_u_arrmul24_and21_7_y0 ^ f_u_arrmul24_fa21_7_f_u_arrmul24_fa22_6_y2;
  assign f_u_arrmul24_fa21_7_y1 = f_u_arrmul24_fa21_7_f_u_arrmul24_and21_7_y0 & f_u_arrmul24_fa21_7_f_u_arrmul24_fa22_6_y2;
  assign f_u_arrmul24_fa21_7_y2 = f_u_arrmul24_fa21_7_y0 ^ f_u_arrmul24_fa21_7_f_u_arrmul24_fa20_7_y4;
  assign f_u_arrmul24_fa21_7_y3 = f_u_arrmul24_fa21_7_y0 & f_u_arrmul24_fa21_7_f_u_arrmul24_fa20_7_y4;
  assign f_u_arrmul24_fa21_7_y4 = f_u_arrmul24_fa21_7_y1 | f_u_arrmul24_fa21_7_y3;
  assign f_u_arrmul24_and22_7_a_22 = a_22;
  assign f_u_arrmul24_and22_7_b_7 = b_7;
  assign f_u_arrmul24_and22_7_y0 = f_u_arrmul24_and22_7_a_22 & f_u_arrmul24_and22_7_b_7;
  assign f_u_arrmul24_fa22_7_f_u_arrmul24_and22_7_y0 = f_u_arrmul24_and22_7_y0;
  assign f_u_arrmul24_fa22_7_f_u_arrmul24_fa23_6_y2 = f_u_arrmul24_fa23_6_y2;
  assign f_u_arrmul24_fa22_7_f_u_arrmul24_fa21_7_y4 = f_u_arrmul24_fa21_7_y4;
  assign f_u_arrmul24_fa22_7_y0 = f_u_arrmul24_fa22_7_f_u_arrmul24_and22_7_y0 ^ f_u_arrmul24_fa22_7_f_u_arrmul24_fa23_6_y2;
  assign f_u_arrmul24_fa22_7_y1 = f_u_arrmul24_fa22_7_f_u_arrmul24_and22_7_y0 & f_u_arrmul24_fa22_7_f_u_arrmul24_fa23_6_y2;
  assign f_u_arrmul24_fa22_7_y2 = f_u_arrmul24_fa22_7_y0 ^ f_u_arrmul24_fa22_7_f_u_arrmul24_fa21_7_y4;
  assign f_u_arrmul24_fa22_7_y3 = f_u_arrmul24_fa22_7_y0 & f_u_arrmul24_fa22_7_f_u_arrmul24_fa21_7_y4;
  assign f_u_arrmul24_fa22_7_y4 = f_u_arrmul24_fa22_7_y1 | f_u_arrmul24_fa22_7_y3;
  assign f_u_arrmul24_and23_7_a_23 = a_23;
  assign f_u_arrmul24_and23_7_b_7 = b_7;
  assign f_u_arrmul24_and23_7_y0 = f_u_arrmul24_and23_7_a_23 & f_u_arrmul24_and23_7_b_7;
  assign f_u_arrmul24_fa23_7_f_u_arrmul24_and23_7_y0 = f_u_arrmul24_and23_7_y0;
  assign f_u_arrmul24_fa23_7_f_u_arrmul24_fa23_6_y4 = f_u_arrmul24_fa23_6_y4;
  assign f_u_arrmul24_fa23_7_f_u_arrmul24_fa22_7_y4 = f_u_arrmul24_fa22_7_y4;
  assign f_u_arrmul24_fa23_7_y0 = f_u_arrmul24_fa23_7_f_u_arrmul24_and23_7_y0 ^ f_u_arrmul24_fa23_7_f_u_arrmul24_fa23_6_y4;
  assign f_u_arrmul24_fa23_7_y1 = f_u_arrmul24_fa23_7_f_u_arrmul24_and23_7_y0 & f_u_arrmul24_fa23_7_f_u_arrmul24_fa23_6_y4;
  assign f_u_arrmul24_fa23_7_y2 = f_u_arrmul24_fa23_7_y0 ^ f_u_arrmul24_fa23_7_f_u_arrmul24_fa22_7_y4;
  assign f_u_arrmul24_fa23_7_y3 = f_u_arrmul24_fa23_7_y0 & f_u_arrmul24_fa23_7_f_u_arrmul24_fa22_7_y4;
  assign f_u_arrmul24_fa23_7_y4 = f_u_arrmul24_fa23_7_y1 | f_u_arrmul24_fa23_7_y3;
  assign f_u_arrmul24_and0_8_a_0 = a_0;
  assign f_u_arrmul24_and0_8_b_8 = b_8;
  assign f_u_arrmul24_and0_8_y0 = f_u_arrmul24_and0_8_a_0 & f_u_arrmul24_and0_8_b_8;
  assign f_u_arrmul24_ha0_8_f_u_arrmul24_and0_8_y0 = f_u_arrmul24_and0_8_y0;
  assign f_u_arrmul24_ha0_8_f_u_arrmul24_fa1_7_y2 = f_u_arrmul24_fa1_7_y2;
  assign f_u_arrmul24_ha0_8_y0 = f_u_arrmul24_ha0_8_f_u_arrmul24_and0_8_y0 ^ f_u_arrmul24_ha0_8_f_u_arrmul24_fa1_7_y2;
  assign f_u_arrmul24_ha0_8_y1 = f_u_arrmul24_ha0_8_f_u_arrmul24_and0_8_y0 & f_u_arrmul24_ha0_8_f_u_arrmul24_fa1_7_y2;
  assign f_u_arrmul24_and1_8_a_1 = a_1;
  assign f_u_arrmul24_and1_8_b_8 = b_8;
  assign f_u_arrmul24_and1_8_y0 = f_u_arrmul24_and1_8_a_1 & f_u_arrmul24_and1_8_b_8;
  assign f_u_arrmul24_fa1_8_f_u_arrmul24_and1_8_y0 = f_u_arrmul24_and1_8_y0;
  assign f_u_arrmul24_fa1_8_f_u_arrmul24_fa2_7_y2 = f_u_arrmul24_fa2_7_y2;
  assign f_u_arrmul24_fa1_8_f_u_arrmul24_ha0_8_y1 = f_u_arrmul24_ha0_8_y1;
  assign f_u_arrmul24_fa1_8_y0 = f_u_arrmul24_fa1_8_f_u_arrmul24_and1_8_y0 ^ f_u_arrmul24_fa1_8_f_u_arrmul24_fa2_7_y2;
  assign f_u_arrmul24_fa1_8_y1 = f_u_arrmul24_fa1_8_f_u_arrmul24_and1_8_y0 & f_u_arrmul24_fa1_8_f_u_arrmul24_fa2_7_y2;
  assign f_u_arrmul24_fa1_8_y2 = f_u_arrmul24_fa1_8_y0 ^ f_u_arrmul24_fa1_8_f_u_arrmul24_ha0_8_y1;
  assign f_u_arrmul24_fa1_8_y3 = f_u_arrmul24_fa1_8_y0 & f_u_arrmul24_fa1_8_f_u_arrmul24_ha0_8_y1;
  assign f_u_arrmul24_fa1_8_y4 = f_u_arrmul24_fa1_8_y1 | f_u_arrmul24_fa1_8_y3;
  assign f_u_arrmul24_and2_8_a_2 = a_2;
  assign f_u_arrmul24_and2_8_b_8 = b_8;
  assign f_u_arrmul24_and2_8_y0 = f_u_arrmul24_and2_8_a_2 & f_u_arrmul24_and2_8_b_8;
  assign f_u_arrmul24_fa2_8_f_u_arrmul24_and2_8_y0 = f_u_arrmul24_and2_8_y0;
  assign f_u_arrmul24_fa2_8_f_u_arrmul24_fa3_7_y2 = f_u_arrmul24_fa3_7_y2;
  assign f_u_arrmul24_fa2_8_f_u_arrmul24_fa1_8_y4 = f_u_arrmul24_fa1_8_y4;
  assign f_u_arrmul24_fa2_8_y0 = f_u_arrmul24_fa2_8_f_u_arrmul24_and2_8_y0 ^ f_u_arrmul24_fa2_8_f_u_arrmul24_fa3_7_y2;
  assign f_u_arrmul24_fa2_8_y1 = f_u_arrmul24_fa2_8_f_u_arrmul24_and2_8_y0 & f_u_arrmul24_fa2_8_f_u_arrmul24_fa3_7_y2;
  assign f_u_arrmul24_fa2_8_y2 = f_u_arrmul24_fa2_8_y0 ^ f_u_arrmul24_fa2_8_f_u_arrmul24_fa1_8_y4;
  assign f_u_arrmul24_fa2_8_y3 = f_u_arrmul24_fa2_8_y0 & f_u_arrmul24_fa2_8_f_u_arrmul24_fa1_8_y4;
  assign f_u_arrmul24_fa2_8_y4 = f_u_arrmul24_fa2_8_y1 | f_u_arrmul24_fa2_8_y3;
  assign f_u_arrmul24_and3_8_a_3 = a_3;
  assign f_u_arrmul24_and3_8_b_8 = b_8;
  assign f_u_arrmul24_and3_8_y0 = f_u_arrmul24_and3_8_a_3 & f_u_arrmul24_and3_8_b_8;
  assign f_u_arrmul24_fa3_8_f_u_arrmul24_and3_8_y0 = f_u_arrmul24_and3_8_y0;
  assign f_u_arrmul24_fa3_8_f_u_arrmul24_fa4_7_y2 = f_u_arrmul24_fa4_7_y2;
  assign f_u_arrmul24_fa3_8_f_u_arrmul24_fa2_8_y4 = f_u_arrmul24_fa2_8_y4;
  assign f_u_arrmul24_fa3_8_y0 = f_u_arrmul24_fa3_8_f_u_arrmul24_and3_8_y0 ^ f_u_arrmul24_fa3_8_f_u_arrmul24_fa4_7_y2;
  assign f_u_arrmul24_fa3_8_y1 = f_u_arrmul24_fa3_8_f_u_arrmul24_and3_8_y0 & f_u_arrmul24_fa3_8_f_u_arrmul24_fa4_7_y2;
  assign f_u_arrmul24_fa3_8_y2 = f_u_arrmul24_fa3_8_y0 ^ f_u_arrmul24_fa3_8_f_u_arrmul24_fa2_8_y4;
  assign f_u_arrmul24_fa3_8_y3 = f_u_arrmul24_fa3_8_y0 & f_u_arrmul24_fa3_8_f_u_arrmul24_fa2_8_y4;
  assign f_u_arrmul24_fa3_8_y4 = f_u_arrmul24_fa3_8_y1 | f_u_arrmul24_fa3_8_y3;
  assign f_u_arrmul24_and4_8_a_4 = a_4;
  assign f_u_arrmul24_and4_8_b_8 = b_8;
  assign f_u_arrmul24_and4_8_y0 = f_u_arrmul24_and4_8_a_4 & f_u_arrmul24_and4_8_b_8;
  assign f_u_arrmul24_fa4_8_f_u_arrmul24_and4_8_y0 = f_u_arrmul24_and4_8_y0;
  assign f_u_arrmul24_fa4_8_f_u_arrmul24_fa5_7_y2 = f_u_arrmul24_fa5_7_y2;
  assign f_u_arrmul24_fa4_8_f_u_arrmul24_fa3_8_y4 = f_u_arrmul24_fa3_8_y4;
  assign f_u_arrmul24_fa4_8_y0 = f_u_arrmul24_fa4_8_f_u_arrmul24_and4_8_y0 ^ f_u_arrmul24_fa4_8_f_u_arrmul24_fa5_7_y2;
  assign f_u_arrmul24_fa4_8_y1 = f_u_arrmul24_fa4_8_f_u_arrmul24_and4_8_y0 & f_u_arrmul24_fa4_8_f_u_arrmul24_fa5_7_y2;
  assign f_u_arrmul24_fa4_8_y2 = f_u_arrmul24_fa4_8_y0 ^ f_u_arrmul24_fa4_8_f_u_arrmul24_fa3_8_y4;
  assign f_u_arrmul24_fa4_8_y3 = f_u_arrmul24_fa4_8_y0 & f_u_arrmul24_fa4_8_f_u_arrmul24_fa3_8_y4;
  assign f_u_arrmul24_fa4_8_y4 = f_u_arrmul24_fa4_8_y1 | f_u_arrmul24_fa4_8_y3;
  assign f_u_arrmul24_and5_8_a_5 = a_5;
  assign f_u_arrmul24_and5_8_b_8 = b_8;
  assign f_u_arrmul24_and5_8_y0 = f_u_arrmul24_and5_8_a_5 & f_u_arrmul24_and5_8_b_8;
  assign f_u_arrmul24_fa5_8_f_u_arrmul24_and5_8_y0 = f_u_arrmul24_and5_8_y0;
  assign f_u_arrmul24_fa5_8_f_u_arrmul24_fa6_7_y2 = f_u_arrmul24_fa6_7_y2;
  assign f_u_arrmul24_fa5_8_f_u_arrmul24_fa4_8_y4 = f_u_arrmul24_fa4_8_y4;
  assign f_u_arrmul24_fa5_8_y0 = f_u_arrmul24_fa5_8_f_u_arrmul24_and5_8_y0 ^ f_u_arrmul24_fa5_8_f_u_arrmul24_fa6_7_y2;
  assign f_u_arrmul24_fa5_8_y1 = f_u_arrmul24_fa5_8_f_u_arrmul24_and5_8_y0 & f_u_arrmul24_fa5_8_f_u_arrmul24_fa6_7_y2;
  assign f_u_arrmul24_fa5_8_y2 = f_u_arrmul24_fa5_8_y0 ^ f_u_arrmul24_fa5_8_f_u_arrmul24_fa4_8_y4;
  assign f_u_arrmul24_fa5_8_y3 = f_u_arrmul24_fa5_8_y0 & f_u_arrmul24_fa5_8_f_u_arrmul24_fa4_8_y4;
  assign f_u_arrmul24_fa5_8_y4 = f_u_arrmul24_fa5_8_y1 | f_u_arrmul24_fa5_8_y3;
  assign f_u_arrmul24_and6_8_a_6 = a_6;
  assign f_u_arrmul24_and6_8_b_8 = b_8;
  assign f_u_arrmul24_and6_8_y0 = f_u_arrmul24_and6_8_a_6 & f_u_arrmul24_and6_8_b_8;
  assign f_u_arrmul24_fa6_8_f_u_arrmul24_and6_8_y0 = f_u_arrmul24_and6_8_y0;
  assign f_u_arrmul24_fa6_8_f_u_arrmul24_fa7_7_y2 = f_u_arrmul24_fa7_7_y2;
  assign f_u_arrmul24_fa6_8_f_u_arrmul24_fa5_8_y4 = f_u_arrmul24_fa5_8_y4;
  assign f_u_arrmul24_fa6_8_y0 = f_u_arrmul24_fa6_8_f_u_arrmul24_and6_8_y0 ^ f_u_arrmul24_fa6_8_f_u_arrmul24_fa7_7_y2;
  assign f_u_arrmul24_fa6_8_y1 = f_u_arrmul24_fa6_8_f_u_arrmul24_and6_8_y0 & f_u_arrmul24_fa6_8_f_u_arrmul24_fa7_7_y2;
  assign f_u_arrmul24_fa6_8_y2 = f_u_arrmul24_fa6_8_y0 ^ f_u_arrmul24_fa6_8_f_u_arrmul24_fa5_8_y4;
  assign f_u_arrmul24_fa6_8_y3 = f_u_arrmul24_fa6_8_y0 & f_u_arrmul24_fa6_8_f_u_arrmul24_fa5_8_y4;
  assign f_u_arrmul24_fa6_8_y4 = f_u_arrmul24_fa6_8_y1 | f_u_arrmul24_fa6_8_y3;
  assign f_u_arrmul24_and7_8_a_7 = a_7;
  assign f_u_arrmul24_and7_8_b_8 = b_8;
  assign f_u_arrmul24_and7_8_y0 = f_u_arrmul24_and7_8_a_7 & f_u_arrmul24_and7_8_b_8;
  assign f_u_arrmul24_fa7_8_f_u_arrmul24_and7_8_y0 = f_u_arrmul24_and7_8_y0;
  assign f_u_arrmul24_fa7_8_f_u_arrmul24_fa8_7_y2 = f_u_arrmul24_fa8_7_y2;
  assign f_u_arrmul24_fa7_8_f_u_arrmul24_fa6_8_y4 = f_u_arrmul24_fa6_8_y4;
  assign f_u_arrmul24_fa7_8_y0 = f_u_arrmul24_fa7_8_f_u_arrmul24_and7_8_y0 ^ f_u_arrmul24_fa7_8_f_u_arrmul24_fa8_7_y2;
  assign f_u_arrmul24_fa7_8_y1 = f_u_arrmul24_fa7_8_f_u_arrmul24_and7_8_y0 & f_u_arrmul24_fa7_8_f_u_arrmul24_fa8_7_y2;
  assign f_u_arrmul24_fa7_8_y2 = f_u_arrmul24_fa7_8_y0 ^ f_u_arrmul24_fa7_8_f_u_arrmul24_fa6_8_y4;
  assign f_u_arrmul24_fa7_8_y3 = f_u_arrmul24_fa7_8_y0 & f_u_arrmul24_fa7_8_f_u_arrmul24_fa6_8_y4;
  assign f_u_arrmul24_fa7_8_y4 = f_u_arrmul24_fa7_8_y1 | f_u_arrmul24_fa7_8_y3;
  assign f_u_arrmul24_and8_8_a_8 = a_8;
  assign f_u_arrmul24_and8_8_b_8 = b_8;
  assign f_u_arrmul24_and8_8_y0 = f_u_arrmul24_and8_8_a_8 & f_u_arrmul24_and8_8_b_8;
  assign f_u_arrmul24_fa8_8_f_u_arrmul24_and8_8_y0 = f_u_arrmul24_and8_8_y0;
  assign f_u_arrmul24_fa8_8_f_u_arrmul24_fa9_7_y2 = f_u_arrmul24_fa9_7_y2;
  assign f_u_arrmul24_fa8_8_f_u_arrmul24_fa7_8_y4 = f_u_arrmul24_fa7_8_y4;
  assign f_u_arrmul24_fa8_8_y0 = f_u_arrmul24_fa8_8_f_u_arrmul24_and8_8_y0 ^ f_u_arrmul24_fa8_8_f_u_arrmul24_fa9_7_y2;
  assign f_u_arrmul24_fa8_8_y1 = f_u_arrmul24_fa8_8_f_u_arrmul24_and8_8_y0 & f_u_arrmul24_fa8_8_f_u_arrmul24_fa9_7_y2;
  assign f_u_arrmul24_fa8_8_y2 = f_u_arrmul24_fa8_8_y0 ^ f_u_arrmul24_fa8_8_f_u_arrmul24_fa7_8_y4;
  assign f_u_arrmul24_fa8_8_y3 = f_u_arrmul24_fa8_8_y0 & f_u_arrmul24_fa8_8_f_u_arrmul24_fa7_8_y4;
  assign f_u_arrmul24_fa8_8_y4 = f_u_arrmul24_fa8_8_y1 | f_u_arrmul24_fa8_8_y3;
  assign f_u_arrmul24_and9_8_a_9 = a_9;
  assign f_u_arrmul24_and9_8_b_8 = b_8;
  assign f_u_arrmul24_and9_8_y0 = f_u_arrmul24_and9_8_a_9 & f_u_arrmul24_and9_8_b_8;
  assign f_u_arrmul24_fa9_8_f_u_arrmul24_and9_8_y0 = f_u_arrmul24_and9_8_y0;
  assign f_u_arrmul24_fa9_8_f_u_arrmul24_fa10_7_y2 = f_u_arrmul24_fa10_7_y2;
  assign f_u_arrmul24_fa9_8_f_u_arrmul24_fa8_8_y4 = f_u_arrmul24_fa8_8_y4;
  assign f_u_arrmul24_fa9_8_y0 = f_u_arrmul24_fa9_8_f_u_arrmul24_and9_8_y0 ^ f_u_arrmul24_fa9_8_f_u_arrmul24_fa10_7_y2;
  assign f_u_arrmul24_fa9_8_y1 = f_u_arrmul24_fa9_8_f_u_arrmul24_and9_8_y0 & f_u_arrmul24_fa9_8_f_u_arrmul24_fa10_7_y2;
  assign f_u_arrmul24_fa9_8_y2 = f_u_arrmul24_fa9_8_y0 ^ f_u_arrmul24_fa9_8_f_u_arrmul24_fa8_8_y4;
  assign f_u_arrmul24_fa9_8_y3 = f_u_arrmul24_fa9_8_y0 & f_u_arrmul24_fa9_8_f_u_arrmul24_fa8_8_y4;
  assign f_u_arrmul24_fa9_8_y4 = f_u_arrmul24_fa9_8_y1 | f_u_arrmul24_fa9_8_y3;
  assign f_u_arrmul24_and10_8_a_10 = a_10;
  assign f_u_arrmul24_and10_8_b_8 = b_8;
  assign f_u_arrmul24_and10_8_y0 = f_u_arrmul24_and10_8_a_10 & f_u_arrmul24_and10_8_b_8;
  assign f_u_arrmul24_fa10_8_f_u_arrmul24_and10_8_y0 = f_u_arrmul24_and10_8_y0;
  assign f_u_arrmul24_fa10_8_f_u_arrmul24_fa11_7_y2 = f_u_arrmul24_fa11_7_y2;
  assign f_u_arrmul24_fa10_8_f_u_arrmul24_fa9_8_y4 = f_u_arrmul24_fa9_8_y4;
  assign f_u_arrmul24_fa10_8_y0 = f_u_arrmul24_fa10_8_f_u_arrmul24_and10_8_y0 ^ f_u_arrmul24_fa10_8_f_u_arrmul24_fa11_7_y2;
  assign f_u_arrmul24_fa10_8_y1 = f_u_arrmul24_fa10_8_f_u_arrmul24_and10_8_y0 & f_u_arrmul24_fa10_8_f_u_arrmul24_fa11_7_y2;
  assign f_u_arrmul24_fa10_8_y2 = f_u_arrmul24_fa10_8_y0 ^ f_u_arrmul24_fa10_8_f_u_arrmul24_fa9_8_y4;
  assign f_u_arrmul24_fa10_8_y3 = f_u_arrmul24_fa10_8_y0 & f_u_arrmul24_fa10_8_f_u_arrmul24_fa9_8_y4;
  assign f_u_arrmul24_fa10_8_y4 = f_u_arrmul24_fa10_8_y1 | f_u_arrmul24_fa10_8_y3;
  assign f_u_arrmul24_and11_8_a_11 = a_11;
  assign f_u_arrmul24_and11_8_b_8 = b_8;
  assign f_u_arrmul24_and11_8_y0 = f_u_arrmul24_and11_8_a_11 & f_u_arrmul24_and11_8_b_8;
  assign f_u_arrmul24_fa11_8_f_u_arrmul24_and11_8_y0 = f_u_arrmul24_and11_8_y0;
  assign f_u_arrmul24_fa11_8_f_u_arrmul24_fa12_7_y2 = f_u_arrmul24_fa12_7_y2;
  assign f_u_arrmul24_fa11_8_f_u_arrmul24_fa10_8_y4 = f_u_arrmul24_fa10_8_y4;
  assign f_u_arrmul24_fa11_8_y0 = f_u_arrmul24_fa11_8_f_u_arrmul24_and11_8_y0 ^ f_u_arrmul24_fa11_8_f_u_arrmul24_fa12_7_y2;
  assign f_u_arrmul24_fa11_8_y1 = f_u_arrmul24_fa11_8_f_u_arrmul24_and11_8_y0 & f_u_arrmul24_fa11_8_f_u_arrmul24_fa12_7_y2;
  assign f_u_arrmul24_fa11_8_y2 = f_u_arrmul24_fa11_8_y0 ^ f_u_arrmul24_fa11_8_f_u_arrmul24_fa10_8_y4;
  assign f_u_arrmul24_fa11_8_y3 = f_u_arrmul24_fa11_8_y0 & f_u_arrmul24_fa11_8_f_u_arrmul24_fa10_8_y4;
  assign f_u_arrmul24_fa11_8_y4 = f_u_arrmul24_fa11_8_y1 | f_u_arrmul24_fa11_8_y3;
  assign f_u_arrmul24_and12_8_a_12 = a_12;
  assign f_u_arrmul24_and12_8_b_8 = b_8;
  assign f_u_arrmul24_and12_8_y0 = f_u_arrmul24_and12_8_a_12 & f_u_arrmul24_and12_8_b_8;
  assign f_u_arrmul24_fa12_8_f_u_arrmul24_and12_8_y0 = f_u_arrmul24_and12_8_y0;
  assign f_u_arrmul24_fa12_8_f_u_arrmul24_fa13_7_y2 = f_u_arrmul24_fa13_7_y2;
  assign f_u_arrmul24_fa12_8_f_u_arrmul24_fa11_8_y4 = f_u_arrmul24_fa11_8_y4;
  assign f_u_arrmul24_fa12_8_y0 = f_u_arrmul24_fa12_8_f_u_arrmul24_and12_8_y0 ^ f_u_arrmul24_fa12_8_f_u_arrmul24_fa13_7_y2;
  assign f_u_arrmul24_fa12_8_y1 = f_u_arrmul24_fa12_8_f_u_arrmul24_and12_8_y0 & f_u_arrmul24_fa12_8_f_u_arrmul24_fa13_7_y2;
  assign f_u_arrmul24_fa12_8_y2 = f_u_arrmul24_fa12_8_y0 ^ f_u_arrmul24_fa12_8_f_u_arrmul24_fa11_8_y4;
  assign f_u_arrmul24_fa12_8_y3 = f_u_arrmul24_fa12_8_y0 & f_u_arrmul24_fa12_8_f_u_arrmul24_fa11_8_y4;
  assign f_u_arrmul24_fa12_8_y4 = f_u_arrmul24_fa12_8_y1 | f_u_arrmul24_fa12_8_y3;
  assign f_u_arrmul24_and13_8_a_13 = a_13;
  assign f_u_arrmul24_and13_8_b_8 = b_8;
  assign f_u_arrmul24_and13_8_y0 = f_u_arrmul24_and13_8_a_13 & f_u_arrmul24_and13_8_b_8;
  assign f_u_arrmul24_fa13_8_f_u_arrmul24_and13_8_y0 = f_u_arrmul24_and13_8_y0;
  assign f_u_arrmul24_fa13_8_f_u_arrmul24_fa14_7_y2 = f_u_arrmul24_fa14_7_y2;
  assign f_u_arrmul24_fa13_8_f_u_arrmul24_fa12_8_y4 = f_u_arrmul24_fa12_8_y4;
  assign f_u_arrmul24_fa13_8_y0 = f_u_arrmul24_fa13_8_f_u_arrmul24_and13_8_y0 ^ f_u_arrmul24_fa13_8_f_u_arrmul24_fa14_7_y2;
  assign f_u_arrmul24_fa13_8_y1 = f_u_arrmul24_fa13_8_f_u_arrmul24_and13_8_y0 & f_u_arrmul24_fa13_8_f_u_arrmul24_fa14_7_y2;
  assign f_u_arrmul24_fa13_8_y2 = f_u_arrmul24_fa13_8_y0 ^ f_u_arrmul24_fa13_8_f_u_arrmul24_fa12_8_y4;
  assign f_u_arrmul24_fa13_8_y3 = f_u_arrmul24_fa13_8_y0 & f_u_arrmul24_fa13_8_f_u_arrmul24_fa12_8_y4;
  assign f_u_arrmul24_fa13_8_y4 = f_u_arrmul24_fa13_8_y1 | f_u_arrmul24_fa13_8_y3;
  assign f_u_arrmul24_and14_8_a_14 = a_14;
  assign f_u_arrmul24_and14_8_b_8 = b_8;
  assign f_u_arrmul24_and14_8_y0 = f_u_arrmul24_and14_8_a_14 & f_u_arrmul24_and14_8_b_8;
  assign f_u_arrmul24_fa14_8_f_u_arrmul24_and14_8_y0 = f_u_arrmul24_and14_8_y0;
  assign f_u_arrmul24_fa14_8_f_u_arrmul24_fa15_7_y2 = f_u_arrmul24_fa15_7_y2;
  assign f_u_arrmul24_fa14_8_f_u_arrmul24_fa13_8_y4 = f_u_arrmul24_fa13_8_y4;
  assign f_u_arrmul24_fa14_8_y0 = f_u_arrmul24_fa14_8_f_u_arrmul24_and14_8_y0 ^ f_u_arrmul24_fa14_8_f_u_arrmul24_fa15_7_y2;
  assign f_u_arrmul24_fa14_8_y1 = f_u_arrmul24_fa14_8_f_u_arrmul24_and14_8_y0 & f_u_arrmul24_fa14_8_f_u_arrmul24_fa15_7_y2;
  assign f_u_arrmul24_fa14_8_y2 = f_u_arrmul24_fa14_8_y0 ^ f_u_arrmul24_fa14_8_f_u_arrmul24_fa13_8_y4;
  assign f_u_arrmul24_fa14_8_y3 = f_u_arrmul24_fa14_8_y0 & f_u_arrmul24_fa14_8_f_u_arrmul24_fa13_8_y4;
  assign f_u_arrmul24_fa14_8_y4 = f_u_arrmul24_fa14_8_y1 | f_u_arrmul24_fa14_8_y3;
  assign f_u_arrmul24_and15_8_a_15 = a_15;
  assign f_u_arrmul24_and15_8_b_8 = b_8;
  assign f_u_arrmul24_and15_8_y0 = f_u_arrmul24_and15_8_a_15 & f_u_arrmul24_and15_8_b_8;
  assign f_u_arrmul24_fa15_8_f_u_arrmul24_and15_8_y0 = f_u_arrmul24_and15_8_y0;
  assign f_u_arrmul24_fa15_8_f_u_arrmul24_fa16_7_y2 = f_u_arrmul24_fa16_7_y2;
  assign f_u_arrmul24_fa15_8_f_u_arrmul24_fa14_8_y4 = f_u_arrmul24_fa14_8_y4;
  assign f_u_arrmul24_fa15_8_y0 = f_u_arrmul24_fa15_8_f_u_arrmul24_and15_8_y0 ^ f_u_arrmul24_fa15_8_f_u_arrmul24_fa16_7_y2;
  assign f_u_arrmul24_fa15_8_y1 = f_u_arrmul24_fa15_8_f_u_arrmul24_and15_8_y0 & f_u_arrmul24_fa15_8_f_u_arrmul24_fa16_7_y2;
  assign f_u_arrmul24_fa15_8_y2 = f_u_arrmul24_fa15_8_y0 ^ f_u_arrmul24_fa15_8_f_u_arrmul24_fa14_8_y4;
  assign f_u_arrmul24_fa15_8_y3 = f_u_arrmul24_fa15_8_y0 & f_u_arrmul24_fa15_8_f_u_arrmul24_fa14_8_y4;
  assign f_u_arrmul24_fa15_8_y4 = f_u_arrmul24_fa15_8_y1 | f_u_arrmul24_fa15_8_y3;
  assign f_u_arrmul24_and16_8_a_16 = a_16;
  assign f_u_arrmul24_and16_8_b_8 = b_8;
  assign f_u_arrmul24_and16_8_y0 = f_u_arrmul24_and16_8_a_16 & f_u_arrmul24_and16_8_b_8;
  assign f_u_arrmul24_fa16_8_f_u_arrmul24_and16_8_y0 = f_u_arrmul24_and16_8_y0;
  assign f_u_arrmul24_fa16_8_f_u_arrmul24_fa17_7_y2 = f_u_arrmul24_fa17_7_y2;
  assign f_u_arrmul24_fa16_8_f_u_arrmul24_fa15_8_y4 = f_u_arrmul24_fa15_8_y4;
  assign f_u_arrmul24_fa16_8_y0 = f_u_arrmul24_fa16_8_f_u_arrmul24_and16_8_y0 ^ f_u_arrmul24_fa16_8_f_u_arrmul24_fa17_7_y2;
  assign f_u_arrmul24_fa16_8_y1 = f_u_arrmul24_fa16_8_f_u_arrmul24_and16_8_y0 & f_u_arrmul24_fa16_8_f_u_arrmul24_fa17_7_y2;
  assign f_u_arrmul24_fa16_8_y2 = f_u_arrmul24_fa16_8_y0 ^ f_u_arrmul24_fa16_8_f_u_arrmul24_fa15_8_y4;
  assign f_u_arrmul24_fa16_8_y3 = f_u_arrmul24_fa16_8_y0 & f_u_arrmul24_fa16_8_f_u_arrmul24_fa15_8_y4;
  assign f_u_arrmul24_fa16_8_y4 = f_u_arrmul24_fa16_8_y1 | f_u_arrmul24_fa16_8_y3;
  assign f_u_arrmul24_and17_8_a_17 = a_17;
  assign f_u_arrmul24_and17_8_b_8 = b_8;
  assign f_u_arrmul24_and17_8_y0 = f_u_arrmul24_and17_8_a_17 & f_u_arrmul24_and17_8_b_8;
  assign f_u_arrmul24_fa17_8_f_u_arrmul24_and17_8_y0 = f_u_arrmul24_and17_8_y0;
  assign f_u_arrmul24_fa17_8_f_u_arrmul24_fa18_7_y2 = f_u_arrmul24_fa18_7_y2;
  assign f_u_arrmul24_fa17_8_f_u_arrmul24_fa16_8_y4 = f_u_arrmul24_fa16_8_y4;
  assign f_u_arrmul24_fa17_8_y0 = f_u_arrmul24_fa17_8_f_u_arrmul24_and17_8_y0 ^ f_u_arrmul24_fa17_8_f_u_arrmul24_fa18_7_y2;
  assign f_u_arrmul24_fa17_8_y1 = f_u_arrmul24_fa17_8_f_u_arrmul24_and17_8_y0 & f_u_arrmul24_fa17_8_f_u_arrmul24_fa18_7_y2;
  assign f_u_arrmul24_fa17_8_y2 = f_u_arrmul24_fa17_8_y0 ^ f_u_arrmul24_fa17_8_f_u_arrmul24_fa16_8_y4;
  assign f_u_arrmul24_fa17_8_y3 = f_u_arrmul24_fa17_8_y0 & f_u_arrmul24_fa17_8_f_u_arrmul24_fa16_8_y4;
  assign f_u_arrmul24_fa17_8_y4 = f_u_arrmul24_fa17_8_y1 | f_u_arrmul24_fa17_8_y3;
  assign f_u_arrmul24_and18_8_a_18 = a_18;
  assign f_u_arrmul24_and18_8_b_8 = b_8;
  assign f_u_arrmul24_and18_8_y0 = f_u_arrmul24_and18_8_a_18 & f_u_arrmul24_and18_8_b_8;
  assign f_u_arrmul24_fa18_8_f_u_arrmul24_and18_8_y0 = f_u_arrmul24_and18_8_y0;
  assign f_u_arrmul24_fa18_8_f_u_arrmul24_fa19_7_y2 = f_u_arrmul24_fa19_7_y2;
  assign f_u_arrmul24_fa18_8_f_u_arrmul24_fa17_8_y4 = f_u_arrmul24_fa17_8_y4;
  assign f_u_arrmul24_fa18_8_y0 = f_u_arrmul24_fa18_8_f_u_arrmul24_and18_8_y0 ^ f_u_arrmul24_fa18_8_f_u_arrmul24_fa19_7_y2;
  assign f_u_arrmul24_fa18_8_y1 = f_u_arrmul24_fa18_8_f_u_arrmul24_and18_8_y0 & f_u_arrmul24_fa18_8_f_u_arrmul24_fa19_7_y2;
  assign f_u_arrmul24_fa18_8_y2 = f_u_arrmul24_fa18_8_y0 ^ f_u_arrmul24_fa18_8_f_u_arrmul24_fa17_8_y4;
  assign f_u_arrmul24_fa18_8_y3 = f_u_arrmul24_fa18_8_y0 & f_u_arrmul24_fa18_8_f_u_arrmul24_fa17_8_y4;
  assign f_u_arrmul24_fa18_8_y4 = f_u_arrmul24_fa18_8_y1 | f_u_arrmul24_fa18_8_y3;
  assign f_u_arrmul24_and19_8_a_19 = a_19;
  assign f_u_arrmul24_and19_8_b_8 = b_8;
  assign f_u_arrmul24_and19_8_y0 = f_u_arrmul24_and19_8_a_19 & f_u_arrmul24_and19_8_b_8;
  assign f_u_arrmul24_fa19_8_f_u_arrmul24_and19_8_y0 = f_u_arrmul24_and19_8_y0;
  assign f_u_arrmul24_fa19_8_f_u_arrmul24_fa20_7_y2 = f_u_arrmul24_fa20_7_y2;
  assign f_u_arrmul24_fa19_8_f_u_arrmul24_fa18_8_y4 = f_u_arrmul24_fa18_8_y4;
  assign f_u_arrmul24_fa19_8_y0 = f_u_arrmul24_fa19_8_f_u_arrmul24_and19_8_y0 ^ f_u_arrmul24_fa19_8_f_u_arrmul24_fa20_7_y2;
  assign f_u_arrmul24_fa19_8_y1 = f_u_arrmul24_fa19_8_f_u_arrmul24_and19_8_y0 & f_u_arrmul24_fa19_8_f_u_arrmul24_fa20_7_y2;
  assign f_u_arrmul24_fa19_8_y2 = f_u_arrmul24_fa19_8_y0 ^ f_u_arrmul24_fa19_8_f_u_arrmul24_fa18_8_y4;
  assign f_u_arrmul24_fa19_8_y3 = f_u_arrmul24_fa19_8_y0 & f_u_arrmul24_fa19_8_f_u_arrmul24_fa18_8_y4;
  assign f_u_arrmul24_fa19_8_y4 = f_u_arrmul24_fa19_8_y1 | f_u_arrmul24_fa19_8_y3;
  assign f_u_arrmul24_and20_8_a_20 = a_20;
  assign f_u_arrmul24_and20_8_b_8 = b_8;
  assign f_u_arrmul24_and20_8_y0 = f_u_arrmul24_and20_8_a_20 & f_u_arrmul24_and20_8_b_8;
  assign f_u_arrmul24_fa20_8_f_u_arrmul24_and20_8_y0 = f_u_arrmul24_and20_8_y0;
  assign f_u_arrmul24_fa20_8_f_u_arrmul24_fa21_7_y2 = f_u_arrmul24_fa21_7_y2;
  assign f_u_arrmul24_fa20_8_f_u_arrmul24_fa19_8_y4 = f_u_arrmul24_fa19_8_y4;
  assign f_u_arrmul24_fa20_8_y0 = f_u_arrmul24_fa20_8_f_u_arrmul24_and20_8_y0 ^ f_u_arrmul24_fa20_8_f_u_arrmul24_fa21_7_y2;
  assign f_u_arrmul24_fa20_8_y1 = f_u_arrmul24_fa20_8_f_u_arrmul24_and20_8_y0 & f_u_arrmul24_fa20_8_f_u_arrmul24_fa21_7_y2;
  assign f_u_arrmul24_fa20_8_y2 = f_u_arrmul24_fa20_8_y0 ^ f_u_arrmul24_fa20_8_f_u_arrmul24_fa19_8_y4;
  assign f_u_arrmul24_fa20_8_y3 = f_u_arrmul24_fa20_8_y0 & f_u_arrmul24_fa20_8_f_u_arrmul24_fa19_8_y4;
  assign f_u_arrmul24_fa20_8_y4 = f_u_arrmul24_fa20_8_y1 | f_u_arrmul24_fa20_8_y3;
  assign f_u_arrmul24_and21_8_a_21 = a_21;
  assign f_u_arrmul24_and21_8_b_8 = b_8;
  assign f_u_arrmul24_and21_8_y0 = f_u_arrmul24_and21_8_a_21 & f_u_arrmul24_and21_8_b_8;
  assign f_u_arrmul24_fa21_8_f_u_arrmul24_and21_8_y0 = f_u_arrmul24_and21_8_y0;
  assign f_u_arrmul24_fa21_8_f_u_arrmul24_fa22_7_y2 = f_u_arrmul24_fa22_7_y2;
  assign f_u_arrmul24_fa21_8_f_u_arrmul24_fa20_8_y4 = f_u_arrmul24_fa20_8_y4;
  assign f_u_arrmul24_fa21_8_y0 = f_u_arrmul24_fa21_8_f_u_arrmul24_and21_8_y0 ^ f_u_arrmul24_fa21_8_f_u_arrmul24_fa22_7_y2;
  assign f_u_arrmul24_fa21_8_y1 = f_u_arrmul24_fa21_8_f_u_arrmul24_and21_8_y0 & f_u_arrmul24_fa21_8_f_u_arrmul24_fa22_7_y2;
  assign f_u_arrmul24_fa21_8_y2 = f_u_arrmul24_fa21_8_y0 ^ f_u_arrmul24_fa21_8_f_u_arrmul24_fa20_8_y4;
  assign f_u_arrmul24_fa21_8_y3 = f_u_arrmul24_fa21_8_y0 & f_u_arrmul24_fa21_8_f_u_arrmul24_fa20_8_y4;
  assign f_u_arrmul24_fa21_8_y4 = f_u_arrmul24_fa21_8_y1 | f_u_arrmul24_fa21_8_y3;
  assign f_u_arrmul24_and22_8_a_22 = a_22;
  assign f_u_arrmul24_and22_8_b_8 = b_8;
  assign f_u_arrmul24_and22_8_y0 = f_u_arrmul24_and22_8_a_22 & f_u_arrmul24_and22_8_b_8;
  assign f_u_arrmul24_fa22_8_f_u_arrmul24_and22_8_y0 = f_u_arrmul24_and22_8_y0;
  assign f_u_arrmul24_fa22_8_f_u_arrmul24_fa23_7_y2 = f_u_arrmul24_fa23_7_y2;
  assign f_u_arrmul24_fa22_8_f_u_arrmul24_fa21_8_y4 = f_u_arrmul24_fa21_8_y4;
  assign f_u_arrmul24_fa22_8_y0 = f_u_arrmul24_fa22_8_f_u_arrmul24_and22_8_y0 ^ f_u_arrmul24_fa22_8_f_u_arrmul24_fa23_7_y2;
  assign f_u_arrmul24_fa22_8_y1 = f_u_arrmul24_fa22_8_f_u_arrmul24_and22_8_y0 & f_u_arrmul24_fa22_8_f_u_arrmul24_fa23_7_y2;
  assign f_u_arrmul24_fa22_8_y2 = f_u_arrmul24_fa22_8_y0 ^ f_u_arrmul24_fa22_8_f_u_arrmul24_fa21_8_y4;
  assign f_u_arrmul24_fa22_8_y3 = f_u_arrmul24_fa22_8_y0 & f_u_arrmul24_fa22_8_f_u_arrmul24_fa21_8_y4;
  assign f_u_arrmul24_fa22_8_y4 = f_u_arrmul24_fa22_8_y1 | f_u_arrmul24_fa22_8_y3;
  assign f_u_arrmul24_and23_8_a_23 = a_23;
  assign f_u_arrmul24_and23_8_b_8 = b_8;
  assign f_u_arrmul24_and23_8_y0 = f_u_arrmul24_and23_8_a_23 & f_u_arrmul24_and23_8_b_8;
  assign f_u_arrmul24_fa23_8_f_u_arrmul24_and23_8_y0 = f_u_arrmul24_and23_8_y0;
  assign f_u_arrmul24_fa23_8_f_u_arrmul24_fa23_7_y4 = f_u_arrmul24_fa23_7_y4;
  assign f_u_arrmul24_fa23_8_f_u_arrmul24_fa22_8_y4 = f_u_arrmul24_fa22_8_y4;
  assign f_u_arrmul24_fa23_8_y0 = f_u_arrmul24_fa23_8_f_u_arrmul24_and23_8_y0 ^ f_u_arrmul24_fa23_8_f_u_arrmul24_fa23_7_y4;
  assign f_u_arrmul24_fa23_8_y1 = f_u_arrmul24_fa23_8_f_u_arrmul24_and23_8_y0 & f_u_arrmul24_fa23_8_f_u_arrmul24_fa23_7_y4;
  assign f_u_arrmul24_fa23_8_y2 = f_u_arrmul24_fa23_8_y0 ^ f_u_arrmul24_fa23_8_f_u_arrmul24_fa22_8_y4;
  assign f_u_arrmul24_fa23_8_y3 = f_u_arrmul24_fa23_8_y0 & f_u_arrmul24_fa23_8_f_u_arrmul24_fa22_8_y4;
  assign f_u_arrmul24_fa23_8_y4 = f_u_arrmul24_fa23_8_y1 | f_u_arrmul24_fa23_8_y3;
  assign f_u_arrmul24_and0_9_a_0 = a_0;
  assign f_u_arrmul24_and0_9_b_9 = b_9;
  assign f_u_arrmul24_and0_9_y0 = f_u_arrmul24_and0_9_a_0 & f_u_arrmul24_and0_9_b_9;
  assign f_u_arrmul24_ha0_9_f_u_arrmul24_and0_9_y0 = f_u_arrmul24_and0_9_y0;
  assign f_u_arrmul24_ha0_9_f_u_arrmul24_fa1_8_y2 = f_u_arrmul24_fa1_8_y2;
  assign f_u_arrmul24_ha0_9_y0 = f_u_arrmul24_ha0_9_f_u_arrmul24_and0_9_y0 ^ f_u_arrmul24_ha0_9_f_u_arrmul24_fa1_8_y2;
  assign f_u_arrmul24_ha0_9_y1 = f_u_arrmul24_ha0_9_f_u_arrmul24_and0_9_y0 & f_u_arrmul24_ha0_9_f_u_arrmul24_fa1_8_y2;
  assign f_u_arrmul24_and1_9_a_1 = a_1;
  assign f_u_arrmul24_and1_9_b_9 = b_9;
  assign f_u_arrmul24_and1_9_y0 = f_u_arrmul24_and1_9_a_1 & f_u_arrmul24_and1_9_b_9;
  assign f_u_arrmul24_fa1_9_f_u_arrmul24_and1_9_y0 = f_u_arrmul24_and1_9_y0;
  assign f_u_arrmul24_fa1_9_f_u_arrmul24_fa2_8_y2 = f_u_arrmul24_fa2_8_y2;
  assign f_u_arrmul24_fa1_9_f_u_arrmul24_ha0_9_y1 = f_u_arrmul24_ha0_9_y1;
  assign f_u_arrmul24_fa1_9_y0 = f_u_arrmul24_fa1_9_f_u_arrmul24_and1_9_y0 ^ f_u_arrmul24_fa1_9_f_u_arrmul24_fa2_8_y2;
  assign f_u_arrmul24_fa1_9_y1 = f_u_arrmul24_fa1_9_f_u_arrmul24_and1_9_y0 & f_u_arrmul24_fa1_9_f_u_arrmul24_fa2_8_y2;
  assign f_u_arrmul24_fa1_9_y2 = f_u_arrmul24_fa1_9_y0 ^ f_u_arrmul24_fa1_9_f_u_arrmul24_ha0_9_y1;
  assign f_u_arrmul24_fa1_9_y3 = f_u_arrmul24_fa1_9_y0 & f_u_arrmul24_fa1_9_f_u_arrmul24_ha0_9_y1;
  assign f_u_arrmul24_fa1_9_y4 = f_u_arrmul24_fa1_9_y1 | f_u_arrmul24_fa1_9_y3;
  assign f_u_arrmul24_and2_9_a_2 = a_2;
  assign f_u_arrmul24_and2_9_b_9 = b_9;
  assign f_u_arrmul24_and2_9_y0 = f_u_arrmul24_and2_9_a_2 & f_u_arrmul24_and2_9_b_9;
  assign f_u_arrmul24_fa2_9_f_u_arrmul24_and2_9_y0 = f_u_arrmul24_and2_9_y0;
  assign f_u_arrmul24_fa2_9_f_u_arrmul24_fa3_8_y2 = f_u_arrmul24_fa3_8_y2;
  assign f_u_arrmul24_fa2_9_f_u_arrmul24_fa1_9_y4 = f_u_arrmul24_fa1_9_y4;
  assign f_u_arrmul24_fa2_9_y0 = f_u_arrmul24_fa2_9_f_u_arrmul24_and2_9_y0 ^ f_u_arrmul24_fa2_9_f_u_arrmul24_fa3_8_y2;
  assign f_u_arrmul24_fa2_9_y1 = f_u_arrmul24_fa2_9_f_u_arrmul24_and2_9_y0 & f_u_arrmul24_fa2_9_f_u_arrmul24_fa3_8_y2;
  assign f_u_arrmul24_fa2_9_y2 = f_u_arrmul24_fa2_9_y0 ^ f_u_arrmul24_fa2_9_f_u_arrmul24_fa1_9_y4;
  assign f_u_arrmul24_fa2_9_y3 = f_u_arrmul24_fa2_9_y0 & f_u_arrmul24_fa2_9_f_u_arrmul24_fa1_9_y4;
  assign f_u_arrmul24_fa2_9_y4 = f_u_arrmul24_fa2_9_y1 | f_u_arrmul24_fa2_9_y3;
  assign f_u_arrmul24_and3_9_a_3 = a_3;
  assign f_u_arrmul24_and3_9_b_9 = b_9;
  assign f_u_arrmul24_and3_9_y0 = f_u_arrmul24_and3_9_a_3 & f_u_arrmul24_and3_9_b_9;
  assign f_u_arrmul24_fa3_9_f_u_arrmul24_and3_9_y0 = f_u_arrmul24_and3_9_y0;
  assign f_u_arrmul24_fa3_9_f_u_arrmul24_fa4_8_y2 = f_u_arrmul24_fa4_8_y2;
  assign f_u_arrmul24_fa3_9_f_u_arrmul24_fa2_9_y4 = f_u_arrmul24_fa2_9_y4;
  assign f_u_arrmul24_fa3_9_y0 = f_u_arrmul24_fa3_9_f_u_arrmul24_and3_9_y0 ^ f_u_arrmul24_fa3_9_f_u_arrmul24_fa4_8_y2;
  assign f_u_arrmul24_fa3_9_y1 = f_u_arrmul24_fa3_9_f_u_arrmul24_and3_9_y0 & f_u_arrmul24_fa3_9_f_u_arrmul24_fa4_8_y2;
  assign f_u_arrmul24_fa3_9_y2 = f_u_arrmul24_fa3_9_y0 ^ f_u_arrmul24_fa3_9_f_u_arrmul24_fa2_9_y4;
  assign f_u_arrmul24_fa3_9_y3 = f_u_arrmul24_fa3_9_y0 & f_u_arrmul24_fa3_9_f_u_arrmul24_fa2_9_y4;
  assign f_u_arrmul24_fa3_9_y4 = f_u_arrmul24_fa3_9_y1 | f_u_arrmul24_fa3_9_y3;
  assign f_u_arrmul24_and4_9_a_4 = a_4;
  assign f_u_arrmul24_and4_9_b_9 = b_9;
  assign f_u_arrmul24_and4_9_y0 = f_u_arrmul24_and4_9_a_4 & f_u_arrmul24_and4_9_b_9;
  assign f_u_arrmul24_fa4_9_f_u_arrmul24_and4_9_y0 = f_u_arrmul24_and4_9_y0;
  assign f_u_arrmul24_fa4_9_f_u_arrmul24_fa5_8_y2 = f_u_arrmul24_fa5_8_y2;
  assign f_u_arrmul24_fa4_9_f_u_arrmul24_fa3_9_y4 = f_u_arrmul24_fa3_9_y4;
  assign f_u_arrmul24_fa4_9_y0 = f_u_arrmul24_fa4_9_f_u_arrmul24_and4_9_y0 ^ f_u_arrmul24_fa4_9_f_u_arrmul24_fa5_8_y2;
  assign f_u_arrmul24_fa4_9_y1 = f_u_arrmul24_fa4_9_f_u_arrmul24_and4_9_y0 & f_u_arrmul24_fa4_9_f_u_arrmul24_fa5_8_y2;
  assign f_u_arrmul24_fa4_9_y2 = f_u_arrmul24_fa4_9_y0 ^ f_u_arrmul24_fa4_9_f_u_arrmul24_fa3_9_y4;
  assign f_u_arrmul24_fa4_9_y3 = f_u_arrmul24_fa4_9_y0 & f_u_arrmul24_fa4_9_f_u_arrmul24_fa3_9_y4;
  assign f_u_arrmul24_fa4_9_y4 = f_u_arrmul24_fa4_9_y1 | f_u_arrmul24_fa4_9_y3;
  assign f_u_arrmul24_and5_9_a_5 = a_5;
  assign f_u_arrmul24_and5_9_b_9 = b_9;
  assign f_u_arrmul24_and5_9_y0 = f_u_arrmul24_and5_9_a_5 & f_u_arrmul24_and5_9_b_9;
  assign f_u_arrmul24_fa5_9_f_u_arrmul24_and5_9_y0 = f_u_arrmul24_and5_9_y0;
  assign f_u_arrmul24_fa5_9_f_u_arrmul24_fa6_8_y2 = f_u_arrmul24_fa6_8_y2;
  assign f_u_arrmul24_fa5_9_f_u_arrmul24_fa4_9_y4 = f_u_arrmul24_fa4_9_y4;
  assign f_u_arrmul24_fa5_9_y0 = f_u_arrmul24_fa5_9_f_u_arrmul24_and5_9_y0 ^ f_u_arrmul24_fa5_9_f_u_arrmul24_fa6_8_y2;
  assign f_u_arrmul24_fa5_9_y1 = f_u_arrmul24_fa5_9_f_u_arrmul24_and5_9_y0 & f_u_arrmul24_fa5_9_f_u_arrmul24_fa6_8_y2;
  assign f_u_arrmul24_fa5_9_y2 = f_u_arrmul24_fa5_9_y0 ^ f_u_arrmul24_fa5_9_f_u_arrmul24_fa4_9_y4;
  assign f_u_arrmul24_fa5_9_y3 = f_u_arrmul24_fa5_9_y0 & f_u_arrmul24_fa5_9_f_u_arrmul24_fa4_9_y4;
  assign f_u_arrmul24_fa5_9_y4 = f_u_arrmul24_fa5_9_y1 | f_u_arrmul24_fa5_9_y3;
  assign f_u_arrmul24_and6_9_a_6 = a_6;
  assign f_u_arrmul24_and6_9_b_9 = b_9;
  assign f_u_arrmul24_and6_9_y0 = f_u_arrmul24_and6_9_a_6 & f_u_arrmul24_and6_9_b_9;
  assign f_u_arrmul24_fa6_9_f_u_arrmul24_and6_9_y0 = f_u_arrmul24_and6_9_y0;
  assign f_u_arrmul24_fa6_9_f_u_arrmul24_fa7_8_y2 = f_u_arrmul24_fa7_8_y2;
  assign f_u_arrmul24_fa6_9_f_u_arrmul24_fa5_9_y4 = f_u_arrmul24_fa5_9_y4;
  assign f_u_arrmul24_fa6_9_y0 = f_u_arrmul24_fa6_9_f_u_arrmul24_and6_9_y0 ^ f_u_arrmul24_fa6_9_f_u_arrmul24_fa7_8_y2;
  assign f_u_arrmul24_fa6_9_y1 = f_u_arrmul24_fa6_9_f_u_arrmul24_and6_9_y0 & f_u_arrmul24_fa6_9_f_u_arrmul24_fa7_8_y2;
  assign f_u_arrmul24_fa6_9_y2 = f_u_arrmul24_fa6_9_y0 ^ f_u_arrmul24_fa6_9_f_u_arrmul24_fa5_9_y4;
  assign f_u_arrmul24_fa6_9_y3 = f_u_arrmul24_fa6_9_y0 & f_u_arrmul24_fa6_9_f_u_arrmul24_fa5_9_y4;
  assign f_u_arrmul24_fa6_9_y4 = f_u_arrmul24_fa6_9_y1 | f_u_arrmul24_fa6_9_y3;
  assign f_u_arrmul24_and7_9_a_7 = a_7;
  assign f_u_arrmul24_and7_9_b_9 = b_9;
  assign f_u_arrmul24_and7_9_y0 = f_u_arrmul24_and7_9_a_7 & f_u_arrmul24_and7_9_b_9;
  assign f_u_arrmul24_fa7_9_f_u_arrmul24_and7_9_y0 = f_u_arrmul24_and7_9_y0;
  assign f_u_arrmul24_fa7_9_f_u_arrmul24_fa8_8_y2 = f_u_arrmul24_fa8_8_y2;
  assign f_u_arrmul24_fa7_9_f_u_arrmul24_fa6_9_y4 = f_u_arrmul24_fa6_9_y4;
  assign f_u_arrmul24_fa7_9_y0 = f_u_arrmul24_fa7_9_f_u_arrmul24_and7_9_y0 ^ f_u_arrmul24_fa7_9_f_u_arrmul24_fa8_8_y2;
  assign f_u_arrmul24_fa7_9_y1 = f_u_arrmul24_fa7_9_f_u_arrmul24_and7_9_y0 & f_u_arrmul24_fa7_9_f_u_arrmul24_fa8_8_y2;
  assign f_u_arrmul24_fa7_9_y2 = f_u_arrmul24_fa7_9_y0 ^ f_u_arrmul24_fa7_9_f_u_arrmul24_fa6_9_y4;
  assign f_u_arrmul24_fa7_9_y3 = f_u_arrmul24_fa7_9_y0 & f_u_arrmul24_fa7_9_f_u_arrmul24_fa6_9_y4;
  assign f_u_arrmul24_fa7_9_y4 = f_u_arrmul24_fa7_9_y1 | f_u_arrmul24_fa7_9_y3;
  assign f_u_arrmul24_and8_9_a_8 = a_8;
  assign f_u_arrmul24_and8_9_b_9 = b_9;
  assign f_u_arrmul24_and8_9_y0 = f_u_arrmul24_and8_9_a_8 & f_u_arrmul24_and8_9_b_9;
  assign f_u_arrmul24_fa8_9_f_u_arrmul24_and8_9_y0 = f_u_arrmul24_and8_9_y0;
  assign f_u_arrmul24_fa8_9_f_u_arrmul24_fa9_8_y2 = f_u_arrmul24_fa9_8_y2;
  assign f_u_arrmul24_fa8_9_f_u_arrmul24_fa7_9_y4 = f_u_arrmul24_fa7_9_y4;
  assign f_u_arrmul24_fa8_9_y0 = f_u_arrmul24_fa8_9_f_u_arrmul24_and8_9_y0 ^ f_u_arrmul24_fa8_9_f_u_arrmul24_fa9_8_y2;
  assign f_u_arrmul24_fa8_9_y1 = f_u_arrmul24_fa8_9_f_u_arrmul24_and8_9_y0 & f_u_arrmul24_fa8_9_f_u_arrmul24_fa9_8_y2;
  assign f_u_arrmul24_fa8_9_y2 = f_u_arrmul24_fa8_9_y0 ^ f_u_arrmul24_fa8_9_f_u_arrmul24_fa7_9_y4;
  assign f_u_arrmul24_fa8_9_y3 = f_u_arrmul24_fa8_9_y0 & f_u_arrmul24_fa8_9_f_u_arrmul24_fa7_9_y4;
  assign f_u_arrmul24_fa8_9_y4 = f_u_arrmul24_fa8_9_y1 | f_u_arrmul24_fa8_9_y3;
  assign f_u_arrmul24_and9_9_a_9 = a_9;
  assign f_u_arrmul24_and9_9_b_9 = b_9;
  assign f_u_arrmul24_and9_9_y0 = f_u_arrmul24_and9_9_a_9 & f_u_arrmul24_and9_9_b_9;
  assign f_u_arrmul24_fa9_9_f_u_arrmul24_and9_9_y0 = f_u_arrmul24_and9_9_y0;
  assign f_u_arrmul24_fa9_9_f_u_arrmul24_fa10_8_y2 = f_u_arrmul24_fa10_8_y2;
  assign f_u_arrmul24_fa9_9_f_u_arrmul24_fa8_9_y4 = f_u_arrmul24_fa8_9_y4;
  assign f_u_arrmul24_fa9_9_y0 = f_u_arrmul24_fa9_9_f_u_arrmul24_and9_9_y0 ^ f_u_arrmul24_fa9_9_f_u_arrmul24_fa10_8_y2;
  assign f_u_arrmul24_fa9_9_y1 = f_u_arrmul24_fa9_9_f_u_arrmul24_and9_9_y0 & f_u_arrmul24_fa9_9_f_u_arrmul24_fa10_8_y2;
  assign f_u_arrmul24_fa9_9_y2 = f_u_arrmul24_fa9_9_y0 ^ f_u_arrmul24_fa9_9_f_u_arrmul24_fa8_9_y4;
  assign f_u_arrmul24_fa9_9_y3 = f_u_arrmul24_fa9_9_y0 & f_u_arrmul24_fa9_9_f_u_arrmul24_fa8_9_y4;
  assign f_u_arrmul24_fa9_9_y4 = f_u_arrmul24_fa9_9_y1 | f_u_arrmul24_fa9_9_y3;
  assign f_u_arrmul24_and10_9_a_10 = a_10;
  assign f_u_arrmul24_and10_9_b_9 = b_9;
  assign f_u_arrmul24_and10_9_y0 = f_u_arrmul24_and10_9_a_10 & f_u_arrmul24_and10_9_b_9;
  assign f_u_arrmul24_fa10_9_f_u_arrmul24_and10_9_y0 = f_u_arrmul24_and10_9_y0;
  assign f_u_arrmul24_fa10_9_f_u_arrmul24_fa11_8_y2 = f_u_arrmul24_fa11_8_y2;
  assign f_u_arrmul24_fa10_9_f_u_arrmul24_fa9_9_y4 = f_u_arrmul24_fa9_9_y4;
  assign f_u_arrmul24_fa10_9_y0 = f_u_arrmul24_fa10_9_f_u_arrmul24_and10_9_y0 ^ f_u_arrmul24_fa10_9_f_u_arrmul24_fa11_8_y2;
  assign f_u_arrmul24_fa10_9_y1 = f_u_arrmul24_fa10_9_f_u_arrmul24_and10_9_y0 & f_u_arrmul24_fa10_9_f_u_arrmul24_fa11_8_y2;
  assign f_u_arrmul24_fa10_9_y2 = f_u_arrmul24_fa10_9_y0 ^ f_u_arrmul24_fa10_9_f_u_arrmul24_fa9_9_y4;
  assign f_u_arrmul24_fa10_9_y3 = f_u_arrmul24_fa10_9_y0 & f_u_arrmul24_fa10_9_f_u_arrmul24_fa9_9_y4;
  assign f_u_arrmul24_fa10_9_y4 = f_u_arrmul24_fa10_9_y1 | f_u_arrmul24_fa10_9_y3;
  assign f_u_arrmul24_and11_9_a_11 = a_11;
  assign f_u_arrmul24_and11_9_b_9 = b_9;
  assign f_u_arrmul24_and11_9_y0 = f_u_arrmul24_and11_9_a_11 & f_u_arrmul24_and11_9_b_9;
  assign f_u_arrmul24_fa11_9_f_u_arrmul24_and11_9_y0 = f_u_arrmul24_and11_9_y0;
  assign f_u_arrmul24_fa11_9_f_u_arrmul24_fa12_8_y2 = f_u_arrmul24_fa12_8_y2;
  assign f_u_arrmul24_fa11_9_f_u_arrmul24_fa10_9_y4 = f_u_arrmul24_fa10_9_y4;
  assign f_u_arrmul24_fa11_9_y0 = f_u_arrmul24_fa11_9_f_u_arrmul24_and11_9_y0 ^ f_u_arrmul24_fa11_9_f_u_arrmul24_fa12_8_y2;
  assign f_u_arrmul24_fa11_9_y1 = f_u_arrmul24_fa11_9_f_u_arrmul24_and11_9_y0 & f_u_arrmul24_fa11_9_f_u_arrmul24_fa12_8_y2;
  assign f_u_arrmul24_fa11_9_y2 = f_u_arrmul24_fa11_9_y0 ^ f_u_arrmul24_fa11_9_f_u_arrmul24_fa10_9_y4;
  assign f_u_arrmul24_fa11_9_y3 = f_u_arrmul24_fa11_9_y0 & f_u_arrmul24_fa11_9_f_u_arrmul24_fa10_9_y4;
  assign f_u_arrmul24_fa11_9_y4 = f_u_arrmul24_fa11_9_y1 | f_u_arrmul24_fa11_9_y3;
  assign f_u_arrmul24_and12_9_a_12 = a_12;
  assign f_u_arrmul24_and12_9_b_9 = b_9;
  assign f_u_arrmul24_and12_9_y0 = f_u_arrmul24_and12_9_a_12 & f_u_arrmul24_and12_9_b_9;
  assign f_u_arrmul24_fa12_9_f_u_arrmul24_and12_9_y0 = f_u_arrmul24_and12_9_y0;
  assign f_u_arrmul24_fa12_9_f_u_arrmul24_fa13_8_y2 = f_u_arrmul24_fa13_8_y2;
  assign f_u_arrmul24_fa12_9_f_u_arrmul24_fa11_9_y4 = f_u_arrmul24_fa11_9_y4;
  assign f_u_arrmul24_fa12_9_y0 = f_u_arrmul24_fa12_9_f_u_arrmul24_and12_9_y0 ^ f_u_arrmul24_fa12_9_f_u_arrmul24_fa13_8_y2;
  assign f_u_arrmul24_fa12_9_y1 = f_u_arrmul24_fa12_9_f_u_arrmul24_and12_9_y0 & f_u_arrmul24_fa12_9_f_u_arrmul24_fa13_8_y2;
  assign f_u_arrmul24_fa12_9_y2 = f_u_arrmul24_fa12_9_y0 ^ f_u_arrmul24_fa12_9_f_u_arrmul24_fa11_9_y4;
  assign f_u_arrmul24_fa12_9_y3 = f_u_arrmul24_fa12_9_y0 & f_u_arrmul24_fa12_9_f_u_arrmul24_fa11_9_y4;
  assign f_u_arrmul24_fa12_9_y4 = f_u_arrmul24_fa12_9_y1 | f_u_arrmul24_fa12_9_y3;
  assign f_u_arrmul24_and13_9_a_13 = a_13;
  assign f_u_arrmul24_and13_9_b_9 = b_9;
  assign f_u_arrmul24_and13_9_y0 = f_u_arrmul24_and13_9_a_13 & f_u_arrmul24_and13_9_b_9;
  assign f_u_arrmul24_fa13_9_f_u_arrmul24_and13_9_y0 = f_u_arrmul24_and13_9_y0;
  assign f_u_arrmul24_fa13_9_f_u_arrmul24_fa14_8_y2 = f_u_arrmul24_fa14_8_y2;
  assign f_u_arrmul24_fa13_9_f_u_arrmul24_fa12_9_y4 = f_u_arrmul24_fa12_9_y4;
  assign f_u_arrmul24_fa13_9_y0 = f_u_arrmul24_fa13_9_f_u_arrmul24_and13_9_y0 ^ f_u_arrmul24_fa13_9_f_u_arrmul24_fa14_8_y2;
  assign f_u_arrmul24_fa13_9_y1 = f_u_arrmul24_fa13_9_f_u_arrmul24_and13_9_y0 & f_u_arrmul24_fa13_9_f_u_arrmul24_fa14_8_y2;
  assign f_u_arrmul24_fa13_9_y2 = f_u_arrmul24_fa13_9_y0 ^ f_u_arrmul24_fa13_9_f_u_arrmul24_fa12_9_y4;
  assign f_u_arrmul24_fa13_9_y3 = f_u_arrmul24_fa13_9_y0 & f_u_arrmul24_fa13_9_f_u_arrmul24_fa12_9_y4;
  assign f_u_arrmul24_fa13_9_y4 = f_u_arrmul24_fa13_9_y1 | f_u_arrmul24_fa13_9_y3;
  assign f_u_arrmul24_and14_9_a_14 = a_14;
  assign f_u_arrmul24_and14_9_b_9 = b_9;
  assign f_u_arrmul24_and14_9_y0 = f_u_arrmul24_and14_9_a_14 & f_u_arrmul24_and14_9_b_9;
  assign f_u_arrmul24_fa14_9_f_u_arrmul24_and14_9_y0 = f_u_arrmul24_and14_9_y0;
  assign f_u_arrmul24_fa14_9_f_u_arrmul24_fa15_8_y2 = f_u_arrmul24_fa15_8_y2;
  assign f_u_arrmul24_fa14_9_f_u_arrmul24_fa13_9_y4 = f_u_arrmul24_fa13_9_y4;
  assign f_u_arrmul24_fa14_9_y0 = f_u_arrmul24_fa14_9_f_u_arrmul24_and14_9_y0 ^ f_u_arrmul24_fa14_9_f_u_arrmul24_fa15_8_y2;
  assign f_u_arrmul24_fa14_9_y1 = f_u_arrmul24_fa14_9_f_u_arrmul24_and14_9_y0 & f_u_arrmul24_fa14_9_f_u_arrmul24_fa15_8_y2;
  assign f_u_arrmul24_fa14_9_y2 = f_u_arrmul24_fa14_9_y0 ^ f_u_arrmul24_fa14_9_f_u_arrmul24_fa13_9_y4;
  assign f_u_arrmul24_fa14_9_y3 = f_u_arrmul24_fa14_9_y0 & f_u_arrmul24_fa14_9_f_u_arrmul24_fa13_9_y4;
  assign f_u_arrmul24_fa14_9_y4 = f_u_arrmul24_fa14_9_y1 | f_u_arrmul24_fa14_9_y3;
  assign f_u_arrmul24_and15_9_a_15 = a_15;
  assign f_u_arrmul24_and15_9_b_9 = b_9;
  assign f_u_arrmul24_and15_9_y0 = f_u_arrmul24_and15_9_a_15 & f_u_arrmul24_and15_9_b_9;
  assign f_u_arrmul24_fa15_9_f_u_arrmul24_and15_9_y0 = f_u_arrmul24_and15_9_y0;
  assign f_u_arrmul24_fa15_9_f_u_arrmul24_fa16_8_y2 = f_u_arrmul24_fa16_8_y2;
  assign f_u_arrmul24_fa15_9_f_u_arrmul24_fa14_9_y4 = f_u_arrmul24_fa14_9_y4;
  assign f_u_arrmul24_fa15_9_y0 = f_u_arrmul24_fa15_9_f_u_arrmul24_and15_9_y0 ^ f_u_arrmul24_fa15_9_f_u_arrmul24_fa16_8_y2;
  assign f_u_arrmul24_fa15_9_y1 = f_u_arrmul24_fa15_9_f_u_arrmul24_and15_9_y0 & f_u_arrmul24_fa15_9_f_u_arrmul24_fa16_8_y2;
  assign f_u_arrmul24_fa15_9_y2 = f_u_arrmul24_fa15_9_y0 ^ f_u_arrmul24_fa15_9_f_u_arrmul24_fa14_9_y4;
  assign f_u_arrmul24_fa15_9_y3 = f_u_arrmul24_fa15_9_y0 & f_u_arrmul24_fa15_9_f_u_arrmul24_fa14_9_y4;
  assign f_u_arrmul24_fa15_9_y4 = f_u_arrmul24_fa15_9_y1 | f_u_arrmul24_fa15_9_y3;
  assign f_u_arrmul24_and16_9_a_16 = a_16;
  assign f_u_arrmul24_and16_9_b_9 = b_9;
  assign f_u_arrmul24_and16_9_y0 = f_u_arrmul24_and16_9_a_16 & f_u_arrmul24_and16_9_b_9;
  assign f_u_arrmul24_fa16_9_f_u_arrmul24_and16_9_y0 = f_u_arrmul24_and16_9_y0;
  assign f_u_arrmul24_fa16_9_f_u_arrmul24_fa17_8_y2 = f_u_arrmul24_fa17_8_y2;
  assign f_u_arrmul24_fa16_9_f_u_arrmul24_fa15_9_y4 = f_u_arrmul24_fa15_9_y4;
  assign f_u_arrmul24_fa16_9_y0 = f_u_arrmul24_fa16_9_f_u_arrmul24_and16_9_y0 ^ f_u_arrmul24_fa16_9_f_u_arrmul24_fa17_8_y2;
  assign f_u_arrmul24_fa16_9_y1 = f_u_arrmul24_fa16_9_f_u_arrmul24_and16_9_y0 & f_u_arrmul24_fa16_9_f_u_arrmul24_fa17_8_y2;
  assign f_u_arrmul24_fa16_9_y2 = f_u_arrmul24_fa16_9_y0 ^ f_u_arrmul24_fa16_9_f_u_arrmul24_fa15_9_y4;
  assign f_u_arrmul24_fa16_9_y3 = f_u_arrmul24_fa16_9_y0 & f_u_arrmul24_fa16_9_f_u_arrmul24_fa15_9_y4;
  assign f_u_arrmul24_fa16_9_y4 = f_u_arrmul24_fa16_9_y1 | f_u_arrmul24_fa16_9_y3;
  assign f_u_arrmul24_and17_9_a_17 = a_17;
  assign f_u_arrmul24_and17_9_b_9 = b_9;
  assign f_u_arrmul24_and17_9_y0 = f_u_arrmul24_and17_9_a_17 & f_u_arrmul24_and17_9_b_9;
  assign f_u_arrmul24_fa17_9_f_u_arrmul24_and17_9_y0 = f_u_arrmul24_and17_9_y0;
  assign f_u_arrmul24_fa17_9_f_u_arrmul24_fa18_8_y2 = f_u_arrmul24_fa18_8_y2;
  assign f_u_arrmul24_fa17_9_f_u_arrmul24_fa16_9_y4 = f_u_arrmul24_fa16_9_y4;
  assign f_u_arrmul24_fa17_9_y0 = f_u_arrmul24_fa17_9_f_u_arrmul24_and17_9_y0 ^ f_u_arrmul24_fa17_9_f_u_arrmul24_fa18_8_y2;
  assign f_u_arrmul24_fa17_9_y1 = f_u_arrmul24_fa17_9_f_u_arrmul24_and17_9_y0 & f_u_arrmul24_fa17_9_f_u_arrmul24_fa18_8_y2;
  assign f_u_arrmul24_fa17_9_y2 = f_u_arrmul24_fa17_9_y0 ^ f_u_arrmul24_fa17_9_f_u_arrmul24_fa16_9_y4;
  assign f_u_arrmul24_fa17_9_y3 = f_u_arrmul24_fa17_9_y0 & f_u_arrmul24_fa17_9_f_u_arrmul24_fa16_9_y4;
  assign f_u_arrmul24_fa17_9_y4 = f_u_arrmul24_fa17_9_y1 | f_u_arrmul24_fa17_9_y3;
  assign f_u_arrmul24_and18_9_a_18 = a_18;
  assign f_u_arrmul24_and18_9_b_9 = b_9;
  assign f_u_arrmul24_and18_9_y0 = f_u_arrmul24_and18_9_a_18 & f_u_arrmul24_and18_9_b_9;
  assign f_u_arrmul24_fa18_9_f_u_arrmul24_and18_9_y0 = f_u_arrmul24_and18_9_y0;
  assign f_u_arrmul24_fa18_9_f_u_arrmul24_fa19_8_y2 = f_u_arrmul24_fa19_8_y2;
  assign f_u_arrmul24_fa18_9_f_u_arrmul24_fa17_9_y4 = f_u_arrmul24_fa17_9_y4;
  assign f_u_arrmul24_fa18_9_y0 = f_u_arrmul24_fa18_9_f_u_arrmul24_and18_9_y0 ^ f_u_arrmul24_fa18_9_f_u_arrmul24_fa19_8_y2;
  assign f_u_arrmul24_fa18_9_y1 = f_u_arrmul24_fa18_9_f_u_arrmul24_and18_9_y0 & f_u_arrmul24_fa18_9_f_u_arrmul24_fa19_8_y2;
  assign f_u_arrmul24_fa18_9_y2 = f_u_arrmul24_fa18_9_y0 ^ f_u_arrmul24_fa18_9_f_u_arrmul24_fa17_9_y4;
  assign f_u_arrmul24_fa18_9_y3 = f_u_arrmul24_fa18_9_y0 & f_u_arrmul24_fa18_9_f_u_arrmul24_fa17_9_y4;
  assign f_u_arrmul24_fa18_9_y4 = f_u_arrmul24_fa18_9_y1 | f_u_arrmul24_fa18_9_y3;
  assign f_u_arrmul24_and19_9_a_19 = a_19;
  assign f_u_arrmul24_and19_9_b_9 = b_9;
  assign f_u_arrmul24_and19_9_y0 = f_u_arrmul24_and19_9_a_19 & f_u_arrmul24_and19_9_b_9;
  assign f_u_arrmul24_fa19_9_f_u_arrmul24_and19_9_y0 = f_u_arrmul24_and19_9_y0;
  assign f_u_arrmul24_fa19_9_f_u_arrmul24_fa20_8_y2 = f_u_arrmul24_fa20_8_y2;
  assign f_u_arrmul24_fa19_9_f_u_arrmul24_fa18_9_y4 = f_u_arrmul24_fa18_9_y4;
  assign f_u_arrmul24_fa19_9_y0 = f_u_arrmul24_fa19_9_f_u_arrmul24_and19_9_y0 ^ f_u_arrmul24_fa19_9_f_u_arrmul24_fa20_8_y2;
  assign f_u_arrmul24_fa19_9_y1 = f_u_arrmul24_fa19_9_f_u_arrmul24_and19_9_y0 & f_u_arrmul24_fa19_9_f_u_arrmul24_fa20_8_y2;
  assign f_u_arrmul24_fa19_9_y2 = f_u_arrmul24_fa19_9_y0 ^ f_u_arrmul24_fa19_9_f_u_arrmul24_fa18_9_y4;
  assign f_u_arrmul24_fa19_9_y3 = f_u_arrmul24_fa19_9_y0 & f_u_arrmul24_fa19_9_f_u_arrmul24_fa18_9_y4;
  assign f_u_arrmul24_fa19_9_y4 = f_u_arrmul24_fa19_9_y1 | f_u_arrmul24_fa19_9_y3;
  assign f_u_arrmul24_and20_9_a_20 = a_20;
  assign f_u_arrmul24_and20_9_b_9 = b_9;
  assign f_u_arrmul24_and20_9_y0 = f_u_arrmul24_and20_9_a_20 & f_u_arrmul24_and20_9_b_9;
  assign f_u_arrmul24_fa20_9_f_u_arrmul24_and20_9_y0 = f_u_arrmul24_and20_9_y0;
  assign f_u_arrmul24_fa20_9_f_u_arrmul24_fa21_8_y2 = f_u_arrmul24_fa21_8_y2;
  assign f_u_arrmul24_fa20_9_f_u_arrmul24_fa19_9_y4 = f_u_arrmul24_fa19_9_y4;
  assign f_u_arrmul24_fa20_9_y0 = f_u_arrmul24_fa20_9_f_u_arrmul24_and20_9_y0 ^ f_u_arrmul24_fa20_9_f_u_arrmul24_fa21_8_y2;
  assign f_u_arrmul24_fa20_9_y1 = f_u_arrmul24_fa20_9_f_u_arrmul24_and20_9_y0 & f_u_arrmul24_fa20_9_f_u_arrmul24_fa21_8_y2;
  assign f_u_arrmul24_fa20_9_y2 = f_u_arrmul24_fa20_9_y0 ^ f_u_arrmul24_fa20_9_f_u_arrmul24_fa19_9_y4;
  assign f_u_arrmul24_fa20_9_y3 = f_u_arrmul24_fa20_9_y0 & f_u_arrmul24_fa20_9_f_u_arrmul24_fa19_9_y4;
  assign f_u_arrmul24_fa20_9_y4 = f_u_arrmul24_fa20_9_y1 | f_u_arrmul24_fa20_9_y3;
  assign f_u_arrmul24_and21_9_a_21 = a_21;
  assign f_u_arrmul24_and21_9_b_9 = b_9;
  assign f_u_arrmul24_and21_9_y0 = f_u_arrmul24_and21_9_a_21 & f_u_arrmul24_and21_9_b_9;
  assign f_u_arrmul24_fa21_9_f_u_arrmul24_and21_9_y0 = f_u_arrmul24_and21_9_y0;
  assign f_u_arrmul24_fa21_9_f_u_arrmul24_fa22_8_y2 = f_u_arrmul24_fa22_8_y2;
  assign f_u_arrmul24_fa21_9_f_u_arrmul24_fa20_9_y4 = f_u_arrmul24_fa20_9_y4;
  assign f_u_arrmul24_fa21_9_y0 = f_u_arrmul24_fa21_9_f_u_arrmul24_and21_9_y0 ^ f_u_arrmul24_fa21_9_f_u_arrmul24_fa22_8_y2;
  assign f_u_arrmul24_fa21_9_y1 = f_u_arrmul24_fa21_9_f_u_arrmul24_and21_9_y0 & f_u_arrmul24_fa21_9_f_u_arrmul24_fa22_8_y2;
  assign f_u_arrmul24_fa21_9_y2 = f_u_arrmul24_fa21_9_y0 ^ f_u_arrmul24_fa21_9_f_u_arrmul24_fa20_9_y4;
  assign f_u_arrmul24_fa21_9_y3 = f_u_arrmul24_fa21_9_y0 & f_u_arrmul24_fa21_9_f_u_arrmul24_fa20_9_y4;
  assign f_u_arrmul24_fa21_9_y4 = f_u_arrmul24_fa21_9_y1 | f_u_arrmul24_fa21_9_y3;
  assign f_u_arrmul24_and22_9_a_22 = a_22;
  assign f_u_arrmul24_and22_9_b_9 = b_9;
  assign f_u_arrmul24_and22_9_y0 = f_u_arrmul24_and22_9_a_22 & f_u_arrmul24_and22_9_b_9;
  assign f_u_arrmul24_fa22_9_f_u_arrmul24_and22_9_y0 = f_u_arrmul24_and22_9_y0;
  assign f_u_arrmul24_fa22_9_f_u_arrmul24_fa23_8_y2 = f_u_arrmul24_fa23_8_y2;
  assign f_u_arrmul24_fa22_9_f_u_arrmul24_fa21_9_y4 = f_u_arrmul24_fa21_9_y4;
  assign f_u_arrmul24_fa22_9_y0 = f_u_arrmul24_fa22_9_f_u_arrmul24_and22_9_y0 ^ f_u_arrmul24_fa22_9_f_u_arrmul24_fa23_8_y2;
  assign f_u_arrmul24_fa22_9_y1 = f_u_arrmul24_fa22_9_f_u_arrmul24_and22_9_y0 & f_u_arrmul24_fa22_9_f_u_arrmul24_fa23_8_y2;
  assign f_u_arrmul24_fa22_9_y2 = f_u_arrmul24_fa22_9_y0 ^ f_u_arrmul24_fa22_9_f_u_arrmul24_fa21_9_y4;
  assign f_u_arrmul24_fa22_9_y3 = f_u_arrmul24_fa22_9_y0 & f_u_arrmul24_fa22_9_f_u_arrmul24_fa21_9_y4;
  assign f_u_arrmul24_fa22_9_y4 = f_u_arrmul24_fa22_9_y1 | f_u_arrmul24_fa22_9_y3;
  assign f_u_arrmul24_and23_9_a_23 = a_23;
  assign f_u_arrmul24_and23_9_b_9 = b_9;
  assign f_u_arrmul24_and23_9_y0 = f_u_arrmul24_and23_9_a_23 & f_u_arrmul24_and23_9_b_9;
  assign f_u_arrmul24_fa23_9_f_u_arrmul24_and23_9_y0 = f_u_arrmul24_and23_9_y0;
  assign f_u_arrmul24_fa23_9_f_u_arrmul24_fa23_8_y4 = f_u_arrmul24_fa23_8_y4;
  assign f_u_arrmul24_fa23_9_f_u_arrmul24_fa22_9_y4 = f_u_arrmul24_fa22_9_y4;
  assign f_u_arrmul24_fa23_9_y0 = f_u_arrmul24_fa23_9_f_u_arrmul24_and23_9_y0 ^ f_u_arrmul24_fa23_9_f_u_arrmul24_fa23_8_y4;
  assign f_u_arrmul24_fa23_9_y1 = f_u_arrmul24_fa23_9_f_u_arrmul24_and23_9_y0 & f_u_arrmul24_fa23_9_f_u_arrmul24_fa23_8_y4;
  assign f_u_arrmul24_fa23_9_y2 = f_u_arrmul24_fa23_9_y0 ^ f_u_arrmul24_fa23_9_f_u_arrmul24_fa22_9_y4;
  assign f_u_arrmul24_fa23_9_y3 = f_u_arrmul24_fa23_9_y0 & f_u_arrmul24_fa23_9_f_u_arrmul24_fa22_9_y4;
  assign f_u_arrmul24_fa23_9_y4 = f_u_arrmul24_fa23_9_y1 | f_u_arrmul24_fa23_9_y3;
  assign f_u_arrmul24_and0_10_a_0 = a_0;
  assign f_u_arrmul24_and0_10_b_10 = b_10;
  assign f_u_arrmul24_and0_10_y0 = f_u_arrmul24_and0_10_a_0 & f_u_arrmul24_and0_10_b_10;
  assign f_u_arrmul24_ha0_10_f_u_arrmul24_and0_10_y0 = f_u_arrmul24_and0_10_y0;
  assign f_u_arrmul24_ha0_10_f_u_arrmul24_fa1_9_y2 = f_u_arrmul24_fa1_9_y2;
  assign f_u_arrmul24_ha0_10_y0 = f_u_arrmul24_ha0_10_f_u_arrmul24_and0_10_y0 ^ f_u_arrmul24_ha0_10_f_u_arrmul24_fa1_9_y2;
  assign f_u_arrmul24_ha0_10_y1 = f_u_arrmul24_ha0_10_f_u_arrmul24_and0_10_y0 & f_u_arrmul24_ha0_10_f_u_arrmul24_fa1_9_y2;
  assign f_u_arrmul24_and1_10_a_1 = a_1;
  assign f_u_arrmul24_and1_10_b_10 = b_10;
  assign f_u_arrmul24_and1_10_y0 = f_u_arrmul24_and1_10_a_1 & f_u_arrmul24_and1_10_b_10;
  assign f_u_arrmul24_fa1_10_f_u_arrmul24_and1_10_y0 = f_u_arrmul24_and1_10_y0;
  assign f_u_arrmul24_fa1_10_f_u_arrmul24_fa2_9_y2 = f_u_arrmul24_fa2_9_y2;
  assign f_u_arrmul24_fa1_10_f_u_arrmul24_ha0_10_y1 = f_u_arrmul24_ha0_10_y1;
  assign f_u_arrmul24_fa1_10_y0 = f_u_arrmul24_fa1_10_f_u_arrmul24_and1_10_y0 ^ f_u_arrmul24_fa1_10_f_u_arrmul24_fa2_9_y2;
  assign f_u_arrmul24_fa1_10_y1 = f_u_arrmul24_fa1_10_f_u_arrmul24_and1_10_y0 & f_u_arrmul24_fa1_10_f_u_arrmul24_fa2_9_y2;
  assign f_u_arrmul24_fa1_10_y2 = f_u_arrmul24_fa1_10_y0 ^ f_u_arrmul24_fa1_10_f_u_arrmul24_ha0_10_y1;
  assign f_u_arrmul24_fa1_10_y3 = f_u_arrmul24_fa1_10_y0 & f_u_arrmul24_fa1_10_f_u_arrmul24_ha0_10_y1;
  assign f_u_arrmul24_fa1_10_y4 = f_u_arrmul24_fa1_10_y1 | f_u_arrmul24_fa1_10_y3;
  assign f_u_arrmul24_and2_10_a_2 = a_2;
  assign f_u_arrmul24_and2_10_b_10 = b_10;
  assign f_u_arrmul24_and2_10_y0 = f_u_arrmul24_and2_10_a_2 & f_u_arrmul24_and2_10_b_10;
  assign f_u_arrmul24_fa2_10_f_u_arrmul24_and2_10_y0 = f_u_arrmul24_and2_10_y0;
  assign f_u_arrmul24_fa2_10_f_u_arrmul24_fa3_9_y2 = f_u_arrmul24_fa3_9_y2;
  assign f_u_arrmul24_fa2_10_f_u_arrmul24_fa1_10_y4 = f_u_arrmul24_fa1_10_y4;
  assign f_u_arrmul24_fa2_10_y0 = f_u_arrmul24_fa2_10_f_u_arrmul24_and2_10_y0 ^ f_u_arrmul24_fa2_10_f_u_arrmul24_fa3_9_y2;
  assign f_u_arrmul24_fa2_10_y1 = f_u_arrmul24_fa2_10_f_u_arrmul24_and2_10_y0 & f_u_arrmul24_fa2_10_f_u_arrmul24_fa3_9_y2;
  assign f_u_arrmul24_fa2_10_y2 = f_u_arrmul24_fa2_10_y0 ^ f_u_arrmul24_fa2_10_f_u_arrmul24_fa1_10_y4;
  assign f_u_arrmul24_fa2_10_y3 = f_u_arrmul24_fa2_10_y0 & f_u_arrmul24_fa2_10_f_u_arrmul24_fa1_10_y4;
  assign f_u_arrmul24_fa2_10_y4 = f_u_arrmul24_fa2_10_y1 | f_u_arrmul24_fa2_10_y3;
  assign f_u_arrmul24_and3_10_a_3 = a_3;
  assign f_u_arrmul24_and3_10_b_10 = b_10;
  assign f_u_arrmul24_and3_10_y0 = f_u_arrmul24_and3_10_a_3 & f_u_arrmul24_and3_10_b_10;
  assign f_u_arrmul24_fa3_10_f_u_arrmul24_and3_10_y0 = f_u_arrmul24_and3_10_y0;
  assign f_u_arrmul24_fa3_10_f_u_arrmul24_fa4_9_y2 = f_u_arrmul24_fa4_9_y2;
  assign f_u_arrmul24_fa3_10_f_u_arrmul24_fa2_10_y4 = f_u_arrmul24_fa2_10_y4;
  assign f_u_arrmul24_fa3_10_y0 = f_u_arrmul24_fa3_10_f_u_arrmul24_and3_10_y0 ^ f_u_arrmul24_fa3_10_f_u_arrmul24_fa4_9_y2;
  assign f_u_arrmul24_fa3_10_y1 = f_u_arrmul24_fa3_10_f_u_arrmul24_and3_10_y0 & f_u_arrmul24_fa3_10_f_u_arrmul24_fa4_9_y2;
  assign f_u_arrmul24_fa3_10_y2 = f_u_arrmul24_fa3_10_y0 ^ f_u_arrmul24_fa3_10_f_u_arrmul24_fa2_10_y4;
  assign f_u_arrmul24_fa3_10_y3 = f_u_arrmul24_fa3_10_y0 & f_u_arrmul24_fa3_10_f_u_arrmul24_fa2_10_y4;
  assign f_u_arrmul24_fa3_10_y4 = f_u_arrmul24_fa3_10_y1 | f_u_arrmul24_fa3_10_y3;
  assign f_u_arrmul24_and4_10_a_4 = a_4;
  assign f_u_arrmul24_and4_10_b_10 = b_10;
  assign f_u_arrmul24_and4_10_y0 = f_u_arrmul24_and4_10_a_4 & f_u_arrmul24_and4_10_b_10;
  assign f_u_arrmul24_fa4_10_f_u_arrmul24_and4_10_y0 = f_u_arrmul24_and4_10_y0;
  assign f_u_arrmul24_fa4_10_f_u_arrmul24_fa5_9_y2 = f_u_arrmul24_fa5_9_y2;
  assign f_u_arrmul24_fa4_10_f_u_arrmul24_fa3_10_y4 = f_u_arrmul24_fa3_10_y4;
  assign f_u_arrmul24_fa4_10_y0 = f_u_arrmul24_fa4_10_f_u_arrmul24_and4_10_y0 ^ f_u_arrmul24_fa4_10_f_u_arrmul24_fa5_9_y2;
  assign f_u_arrmul24_fa4_10_y1 = f_u_arrmul24_fa4_10_f_u_arrmul24_and4_10_y0 & f_u_arrmul24_fa4_10_f_u_arrmul24_fa5_9_y2;
  assign f_u_arrmul24_fa4_10_y2 = f_u_arrmul24_fa4_10_y0 ^ f_u_arrmul24_fa4_10_f_u_arrmul24_fa3_10_y4;
  assign f_u_arrmul24_fa4_10_y3 = f_u_arrmul24_fa4_10_y0 & f_u_arrmul24_fa4_10_f_u_arrmul24_fa3_10_y4;
  assign f_u_arrmul24_fa4_10_y4 = f_u_arrmul24_fa4_10_y1 | f_u_arrmul24_fa4_10_y3;
  assign f_u_arrmul24_and5_10_a_5 = a_5;
  assign f_u_arrmul24_and5_10_b_10 = b_10;
  assign f_u_arrmul24_and5_10_y0 = f_u_arrmul24_and5_10_a_5 & f_u_arrmul24_and5_10_b_10;
  assign f_u_arrmul24_fa5_10_f_u_arrmul24_and5_10_y0 = f_u_arrmul24_and5_10_y0;
  assign f_u_arrmul24_fa5_10_f_u_arrmul24_fa6_9_y2 = f_u_arrmul24_fa6_9_y2;
  assign f_u_arrmul24_fa5_10_f_u_arrmul24_fa4_10_y4 = f_u_arrmul24_fa4_10_y4;
  assign f_u_arrmul24_fa5_10_y0 = f_u_arrmul24_fa5_10_f_u_arrmul24_and5_10_y0 ^ f_u_arrmul24_fa5_10_f_u_arrmul24_fa6_9_y2;
  assign f_u_arrmul24_fa5_10_y1 = f_u_arrmul24_fa5_10_f_u_arrmul24_and5_10_y0 & f_u_arrmul24_fa5_10_f_u_arrmul24_fa6_9_y2;
  assign f_u_arrmul24_fa5_10_y2 = f_u_arrmul24_fa5_10_y0 ^ f_u_arrmul24_fa5_10_f_u_arrmul24_fa4_10_y4;
  assign f_u_arrmul24_fa5_10_y3 = f_u_arrmul24_fa5_10_y0 & f_u_arrmul24_fa5_10_f_u_arrmul24_fa4_10_y4;
  assign f_u_arrmul24_fa5_10_y4 = f_u_arrmul24_fa5_10_y1 | f_u_arrmul24_fa5_10_y3;
  assign f_u_arrmul24_and6_10_a_6 = a_6;
  assign f_u_arrmul24_and6_10_b_10 = b_10;
  assign f_u_arrmul24_and6_10_y0 = f_u_arrmul24_and6_10_a_6 & f_u_arrmul24_and6_10_b_10;
  assign f_u_arrmul24_fa6_10_f_u_arrmul24_and6_10_y0 = f_u_arrmul24_and6_10_y0;
  assign f_u_arrmul24_fa6_10_f_u_arrmul24_fa7_9_y2 = f_u_arrmul24_fa7_9_y2;
  assign f_u_arrmul24_fa6_10_f_u_arrmul24_fa5_10_y4 = f_u_arrmul24_fa5_10_y4;
  assign f_u_arrmul24_fa6_10_y0 = f_u_arrmul24_fa6_10_f_u_arrmul24_and6_10_y0 ^ f_u_arrmul24_fa6_10_f_u_arrmul24_fa7_9_y2;
  assign f_u_arrmul24_fa6_10_y1 = f_u_arrmul24_fa6_10_f_u_arrmul24_and6_10_y0 & f_u_arrmul24_fa6_10_f_u_arrmul24_fa7_9_y2;
  assign f_u_arrmul24_fa6_10_y2 = f_u_arrmul24_fa6_10_y0 ^ f_u_arrmul24_fa6_10_f_u_arrmul24_fa5_10_y4;
  assign f_u_arrmul24_fa6_10_y3 = f_u_arrmul24_fa6_10_y0 & f_u_arrmul24_fa6_10_f_u_arrmul24_fa5_10_y4;
  assign f_u_arrmul24_fa6_10_y4 = f_u_arrmul24_fa6_10_y1 | f_u_arrmul24_fa6_10_y3;
  assign f_u_arrmul24_and7_10_a_7 = a_7;
  assign f_u_arrmul24_and7_10_b_10 = b_10;
  assign f_u_arrmul24_and7_10_y0 = f_u_arrmul24_and7_10_a_7 & f_u_arrmul24_and7_10_b_10;
  assign f_u_arrmul24_fa7_10_f_u_arrmul24_and7_10_y0 = f_u_arrmul24_and7_10_y0;
  assign f_u_arrmul24_fa7_10_f_u_arrmul24_fa8_9_y2 = f_u_arrmul24_fa8_9_y2;
  assign f_u_arrmul24_fa7_10_f_u_arrmul24_fa6_10_y4 = f_u_arrmul24_fa6_10_y4;
  assign f_u_arrmul24_fa7_10_y0 = f_u_arrmul24_fa7_10_f_u_arrmul24_and7_10_y0 ^ f_u_arrmul24_fa7_10_f_u_arrmul24_fa8_9_y2;
  assign f_u_arrmul24_fa7_10_y1 = f_u_arrmul24_fa7_10_f_u_arrmul24_and7_10_y0 & f_u_arrmul24_fa7_10_f_u_arrmul24_fa8_9_y2;
  assign f_u_arrmul24_fa7_10_y2 = f_u_arrmul24_fa7_10_y0 ^ f_u_arrmul24_fa7_10_f_u_arrmul24_fa6_10_y4;
  assign f_u_arrmul24_fa7_10_y3 = f_u_arrmul24_fa7_10_y0 & f_u_arrmul24_fa7_10_f_u_arrmul24_fa6_10_y4;
  assign f_u_arrmul24_fa7_10_y4 = f_u_arrmul24_fa7_10_y1 | f_u_arrmul24_fa7_10_y3;
  assign f_u_arrmul24_and8_10_a_8 = a_8;
  assign f_u_arrmul24_and8_10_b_10 = b_10;
  assign f_u_arrmul24_and8_10_y0 = f_u_arrmul24_and8_10_a_8 & f_u_arrmul24_and8_10_b_10;
  assign f_u_arrmul24_fa8_10_f_u_arrmul24_and8_10_y0 = f_u_arrmul24_and8_10_y0;
  assign f_u_arrmul24_fa8_10_f_u_arrmul24_fa9_9_y2 = f_u_arrmul24_fa9_9_y2;
  assign f_u_arrmul24_fa8_10_f_u_arrmul24_fa7_10_y4 = f_u_arrmul24_fa7_10_y4;
  assign f_u_arrmul24_fa8_10_y0 = f_u_arrmul24_fa8_10_f_u_arrmul24_and8_10_y0 ^ f_u_arrmul24_fa8_10_f_u_arrmul24_fa9_9_y2;
  assign f_u_arrmul24_fa8_10_y1 = f_u_arrmul24_fa8_10_f_u_arrmul24_and8_10_y0 & f_u_arrmul24_fa8_10_f_u_arrmul24_fa9_9_y2;
  assign f_u_arrmul24_fa8_10_y2 = f_u_arrmul24_fa8_10_y0 ^ f_u_arrmul24_fa8_10_f_u_arrmul24_fa7_10_y4;
  assign f_u_arrmul24_fa8_10_y3 = f_u_arrmul24_fa8_10_y0 & f_u_arrmul24_fa8_10_f_u_arrmul24_fa7_10_y4;
  assign f_u_arrmul24_fa8_10_y4 = f_u_arrmul24_fa8_10_y1 | f_u_arrmul24_fa8_10_y3;
  assign f_u_arrmul24_and9_10_a_9 = a_9;
  assign f_u_arrmul24_and9_10_b_10 = b_10;
  assign f_u_arrmul24_and9_10_y0 = f_u_arrmul24_and9_10_a_9 & f_u_arrmul24_and9_10_b_10;
  assign f_u_arrmul24_fa9_10_f_u_arrmul24_and9_10_y0 = f_u_arrmul24_and9_10_y0;
  assign f_u_arrmul24_fa9_10_f_u_arrmul24_fa10_9_y2 = f_u_arrmul24_fa10_9_y2;
  assign f_u_arrmul24_fa9_10_f_u_arrmul24_fa8_10_y4 = f_u_arrmul24_fa8_10_y4;
  assign f_u_arrmul24_fa9_10_y0 = f_u_arrmul24_fa9_10_f_u_arrmul24_and9_10_y0 ^ f_u_arrmul24_fa9_10_f_u_arrmul24_fa10_9_y2;
  assign f_u_arrmul24_fa9_10_y1 = f_u_arrmul24_fa9_10_f_u_arrmul24_and9_10_y0 & f_u_arrmul24_fa9_10_f_u_arrmul24_fa10_9_y2;
  assign f_u_arrmul24_fa9_10_y2 = f_u_arrmul24_fa9_10_y0 ^ f_u_arrmul24_fa9_10_f_u_arrmul24_fa8_10_y4;
  assign f_u_arrmul24_fa9_10_y3 = f_u_arrmul24_fa9_10_y0 & f_u_arrmul24_fa9_10_f_u_arrmul24_fa8_10_y4;
  assign f_u_arrmul24_fa9_10_y4 = f_u_arrmul24_fa9_10_y1 | f_u_arrmul24_fa9_10_y3;
  assign f_u_arrmul24_and10_10_a_10 = a_10;
  assign f_u_arrmul24_and10_10_b_10 = b_10;
  assign f_u_arrmul24_and10_10_y0 = f_u_arrmul24_and10_10_a_10 & f_u_arrmul24_and10_10_b_10;
  assign f_u_arrmul24_fa10_10_f_u_arrmul24_and10_10_y0 = f_u_arrmul24_and10_10_y0;
  assign f_u_arrmul24_fa10_10_f_u_arrmul24_fa11_9_y2 = f_u_arrmul24_fa11_9_y2;
  assign f_u_arrmul24_fa10_10_f_u_arrmul24_fa9_10_y4 = f_u_arrmul24_fa9_10_y4;
  assign f_u_arrmul24_fa10_10_y0 = f_u_arrmul24_fa10_10_f_u_arrmul24_and10_10_y0 ^ f_u_arrmul24_fa10_10_f_u_arrmul24_fa11_9_y2;
  assign f_u_arrmul24_fa10_10_y1 = f_u_arrmul24_fa10_10_f_u_arrmul24_and10_10_y0 & f_u_arrmul24_fa10_10_f_u_arrmul24_fa11_9_y2;
  assign f_u_arrmul24_fa10_10_y2 = f_u_arrmul24_fa10_10_y0 ^ f_u_arrmul24_fa10_10_f_u_arrmul24_fa9_10_y4;
  assign f_u_arrmul24_fa10_10_y3 = f_u_arrmul24_fa10_10_y0 & f_u_arrmul24_fa10_10_f_u_arrmul24_fa9_10_y4;
  assign f_u_arrmul24_fa10_10_y4 = f_u_arrmul24_fa10_10_y1 | f_u_arrmul24_fa10_10_y3;
  assign f_u_arrmul24_and11_10_a_11 = a_11;
  assign f_u_arrmul24_and11_10_b_10 = b_10;
  assign f_u_arrmul24_and11_10_y0 = f_u_arrmul24_and11_10_a_11 & f_u_arrmul24_and11_10_b_10;
  assign f_u_arrmul24_fa11_10_f_u_arrmul24_and11_10_y0 = f_u_arrmul24_and11_10_y0;
  assign f_u_arrmul24_fa11_10_f_u_arrmul24_fa12_9_y2 = f_u_arrmul24_fa12_9_y2;
  assign f_u_arrmul24_fa11_10_f_u_arrmul24_fa10_10_y4 = f_u_arrmul24_fa10_10_y4;
  assign f_u_arrmul24_fa11_10_y0 = f_u_arrmul24_fa11_10_f_u_arrmul24_and11_10_y0 ^ f_u_arrmul24_fa11_10_f_u_arrmul24_fa12_9_y2;
  assign f_u_arrmul24_fa11_10_y1 = f_u_arrmul24_fa11_10_f_u_arrmul24_and11_10_y0 & f_u_arrmul24_fa11_10_f_u_arrmul24_fa12_9_y2;
  assign f_u_arrmul24_fa11_10_y2 = f_u_arrmul24_fa11_10_y0 ^ f_u_arrmul24_fa11_10_f_u_arrmul24_fa10_10_y4;
  assign f_u_arrmul24_fa11_10_y3 = f_u_arrmul24_fa11_10_y0 & f_u_arrmul24_fa11_10_f_u_arrmul24_fa10_10_y4;
  assign f_u_arrmul24_fa11_10_y4 = f_u_arrmul24_fa11_10_y1 | f_u_arrmul24_fa11_10_y3;
  assign f_u_arrmul24_and12_10_a_12 = a_12;
  assign f_u_arrmul24_and12_10_b_10 = b_10;
  assign f_u_arrmul24_and12_10_y0 = f_u_arrmul24_and12_10_a_12 & f_u_arrmul24_and12_10_b_10;
  assign f_u_arrmul24_fa12_10_f_u_arrmul24_and12_10_y0 = f_u_arrmul24_and12_10_y0;
  assign f_u_arrmul24_fa12_10_f_u_arrmul24_fa13_9_y2 = f_u_arrmul24_fa13_9_y2;
  assign f_u_arrmul24_fa12_10_f_u_arrmul24_fa11_10_y4 = f_u_arrmul24_fa11_10_y4;
  assign f_u_arrmul24_fa12_10_y0 = f_u_arrmul24_fa12_10_f_u_arrmul24_and12_10_y0 ^ f_u_arrmul24_fa12_10_f_u_arrmul24_fa13_9_y2;
  assign f_u_arrmul24_fa12_10_y1 = f_u_arrmul24_fa12_10_f_u_arrmul24_and12_10_y0 & f_u_arrmul24_fa12_10_f_u_arrmul24_fa13_9_y2;
  assign f_u_arrmul24_fa12_10_y2 = f_u_arrmul24_fa12_10_y0 ^ f_u_arrmul24_fa12_10_f_u_arrmul24_fa11_10_y4;
  assign f_u_arrmul24_fa12_10_y3 = f_u_arrmul24_fa12_10_y0 & f_u_arrmul24_fa12_10_f_u_arrmul24_fa11_10_y4;
  assign f_u_arrmul24_fa12_10_y4 = f_u_arrmul24_fa12_10_y1 | f_u_arrmul24_fa12_10_y3;
  assign f_u_arrmul24_and13_10_a_13 = a_13;
  assign f_u_arrmul24_and13_10_b_10 = b_10;
  assign f_u_arrmul24_and13_10_y0 = f_u_arrmul24_and13_10_a_13 & f_u_arrmul24_and13_10_b_10;
  assign f_u_arrmul24_fa13_10_f_u_arrmul24_and13_10_y0 = f_u_arrmul24_and13_10_y0;
  assign f_u_arrmul24_fa13_10_f_u_arrmul24_fa14_9_y2 = f_u_arrmul24_fa14_9_y2;
  assign f_u_arrmul24_fa13_10_f_u_arrmul24_fa12_10_y4 = f_u_arrmul24_fa12_10_y4;
  assign f_u_arrmul24_fa13_10_y0 = f_u_arrmul24_fa13_10_f_u_arrmul24_and13_10_y0 ^ f_u_arrmul24_fa13_10_f_u_arrmul24_fa14_9_y2;
  assign f_u_arrmul24_fa13_10_y1 = f_u_arrmul24_fa13_10_f_u_arrmul24_and13_10_y0 & f_u_arrmul24_fa13_10_f_u_arrmul24_fa14_9_y2;
  assign f_u_arrmul24_fa13_10_y2 = f_u_arrmul24_fa13_10_y0 ^ f_u_arrmul24_fa13_10_f_u_arrmul24_fa12_10_y4;
  assign f_u_arrmul24_fa13_10_y3 = f_u_arrmul24_fa13_10_y0 & f_u_arrmul24_fa13_10_f_u_arrmul24_fa12_10_y4;
  assign f_u_arrmul24_fa13_10_y4 = f_u_arrmul24_fa13_10_y1 | f_u_arrmul24_fa13_10_y3;
  assign f_u_arrmul24_and14_10_a_14 = a_14;
  assign f_u_arrmul24_and14_10_b_10 = b_10;
  assign f_u_arrmul24_and14_10_y0 = f_u_arrmul24_and14_10_a_14 & f_u_arrmul24_and14_10_b_10;
  assign f_u_arrmul24_fa14_10_f_u_arrmul24_and14_10_y0 = f_u_arrmul24_and14_10_y0;
  assign f_u_arrmul24_fa14_10_f_u_arrmul24_fa15_9_y2 = f_u_arrmul24_fa15_9_y2;
  assign f_u_arrmul24_fa14_10_f_u_arrmul24_fa13_10_y4 = f_u_arrmul24_fa13_10_y4;
  assign f_u_arrmul24_fa14_10_y0 = f_u_arrmul24_fa14_10_f_u_arrmul24_and14_10_y0 ^ f_u_arrmul24_fa14_10_f_u_arrmul24_fa15_9_y2;
  assign f_u_arrmul24_fa14_10_y1 = f_u_arrmul24_fa14_10_f_u_arrmul24_and14_10_y0 & f_u_arrmul24_fa14_10_f_u_arrmul24_fa15_9_y2;
  assign f_u_arrmul24_fa14_10_y2 = f_u_arrmul24_fa14_10_y0 ^ f_u_arrmul24_fa14_10_f_u_arrmul24_fa13_10_y4;
  assign f_u_arrmul24_fa14_10_y3 = f_u_arrmul24_fa14_10_y0 & f_u_arrmul24_fa14_10_f_u_arrmul24_fa13_10_y4;
  assign f_u_arrmul24_fa14_10_y4 = f_u_arrmul24_fa14_10_y1 | f_u_arrmul24_fa14_10_y3;
  assign f_u_arrmul24_and15_10_a_15 = a_15;
  assign f_u_arrmul24_and15_10_b_10 = b_10;
  assign f_u_arrmul24_and15_10_y0 = f_u_arrmul24_and15_10_a_15 & f_u_arrmul24_and15_10_b_10;
  assign f_u_arrmul24_fa15_10_f_u_arrmul24_and15_10_y0 = f_u_arrmul24_and15_10_y0;
  assign f_u_arrmul24_fa15_10_f_u_arrmul24_fa16_9_y2 = f_u_arrmul24_fa16_9_y2;
  assign f_u_arrmul24_fa15_10_f_u_arrmul24_fa14_10_y4 = f_u_arrmul24_fa14_10_y4;
  assign f_u_arrmul24_fa15_10_y0 = f_u_arrmul24_fa15_10_f_u_arrmul24_and15_10_y0 ^ f_u_arrmul24_fa15_10_f_u_arrmul24_fa16_9_y2;
  assign f_u_arrmul24_fa15_10_y1 = f_u_arrmul24_fa15_10_f_u_arrmul24_and15_10_y0 & f_u_arrmul24_fa15_10_f_u_arrmul24_fa16_9_y2;
  assign f_u_arrmul24_fa15_10_y2 = f_u_arrmul24_fa15_10_y0 ^ f_u_arrmul24_fa15_10_f_u_arrmul24_fa14_10_y4;
  assign f_u_arrmul24_fa15_10_y3 = f_u_arrmul24_fa15_10_y0 & f_u_arrmul24_fa15_10_f_u_arrmul24_fa14_10_y4;
  assign f_u_arrmul24_fa15_10_y4 = f_u_arrmul24_fa15_10_y1 | f_u_arrmul24_fa15_10_y3;
  assign f_u_arrmul24_and16_10_a_16 = a_16;
  assign f_u_arrmul24_and16_10_b_10 = b_10;
  assign f_u_arrmul24_and16_10_y0 = f_u_arrmul24_and16_10_a_16 & f_u_arrmul24_and16_10_b_10;
  assign f_u_arrmul24_fa16_10_f_u_arrmul24_and16_10_y0 = f_u_arrmul24_and16_10_y0;
  assign f_u_arrmul24_fa16_10_f_u_arrmul24_fa17_9_y2 = f_u_arrmul24_fa17_9_y2;
  assign f_u_arrmul24_fa16_10_f_u_arrmul24_fa15_10_y4 = f_u_arrmul24_fa15_10_y4;
  assign f_u_arrmul24_fa16_10_y0 = f_u_arrmul24_fa16_10_f_u_arrmul24_and16_10_y0 ^ f_u_arrmul24_fa16_10_f_u_arrmul24_fa17_9_y2;
  assign f_u_arrmul24_fa16_10_y1 = f_u_arrmul24_fa16_10_f_u_arrmul24_and16_10_y0 & f_u_arrmul24_fa16_10_f_u_arrmul24_fa17_9_y2;
  assign f_u_arrmul24_fa16_10_y2 = f_u_arrmul24_fa16_10_y0 ^ f_u_arrmul24_fa16_10_f_u_arrmul24_fa15_10_y4;
  assign f_u_arrmul24_fa16_10_y3 = f_u_arrmul24_fa16_10_y0 & f_u_arrmul24_fa16_10_f_u_arrmul24_fa15_10_y4;
  assign f_u_arrmul24_fa16_10_y4 = f_u_arrmul24_fa16_10_y1 | f_u_arrmul24_fa16_10_y3;
  assign f_u_arrmul24_and17_10_a_17 = a_17;
  assign f_u_arrmul24_and17_10_b_10 = b_10;
  assign f_u_arrmul24_and17_10_y0 = f_u_arrmul24_and17_10_a_17 & f_u_arrmul24_and17_10_b_10;
  assign f_u_arrmul24_fa17_10_f_u_arrmul24_and17_10_y0 = f_u_arrmul24_and17_10_y0;
  assign f_u_arrmul24_fa17_10_f_u_arrmul24_fa18_9_y2 = f_u_arrmul24_fa18_9_y2;
  assign f_u_arrmul24_fa17_10_f_u_arrmul24_fa16_10_y4 = f_u_arrmul24_fa16_10_y4;
  assign f_u_arrmul24_fa17_10_y0 = f_u_arrmul24_fa17_10_f_u_arrmul24_and17_10_y0 ^ f_u_arrmul24_fa17_10_f_u_arrmul24_fa18_9_y2;
  assign f_u_arrmul24_fa17_10_y1 = f_u_arrmul24_fa17_10_f_u_arrmul24_and17_10_y0 & f_u_arrmul24_fa17_10_f_u_arrmul24_fa18_9_y2;
  assign f_u_arrmul24_fa17_10_y2 = f_u_arrmul24_fa17_10_y0 ^ f_u_arrmul24_fa17_10_f_u_arrmul24_fa16_10_y4;
  assign f_u_arrmul24_fa17_10_y3 = f_u_arrmul24_fa17_10_y0 & f_u_arrmul24_fa17_10_f_u_arrmul24_fa16_10_y4;
  assign f_u_arrmul24_fa17_10_y4 = f_u_arrmul24_fa17_10_y1 | f_u_arrmul24_fa17_10_y3;
  assign f_u_arrmul24_and18_10_a_18 = a_18;
  assign f_u_arrmul24_and18_10_b_10 = b_10;
  assign f_u_arrmul24_and18_10_y0 = f_u_arrmul24_and18_10_a_18 & f_u_arrmul24_and18_10_b_10;
  assign f_u_arrmul24_fa18_10_f_u_arrmul24_and18_10_y0 = f_u_arrmul24_and18_10_y0;
  assign f_u_arrmul24_fa18_10_f_u_arrmul24_fa19_9_y2 = f_u_arrmul24_fa19_9_y2;
  assign f_u_arrmul24_fa18_10_f_u_arrmul24_fa17_10_y4 = f_u_arrmul24_fa17_10_y4;
  assign f_u_arrmul24_fa18_10_y0 = f_u_arrmul24_fa18_10_f_u_arrmul24_and18_10_y0 ^ f_u_arrmul24_fa18_10_f_u_arrmul24_fa19_9_y2;
  assign f_u_arrmul24_fa18_10_y1 = f_u_arrmul24_fa18_10_f_u_arrmul24_and18_10_y0 & f_u_arrmul24_fa18_10_f_u_arrmul24_fa19_9_y2;
  assign f_u_arrmul24_fa18_10_y2 = f_u_arrmul24_fa18_10_y0 ^ f_u_arrmul24_fa18_10_f_u_arrmul24_fa17_10_y4;
  assign f_u_arrmul24_fa18_10_y3 = f_u_arrmul24_fa18_10_y0 & f_u_arrmul24_fa18_10_f_u_arrmul24_fa17_10_y4;
  assign f_u_arrmul24_fa18_10_y4 = f_u_arrmul24_fa18_10_y1 | f_u_arrmul24_fa18_10_y3;
  assign f_u_arrmul24_and19_10_a_19 = a_19;
  assign f_u_arrmul24_and19_10_b_10 = b_10;
  assign f_u_arrmul24_and19_10_y0 = f_u_arrmul24_and19_10_a_19 & f_u_arrmul24_and19_10_b_10;
  assign f_u_arrmul24_fa19_10_f_u_arrmul24_and19_10_y0 = f_u_arrmul24_and19_10_y0;
  assign f_u_arrmul24_fa19_10_f_u_arrmul24_fa20_9_y2 = f_u_arrmul24_fa20_9_y2;
  assign f_u_arrmul24_fa19_10_f_u_arrmul24_fa18_10_y4 = f_u_arrmul24_fa18_10_y4;
  assign f_u_arrmul24_fa19_10_y0 = f_u_arrmul24_fa19_10_f_u_arrmul24_and19_10_y0 ^ f_u_arrmul24_fa19_10_f_u_arrmul24_fa20_9_y2;
  assign f_u_arrmul24_fa19_10_y1 = f_u_arrmul24_fa19_10_f_u_arrmul24_and19_10_y0 & f_u_arrmul24_fa19_10_f_u_arrmul24_fa20_9_y2;
  assign f_u_arrmul24_fa19_10_y2 = f_u_arrmul24_fa19_10_y0 ^ f_u_arrmul24_fa19_10_f_u_arrmul24_fa18_10_y4;
  assign f_u_arrmul24_fa19_10_y3 = f_u_arrmul24_fa19_10_y0 & f_u_arrmul24_fa19_10_f_u_arrmul24_fa18_10_y4;
  assign f_u_arrmul24_fa19_10_y4 = f_u_arrmul24_fa19_10_y1 | f_u_arrmul24_fa19_10_y3;
  assign f_u_arrmul24_and20_10_a_20 = a_20;
  assign f_u_arrmul24_and20_10_b_10 = b_10;
  assign f_u_arrmul24_and20_10_y0 = f_u_arrmul24_and20_10_a_20 & f_u_arrmul24_and20_10_b_10;
  assign f_u_arrmul24_fa20_10_f_u_arrmul24_and20_10_y0 = f_u_arrmul24_and20_10_y0;
  assign f_u_arrmul24_fa20_10_f_u_arrmul24_fa21_9_y2 = f_u_arrmul24_fa21_9_y2;
  assign f_u_arrmul24_fa20_10_f_u_arrmul24_fa19_10_y4 = f_u_arrmul24_fa19_10_y4;
  assign f_u_arrmul24_fa20_10_y0 = f_u_arrmul24_fa20_10_f_u_arrmul24_and20_10_y0 ^ f_u_arrmul24_fa20_10_f_u_arrmul24_fa21_9_y2;
  assign f_u_arrmul24_fa20_10_y1 = f_u_arrmul24_fa20_10_f_u_arrmul24_and20_10_y0 & f_u_arrmul24_fa20_10_f_u_arrmul24_fa21_9_y2;
  assign f_u_arrmul24_fa20_10_y2 = f_u_arrmul24_fa20_10_y0 ^ f_u_arrmul24_fa20_10_f_u_arrmul24_fa19_10_y4;
  assign f_u_arrmul24_fa20_10_y3 = f_u_arrmul24_fa20_10_y0 & f_u_arrmul24_fa20_10_f_u_arrmul24_fa19_10_y4;
  assign f_u_arrmul24_fa20_10_y4 = f_u_arrmul24_fa20_10_y1 | f_u_arrmul24_fa20_10_y3;
  assign f_u_arrmul24_and21_10_a_21 = a_21;
  assign f_u_arrmul24_and21_10_b_10 = b_10;
  assign f_u_arrmul24_and21_10_y0 = f_u_arrmul24_and21_10_a_21 & f_u_arrmul24_and21_10_b_10;
  assign f_u_arrmul24_fa21_10_f_u_arrmul24_and21_10_y0 = f_u_arrmul24_and21_10_y0;
  assign f_u_arrmul24_fa21_10_f_u_arrmul24_fa22_9_y2 = f_u_arrmul24_fa22_9_y2;
  assign f_u_arrmul24_fa21_10_f_u_arrmul24_fa20_10_y4 = f_u_arrmul24_fa20_10_y4;
  assign f_u_arrmul24_fa21_10_y0 = f_u_arrmul24_fa21_10_f_u_arrmul24_and21_10_y0 ^ f_u_arrmul24_fa21_10_f_u_arrmul24_fa22_9_y2;
  assign f_u_arrmul24_fa21_10_y1 = f_u_arrmul24_fa21_10_f_u_arrmul24_and21_10_y0 & f_u_arrmul24_fa21_10_f_u_arrmul24_fa22_9_y2;
  assign f_u_arrmul24_fa21_10_y2 = f_u_arrmul24_fa21_10_y0 ^ f_u_arrmul24_fa21_10_f_u_arrmul24_fa20_10_y4;
  assign f_u_arrmul24_fa21_10_y3 = f_u_arrmul24_fa21_10_y0 & f_u_arrmul24_fa21_10_f_u_arrmul24_fa20_10_y4;
  assign f_u_arrmul24_fa21_10_y4 = f_u_arrmul24_fa21_10_y1 | f_u_arrmul24_fa21_10_y3;
  assign f_u_arrmul24_and22_10_a_22 = a_22;
  assign f_u_arrmul24_and22_10_b_10 = b_10;
  assign f_u_arrmul24_and22_10_y0 = f_u_arrmul24_and22_10_a_22 & f_u_arrmul24_and22_10_b_10;
  assign f_u_arrmul24_fa22_10_f_u_arrmul24_and22_10_y0 = f_u_arrmul24_and22_10_y0;
  assign f_u_arrmul24_fa22_10_f_u_arrmul24_fa23_9_y2 = f_u_arrmul24_fa23_9_y2;
  assign f_u_arrmul24_fa22_10_f_u_arrmul24_fa21_10_y4 = f_u_arrmul24_fa21_10_y4;
  assign f_u_arrmul24_fa22_10_y0 = f_u_arrmul24_fa22_10_f_u_arrmul24_and22_10_y0 ^ f_u_arrmul24_fa22_10_f_u_arrmul24_fa23_9_y2;
  assign f_u_arrmul24_fa22_10_y1 = f_u_arrmul24_fa22_10_f_u_arrmul24_and22_10_y0 & f_u_arrmul24_fa22_10_f_u_arrmul24_fa23_9_y2;
  assign f_u_arrmul24_fa22_10_y2 = f_u_arrmul24_fa22_10_y0 ^ f_u_arrmul24_fa22_10_f_u_arrmul24_fa21_10_y4;
  assign f_u_arrmul24_fa22_10_y3 = f_u_arrmul24_fa22_10_y0 & f_u_arrmul24_fa22_10_f_u_arrmul24_fa21_10_y4;
  assign f_u_arrmul24_fa22_10_y4 = f_u_arrmul24_fa22_10_y1 | f_u_arrmul24_fa22_10_y3;
  assign f_u_arrmul24_and23_10_a_23 = a_23;
  assign f_u_arrmul24_and23_10_b_10 = b_10;
  assign f_u_arrmul24_and23_10_y0 = f_u_arrmul24_and23_10_a_23 & f_u_arrmul24_and23_10_b_10;
  assign f_u_arrmul24_fa23_10_f_u_arrmul24_and23_10_y0 = f_u_arrmul24_and23_10_y0;
  assign f_u_arrmul24_fa23_10_f_u_arrmul24_fa23_9_y4 = f_u_arrmul24_fa23_9_y4;
  assign f_u_arrmul24_fa23_10_f_u_arrmul24_fa22_10_y4 = f_u_arrmul24_fa22_10_y4;
  assign f_u_arrmul24_fa23_10_y0 = f_u_arrmul24_fa23_10_f_u_arrmul24_and23_10_y0 ^ f_u_arrmul24_fa23_10_f_u_arrmul24_fa23_9_y4;
  assign f_u_arrmul24_fa23_10_y1 = f_u_arrmul24_fa23_10_f_u_arrmul24_and23_10_y0 & f_u_arrmul24_fa23_10_f_u_arrmul24_fa23_9_y4;
  assign f_u_arrmul24_fa23_10_y2 = f_u_arrmul24_fa23_10_y0 ^ f_u_arrmul24_fa23_10_f_u_arrmul24_fa22_10_y4;
  assign f_u_arrmul24_fa23_10_y3 = f_u_arrmul24_fa23_10_y0 & f_u_arrmul24_fa23_10_f_u_arrmul24_fa22_10_y4;
  assign f_u_arrmul24_fa23_10_y4 = f_u_arrmul24_fa23_10_y1 | f_u_arrmul24_fa23_10_y3;
  assign f_u_arrmul24_and0_11_a_0 = a_0;
  assign f_u_arrmul24_and0_11_b_11 = b_11;
  assign f_u_arrmul24_and0_11_y0 = f_u_arrmul24_and0_11_a_0 & f_u_arrmul24_and0_11_b_11;
  assign f_u_arrmul24_ha0_11_f_u_arrmul24_and0_11_y0 = f_u_arrmul24_and0_11_y0;
  assign f_u_arrmul24_ha0_11_f_u_arrmul24_fa1_10_y2 = f_u_arrmul24_fa1_10_y2;
  assign f_u_arrmul24_ha0_11_y0 = f_u_arrmul24_ha0_11_f_u_arrmul24_and0_11_y0 ^ f_u_arrmul24_ha0_11_f_u_arrmul24_fa1_10_y2;
  assign f_u_arrmul24_ha0_11_y1 = f_u_arrmul24_ha0_11_f_u_arrmul24_and0_11_y0 & f_u_arrmul24_ha0_11_f_u_arrmul24_fa1_10_y2;
  assign f_u_arrmul24_and1_11_a_1 = a_1;
  assign f_u_arrmul24_and1_11_b_11 = b_11;
  assign f_u_arrmul24_and1_11_y0 = f_u_arrmul24_and1_11_a_1 & f_u_arrmul24_and1_11_b_11;
  assign f_u_arrmul24_fa1_11_f_u_arrmul24_and1_11_y0 = f_u_arrmul24_and1_11_y0;
  assign f_u_arrmul24_fa1_11_f_u_arrmul24_fa2_10_y2 = f_u_arrmul24_fa2_10_y2;
  assign f_u_arrmul24_fa1_11_f_u_arrmul24_ha0_11_y1 = f_u_arrmul24_ha0_11_y1;
  assign f_u_arrmul24_fa1_11_y0 = f_u_arrmul24_fa1_11_f_u_arrmul24_and1_11_y0 ^ f_u_arrmul24_fa1_11_f_u_arrmul24_fa2_10_y2;
  assign f_u_arrmul24_fa1_11_y1 = f_u_arrmul24_fa1_11_f_u_arrmul24_and1_11_y0 & f_u_arrmul24_fa1_11_f_u_arrmul24_fa2_10_y2;
  assign f_u_arrmul24_fa1_11_y2 = f_u_arrmul24_fa1_11_y0 ^ f_u_arrmul24_fa1_11_f_u_arrmul24_ha0_11_y1;
  assign f_u_arrmul24_fa1_11_y3 = f_u_arrmul24_fa1_11_y0 & f_u_arrmul24_fa1_11_f_u_arrmul24_ha0_11_y1;
  assign f_u_arrmul24_fa1_11_y4 = f_u_arrmul24_fa1_11_y1 | f_u_arrmul24_fa1_11_y3;
  assign f_u_arrmul24_and2_11_a_2 = a_2;
  assign f_u_arrmul24_and2_11_b_11 = b_11;
  assign f_u_arrmul24_and2_11_y0 = f_u_arrmul24_and2_11_a_2 & f_u_arrmul24_and2_11_b_11;
  assign f_u_arrmul24_fa2_11_f_u_arrmul24_and2_11_y0 = f_u_arrmul24_and2_11_y0;
  assign f_u_arrmul24_fa2_11_f_u_arrmul24_fa3_10_y2 = f_u_arrmul24_fa3_10_y2;
  assign f_u_arrmul24_fa2_11_f_u_arrmul24_fa1_11_y4 = f_u_arrmul24_fa1_11_y4;
  assign f_u_arrmul24_fa2_11_y0 = f_u_arrmul24_fa2_11_f_u_arrmul24_and2_11_y0 ^ f_u_arrmul24_fa2_11_f_u_arrmul24_fa3_10_y2;
  assign f_u_arrmul24_fa2_11_y1 = f_u_arrmul24_fa2_11_f_u_arrmul24_and2_11_y0 & f_u_arrmul24_fa2_11_f_u_arrmul24_fa3_10_y2;
  assign f_u_arrmul24_fa2_11_y2 = f_u_arrmul24_fa2_11_y0 ^ f_u_arrmul24_fa2_11_f_u_arrmul24_fa1_11_y4;
  assign f_u_arrmul24_fa2_11_y3 = f_u_arrmul24_fa2_11_y0 & f_u_arrmul24_fa2_11_f_u_arrmul24_fa1_11_y4;
  assign f_u_arrmul24_fa2_11_y4 = f_u_arrmul24_fa2_11_y1 | f_u_arrmul24_fa2_11_y3;
  assign f_u_arrmul24_and3_11_a_3 = a_3;
  assign f_u_arrmul24_and3_11_b_11 = b_11;
  assign f_u_arrmul24_and3_11_y0 = f_u_arrmul24_and3_11_a_3 & f_u_arrmul24_and3_11_b_11;
  assign f_u_arrmul24_fa3_11_f_u_arrmul24_and3_11_y0 = f_u_arrmul24_and3_11_y0;
  assign f_u_arrmul24_fa3_11_f_u_arrmul24_fa4_10_y2 = f_u_arrmul24_fa4_10_y2;
  assign f_u_arrmul24_fa3_11_f_u_arrmul24_fa2_11_y4 = f_u_arrmul24_fa2_11_y4;
  assign f_u_arrmul24_fa3_11_y0 = f_u_arrmul24_fa3_11_f_u_arrmul24_and3_11_y0 ^ f_u_arrmul24_fa3_11_f_u_arrmul24_fa4_10_y2;
  assign f_u_arrmul24_fa3_11_y1 = f_u_arrmul24_fa3_11_f_u_arrmul24_and3_11_y0 & f_u_arrmul24_fa3_11_f_u_arrmul24_fa4_10_y2;
  assign f_u_arrmul24_fa3_11_y2 = f_u_arrmul24_fa3_11_y0 ^ f_u_arrmul24_fa3_11_f_u_arrmul24_fa2_11_y4;
  assign f_u_arrmul24_fa3_11_y3 = f_u_arrmul24_fa3_11_y0 & f_u_arrmul24_fa3_11_f_u_arrmul24_fa2_11_y4;
  assign f_u_arrmul24_fa3_11_y4 = f_u_arrmul24_fa3_11_y1 | f_u_arrmul24_fa3_11_y3;
  assign f_u_arrmul24_and4_11_a_4 = a_4;
  assign f_u_arrmul24_and4_11_b_11 = b_11;
  assign f_u_arrmul24_and4_11_y0 = f_u_arrmul24_and4_11_a_4 & f_u_arrmul24_and4_11_b_11;
  assign f_u_arrmul24_fa4_11_f_u_arrmul24_and4_11_y0 = f_u_arrmul24_and4_11_y0;
  assign f_u_arrmul24_fa4_11_f_u_arrmul24_fa5_10_y2 = f_u_arrmul24_fa5_10_y2;
  assign f_u_arrmul24_fa4_11_f_u_arrmul24_fa3_11_y4 = f_u_arrmul24_fa3_11_y4;
  assign f_u_arrmul24_fa4_11_y0 = f_u_arrmul24_fa4_11_f_u_arrmul24_and4_11_y0 ^ f_u_arrmul24_fa4_11_f_u_arrmul24_fa5_10_y2;
  assign f_u_arrmul24_fa4_11_y1 = f_u_arrmul24_fa4_11_f_u_arrmul24_and4_11_y0 & f_u_arrmul24_fa4_11_f_u_arrmul24_fa5_10_y2;
  assign f_u_arrmul24_fa4_11_y2 = f_u_arrmul24_fa4_11_y0 ^ f_u_arrmul24_fa4_11_f_u_arrmul24_fa3_11_y4;
  assign f_u_arrmul24_fa4_11_y3 = f_u_arrmul24_fa4_11_y0 & f_u_arrmul24_fa4_11_f_u_arrmul24_fa3_11_y4;
  assign f_u_arrmul24_fa4_11_y4 = f_u_arrmul24_fa4_11_y1 | f_u_arrmul24_fa4_11_y3;
  assign f_u_arrmul24_and5_11_a_5 = a_5;
  assign f_u_arrmul24_and5_11_b_11 = b_11;
  assign f_u_arrmul24_and5_11_y0 = f_u_arrmul24_and5_11_a_5 & f_u_arrmul24_and5_11_b_11;
  assign f_u_arrmul24_fa5_11_f_u_arrmul24_and5_11_y0 = f_u_arrmul24_and5_11_y0;
  assign f_u_arrmul24_fa5_11_f_u_arrmul24_fa6_10_y2 = f_u_arrmul24_fa6_10_y2;
  assign f_u_arrmul24_fa5_11_f_u_arrmul24_fa4_11_y4 = f_u_arrmul24_fa4_11_y4;
  assign f_u_arrmul24_fa5_11_y0 = f_u_arrmul24_fa5_11_f_u_arrmul24_and5_11_y0 ^ f_u_arrmul24_fa5_11_f_u_arrmul24_fa6_10_y2;
  assign f_u_arrmul24_fa5_11_y1 = f_u_arrmul24_fa5_11_f_u_arrmul24_and5_11_y0 & f_u_arrmul24_fa5_11_f_u_arrmul24_fa6_10_y2;
  assign f_u_arrmul24_fa5_11_y2 = f_u_arrmul24_fa5_11_y0 ^ f_u_arrmul24_fa5_11_f_u_arrmul24_fa4_11_y4;
  assign f_u_arrmul24_fa5_11_y3 = f_u_arrmul24_fa5_11_y0 & f_u_arrmul24_fa5_11_f_u_arrmul24_fa4_11_y4;
  assign f_u_arrmul24_fa5_11_y4 = f_u_arrmul24_fa5_11_y1 | f_u_arrmul24_fa5_11_y3;
  assign f_u_arrmul24_and6_11_a_6 = a_6;
  assign f_u_arrmul24_and6_11_b_11 = b_11;
  assign f_u_arrmul24_and6_11_y0 = f_u_arrmul24_and6_11_a_6 & f_u_arrmul24_and6_11_b_11;
  assign f_u_arrmul24_fa6_11_f_u_arrmul24_and6_11_y0 = f_u_arrmul24_and6_11_y0;
  assign f_u_arrmul24_fa6_11_f_u_arrmul24_fa7_10_y2 = f_u_arrmul24_fa7_10_y2;
  assign f_u_arrmul24_fa6_11_f_u_arrmul24_fa5_11_y4 = f_u_arrmul24_fa5_11_y4;
  assign f_u_arrmul24_fa6_11_y0 = f_u_arrmul24_fa6_11_f_u_arrmul24_and6_11_y0 ^ f_u_arrmul24_fa6_11_f_u_arrmul24_fa7_10_y2;
  assign f_u_arrmul24_fa6_11_y1 = f_u_arrmul24_fa6_11_f_u_arrmul24_and6_11_y0 & f_u_arrmul24_fa6_11_f_u_arrmul24_fa7_10_y2;
  assign f_u_arrmul24_fa6_11_y2 = f_u_arrmul24_fa6_11_y0 ^ f_u_arrmul24_fa6_11_f_u_arrmul24_fa5_11_y4;
  assign f_u_arrmul24_fa6_11_y3 = f_u_arrmul24_fa6_11_y0 & f_u_arrmul24_fa6_11_f_u_arrmul24_fa5_11_y4;
  assign f_u_arrmul24_fa6_11_y4 = f_u_arrmul24_fa6_11_y1 | f_u_arrmul24_fa6_11_y3;
  assign f_u_arrmul24_and7_11_a_7 = a_7;
  assign f_u_arrmul24_and7_11_b_11 = b_11;
  assign f_u_arrmul24_and7_11_y0 = f_u_arrmul24_and7_11_a_7 & f_u_arrmul24_and7_11_b_11;
  assign f_u_arrmul24_fa7_11_f_u_arrmul24_and7_11_y0 = f_u_arrmul24_and7_11_y0;
  assign f_u_arrmul24_fa7_11_f_u_arrmul24_fa8_10_y2 = f_u_arrmul24_fa8_10_y2;
  assign f_u_arrmul24_fa7_11_f_u_arrmul24_fa6_11_y4 = f_u_arrmul24_fa6_11_y4;
  assign f_u_arrmul24_fa7_11_y0 = f_u_arrmul24_fa7_11_f_u_arrmul24_and7_11_y0 ^ f_u_arrmul24_fa7_11_f_u_arrmul24_fa8_10_y2;
  assign f_u_arrmul24_fa7_11_y1 = f_u_arrmul24_fa7_11_f_u_arrmul24_and7_11_y0 & f_u_arrmul24_fa7_11_f_u_arrmul24_fa8_10_y2;
  assign f_u_arrmul24_fa7_11_y2 = f_u_arrmul24_fa7_11_y0 ^ f_u_arrmul24_fa7_11_f_u_arrmul24_fa6_11_y4;
  assign f_u_arrmul24_fa7_11_y3 = f_u_arrmul24_fa7_11_y0 & f_u_arrmul24_fa7_11_f_u_arrmul24_fa6_11_y4;
  assign f_u_arrmul24_fa7_11_y4 = f_u_arrmul24_fa7_11_y1 | f_u_arrmul24_fa7_11_y3;
  assign f_u_arrmul24_and8_11_a_8 = a_8;
  assign f_u_arrmul24_and8_11_b_11 = b_11;
  assign f_u_arrmul24_and8_11_y0 = f_u_arrmul24_and8_11_a_8 & f_u_arrmul24_and8_11_b_11;
  assign f_u_arrmul24_fa8_11_f_u_arrmul24_and8_11_y0 = f_u_arrmul24_and8_11_y0;
  assign f_u_arrmul24_fa8_11_f_u_arrmul24_fa9_10_y2 = f_u_arrmul24_fa9_10_y2;
  assign f_u_arrmul24_fa8_11_f_u_arrmul24_fa7_11_y4 = f_u_arrmul24_fa7_11_y4;
  assign f_u_arrmul24_fa8_11_y0 = f_u_arrmul24_fa8_11_f_u_arrmul24_and8_11_y0 ^ f_u_arrmul24_fa8_11_f_u_arrmul24_fa9_10_y2;
  assign f_u_arrmul24_fa8_11_y1 = f_u_arrmul24_fa8_11_f_u_arrmul24_and8_11_y0 & f_u_arrmul24_fa8_11_f_u_arrmul24_fa9_10_y2;
  assign f_u_arrmul24_fa8_11_y2 = f_u_arrmul24_fa8_11_y0 ^ f_u_arrmul24_fa8_11_f_u_arrmul24_fa7_11_y4;
  assign f_u_arrmul24_fa8_11_y3 = f_u_arrmul24_fa8_11_y0 & f_u_arrmul24_fa8_11_f_u_arrmul24_fa7_11_y4;
  assign f_u_arrmul24_fa8_11_y4 = f_u_arrmul24_fa8_11_y1 | f_u_arrmul24_fa8_11_y3;
  assign f_u_arrmul24_and9_11_a_9 = a_9;
  assign f_u_arrmul24_and9_11_b_11 = b_11;
  assign f_u_arrmul24_and9_11_y0 = f_u_arrmul24_and9_11_a_9 & f_u_arrmul24_and9_11_b_11;
  assign f_u_arrmul24_fa9_11_f_u_arrmul24_and9_11_y0 = f_u_arrmul24_and9_11_y0;
  assign f_u_arrmul24_fa9_11_f_u_arrmul24_fa10_10_y2 = f_u_arrmul24_fa10_10_y2;
  assign f_u_arrmul24_fa9_11_f_u_arrmul24_fa8_11_y4 = f_u_arrmul24_fa8_11_y4;
  assign f_u_arrmul24_fa9_11_y0 = f_u_arrmul24_fa9_11_f_u_arrmul24_and9_11_y0 ^ f_u_arrmul24_fa9_11_f_u_arrmul24_fa10_10_y2;
  assign f_u_arrmul24_fa9_11_y1 = f_u_arrmul24_fa9_11_f_u_arrmul24_and9_11_y0 & f_u_arrmul24_fa9_11_f_u_arrmul24_fa10_10_y2;
  assign f_u_arrmul24_fa9_11_y2 = f_u_arrmul24_fa9_11_y0 ^ f_u_arrmul24_fa9_11_f_u_arrmul24_fa8_11_y4;
  assign f_u_arrmul24_fa9_11_y3 = f_u_arrmul24_fa9_11_y0 & f_u_arrmul24_fa9_11_f_u_arrmul24_fa8_11_y4;
  assign f_u_arrmul24_fa9_11_y4 = f_u_arrmul24_fa9_11_y1 | f_u_arrmul24_fa9_11_y3;
  assign f_u_arrmul24_and10_11_a_10 = a_10;
  assign f_u_arrmul24_and10_11_b_11 = b_11;
  assign f_u_arrmul24_and10_11_y0 = f_u_arrmul24_and10_11_a_10 & f_u_arrmul24_and10_11_b_11;
  assign f_u_arrmul24_fa10_11_f_u_arrmul24_and10_11_y0 = f_u_arrmul24_and10_11_y0;
  assign f_u_arrmul24_fa10_11_f_u_arrmul24_fa11_10_y2 = f_u_arrmul24_fa11_10_y2;
  assign f_u_arrmul24_fa10_11_f_u_arrmul24_fa9_11_y4 = f_u_arrmul24_fa9_11_y4;
  assign f_u_arrmul24_fa10_11_y0 = f_u_arrmul24_fa10_11_f_u_arrmul24_and10_11_y0 ^ f_u_arrmul24_fa10_11_f_u_arrmul24_fa11_10_y2;
  assign f_u_arrmul24_fa10_11_y1 = f_u_arrmul24_fa10_11_f_u_arrmul24_and10_11_y0 & f_u_arrmul24_fa10_11_f_u_arrmul24_fa11_10_y2;
  assign f_u_arrmul24_fa10_11_y2 = f_u_arrmul24_fa10_11_y0 ^ f_u_arrmul24_fa10_11_f_u_arrmul24_fa9_11_y4;
  assign f_u_arrmul24_fa10_11_y3 = f_u_arrmul24_fa10_11_y0 & f_u_arrmul24_fa10_11_f_u_arrmul24_fa9_11_y4;
  assign f_u_arrmul24_fa10_11_y4 = f_u_arrmul24_fa10_11_y1 | f_u_arrmul24_fa10_11_y3;
  assign f_u_arrmul24_and11_11_a_11 = a_11;
  assign f_u_arrmul24_and11_11_b_11 = b_11;
  assign f_u_arrmul24_and11_11_y0 = f_u_arrmul24_and11_11_a_11 & f_u_arrmul24_and11_11_b_11;
  assign f_u_arrmul24_fa11_11_f_u_arrmul24_and11_11_y0 = f_u_arrmul24_and11_11_y0;
  assign f_u_arrmul24_fa11_11_f_u_arrmul24_fa12_10_y2 = f_u_arrmul24_fa12_10_y2;
  assign f_u_arrmul24_fa11_11_f_u_arrmul24_fa10_11_y4 = f_u_arrmul24_fa10_11_y4;
  assign f_u_arrmul24_fa11_11_y0 = f_u_arrmul24_fa11_11_f_u_arrmul24_and11_11_y0 ^ f_u_arrmul24_fa11_11_f_u_arrmul24_fa12_10_y2;
  assign f_u_arrmul24_fa11_11_y1 = f_u_arrmul24_fa11_11_f_u_arrmul24_and11_11_y0 & f_u_arrmul24_fa11_11_f_u_arrmul24_fa12_10_y2;
  assign f_u_arrmul24_fa11_11_y2 = f_u_arrmul24_fa11_11_y0 ^ f_u_arrmul24_fa11_11_f_u_arrmul24_fa10_11_y4;
  assign f_u_arrmul24_fa11_11_y3 = f_u_arrmul24_fa11_11_y0 & f_u_arrmul24_fa11_11_f_u_arrmul24_fa10_11_y4;
  assign f_u_arrmul24_fa11_11_y4 = f_u_arrmul24_fa11_11_y1 | f_u_arrmul24_fa11_11_y3;
  assign f_u_arrmul24_and12_11_a_12 = a_12;
  assign f_u_arrmul24_and12_11_b_11 = b_11;
  assign f_u_arrmul24_and12_11_y0 = f_u_arrmul24_and12_11_a_12 & f_u_arrmul24_and12_11_b_11;
  assign f_u_arrmul24_fa12_11_f_u_arrmul24_and12_11_y0 = f_u_arrmul24_and12_11_y0;
  assign f_u_arrmul24_fa12_11_f_u_arrmul24_fa13_10_y2 = f_u_arrmul24_fa13_10_y2;
  assign f_u_arrmul24_fa12_11_f_u_arrmul24_fa11_11_y4 = f_u_arrmul24_fa11_11_y4;
  assign f_u_arrmul24_fa12_11_y0 = f_u_arrmul24_fa12_11_f_u_arrmul24_and12_11_y0 ^ f_u_arrmul24_fa12_11_f_u_arrmul24_fa13_10_y2;
  assign f_u_arrmul24_fa12_11_y1 = f_u_arrmul24_fa12_11_f_u_arrmul24_and12_11_y0 & f_u_arrmul24_fa12_11_f_u_arrmul24_fa13_10_y2;
  assign f_u_arrmul24_fa12_11_y2 = f_u_arrmul24_fa12_11_y0 ^ f_u_arrmul24_fa12_11_f_u_arrmul24_fa11_11_y4;
  assign f_u_arrmul24_fa12_11_y3 = f_u_arrmul24_fa12_11_y0 & f_u_arrmul24_fa12_11_f_u_arrmul24_fa11_11_y4;
  assign f_u_arrmul24_fa12_11_y4 = f_u_arrmul24_fa12_11_y1 | f_u_arrmul24_fa12_11_y3;
  assign f_u_arrmul24_and13_11_a_13 = a_13;
  assign f_u_arrmul24_and13_11_b_11 = b_11;
  assign f_u_arrmul24_and13_11_y0 = f_u_arrmul24_and13_11_a_13 & f_u_arrmul24_and13_11_b_11;
  assign f_u_arrmul24_fa13_11_f_u_arrmul24_and13_11_y0 = f_u_arrmul24_and13_11_y0;
  assign f_u_arrmul24_fa13_11_f_u_arrmul24_fa14_10_y2 = f_u_arrmul24_fa14_10_y2;
  assign f_u_arrmul24_fa13_11_f_u_arrmul24_fa12_11_y4 = f_u_arrmul24_fa12_11_y4;
  assign f_u_arrmul24_fa13_11_y0 = f_u_arrmul24_fa13_11_f_u_arrmul24_and13_11_y0 ^ f_u_arrmul24_fa13_11_f_u_arrmul24_fa14_10_y2;
  assign f_u_arrmul24_fa13_11_y1 = f_u_arrmul24_fa13_11_f_u_arrmul24_and13_11_y0 & f_u_arrmul24_fa13_11_f_u_arrmul24_fa14_10_y2;
  assign f_u_arrmul24_fa13_11_y2 = f_u_arrmul24_fa13_11_y0 ^ f_u_arrmul24_fa13_11_f_u_arrmul24_fa12_11_y4;
  assign f_u_arrmul24_fa13_11_y3 = f_u_arrmul24_fa13_11_y0 & f_u_arrmul24_fa13_11_f_u_arrmul24_fa12_11_y4;
  assign f_u_arrmul24_fa13_11_y4 = f_u_arrmul24_fa13_11_y1 | f_u_arrmul24_fa13_11_y3;
  assign f_u_arrmul24_and14_11_a_14 = a_14;
  assign f_u_arrmul24_and14_11_b_11 = b_11;
  assign f_u_arrmul24_and14_11_y0 = f_u_arrmul24_and14_11_a_14 & f_u_arrmul24_and14_11_b_11;
  assign f_u_arrmul24_fa14_11_f_u_arrmul24_and14_11_y0 = f_u_arrmul24_and14_11_y0;
  assign f_u_arrmul24_fa14_11_f_u_arrmul24_fa15_10_y2 = f_u_arrmul24_fa15_10_y2;
  assign f_u_arrmul24_fa14_11_f_u_arrmul24_fa13_11_y4 = f_u_arrmul24_fa13_11_y4;
  assign f_u_arrmul24_fa14_11_y0 = f_u_arrmul24_fa14_11_f_u_arrmul24_and14_11_y0 ^ f_u_arrmul24_fa14_11_f_u_arrmul24_fa15_10_y2;
  assign f_u_arrmul24_fa14_11_y1 = f_u_arrmul24_fa14_11_f_u_arrmul24_and14_11_y0 & f_u_arrmul24_fa14_11_f_u_arrmul24_fa15_10_y2;
  assign f_u_arrmul24_fa14_11_y2 = f_u_arrmul24_fa14_11_y0 ^ f_u_arrmul24_fa14_11_f_u_arrmul24_fa13_11_y4;
  assign f_u_arrmul24_fa14_11_y3 = f_u_arrmul24_fa14_11_y0 & f_u_arrmul24_fa14_11_f_u_arrmul24_fa13_11_y4;
  assign f_u_arrmul24_fa14_11_y4 = f_u_arrmul24_fa14_11_y1 | f_u_arrmul24_fa14_11_y3;
  assign f_u_arrmul24_and15_11_a_15 = a_15;
  assign f_u_arrmul24_and15_11_b_11 = b_11;
  assign f_u_arrmul24_and15_11_y0 = f_u_arrmul24_and15_11_a_15 & f_u_arrmul24_and15_11_b_11;
  assign f_u_arrmul24_fa15_11_f_u_arrmul24_and15_11_y0 = f_u_arrmul24_and15_11_y0;
  assign f_u_arrmul24_fa15_11_f_u_arrmul24_fa16_10_y2 = f_u_arrmul24_fa16_10_y2;
  assign f_u_arrmul24_fa15_11_f_u_arrmul24_fa14_11_y4 = f_u_arrmul24_fa14_11_y4;
  assign f_u_arrmul24_fa15_11_y0 = f_u_arrmul24_fa15_11_f_u_arrmul24_and15_11_y0 ^ f_u_arrmul24_fa15_11_f_u_arrmul24_fa16_10_y2;
  assign f_u_arrmul24_fa15_11_y1 = f_u_arrmul24_fa15_11_f_u_arrmul24_and15_11_y0 & f_u_arrmul24_fa15_11_f_u_arrmul24_fa16_10_y2;
  assign f_u_arrmul24_fa15_11_y2 = f_u_arrmul24_fa15_11_y0 ^ f_u_arrmul24_fa15_11_f_u_arrmul24_fa14_11_y4;
  assign f_u_arrmul24_fa15_11_y3 = f_u_arrmul24_fa15_11_y0 & f_u_arrmul24_fa15_11_f_u_arrmul24_fa14_11_y4;
  assign f_u_arrmul24_fa15_11_y4 = f_u_arrmul24_fa15_11_y1 | f_u_arrmul24_fa15_11_y3;
  assign f_u_arrmul24_and16_11_a_16 = a_16;
  assign f_u_arrmul24_and16_11_b_11 = b_11;
  assign f_u_arrmul24_and16_11_y0 = f_u_arrmul24_and16_11_a_16 & f_u_arrmul24_and16_11_b_11;
  assign f_u_arrmul24_fa16_11_f_u_arrmul24_and16_11_y0 = f_u_arrmul24_and16_11_y0;
  assign f_u_arrmul24_fa16_11_f_u_arrmul24_fa17_10_y2 = f_u_arrmul24_fa17_10_y2;
  assign f_u_arrmul24_fa16_11_f_u_arrmul24_fa15_11_y4 = f_u_arrmul24_fa15_11_y4;
  assign f_u_arrmul24_fa16_11_y0 = f_u_arrmul24_fa16_11_f_u_arrmul24_and16_11_y0 ^ f_u_arrmul24_fa16_11_f_u_arrmul24_fa17_10_y2;
  assign f_u_arrmul24_fa16_11_y1 = f_u_arrmul24_fa16_11_f_u_arrmul24_and16_11_y0 & f_u_arrmul24_fa16_11_f_u_arrmul24_fa17_10_y2;
  assign f_u_arrmul24_fa16_11_y2 = f_u_arrmul24_fa16_11_y0 ^ f_u_arrmul24_fa16_11_f_u_arrmul24_fa15_11_y4;
  assign f_u_arrmul24_fa16_11_y3 = f_u_arrmul24_fa16_11_y0 & f_u_arrmul24_fa16_11_f_u_arrmul24_fa15_11_y4;
  assign f_u_arrmul24_fa16_11_y4 = f_u_arrmul24_fa16_11_y1 | f_u_arrmul24_fa16_11_y3;
  assign f_u_arrmul24_and17_11_a_17 = a_17;
  assign f_u_arrmul24_and17_11_b_11 = b_11;
  assign f_u_arrmul24_and17_11_y0 = f_u_arrmul24_and17_11_a_17 & f_u_arrmul24_and17_11_b_11;
  assign f_u_arrmul24_fa17_11_f_u_arrmul24_and17_11_y0 = f_u_arrmul24_and17_11_y0;
  assign f_u_arrmul24_fa17_11_f_u_arrmul24_fa18_10_y2 = f_u_arrmul24_fa18_10_y2;
  assign f_u_arrmul24_fa17_11_f_u_arrmul24_fa16_11_y4 = f_u_arrmul24_fa16_11_y4;
  assign f_u_arrmul24_fa17_11_y0 = f_u_arrmul24_fa17_11_f_u_arrmul24_and17_11_y0 ^ f_u_arrmul24_fa17_11_f_u_arrmul24_fa18_10_y2;
  assign f_u_arrmul24_fa17_11_y1 = f_u_arrmul24_fa17_11_f_u_arrmul24_and17_11_y0 & f_u_arrmul24_fa17_11_f_u_arrmul24_fa18_10_y2;
  assign f_u_arrmul24_fa17_11_y2 = f_u_arrmul24_fa17_11_y0 ^ f_u_arrmul24_fa17_11_f_u_arrmul24_fa16_11_y4;
  assign f_u_arrmul24_fa17_11_y3 = f_u_arrmul24_fa17_11_y0 & f_u_arrmul24_fa17_11_f_u_arrmul24_fa16_11_y4;
  assign f_u_arrmul24_fa17_11_y4 = f_u_arrmul24_fa17_11_y1 | f_u_arrmul24_fa17_11_y3;
  assign f_u_arrmul24_and18_11_a_18 = a_18;
  assign f_u_arrmul24_and18_11_b_11 = b_11;
  assign f_u_arrmul24_and18_11_y0 = f_u_arrmul24_and18_11_a_18 & f_u_arrmul24_and18_11_b_11;
  assign f_u_arrmul24_fa18_11_f_u_arrmul24_and18_11_y0 = f_u_arrmul24_and18_11_y0;
  assign f_u_arrmul24_fa18_11_f_u_arrmul24_fa19_10_y2 = f_u_arrmul24_fa19_10_y2;
  assign f_u_arrmul24_fa18_11_f_u_arrmul24_fa17_11_y4 = f_u_arrmul24_fa17_11_y4;
  assign f_u_arrmul24_fa18_11_y0 = f_u_arrmul24_fa18_11_f_u_arrmul24_and18_11_y0 ^ f_u_arrmul24_fa18_11_f_u_arrmul24_fa19_10_y2;
  assign f_u_arrmul24_fa18_11_y1 = f_u_arrmul24_fa18_11_f_u_arrmul24_and18_11_y0 & f_u_arrmul24_fa18_11_f_u_arrmul24_fa19_10_y2;
  assign f_u_arrmul24_fa18_11_y2 = f_u_arrmul24_fa18_11_y0 ^ f_u_arrmul24_fa18_11_f_u_arrmul24_fa17_11_y4;
  assign f_u_arrmul24_fa18_11_y3 = f_u_arrmul24_fa18_11_y0 & f_u_arrmul24_fa18_11_f_u_arrmul24_fa17_11_y4;
  assign f_u_arrmul24_fa18_11_y4 = f_u_arrmul24_fa18_11_y1 | f_u_arrmul24_fa18_11_y3;
  assign f_u_arrmul24_and19_11_a_19 = a_19;
  assign f_u_arrmul24_and19_11_b_11 = b_11;
  assign f_u_arrmul24_and19_11_y0 = f_u_arrmul24_and19_11_a_19 & f_u_arrmul24_and19_11_b_11;
  assign f_u_arrmul24_fa19_11_f_u_arrmul24_and19_11_y0 = f_u_arrmul24_and19_11_y0;
  assign f_u_arrmul24_fa19_11_f_u_arrmul24_fa20_10_y2 = f_u_arrmul24_fa20_10_y2;
  assign f_u_arrmul24_fa19_11_f_u_arrmul24_fa18_11_y4 = f_u_arrmul24_fa18_11_y4;
  assign f_u_arrmul24_fa19_11_y0 = f_u_arrmul24_fa19_11_f_u_arrmul24_and19_11_y0 ^ f_u_arrmul24_fa19_11_f_u_arrmul24_fa20_10_y2;
  assign f_u_arrmul24_fa19_11_y1 = f_u_arrmul24_fa19_11_f_u_arrmul24_and19_11_y0 & f_u_arrmul24_fa19_11_f_u_arrmul24_fa20_10_y2;
  assign f_u_arrmul24_fa19_11_y2 = f_u_arrmul24_fa19_11_y0 ^ f_u_arrmul24_fa19_11_f_u_arrmul24_fa18_11_y4;
  assign f_u_arrmul24_fa19_11_y3 = f_u_arrmul24_fa19_11_y0 & f_u_arrmul24_fa19_11_f_u_arrmul24_fa18_11_y4;
  assign f_u_arrmul24_fa19_11_y4 = f_u_arrmul24_fa19_11_y1 | f_u_arrmul24_fa19_11_y3;
  assign f_u_arrmul24_and20_11_a_20 = a_20;
  assign f_u_arrmul24_and20_11_b_11 = b_11;
  assign f_u_arrmul24_and20_11_y0 = f_u_arrmul24_and20_11_a_20 & f_u_arrmul24_and20_11_b_11;
  assign f_u_arrmul24_fa20_11_f_u_arrmul24_and20_11_y0 = f_u_arrmul24_and20_11_y0;
  assign f_u_arrmul24_fa20_11_f_u_arrmul24_fa21_10_y2 = f_u_arrmul24_fa21_10_y2;
  assign f_u_arrmul24_fa20_11_f_u_arrmul24_fa19_11_y4 = f_u_arrmul24_fa19_11_y4;
  assign f_u_arrmul24_fa20_11_y0 = f_u_arrmul24_fa20_11_f_u_arrmul24_and20_11_y0 ^ f_u_arrmul24_fa20_11_f_u_arrmul24_fa21_10_y2;
  assign f_u_arrmul24_fa20_11_y1 = f_u_arrmul24_fa20_11_f_u_arrmul24_and20_11_y0 & f_u_arrmul24_fa20_11_f_u_arrmul24_fa21_10_y2;
  assign f_u_arrmul24_fa20_11_y2 = f_u_arrmul24_fa20_11_y0 ^ f_u_arrmul24_fa20_11_f_u_arrmul24_fa19_11_y4;
  assign f_u_arrmul24_fa20_11_y3 = f_u_arrmul24_fa20_11_y0 & f_u_arrmul24_fa20_11_f_u_arrmul24_fa19_11_y4;
  assign f_u_arrmul24_fa20_11_y4 = f_u_arrmul24_fa20_11_y1 | f_u_arrmul24_fa20_11_y3;
  assign f_u_arrmul24_and21_11_a_21 = a_21;
  assign f_u_arrmul24_and21_11_b_11 = b_11;
  assign f_u_arrmul24_and21_11_y0 = f_u_arrmul24_and21_11_a_21 & f_u_arrmul24_and21_11_b_11;
  assign f_u_arrmul24_fa21_11_f_u_arrmul24_and21_11_y0 = f_u_arrmul24_and21_11_y0;
  assign f_u_arrmul24_fa21_11_f_u_arrmul24_fa22_10_y2 = f_u_arrmul24_fa22_10_y2;
  assign f_u_arrmul24_fa21_11_f_u_arrmul24_fa20_11_y4 = f_u_arrmul24_fa20_11_y4;
  assign f_u_arrmul24_fa21_11_y0 = f_u_arrmul24_fa21_11_f_u_arrmul24_and21_11_y0 ^ f_u_arrmul24_fa21_11_f_u_arrmul24_fa22_10_y2;
  assign f_u_arrmul24_fa21_11_y1 = f_u_arrmul24_fa21_11_f_u_arrmul24_and21_11_y0 & f_u_arrmul24_fa21_11_f_u_arrmul24_fa22_10_y2;
  assign f_u_arrmul24_fa21_11_y2 = f_u_arrmul24_fa21_11_y0 ^ f_u_arrmul24_fa21_11_f_u_arrmul24_fa20_11_y4;
  assign f_u_arrmul24_fa21_11_y3 = f_u_arrmul24_fa21_11_y0 & f_u_arrmul24_fa21_11_f_u_arrmul24_fa20_11_y4;
  assign f_u_arrmul24_fa21_11_y4 = f_u_arrmul24_fa21_11_y1 | f_u_arrmul24_fa21_11_y3;
  assign f_u_arrmul24_and22_11_a_22 = a_22;
  assign f_u_arrmul24_and22_11_b_11 = b_11;
  assign f_u_arrmul24_and22_11_y0 = f_u_arrmul24_and22_11_a_22 & f_u_arrmul24_and22_11_b_11;
  assign f_u_arrmul24_fa22_11_f_u_arrmul24_and22_11_y0 = f_u_arrmul24_and22_11_y0;
  assign f_u_arrmul24_fa22_11_f_u_arrmul24_fa23_10_y2 = f_u_arrmul24_fa23_10_y2;
  assign f_u_arrmul24_fa22_11_f_u_arrmul24_fa21_11_y4 = f_u_arrmul24_fa21_11_y4;
  assign f_u_arrmul24_fa22_11_y0 = f_u_arrmul24_fa22_11_f_u_arrmul24_and22_11_y0 ^ f_u_arrmul24_fa22_11_f_u_arrmul24_fa23_10_y2;
  assign f_u_arrmul24_fa22_11_y1 = f_u_arrmul24_fa22_11_f_u_arrmul24_and22_11_y0 & f_u_arrmul24_fa22_11_f_u_arrmul24_fa23_10_y2;
  assign f_u_arrmul24_fa22_11_y2 = f_u_arrmul24_fa22_11_y0 ^ f_u_arrmul24_fa22_11_f_u_arrmul24_fa21_11_y4;
  assign f_u_arrmul24_fa22_11_y3 = f_u_arrmul24_fa22_11_y0 & f_u_arrmul24_fa22_11_f_u_arrmul24_fa21_11_y4;
  assign f_u_arrmul24_fa22_11_y4 = f_u_arrmul24_fa22_11_y1 | f_u_arrmul24_fa22_11_y3;
  assign f_u_arrmul24_and23_11_a_23 = a_23;
  assign f_u_arrmul24_and23_11_b_11 = b_11;
  assign f_u_arrmul24_and23_11_y0 = f_u_arrmul24_and23_11_a_23 & f_u_arrmul24_and23_11_b_11;
  assign f_u_arrmul24_fa23_11_f_u_arrmul24_and23_11_y0 = f_u_arrmul24_and23_11_y0;
  assign f_u_arrmul24_fa23_11_f_u_arrmul24_fa23_10_y4 = f_u_arrmul24_fa23_10_y4;
  assign f_u_arrmul24_fa23_11_f_u_arrmul24_fa22_11_y4 = f_u_arrmul24_fa22_11_y4;
  assign f_u_arrmul24_fa23_11_y0 = f_u_arrmul24_fa23_11_f_u_arrmul24_and23_11_y0 ^ f_u_arrmul24_fa23_11_f_u_arrmul24_fa23_10_y4;
  assign f_u_arrmul24_fa23_11_y1 = f_u_arrmul24_fa23_11_f_u_arrmul24_and23_11_y0 & f_u_arrmul24_fa23_11_f_u_arrmul24_fa23_10_y4;
  assign f_u_arrmul24_fa23_11_y2 = f_u_arrmul24_fa23_11_y0 ^ f_u_arrmul24_fa23_11_f_u_arrmul24_fa22_11_y4;
  assign f_u_arrmul24_fa23_11_y3 = f_u_arrmul24_fa23_11_y0 & f_u_arrmul24_fa23_11_f_u_arrmul24_fa22_11_y4;
  assign f_u_arrmul24_fa23_11_y4 = f_u_arrmul24_fa23_11_y1 | f_u_arrmul24_fa23_11_y3;
  assign f_u_arrmul24_and0_12_a_0 = a_0;
  assign f_u_arrmul24_and0_12_b_12 = b_12;
  assign f_u_arrmul24_and0_12_y0 = f_u_arrmul24_and0_12_a_0 & f_u_arrmul24_and0_12_b_12;
  assign f_u_arrmul24_ha0_12_f_u_arrmul24_and0_12_y0 = f_u_arrmul24_and0_12_y0;
  assign f_u_arrmul24_ha0_12_f_u_arrmul24_fa1_11_y2 = f_u_arrmul24_fa1_11_y2;
  assign f_u_arrmul24_ha0_12_y0 = f_u_arrmul24_ha0_12_f_u_arrmul24_and0_12_y0 ^ f_u_arrmul24_ha0_12_f_u_arrmul24_fa1_11_y2;
  assign f_u_arrmul24_ha0_12_y1 = f_u_arrmul24_ha0_12_f_u_arrmul24_and0_12_y0 & f_u_arrmul24_ha0_12_f_u_arrmul24_fa1_11_y2;
  assign f_u_arrmul24_and1_12_a_1 = a_1;
  assign f_u_arrmul24_and1_12_b_12 = b_12;
  assign f_u_arrmul24_and1_12_y0 = f_u_arrmul24_and1_12_a_1 & f_u_arrmul24_and1_12_b_12;
  assign f_u_arrmul24_fa1_12_f_u_arrmul24_and1_12_y0 = f_u_arrmul24_and1_12_y0;
  assign f_u_arrmul24_fa1_12_f_u_arrmul24_fa2_11_y2 = f_u_arrmul24_fa2_11_y2;
  assign f_u_arrmul24_fa1_12_f_u_arrmul24_ha0_12_y1 = f_u_arrmul24_ha0_12_y1;
  assign f_u_arrmul24_fa1_12_y0 = f_u_arrmul24_fa1_12_f_u_arrmul24_and1_12_y0 ^ f_u_arrmul24_fa1_12_f_u_arrmul24_fa2_11_y2;
  assign f_u_arrmul24_fa1_12_y1 = f_u_arrmul24_fa1_12_f_u_arrmul24_and1_12_y0 & f_u_arrmul24_fa1_12_f_u_arrmul24_fa2_11_y2;
  assign f_u_arrmul24_fa1_12_y2 = f_u_arrmul24_fa1_12_y0 ^ f_u_arrmul24_fa1_12_f_u_arrmul24_ha0_12_y1;
  assign f_u_arrmul24_fa1_12_y3 = f_u_arrmul24_fa1_12_y0 & f_u_arrmul24_fa1_12_f_u_arrmul24_ha0_12_y1;
  assign f_u_arrmul24_fa1_12_y4 = f_u_arrmul24_fa1_12_y1 | f_u_arrmul24_fa1_12_y3;
  assign f_u_arrmul24_and2_12_a_2 = a_2;
  assign f_u_arrmul24_and2_12_b_12 = b_12;
  assign f_u_arrmul24_and2_12_y0 = f_u_arrmul24_and2_12_a_2 & f_u_arrmul24_and2_12_b_12;
  assign f_u_arrmul24_fa2_12_f_u_arrmul24_and2_12_y0 = f_u_arrmul24_and2_12_y0;
  assign f_u_arrmul24_fa2_12_f_u_arrmul24_fa3_11_y2 = f_u_arrmul24_fa3_11_y2;
  assign f_u_arrmul24_fa2_12_f_u_arrmul24_fa1_12_y4 = f_u_arrmul24_fa1_12_y4;
  assign f_u_arrmul24_fa2_12_y0 = f_u_arrmul24_fa2_12_f_u_arrmul24_and2_12_y0 ^ f_u_arrmul24_fa2_12_f_u_arrmul24_fa3_11_y2;
  assign f_u_arrmul24_fa2_12_y1 = f_u_arrmul24_fa2_12_f_u_arrmul24_and2_12_y0 & f_u_arrmul24_fa2_12_f_u_arrmul24_fa3_11_y2;
  assign f_u_arrmul24_fa2_12_y2 = f_u_arrmul24_fa2_12_y0 ^ f_u_arrmul24_fa2_12_f_u_arrmul24_fa1_12_y4;
  assign f_u_arrmul24_fa2_12_y3 = f_u_arrmul24_fa2_12_y0 & f_u_arrmul24_fa2_12_f_u_arrmul24_fa1_12_y4;
  assign f_u_arrmul24_fa2_12_y4 = f_u_arrmul24_fa2_12_y1 | f_u_arrmul24_fa2_12_y3;
  assign f_u_arrmul24_and3_12_a_3 = a_3;
  assign f_u_arrmul24_and3_12_b_12 = b_12;
  assign f_u_arrmul24_and3_12_y0 = f_u_arrmul24_and3_12_a_3 & f_u_arrmul24_and3_12_b_12;
  assign f_u_arrmul24_fa3_12_f_u_arrmul24_and3_12_y0 = f_u_arrmul24_and3_12_y0;
  assign f_u_arrmul24_fa3_12_f_u_arrmul24_fa4_11_y2 = f_u_arrmul24_fa4_11_y2;
  assign f_u_arrmul24_fa3_12_f_u_arrmul24_fa2_12_y4 = f_u_arrmul24_fa2_12_y4;
  assign f_u_arrmul24_fa3_12_y0 = f_u_arrmul24_fa3_12_f_u_arrmul24_and3_12_y0 ^ f_u_arrmul24_fa3_12_f_u_arrmul24_fa4_11_y2;
  assign f_u_arrmul24_fa3_12_y1 = f_u_arrmul24_fa3_12_f_u_arrmul24_and3_12_y0 & f_u_arrmul24_fa3_12_f_u_arrmul24_fa4_11_y2;
  assign f_u_arrmul24_fa3_12_y2 = f_u_arrmul24_fa3_12_y0 ^ f_u_arrmul24_fa3_12_f_u_arrmul24_fa2_12_y4;
  assign f_u_arrmul24_fa3_12_y3 = f_u_arrmul24_fa3_12_y0 & f_u_arrmul24_fa3_12_f_u_arrmul24_fa2_12_y4;
  assign f_u_arrmul24_fa3_12_y4 = f_u_arrmul24_fa3_12_y1 | f_u_arrmul24_fa3_12_y3;
  assign f_u_arrmul24_and4_12_a_4 = a_4;
  assign f_u_arrmul24_and4_12_b_12 = b_12;
  assign f_u_arrmul24_and4_12_y0 = f_u_arrmul24_and4_12_a_4 & f_u_arrmul24_and4_12_b_12;
  assign f_u_arrmul24_fa4_12_f_u_arrmul24_and4_12_y0 = f_u_arrmul24_and4_12_y0;
  assign f_u_arrmul24_fa4_12_f_u_arrmul24_fa5_11_y2 = f_u_arrmul24_fa5_11_y2;
  assign f_u_arrmul24_fa4_12_f_u_arrmul24_fa3_12_y4 = f_u_arrmul24_fa3_12_y4;
  assign f_u_arrmul24_fa4_12_y0 = f_u_arrmul24_fa4_12_f_u_arrmul24_and4_12_y0 ^ f_u_arrmul24_fa4_12_f_u_arrmul24_fa5_11_y2;
  assign f_u_arrmul24_fa4_12_y1 = f_u_arrmul24_fa4_12_f_u_arrmul24_and4_12_y0 & f_u_arrmul24_fa4_12_f_u_arrmul24_fa5_11_y2;
  assign f_u_arrmul24_fa4_12_y2 = f_u_arrmul24_fa4_12_y0 ^ f_u_arrmul24_fa4_12_f_u_arrmul24_fa3_12_y4;
  assign f_u_arrmul24_fa4_12_y3 = f_u_arrmul24_fa4_12_y0 & f_u_arrmul24_fa4_12_f_u_arrmul24_fa3_12_y4;
  assign f_u_arrmul24_fa4_12_y4 = f_u_arrmul24_fa4_12_y1 | f_u_arrmul24_fa4_12_y3;
  assign f_u_arrmul24_and5_12_a_5 = a_5;
  assign f_u_arrmul24_and5_12_b_12 = b_12;
  assign f_u_arrmul24_and5_12_y0 = f_u_arrmul24_and5_12_a_5 & f_u_arrmul24_and5_12_b_12;
  assign f_u_arrmul24_fa5_12_f_u_arrmul24_and5_12_y0 = f_u_arrmul24_and5_12_y0;
  assign f_u_arrmul24_fa5_12_f_u_arrmul24_fa6_11_y2 = f_u_arrmul24_fa6_11_y2;
  assign f_u_arrmul24_fa5_12_f_u_arrmul24_fa4_12_y4 = f_u_arrmul24_fa4_12_y4;
  assign f_u_arrmul24_fa5_12_y0 = f_u_arrmul24_fa5_12_f_u_arrmul24_and5_12_y0 ^ f_u_arrmul24_fa5_12_f_u_arrmul24_fa6_11_y2;
  assign f_u_arrmul24_fa5_12_y1 = f_u_arrmul24_fa5_12_f_u_arrmul24_and5_12_y0 & f_u_arrmul24_fa5_12_f_u_arrmul24_fa6_11_y2;
  assign f_u_arrmul24_fa5_12_y2 = f_u_arrmul24_fa5_12_y0 ^ f_u_arrmul24_fa5_12_f_u_arrmul24_fa4_12_y4;
  assign f_u_arrmul24_fa5_12_y3 = f_u_arrmul24_fa5_12_y0 & f_u_arrmul24_fa5_12_f_u_arrmul24_fa4_12_y4;
  assign f_u_arrmul24_fa5_12_y4 = f_u_arrmul24_fa5_12_y1 | f_u_arrmul24_fa5_12_y3;
  assign f_u_arrmul24_and6_12_a_6 = a_6;
  assign f_u_arrmul24_and6_12_b_12 = b_12;
  assign f_u_arrmul24_and6_12_y0 = f_u_arrmul24_and6_12_a_6 & f_u_arrmul24_and6_12_b_12;
  assign f_u_arrmul24_fa6_12_f_u_arrmul24_and6_12_y0 = f_u_arrmul24_and6_12_y0;
  assign f_u_arrmul24_fa6_12_f_u_arrmul24_fa7_11_y2 = f_u_arrmul24_fa7_11_y2;
  assign f_u_arrmul24_fa6_12_f_u_arrmul24_fa5_12_y4 = f_u_arrmul24_fa5_12_y4;
  assign f_u_arrmul24_fa6_12_y0 = f_u_arrmul24_fa6_12_f_u_arrmul24_and6_12_y0 ^ f_u_arrmul24_fa6_12_f_u_arrmul24_fa7_11_y2;
  assign f_u_arrmul24_fa6_12_y1 = f_u_arrmul24_fa6_12_f_u_arrmul24_and6_12_y0 & f_u_arrmul24_fa6_12_f_u_arrmul24_fa7_11_y2;
  assign f_u_arrmul24_fa6_12_y2 = f_u_arrmul24_fa6_12_y0 ^ f_u_arrmul24_fa6_12_f_u_arrmul24_fa5_12_y4;
  assign f_u_arrmul24_fa6_12_y3 = f_u_arrmul24_fa6_12_y0 & f_u_arrmul24_fa6_12_f_u_arrmul24_fa5_12_y4;
  assign f_u_arrmul24_fa6_12_y4 = f_u_arrmul24_fa6_12_y1 | f_u_arrmul24_fa6_12_y3;
  assign f_u_arrmul24_and7_12_a_7 = a_7;
  assign f_u_arrmul24_and7_12_b_12 = b_12;
  assign f_u_arrmul24_and7_12_y0 = f_u_arrmul24_and7_12_a_7 & f_u_arrmul24_and7_12_b_12;
  assign f_u_arrmul24_fa7_12_f_u_arrmul24_and7_12_y0 = f_u_arrmul24_and7_12_y0;
  assign f_u_arrmul24_fa7_12_f_u_arrmul24_fa8_11_y2 = f_u_arrmul24_fa8_11_y2;
  assign f_u_arrmul24_fa7_12_f_u_arrmul24_fa6_12_y4 = f_u_arrmul24_fa6_12_y4;
  assign f_u_arrmul24_fa7_12_y0 = f_u_arrmul24_fa7_12_f_u_arrmul24_and7_12_y0 ^ f_u_arrmul24_fa7_12_f_u_arrmul24_fa8_11_y2;
  assign f_u_arrmul24_fa7_12_y1 = f_u_arrmul24_fa7_12_f_u_arrmul24_and7_12_y0 & f_u_arrmul24_fa7_12_f_u_arrmul24_fa8_11_y2;
  assign f_u_arrmul24_fa7_12_y2 = f_u_arrmul24_fa7_12_y0 ^ f_u_arrmul24_fa7_12_f_u_arrmul24_fa6_12_y4;
  assign f_u_arrmul24_fa7_12_y3 = f_u_arrmul24_fa7_12_y0 & f_u_arrmul24_fa7_12_f_u_arrmul24_fa6_12_y4;
  assign f_u_arrmul24_fa7_12_y4 = f_u_arrmul24_fa7_12_y1 | f_u_arrmul24_fa7_12_y3;
  assign f_u_arrmul24_and8_12_a_8 = a_8;
  assign f_u_arrmul24_and8_12_b_12 = b_12;
  assign f_u_arrmul24_and8_12_y0 = f_u_arrmul24_and8_12_a_8 & f_u_arrmul24_and8_12_b_12;
  assign f_u_arrmul24_fa8_12_f_u_arrmul24_and8_12_y0 = f_u_arrmul24_and8_12_y0;
  assign f_u_arrmul24_fa8_12_f_u_arrmul24_fa9_11_y2 = f_u_arrmul24_fa9_11_y2;
  assign f_u_arrmul24_fa8_12_f_u_arrmul24_fa7_12_y4 = f_u_arrmul24_fa7_12_y4;
  assign f_u_arrmul24_fa8_12_y0 = f_u_arrmul24_fa8_12_f_u_arrmul24_and8_12_y0 ^ f_u_arrmul24_fa8_12_f_u_arrmul24_fa9_11_y2;
  assign f_u_arrmul24_fa8_12_y1 = f_u_arrmul24_fa8_12_f_u_arrmul24_and8_12_y0 & f_u_arrmul24_fa8_12_f_u_arrmul24_fa9_11_y2;
  assign f_u_arrmul24_fa8_12_y2 = f_u_arrmul24_fa8_12_y0 ^ f_u_arrmul24_fa8_12_f_u_arrmul24_fa7_12_y4;
  assign f_u_arrmul24_fa8_12_y3 = f_u_arrmul24_fa8_12_y0 & f_u_arrmul24_fa8_12_f_u_arrmul24_fa7_12_y4;
  assign f_u_arrmul24_fa8_12_y4 = f_u_arrmul24_fa8_12_y1 | f_u_arrmul24_fa8_12_y3;
  assign f_u_arrmul24_and9_12_a_9 = a_9;
  assign f_u_arrmul24_and9_12_b_12 = b_12;
  assign f_u_arrmul24_and9_12_y0 = f_u_arrmul24_and9_12_a_9 & f_u_arrmul24_and9_12_b_12;
  assign f_u_arrmul24_fa9_12_f_u_arrmul24_and9_12_y0 = f_u_arrmul24_and9_12_y0;
  assign f_u_arrmul24_fa9_12_f_u_arrmul24_fa10_11_y2 = f_u_arrmul24_fa10_11_y2;
  assign f_u_arrmul24_fa9_12_f_u_arrmul24_fa8_12_y4 = f_u_arrmul24_fa8_12_y4;
  assign f_u_arrmul24_fa9_12_y0 = f_u_arrmul24_fa9_12_f_u_arrmul24_and9_12_y0 ^ f_u_arrmul24_fa9_12_f_u_arrmul24_fa10_11_y2;
  assign f_u_arrmul24_fa9_12_y1 = f_u_arrmul24_fa9_12_f_u_arrmul24_and9_12_y0 & f_u_arrmul24_fa9_12_f_u_arrmul24_fa10_11_y2;
  assign f_u_arrmul24_fa9_12_y2 = f_u_arrmul24_fa9_12_y0 ^ f_u_arrmul24_fa9_12_f_u_arrmul24_fa8_12_y4;
  assign f_u_arrmul24_fa9_12_y3 = f_u_arrmul24_fa9_12_y0 & f_u_arrmul24_fa9_12_f_u_arrmul24_fa8_12_y4;
  assign f_u_arrmul24_fa9_12_y4 = f_u_arrmul24_fa9_12_y1 | f_u_arrmul24_fa9_12_y3;
  assign f_u_arrmul24_and10_12_a_10 = a_10;
  assign f_u_arrmul24_and10_12_b_12 = b_12;
  assign f_u_arrmul24_and10_12_y0 = f_u_arrmul24_and10_12_a_10 & f_u_arrmul24_and10_12_b_12;
  assign f_u_arrmul24_fa10_12_f_u_arrmul24_and10_12_y0 = f_u_arrmul24_and10_12_y0;
  assign f_u_arrmul24_fa10_12_f_u_arrmul24_fa11_11_y2 = f_u_arrmul24_fa11_11_y2;
  assign f_u_arrmul24_fa10_12_f_u_arrmul24_fa9_12_y4 = f_u_arrmul24_fa9_12_y4;
  assign f_u_arrmul24_fa10_12_y0 = f_u_arrmul24_fa10_12_f_u_arrmul24_and10_12_y0 ^ f_u_arrmul24_fa10_12_f_u_arrmul24_fa11_11_y2;
  assign f_u_arrmul24_fa10_12_y1 = f_u_arrmul24_fa10_12_f_u_arrmul24_and10_12_y0 & f_u_arrmul24_fa10_12_f_u_arrmul24_fa11_11_y2;
  assign f_u_arrmul24_fa10_12_y2 = f_u_arrmul24_fa10_12_y0 ^ f_u_arrmul24_fa10_12_f_u_arrmul24_fa9_12_y4;
  assign f_u_arrmul24_fa10_12_y3 = f_u_arrmul24_fa10_12_y0 & f_u_arrmul24_fa10_12_f_u_arrmul24_fa9_12_y4;
  assign f_u_arrmul24_fa10_12_y4 = f_u_arrmul24_fa10_12_y1 | f_u_arrmul24_fa10_12_y3;
  assign f_u_arrmul24_and11_12_a_11 = a_11;
  assign f_u_arrmul24_and11_12_b_12 = b_12;
  assign f_u_arrmul24_and11_12_y0 = f_u_arrmul24_and11_12_a_11 & f_u_arrmul24_and11_12_b_12;
  assign f_u_arrmul24_fa11_12_f_u_arrmul24_and11_12_y0 = f_u_arrmul24_and11_12_y0;
  assign f_u_arrmul24_fa11_12_f_u_arrmul24_fa12_11_y2 = f_u_arrmul24_fa12_11_y2;
  assign f_u_arrmul24_fa11_12_f_u_arrmul24_fa10_12_y4 = f_u_arrmul24_fa10_12_y4;
  assign f_u_arrmul24_fa11_12_y0 = f_u_arrmul24_fa11_12_f_u_arrmul24_and11_12_y0 ^ f_u_arrmul24_fa11_12_f_u_arrmul24_fa12_11_y2;
  assign f_u_arrmul24_fa11_12_y1 = f_u_arrmul24_fa11_12_f_u_arrmul24_and11_12_y0 & f_u_arrmul24_fa11_12_f_u_arrmul24_fa12_11_y2;
  assign f_u_arrmul24_fa11_12_y2 = f_u_arrmul24_fa11_12_y0 ^ f_u_arrmul24_fa11_12_f_u_arrmul24_fa10_12_y4;
  assign f_u_arrmul24_fa11_12_y3 = f_u_arrmul24_fa11_12_y0 & f_u_arrmul24_fa11_12_f_u_arrmul24_fa10_12_y4;
  assign f_u_arrmul24_fa11_12_y4 = f_u_arrmul24_fa11_12_y1 | f_u_arrmul24_fa11_12_y3;
  assign f_u_arrmul24_and12_12_a_12 = a_12;
  assign f_u_arrmul24_and12_12_b_12 = b_12;
  assign f_u_arrmul24_and12_12_y0 = f_u_arrmul24_and12_12_a_12 & f_u_arrmul24_and12_12_b_12;
  assign f_u_arrmul24_fa12_12_f_u_arrmul24_and12_12_y0 = f_u_arrmul24_and12_12_y0;
  assign f_u_arrmul24_fa12_12_f_u_arrmul24_fa13_11_y2 = f_u_arrmul24_fa13_11_y2;
  assign f_u_arrmul24_fa12_12_f_u_arrmul24_fa11_12_y4 = f_u_arrmul24_fa11_12_y4;
  assign f_u_arrmul24_fa12_12_y0 = f_u_arrmul24_fa12_12_f_u_arrmul24_and12_12_y0 ^ f_u_arrmul24_fa12_12_f_u_arrmul24_fa13_11_y2;
  assign f_u_arrmul24_fa12_12_y1 = f_u_arrmul24_fa12_12_f_u_arrmul24_and12_12_y0 & f_u_arrmul24_fa12_12_f_u_arrmul24_fa13_11_y2;
  assign f_u_arrmul24_fa12_12_y2 = f_u_arrmul24_fa12_12_y0 ^ f_u_arrmul24_fa12_12_f_u_arrmul24_fa11_12_y4;
  assign f_u_arrmul24_fa12_12_y3 = f_u_arrmul24_fa12_12_y0 & f_u_arrmul24_fa12_12_f_u_arrmul24_fa11_12_y4;
  assign f_u_arrmul24_fa12_12_y4 = f_u_arrmul24_fa12_12_y1 | f_u_arrmul24_fa12_12_y3;
  assign f_u_arrmul24_and13_12_a_13 = a_13;
  assign f_u_arrmul24_and13_12_b_12 = b_12;
  assign f_u_arrmul24_and13_12_y0 = f_u_arrmul24_and13_12_a_13 & f_u_arrmul24_and13_12_b_12;
  assign f_u_arrmul24_fa13_12_f_u_arrmul24_and13_12_y0 = f_u_arrmul24_and13_12_y0;
  assign f_u_arrmul24_fa13_12_f_u_arrmul24_fa14_11_y2 = f_u_arrmul24_fa14_11_y2;
  assign f_u_arrmul24_fa13_12_f_u_arrmul24_fa12_12_y4 = f_u_arrmul24_fa12_12_y4;
  assign f_u_arrmul24_fa13_12_y0 = f_u_arrmul24_fa13_12_f_u_arrmul24_and13_12_y0 ^ f_u_arrmul24_fa13_12_f_u_arrmul24_fa14_11_y2;
  assign f_u_arrmul24_fa13_12_y1 = f_u_arrmul24_fa13_12_f_u_arrmul24_and13_12_y0 & f_u_arrmul24_fa13_12_f_u_arrmul24_fa14_11_y2;
  assign f_u_arrmul24_fa13_12_y2 = f_u_arrmul24_fa13_12_y0 ^ f_u_arrmul24_fa13_12_f_u_arrmul24_fa12_12_y4;
  assign f_u_arrmul24_fa13_12_y3 = f_u_arrmul24_fa13_12_y0 & f_u_arrmul24_fa13_12_f_u_arrmul24_fa12_12_y4;
  assign f_u_arrmul24_fa13_12_y4 = f_u_arrmul24_fa13_12_y1 | f_u_arrmul24_fa13_12_y3;
  assign f_u_arrmul24_and14_12_a_14 = a_14;
  assign f_u_arrmul24_and14_12_b_12 = b_12;
  assign f_u_arrmul24_and14_12_y0 = f_u_arrmul24_and14_12_a_14 & f_u_arrmul24_and14_12_b_12;
  assign f_u_arrmul24_fa14_12_f_u_arrmul24_and14_12_y0 = f_u_arrmul24_and14_12_y0;
  assign f_u_arrmul24_fa14_12_f_u_arrmul24_fa15_11_y2 = f_u_arrmul24_fa15_11_y2;
  assign f_u_arrmul24_fa14_12_f_u_arrmul24_fa13_12_y4 = f_u_arrmul24_fa13_12_y4;
  assign f_u_arrmul24_fa14_12_y0 = f_u_arrmul24_fa14_12_f_u_arrmul24_and14_12_y0 ^ f_u_arrmul24_fa14_12_f_u_arrmul24_fa15_11_y2;
  assign f_u_arrmul24_fa14_12_y1 = f_u_arrmul24_fa14_12_f_u_arrmul24_and14_12_y0 & f_u_arrmul24_fa14_12_f_u_arrmul24_fa15_11_y2;
  assign f_u_arrmul24_fa14_12_y2 = f_u_arrmul24_fa14_12_y0 ^ f_u_arrmul24_fa14_12_f_u_arrmul24_fa13_12_y4;
  assign f_u_arrmul24_fa14_12_y3 = f_u_arrmul24_fa14_12_y0 & f_u_arrmul24_fa14_12_f_u_arrmul24_fa13_12_y4;
  assign f_u_arrmul24_fa14_12_y4 = f_u_arrmul24_fa14_12_y1 | f_u_arrmul24_fa14_12_y3;
  assign f_u_arrmul24_and15_12_a_15 = a_15;
  assign f_u_arrmul24_and15_12_b_12 = b_12;
  assign f_u_arrmul24_and15_12_y0 = f_u_arrmul24_and15_12_a_15 & f_u_arrmul24_and15_12_b_12;
  assign f_u_arrmul24_fa15_12_f_u_arrmul24_and15_12_y0 = f_u_arrmul24_and15_12_y0;
  assign f_u_arrmul24_fa15_12_f_u_arrmul24_fa16_11_y2 = f_u_arrmul24_fa16_11_y2;
  assign f_u_arrmul24_fa15_12_f_u_arrmul24_fa14_12_y4 = f_u_arrmul24_fa14_12_y4;
  assign f_u_arrmul24_fa15_12_y0 = f_u_arrmul24_fa15_12_f_u_arrmul24_and15_12_y0 ^ f_u_arrmul24_fa15_12_f_u_arrmul24_fa16_11_y2;
  assign f_u_arrmul24_fa15_12_y1 = f_u_arrmul24_fa15_12_f_u_arrmul24_and15_12_y0 & f_u_arrmul24_fa15_12_f_u_arrmul24_fa16_11_y2;
  assign f_u_arrmul24_fa15_12_y2 = f_u_arrmul24_fa15_12_y0 ^ f_u_arrmul24_fa15_12_f_u_arrmul24_fa14_12_y4;
  assign f_u_arrmul24_fa15_12_y3 = f_u_arrmul24_fa15_12_y0 & f_u_arrmul24_fa15_12_f_u_arrmul24_fa14_12_y4;
  assign f_u_arrmul24_fa15_12_y4 = f_u_arrmul24_fa15_12_y1 | f_u_arrmul24_fa15_12_y3;
  assign f_u_arrmul24_and16_12_a_16 = a_16;
  assign f_u_arrmul24_and16_12_b_12 = b_12;
  assign f_u_arrmul24_and16_12_y0 = f_u_arrmul24_and16_12_a_16 & f_u_arrmul24_and16_12_b_12;
  assign f_u_arrmul24_fa16_12_f_u_arrmul24_and16_12_y0 = f_u_arrmul24_and16_12_y0;
  assign f_u_arrmul24_fa16_12_f_u_arrmul24_fa17_11_y2 = f_u_arrmul24_fa17_11_y2;
  assign f_u_arrmul24_fa16_12_f_u_arrmul24_fa15_12_y4 = f_u_arrmul24_fa15_12_y4;
  assign f_u_arrmul24_fa16_12_y0 = f_u_arrmul24_fa16_12_f_u_arrmul24_and16_12_y0 ^ f_u_arrmul24_fa16_12_f_u_arrmul24_fa17_11_y2;
  assign f_u_arrmul24_fa16_12_y1 = f_u_arrmul24_fa16_12_f_u_arrmul24_and16_12_y0 & f_u_arrmul24_fa16_12_f_u_arrmul24_fa17_11_y2;
  assign f_u_arrmul24_fa16_12_y2 = f_u_arrmul24_fa16_12_y0 ^ f_u_arrmul24_fa16_12_f_u_arrmul24_fa15_12_y4;
  assign f_u_arrmul24_fa16_12_y3 = f_u_arrmul24_fa16_12_y0 & f_u_arrmul24_fa16_12_f_u_arrmul24_fa15_12_y4;
  assign f_u_arrmul24_fa16_12_y4 = f_u_arrmul24_fa16_12_y1 | f_u_arrmul24_fa16_12_y3;
  assign f_u_arrmul24_and17_12_a_17 = a_17;
  assign f_u_arrmul24_and17_12_b_12 = b_12;
  assign f_u_arrmul24_and17_12_y0 = f_u_arrmul24_and17_12_a_17 & f_u_arrmul24_and17_12_b_12;
  assign f_u_arrmul24_fa17_12_f_u_arrmul24_and17_12_y0 = f_u_arrmul24_and17_12_y0;
  assign f_u_arrmul24_fa17_12_f_u_arrmul24_fa18_11_y2 = f_u_arrmul24_fa18_11_y2;
  assign f_u_arrmul24_fa17_12_f_u_arrmul24_fa16_12_y4 = f_u_arrmul24_fa16_12_y4;
  assign f_u_arrmul24_fa17_12_y0 = f_u_arrmul24_fa17_12_f_u_arrmul24_and17_12_y0 ^ f_u_arrmul24_fa17_12_f_u_arrmul24_fa18_11_y2;
  assign f_u_arrmul24_fa17_12_y1 = f_u_arrmul24_fa17_12_f_u_arrmul24_and17_12_y0 & f_u_arrmul24_fa17_12_f_u_arrmul24_fa18_11_y2;
  assign f_u_arrmul24_fa17_12_y2 = f_u_arrmul24_fa17_12_y0 ^ f_u_arrmul24_fa17_12_f_u_arrmul24_fa16_12_y4;
  assign f_u_arrmul24_fa17_12_y3 = f_u_arrmul24_fa17_12_y0 & f_u_arrmul24_fa17_12_f_u_arrmul24_fa16_12_y4;
  assign f_u_arrmul24_fa17_12_y4 = f_u_arrmul24_fa17_12_y1 | f_u_arrmul24_fa17_12_y3;
  assign f_u_arrmul24_and18_12_a_18 = a_18;
  assign f_u_arrmul24_and18_12_b_12 = b_12;
  assign f_u_arrmul24_and18_12_y0 = f_u_arrmul24_and18_12_a_18 & f_u_arrmul24_and18_12_b_12;
  assign f_u_arrmul24_fa18_12_f_u_arrmul24_and18_12_y0 = f_u_arrmul24_and18_12_y0;
  assign f_u_arrmul24_fa18_12_f_u_arrmul24_fa19_11_y2 = f_u_arrmul24_fa19_11_y2;
  assign f_u_arrmul24_fa18_12_f_u_arrmul24_fa17_12_y4 = f_u_arrmul24_fa17_12_y4;
  assign f_u_arrmul24_fa18_12_y0 = f_u_arrmul24_fa18_12_f_u_arrmul24_and18_12_y0 ^ f_u_arrmul24_fa18_12_f_u_arrmul24_fa19_11_y2;
  assign f_u_arrmul24_fa18_12_y1 = f_u_arrmul24_fa18_12_f_u_arrmul24_and18_12_y0 & f_u_arrmul24_fa18_12_f_u_arrmul24_fa19_11_y2;
  assign f_u_arrmul24_fa18_12_y2 = f_u_arrmul24_fa18_12_y0 ^ f_u_arrmul24_fa18_12_f_u_arrmul24_fa17_12_y4;
  assign f_u_arrmul24_fa18_12_y3 = f_u_arrmul24_fa18_12_y0 & f_u_arrmul24_fa18_12_f_u_arrmul24_fa17_12_y4;
  assign f_u_arrmul24_fa18_12_y4 = f_u_arrmul24_fa18_12_y1 | f_u_arrmul24_fa18_12_y3;
  assign f_u_arrmul24_and19_12_a_19 = a_19;
  assign f_u_arrmul24_and19_12_b_12 = b_12;
  assign f_u_arrmul24_and19_12_y0 = f_u_arrmul24_and19_12_a_19 & f_u_arrmul24_and19_12_b_12;
  assign f_u_arrmul24_fa19_12_f_u_arrmul24_and19_12_y0 = f_u_arrmul24_and19_12_y0;
  assign f_u_arrmul24_fa19_12_f_u_arrmul24_fa20_11_y2 = f_u_arrmul24_fa20_11_y2;
  assign f_u_arrmul24_fa19_12_f_u_arrmul24_fa18_12_y4 = f_u_arrmul24_fa18_12_y4;
  assign f_u_arrmul24_fa19_12_y0 = f_u_arrmul24_fa19_12_f_u_arrmul24_and19_12_y0 ^ f_u_arrmul24_fa19_12_f_u_arrmul24_fa20_11_y2;
  assign f_u_arrmul24_fa19_12_y1 = f_u_arrmul24_fa19_12_f_u_arrmul24_and19_12_y0 & f_u_arrmul24_fa19_12_f_u_arrmul24_fa20_11_y2;
  assign f_u_arrmul24_fa19_12_y2 = f_u_arrmul24_fa19_12_y0 ^ f_u_arrmul24_fa19_12_f_u_arrmul24_fa18_12_y4;
  assign f_u_arrmul24_fa19_12_y3 = f_u_arrmul24_fa19_12_y0 & f_u_arrmul24_fa19_12_f_u_arrmul24_fa18_12_y4;
  assign f_u_arrmul24_fa19_12_y4 = f_u_arrmul24_fa19_12_y1 | f_u_arrmul24_fa19_12_y3;
  assign f_u_arrmul24_and20_12_a_20 = a_20;
  assign f_u_arrmul24_and20_12_b_12 = b_12;
  assign f_u_arrmul24_and20_12_y0 = f_u_arrmul24_and20_12_a_20 & f_u_arrmul24_and20_12_b_12;
  assign f_u_arrmul24_fa20_12_f_u_arrmul24_and20_12_y0 = f_u_arrmul24_and20_12_y0;
  assign f_u_arrmul24_fa20_12_f_u_arrmul24_fa21_11_y2 = f_u_arrmul24_fa21_11_y2;
  assign f_u_arrmul24_fa20_12_f_u_arrmul24_fa19_12_y4 = f_u_arrmul24_fa19_12_y4;
  assign f_u_arrmul24_fa20_12_y0 = f_u_arrmul24_fa20_12_f_u_arrmul24_and20_12_y0 ^ f_u_arrmul24_fa20_12_f_u_arrmul24_fa21_11_y2;
  assign f_u_arrmul24_fa20_12_y1 = f_u_arrmul24_fa20_12_f_u_arrmul24_and20_12_y0 & f_u_arrmul24_fa20_12_f_u_arrmul24_fa21_11_y2;
  assign f_u_arrmul24_fa20_12_y2 = f_u_arrmul24_fa20_12_y0 ^ f_u_arrmul24_fa20_12_f_u_arrmul24_fa19_12_y4;
  assign f_u_arrmul24_fa20_12_y3 = f_u_arrmul24_fa20_12_y0 & f_u_arrmul24_fa20_12_f_u_arrmul24_fa19_12_y4;
  assign f_u_arrmul24_fa20_12_y4 = f_u_arrmul24_fa20_12_y1 | f_u_arrmul24_fa20_12_y3;
  assign f_u_arrmul24_and21_12_a_21 = a_21;
  assign f_u_arrmul24_and21_12_b_12 = b_12;
  assign f_u_arrmul24_and21_12_y0 = f_u_arrmul24_and21_12_a_21 & f_u_arrmul24_and21_12_b_12;
  assign f_u_arrmul24_fa21_12_f_u_arrmul24_and21_12_y0 = f_u_arrmul24_and21_12_y0;
  assign f_u_arrmul24_fa21_12_f_u_arrmul24_fa22_11_y2 = f_u_arrmul24_fa22_11_y2;
  assign f_u_arrmul24_fa21_12_f_u_arrmul24_fa20_12_y4 = f_u_arrmul24_fa20_12_y4;
  assign f_u_arrmul24_fa21_12_y0 = f_u_arrmul24_fa21_12_f_u_arrmul24_and21_12_y0 ^ f_u_arrmul24_fa21_12_f_u_arrmul24_fa22_11_y2;
  assign f_u_arrmul24_fa21_12_y1 = f_u_arrmul24_fa21_12_f_u_arrmul24_and21_12_y0 & f_u_arrmul24_fa21_12_f_u_arrmul24_fa22_11_y2;
  assign f_u_arrmul24_fa21_12_y2 = f_u_arrmul24_fa21_12_y0 ^ f_u_arrmul24_fa21_12_f_u_arrmul24_fa20_12_y4;
  assign f_u_arrmul24_fa21_12_y3 = f_u_arrmul24_fa21_12_y0 & f_u_arrmul24_fa21_12_f_u_arrmul24_fa20_12_y4;
  assign f_u_arrmul24_fa21_12_y4 = f_u_arrmul24_fa21_12_y1 | f_u_arrmul24_fa21_12_y3;
  assign f_u_arrmul24_and22_12_a_22 = a_22;
  assign f_u_arrmul24_and22_12_b_12 = b_12;
  assign f_u_arrmul24_and22_12_y0 = f_u_arrmul24_and22_12_a_22 & f_u_arrmul24_and22_12_b_12;
  assign f_u_arrmul24_fa22_12_f_u_arrmul24_and22_12_y0 = f_u_arrmul24_and22_12_y0;
  assign f_u_arrmul24_fa22_12_f_u_arrmul24_fa23_11_y2 = f_u_arrmul24_fa23_11_y2;
  assign f_u_arrmul24_fa22_12_f_u_arrmul24_fa21_12_y4 = f_u_arrmul24_fa21_12_y4;
  assign f_u_arrmul24_fa22_12_y0 = f_u_arrmul24_fa22_12_f_u_arrmul24_and22_12_y0 ^ f_u_arrmul24_fa22_12_f_u_arrmul24_fa23_11_y2;
  assign f_u_arrmul24_fa22_12_y1 = f_u_arrmul24_fa22_12_f_u_arrmul24_and22_12_y0 & f_u_arrmul24_fa22_12_f_u_arrmul24_fa23_11_y2;
  assign f_u_arrmul24_fa22_12_y2 = f_u_arrmul24_fa22_12_y0 ^ f_u_arrmul24_fa22_12_f_u_arrmul24_fa21_12_y4;
  assign f_u_arrmul24_fa22_12_y3 = f_u_arrmul24_fa22_12_y0 & f_u_arrmul24_fa22_12_f_u_arrmul24_fa21_12_y4;
  assign f_u_arrmul24_fa22_12_y4 = f_u_arrmul24_fa22_12_y1 | f_u_arrmul24_fa22_12_y3;
  assign f_u_arrmul24_and23_12_a_23 = a_23;
  assign f_u_arrmul24_and23_12_b_12 = b_12;
  assign f_u_arrmul24_and23_12_y0 = f_u_arrmul24_and23_12_a_23 & f_u_arrmul24_and23_12_b_12;
  assign f_u_arrmul24_fa23_12_f_u_arrmul24_and23_12_y0 = f_u_arrmul24_and23_12_y0;
  assign f_u_arrmul24_fa23_12_f_u_arrmul24_fa23_11_y4 = f_u_arrmul24_fa23_11_y4;
  assign f_u_arrmul24_fa23_12_f_u_arrmul24_fa22_12_y4 = f_u_arrmul24_fa22_12_y4;
  assign f_u_arrmul24_fa23_12_y0 = f_u_arrmul24_fa23_12_f_u_arrmul24_and23_12_y0 ^ f_u_arrmul24_fa23_12_f_u_arrmul24_fa23_11_y4;
  assign f_u_arrmul24_fa23_12_y1 = f_u_arrmul24_fa23_12_f_u_arrmul24_and23_12_y0 & f_u_arrmul24_fa23_12_f_u_arrmul24_fa23_11_y4;
  assign f_u_arrmul24_fa23_12_y2 = f_u_arrmul24_fa23_12_y0 ^ f_u_arrmul24_fa23_12_f_u_arrmul24_fa22_12_y4;
  assign f_u_arrmul24_fa23_12_y3 = f_u_arrmul24_fa23_12_y0 & f_u_arrmul24_fa23_12_f_u_arrmul24_fa22_12_y4;
  assign f_u_arrmul24_fa23_12_y4 = f_u_arrmul24_fa23_12_y1 | f_u_arrmul24_fa23_12_y3;
  assign f_u_arrmul24_and0_13_a_0 = a_0;
  assign f_u_arrmul24_and0_13_b_13 = b_13;
  assign f_u_arrmul24_and0_13_y0 = f_u_arrmul24_and0_13_a_0 & f_u_arrmul24_and0_13_b_13;
  assign f_u_arrmul24_ha0_13_f_u_arrmul24_and0_13_y0 = f_u_arrmul24_and0_13_y0;
  assign f_u_arrmul24_ha0_13_f_u_arrmul24_fa1_12_y2 = f_u_arrmul24_fa1_12_y2;
  assign f_u_arrmul24_ha0_13_y0 = f_u_arrmul24_ha0_13_f_u_arrmul24_and0_13_y0 ^ f_u_arrmul24_ha0_13_f_u_arrmul24_fa1_12_y2;
  assign f_u_arrmul24_ha0_13_y1 = f_u_arrmul24_ha0_13_f_u_arrmul24_and0_13_y0 & f_u_arrmul24_ha0_13_f_u_arrmul24_fa1_12_y2;
  assign f_u_arrmul24_and1_13_a_1 = a_1;
  assign f_u_arrmul24_and1_13_b_13 = b_13;
  assign f_u_arrmul24_and1_13_y0 = f_u_arrmul24_and1_13_a_1 & f_u_arrmul24_and1_13_b_13;
  assign f_u_arrmul24_fa1_13_f_u_arrmul24_and1_13_y0 = f_u_arrmul24_and1_13_y0;
  assign f_u_arrmul24_fa1_13_f_u_arrmul24_fa2_12_y2 = f_u_arrmul24_fa2_12_y2;
  assign f_u_arrmul24_fa1_13_f_u_arrmul24_ha0_13_y1 = f_u_arrmul24_ha0_13_y1;
  assign f_u_arrmul24_fa1_13_y0 = f_u_arrmul24_fa1_13_f_u_arrmul24_and1_13_y0 ^ f_u_arrmul24_fa1_13_f_u_arrmul24_fa2_12_y2;
  assign f_u_arrmul24_fa1_13_y1 = f_u_arrmul24_fa1_13_f_u_arrmul24_and1_13_y0 & f_u_arrmul24_fa1_13_f_u_arrmul24_fa2_12_y2;
  assign f_u_arrmul24_fa1_13_y2 = f_u_arrmul24_fa1_13_y0 ^ f_u_arrmul24_fa1_13_f_u_arrmul24_ha0_13_y1;
  assign f_u_arrmul24_fa1_13_y3 = f_u_arrmul24_fa1_13_y0 & f_u_arrmul24_fa1_13_f_u_arrmul24_ha0_13_y1;
  assign f_u_arrmul24_fa1_13_y4 = f_u_arrmul24_fa1_13_y1 | f_u_arrmul24_fa1_13_y3;
  assign f_u_arrmul24_and2_13_a_2 = a_2;
  assign f_u_arrmul24_and2_13_b_13 = b_13;
  assign f_u_arrmul24_and2_13_y0 = f_u_arrmul24_and2_13_a_2 & f_u_arrmul24_and2_13_b_13;
  assign f_u_arrmul24_fa2_13_f_u_arrmul24_and2_13_y0 = f_u_arrmul24_and2_13_y0;
  assign f_u_arrmul24_fa2_13_f_u_arrmul24_fa3_12_y2 = f_u_arrmul24_fa3_12_y2;
  assign f_u_arrmul24_fa2_13_f_u_arrmul24_fa1_13_y4 = f_u_arrmul24_fa1_13_y4;
  assign f_u_arrmul24_fa2_13_y0 = f_u_arrmul24_fa2_13_f_u_arrmul24_and2_13_y0 ^ f_u_arrmul24_fa2_13_f_u_arrmul24_fa3_12_y2;
  assign f_u_arrmul24_fa2_13_y1 = f_u_arrmul24_fa2_13_f_u_arrmul24_and2_13_y0 & f_u_arrmul24_fa2_13_f_u_arrmul24_fa3_12_y2;
  assign f_u_arrmul24_fa2_13_y2 = f_u_arrmul24_fa2_13_y0 ^ f_u_arrmul24_fa2_13_f_u_arrmul24_fa1_13_y4;
  assign f_u_arrmul24_fa2_13_y3 = f_u_arrmul24_fa2_13_y0 & f_u_arrmul24_fa2_13_f_u_arrmul24_fa1_13_y4;
  assign f_u_arrmul24_fa2_13_y4 = f_u_arrmul24_fa2_13_y1 | f_u_arrmul24_fa2_13_y3;
  assign f_u_arrmul24_and3_13_a_3 = a_3;
  assign f_u_arrmul24_and3_13_b_13 = b_13;
  assign f_u_arrmul24_and3_13_y0 = f_u_arrmul24_and3_13_a_3 & f_u_arrmul24_and3_13_b_13;
  assign f_u_arrmul24_fa3_13_f_u_arrmul24_and3_13_y0 = f_u_arrmul24_and3_13_y0;
  assign f_u_arrmul24_fa3_13_f_u_arrmul24_fa4_12_y2 = f_u_arrmul24_fa4_12_y2;
  assign f_u_arrmul24_fa3_13_f_u_arrmul24_fa2_13_y4 = f_u_arrmul24_fa2_13_y4;
  assign f_u_arrmul24_fa3_13_y0 = f_u_arrmul24_fa3_13_f_u_arrmul24_and3_13_y0 ^ f_u_arrmul24_fa3_13_f_u_arrmul24_fa4_12_y2;
  assign f_u_arrmul24_fa3_13_y1 = f_u_arrmul24_fa3_13_f_u_arrmul24_and3_13_y0 & f_u_arrmul24_fa3_13_f_u_arrmul24_fa4_12_y2;
  assign f_u_arrmul24_fa3_13_y2 = f_u_arrmul24_fa3_13_y0 ^ f_u_arrmul24_fa3_13_f_u_arrmul24_fa2_13_y4;
  assign f_u_arrmul24_fa3_13_y3 = f_u_arrmul24_fa3_13_y0 & f_u_arrmul24_fa3_13_f_u_arrmul24_fa2_13_y4;
  assign f_u_arrmul24_fa3_13_y4 = f_u_arrmul24_fa3_13_y1 | f_u_arrmul24_fa3_13_y3;
  assign f_u_arrmul24_and4_13_a_4 = a_4;
  assign f_u_arrmul24_and4_13_b_13 = b_13;
  assign f_u_arrmul24_and4_13_y0 = f_u_arrmul24_and4_13_a_4 & f_u_arrmul24_and4_13_b_13;
  assign f_u_arrmul24_fa4_13_f_u_arrmul24_and4_13_y0 = f_u_arrmul24_and4_13_y0;
  assign f_u_arrmul24_fa4_13_f_u_arrmul24_fa5_12_y2 = f_u_arrmul24_fa5_12_y2;
  assign f_u_arrmul24_fa4_13_f_u_arrmul24_fa3_13_y4 = f_u_arrmul24_fa3_13_y4;
  assign f_u_arrmul24_fa4_13_y0 = f_u_arrmul24_fa4_13_f_u_arrmul24_and4_13_y0 ^ f_u_arrmul24_fa4_13_f_u_arrmul24_fa5_12_y2;
  assign f_u_arrmul24_fa4_13_y1 = f_u_arrmul24_fa4_13_f_u_arrmul24_and4_13_y0 & f_u_arrmul24_fa4_13_f_u_arrmul24_fa5_12_y2;
  assign f_u_arrmul24_fa4_13_y2 = f_u_arrmul24_fa4_13_y0 ^ f_u_arrmul24_fa4_13_f_u_arrmul24_fa3_13_y4;
  assign f_u_arrmul24_fa4_13_y3 = f_u_arrmul24_fa4_13_y0 & f_u_arrmul24_fa4_13_f_u_arrmul24_fa3_13_y4;
  assign f_u_arrmul24_fa4_13_y4 = f_u_arrmul24_fa4_13_y1 | f_u_arrmul24_fa4_13_y3;
  assign f_u_arrmul24_and5_13_a_5 = a_5;
  assign f_u_arrmul24_and5_13_b_13 = b_13;
  assign f_u_arrmul24_and5_13_y0 = f_u_arrmul24_and5_13_a_5 & f_u_arrmul24_and5_13_b_13;
  assign f_u_arrmul24_fa5_13_f_u_arrmul24_and5_13_y0 = f_u_arrmul24_and5_13_y0;
  assign f_u_arrmul24_fa5_13_f_u_arrmul24_fa6_12_y2 = f_u_arrmul24_fa6_12_y2;
  assign f_u_arrmul24_fa5_13_f_u_arrmul24_fa4_13_y4 = f_u_arrmul24_fa4_13_y4;
  assign f_u_arrmul24_fa5_13_y0 = f_u_arrmul24_fa5_13_f_u_arrmul24_and5_13_y0 ^ f_u_arrmul24_fa5_13_f_u_arrmul24_fa6_12_y2;
  assign f_u_arrmul24_fa5_13_y1 = f_u_arrmul24_fa5_13_f_u_arrmul24_and5_13_y0 & f_u_arrmul24_fa5_13_f_u_arrmul24_fa6_12_y2;
  assign f_u_arrmul24_fa5_13_y2 = f_u_arrmul24_fa5_13_y0 ^ f_u_arrmul24_fa5_13_f_u_arrmul24_fa4_13_y4;
  assign f_u_arrmul24_fa5_13_y3 = f_u_arrmul24_fa5_13_y0 & f_u_arrmul24_fa5_13_f_u_arrmul24_fa4_13_y4;
  assign f_u_arrmul24_fa5_13_y4 = f_u_arrmul24_fa5_13_y1 | f_u_arrmul24_fa5_13_y3;
  assign f_u_arrmul24_and6_13_a_6 = a_6;
  assign f_u_arrmul24_and6_13_b_13 = b_13;
  assign f_u_arrmul24_and6_13_y0 = f_u_arrmul24_and6_13_a_6 & f_u_arrmul24_and6_13_b_13;
  assign f_u_arrmul24_fa6_13_f_u_arrmul24_and6_13_y0 = f_u_arrmul24_and6_13_y0;
  assign f_u_arrmul24_fa6_13_f_u_arrmul24_fa7_12_y2 = f_u_arrmul24_fa7_12_y2;
  assign f_u_arrmul24_fa6_13_f_u_arrmul24_fa5_13_y4 = f_u_arrmul24_fa5_13_y4;
  assign f_u_arrmul24_fa6_13_y0 = f_u_arrmul24_fa6_13_f_u_arrmul24_and6_13_y0 ^ f_u_arrmul24_fa6_13_f_u_arrmul24_fa7_12_y2;
  assign f_u_arrmul24_fa6_13_y1 = f_u_arrmul24_fa6_13_f_u_arrmul24_and6_13_y0 & f_u_arrmul24_fa6_13_f_u_arrmul24_fa7_12_y2;
  assign f_u_arrmul24_fa6_13_y2 = f_u_arrmul24_fa6_13_y0 ^ f_u_arrmul24_fa6_13_f_u_arrmul24_fa5_13_y4;
  assign f_u_arrmul24_fa6_13_y3 = f_u_arrmul24_fa6_13_y0 & f_u_arrmul24_fa6_13_f_u_arrmul24_fa5_13_y4;
  assign f_u_arrmul24_fa6_13_y4 = f_u_arrmul24_fa6_13_y1 | f_u_arrmul24_fa6_13_y3;
  assign f_u_arrmul24_and7_13_a_7 = a_7;
  assign f_u_arrmul24_and7_13_b_13 = b_13;
  assign f_u_arrmul24_and7_13_y0 = f_u_arrmul24_and7_13_a_7 & f_u_arrmul24_and7_13_b_13;
  assign f_u_arrmul24_fa7_13_f_u_arrmul24_and7_13_y0 = f_u_arrmul24_and7_13_y0;
  assign f_u_arrmul24_fa7_13_f_u_arrmul24_fa8_12_y2 = f_u_arrmul24_fa8_12_y2;
  assign f_u_arrmul24_fa7_13_f_u_arrmul24_fa6_13_y4 = f_u_arrmul24_fa6_13_y4;
  assign f_u_arrmul24_fa7_13_y0 = f_u_arrmul24_fa7_13_f_u_arrmul24_and7_13_y0 ^ f_u_arrmul24_fa7_13_f_u_arrmul24_fa8_12_y2;
  assign f_u_arrmul24_fa7_13_y1 = f_u_arrmul24_fa7_13_f_u_arrmul24_and7_13_y0 & f_u_arrmul24_fa7_13_f_u_arrmul24_fa8_12_y2;
  assign f_u_arrmul24_fa7_13_y2 = f_u_arrmul24_fa7_13_y0 ^ f_u_arrmul24_fa7_13_f_u_arrmul24_fa6_13_y4;
  assign f_u_arrmul24_fa7_13_y3 = f_u_arrmul24_fa7_13_y0 & f_u_arrmul24_fa7_13_f_u_arrmul24_fa6_13_y4;
  assign f_u_arrmul24_fa7_13_y4 = f_u_arrmul24_fa7_13_y1 | f_u_arrmul24_fa7_13_y3;
  assign f_u_arrmul24_and8_13_a_8 = a_8;
  assign f_u_arrmul24_and8_13_b_13 = b_13;
  assign f_u_arrmul24_and8_13_y0 = f_u_arrmul24_and8_13_a_8 & f_u_arrmul24_and8_13_b_13;
  assign f_u_arrmul24_fa8_13_f_u_arrmul24_and8_13_y0 = f_u_arrmul24_and8_13_y0;
  assign f_u_arrmul24_fa8_13_f_u_arrmul24_fa9_12_y2 = f_u_arrmul24_fa9_12_y2;
  assign f_u_arrmul24_fa8_13_f_u_arrmul24_fa7_13_y4 = f_u_arrmul24_fa7_13_y4;
  assign f_u_arrmul24_fa8_13_y0 = f_u_arrmul24_fa8_13_f_u_arrmul24_and8_13_y0 ^ f_u_arrmul24_fa8_13_f_u_arrmul24_fa9_12_y2;
  assign f_u_arrmul24_fa8_13_y1 = f_u_arrmul24_fa8_13_f_u_arrmul24_and8_13_y0 & f_u_arrmul24_fa8_13_f_u_arrmul24_fa9_12_y2;
  assign f_u_arrmul24_fa8_13_y2 = f_u_arrmul24_fa8_13_y0 ^ f_u_arrmul24_fa8_13_f_u_arrmul24_fa7_13_y4;
  assign f_u_arrmul24_fa8_13_y3 = f_u_arrmul24_fa8_13_y0 & f_u_arrmul24_fa8_13_f_u_arrmul24_fa7_13_y4;
  assign f_u_arrmul24_fa8_13_y4 = f_u_arrmul24_fa8_13_y1 | f_u_arrmul24_fa8_13_y3;
  assign f_u_arrmul24_and9_13_a_9 = a_9;
  assign f_u_arrmul24_and9_13_b_13 = b_13;
  assign f_u_arrmul24_and9_13_y0 = f_u_arrmul24_and9_13_a_9 & f_u_arrmul24_and9_13_b_13;
  assign f_u_arrmul24_fa9_13_f_u_arrmul24_and9_13_y0 = f_u_arrmul24_and9_13_y0;
  assign f_u_arrmul24_fa9_13_f_u_arrmul24_fa10_12_y2 = f_u_arrmul24_fa10_12_y2;
  assign f_u_arrmul24_fa9_13_f_u_arrmul24_fa8_13_y4 = f_u_arrmul24_fa8_13_y4;
  assign f_u_arrmul24_fa9_13_y0 = f_u_arrmul24_fa9_13_f_u_arrmul24_and9_13_y0 ^ f_u_arrmul24_fa9_13_f_u_arrmul24_fa10_12_y2;
  assign f_u_arrmul24_fa9_13_y1 = f_u_arrmul24_fa9_13_f_u_arrmul24_and9_13_y0 & f_u_arrmul24_fa9_13_f_u_arrmul24_fa10_12_y2;
  assign f_u_arrmul24_fa9_13_y2 = f_u_arrmul24_fa9_13_y0 ^ f_u_arrmul24_fa9_13_f_u_arrmul24_fa8_13_y4;
  assign f_u_arrmul24_fa9_13_y3 = f_u_arrmul24_fa9_13_y0 & f_u_arrmul24_fa9_13_f_u_arrmul24_fa8_13_y4;
  assign f_u_arrmul24_fa9_13_y4 = f_u_arrmul24_fa9_13_y1 | f_u_arrmul24_fa9_13_y3;
  assign f_u_arrmul24_and10_13_a_10 = a_10;
  assign f_u_arrmul24_and10_13_b_13 = b_13;
  assign f_u_arrmul24_and10_13_y0 = f_u_arrmul24_and10_13_a_10 & f_u_arrmul24_and10_13_b_13;
  assign f_u_arrmul24_fa10_13_f_u_arrmul24_and10_13_y0 = f_u_arrmul24_and10_13_y0;
  assign f_u_arrmul24_fa10_13_f_u_arrmul24_fa11_12_y2 = f_u_arrmul24_fa11_12_y2;
  assign f_u_arrmul24_fa10_13_f_u_arrmul24_fa9_13_y4 = f_u_arrmul24_fa9_13_y4;
  assign f_u_arrmul24_fa10_13_y0 = f_u_arrmul24_fa10_13_f_u_arrmul24_and10_13_y0 ^ f_u_arrmul24_fa10_13_f_u_arrmul24_fa11_12_y2;
  assign f_u_arrmul24_fa10_13_y1 = f_u_arrmul24_fa10_13_f_u_arrmul24_and10_13_y0 & f_u_arrmul24_fa10_13_f_u_arrmul24_fa11_12_y2;
  assign f_u_arrmul24_fa10_13_y2 = f_u_arrmul24_fa10_13_y0 ^ f_u_arrmul24_fa10_13_f_u_arrmul24_fa9_13_y4;
  assign f_u_arrmul24_fa10_13_y3 = f_u_arrmul24_fa10_13_y0 & f_u_arrmul24_fa10_13_f_u_arrmul24_fa9_13_y4;
  assign f_u_arrmul24_fa10_13_y4 = f_u_arrmul24_fa10_13_y1 | f_u_arrmul24_fa10_13_y3;
  assign f_u_arrmul24_and11_13_a_11 = a_11;
  assign f_u_arrmul24_and11_13_b_13 = b_13;
  assign f_u_arrmul24_and11_13_y0 = f_u_arrmul24_and11_13_a_11 & f_u_arrmul24_and11_13_b_13;
  assign f_u_arrmul24_fa11_13_f_u_arrmul24_and11_13_y0 = f_u_arrmul24_and11_13_y0;
  assign f_u_arrmul24_fa11_13_f_u_arrmul24_fa12_12_y2 = f_u_arrmul24_fa12_12_y2;
  assign f_u_arrmul24_fa11_13_f_u_arrmul24_fa10_13_y4 = f_u_arrmul24_fa10_13_y4;
  assign f_u_arrmul24_fa11_13_y0 = f_u_arrmul24_fa11_13_f_u_arrmul24_and11_13_y0 ^ f_u_arrmul24_fa11_13_f_u_arrmul24_fa12_12_y2;
  assign f_u_arrmul24_fa11_13_y1 = f_u_arrmul24_fa11_13_f_u_arrmul24_and11_13_y0 & f_u_arrmul24_fa11_13_f_u_arrmul24_fa12_12_y2;
  assign f_u_arrmul24_fa11_13_y2 = f_u_arrmul24_fa11_13_y0 ^ f_u_arrmul24_fa11_13_f_u_arrmul24_fa10_13_y4;
  assign f_u_arrmul24_fa11_13_y3 = f_u_arrmul24_fa11_13_y0 & f_u_arrmul24_fa11_13_f_u_arrmul24_fa10_13_y4;
  assign f_u_arrmul24_fa11_13_y4 = f_u_arrmul24_fa11_13_y1 | f_u_arrmul24_fa11_13_y3;
  assign f_u_arrmul24_and12_13_a_12 = a_12;
  assign f_u_arrmul24_and12_13_b_13 = b_13;
  assign f_u_arrmul24_and12_13_y0 = f_u_arrmul24_and12_13_a_12 & f_u_arrmul24_and12_13_b_13;
  assign f_u_arrmul24_fa12_13_f_u_arrmul24_and12_13_y0 = f_u_arrmul24_and12_13_y0;
  assign f_u_arrmul24_fa12_13_f_u_arrmul24_fa13_12_y2 = f_u_arrmul24_fa13_12_y2;
  assign f_u_arrmul24_fa12_13_f_u_arrmul24_fa11_13_y4 = f_u_arrmul24_fa11_13_y4;
  assign f_u_arrmul24_fa12_13_y0 = f_u_arrmul24_fa12_13_f_u_arrmul24_and12_13_y0 ^ f_u_arrmul24_fa12_13_f_u_arrmul24_fa13_12_y2;
  assign f_u_arrmul24_fa12_13_y1 = f_u_arrmul24_fa12_13_f_u_arrmul24_and12_13_y0 & f_u_arrmul24_fa12_13_f_u_arrmul24_fa13_12_y2;
  assign f_u_arrmul24_fa12_13_y2 = f_u_arrmul24_fa12_13_y0 ^ f_u_arrmul24_fa12_13_f_u_arrmul24_fa11_13_y4;
  assign f_u_arrmul24_fa12_13_y3 = f_u_arrmul24_fa12_13_y0 & f_u_arrmul24_fa12_13_f_u_arrmul24_fa11_13_y4;
  assign f_u_arrmul24_fa12_13_y4 = f_u_arrmul24_fa12_13_y1 | f_u_arrmul24_fa12_13_y3;
  assign f_u_arrmul24_and13_13_a_13 = a_13;
  assign f_u_arrmul24_and13_13_b_13 = b_13;
  assign f_u_arrmul24_and13_13_y0 = f_u_arrmul24_and13_13_a_13 & f_u_arrmul24_and13_13_b_13;
  assign f_u_arrmul24_fa13_13_f_u_arrmul24_and13_13_y0 = f_u_arrmul24_and13_13_y0;
  assign f_u_arrmul24_fa13_13_f_u_arrmul24_fa14_12_y2 = f_u_arrmul24_fa14_12_y2;
  assign f_u_arrmul24_fa13_13_f_u_arrmul24_fa12_13_y4 = f_u_arrmul24_fa12_13_y4;
  assign f_u_arrmul24_fa13_13_y0 = f_u_arrmul24_fa13_13_f_u_arrmul24_and13_13_y0 ^ f_u_arrmul24_fa13_13_f_u_arrmul24_fa14_12_y2;
  assign f_u_arrmul24_fa13_13_y1 = f_u_arrmul24_fa13_13_f_u_arrmul24_and13_13_y0 & f_u_arrmul24_fa13_13_f_u_arrmul24_fa14_12_y2;
  assign f_u_arrmul24_fa13_13_y2 = f_u_arrmul24_fa13_13_y0 ^ f_u_arrmul24_fa13_13_f_u_arrmul24_fa12_13_y4;
  assign f_u_arrmul24_fa13_13_y3 = f_u_arrmul24_fa13_13_y0 & f_u_arrmul24_fa13_13_f_u_arrmul24_fa12_13_y4;
  assign f_u_arrmul24_fa13_13_y4 = f_u_arrmul24_fa13_13_y1 | f_u_arrmul24_fa13_13_y3;
  assign f_u_arrmul24_and14_13_a_14 = a_14;
  assign f_u_arrmul24_and14_13_b_13 = b_13;
  assign f_u_arrmul24_and14_13_y0 = f_u_arrmul24_and14_13_a_14 & f_u_arrmul24_and14_13_b_13;
  assign f_u_arrmul24_fa14_13_f_u_arrmul24_and14_13_y0 = f_u_arrmul24_and14_13_y0;
  assign f_u_arrmul24_fa14_13_f_u_arrmul24_fa15_12_y2 = f_u_arrmul24_fa15_12_y2;
  assign f_u_arrmul24_fa14_13_f_u_arrmul24_fa13_13_y4 = f_u_arrmul24_fa13_13_y4;
  assign f_u_arrmul24_fa14_13_y0 = f_u_arrmul24_fa14_13_f_u_arrmul24_and14_13_y0 ^ f_u_arrmul24_fa14_13_f_u_arrmul24_fa15_12_y2;
  assign f_u_arrmul24_fa14_13_y1 = f_u_arrmul24_fa14_13_f_u_arrmul24_and14_13_y0 & f_u_arrmul24_fa14_13_f_u_arrmul24_fa15_12_y2;
  assign f_u_arrmul24_fa14_13_y2 = f_u_arrmul24_fa14_13_y0 ^ f_u_arrmul24_fa14_13_f_u_arrmul24_fa13_13_y4;
  assign f_u_arrmul24_fa14_13_y3 = f_u_arrmul24_fa14_13_y0 & f_u_arrmul24_fa14_13_f_u_arrmul24_fa13_13_y4;
  assign f_u_arrmul24_fa14_13_y4 = f_u_arrmul24_fa14_13_y1 | f_u_arrmul24_fa14_13_y3;
  assign f_u_arrmul24_and15_13_a_15 = a_15;
  assign f_u_arrmul24_and15_13_b_13 = b_13;
  assign f_u_arrmul24_and15_13_y0 = f_u_arrmul24_and15_13_a_15 & f_u_arrmul24_and15_13_b_13;
  assign f_u_arrmul24_fa15_13_f_u_arrmul24_and15_13_y0 = f_u_arrmul24_and15_13_y0;
  assign f_u_arrmul24_fa15_13_f_u_arrmul24_fa16_12_y2 = f_u_arrmul24_fa16_12_y2;
  assign f_u_arrmul24_fa15_13_f_u_arrmul24_fa14_13_y4 = f_u_arrmul24_fa14_13_y4;
  assign f_u_arrmul24_fa15_13_y0 = f_u_arrmul24_fa15_13_f_u_arrmul24_and15_13_y0 ^ f_u_arrmul24_fa15_13_f_u_arrmul24_fa16_12_y2;
  assign f_u_arrmul24_fa15_13_y1 = f_u_arrmul24_fa15_13_f_u_arrmul24_and15_13_y0 & f_u_arrmul24_fa15_13_f_u_arrmul24_fa16_12_y2;
  assign f_u_arrmul24_fa15_13_y2 = f_u_arrmul24_fa15_13_y0 ^ f_u_arrmul24_fa15_13_f_u_arrmul24_fa14_13_y4;
  assign f_u_arrmul24_fa15_13_y3 = f_u_arrmul24_fa15_13_y0 & f_u_arrmul24_fa15_13_f_u_arrmul24_fa14_13_y4;
  assign f_u_arrmul24_fa15_13_y4 = f_u_arrmul24_fa15_13_y1 | f_u_arrmul24_fa15_13_y3;
  assign f_u_arrmul24_and16_13_a_16 = a_16;
  assign f_u_arrmul24_and16_13_b_13 = b_13;
  assign f_u_arrmul24_and16_13_y0 = f_u_arrmul24_and16_13_a_16 & f_u_arrmul24_and16_13_b_13;
  assign f_u_arrmul24_fa16_13_f_u_arrmul24_and16_13_y0 = f_u_arrmul24_and16_13_y0;
  assign f_u_arrmul24_fa16_13_f_u_arrmul24_fa17_12_y2 = f_u_arrmul24_fa17_12_y2;
  assign f_u_arrmul24_fa16_13_f_u_arrmul24_fa15_13_y4 = f_u_arrmul24_fa15_13_y4;
  assign f_u_arrmul24_fa16_13_y0 = f_u_arrmul24_fa16_13_f_u_arrmul24_and16_13_y0 ^ f_u_arrmul24_fa16_13_f_u_arrmul24_fa17_12_y2;
  assign f_u_arrmul24_fa16_13_y1 = f_u_arrmul24_fa16_13_f_u_arrmul24_and16_13_y0 & f_u_arrmul24_fa16_13_f_u_arrmul24_fa17_12_y2;
  assign f_u_arrmul24_fa16_13_y2 = f_u_arrmul24_fa16_13_y0 ^ f_u_arrmul24_fa16_13_f_u_arrmul24_fa15_13_y4;
  assign f_u_arrmul24_fa16_13_y3 = f_u_arrmul24_fa16_13_y0 & f_u_arrmul24_fa16_13_f_u_arrmul24_fa15_13_y4;
  assign f_u_arrmul24_fa16_13_y4 = f_u_arrmul24_fa16_13_y1 | f_u_arrmul24_fa16_13_y3;
  assign f_u_arrmul24_and17_13_a_17 = a_17;
  assign f_u_arrmul24_and17_13_b_13 = b_13;
  assign f_u_arrmul24_and17_13_y0 = f_u_arrmul24_and17_13_a_17 & f_u_arrmul24_and17_13_b_13;
  assign f_u_arrmul24_fa17_13_f_u_arrmul24_and17_13_y0 = f_u_arrmul24_and17_13_y0;
  assign f_u_arrmul24_fa17_13_f_u_arrmul24_fa18_12_y2 = f_u_arrmul24_fa18_12_y2;
  assign f_u_arrmul24_fa17_13_f_u_arrmul24_fa16_13_y4 = f_u_arrmul24_fa16_13_y4;
  assign f_u_arrmul24_fa17_13_y0 = f_u_arrmul24_fa17_13_f_u_arrmul24_and17_13_y0 ^ f_u_arrmul24_fa17_13_f_u_arrmul24_fa18_12_y2;
  assign f_u_arrmul24_fa17_13_y1 = f_u_arrmul24_fa17_13_f_u_arrmul24_and17_13_y0 & f_u_arrmul24_fa17_13_f_u_arrmul24_fa18_12_y2;
  assign f_u_arrmul24_fa17_13_y2 = f_u_arrmul24_fa17_13_y0 ^ f_u_arrmul24_fa17_13_f_u_arrmul24_fa16_13_y4;
  assign f_u_arrmul24_fa17_13_y3 = f_u_arrmul24_fa17_13_y0 & f_u_arrmul24_fa17_13_f_u_arrmul24_fa16_13_y4;
  assign f_u_arrmul24_fa17_13_y4 = f_u_arrmul24_fa17_13_y1 | f_u_arrmul24_fa17_13_y3;
  assign f_u_arrmul24_and18_13_a_18 = a_18;
  assign f_u_arrmul24_and18_13_b_13 = b_13;
  assign f_u_arrmul24_and18_13_y0 = f_u_arrmul24_and18_13_a_18 & f_u_arrmul24_and18_13_b_13;
  assign f_u_arrmul24_fa18_13_f_u_arrmul24_and18_13_y0 = f_u_arrmul24_and18_13_y0;
  assign f_u_arrmul24_fa18_13_f_u_arrmul24_fa19_12_y2 = f_u_arrmul24_fa19_12_y2;
  assign f_u_arrmul24_fa18_13_f_u_arrmul24_fa17_13_y4 = f_u_arrmul24_fa17_13_y4;
  assign f_u_arrmul24_fa18_13_y0 = f_u_arrmul24_fa18_13_f_u_arrmul24_and18_13_y0 ^ f_u_arrmul24_fa18_13_f_u_arrmul24_fa19_12_y2;
  assign f_u_arrmul24_fa18_13_y1 = f_u_arrmul24_fa18_13_f_u_arrmul24_and18_13_y0 & f_u_arrmul24_fa18_13_f_u_arrmul24_fa19_12_y2;
  assign f_u_arrmul24_fa18_13_y2 = f_u_arrmul24_fa18_13_y0 ^ f_u_arrmul24_fa18_13_f_u_arrmul24_fa17_13_y4;
  assign f_u_arrmul24_fa18_13_y3 = f_u_arrmul24_fa18_13_y0 & f_u_arrmul24_fa18_13_f_u_arrmul24_fa17_13_y4;
  assign f_u_arrmul24_fa18_13_y4 = f_u_arrmul24_fa18_13_y1 | f_u_arrmul24_fa18_13_y3;
  assign f_u_arrmul24_and19_13_a_19 = a_19;
  assign f_u_arrmul24_and19_13_b_13 = b_13;
  assign f_u_arrmul24_and19_13_y0 = f_u_arrmul24_and19_13_a_19 & f_u_arrmul24_and19_13_b_13;
  assign f_u_arrmul24_fa19_13_f_u_arrmul24_and19_13_y0 = f_u_arrmul24_and19_13_y0;
  assign f_u_arrmul24_fa19_13_f_u_arrmul24_fa20_12_y2 = f_u_arrmul24_fa20_12_y2;
  assign f_u_arrmul24_fa19_13_f_u_arrmul24_fa18_13_y4 = f_u_arrmul24_fa18_13_y4;
  assign f_u_arrmul24_fa19_13_y0 = f_u_arrmul24_fa19_13_f_u_arrmul24_and19_13_y0 ^ f_u_arrmul24_fa19_13_f_u_arrmul24_fa20_12_y2;
  assign f_u_arrmul24_fa19_13_y1 = f_u_arrmul24_fa19_13_f_u_arrmul24_and19_13_y0 & f_u_arrmul24_fa19_13_f_u_arrmul24_fa20_12_y2;
  assign f_u_arrmul24_fa19_13_y2 = f_u_arrmul24_fa19_13_y0 ^ f_u_arrmul24_fa19_13_f_u_arrmul24_fa18_13_y4;
  assign f_u_arrmul24_fa19_13_y3 = f_u_arrmul24_fa19_13_y0 & f_u_arrmul24_fa19_13_f_u_arrmul24_fa18_13_y4;
  assign f_u_arrmul24_fa19_13_y4 = f_u_arrmul24_fa19_13_y1 | f_u_arrmul24_fa19_13_y3;
  assign f_u_arrmul24_and20_13_a_20 = a_20;
  assign f_u_arrmul24_and20_13_b_13 = b_13;
  assign f_u_arrmul24_and20_13_y0 = f_u_arrmul24_and20_13_a_20 & f_u_arrmul24_and20_13_b_13;
  assign f_u_arrmul24_fa20_13_f_u_arrmul24_and20_13_y0 = f_u_arrmul24_and20_13_y0;
  assign f_u_arrmul24_fa20_13_f_u_arrmul24_fa21_12_y2 = f_u_arrmul24_fa21_12_y2;
  assign f_u_arrmul24_fa20_13_f_u_arrmul24_fa19_13_y4 = f_u_arrmul24_fa19_13_y4;
  assign f_u_arrmul24_fa20_13_y0 = f_u_arrmul24_fa20_13_f_u_arrmul24_and20_13_y0 ^ f_u_arrmul24_fa20_13_f_u_arrmul24_fa21_12_y2;
  assign f_u_arrmul24_fa20_13_y1 = f_u_arrmul24_fa20_13_f_u_arrmul24_and20_13_y0 & f_u_arrmul24_fa20_13_f_u_arrmul24_fa21_12_y2;
  assign f_u_arrmul24_fa20_13_y2 = f_u_arrmul24_fa20_13_y0 ^ f_u_arrmul24_fa20_13_f_u_arrmul24_fa19_13_y4;
  assign f_u_arrmul24_fa20_13_y3 = f_u_arrmul24_fa20_13_y0 & f_u_arrmul24_fa20_13_f_u_arrmul24_fa19_13_y4;
  assign f_u_arrmul24_fa20_13_y4 = f_u_arrmul24_fa20_13_y1 | f_u_arrmul24_fa20_13_y3;
  assign f_u_arrmul24_and21_13_a_21 = a_21;
  assign f_u_arrmul24_and21_13_b_13 = b_13;
  assign f_u_arrmul24_and21_13_y0 = f_u_arrmul24_and21_13_a_21 & f_u_arrmul24_and21_13_b_13;
  assign f_u_arrmul24_fa21_13_f_u_arrmul24_and21_13_y0 = f_u_arrmul24_and21_13_y0;
  assign f_u_arrmul24_fa21_13_f_u_arrmul24_fa22_12_y2 = f_u_arrmul24_fa22_12_y2;
  assign f_u_arrmul24_fa21_13_f_u_arrmul24_fa20_13_y4 = f_u_arrmul24_fa20_13_y4;
  assign f_u_arrmul24_fa21_13_y0 = f_u_arrmul24_fa21_13_f_u_arrmul24_and21_13_y0 ^ f_u_arrmul24_fa21_13_f_u_arrmul24_fa22_12_y2;
  assign f_u_arrmul24_fa21_13_y1 = f_u_arrmul24_fa21_13_f_u_arrmul24_and21_13_y0 & f_u_arrmul24_fa21_13_f_u_arrmul24_fa22_12_y2;
  assign f_u_arrmul24_fa21_13_y2 = f_u_arrmul24_fa21_13_y0 ^ f_u_arrmul24_fa21_13_f_u_arrmul24_fa20_13_y4;
  assign f_u_arrmul24_fa21_13_y3 = f_u_arrmul24_fa21_13_y0 & f_u_arrmul24_fa21_13_f_u_arrmul24_fa20_13_y4;
  assign f_u_arrmul24_fa21_13_y4 = f_u_arrmul24_fa21_13_y1 | f_u_arrmul24_fa21_13_y3;
  assign f_u_arrmul24_and22_13_a_22 = a_22;
  assign f_u_arrmul24_and22_13_b_13 = b_13;
  assign f_u_arrmul24_and22_13_y0 = f_u_arrmul24_and22_13_a_22 & f_u_arrmul24_and22_13_b_13;
  assign f_u_arrmul24_fa22_13_f_u_arrmul24_and22_13_y0 = f_u_arrmul24_and22_13_y0;
  assign f_u_arrmul24_fa22_13_f_u_arrmul24_fa23_12_y2 = f_u_arrmul24_fa23_12_y2;
  assign f_u_arrmul24_fa22_13_f_u_arrmul24_fa21_13_y4 = f_u_arrmul24_fa21_13_y4;
  assign f_u_arrmul24_fa22_13_y0 = f_u_arrmul24_fa22_13_f_u_arrmul24_and22_13_y0 ^ f_u_arrmul24_fa22_13_f_u_arrmul24_fa23_12_y2;
  assign f_u_arrmul24_fa22_13_y1 = f_u_arrmul24_fa22_13_f_u_arrmul24_and22_13_y0 & f_u_arrmul24_fa22_13_f_u_arrmul24_fa23_12_y2;
  assign f_u_arrmul24_fa22_13_y2 = f_u_arrmul24_fa22_13_y0 ^ f_u_arrmul24_fa22_13_f_u_arrmul24_fa21_13_y4;
  assign f_u_arrmul24_fa22_13_y3 = f_u_arrmul24_fa22_13_y0 & f_u_arrmul24_fa22_13_f_u_arrmul24_fa21_13_y4;
  assign f_u_arrmul24_fa22_13_y4 = f_u_arrmul24_fa22_13_y1 | f_u_arrmul24_fa22_13_y3;
  assign f_u_arrmul24_and23_13_a_23 = a_23;
  assign f_u_arrmul24_and23_13_b_13 = b_13;
  assign f_u_arrmul24_and23_13_y0 = f_u_arrmul24_and23_13_a_23 & f_u_arrmul24_and23_13_b_13;
  assign f_u_arrmul24_fa23_13_f_u_arrmul24_and23_13_y0 = f_u_arrmul24_and23_13_y0;
  assign f_u_arrmul24_fa23_13_f_u_arrmul24_fa23_12_y4 = f_u_arrmul24_fa23_12_y4;
  assign f_u_arrmul24_fa23_13_f_u_arrmul24_fa22_13_y4 = f_u_arrmul24_fa22_13_y4;
  assign f_u_arrmul24_fa23_13_y0 = f_u_arrmul24_fa23_13_f_u_arrmul24_and23_13_y0 ^ f_u_arrmul24_fa23_13_f_u_arrmul24_fa23_12_y4;
  assign f_u_arrmul24_fa23_13_y1 = f_u_arrmul24_fa23_13_f_u_arrmul24_and23_13_y0 & f_u_arrmul24_fa23_13_f_u_arrmul24_fa23_12_y4;
  assign f_u_arrmul24_fa23_13_y2 = f_u_arrmul24_fa23_13_y0 ^ f_u_arrmul24_fa23_13_f_u_arrmul24_fa22_13_y4;
  assign f_u_arrmul24_fa23_13_y3 = f_u_arrmul24_fa23_13_y0 & f_u_arrmul24_fa23_13_f_u_arrmul24_fa22_13_y4;
  assign f_u_arrmul24_fa23_13_y4 = f_u_arrmul24_fa23_13_y1 | f_u_arrmul24_fa23_13_y3;
  assign f_u_arrmul24_and0_14_a_0 = a_0;
  assign f_u_arrmul24_and0_14_b_14 = b_14;
  assign f_u_arrmul24_and0_14_y0 = f_u_arrmul24_and0_14_a_0 & f_u_arrmul24_and0_14_b_14;
  assign f_u_arrmul24_ha0_14_f_u_arrmul24_and0_14_y0 = f_u_arrmul24_and0_14_y0;
  assign f_u_arrmul24_ha0_14_f_u_arrmul24_fa1_13_y2 = f_u_arrmul24_fa1_13_y2;
  assign f_u_arrmul24_ha0_14_y0 = f_u_arrmul24_ha0_14_f_u_arrmul24_and0_14_y0 ^ f_u_arrmul24_ha0_14_f_u_arrmul24_fa1_13_y2;
  assign f_u_arrmul24_ha0_14_y1 = f_u_arrmul24_ha0_14_f_u_arrmul24_and0_14_y0 & f_u_arrmul24_ha0_14_f_u_arrmul24_fa1_13_y2;
  assign f_u_arrmul24_and1_14_a_1 = a_1;
  assign f_u_arrmul24_and1_14_b_14 = b_14;
  assign f_u_arrmul24_and1_14_y0 = f_u_arrmul24_and1_14_a_1 & f_u_arrmul24_and1_14_b_14;
  assign f_u_arrmul24_fa1_14_f_u_arrmul24_and1_14_y0 = f_u_arrmul24_and1_14_y0;
  assign f_u_arrmul24_fa1_14_f_u_arrmul24_fa2_13_y2 = f_u_arrmul24_fa2_13_y2;
  assign f_u_arrmul24_fa1_14_f_u_arrmul24_ha0_14_y1 = f_u_arrmul24_ha0_14_y1;
  assign f_u_arrmul24_fa1_14_y0 = f_u_arrmul24_fa1_14_f_u_arrmul24_and1_14_y0 ^ f_u_arrmul24_fa1_14_f_u_arrmul24_fa2_13_y2;
  assign f_u_arrmul24_fa1_14_y1 = f_u_arrmul24_fa1_14_f_u_arrmul24_and1_14_y0 & f_u_arrmul24_fa1_14_f_u_arrmul24_fa2_13_y2;
  assign f_u_arrmul24_fa1_14_y2 = f_u_arrmul24_fa1_14_y0 ^ f_u_arrmul24_fa1_14_f_u_arrmul24_ha0_14_y1;
  assign f_u_arrmul24_fa1_14_y3 = f_u_arrmul24_fa1_14_y0 & f_u_arrmul24_fa1_14_f_u_arrmul24_ha0_14_y1;
  assign f_u_arrmul24_fa1_14_y4 = f_u_arrmul24_fa1_14_y1 | f_u_arrmul24_fa1_14_y3;
  assign f_u_arrmul24_and2_14_a_2 = a_2;
  assign f_u_arrmul24_and2_14_b_14 = b_14;
  assign f_u_arrmul24_and2_14_y0 = f_u_arrmul24_and2_14_a_2 & f_u_arrmul24_and2_14_b_14;
  assign f_u_arrmul24_fa2_14_f_u_arrmul24_and2_14_y0 = f_u_arrmul24_and2_14_y0;
  assign f_u_arrmul24_fa2_14_f_u_arrmul24_fa3_13_y2 = f_u_arrmul24_fa3_13_y2;
  assign f_u_arrmul24_fa2_14_f_u_arrmul24_fa1_14_y4 = f_u_arrmul24_fa1_14_y4;
  assign f_u_arrmul24_fa2_14_y0 = f_u_arrmul24_fa2_14_f_u_arrmul24_and2_14_y0 ^ f_u_arrmul24_fa2_14_f_u_arrmul24_fa3_13_y2;
  assign f_u_arrmul24_fa2_14_y1 = f_u_arrmul24_fa2_14_f_u_arrmul24_and2_14_y0 & f_u_arrmul24_fa2_14_f_u_arrmul24_fa3_13_y2;
  assign f_u_arrmul24_fa2_14_y2 = f_u_arrmul24_fa2_14_y0 ^ f_u_arrmul24_fa2_14_f_u_arrmul24_fa1_14_y4;
  assign f_u_arrmul24_fa2_14_y3 = f_u_arrmul24_fa2_14_y0 & f_u_arrmul24_fa2_14_f_u_arrmul24_fa1_14_y4;
  assign f_u_arrmul24_fa2_14_y4 = f_u_arrmul24_fa2_14_y1 | f_u_arrmul24_fa2_14_y3;
  assign f_u_arrmul24_and3_14_a_3 = a_3;
  assign f_u_arrmul24_and3_14_b_14 = b_14;
  assign f_u_arrmul24_and3_14_y0 = f_u_arrmul24_and3_14_a_3 & f_u_arrmul24_and3_14_b_14;
  assign f_u_arrmul24_fa3_14_f_u_arrmul24_and3_14_y0 = f_u_arrmul24_and3_14_y0;
  assign f_u_arrmul24_fa3_14_f_u_arrmul24_fa4_13_y2 = f_u_arrmul24_fa4_13_y2;
  assign f_u_arrmul24_fa3_14_f_u_arrmul24_fa2_14_y4 = f_u_arrmul24_fa2_14_y4;
  assign f_u_arrmul24_fa3_14_y0 = f_u_arrmul24_fa3_14_f_u_arrmul24_and3_14_y0 ^ f_u_arrmul24_fa3_14_f_u_arrmul24_fa4_13_y2;
  assign f_u_arrmul24_fa3_14_y1 = f_u_arrmul24_fa3_14_f_u_arrmul24_and3_14_y0 & f_u_arrmul24_fa3_14_f_u_arrmul24_fa4_13_y2;
  assign f_u_arrmul24_fa3_14_y2 = f_u_arrmul24_fa3_14_y0 ^ f_u_arrmul24_fa3_14_f_u_arrmul24_fa2_14_y4;
  assign f_u_arrmul24_fa3_14_y3 = f_u_arrmul24_fa3_14_y0 & f_u_arrmul24_fa3_14_f_u_arrmul24_fa2_14_y4;
  assign f_u_arrmul24_fa3_14_y4 = f_u_arrmul24_fa3_14_y1 | f_u_arrmul24_fa3_14_y3;
  assign f_u_arrmul24_and4_14_a_4 = a_4;
  assign f_u_arrmul24_and4_14_b_14 = b_14;
  assign f_u_arrmul24_and4_14_y0 = f_u_arrmul24_and4_14_a_4 & f_u_arrmul24_and4_14_b_14;
  assign f_u_arrmul24_fa4_14_f_u_arrmul24_and4_14_y0 = f_u_arrmul24_and4_14_y0;
  assign f_u_arrmul24_fa4_14_f_u_arrmul24_fa5_13_y2 = f_u_arrmul24_fa5_13_y2;
  assign f_u_arrmul24_fa4_14_f_u_arrmul24_fa3_14_y4 = f_u_arrmul24_fa3_14_y4;
  assign f_u_arrmul24_fa4_14_y0 = f_u_arrmul24_fa4_14_f_u_arrmul24_and4_14_y0 ^ f_u_arrmul24_fa4_14_f_u_arrmul24_fa5_13_y2;
  assign f_u_arrmul24_fa4_14_y1 = f_u_arrmul24_fa4_14_f_u_arrmul24_and4_14_y0 & f_u_arrmul24_fa4_14_f_u_arrmul24_fa5_13_y2;
  assign f_u_arrmul24_fa4_14_y2 = f_u_arrmul24_fa4_14_y0 ^ f_u_arrmul24_fa4_14_f_u_arrmul24_fa3_14_y4;
  assign f_u_arrmul24_fa4_14_y3 = f_u_arrmul24_fa4_14_y0 & f_u_arrmul24_fa4_14_f_u_arrmul24_fa3_14_y4;
  assign f_u_arrmul24_fa4_14_y4 = f_u_arrmul24_fa4_14_y1 | f_u_arrmul24_fa4_14_y3;
  assign f_u_arrmul24_and5_14_a_5 = a_5;
  assign f_u_arrmul24_and5_14_b_14 = b_14;
  assign f_u_arrmul24_and5_14_y0 = f_u_arrmul24_and5_14_a_5 & f_u_arrmul24_and5_14_b_14;
  assign f_u_arrmul24_fa5_14_f_u_arrmul24_and5_14_y0 = f_u_arrmul24_and5_14_y0;
  assign f_u_arrmul24_fa5_14_f_u_arrmul24_fa6_13_y2 = f_u_arrmul24_fa6_13_y2;
  assign f_u_arrmul24_fa5_14_f_u_arrmul24_fa4_14_y4 = f_u_arrmul24_fa4_14_y4;
  assign f_u_arrmul24_fa5_14_y0 = f_u_arrmul24_fa5_14_f_u_arrmul24_and5_14_y0 ^ f_u_arrmul24_fa5_14_f_u_arrmul24_fa6_13_y2;
  assign f_u_arrmul24_fa5_14_y1 = f_u_arrmul24_fa5_14_f_u_arrmul24_and5_14_y0 & f_u_arrmul24_fa5_14_f_u_arrmul24_fa6_13_y2;
  assign f_u_arrmul24_fa5_14_y2 = f_u_arrmul24_fa5_14_y0 ^ f_u_arrmul24_fa5_14_f_u_arrmul24_fa4_14_y4;
  assign f_u_arrmul24_fa5_14_y3 = f_u_arrmul24_fa5_14_y0 & f_u_arrmul24_fa5_14_f_u_arrmul24_fa4_14_y4;
  assign f_u_arrmul24_fa5_14_y4 = f_u_arrmul24_fa5_14_y1 | f_u_arrmul24_fa5_14_y3;
  assign f_u_arrmul24_and6_14_a_6 = a_6;
  assign f_u_arrmul24_and6_14_b_14 = b_14;
  assign f_u_arrmul24_and6_14_y0 = f_u_arrmul24_and6_14_a_6 & f_u_arrmul24_and6_14_b_14;
  assign f_u_arrmul24_fa6_14_f_u_arrmul24_and6_14_y0 = f_u_arrmul24_and6_14_y0;
  assign f_u_arrmul24_fa6_14_f_u_arrmul24_fa7_13_y2 = f_u_arrmul24_fa7_13_y2;
  assign f_u_arrmul24_fa6_14_f_u_arrmul24_fa5_14_y4 = f_u_arrmul24_fa5_14_y4;
  assign f_u_arrmul24_fa6_14_y0 = f_u_arrmul24_fa6_14_f_u_arrmul24_and6_14_y0 ^ f_u_arrmul24_fa6_14_f_u_arrmul24_fa7_13_y2;
  assign f_u_arrmul24_fa6_14_y1 = f_u_arrmul24_fa6_14_f_u_arrmul24_and6_14_y0 & f_u_arrmul24_fa6_14_f_u_arrmul24_fa7_13_y2;
  assign f_u_arrmul24_fa6_14_y2 = f_u_arrmul24_fa6_14_y0 ^ f_u_arrmul24_fa6_14_f_u_arrmul24_fa5_14_y4;
  assign f_u_arrmul24_fa6_14_y3 = f_u_arrmul24_fa6_14_y0 & f_u_arrmul24_fa6_14_f_u_arrmul24_fa5_14_y4;
  assign f_u_arrmul24_fa6_14_y4 = f_u_arrmul24_fa6_14_y1 | f_u_arrmul24_fa6_14_y3;
  assign f_u_arrmul24_and7_14_a_7 = a_7;
  assign f_u_arrmul24_and7_14_b_14 = b_14;
  assign f_u_arrmul24_and7_14_y0 = f_u_arrmul24_and7_14_a_7 & f_u_arrmul24_and7_14_b_14;
  assign f_u_arrmul24_fa7_14_f_u_arrmul24_and7_14_y0 = f_u_arrmul24_and7_14_y0;
  assign f_u_arrmul24_fa7_14_f_u_arrmul24_fa8_13_y2 = f_u_arrmul24_fa8_13_y2;
  assign f_u_arrmul24_fa7_14_f_u_arrmul24_fa6_14_y4 = f_u_arrmul24_fa6_14_y4;
  assign f_u_arrmul24_fa7_14_y0 = f_u_arrmul24_fa7_14_f_u_arrmul24_and7_14_y0 ^ f_u_arrmul24_fa7_14_f_u_arrmul24_fa8_13_y2;
  assign f_u_arrmul24_fa7_14_y1 = f_u_arrmul24_fa7_14_f_u_arrmul24_and7_14_y0 & f_u_arrmul24_fa7_14_f_u_arrmul24_fa8_13_y2;
  assign f_u_arrmul24_fa7_14_y2 = f_u_arrmul24_fa7_14_y0 ^ f_u_arrmul24_fa7_14_f_u_arrmul24_fa6_14_y4;
  assign f_u_arrmul24_fa7_14_y3 = f_u_arrmul24_fa7_14_y0 & f_u_arrmul24_fa7_14_f_u_arrmul24_fa6_14_y4;
  assign f_u_arrmul24_fa7_14_y4 = f_u_arrmul24_fa7_14_y1 | f_u_arrmul24_fa7_14_y3;
  assign f_u_arrmul24_and8_14_a_8 = a_8;
  assign f_u_arrmul24_and8_14_b_14 = b_14;
  assign f_u_arrmul24_and8_14_y0 = f_u_arrmul24_and8_14_a_8 & f_u_arrmul24_and8_14_b_14;
  assign f_u_arrmul24_fa8_14_f_u_arrmul24_and8_14_y0 = f_u_arrmul24_and8_14_y0;
  assign f_u_arrmul24_fa8_14_f_u_arrmul24_fa9_13_y2 = f_u_arrmul24_fa9_13_y2;
  assign f_u_arrmul24_fa8_14_f_u_arrmul24_fa7_14_y4 = f_u_arrmul24_fa7_14_y4;
  assign f_u_arrmul24_fa8_14_y0 = f_u_arrmul24_fa8_14_f_u_arrmul24_and8_14_y0 ^ f_u_arrmul24_fa8_14_f_u_arrmul24_fa9_13_y2;
  assign f_u_arrmul24_fa8_14_y1 = f_u_arrmul24_fa8_14_f_u_arrmul24_and8_14_y0 & f_u_arrmul24_fa8_14_f_u_arrmul24_fa9_13_y2;
  assign f_u_arrmul24_fa8_14_y2 = f_u_arrmul24_fa8_14_y0 ^ f_u_arrmul24_fa8_14_f_u_arrmul24_fa7_14_y4;
  assign f_u_arrmul24_fa8_14_y3 = f_u_arrmul24_fa8_14_y0 & f_u_arrmul24_fa8_14_f_u_arrmul24_fa7_14_y4;
  assign f_u_arrmul24_fa8_14_y4 = f_u_arrmul24_fa8_14_y1 | f_u_arrmul24_fa8_14_y3;
  assign f_u_arrmul24_and9_14_a_9 = a_9;
  assign f_u_arrmul24_and9_14_b_14 = b_14;
  assign f_u_arrmul24_and9_14_y0 = f_u_arrmul24_and9_14_a_9 & f_u_arrmul24_and9_14_b_14;
  assign f_u_arrmul24_fa9_14_f_u_arrmul24_and9_14_y0 = f_u_arrmul24_and9_14_y0;
  assign f_u_arrmul24_fa9_14_f_u_arrmul24_fa10_13_y2 = f_u_arrmul24_fa10_13_y2;
  assign f_u_arrmul24_fa9_14_f_u_arrmul24_fa8_14_y4 = f_u_arrmul24_fa8_14_y4;
  assign f_u_arrmul24_fa9_14_y0 = f_u_arrmul24_fa9_14_f_u_arrmul24_and9_14_y0 ^ f_u_arrmul24_fa9_14_f_u_arrmul24_fa10_13_y2;
  assign f_u_arrmul24_fa9_14_y1 = f_u_arrmul24_fa9_14_f_u_arrmul24_and9_14_y0 & f_u_arrmul24_fa9_14_f_u_arrmul24_fa10_13_y2;
  assign f_u_arrmul24_fa9_14_y2 = f_u_arrmul24_fa9_14_y0 ^ f_u_arrmul24_fa9_14_f_u_arrmul24_fa8_14_y4;
  assign f_u_arrmul24_fa9_14_y3 = f_u_arrmul24_fa9_14_y0 & f_u_arrmul24_fa9_14_f_u_arrmul24_fa8_14_y4;
  assign f_u_arrmul24_fa9_14_y4 = f_u_arrmul24_fa9_14_y1 | f_u_arrmul24_fa9_14_y3;
  assign f_u_arrmul24_and10_14_a_10 = a_10;
  assign f_u_arrmul24_and10_14_b_14 = b_14;
  assign f_u_arrmul24_and10_14_y0 = f_u_arrmul24_and10_14_a_10 & f_u_arrmul24_and10_14_b_14;
  assign f_u_arrmul24_fa10_14_f_u_arrmul24_and10_14_y0 = f_u_arrmul24_and10_14_y0;
  assign f_u_arrmul24_fa10_14_f_u_arrmul24_fa11_13_y2 = f_u_arrmul24_fa11_13_y2;
  assign f_u_arrmul24_fa10_14_f_u_arrmul24_fa9_14_y4 = f_u_arrmul24_fa9_14_y4;
  assign f_u_arrmul24_fa10_14_y0 = f_u_arrmul24_fa10_14_f_u_arrmul24_and10_14_y0 ^ f_u_arrmul24_fa10_14_f_u_arrmul24_fa11_13_y2;
  assign f_u_arrmul24_fa10_14_y1 = f_u_arrmul24_fa10_14_f_u_arrmul24_and10_14_y0 & f_u_arrmul24_fa10_14_f_u_arrmul24_fa11_13_y2;
  assign f_u_arrmul24_fa10_14_y2 = f_u_arrmul24_fa10_14_y0 ^ f_u_arrmul24_fa10_14_f_u_arrmul24_fa9_14_y4;
  assign f_u_arrmul24_fa10_14_y3 = f_u_arrmul24_fa10_14_y0 & f_u_arrmul24_fa10_14_f_u_arrmul24_fa9_14_y4;
  assign f_u_arrmul24_fa10_14_y4 = f_u_arrmul24_fa10_14_y1 | f_u_arrmul24_fa10_14_y3;
  assign f_u_arrmul24_and11_14_a_11 = a_11;
  assign f_u_arrmul24_and11_14_b_14 = b_14;
  assign f_u_arrmul24_and11_14_y0 = f_u_arrmul24_and11_14_a_11 & f_u_arrmul24_and11_14_b_14;
  assign f_u_arrmul24_fa11_14_f_u_arrmul24_and11_14_y0 = f_u_arrmul24_and11_14_y0;
  assign f_u_arrmul24_fa11_14_f_u_arrmul24_fa12_13_y2 = f_u_arrmul24_fa12_13_y2;
  assign f_u_arrmul24_fa11_14_f_u_arrmul24_fa10_14_y4 = f_u_arrmul24_fa10_14_y4;
  assign f_u_arrmul24_fa11_14_y0 = f_u_arrmul24_fa11_14_f_u_arrmul24_and11_14_y0 ^ f_u_arrmul24_fa11_14_f_u_arrmul24_fa12_13_y2;
  assign f_u_arrmul24_fa11_14_y1 = f_u_arrmul24_fa11_14_f_u_arrmul24_and11_14_y0 & f_u_arrmul24_fa11_14_f_u_arrmul24_fa12_13_y2;
  assign f_u_arrmul24_fa11_14_y2 = f_u_arrmul24_fa11_14_y0 ^ f_u_arrmul24_fa11_14_f_u_arrmul24_fa10_14_y4;
  assign f_u_arrmul24_fa11_14_y3 = f_u_arrmul24_fa11_14_y0 & f_u_arrmul24_fa11_14_f_u_arrmul24_fa10_14_y4;
  assign f_u_arrmul24_fa11_14_y4 = f_u_arrmul24_fa11_14_y1 | f_u_arrmul24_fa11_14_y3;
  assign f_u_arrmul24_and12_14_a_12 = a_12;
  assign f_u_arrmul24_and12_14_b_14 = b_14;
  assign f_u_arrmul24_and12_14_y0 = f_u_arrmul24_and12_14_a_12 & f_u_arrmul24_and12_14_b_14;
  assign f_u_arrmul24_fa12_14_f_u_arrmul24_and12_14_y0 = f_u_arrmul24_and12_14_y0;
  assign f_u_arrmul24_fa12_14_f_u_arrmul24_fa13_13_y2 = f_u_arrmul24_fa13_13_y2;
  assign f_u_arrmul24_fa12_14_f_u_arrmul24_fa11_14_y4 = f_u_arrmul24_fa11_14_y4;
  assign f_u_arrmul24_fa12_14_y0 = f_u_arrmul24_fa12_14_f_u_arrmul24_and12_14_y0 ^ f_u_arrmul24_fa12_14_f_u_arrmul24_fa13_13_y2;
  assign f_u_arrmul24_fa12_14_y1 = f_u_arrmul24_fa12_14_f_u_arrmul24_and12_14_y0 & f_u_arrmul24_fa12_14_f_u_arrmul24_fa13_13_y2;
  assign f_u_arrmul24_fa12_14_y2 = f_u_arrmul24_fa12_14_y0 ^ f_u_arrmul24_fa12_14_f_u_arrmul24_fa11_14_y4;
  assign f_u_arrmul24_fa12_14_y3 = f_u_arrmul24_fa12_14_y0 & f_u_arrmul24_fa12_14_f_u_arrmul24_fa11_14_y4;
  assign f_u_arrmul24_fa12_14_y4 = f_u_arrmul24_fa12_14_y1 | f_u_arrmul24_fa12_14_y3;
  assign f_u_arrmul24_and13_14_a_13 = a_13;
  assign f_u_arrmul24_and13_14_b_14 = b_14;
  assign f_u_arrmul24_and13_14_y0 = f_u_arrmul24_and13_14_a_13 & f_u_arrmul24_and13_14_b_14;
  assign f_u_arrmul24_fa13_14_f_u_arrmul24_and13_14_y0 = f_u_arrmul24_and13_14_y0;
  assign f_u_arrmul24_fa13_14_f_u_arrmul24_fa14_13_y2 = f_u_arrmul24_fa14_13_y2;
  assign f_u_arrmul24_fa13_14_f_u_arrmul24_fa12_14_y4 = f_u_arrmul24_fa12_14_y4;
  assign f_u_arrmul24_fa13_14_y0 = f_u_arrmul24_fa13_14_f_u_arrmul24_and13_14_y0 ^ f_u_arrmul24_fa13_14_f_u_arrmul24_fa14_13_y2;
  assign f_u_arrmul24_fa13_14_y1 = f_u_arrmul24_fa13_14_f_u_arrmul24_and13_14_y0 & f_u_arrmul24_fa13_14_f_u_arrmul24_fa14_13_y2;
  assign f_u_arrmul24_fa13_14_y2 = f_u_arrmul24_fa13_14_y0 ^ f_u_arrmul24_fa13_14_f_u_arrmul24_fa12_14_y4;
  assign f_u_arrmul24_fa13_14_y3 = f_u_arrmul24_fa13_14_y0 & f_u_arrmul24_fa13_14_f_u_arrmul24_fa12_14_y4;
  assign f_u_arrmul24_fa13_14_y4 = f_u_arrmul24_fa13_14_y1 | f_u_arrmul24_fa13_14_y3;
  assign f_u_arrmul24_and14_14_a_14 = a_14;
  assign f_u_arrmul24_and14_14_b_14 = b_14;
  assign f_u_arrmul24_and14_14_y0 = f_u_arrmul24_and14_14_a_14 & f_u_arrmul24_and14_14_b_14;
  assign f_u_arrmul24_fa14_14_f_u_arrmul24_and14_14_y0 = f_u_arrmul24_and14_14_y0;
  assign f_u_arrmul24_fa14_14_f_u_arrmul24_fa15_13_y2 = f_u_arrmul24_fa15_13_y2;
  assign f_u_arrmul24_fa14_14_f_u_arrmul24_fa13_14_y4 = f_u_arrmul24_fa13_14_y4;
  assign f_u_arrmul24_fa14_14_y0 = f_u_arrmul24_fa14_14_f_u_arrmul24_and14_14_y0 ^ f_u_arrmul24_fa14_14_f_u_arrmul24_fa15_13_y2;
  assign f_u_arrmul24_fa14_14_y1 = f_u_arrmul24_fa14_14_f_u_arrmul24_and14_14_y0 & f_u_arrmul24_fa14_14_f_u_arrmul24_fa15_13_y2;
  assign f_u_arrmul24_fa14_14_y2 = f_u_arrmul24_fa14_14_y0 ^ f_u_arrmul24_fa14_14_f_u_arrmul24_fa13_14_y4;
  assign f_u_arrmul24_fa14_14_y3 = f_u_arrmul24_fa14_14_y0 & f_u_arrmul24_fa14_14_f_u_arrmul24_fa13_14_y4;
  assign f_u_arrmul24_fa14_14_y4 = f_u_arrmul24_fa14_14_y1 | f_u_arrmul24_fa14_14_y3;
  assign f_u_arrmul24_and15_14_a_15 = a_15;
  assign f_u_arrmul24_and15_14_b_14 = b_14;
  assign f_u_arrmul24_and15_14_y0 = f_u_arrmul24_and15_14_a_15 & f_u_arrmul24_and15_14_b_14;
  assign f_u_arrmul24_fa15_14_f_u_arrmul24_and15_14_y0 = f_u_arrmul24_and15_14_y0;
  assign f_u_arrmul24_fa15_14_f_u_arrmul24_fa16_13_y2 = f_u_arrmul24_fa16_13_y2;
  assign f_u_arrmul24_fa15_14_f_u_arrmul24_fa14_14_y4 = f_u_arrmul24_fa14_14_y4;
  assign f_u_arrmul24_fa15_14_y0 = f_u_arrmul24_fa15_14_f_u_arrmul24_and15_14_y0 ^ f_u_arrmul24_fa15_14_f_u_arrmul24_fa16_13_y2;
  assign f_u_arrmul24_fa15_14_y1 = f_u_arrmul24_fa15_14_f_u_arrmul24_and15_14_y0 & f_u_arrmul24_fa15_14_f_u_arrmul24_fa16_13_y2;
  assign f_u_arrmul24_fa15_14_y2 = f_u_arrmul24_fa15_14_y0 ^ f_u_arrmul24_fa15_14_f_u_arrmul24_fa14_14_y4;
  assign f_u_arrmul24_fa15_14_y3 = f_u_arrmul24_fa15_14_y0 & f_u_arrmul24_fa15_14_f_u_arrmul24_fa14_14_y4;
  assign f_u_arrmul24_fa15_14_y4 = f_u_arrmul24_fa15_14_y1 | f_u_arrmul24_fa15_14_y3;
  assign f_u_arrmul24_and16_14_a_16 = a_16;
  assign f_u_arrmul24_and16_14_b_14 = b_14;
  assign f_u_arrmul24_and16_14_y0 = f_u_arrmul24_and16_14_a_16 & f_u_arrmul24_and16_14_b_14;
  assign f_u_arrmul24_fa16_14_f_u_arrmul24_and16_14_y0 = f_u_arrmul24_and16_14_y0;
  assign f_u_arrmul24_fa16_14_f_u_arrmul24_fa17_13_y2 = f_u_arrmul24_fa17_13_y2;
  assign f_u_arrmul24_fa16_14_f_u_arrmul24_fa15_14_y4 = f_u_arrmul24_fa15_14_y4;
  assign f_u_arrmul24_fa16_14_y0 = f_u_arrmul24_fa16_14_f_u_arrmul24_and16_14_y0 ^ f_u_arrmul24_fa16_14_f_u_arrmul24_fa17_13_y2;
  assign f_u_arrmul24_fa16_14_y1 = f_u_arrmul24_fa16_14_f_u_arrmul24_and16_14_y0 & f_u_arrmul24_fa16_14_f_u_arrmul24_fa17_13_y2;
  assign f_u_arrmul24_fa16_14_y2 = f_u_arrmul24_fa16_14_y0 ^ f_u_arrmul24_fa16_14_f_u_arrmul24_fa15_14_y4;
  assign f_u_arrmul24_fa16_14_y3 = f_u_arrmul24_fa16_14_y0 & f_u_arrmul24_fa16_14_f_u_arrmul24_fa15_14_y4;
  assign f_u_arrmul24_fa16_14_y4 = f_u_arrmul24_fa16_14_y1 | f_u_arrmul24_fa16_14_y3;
  assign f_u_arrmul24_and17_14_a_17 = a_17;
  assign f_u_arrmul24_and17_14_b_14 = b_14;
  assign f_u_arrmul24_and17_14_y0 = f_u_arrmul24_and17_14_a_17 & f_u_arrmul24_and17_14_b_14;
  assign f_u_arrmul24_fa17_14_f_u_arrmul24_and17_14_y0 = f_u_arrmul24_and17_14_y0;
  assign f_u_arrmul24_fa17_14_f_u_arrmul24_fa18_13_y2 = f_u_arrmul24_fa18_13_y2;
  assign f_u_arrmul24_fa17_14_f_u_arrmul24_fa16_14_y4 = f_u_arrmul24_fa16_14_y4;
  assign f_u_arrmul24_fa17_14_y0 = f_u_arrmul24_fa17_14_f_u_arrmul24_and17_14_y0 ^ f_u_arrmul24_fa17_14_f_u_arrmul24_fa18_13_y2;
  assign f_u_arrmul24_fa17_14_y1 = f_u_arrmul24_fa17_14_f_u_arrmul24_and17_14_y0 & f_u_arrmul24_fa17_14_f_u_arrmul24_fa18_13_y2;
  assign f_u_arrmul24_fa17_14_y2 = f_u_arrmul24_fa17_14_y0 ^ f_u_arrmul24_fa17_14_f_u_arrmul24_fa16_14_y4;
  assign f_u_arrmul24_fa17_14_y3 = f_u_arrmul24_fa17_14_y0 & f_u_arrmul24_fa17_14_f_u_arrmul24_fa16_14_y4;
  assign f_u_arrmul24_fa17_14_y4 = f_u_arrmul24_fa17_14_y1 | f_u_arrmul24_fa17_14_y3;
  assign f_u_arrmul24_and18_14_a_18 = a_18;
  assign f_u_arrmul24_and18_14_b_14 = b_14;
  assign f_u_arrmul24_and18_14_y0 = f_u_arrmul24_and18_14_a_18 & f_u_arrmul24_and18_14_b_14;
  assign f_u_arrmul24_fa18_14_f_u_arrmul24_and18_14_y0 = f_u_arrmul24_and18_14_y0;
  assign f_u_arrmul24_fa18_14_f_u_arrmul24_fa19_13_y2 = f_u_arrmul24_fa19_13_y2;
  assign f_u_arrmul24_fa18_14_f_u_arrmul24_fa17_14_y4 = f_u_arrmul24_fa17_14_y4;
  assign f_u_arrmul24_fa18_14_y0 = f_u_arrmul24_fa18_14_f_u_arrmul24_and18_14_y0 ^ f_u_arrmul24_fa18_14_f_u_arrmul24_fa19_13_y2;
  assign f_u_arrmul24_fa18_14_y1 = f_u_arrmul24_fa18_14_f_u_arrmul24_and18_14_y0 & f_u_arrmul24_fa18_14_f_u_arrmul24_fa19_13_y2;
  assign f_u_arrmul24_fa18_14_y2 = f_u_arrmul24_fa18_14_y0 ^ f_u_arrmul24_fa18_14_f_u_arrmul24_fa17_14_y4;
  assign f_u_arrmul24_fa18_14_y3 = f_u_arrmul24_fa18_14_y0 & f_u_arrmul24_fa18_14_f_u_arrmul24_fa17_14_y4;
  assign f_u_arrmul24_fa18_14_y4 = f_u_arrmul24_fa18_14_y1 | f_u_arrmul24_fa18_14_y3;
  assign f_u_arrmul24_and19_14_a_19 = a_19;
  assign f_u_arrmul24_and19_14_b_14 = b_14;
  assign f_u_arrmul24_and19_14_y0 = f_u_arrmul24_and19_14_a_19 & f_u_arrmul24_and19_14_b_14;
  assign f_u_arrmul24_fa19_14_f_u_arrmul24_and19_14_y0 = f_u_arrmul24_and19_14_y0;
  assign f_u_arrmul24_fa19_14_f_u_arrmul24_fa20_13_y2 = f_u_arrmul24_fa20_13_y2;
  assign f_u_arrmul24_fa19_14_f_u_arrmul24_fa18_14_y4 = f_u_arrmul24_fa18_14_y4;
  assign f_u_arrmul24_fa19_14_y0 = f_u_arrmul24_fa19_14_f_u_arrmul24_and19_14_y0 ^ f_u_arrmul24_fa19_14_f_u_arrmul24_fa20_13_y2;
  assign f_u_arrmul24_fa19_14_y1 = f_u_arrmul24_fa19_14_f_u_arrmul24_and19_14_y0 & f_u_arrmul24_fa19_14_f_u_arrmul24_fa20_13_y2;
  assign f_u_arrmul24_fa19_14_y2 = f_u_arrmul24_fa19_14_y0 ^ f_u_arrmul24_fa19_14_f_u_arrmul24_fa18_14_y4;
  assign f_u_arrmul24_fa19_14_y3 = f_u_arrmul24_fa19_14_y0 & f_u_arrmul24_fa19_14_f_u_arrmul24_fa18_14_y4;
  assign f_u_arrmul24_fa19_14_y4 = f_u_arrmul24_fa19_14_y1 | f_u_arrmul24_fa19_14_y3;
  assign f_u_arrmul24_and20_14_a_20 = a_20;
  assign f_u_arrmul24_and20_14_b_14 = b_14;
  assign f_u_arrmul24_and20_14_y0 = f_u_arrmul24_and20_14_a_20 & f_u_arrmul24_and20_14_b_14;
  assign f_u_arrmul24_fa20_14_f_u_arrmul24_and20_14_y0 = f_u_arrmul24_and20_14_y0;
  assign f_u_arrmul24_fa20_14_f_u_arrmul24_fa21_13_y2 = f_u_arrmul24_fa21_13_y2;
  assign f_u_arrmul24_fa20_14_f_u_arrmul24_fa19_14_y4 = f_u_arrmul24_fa19_14_y4;
  assign f_u_arrmul24_fa20_14_y0 = f_u_arrmul24_fa20_14_f_u_arrmul24_and20_14_y0 ^ f_u_arrmul24_fa20_14_f_u_arrmul24_fa21_13_y2;
  assign f_u_arrmul24_fa20_14_y1 = f_u_arrmul24_fa20_14_f_u_arrmul24_and20_14_y0 & f_u_arrmul24_fa20_14_f_u_arrmul24_fa21_13_y2;
  assign f_u_arrmul24_fa20_14_y2 = f_u_arrmul24_fa20_14_y0 ^ f_u_arrmul24_fa20_14_f_u_arrmul24_fa19_14_y4;
  assign f_u_arrmul24_fa20_14_y3 = f_u_arrmul24_fa20_14_y0 & f_u_arrmul24_fa20_14_f_u_arrmul24_fa19_14_y4;
  assign f_u_arrmul24_fa20_14_y4 = f_u_arrmul24_fa20_14_y1 | f_u_arrmul24_fa20_14_y3;
  assign f_u_arrmul24_and21_14_a_21 = a_21;
  assign f_u_arrmul24_and21_14_b_14 = b_14;
  assign f_u_arrmul24_and21_14_y0 = f_u_arrmul24_and21_14_a_21 & f_u_arrmul24_and21_14_b_14;
  assign f_u_arrmul24_fa21_14_f_u_arrmul24_and21_14_y0 = f_u_arrmul24_and21_14_y0;
  assign f_u_arrmul24_fa21_14_f_u_arrmul24_fa22_13_y2 = f_u_arrmul24_fa22_13_y2;
  assign f_u_arrmul24_fa21_14_f_u_arrmul24_fa20_14_y4 = f_u_arrmul24_fa20_14_y4;
  assign f_u_arrmul24_fa21_14_y0 = f_u_arrmul24_fa21_14_f_u_arrmul24_and21_14_y0 ^ f_u_arrmul24_fa21_14_f_u_arrmul24_fa22_13_y2;
  assign f_u_arrmul24_fa21_14_y1 = f_u_arrmul24_fa21_14_f_u_arrmul24_and21_14_y0 & f_u_arrmul24_fa21_14_f_u_arrmul24_fa22_13_y2;
  assign f_u_arrmul24_fa21_14_y2 = f_u_arrmul24_fa21_14_y0 ^ f_u_arrmul24_fa21_14_f_u_arrmul24_fa20_14_y4;
  assign f_u_arrmul24_fa21_14_y3 = f_u_arrmul24_fa21_14_y0 & f_u_arrmul24_fa21_14_f_u_arrmul24_fa20_14_y4;
  assign f_u_arrmul24_fa21_14_y4 = f_u_arrmul24_fa21_14_y1 | f_u_arrmul24_fa21_14_y3;
  assign f_u_arrmul24_and22_14_a_22 = a_22;
  assign f_u_arrmul24_and22_14_b_14 = b_14;
  assign f_u_arrmul24_and22_14_y0 = f_u_arrmul24_and22_14_a_22 & f_u_arrmul24_and22_14_b_14;
  assign f_u_arrmul24_fa22_14_f_u_arrmul24_and22_14_y0 = f_u_arrmul24_and22_14_y0;
  assign f_u_arrmul24_fa22_14_f_u_arrmul24_fa23_13_y2 = f_u_arrmul24_fa23_13_y2;
  assign f_u_arrmul24_fa22_14_f_u_arrmul24_fa21_14_y4 = f_u_arrmul24_fa21_14_y4;
  assign f_u_arrmul24_fa22_14_y0 = f_u_arrmul24_fa22_14_f_u_arrmul24_and22_14_y0 ^ f_u_arrmul24_fa22_14_f_u_arrmul24_fa23_13_y2;
  assign f_u_arrmul24_fa22_14_y1 = f_u_arrmul24_fa22_14_f_u_arrmul24_and22_14_y0 & f_u_arrmul24_fa22_14_f_u_arrmul24_fa23_13_y2;
  assign f_u_arrmul24_fa22_14_y2 = f_u_arrmul24_fa22_14_y0 ^ f_u_arrmul24_fa22_14_f_u_arrmul24_fa21_14_y4;
  assign f_u_arrmul24_fa22_14_y3 = f_u_arrmul24_fa22_14_y0 & f_u_arrmul24_fa22_14_f_u_arrmul24_fa21_14_y4;
  assign f_u_arrmul24_fa22_14_y4 = f_u_arrmul24_fa22_14_y1 | f_u_arrmul24_fa22_14_y3;
  assign f_u_arrmul24_and23_14_a_23 = a_23;
  assign f_u_arrmul24_and23_14_b_14 = b_14;
  assign f_u_arrmul24_and23_14_y0 = f_u_arrmul24_and23_14_a_23 & f_u_arrmul24_and23_14_b_14;
  assign f_u_arrmul24_fa23_14_f_u_arrmul24_and23_14_y0 = f_u_arrmul24_and23_14_y0;
  assign f_u_arrmul24_fa23_14_f_u_arrmul24_fa23_13_y4 = f_u_arrmul24_fa23_13_y4;
  assign f_u_arrmul24_fa23_14_f_u_arrmul24_fa22_14_y4 = f_u_arrmul24_fa22_14_y4;
  assign f_u_arrmul24_fa23_14_y0 = f_u_arrmul24_fa23_14_f_u_arrmul24_and23_14_y0 ^ f_u_arrmul24_fa23_14_f_u_arrmul24_fa23_13_y4;
  assign f_u_arrmul24_fa23_14_y1 = f_u_arrmul24_fa23_14_f_u_arrmul24_and23_14_y0 & f_u_arrmul24_fa23_14_f_u_arrmul24_fa23_13_y4;
  assign f_u_arrmul24_fa23_14_y2 = f_u_arrmul24_fa23_14_y0 ^ f_u_arrmul24_fa23_14_f_u_arrmul24_fa22_14_y4;
  assign f_u_arrmul24_fa23_14_y3 = f_u_arrmul24_fa23_14_y0 & f_u_arrmul24_fa23_14_f_u_arrmul24_fa22_14_y4;
  assign f_u_arrmul24_fa23_14_y4 = f_u_arrmul24_fa23_14_y1 | f_u_arrmul24_fa23_14_y3;
  assign f_u_arrmul24_and0_15_a_0 = a_0;
  assign f_u_arrmul24_and0_15_b_15 = b_15;
  assign f_u_arrmul24_and0_15_y0 = f_u_arrmul24_and0_15_a_0 & f_u_arrmul24_and0_15_b_15;
  assign f_u_arrmul24_ha0_15_f_u_arrmul24_and0_15_y0 = f_u_arrmul24_and0_15_y0;
  assign f_u_arrmul24_ha0_15_f_u_arrmul24_fa1_14_y2 = f_u_arrmul24_fa1_14_y2;
  assign f_u_arrmul24_ha0_15_y0 = f_u_arrmul24_ha0_15_f_u_arrmul24_and0_15_y0 ^ f_u_arrmul24_ha0_15_f_u_arrmul24_fa1_14_y2;
  assign f_u_arrmul24_ha0_15_y1 = f_u_arrmul24_ha0_15_f_u_arrmul24_and0_15_y0 & f_u_arrmul24_ha0_15_f_u_arrmul24_fa1_14_y2;
  assign f_u_arrmul24_and1_15_a_1 = a_1;
  assign f_u_arrmul24_and1_15_b_15 = b_15;
  assign f_u_arrmul24_and1_15_y0 = f_u_arrmul24_and1_15_a_1 & f_u_arrmul24_and1_15_b_15;
  assign f_u_arrmul24_fa1_15_f_u_arrmul24_and1_15_y0 = f_u_arrmul24_and1_15_y0;
  assign f_u_arrmul24_fa1_15_f_u_arrmul24_fa2_14_y2 = f_u_arrmul24_fa2_14_y2;
  assign f_u_arrmul24_fa1_15_f_u_arrmul24_ha0_15_y1 = f_u_arrmul24_ha0_15_y1;
  assign f_u_arrmul24_fa1_15_y0 = f_u_arrmul24_fa1_15_f_u_arrmul24_and1_15_y0 ^ f_u_arrmul24_fa1_15_f_u_arrmul24_fa2_14_y2;
  assign f_u_arrmul24_fa1_15_y1 = f_u_arrmul24_fa1_15_f_u_arrmul24_and1_15_y0 & f_u_arrmul24_fa1_15_f_u_arrmul24_fa2_14_y2;
  assign f_u_arrmul24_fa1_15_y2 = f_u_arrmul24_fa1_15_y0 ^ f_u_arrmul24_fa1_15_f_u_arrmul24_ha0_15_y1;
  assign f_u_arrmul24_fa1_15_y3 = f_u_arrmul24_fa1_15_y0 & f_u_arrmul24_fa1_15_f_u_arrmul24_ha0_15_y1;
  assign f_u_arrmul24_fa1_15_y4 = f_u_arrmul24_fa1_15_y1 | f_u_arrmul24_fa1_15_y3;
  assign f_u_arrmul24_and2_15_a_2 = a_2;
  assign f_u_arrmul24_and2_15_b_15 = b_15;
  assign f_u_arrmul24_and2_15_y0 = f_u_arrmul24_and2_15_a_2 & f_u_arrmul24_and2_15_b_15;
  assign f_u_arrmul24_fa2_15_f_u_arrmul24_and2_15_y0 = f_u_arrmul24_and2_15_y0;
  assign f_u_arrmul24_fa2_15_f_u_arrmul24_fa3_14_y2 = f_u_arrmul24_fa3_14_y2;
  assign f_u_arrmul24_fa2_15_f_u_arrmul24_fa1_15_y4 = f_u_arrmul24_fa1_15_y4;
  assign f_u_arrmul24_fa2_15_y0 = f_u_arrmul24_fa2_15_f_u_arrmul24_and2_15_y0 ^ f_u_arrmul24_fa2_15_f_u_arrmul24_fa3_14_y2;
  assign f_u_arrmul24_fa2_15_y1 = f_u_arrmul24_fa2_15_f_u_arrmul24_and2_15_y0 & f_u_arrmul24_fa2_15_f_u_arrmul24_fa3_14_y2;
  assign f_u_arrmul24_fa2_15_y2 = f_u_arrmul24_fa2_15_y0 ^ f_u_arrmul24_fa2_15_f_u_arrmul24_fa1_15_y4;
  assign f_u_arrmul24_fa2_15_y3 = f_u_arrmul24_fa2_15_y0 & f_u_arrmul24_fa2_15_f_u_arrmul24_fa1_15_y4;
  assign f_u_arrmul24_fa2_15_y4 = f_u_arrmul24_fa2_15_y1 | f_u_arrmul24_fa2_15_y3;
  assign f_u_arrmul24_and3_15_a_3 = a_3;
  assign f_u_arrmul24_and3_15_b_15 = b_15;
  assign f_u_arrmul24_and3_15_y0 = f_u_arrmul24_and3_15_a_3 & f_u_arrmul24_and3_15_b_15;
  assign f_u_arrmul24_fa3_15_f_u_arrmul24_and3_15_y0 = f_u_arrmul24_and3_15_y0;
  assign f_u_arrmul24_fa3_15_f_u_arrmul24_fa4_14_y2 = f_u_arrmul24_fa4_14_y2;
  assign f_u_arrmul24_fa3_15_f_u_arrmul24_fa2_15_y4 = f_u_arrmul24_fa2_15_y4;
  assign f_u_arrmul24_fa3_15_y0 = f_u_arrmul24_fa3_15_f_u_arrmul24_and3_15_y0 ^ f_u_arrmul24_fa3_15_f_u_arrmul24_fa4_14_y2;
  assign f_u_arrmul24_fa3_15_y1 = f_u_arrmul24_fa3_15_f_u_arrmul24_and3_15_y0 & f_u_arrmul24_fa3_15_f_u_arrmul24_fa4_14_y2;
  assign f_u_arrmul24_fa3_15_y2 = f_u_arrmul24_fa3_15_y0 ^ f_u_arrmul24_fa3_15_f_u_arrmul24_fa2_15_y4;
  assign f_u_arrmul24_fa3_15_y3 = f_u_arrmul24_fa3_15_y0 & f_u_arrmul24_fa3_15_f_u_arrmul24_fa2_15_y4;
  assign f_u_arrmul24_fa3_15_y4 = f_u_arrmul24_fa3_15_y1 | f_u_arrmul24_fa3_15_y3;
  assign f_u_arrmul24_and4_15_a_4 = a_4;
  assign f_u_arrmul24_and4_15_b_15 = b_15;
  assign f_u_arrmul24_and4_15_y0 = f_u_arrmul24_and4_15_a_4 & f_u_arrmul24_and4_15_b_15;
  assign f_u_arrmul24_fa4_15_f_u_arrmul24_and4_15_y0 = f_u_arrmul24_and4_15_y0;
  assign f_u_arrmul24_fa4_15_f_u_arrmul24_fa5_14_y2 = f_u_arrmul24_fa5_14_y2;
  assign f_u_arrmul24_fa4_15_f_u_arrmul24_fa3_15_y4 = f_u_arrmul24_fa3_15_y4;
  assign f_u_arrmul24_fa4_15_y0 = f_u_arrmul24_fa4_15_f_u_arrmul24_and4_15_y0 ^ f_u_arrmul24_fa4_15_f_u_arrmul24_fa5_14_y2;
  assign f_u_arrmul24_fa4_15_y1 = f_u_arrmul24_fa4_15_f_u_arrmul24_and4_15_y0 & f_u_arrmul24_fa4_15_f_u_arrmul24_fa5_14_y2;
  assign f_u_arrmul24_fa4_15_y2 = f_u_arrmul24_fa4_15_y0 ^ f_u_arrmul24_fa4_15_f_u_arrmul24_fa3_15_y4;
  assign f_u_arrmul24_fa4_15_y3 = f_u_arrmul24_fa4_15_y0 & f_u_arrmul24_fa4_15_f_u_arrmul24_fa3_15_y4;
  assign f_u_arrmul24_fa4_15_y4 = f_u_arrmul24_fa4_15_y1 | f_u_arrmul24_fa4_15_y3;
  assign f_u_arrmul24_and5_15_a_5 = a_5;
  assign f_u_arrmul24_and5_15_b_15 = b_15;
  assign f_u_arrmul24_and5_15_y0 = f_u_arrmul24_and5_15_a_5 & f_u_arrmul24_and5_15_b_15;
  assign f_u_arrmul24_fa5_15_f_u_arrmul24_and5_15_y0 = f_u_arrmul24_and5_15_y0;
  assign f_u_arrmul24_fa5_15_f_u_arrmul24_fa6_14_y2 = f_u_arrmul24_fa6_14_y2;
  assign f_u_arrmul24_fa5_15_f_u_arrmul24_fa4_15_y4 = f_u_arrmul24_fa4_15_y4;
  assign f_u_arrmul24_fa5_15_y0 = f_u_arrmul24_fa5_15_f_u_arrmul24_and5_15_y0 ^ f_u_arrmul24_fa5_15_f_u_arrmul24_fa6_14_y2;
  assign f_u_arrmul24_fa5_15_y1 = f_u_arrmul24_fa5_15_f_u_arrmul24_and5_15_y0 & f_u_arrmul24_fa5_15_f_u_arrmul24_fa6_14_y2;
  assign f_u_arrmul24_fa5_15_y2 = f_u_arrmul24_fa5_15_y0 ^ f_u_arrmul24_fa5_15_f_u_arrmul24_fa4_15_y4;
  assign f_u_arrmul24_fa5_15_y3 = f_u_arrmul24_fa5_15_y0 & f_u_arrmul24_fa5_15_f_u_arrmul24_fa4_15_y4;
  assign f_u_arrmul24_fa5_15_y4 = f_u_arrmul24_fa5_15_y1 | f_u_arrmul24_fa5_15_y3;
  assign f_u_arrmul24_and6_15_a_6 = a_6;
  assign f_u_arrmul24_and6_15_b_15 = b_15;
  assign f_u_arrmul24_and6_15_y0 = f_u_arrmul24_and6_15_a_6 & f_u_arrmul24_and6_15_b_15;
  assign f_u_arrmul24_fa6_15_f_u_arrmul24_and6_15_y0 = f_u_arrmul24_and6_15_y0;
  assign f_u_arrmul24_fa6_15_f_u_arrmul24_fa7_14_y2 = f_u_arrmul24_fa7_14_y2;
  assign f_u_arrmul24_fa6_15_f_u_arrmul24_fa5_15_y4 = f_u_arrmul24_fa5_15_y4;
  assign f_u_arrmul24_fa6_15_y0 = f_u_arrmul24_fa6_15_f_u_arrmul24_and6_15_y0 ^ f_u_arrmul24_fa6_15_f_u_arrmul24_fa7_14_y2;
  assign f_u_arrmul24_fa6_15_y1 = f_u_arrmul24_fa6_15_f_u_arrmul24_and6_15_y0 & f_u_arrmul24_fa6_15_f_u_arrmul24_fa7_14_y2;
  assign f_u_arrmul24_fa6_15_y2 = f_u_arrmul24_fa6_15_y0 ^ f_u_arrmul24_fa6_15_f_u_arrmul24_fa5_15_y4;
  assign f_u_arrmul24_fa6_15_y3 = f_u_arrmul24_fa6_15_y0 & f_u_arrmul24_fa6_15_f_u_arrmul24_fa5_15_y4;
  assign f_u_arrmul24_fa6_15_y4 = f_u_arrmul24_fa6_15_y1 | f_u_arrmul24_fa6_15_y3;
  assign f_u_arrmul24_and7_15_a_7 = a_7;
  assign f_u_arrmul24_and7_15_b_15 = b_15;
  assign f_u_arrmul24_and7_15_y0 = f_u_arrmul24_and7_15_a_7 & f_u_arrmul24_and7_15_b_15;
  assign f_u_arrmul24_fa7_15_f_u_arrmul24_and7_15_y0 = f_u_arrmul24_and7_15_y0;
  assign f_u_arrmul24_fa7_15_f_u_arrmul24_fa8_14_y2 = f_u_arrmul24_fa8_14_y2;
  assign f_u_arrmul24_fa7_15_f_u_arrmul24_fa6_15_y4 = f_u_arrmul24_fa6_15_y4;
  assign f_u_arrmul24_fa7_15_y0 = f_u_arrmul24_fa7_15_f_u_arrmul24_and7_15_y0 ^ f_u_arrmul24_fa7_15_f_u_arrmul24_fa8_14_y2;
  assign f_u_arrmul24_fa7_15_y1 = f_u_arrmul24_fa7_15_f_u_arrmul24_and7_15_y0 & f_u_arrmul24_fa7_15_f_u_arrmul24_fa8_14_y2;
  assign f_u_arrmul24_fa7_15_y2 = f_u_arrmul24_fa7_15_y0 ^ f_u_arrmul24_fa7_15_f_u_arrmul24_fa6_15_y4;
  assign f_u_arrmul24_fa7_15_y3 = f_u_arrmul24_fa7_15_y0 & f_u_arrmul24_fa7_15_f_u_arrmul24_fa6_15_y4;
  assign f_u_arrmul24_fa7_15_y4 = f_u_arrmul24_fa7_15_y1 | f_u_arrmul24_fa7_15_y3;
  assign f_u_arrmul24_and8_15_a_8 = a_8;
  assign f_u_arrmul24_and8_15_b_15 = b_15;
  assign f_u_arrmul24_and8_15_y0 = f_u_arrmul24_and8_15_a_8 & f_u_arrmul24_and8_15_b_15;
  assign f_u_arrmul24_fa8_15_f_u_arrmul24_and8_15_y0 = f_u_arrmul24_and8_15_y0;
  assign f_u_arrmul24_fa8_15_f_u_arrmul24_fa9_14_y2 = f_u_arrmul24_fa9_14_y2;
  assign f_u_arrmul24_fa8_15_f_u_arrmul24_fa7_15_y4 = f_u_arrmul24_fa7_15_y4;
  assign f_u_arrmul24_fa8_15_y0 = f_u_arrmul24_fa8_15_f_u_arrmul24_and8_15_y0 ^ f_u_arrmul24_fa8_15_f_u_arrmul24_fa9_14_y2;
  assign f_u_arrmul24_fa8_15_y1 = f_u_arrmul24_fa8_15_f_u_arrmul24_and8_15_y0 & f_u_arrmul24_fa8_15_f_u_arrmul24_fa9_14_y2;
  assign f_u_arrmul24_fa8_15_y2 = f_u_arrmul24_fa8_15_y0 ^ f_u_arrmul24_fa8_15_f_u_arrmul24_fa7_15_y4;
  assign f_u_arrmul24_fa8_15_y3 = f_u_arrmul24_fa8_15_y0 & f_u_arrmul24_fa8_15_f_u_arrmul24_fa7_15_y4;
  assign f_u_arrmul24_fa8_15_y4 = f_u_arrmul24_fa8_15_y1 | f_u_arrmul24_fa8_15_y3;
  assign f_u_arrmul24_and9_15_a_9 = a_9;
  assign f_u_arrmul24_and9_15_b_15 = b_15;
  assign f_u_arrmul24_and9_15_y0 = f_u_arrmul24_and9_15_a_9 & f_u_arrmul24_and9_15_b_15;
  assign f_u_arrmul24_fa9_15_f_u_arrmul24_and9_15_y0 = f_u_arrmul24_and9_15_y0;
  assign f_u_arrmul24_fa9_15_f_u_arrmul24_fa10_14_y2 = f_u_arrmul24_fa10_14_y2;
  assign f_u_arrmul24_fa9_15_f_u_arrmul24_fa8_15_y4 = f_u_arrmul24_fa8_15_y4;
  assign f_u_arrmul24_fa9_15_y0 = f_u_arrmul24_fa9_15_f_u_arrmul24_and9_15_y0 ^ f_u_arrmul24_fa9_15_f_u_arrmul24_fa10_14_y2;
  assign f_u_arrmul24_fa9_15_y1 = f_u_arrmul24_fa9_15_f_u_arrmul24_and9_15_y0 & f_u_arrmul24_fa9_15_f_u_arrmul24_fa10_14_y2;
  assign f_u_arrmul24_fa9_15_y2 = f_u_arrmul24_fa9_15_y0 ^ f_u_arrmul24_fa9_15_f_u_arrmul24_fa8_15_y4;
  assign f_u_arrmul24_fa9_15_y3 = f_u_arrmul24_fa9_15_y0 & f_u_arrmul24_fa9_15_f_u_arrmul24_fa8_15_y4;
  assign f_u_arrmul24_fa9_15_y4 = f_u_arrmul24_fa9_15_y1 | f_u_arrmul24_fa9_15_y3;
  assign f_u_arrmul24_and10_15_a_10 = a_10;
  assign f_u_arrmul24_and10_15_b_15 = b_15;
  assign f_u_arrmul24_and10_15_y0 = f_u_arrmul24_and10_15_a_10 & f_u_arrmul24_and10_15_b_15;
  assign f_u_arrmul24_fa10_15_f_u_arrmul24_and10_15_y0 = f_u_arrmul24_and10_15_y0;
  assign f_u_arrmul24_fa10_15_f_u_arrmul24_fa11_14_y2 = f_u_arrmul24_fa11_14_y2;
  assign f_u_arrmul24_fa10_15_f_u_arrmul24_fa9_15_y4 = f_u_arrmul24_fa9_15_y4;
  assign f_u_arrmul24_fa10_15_y0 = f_u_arrmul24_fa10_15_f_u_arrmul24_and10_15_y0 ^ f_u_arrmul24_fa10_15_f_u_arrmul24_fa11_14_y2;
  assign f_u_arrmul24_fa10_15_y1 = f_u_arrmul24_fa10_15_f_u_arrmul24_and10_15_y0 & f_u_arrmul24_fa10_15_f_u_arrmul24_fa11_14_y2;
  assign f_u_arrmul24_fa10_15_y2 = f_u_arrmul24_fa10_15_y0 ^ f_u_arrmul24_fa10_15_f_u_arrmul24_fa9_15_y4;
  assign f_u_arrmul24_fa10_15_y3 = f_u_arrmul24_fa10_15_y0 & f_u_arrmul24_fa10_15_f_u_arrmul24_fa9_15_y4;
  assign f_u_arrmul24_fa10_15_y4 = f_u_arrmul24_fa10_15_y1 | f_u_arrmul24_fa10_15_y3;
  assign f_u_arrmul24_and11_15_a_11 = a_11;
  assign f_u_arrmul24_and11_15_b_15 = b_15;
  assign f_u_arrmul24_and11_15_y0 = f_u_arrmul24_and11_15_a_11 & f_u_arrmul24_and11_15_b_15;
  assign f_u_arrmul24_fa11_15_f_u_arrmul24_and11_15_y0 = f_u_arrmul24_and11_15_y0;
  assign f_u_arrmul24_fa11_15_f_u_arrmul24_fa12_14_y2 = f_u_arrmul24_fa12_14_y2;
  assign f_u_arrmul24_fa11_15_f_u_arrmul24_fa10_15_y4 = f_u_arrmul24_fa10_15_y4;
  assign f_u_arrmul24_fa11_15_y0 = f_u_arrmul24_fa11_15_f_u_arrmul24_and11_15_y0 ^ f_u_arrmul24_fa11_15_f_u_arrmul24_fa12_14_y2;
  assign f_u_arrmul24_fa11_15_y1 = f_u_arrmul24_fa11_15_f_u_arrmul24_and11_15_y0 & f_u_arrmul24_fa11_15_f_u_arrmul24_fa12_14_y2;
  assign f_u_arrmul24_fa11_15_y2 = f_u_arrmul24_fa11_15_y0 ^ f_u_arrmul24_fa11_15_f_u_arrmul24_fa10_15_y4;
  assign f_u_arrmul24_fa11_15_y3 = f_u_arrmul24_fa11_15_y0 & f_u_arrmul24_fa11_15_f_u_arrmul24_fa10_15_y4;
  assign f_u_arrmul24_fa11_15_y4 = f_u_arrmul24_fa11_15_y1 | f_u_arrmul24_fa11_15_y3;
  assign f_u_arrmul24_and12_15_a_12 = a_12;
  assign f_u_arrmul24_and12_15_b_15 = b_15;
  assign f_u_arrmul24_and12_15_y0 = f_u_arrmul24_and12_15_a_12 & f_u_arrmul24_and12_15_b_15;
  assign f_u_arrmul24_fa12_15_f_u_arrmul24_and12_15_y0 = f_u_arrmul24_and12_15_y0;
  assign f_u_arrmul24_fa12_15_f_u_arrmul24_fa13_14_y2 = f_u_arrmul24_fa13_14_y2;
  assign f_u_arrmul24_fa12_15_f_u_arrmul24_fa11_15_y4 = f_u_arrmul24_fa11_15_y4;
  assign f_u_arrmul24_fa12_15_y0 = f_u_arrmul24_fa12_15_f_u_arrmul24_and12_15_y0 ^ f_u_arrmul24_fa12_15_f_u_arrmul24_fa13_14_y2;
  assign f_u_arrmul24_fa12_15_y1 = f_u_arrmul24_fa12_15_f_u_arrmul24_and12_15_y0 & f_u_arrmul24_fa12_15_f_u_arrmul24_fa13_14_y2;
  assign f_u_arrmul24_fa12_15_y2 = f_u_arrmul24_fa12_15_y0 ^ f_u_arrmul24_fa12_15_f_u_arrmul24_fa11_15_y4;
  assign f_u_arrmul24_fa12_15_y3 = f_u_arrmul24_fa12_15_y0 & f_u_arrmul24_fa12_15_f_u_arrmul24_fa11_15_y4;
  assign f_u_arrmul24_fa12_15_y4 = f_u_arrmul24_fa12_15_y1 | f_u_arrmul24_fa12_15_y3;
  assign f_u_arrmul24_and13_15_a_13 = a_13;
  assign f_u_arrmul24_and13_15_b_15 = b_15;
  assign f_u_arrmul24_and13_15_y0 = f_u_arrmul24_and13_15_a_13 & f_u_arrmul24_and13_15_b_15;
  assign f_u_arrmul24_fa13_15_f_u_arrmul24_and13_15_y0 = f_u_arrmul24_and13_15_y0;
  assign f_u_arrmul24_fa13_15_f_u_arrmul24_fa14_14_y2 = f_u_arrmul24_fa14_14_y2;
  assign f_u_arrmul24_fa13_15_f_u_arrmul24_fa12_15_y4 = f_u_arrmul24_fa12_15_y4;
  assign f_u_arrmul24_fa13_15_y0 = f_u_arrmul24_fa13_15_f_u_arrmul24_and13_15_y0 ^ f_u_arrmul24_fa13_15_f_u_arrmul24_fa14_14_y2;
  assign f_u_arrmul24_fa13_15_y1 = f_u_arrmul24_fa13_15_f_u_arrmul24_and13_15_y0 & f_u_arrmul24_fa13_15_f_u_arrmul24_fa14_14_y2;
  assign f_u_arrmul24_fa13_15_y2 = f_u_arrmul24_fa13_15_y0 ^ f_u_arrmul24_fa13_15_f_u_arrmul24_fa12_15_y4;
  assign f_u_arrmul24_fa13_15_y3 = f_u_arrmul24_fa13_15_y0 & f_u_arrmul24_fa13_15_f_u_arrmul24_fa12_15_y4;
  assign f_u_arrmul24_fa13_15_y4 = f_u_arrmul24_fa13_15_y1 | f_u_arrmul24_fa13_15_y3;
  assign f_u_arrmul24_and14_15_a_14 = a_14;
  assign f_u_arrmul24_and14_15_b_15 = b_15;
  assign f_u_arrmul24_and14_15_y0 = f_u_arrmul24_and14_15_a_14 & f_u_arrmul24_and14_15_b_15;
  assign f_u_arrmul24_fa14_15_f_u_arrmul24_and14_15_y0 = f_u_arrmul24_and14_15_y0;
  assign f_u_arrmul24_fa14_15_f_u_arrmul24_fa15_14_y2 = f_u_arrmul24_fa15_14_y2;
  assign f_u_arrmul24_fa14_15_f_u_arrmul24_fa13_15_y4 = f_u_arrmul24_fa13_15_y4;
  assign f_u_arrmul24_fa14_15_y0 = f_u_arrmul24_fa14_15_f_u_arrmul24_and14_15_y0 ^ f_u_arrmul24_fa14_15_f_u_arrmul24_fa15_14_y2;
  assign f_u_arrmul24_fa14_15_y1 = f_u_arrmul24_fa14_15_f_u_arrmul24_and14_15_y0 & f_u_arrmul24_fa14_15_f_u_arrmul24_fa15_14_y2;
  assign f_u_arrmul24_fa14_15_y2 = f_u_arrmul24_fa14_15_y0 ^ f_u_arrmul24_fa14_15_f_u_arrmul24_fa13_15_y4;
  assign f_u_arrmul24_fa14_15_y3 = f_u_arrmul24_fa14_15_y0 & f_u_arrmul24_fa14_15_f_u_arrmul24_fa13_15_y4;
  assign f_u_arrmul24_fa14_15_y4 = f_u_arrmul24_fa14_15_y1 | f_u_arrmul24_fa14_15_y3;
  assign f_u_arrmul24_and15_15_a_15 = a_15;
  assign f_u_arrmul24_and15_15_b_15 = b_15;
  assign f_u_arrmul24_and15_15_y0 = f_u_arrmul24_and15_15_a_15 & f_u_arrmul24_and15_15_b_15;
  assign f_u_arrmul24_fa15_15_f_u_arrmul24_and15_15_y0 = f_u_arrmul24_and15_15_y0;
  assign f_u_arrmul24_fa15_15_f_u_arrmul24_fa16_14_y2 = f_u_arrmul24_fa16_14_y2;
  assign f_u_arrmul24_fa15_15_f_u_arrmul24_fa14_15_y4 = f_u_arrmul24_fa14_15_y4;
  assign f_u_arrmul24_fa15_15_y0 = f_u_arrmul24_fa15_15_f_u_arrmul24_and15_15_y0 ^ f_u_arrmul24_fa15_15_f_u_arrmul24_fa16_14_y2;
  assign f_u_arrmul24_fa15_15_y1 = f_u_arrmul24_fa15_15_f_u_arrmul24_and15_15_y0 & f_u_arrmul24_fa15_15_f_u_arrmul24_fa16_14_y2;
  assign f_u_arrmul24_fa15_15_y2 = f_u_arrmul24_fa15_15_y0 ^ f_u_arrmul24_fa15_15_f_u_arrmul24_fa14_15_y4;
  assign f_u_arrmul24_fa15_15_y3 = f_u_arrmul24_fa15_15_y0 & f_u_arrmul24_fa15_15_f_u_arrmul24_fa14_15_y4;
  assign f_u_arrmul24_fa15_15_y4 = f_u_arrmul24_fa15_15_y1 | f_u_arrmul24_fa15_15_y3;
  assign f_u_arrmul24_and16_15_a_16 = a_16;
  assign f_u_arrmul24_and16_15_b_15 = b_15;
  assign f_u_arrmul24_and16_15_y0 = f_u_arrmul24_and16_15_a_16 & f_u_arrmul24_and16_15_b_15;
  assign f_u_arrmul24_fa16_15_f_u_arrmul24_and16_15_y0 = f_u_arrmul24_and16_15_y0;
  assign f_u_arrmul24_fa16_15_f_u_arrmul24_fa17_14_y2 = f_u_arrmul24_fa17_14_y2;
  assign f_u_arrmul24_fa16_15_f_u_arrmul24_fa15_15_y4 = f_u_arrmul24_fa15_15_y4;
  assign f_u_arrmul24_fa16_15_y0 = f_u_arrmul24_fa16_15_f_u_arrmul24_and16_15_y0 ^ f_u_arrmul24_fa16_15_f_u_arrmul24_fa17_14_y2;
  assign f_u_arrmul24_fa16_15_y1 = f_u_arrmul24_fa16_15_f_u_arrmul24_and16_15_y0 & f_u_arrmul24_fa16_15_f_u_arrmul24_fa17_14_y2;
  assign f_u_arrmul24_fa16_15_y2 = f_u_arrmul24_fa16_15_y0 ^ f_u_arrmul24_fa16_15_f_u_arrmul24_fa15_15_y4;
  assign f_u_arrmul24_fa16_15_y3 = f_u_arrmul24_fa16_15_y0 & f_u_arrmul24_fa16_15_f_u_arrmul24_fa15_15_y4;
  assign f_u_arrmul24_fa16_15_y4 = f_u_arrmul24_fa16_15_y1 | f_u_arrmul24_fa16_15_y3;
  assign f_u_arrmul24_and17_15_a_17 = a_17;
  assign f_u_arrmul24_and17_15_b_15 = b_15;
  assign f_u_arrmul24_and17_15_y0 = f_u_arrmul24_and17_15_a_17 & f_u_arrmul24_and17_15_b_15;
  assign f_u_arrmul24_fa17_15_f_u_arrmul24_and17_15_y0 = f_u_arrmul24_and17_15_y0;
  assign f_u_arrmul24_fa17_15_f_u_arrmul24_fa18_14_y2 = f_u_arrmul24_fa18_14_y2;
  assign f_u_arrmul24_fa17_15_f_u_arrmul24_fa16_15_y4 = f_u_arrmul24_fa16_15_y4;
  assign f_u_arrmul24_fa17_15_y0 = f_u_arrmul24_fa17_15_f_u_arrmul24_and17_15_y0 ^ f_u_arrmul24_fa17_15_f_u_arrmul24_fa18_14_y2;
  assign f_u_arrmul24_fa17_15_y1 = f_u_arrmul24_fa17_15_f_u_arrmul24_and17_15_y0 & f_u_arrmul24_fa17_15_f_u_arrmul24_fa18_14_y2;
  assign f_u_arrmul24_fa17_15_y2 = f_u_arrmul24_fa17_15_y0 ^ f_u_arrmul24_fa17_15_f_u_arrmul24_fa16_15_y4;
  assign f_u_arrmul24_fa17_15_y3 = f_u_arrmul24_fa17_15_y0 & f_u_arrmul24_fa17_15_f_u_arrmul24_fa16_15_y4;
  assign f_u_arrmul24_fa17_15_y4 = f_u_arrmul24_fa17_15_y1 | f_u_arrmul24_fa17_15_y3;
  assign f_u_arrmul24_and18_15_a_18 = a_18;
  assign f_u_arrmul24_and18_15_b_15 = b_15;
  assign f_u_arrmul24_and18_15_y0 = f_u_arrmul24_and18_15_a_18 & f_u_arrmul24_and18_15_b_15;
  assign f_u_arrmul24_fa18_15_f_u_arrmul24_and18_15_y0 = f_u_arrmul24_and18_15_y0;
  assign f_u_arrmul24_fa18_15_f_u_arrmul24_fa19_14_y2 = f_u_arrmul24_fa19_14_y2;
  assign f_u_arrmul24_fa18_15_f_u_arrmul24_fa17_15_y4 = f_u_arrmul24_fa17_15_y4;
  assign f_u_arrmul24_fa18_15_y0 = f_u_arrmul24_fa18_15_f_u_arrmul24_and18_15_y0 ^ f_u_arrmul24_fa18_15_f_u_arrmul24_fa19_14_y2;
  assign f_u_arrmul24_fa18_15_y1 = f_u_arrmul24_fa18_15_f_u_arrmul24_and18_15_y0 & f_u_arrmul24_fa18_15_f_u_arrmul24_fa19_14_y2;
  assign f_u_arrmul24_fa18_15_y2 = f_u_arrmul24_fa18_15_y0 ^ f_u_arrmul24_fa18_15_f_u_arrmul24_fa17_15_y4;
  assign f_u_arrmul24_fa18_15_y3 = f_u_arrmul24_fa18_15_y0 & f_u_arrmul24_fa18_15_f_u_arrmul24_fa17_15_y4;
  assign f_u_arrmul24_fa18_15_y4 = f_u_arrmul24_fa18_15_y1 | f_u_arrmul24_fa18_15_y3;
  assign f_u_arrmul24_and19_15_a_19 = a_19;
  assign f_u_arrmul24_and19_15_b_15 = b_15;
  assign f_u_arrmul24_and19_15_y0 = f_u_arrmul24_and19_15_a_19 & f_u_arrmul24_and19_15_b_15;
  assign f_u_arrmul24_fa19_15_f_u_arrmul24_and19_15_y0 = f_u_arrmul24_and19_15_y0;
  assign f_u_arrmul24_fa19_15_f_u_arrmul24_fa20_14_y2 = f_u_arrmul24_fa20_14_y2;
  assign f_u_arrmul24_fa19_15_f_u_arrmul24_fa18_15_y4 = f_u_arrmul24_fa18_15_y4;
  assign f_u_arrmul24_fa19_15_y0 = f_u_arrmul24_fa19_15_f_u_arrmul24_and19_15_y0 ^ f_u_arrmul24_fa19_15_f_u_arrmul24_fa20_14_y2;
  assign f_u_arrmul24_fa19_15_y1 = f_u_arrmul24_fa19_15_f_u_arrmul24_and19_15_y0 & f_u_arrmul24_fa19_15_f_u_arrmul24_fa20_14_y2;
  assign f_u_arrmul24_fa19_15_y2 = f_u_arrmul24_fa19_15_y0 ^ f_u_arrmul24_fa19_15_f_u_arrmul24_fa18_15_y4;
  assign f_u_arrmul24_fa19_15_y3 = f_u_arrmul24_fa19_15_y0 & f_u_arrmul24_fa19_15_f_u_arrmul24_fa18_15_y4;
  assign f_u_arrmul24_fa19_15_y4 = f_u_arrmul24_fa19_15_y1 | f_u_arrmul24_fa19_15_y3;
  assign f_u_arrmul24_and20_15_a_20 = a_20;
  assign f_u_arrmul24_and20_15_b_15 = b_15;
  assign f_u_arrmul24_and20_15_y0 = f_u_arrmul24_and20_15_a_20 & f_u_arrmul24_and20_15_b_15;
  assign f_u_arrmul24_fa20_15_f_u_arrmul24_and20_15_y0 = f_u_arrmul24_and20_15_y0;
  assign f_u_arrmul24_fa20_15_f_u_arrmul24_fa21_14_y2 = f_u_arrmul24_fa21_14_y2;
  assign f_u_arrmul24_fa20_15_f_u_arrmul24_fa19_15_y4 = f_u_arrmul24_fa19_15_y4;
  assign f_u_arrmul24_fa20_15_y0 = f_u_arrmul24_fa20_15_f_u_arrmul24_and20_15_y0 ^ f_u_arrmul24_fa20_15_f_u_arrmul24_fa21_14_y2;
  assign f_u_arrmul24_fa20_15_y1 = f_u_arrmul24_fa20_15_f_u_arrmul24_and20_15_y0 & f_u_arrmul24_fa20_15_f_u_arrmul24_fa21_14_y2;
  assign f_u_arrmul24_fa20_15_y2 = f_u_arrmul24_fa20_15_y0 ^ f_u_arrmul24_fa20_15_f_u_arrmul24_fa19_15_y4;
  assign f_u_arrmul24_fa20_15_y3 = f_u_arrmul24_fa20_15_y0 & f_u_arrmul24_fa20_15_f_u_arrmul24_fa19_15_y4;
  assign f_u_arrmul24_fa20_15_y4 = f_u_arrmul24_fa20_15_y1 | f_u_arrmul24_fa20_15_y3;
  assign f_u_arrmul24_and21_15_a_21 = a_21;
  assign f_u_arrmul24_and21_15_b_15 = b_15;
  assign f_u_arrmul24_and21_15_y0 = f_u_arrmul24_and21_15_a_21 & f_u_arrmul24_and21_15_b_15;
  assign f_u_arrmul24_fa21_15_f_u_arrmul24_and21_15_y0 = f_u_arrmul24_and21_15_y0;
  assign f_u_arrmul24_fa21_15_f_u_arrmul24_fa22_14_y2 = f_u_arrmul24_fa22_14_y2;
  assign f_u_arrmul24_fa21_15_f_u_arrmul24_fa20_15_y4 = f_u_arrmul24_fa20_15_y4;
  assign f_u_arrmul24_fa21_15_y0 = f_u_arrmul24_fa21_15_f_u_arrmul24_and21_15_y0 ^ f_u_arrmul24_fa21_15_f_u_arrmul24_fa22_14_y2;
  assign f_u_arrmul24_fa21_15_y1 = f_u_arrmul24_fa21_15_f_u_arrmul24_and21_15_y0 & f_u_arrmul24_fa21_15_f_u_arrmul24_fa22_14_y2;
  assign f_u_arrmul24_fa21_15_y2 = f_u_arrmul24_fa21_15_y0 ^ f_u_arrmul24_fa21_15_f_u_arrmul24_fa20_15_y4;
  assign f_u_arrmul24_fa21_15_y3 = f_u_arrmul24_fa21_15_y0 & f_u_arrmul24_fa21_15_f_u_arrmul24_fa20_15_y4;
  assign f_u_arrmul24_fa21_15_y4 = f_u_arrmul24_fa21_15_y1 | f_u_arrmul24_fa21_15_y3;
  assign f_u_arrmul24_and22_15_a_22 = a_22;
  assign f_u_arrmul24_and22_15_b_15 = b_15;
  assign f_u_arrmul24_and22_15_y0 = f_u_arrmul24_and22_15_a_22 & f_u_arrmul24_and22_15_b_15;
  assign f_u_arrmul24_fa22_15_f_u_arrmul24_and22_15_y0 = f_u_arrmul24_and22_15_y0;
  assign f_u_arrmul24_fa22_15_f_u_arrmul24_fa23_14_y2 = f_u_arrmul24_fa23_14_y2;
  assign f_u_arrmul24_fa22_15_f_u_arrmul24_fa21_15_y4 = f_u_arrmul24_fa21_15_y4;
  assign f_u_arrmul24_fa22_15_y0 = f_u_arrmul24_fa22_15_f_u_arrmul24_and22_15_y0 ^ f_u_arrmul24_fa22_15_f_u_arrmul24_fa23_14_y2;
  assign f_u_arrmul24_fa22_15_y1 = f_u_arrmul24_fa22_15_f_u_arrmul24_and22_15_y0 & f_u_arrmul24_fa22_15_f_u_arrmul24_fa23_14_y2;
  assign f_u_arrmul24_fa22_15_y2 = f_u_arrmul24_fa22_15_y0 ^ f_u_arrmul24_fa22_15_f_u_arrmul24_fa21_15_y4;
  assign f_u_arrmul24_fa22_15_y3 = f_u_arrmul24_fa22_15_y0 & f_u_arrmul24_fa22_15_f_u_arrmul24_fa21_15_y4;
  assign f_u_arrmul24_fa22_15_y4 = f_u_arrmul24_fa22_15_y1 | f_u_arrmul24_fa22_15_y3;
  assign f_u_arrmul24_and23_15_a_23 = a_23;
  assign f_u_arrmul24_and23_15_b_15 = b_15;
  assign f_u_arrmul24_and23_15_y0 = f_u_arrmul24_and23_15_a_23 & f_u_arrmul24_and23_15_b_15;
  assign f_u_arrmul24_fa23_15_f_u_arrmul24_and23_15_y0 = f_u_arrmul24_and23_15_y0;
  assign f_u_arrmul24_fa23_15_f_u_arrmul24_fa23_14_y4 = f_u_arrmul24_fa23_14_y4;
  assign f_u_arrmul24_fa23_15_f_u_arrmul24_fa22_15_y4 = f_u_arrmul24_fa22_15_y4;
  assign f_u_arrmul24_fa23_15_y0 = f_u_arrmul24_fa23_15_f_u_arrmul24_and23_15_y0 ^ f_u_arrmul24_fa23_15_f_u_arrmul24_fa23_14_y4;
  assign f_u_arrmul24_fa23_15_y1 = f_u_arrmul24_fa23_15_f_u_arrmul24_and23_15_y0 & f_u_arrmul24_fa23_15_f_u_arrmul24_fa23_14_y4;
  assign f_u_arrmul24_fa23_15_y2 = f_u_arrmul24_fa23_15_y0 ^ f_u_arrmul24_fa23_15_f_u_arrmul24_fa22_15_y4;
  assign f_u_arrmul24_fa23_15_y3 = f_u_arrmul24_fa23_15_y0 & f_u_arrmul24_fa23_15_f_u_arrmul24_fa22_15_y4;
  assign f_u_arrmul24_fa23_15_y4 = f_u_arrmul24_fa23_15_y1 | f_u_arrmul24_fa23_15_y3;
  assign f_u_arrmul24_and0_16_a_0 = a_0;
  assign f_u_arrmul24_and0_16_b_16 = b_16;
  assign f_u_arrmul24_and0_16_y0 = f_u_arrmul24_and0_16_a_0 & f_u_arrmul24_and0_16_b_16;
  assign f_u_arrmul24_ha0_16_f_u_arrmul24_and0_16_y0 = f_u_arrmul24_and0_16_y0;
  assign f_u_arrmul24_ha0_16_f_u_arrmul24_fa1_15_y2 = f_u_arrmul24_fa1_15_y2;
  assign f_u_arrmul24_ha0_16_y0 = f_u_arrmul24_ha0_16_f_u_arrmul24_and0_16_y0 ^ f_u_arrmul24_ha0_16_f_u_arrmul24_fa1_15_y2;
  assign f_u_arrmul24_ha0_16_y1 = f_u_arrmul24_ha0_16_f_u_arrmul24_and0_16_y0 & f_u_arrmul24_ha0_16_f_u_arrmul24_fa1_15_y2;
  assign f_u_arrmul24_and1_16_a_1 = a_1;
  assign f_u_arrmul24_and1_16_b_16 = b_16;
  assign f_u_arrmul24_and1_16_y0 = f_u_arrmul24_and1_16_a_1 & f_u_arrmul24_and1_16_b_16;
  assign f_u_arrmul24_fa1_16_f_u_arrmul24_and1_16_y0 = f_u_arrmul24_and1_16_y0;
  assign f_u_arrmul24_fa1_16_f_u_arrmul24_fa2_15_y2 = f_u_arrmul24_fa2_15_y2;
  assign f_u_arrmul24_fa1_16_f_u_arrmul24_ha0_16_y1 = f_u_arrmul24_ha0_16_y1;
  assign f_u_arrmul24_fa1_16_y0 = f_u_arrmul24_fa1_16_f_u_arrmul24_and1_16_y0 ^ f_u_arrmul24_fa1_16_f_u_arrmul24_fa2_15_y2;
  assign f_u_arrmul24_fa1_16_y1 = f_u_arrmul24_fa1_16_f_u_arrmul24_and1_16_y0 & f_u_arrmul24_fa1_16_f_u_arrmul24_fa2_15_y2;
  assign f_u_arrmul24_fa1_16_y2 = f_u_arrmul24_fa1_16_y0 ^ f_u_arrmul24_fa1_16_f_u_arrmul24_ha0_16_y1;
  assign f_u_arrmul24_fa1_16_y3 = f_u_arrmul24_fa1_16_y0 & f_u_arrmul24_fa1_16_f_u_arrmul24_ha0_16_y1;
  assign f_u_arrmul24_fa1_16_y4 = f_u_arrmul24_fa1_16_y1 | f_u_arrmul24_fa1_16_y3;
  assign f_u_arrmul24_and2_16_a_2 = a_2;
  assign f_u_arrmul24_and2_16_b_16 = b_16;
  assign f_u_arrmul24_and2_16_y0 = f_u_arrmul24_and2_16_a_2 & f_u_arrmul24_and2_16_b_16;
  assign f_u_arrmul24_fa2_16_f_u_arrmul24_and2_16_y0 = f_u_arrmul24_and2_16_y0;
  assign f_u_arrmul24_fa2_16_f_u_arrmul24_fa3_15_y2 = f_u_arrmul24_fa3_15_y2;
  assign f_u_arrmul24_fa2_16_f_u_arrmul24_fa1_16_y4 = f_u_arrmul24_fa1_16_y4;
  assign f_u_arrmul24_fa2_16_y0 = f_u_arrmul24_fa2_16_f_u_arrmul24_and2_16_y0 ^ f_u_arrmul24_fa2_16_f_u_arrmul24_fa3_15_y2;
  assign f_u_arrmul24_fa2_16_y1 = f_u_arrmul24_fa2_16_f_u_arrmul24_and2_16_y0 & f_u_arrmul24_fa2_16_f_u_arrmul24_fa3_15_y2;
  assign f_u_arrmul24_fa2_16_y2 = f_u_arrmul24_fa2_16_y0 ^ f_u_arrmul24_fa2_16_f_u_arrmul24_fa1_16_y4;
  assign f_u_arrmul24_fa2_16_y3 = f_u_arrmul24_fa2_16_y0 & f_u_arrmul24_fa2_16_f_u_arrmul24_fa1_16_y4;
  assign f_u_arrmul24_fa2_16_y4 = f_u_arrmul24_fa2_16_y1 | f_u_arrmul24_fa2_16_y3;
  assign f_u_arrmul24_and3_16_a_3 = a_3;
  assign f_u_arrmul24_and3_16_b_16 = b_16;
  assign f_u_arrmul24_and3_16_y0 = f_u_arrmul24_and3_16_a_3 & f_u_arrmul24_and3_16_b_16;
  assign f_u_arrmul24_fa3_16_f_u_arrmul24_and3_16_y0 = f_u_arrmul24_and3_16_y0;
  assign f_u_arrmul24_fa3_16_f_u_arrmul24_fa4_15_y2 = f_u_arrmul24_fa4_15_y2;
  assign f_u_arrmul24_fa3_16_f_u_arrmul24_fa2_16_y4 = f_u_arrmul24_fa2_16_y4;
  assign f_u_arrmul24_fa3_16_y0 = f_u_arrmul24_fa3_16_f_u_arrmul24_and3_16_y0 ^ f_u_arrmul24_fa3_16_f_u_arrmul24_fa4_15_y2;
  assign f_u_arrmul24_fa3_16_y1 = f_u_arrmul24_fa3_16_f_u_arrmul24_and3_16_y0 & f_u_arrmul24_fa3_16_f_u_arrmul24_fa4_15_y2;
  assign f_u_arrmul24_fa3_16_y2 = f_u_arrmul24_fa3_16_y0 ^ f_u_arrmul24_fa3_16_f_u_arrmul24_fa2_16_y4;
  assign f_u_arrmul24_fa3_16_y3 = f_u_arrmul24_fa3_16_y0 & f_u_arrmul24_fa3_16_f_u_arrmul24_fa2_16_y4;
  assign f_u_arrmul24_fa3_16_y4 = f_u_arrmul24_fa3_16_y1 | f_u_arrmul24_fa3_16_y3;
  assign f_u_arrmul24_and4_16_a_4 = a_4;
  assign f_u_arrmul24_and4_16_b_16 = b_16;
  assign f_u_arrmul24_and4_16_y0 = f_u_arrmul24_and4_16_a_4 & f_u_arrmul24_and4_16_b_16;
  assign f_u_arrmul24_fa4_16_f_u_arrmul24_and4_16_y0 = f_u_arrmul24_and4_16_y0;
  assign f_u_arrmul24_fa4_16_f_u_arrmul24_fa5_15_y2 = f_u_arrmul24_fa5_15_y2;
  assign f_u_arrmul24_fa4_16_f_u_arrmul24_fa3_16_y4 = f_u_arrmul24_fa3_16_y4;
  assign f_u_arrmul24_fa4_16_y0 = f_u_arrmul24_fa4_16_f_u_arrmul24_and4_16_y0 ^ f_u_arrmul24_fa4_16_f_u_arrmul24_fa5_15_y2;
  assign f_u_arrmul24_fa4_16_y1 = f_u_arrmul24_fa4_16_f_u_arrmul24_and4_16_y0 & f_u_arrmul24_fa4_16_f_u_arrmul24_fa5_15_y2;
  assign f_u_arrmul24_fa4_16_y2 = f_u_arrmul24_fa4_16_y0 ^ f_u_arrmul24_fa4_16_f_u_arrmul24_fa3_16_y4;
  assign f_u_arrmul24_fa4_16_y3 = f_u_arrmul24_fa4_16_y0 & f_u_arrmul24_fa4_16_f_u_arrmul24_fa3_16_y4;
  assign f_u_arrmul24_fa4_16_y4 = f_u_arrmul24_fa4_16_y1 | f_u_arrmul24_fa4_16_y3;
  assign f_u_arrmul24_and5_16_a_5 = a_5;
  assign f_u_arrmul24_and5_16_b_16 = b_16;
  assign f_u_arrmul24_and5_16_y0 = f_u_arrmul24_and5_16_a_5 & f_u_arrmul24_and5_16_b_16;
  assign f_u_arrmul24_fa5_16_f_u_arrmul24_and5_16_y0 = f_u_arrmul24_and5_16_y0;
  assign f_u_arrmul24_fa5_16_f_u_arrmul24_fa6_15_y2 = f_u_arrmul24_fa6_15_y2;
  assign f_u_arrmul24_fa5_16_f_u_arrmul24_fa4_16_y4 = f_u_arrmul24_fa4_16_y4;
  assign f_u_arrmul24_fa5_16_y0 = f_u_arrmul24_fa5_16_f_u_arrmul24_and5_16_y0 ^ f_u_arrmul24_fa5_16_f_u_arrmul24_fa6_15_y2;
  assign f_u_arrmul24_fa5_16_y1 = f_u_arrmul24_fa5_16_f_u_arrmul24_and5_16_y0 & f_u_arrmul24_fa5_16_f_u_arrmul24_fa6_15_y2;
  assign f_u_arrmul24_fa5_16_y2 = f_u_arrmul24_fa5_16_y0 ^ f_u_arrmul24_fa5_16_f_u_arrmul24_fa4_16_y4;
  assign f_u_arrmul24_fa5_16_y3 = f_u_arrmul24_fa5_16_y0 & f_u_arrmul24_fa5_16_f_u_arrmul24_fa4_16_y4;
  assign f_u_arrmul24_fa5_16_y4 = f_u_arrmul24_fa5_16_y1 | f_u_arrmul24_fa5_16_y3;
  assign f_u_arrmul24_and6_16_a_6 = a_6;
  assign f_u_arrmul24_and6_16_b_16 = b_16;
  assign f_u_arrmul24_and6_16_y0 = f_u_arrmul24_and6_16_a_6 & f_u_arrmul24_and6_16_b_16;
  assign f_u_arrmul24_fa6_16_f_u_arrmul24_and6_16_y0 = f_u_arrmul24_and6_16_y0;
  assign f_u_arrmul24_fa6_16_f_u_arrmul24_fa7_15_y2 = f_u_arrmul24_fa7_15_y2;
  assign f_u_arrmul24_fa6_16_f_u_arrmul24_fa5_16_y4 = f_u_arrmul24_fa5_16_y4;
  assign f_u_arrmul24_fa6_16_y0 = f_u_arrmul24_fa6_16_f_u_arrmul24_and6_16_y0 ^ f_u_arrmul24_fa6_16_f_u_arrmul24_fa7_15_y2;
  assign f_u_arrmul24_fa6_16_y1 = f_u_arrmul24_fa6_16_f_u_arrmul24_and6_16_y0 & f_u_arrmul24_fa6_16_f_u_arrmul24_fa7_15_y2;
  assign f_u_arrmul24_fa6_16_y2 = f_u_arrmul24_fa6_16_y0 ^ f_u_arrmul24_fa6_16_f_u_arrmul24_fa5_16_y4;
  assign f_u_arrmul24_fa6_16_y3 = f_u_arrmul24_fa6_16_y0 & f_u_arrmul24_fa6_16_f_u_arrmul24_fa5_16_y4;
  assign f_u_arrmul24_fa6_16_y4 = f_u_arrmul24_fa6_16_y1 | f_u_arrmul24_fa6_16_y3;
  assign f_u_arrmul24_and7_16_a_7 = a_7;
  assign f_u_arrmul24_and7_16_b_16 = b_16;
  assign f_u_arrmul24_and7_16_y0 = f_u_arrmul24_and7_16_a_7 & f_u_arrmul24_and7_16_b_16;
  assign f_u_arrmul24_fa7_16_f_u_arrmul24_and7_16_y0 = f_u_arrmul24_and7_16_y0;
  assign f_u_arrmul24_fa7_16_f_u_arrmul24_fa8_15_y2 = f_u_arrmul24_fa8_15_y2;
  assign f_u_arrmul24_fa7_16_f_u_arrmul24_fa6_16_y4 = f_u_arrmul24_fa6_16_y4;
  assign f_u_arrmul24_fa7_16_y0 = f_u_arrmul24_fa7_16_f_u_arrmul24_and7_16_y0 ^ f_u_arrmul24_fa7_16_f_u_arrmul24_fa8_15_y2;
  assign f_u_arrmul24_fa7_16_y1 = f_u_arrmul24_fa7_16_f_u_arrmul24_and7_16_y0 & f_u_arrmul24_fa7_16_f_u_arrmul24_fa8_15_y2;
  assign f_u_arrmul24_fa7_16_y2 = f_u_arrmul24_fa7_16_y0 ^ f_u_arrmul24_fa7_16_f_u_arrmul24_fa6_16_y4;
  assign f_u_arrmul24_fa7_16_y3 = f_u_arrmul24_fa7_16_y0 & f_u_arrmul24_fa7_16_f_u_arrmul24_fa6_16_y4;
  assign f_u_arrmul24_fa7_16_y4 = f_u_arrmul24_fa7_16_y1 | f_u_arrmul24_fa7_16_y3;
  assign f_u_arrmul24_and8_16_a_8 = a_8;
  assign f_u_arrmul24_and8_16_b_16 = b_16;
  assign f_u_arrmul24_and8_16_y0 = f_u_arrmul24_and8_16_a_8 & f_u_arrmul24_and8_16_b_16;
  assign f_u_arrmul24_fa8_16_f_u_arrmul24_and8_16_y0 = f_u_arrmul24_and8_16_y0;
  assign f_u_arrmul24_fa8_16_f_u_arrmul24_fa9_15_y2 = f_u_arrmul24_fa9_15_y2;
  assign f_u_arrmul24_fa8_16_f_u_arrmul24_fa7_16_y4 = f_u_arrmul24_fa7_16_y4;
  assign f_u_arrmul24_fa8_16_y0 = f_u_arrmul24_fa8_16_f_u_arrmul24_and8_16_y0 ^ f_u_arrmul24_fa8_16_f_u_arrmul24_fa9_15_y2;
  assign f_u_arrmul24_fa8_16_y1 = f_u_arrmul24_fa8_16_f_u_arrmul24_and8_16_y0 & f_u_arrmul24_fa8_16_f_u_arrmul24_fa9_15_y2;
  assign f_u_arrmul24_fa8_16_y2 = f_u_arrmul24_fa8_16_y0 ^ f_u_arrmul24_fa8_16_f_u_arrmul24_fa7_16_y4;
  assign f_u_arrmul24_fa8_16_y3 = f_u_arrmul24_fa8_16_y0 & f_u_arrmul24_fa8_16_f_u_arrmul24_fa7_16_y4;
  assign f_u_arrmul24_fa8_16_y4 = f_u_arrmul24_fa8_16_y1 | f_u_arrmul24_fa8_16_y3;
  assign f_u_arrmul24_and9_16_a_9 = a_9;
  assign f_u_arrmul24_and9_16_b_16 = b_16;
  assign f_u_arrmul24_and9_16_y0 = f_u_arrmul24_and9_16_a_9 & f_u_arrmul24_and9_16_b_16;
  assign f_u_arrmul24_fa9_16_f_u_arrmul24_and9_16_y0 = f_u_arrmul24_and9_16_y0;
  assign f_u_arrmul24_fa9_16_f_u_arrmul24_fa10_15_y2 = f_u_arrmul24_fa10_15_y2;
  assign f_u_arrmul24_fa9_16_f_u_arrmul24_fa8_16_y4 = f_u_arrmul24_fa8_16_y4;
  assign f_u_arrmul24_fa9_16_y0 = f_u_arrmul24_fa9_16_f_u_arrmul24_and9_16_y0 ^ f_u_arrmul24_fa9_16_f_u_arrmul24_fa10_15_y2;
  assign f_u_arrmul24_fa9_16_y1 = f_u_arrmul24_fa9_16_f_u_arrmul24_and9_16_y0 & f_u_arrmul24_fa9_16_f_u_arrmul24_fa10_15_y2;
  assign f_u_arrmul24_fa9_16_y2 = f_u_arrmul24_fa9_16_y0 ^ f_u_arrmul24_fa9_16_f_u_arrmul24_fa8_16_y4;
  assign f_u_arrmul24_fa9_16_y3 = f_u_arrmul24_fa9_16_y0 & f_u_arrmul24_fa9_16_f_u_arrmul24_fa8_16_y4;
  assign f_u_arrmul24_fa9_16_y4 = f_u_arrmul24_fa9_16_y1 | f_u_arrmul24_fa9_16_y3;
  assign f_u_arrmul24_and10_16_a_10 = a_10;
  assign f_u_arrmul24_and10_16_b_16 = b_16;
  assign f_u_arrmul24_and10_16_y0 = f_u_arrmul24_and10_16_a_10 & f_u_arrmul24_and10_16_b_16;
  assign f_u_arrmul24_fa10_16_f_u_arrmul24_and10_16_y0 = f_u_arrmul24_and10_16_y0;
  assign f_u_arrmul24_fa10_16_f_u_arrmul24_fa11_15_y2 = f_u_arrmul24_fa11_15_y2;
  assign f_u_arrmul24_fa10_16_f_u_arrmul24_fa9_16_y4 = f_u_arrmul24_fa9_16_y4;
  assign f_u_arrmul24_fa10_16_y0 = f_u_arrmul24_fa10_16_f_u_arrmul24_and10_16_y0 ^ f_u_arrmul24_fa10_16_f_u_arrmul24_fa11_15_y2;
  assign f_u_arrmul24_fa10_16_y1 = f_u_arrmul24_fa10_16_f_u_arrmul24_and10_16_y0 & f_u_arrmul24_fa10_16_f_u_arrmul24_fa11_15_y2;
  assign f_u_arrmul24_fa10_16_y2 = f_u_arrmul24_fa10_16_y0 ^ f_u_arrmul24_fa10_16_f_u_arrmul24_fa9_16_y4;
  assign f_u_arrmul24_fa10_16_y3 = f_u_arrmul24_fa10_16_y0 & f_u_arrmul24_fa10_16_f_u_arrmul24_fa9_16_y4;
  assign f_u_arrmul24_fa10_16_y4 = f_u_arrmul24_fa10_16_y1 | f_u_arrmul24_fa10_16_y3;
  assign f_u_arrmul24_and11_16_a_11 = a_11;
  assign f_u_arrmul24_and11_16_b_16 = b_16;
  assign f_u_arrmul24_and11_16_y0 = f_u_arrmul24_and11_16_a_11 & f_u_arrmul24_and11_16_b_16;
  assign f_u_arrmul24_fa11_16_f_u_arrmul24_and11_16_y0 = f_u_arrmul24_and11_16_y0;
  assign f_u_arrmul24_fa11_16_f_u_arrmul24_fa12_15_y2 = f_u_arrmul24_fa12_15_y2;
  assign f_u_arrmul24_fa11_16_f_u_arrmul24_fa10_16_y4 = f_u_arrmul24_fa10_16_y4;
  assign f_u_arrmul24_fa11_16_y0 = f_u_arrmul24_fa11_16_f_u_arrmul24_and11_16_y0 ^ f_u_arrmul24_fa11_16_f_u_arrmul24_fa12_15_y2;
  assign f_u_arrmul24_fa11_16_y1 = f_u_arrmul24_fa11_16_f_u_arrmul24_and11_16_y0 & f_u_arrmul24_fa11_16_f_u_arrmul24_fa12_15_y2;
  assign f_u_arrmul24_fa11_16_y2 = f_u_arrmul24_fa11_16_y0 ^ f_u_arrmul24_fa11_16_f_u_arrmul24_fa10_16_y4;
  assign f_u_arrmul24_fa11_16_y3 = f_u_arrmul24_fa11_16_y0 & f_u_arrmul24_fa11_16_f_u_arrmul24_fa10_16_y4;
  assign f_u_arrmul24_fa11_16_y4 = f_u_arrmul24_fa11_16_y1 | f_u_arrmul24_fa11_16_y3;
  assign f_u_arrmul24_and12_16_a_12 = a_12;
  assign f_u_arrmul24_and12_16_b_16 = b_16;
  assign f_u_arrmul24_and12_16_y0 = f_u_arrmul24_and12_16_a_12 & f_u_arrmul24_and12_16_b_16;
  assign f_u_arrmul24_fa12_16_f_u_arrmul24_and12_16_y0 = f_u_arrmul24_and12_16_y0;
  assign f_u_arrmul24_fa12_16_f_u_arrmul24_fa13_15_y2 = f_u_arrmul24_fa13_15_y2;
  assign f_u_arrmul24_fa12_16_f_u_arrmul24_fa11_16_y4 = f_u_arrmul24_fa11_16_y4;
  assign f_u_arrmul24_fa12_16_y0 = f_u_arrmul24_fa12_16_f_u_arrmul24_and12_16_y0 ^ f_u_arrmul24_fa12_16_f_u_arrmul24_fa13_15_y2;
  assign f_u_arrmul24_fa12_16_y1 = f_u_arrmul24_fa12_16_f_u_arrmul24_and12_16_y0 & f_u_arrmul24_fa12_16_f_u_arrmul24_fa13_15_y2;
  assign f_u_arrmul24_fa12_16_y2 = f_u_arrmul24_fa12_16_y0 ^ f_u_arrmul24_fa12_16_f_u_arrmul24_fa11_16_y4;
  assign f_u_arrmul24_fa12_16_y3 = f_u_arrmul24_fa12_16_y0 & f_u_arrmul24_fa12_16_f_u_arrmul24_fa11_16_y4;
  assign f_u_arrmul24_fa12_16_y4 = f_u_arrmul24_fa12_16_y1 | f_u_arrmul24_fa12_16_y3;
  assign f_u_arrmul24_and13_16_a_13 = a_13;
  assign f_u_arrmul24_and13_16_b_16 = b_16;
  assign f_u_arrmul24_and13_16_y0 = f_u_arrmul24_and13_16_a_13 & f_u_arrmul24_and13_16_b_16;
  assign f_u_arrmul24_fa13_16_f_u_arrmul24_and13_16_y0 = f_u_arrmul24_and13_16_y0;
  assign f_u_arrmul24_fa13_16_f_u_arrmul24_fa14_15_y2 = f_u_arrmul24_fa14_15_y2;
  assign f_u_arrmul24_fa13_16_f_u_arrmul24_fa12_16_y4 = f_u_arrmul24_fa12_16_y4;
  assign f_u_arrmul24_fa13_16_y0 = f_u_arrmul24_fa13_16_f_u_arrmul24_and13_16_y0 ^ f_u_arrmul24_fa13_16_f_u_arrmul24_fa14_15_y2;
  assign f_u_arrmul24_fa13_16_y1 = f_u_arrmul24_fa13_16_f_u_arrmul24_and13_16_y0 & f_u_arrmul24_fa13_16_f_u_arrmul24_fa14_15_y2;
  assign f_u_arrmul24_fa13_16_y2 = f_u_arrmul24_fa13_16_y0 ^ f_u_arrmul24_fa13_16_f_u_arrmul24_fa12_16_y4;
  assign f_u_arrmul24_fa13_16_y3 = f_u_arrmul24_fa13_16_y0 & f_u_arrmul24_fa13_16_f_u_arrmul24_fa12_16_y4;
  assign f_u_arrmul24_fa13_16_y4 = f_u_arrmul24_fa13_16_y1 | f_u_arrmul24_fa13_16_y3;
  assign f_u_arrmul24_and14_16_a_14 = a_14;
  assign f_u_arrmul24_and14_16_b_16 = b_16;
  assign f_u_arrmul24_and14_16_y0 = f_u_arrmul24_and14_16_a_14 & f_u_arrmul24_and14_16_b_16;
  assign f_u_arrmul24_fa14_16_f_u_arrmul24_and14_16_y0 = f_u_arrmul24_and14_16_y0;
  assign f_u_arrmul24_fa14_16_f_u_arrmul24_fa15_15_y2 = f_u_arrmul24_fa15_15_y2;
  assign f_u_arrmul24_fa14_16_f_u_arrmul24_fa13_16_y4 = f_u_arrmul24_fa13_16_y4;
  assign f_u_arrmul24_fa14_16_y0 = f_u_arrmul24_fa14_16_f_u_arrmul24_and14_16_y0 ^ f_u_arrmul24_fa14_16_f_u_arrmul24_fa15_15_y2;
  assign f_u_arrmul24_fa14_16_y1 = f_u_arrmul24_fa14_16_f_u_arrmul24_and14_16_y0 & f_u_arrmul24_fa14_16_f_u_arrmul24_fa15_15_y2;
  assign f_u_arrmul24_fa14_16_y2 = f_u_arrmul24_fa14_16_y0 ^ f_u_arrmul24_fa14_16_f_u_arrmul24_fa13_16_y4;
  assign f_u_arrmul24_fa14_16_y3 = f_u_arrmul24_fa14_16_y0 & f_u_arrmul24_fa14_16_f_u_arrmul24_fa13_16_y4;
  assign f_u_arrmul24_fa14_16_y4 = f_u_arrmul24_fa14_16_y1 | f_u_arrmul24_fa14_16_y3;
  assign f_u_arrmul24_and15_16_a_15 = a_15;
  assign f_u_arrmul24_and15_16_b_16 = b_16;
  assign f_u_arrmul24_and15_16_y0 = f_u_arrmul24_and15_16_a_15 & f_u_arrmul24_and15_16_b_16;
  assign f_u_arrmul24_fa15_16_f_u_arrmul24_and15_16_y0 = f_u_arrmul24_and15_16_y0;
  assign f_u_arrmul24_fa15_16_f_u_arrmul24_fa16_15_y2 = f_u_arrmul24_fa16_15_y2;
  assign f_u_arrmul24_fa15_16_f_u_arrmul24_fa14_16_y4 = f_u_arrmul24_fa14_16_y4;
  assign f_u_arrmul24_fa15_16_y0 = f_u_arrmul24_fa15_16_f_u_arrmul24_and15_16_y0 ^ f_u_arrmul24_fa15_16_f_u_arrmul24_fa16_15_y2;
  assign f_u_arrmul24_fa15_16_y1 = f_u_arrmul24_fa15_16_f_u_arrmul24_and15_16_y0 & f_u_arrmul24_fa15_16_f_u_arrmul24_fa16_15_y2;
  assign f_u_arrmul24_fa15_16_y2 = f_u_arrmul24_fa15_16_y0 ^ f_u_arrmul24_fa15_16_f_u_arrmul24_fa14_16_y4;
  assign f_u_arrmul24_fa15_16_y3 = f_u_arrmul24_fa15_16_y0 & f_u_arrmul24_fa15_16_f_u_arrmul24_fa14_16_y4;
  assign f_u_arrmul24_fa15_16_y4 = f_u_arrmul24_fa15_16_y1 | f_u_arrmul24_fa15_16_y3;
  assign f_u_arrmul24_and16_16_a_16 = a_16;
  assign f_u_arrmul24_and16_16_b_16 = b_16;
  assign f_u_arrmul24_and16_16_y0 = f_u_arrmul24_and16_16_a_16 & f_u_arrmul24_and16_16_b_16;
  assign f_u_arrmul24_fa16_16_f_u_arrmul24_and16_16_y0 = f_u_arrmul24_and16_16_y0;
  assign f_u_arrmul24_fa16_16_f_u_arrmul24_fa17_15_y2 = f_u_arrmul24_fa17_15_y2;
  assign f_u_arrmul24_fa16_16_f_u_arrmul24_fa15_16_y4 = f_u_arrmul24_fa15_16_y4;
  assign f_u_arrmul24_fa16_16_y0 = f_u_arrmul24_fa16_16_f_u_arrmul24_and16_16_y0 ^ f_u_arrmul24_fa16_16_f_u_arrmul24_fa17_15_y2;
  assign f_u_arrmul24_fa16_16_y1 = f_u_arrmul24_fa16_16_f_u_arrmul24_and16_16_y0 & f_u_arrmul24_fa16_16_f_u_arrmul24_fa17_15_y2;
  assign f_u_arrmul24_fa16_16_y2 = f_u_arrmul24_fa16_16_y0 ^ f_u_arrmul24_fa16_16_f_u_arrmul24_fa15_16_y4;
  assign f_u_arrmul24_fa16_16_y3 = f_u_arrmul24_fa16_16_y0 & f_u_arrmul24_fa16_16_f_u_arrmul24_fa15_16_y4;
  assign f_u_arrmul24_fa16_16_y4 = f_u_arrmul24_fa16_16_y1 | f_u_arrmul24_fa16_16_y3;
  assign f_u_arrmul24_and17_16_a_17 = a_17;
  assign f_u_arrmul24_and17_16_b_16 = b_16;
  assign f_u_arrmul24_and17_16_y0 = f_u_arrmul24_and17_16_a_17 & f_u_arrmul24_and17_16_b_16;
  assign f_u_arrmul24_fa17_16_f_u_arrmul24_and17_16_y0 = f_u_arrmul24_and17_16_y0;
  assign f_u_arrmul24_fa17_16_f_u_arrmul24_fa18_15_y2 = f_u_arrmul24_fa18_15_y2;
  assign f_u_arrmul24_fa17_16_f_u_arrmul24_fa16_16_y4 = f_u_arrmul24_fa16_16_y4;
  assign f_u_arrmul24_fa17_16_y0 = f_u_arrmul24_fa17_16_f_u_arrmul24_and17_16_y0 ^ f_u_arrmul24_fa17_16_f_u_arrmul24_fa18_15_y2;
  assign f_u_arrmul24_fa17_16_y1 = f_u_arrmul24_fa17_16_f_u_arrmul24_and17_16_y0 & f_u_arrmul24_fa17_16_f_u_arrmul24_fa18_15_y2;
  assign f_u_arrmul24_fa17_16_y2 = f_u_arrmul24_fa17_16_y0 ^ f_u_arrmul24_fa17_16_f_u_arrmul24_fa16_16_y4;
  assign f_u_arrmul24_fa17_16_y3 = f_u_arrmul24_fa17_16_y0 & f_u_arrmul24_fa17_16_f_u_arrmul24_fa16_16_y4;
  assign f_u_arrmul24_fa17_16_y4 = f_u_arrmul24_fa17_16_y1 | f_u_arrmul24_fa17_16_y3;
  assign f_u_arrmul24_and18_16_a_18 = a_18;
  assign f_u_arrmul24_and18_16_b_16 = b_16;
  assign f_u_arrmul24_and18_16_y0 = f_u_arrmul24_and18_16_a_18 & f_u_arrmul24_and18_16_b_16;
  assign f_u_arrmul24_fa18_16_f_u_arrmul24_and18_16_y0 = f_u_arrmul24_and18_16_y0;
  assign f_u_arrmul24_fa18_16_f_u_arrmul24_fa19_15_y2 = f_u_arrmul24_fa19_15_y2;
  assign f_u_arrmul24_fa18_16_f_u_arrmul24_fa17_16_y4 = f_u_arrmul24_fa17_16_y4;
  assign f_u_arrmul24_fa18_16_y0 = f_u_arrmul24_fa18_16_f_u_arrmul24_and18_16_y0 ^ f_u_arrmul24_fa18_16_f_u_arrmul24_fa19_15_y2;
  assign f_u_arrmul24_fa18_16_y1 = f_u_arrmul24_fa18_16_f_u_arrmul24_and18_16_y0 & f_u_arrmul24_fa18_16_f_u_arrmul24_fa19_15_y2;
  assign f_u_arrmul24_fa18_16_y2 = f_u_arrmul24_fa18_16_y0 ^ f_u_arrmul24_fa18_16_f_u_arrmul24_fa17_16_y4;
  assign f_u_arrmul24_fa18_16_y3 = f_u_arrmul24_fa18_16_y0 & f_u_arrmul24_fa18_16_f_u_arrmul24_fa17_16_y4;
  assign f_u_arrmul24_fa18_16_y4 = f_u_arrmul24_fa18_16_y1 | f_u_arrmul24_fa18_16_y3;
  assign f_u_arrmul24_and19_16_a_19 = a_19;
  assign f_u_arrmul24_and19_16_b_16 = b_16;
  assign f_u_arrmul24_and19_16_y0 = f_u_arrmul24_and19_16_a_19 & f_u_arrmul24_and19_16_b_16;
  assign f_u_arrmul24_fa19_16_f_u_arrmul24_and19_16_y0 = f_u_arrmul24_and19_16_y0;
  assign f_u_arrmul24_fa19_16_f_u_arrmul24_fa20_15_y2 = f_u_arrmul24_fa20_15_y2;
  assign f_u_arrmul24_fa19_16_f_u_arrmul24_fa18_16_y4 = f_u_arrmul24_fa18_16_y4;
  assign f_u_arrmul24_fa19_16_y0 = f_u_arrmul24_fa19_16_f_u_arrmul24_and19_16_y0 ^ f_u_arrmul24_fa19_16_f_u_arrmul24_fa20_15_y2;
  assign f_u_arrmul24_fa19_16_y1 = f_u_arrmul24_fa19_16_f_u_arrmul24_and19_16_y0 & f_u_arrmul24_fa19_16_f_u_arrmul24_fa20_15_y2;
  assign f_u_arrmul24_fa19_16_y2 = f_u_arrmul24_fa19_16_y0 ^ f_u_arrmul24_fa19_16_f_u_arrmul24_fa18_16_y4;
  assign f_u_arrmul24_fa19_16_y3 = f_u_arrmul24_fa19_16_y0 & f_u_arrmul24_fa19_16_f_u_arrmul24_fa18_16_y4;
  assign f_u_arrmul24_fa19_16_y4 = f_u_arrmul24_fa19_16_y1 | f_u_arrmul24_fa19_16_y3;
  assign f_u_arrmul24_and20_16_a_20 = a_20;
  assign f_u_arrmul24_and20_16_b_16 = b_16;
  assign f_u_arrmul24_and20_16_y0 = f_u_arrmul24_and20_16_a_20 & f_u_arrmul24_and20_16_b_16;
  assign f_u_arrmul24_fa20_16_f_u_arrmul24_and20_16_y0 = f_u_arrmul24_and20_16_y0;
  assign f_u_arrmul24_fa20_16_f_u_arrmul24_fa21_15_y2 = f_u_arrmul24_fa21_15_y2;
  assign f_u_arrmul24_fa20_16_f_u_arrmul24_fa19_16_y4 = f_u_arrmul24_fa19_16_y4;
  assign f_u_arrmul24_fa20_16_y0 = f_u_arrmul24_fa20_16_f_u_arrmul24_and20_16_y0 ^ f_u_arrmul24_fa20_16_f_u_arrmul24_fa21_15_y2;
  assign f_u_arrmul24_fa20_16_y1 = f_u_arrmul24_fa20_16_f_u_arrmul24_and20_16_y0 & f_u_arrmul24_fa20_16_f_u_arrmul24_fa21_15_y2;
  assign f_u_arrmul24_fa20_16_y2 = f_u_arrmul24_fa20_16_y0 ^ f_u_arrmul24_fa20_16_f_u_arrmul24_fa19_16_y4;
  assign f_u_arrmul24_fa20_16_y3 = f_u_arrmul24_fa20_16_y0 & f_u_arrmul24_fa20_16_f_u_arrmul24_fa19_16_y4;
  assign f_u_arrmul24_fa20_16_y4 = f_u_arrmul24_fa20_16_y1 | f_u_arrmul24_fa20_16_y3;
  assign f_u_arrmul24_and21_16_a_21 = a_21;
  assign f_u_arrmul24_and21_16_b_16 = b_16;
  assign f_u_arrmul24_and21_16_y0 = f_u_arrmul24_and21_16_a_21 & f_u_arrmul24_and21_16_b_16;
  assign f_u_arrmul24_fa21_16_f_u_arrmul24_and21_16_y0 = f_u_arrmul24_and21_16_y0;
  assign f_u_arrmul24_fa21_16_f_u_arrmul24_fa22_15_y2 = f_u_arrmul24_fa22_15_y2;
  assign f_u_arrmul24_fa21_16_f_u_arrmul24_fa20_16_y4 = f_u_arrmul24_fa20_16_y4;
  assign f_u_arrmul24_fa21_16_y0 = f_u_arrmul24_fa21_16_f_u_arrmul24_and21_16_y0 ^ f_u_arrmul24_fa21_16_f_u_arrmul24_fa22_15_y2;
  assign f_u_arrmul24_fa21_16_y1 = f_u_arrmul24_fa21_16_f_u_arrmul24_and21_16_y0 & f_u_arrmul24_fa21_16_f_u_arrmul24_fa22_15_y2;
  assign f_u_arrmul24_fa21_16_y2 = f_u_arrmul24_fa21_16_y0 ^ f_u_arrmul24_fa21_16_f_u_arrmul24_fa20_16_y4;
  assign f_u_arrmul24_fa21_16_y3 = f_u_arrmul24_fa21_16_y0 & f_u_arrmul24_fa21_16_f_u_arrmul24_fa20_16_y4;
  assign f_u_arrmul24_fa21_16_y4 = f_u_arrmul24_fa21_16_y1 | f_u_arrmul24_fa21_16_y3;
  assign f_u_arrmul24_and22_16_a_22 = a_22;
  assign f_u_arrmul24_and22_16_b_16 = b_16;
  assign f_u_arrmul24_and22_16_y0 = f_u_arrmul24_and22_16_a_22 & f_u_arrmul24_and22_16_b_16;
  assign f_u_arrmul24_fa22_16_f_u_arrmul24_and22_16_y0 = f_u_arrmul24_and22_16_y0;
  assign f_u_arrmul24_fa22_16_f_u_arrmul24_fa23_15_y2 = f_u_arrmul24_fa23_15_y2;
  assign f_u_arrmul24_fa22_16_f_u_arrmul24_fa21_16_y4 = f_u_arrmul24_fa21_16_y4;
  assign f_u_arrmul24_fa22_16_y0 = f_u_arrmul24_fa22_16_f_u_arrmul24_and22_16_y0 ^ f_u_arrmul24_fa22_16_f_u_arrmul24_fa23_15_y2;
  assign f_u_arrmul24_fa22_16_y1 = f_u_arrmul24_fa22_16_f_u_arrmul24_and22_16_y0 & f_u_arrmul24_fa22_16_f_u_arrmul24_fa23_15_y2;
  assign f_u_arrmul24_fa22_16_y2 = f_u_arrmul24_fa22_16_y0 ^ f_u_arrmul24_fa22_16_f_u_arrmul24_fa21_16_y4;
  assign f_u_arrmul24_fa22_16_y3 = f_u_arrmul24_fa22_16_y0 & f_u_arrmul24_fa22_16_f_u_arrmul24_fa21_16_y4;
  assign f_u_arrmul24_fa22_16_y4 = f_u_arrmul24_fa22_16_y1 | f_u_arrmul24_fa22_16_y3;
  assign f_u_arrmul24_and23_16_a_23 = a_23;
  assign f_u_arrmul24_and23_16_b_16 = b_16;
  assign f_u_arrmul24_and23_16_y0 = f_u_arrmul24_and23_16_a_23 & f_u_arrmul24_and23_16_b_16;
  assign f_u_arrmul24_fa23_16_f_u_arrmul24_and23_16_y0 = f_u_arrmul24_and23_16_y0;
  assign f_u_arrmul24_fa23_16_f_u_arrmul24_fa23_15_y4 = f_u_arrmul24_fa23_15_y4;
  assign f_u_arrmul24_fa23_16_f_u_arrmul24_fa22_16_y4 = f_u_arrmul24_fa22_16_y4;
  assign f_u_arrmul24_fa23_16_y0 = f_u_arrmul24_fa23_16_f_u_arrmul24_and23_16_y0 ^ f_u_arrmul24_fa23_16_f_u_arrmul24_fa23_15_y4;
  assign f_u_arrmul24_fa23_16_y1 = f_u_arrmul24_fa23_16_f_u_arrmul24_and23_16_y0 & f_u_arrmul24_fa23_16_f_u_arrmul24_fa23_15_y4;
  assign f_u_arrmul24_fa23_16_y2 = f_u_arrmul24_fa23_16_y0 ^ f_u_arrmul24_fa23_16_f_u_arrmul24_fa22_16_y4;
  assign f_u_arrmul24_fa23_16_y3 = f_u_arrmul24_fa23_16_y0 & f_u_arrmul24_fa23_16_f_u_arrmul24_fa22_16_y4;
  assign f_u_arrmul24_fa23_16_y4 = f_u_arrmul24_fa23_16_y1 | f_u_arrmul24_fa23_16_y3;
  assign f_u_arrmul24_and0_17_a_0 = a_0;
  assign f_u_arrmul24_and0_17_b_17 = b_17;
  assign f_u_arrmul24_and0_17_y0 = f_u_arrmul24_and0_17_a_0 & f_u_arrmul24_and0_17_b_17;
  assign f_u_arrmul24_ha0_17_f_u_arrmul24_and0_17_y0 = f_u_arrmul24_and0_17_y0;
  assign f_u_arrmul24_ha0_17_f_u_arrmul24_fa1_16_y2 = f_u_arrmul24_fa1_16_y2;
  assign f_u_arrmul24_ha0_17_y0 = f_u_arrmul24_ha0_17_f_u_arrmul24_and0_17_y0 ^ f_u_arrmul24_ha0_17_f_u_arrmul24_fa1_16_y2;
  assign f_u_arrmul24_ha0_17_y1 = f_u_arrmul24_ha0_17_f_u_arrmul24_and0_17_y0 & f_u_arrmul24_ha0_17_f_u_arrmul24_fa1_16_y2;
  assign f_u_arrmul24_and1_17_a_1 = a_1;
  assign f_u_arrmul24_and1_17_b_17 = b_17;
  assign f_u_arrmul24_and1_17_y0 = f_u_arrmul24_and1_17_a_1 & f_u_arrmul24_and1_17_b_17;
  assign f_u_arrmul24_fa1_17_f_u_arrmul24_and1_17_y0 = f_u_arrmul24_and1_17_y0;
  assign f_u_arrmul24_fa1_17_f_u_arrmul24_fa2_16_y2 = f_u_arrmul24_fa2_16_y2;
  assign f_u_arrmul24_fa1_17_f_u_arrmul24_ha0_17_y1 = f_u_arrmul24_ha0_17_y1;
  assign f_u_arrmul24_fa1_17_y0 = f_u_arrmul24_fa1_17_f_u_arrmul24_and1_17_y0 ^ f_u_arrmul24_fa1_17_f_u_arrmul24_fa2_16_y2;
  assign f_u_arrmul24_fa1_17_y1 = f_u_arrmul24_fa1_17_f_u_arrmul24_and1_17_y0 & f_u_arrmul24_fa1_17_f_u_arrmul24_fa2_16_y2;
  assign f_u_arrmul24_fa1_17_y2 = f_u_arrmul24_fa1_17_y0 ^ f_u_arrmul24_fa1_17_f_u_arrmul24_ha0_17_y1;
  assign f_u_arrmul24_fa1_17_y3 = f_u_arrmul24_fa1_17_y0 & f_u_arrmul24_fa1_17_f_u_arrmul24_ha0_17_y1;
  assign f_u_arrmul24_fa1_17_y4 = f_u_arrmul24_fa1_17_y1 | f_u_arrmul24_fa1_17_y3;
  assign f_u_arrmul24_and2_17_a_2 = a_2;
  assign f_u_arrmul24_and2_17_b_17 = b_17;
  assign f_u_arrmul24_and2_17_y0 = f_u_arrmul24_and2_17_a_2 & f_u_arrmul24_and2_17_b_17;
  assign f_u_arrmul24_fa2_17_f_u_arrmul24_and2_17_y0 = f_u_arrmul24_and2_17_y0;
  assign f_u_arrmul24_fa2_17_f_u_arrmul24_fa3_16_y2 = f_u_arrmul24_fa3_16_y2;
  assign f_u_arrmul24_fa2_17_f_u_arrmul24_fa1_17_y4 = f_u_arrmul24_fa1_17_y4;
  assign f_u_arrmul24_fa2_17_y0 = f_u_arrmul24_fa2_17_f_u_arrmul24_and2_17_y0 ^ f_u_arrmul24_fa2_17_f_u_arrmul24_fa3_16_y2;
  assign f_u_arrmul24_fa2_17_y1 = f_u_arrmul24_fa2_17_f_u_arrmul24_and2_17_y0 & f_u_arrmul24_fa2_17_f_u_arrmul24_fa3_16_y2;
  assign f_u_arrmul24_fa2_17_y2 = f_u_arrmul24_fa2_17_y0 ^ f_u_arrmul24_fa2_17_f_u_arrmul24_fa1_17_y4;
  assign f_u_arrmul24_fa2_17_y3 = f_u_arrmul24_fa2_17_y0 & f_u_arrmul24_fa2_17_f_u_arrmul24_fa1_17_y4;
  assign f_u_arrmul24_fa2_17_y4 = f_u_arrmul24_fa2_17_y1 | f_u_arrmul24_fa2_17_y3;
  assign f_u_arrmul24_and3_17_a_3 = a_3;
  assign f_u_arrmul24_and3_17_b_17 = b_17;
  assign f_u_arrmul24_and3_17_y0 = f_u_arrmul24_and3_17_a_3 & f_u_arrmul24_and3_17_b_17;
  assign f_u_arrmul24_fa3_17_f_u_arrmul24_and3_17_y0 = f_u_arrmul24_and3_17_y0;
  assign f_u_arrmul24_fa3_17_f_u_arrmul24_fa4_16_y2 = f_u_arrmul24_fa4_16_y2;
  assign f_u_arrmul24_fa3_17_f_u_arrmul24_fa2_17_y4 = f_u_arrmul24_fa2_17_y4;
  assign f_u_arrmul24_fa3_17_y0 = f_u_arrmul24_fa3_17_f_u_arrmul24_and3_17_y0 ^ f_u_arrmul24_fa3_17_f_u_arrmul24_fa4_16_y2;
  assign f_u_arrmul24_fa3_17_y1 = f_u_arrmul24_fa3_17_f_u_arrmul24_and3_17_y0 & f_u_arrmul24_fa3_17_f_u_arrmul24_fa4_16_y2;
  assign f_u_arrmul24_fa3_17_y2 = f_u_arrmul24_fa3_17_y0 ^ f_u_arrmul24_fa3_17_f_u_arrmul24_fa2_17_y4;
  assign f_u_arrmul24_fa3_17_y3 = f_u_arrmul24_fa3_17_y0 & f_u_arrmul24_fa3_17_f_u_arrmul24_fa2_17_y4;
  assign f_u_arrmul24_fa3_17_y4 = f_u_arrmul24_fa3_17_y1 | f_u_arrmul24_fa3_17_y3;
  assign f_u_arrmul24_and4_17_a_4 = a_4;
  assign f_u_arrmul24_and4_17_b_17 = b_17;
  assign f_u_arrmul24_and4_17_y0 = f_u_arrmul24_and4_17_a_4 & f_u_arrmul24_and4_17_b_17;
  assign f_u_arrmul24_fa4_17_f_u_arrmul24_and4_17_y0 = f_u_arrmul24_and4_17_y0;
  assign f_u_arrmul24_fa4_17_f_u_arrmul24_fa5_16_y2 = f_u_arrmul24_fa5_16_y2;
  assign f_u_arrmul24_fa4_17_f_u_arrmul24_fa3_17_y4 = f_u_arrmul24_fa3_17_y4;
  assign f_u_arrmul24_fa4_17_y0 = f_u_arrmul24_fa4_17_f_u_arrmul24_and4_17_y0 ^ f_u_arrmul24_fa4_17_f_u_arrmul24_fa5_16_y2;
  assign f_u_arrmul24_fa4_17_y1 = f_u_arrmul24_fa4_17_f_u_arrmul24_and4_17_y0 & f_u_arrmul24_fa4_17_f_u_arrmul24_fa5_16_y2;
  assign f_u_arrmul24_fa4_17_y2 = f_u_arrmul24_fa4_17_y0 ^ f_u_arrmul24_fa4_17_f_u_arrmul24_fa3_17_y4;
  assign f_u_arrmul24_fa4_17_y3 = f_u_arrmul24_fa4_17_y0 & f_u_arrmul24_fa4_17_f_u_arrmul24_fa3_17_y4;
  assign f_u_arrmul24_fa4_17_y4 = f_u_arrmul24_fa4_17_y1 | f_u_arrmul24_fa4_17_y3;
  assign f_u_arrmul24_and5_17_a_5 = a_5;
  assign f_u_arrmul24_and5_17_b_17 = b_17;
  assign f_u_arrmul24_and5_17_y0 = f_u_arrmul24_and5_17_a_5 & f_u_arrmul24_and5_17_b_17;
  assign f_u_arrmul24_fa5_17_f_u_arrmul24_and5_17_y0 = f_u_arrmul24_and5_17_y0;
  assign f_u_arrmul24_fa5_17_f_u_arrmul24_fa6_16_y2 = f_u_arrmul24_fa6_16_y2;
  assign f_u_arrmul24_fa5_17_f_u_arrmul24_fa4_17_y4 = f_u_arrmul24_fa4_17_y4;
  assign f_u_arrmul24_fa5_17_y0 = f_u_arrmul24_fa5_17_f_u_arrmul24_and5_17_y0 ^ f_u_arrmul24_fa5_17_f_u_arrmul24_fa6_16_y2;
  assign f_u_arrmul24_fa5_17_y1 = f_u_arrmul24_fa5_17_f_u_arrmul24_and5_17_y0 & f_u_arrmul24_fa5_17_f_u_arrmul24_fa6_16_y2;
  assign f_u_arrmul24_fa5_17_y2 = f_u_arrmul24_fa5_17_y0 ^ f_u_arrmul24_fa5_17_f_u_arrmul24_fa4_17_y4;
  assign f_u_arrmul24_fa5_17_y3 = f_u_arrmul24_fa5_17_y0 & f_u_arrmul24_fa5_17_f_u_arrmul24_fa4_17_y4;
  assign f_u_arrmul24_fa5_17_y4 = f_u_arrmul24_fa5_17_y1 | f_u_arrmul24_fa5_17_y3;
  assign f_u_arrmul24_and6_17_a_6 = a_6;
  assign f_u_arrmul24_and6_17_b_17 = b_17;
  assign f_u_arrmul24_and6_17_y0 = f_u_arrmul24_and6_17_a_6 & f_u_arrmul24_and6_17_b_17;
  assign f_u_arrmul24_fa6_17_f_u_arrmul24_and6_17_y0 = f_u_arrmul24_and6_17_y0;
  assign f_u_arrmul24_fa6_17_f_u_arrmul24_fa7_16_y2 = f_u_arrmul24_fa7_16_y2;
  assign f_u_arrmul24_fa6_17_f_u_arrmul24_fa5_17_y4 = f_u_arrmul24_fa5_17_y4;
  assign f_u_arrmul24_fa6_17_y0 = f_u_arrmul24_fa6_17_f_u_arrmul24_and6_17_y0 ^ f_u_arrmul24_fa6_17_f_u_arrmul24_fa7_16_y2;
  assign f_u_arrmul24_fa6_17_y1 = f_u_arrmul24_fa6_17_f_u_arrmul24_and6_17_y0 & f_u_arrmul24_fa6_17_f_u_arrmul24_fa7_16_y2;
  assign f_u_arrmul24_fa6_17_y2 = f_u_arrmul24_fa6_17_y0 ^ f_u_arrmul24_fa6_17_f_u_arrmul24_fa5_17_y4;
  assign f_u_arrmul24_fa6_17_y3 = f_u_arrmul24_fa6_17_y0 & f_u_arrmul24_fa6_17_f_u_arrmul24_fa5_17_y4;
  assign f_u_arrmul24_fa6_17_y4 = f_u_arrmul24_fa6_17_y1 | f_u_arrmul24_fa6_17_y3;
  assign f_u_arrmul24_and7_17_a_7 = a_7;
  assign f_u_arrmul24_and7_17_b_17 = b_17;
  assign f_u_arrmul24_and7_17_y0 = f_u_arrmul24_and7_17_a_7 & f_u_arrmul24_and7_17_b_17;
  assign f_u_arrmul24_fa7_17_f_u_arrmul24_and7_17_y0 = f_u_arrmul24_and7_17_y0;
  assign f_u_arrmul24_fa7_17_f_u_arrmul24_fa8_16_y2 = f_u_arrmul24_fa8_16_y2;
  assign f_u_arrmul24_fa7_17_f_u_arrmul24_fa6_17_y4 = f_u_arrmul24_fa6_17_y4;
  assign f_u_arrmul24_fa7_17_y0 = f_u_arrmul24_fa7_17_f_u_arrmul24_and7_17_y0 ^ f_u_arrmul24_fa7_17_f_u_arrmul24_fa8_16_y2;
  assign f_u_arrmul24_fa7_17_y1 = f_u_arrmul24_fa7_17_f_u_arrmul24_and7_17_y0 & f_u_arrmul24_fa7_17_f_u_arrmul24_fa8_16_y2;
  assign f_u_arrmul24_fa7_17_y2 = f_u_arrmul24_fa7_17_y0 ^ f_u_arrmul24_fa7_17_f_u_arrmul24_fa6_17_y4;
  assign f_u_arrmul24_fa7_17_y3 = f_u_arrmul24_fa7_17_y0 & f_u_arrmul24_fa7_17_f_u_arrmul24_fa6_17_y4;
  assign f_u_arrmul24_fa7_17_y4 = f_u_arrmul24_fa7_17_y1 | f_u_arrmul24_fa7_17_y3;
  assign f_u_arrmul24_and8_17_a_8 = a_8;
  assign f_u_arrmul24_and8_17_b_17 = b_17;
  assign f_u_arrmul24_and8_17_y0 = f_u_arrmul24_and8_17_a_8 & f_u_arrmul24_and8_17_b_17;
  assign f_u_arrmul24_fa8_17_f_u_arrmul24_and8_17_y0 = f_u_arrmul24_and8_17_y0;
  assign f_u_arrmul24_fa8_17_f_u_arrmul24_fa9_16_y2 = f_u_arrmul24_fa9_16_y2;
  assign f_u_arrmul24_fa8_17_f_u_arrmul24_fa7_17_y4 = f_u_arrmul24_fa7_17_y4;
  assign f_u_arrmul24_fa8_17_y0 = f_u_arrmul24_fa8_17_f_u_arrmul24_and8_17_y0 ^ f_u_arrmul24_fa8_17_f_u_arrmul24_fa9_16_y2;
  assign f_u_arrmul24_fa8_17_y1 = f_u_arrmul24_fa8_17_f_u_arrmul24_and8_17_y0 & f_u_arrmul24_fa8_17_f_u_arrmul24_fa9_16_y2;
  assign f_u_arrmul24_fa8_17_y2 = f_u_arrmul24_fa8_17_y0 ^ f_u_arrmul24_fa8_17_f_u_arrmul24_fa7_17_y4;
  assign f_u_arrmul24_fa8_17_y3 = f_u_arrmul24_fa8_17_y0 & f_u_arrmul24_fa8_17_f_u_arrmul24_fa7_17_y4;
  assign f_u_arrmul24_fa8_17_y4 = f_u_arrmul24_fa8_17_y1 | f_u_arrmul24_fa8_17_y3;
  assign f_u_arrmul24_and9_17_a_9 = a_9;
  assign f_u_arrmul24_and9_17_b_17 = b_17;
  assign f_u_arrmul24_and9_17_y0 = f_u_arrmul24_and9_17_a_9 & f_u_arrmul24_and9_17_b_17;
  assign f_u_arrmul24_fa9_17_f_u_arrmul24_and9_17_y0 = f_u_arrmul24_and9_17_y0;
  assign f_u_arrmul24_fa9_17_f_u_arrmul24_fa10_16_y2 = f_u_arrmul24_fa10_16_y2;
  assign f_u_arrmul24_fa9_17_f_u_arrmul24_fa8_17_y4 = f_u_arrmul24_fa8_17_y4;
  assign f_u_arrmul24_fa9_17_y0 = f_u_arrmul24_fa9_17_f_u_arrmul24_and9_17_y0 ^ f_u_arrmul24_fa9_17_f_u_arrmul24_fa10_16_y2;
  assign f_u_arrmul24_fa9_17_y1 = f_u_arrmul24_fa9_17_f_u_arrmul24_and9_17_y0 & f_u_arrmul24_fa9_17_f_u_arrmul24_fa10_16_y2;
  assign f_u_arrmul24_fa9_17_y2 = f_u_arrmul24_fa9_17_y0 ^ f_u_arrmul24_fa9_17_f_u_arrmul24_fa8_17_y4;
  assign f_u_arrmul24_fa9_17_y3 = f_u_arrmul24_fa9_17_y0 & f_u_arrmul24_fa9_17_f_u_arrmul24_fa8_17_y4;
  assign f_u_arrmul24_fa9_17_y4 = f_u_arrmul24_fa9_17_y1 | f_u_arrmul24_fa9_17_y3;
  assign f_u_arrmul24_and10_17_a_10 = a_10;
  assign f_u_arrmul24_and10_17_b_17 = b_17;
  assign f_u_arrmul24_and10_17_y0 = f_u_arrmul24_and10_17_a_10 & f_u_arrmul24_and10_17_b_17;
  assign f_u_arrmul24_fa10_17_f_u_arrmul24_and10_17_y0 = f_u_arrmul24_and10_17_y0;
  assign f_u_arrmul24_fa10_17_f_u_arrmul24_fa11_16_y2 = f_u_arrmul24_fa11_16_y2;
  assign f_u_arrmul24_fa10_17_f_u_arrmul24_fa9_17_y4 = f_u_arrmul24_fa9_17_y4;
  assign f_u_arrmul24_fa10_17_y0 = f_u_arrmul24_fa10_17_f_u_arrmul24_and10_17_y0 ^ f_u_arrmul24_fa10_17_f_u_arrmul24_fa11_16_y2;
  assign f_u_arrmul24_fa10_17_y1 = f_u_arrmul24_fa10_17_f_u_arrmul24_and10_17_y0 & f_u_arrmul24_fa10_17_f_u_arrmul24_fa11_16_y2;
  assign f_u_arrmul24_fa10_17_y2 = f_u_arrmul24_fa10_17_y0 ^ f_u_arrmul24_fa10_17_f_u_arrmul24_fa9_17_y4;
  assign f_u_arrmul24_fa10_17_y3 = f_u_arrmul24_fa10_17_y0 & f_u_arrmul24_fa10_17_f_u_arrmul24_fa9_17_y4;
  assign f_u_arrmul24_fa10_17_y4 = f_u_arrmul24_fa10_17_y1 | f_u_arrmul24_fa10_17_y3;
  assign f_u_arrmul24_and11_17_a_11 = a_11;
  assign f_u_arrmul24_and11_17_b_17 = b_17;
  assign f_u_arrmul24_and11_17_y0 = f_u_arrmul24_and11_17_a_11 & f_u_arrmul24_and11_17_b_17;
  assign f_u_arrmul24_fa11_17_f_u_arrmul24_and11_17_y0 = f_u_arrmul24_and11_17_y0;
  assign f_u_arrmul24_fa11_17_f_u_arrmul24_fa12_16_y2 = f_u_arrmul24_fa12_16_y2;
  assign f_u_arrmul24_fa11_17_f_u_arrmul24_fa10_17_y4 = f_u_arrmul24_fa10_17_y4;
  assign f_u_arrmul24_fa11_17_y0 = f_u_arrmul24_fa11_17_f_u_arrmul24_and11_17_y0 ^ f_u_arrmul24_fa11_17_f_u_arrmul24_fa12_16_y2;
  assign f_u_arrmul24_fa11_17_y1 = f_u_arrmul24_fa11_17_f_u_arrmul24_and11_17_y0 & f_u_arrmul24_fa11_17_f_u_arrmul24_fa12_16_y2;
  assign f_u_arrmul24_fa11_17_y2 = f_u_arrmul24_fa11_17_y0 ^ f_u_arrmul24_fa11_17_f_u_arrmul24_fa10_17_y4;
  assign f_u_arrmul24_fa11_17_y3 = f_u_arrmul24_fa11_17_y0 & f_u_arrmul24_fa11_17_f_u_arrmul24_fa10_17_y4;
  assign f_u_arrmul24_fa11_17_y4 = f_u_arrmul24_fa11_17_y1 | f_u_arrmul24_fa11_17_y3;
  assign f_u_arrmul24_and12_17_a_12 = a_12;
  assign f_u_arrmul24_and12_17_b_17 = b_17;
  assign f_u_arrmul24_and12_17_y0 = f_u_arrmul24_and12_17_a_12 & f_u_arrmul24_and12_17_b_17;
  assign f_u_arrmul24_fa12_17_f_u_arrmul24_and12_17_y0 = f_u_arrmul24_and12_17_y0;
  assign f_u_arrmul24_fa12_17_f_u_arrmul24_fa13_16_y2 = f_u_arrmul24_fa13_16_y2;
  assign f_u_arrmul24_fa12_17_f_u_arrmul24_fa11_17_y4 = f_u_arrmul24_fa11_17_y4;
  assign f_u_arrmul24_fa12_17_y0 = f_u_arrmul24_fa12_17_f_u_arrmul24_and12_17_y0 ^ f_u_arrmul24_fa12_17_f_u_arrmul24_fa13_16_y2;
  assign f_u_arrmul24_fa12_17_y1 = f_u_arrmul24_fa12_17_f_u_arrmul24_and12_17_y0 & f_u_arrmul24_fa12_17_f_u_arrmul24_fa13_16_y2;
  assign f_u_arrmul24_fa12_17_y2 = f_u_arrmul24_fa12_17_y0 ^ f_u_arrmul24_fa12_17_f_u_arrmul24_fa11_17_y4;
  assign f_u_arrmul24_fa12_17_y3 = f_u_arrmul24_fa12_17_y0 & f_u_arrmul24_fa12_17_f_u_arrmul24_fa11_17_y4;
  assign f_u_arrmul24_fa12_17_y4 = f_u_arrmul24_fa12_17_y1 | f_u_arrmul24_fa12_17_y3;
  assign f_u_arrmul24_and13_17_a_13 = a_13;
  assign f_u_arrmul24_and13_17_b_17 = b_17;
  assign f_u_arrmul24_and13_17_y0 = f_u_arrmul24_and13_17_a_13 & f_u_arrmul24_and13_17_b_17;
  assign f_u_arrmul24_fa13_17_f_u_arrmul24_and13_17_y0 = f_u_arrmul24_and13_17_y0;
  assign f_u_arrmul24_fa13_17_f_u_arrmul24_fa14_16_y2 = f_u_arrmul24_fa14_16_y2;
  assign f_u_arrmul24_fa13_17_f_u_arrmul24_fa12_17_y4 = f_u_arrmul24_fa12_17_y4;
  assign f_u_arrmul24_fa13_17_y0 = f_u_arrmul24_fa13_17_f_u_arrmul24_and13_17_y0 ^ f_u_arrmul24_fa13_17_f_u_arrmul24_fa14_16_y2;
  assign f_u_arrmul24_fa13_17_y1 = f_u_arrmul24_fa13_17_f_u_arrmul24_and13_17_y0 & f_u_arrmul24_fa13_17_f_u_arrmul24_fa14_16_y2;
  assign f_u_arrmul24_fa13_17_y2 = f_u_arrmul24_fa13_17_y0 ^ f_u_arrmul24_fa13_17_f_u_arrmul24_fa12_17_y4;
  assign f_u_arrmul24_fa13_17_y3 = f_u_arrmul24_fa13_17_y0 & f_u_arrmul24_fa13_17_f_u_arrmul24_fa12_17_y4;
  assign f_u_arrmul24_fa13_17_y4 = f_u_arrmul24_fa13_17_y1 | f_u_arrmul24_fa13_17_y3;
  assign f_u_arrmul24_and14_17_a_14 = a_14;
  assign f_u_arrmul24_and14_17_b_17 = b_17;
  assign f_u_arrmul24_and14_17_y0 = f_u_arrmul24_and14_17_a_14 & f_u_arrmul24_and14_17_b_17;
  assign f_u_arrmul24_fa14_17_f_u_arrmul24_and14_17_y0 = f_u_arrmul24_and14_17_y0;
  assign f_u_arrmul24_fa14_17_f_u_arrmul24_fa15_16_y2 = f_u_arrmul24_fa15_16_y2;
  assign f_u_arrmul24_fa14_17_f_u_arrmul24_fa13_17_y4 = f_u_arrmul24_fa13_17_y4;
  assign f_u_arrmul24_fa14_17_y0 = f_u_arrmul24_fa14_17_f_u_arrmul24_and14_17_y0 ^ f_u_arrmul24_fa14_17_f_u_arrmul24_fa15_16_y2;
  assign f_u_arrmul24_fa14_17_y1 = f_u_arrmul24_fa14_17_f_u_arrmul24_and14_17_y0 & f_u_arrmul24_fa14_17_f_u_arrmul24_fa15_16_y2;
  assign f_u_arrmul24_fa14_17_y2 = f_u_arrmul24_fa14_17_y0 ^ f_u_arrmul24_fa14_17_f_u_arrmul24_fa13_17_y4;
  assign f_u_arrmul24_fa14_17_y3 = f_u_arrmul24_fa14_17_y0 & f_u_arrmul24_fa14_17_f_u_arrmul24_fa13_17_y4;
  assign f_u_arrmul24_fa14_17_y4 = f_u_arrmul24_fa14_17_y1 | f_u_arrmul24_fa14_17_y3;
  assign f_u_arrmul24_and15_17_a_15 = a_15;
  assign f_u_arrmul24_and15_17_b_17 = b_17;
  assign f_u_arrmul24_and15_17_y0 = f_u_arrmul24_and15_17_a_15 & f_u_arrmul24_and15_17_b_17;
  assign f_u_arrmul24_fa15_17_f_u_arrmul24_and15_17_y0 = f_u_arrmul24_and15_17_y0;
  assign f_u_arrmul24_fa15_17_f_u_arrmul24_fa16_16_y2 = f_u_arrmul24_fa16_16_y2;
  assign f_u_arrmul24_fa15_17_f_u_arrmul24_fa14_17_y4 = f_u_arrmul24_fa14_17_y4;
  assign f_u_arrmul24_fa15_17_y0 = f_u_arrmul24_fa15_17_f_u_arrmul24_and15_17_y0 ^ f_u_arrmul24_fa15_17_f_u_arrmul24_fa16_16_y2;
  assign f_u_arrmul24_fa15_17_y1 = f_u_arrmul24_fa15_17_f_u_arrmul24_and15_17_y0 & f_u_arrmul24_fa15_17_f_u_arrmul24_fa16_16_y2;
  assign f_u_arrmul24_fa15_17_y2 = f_u_arrmul24_fa15_17_y0 ^ f_u_arrmul24_fa15_17_f_u_arrmul24_fa14_17_y4;
  assign f_u_arrmul24_fa15_17_y3 = f_u_arrmul24_fa15_17_y0 & f_u_arrmul24_fa15_17_f_u_arrmul24_fa14_17_y4;
  assign f_u_arrmul24_fa15_17_y4 = f_u_arrmul24_fa15_17_y1 | f_u_arrmul24_fa15_17_y3;
  assign f_u_arrmul24_and16_17_a_16 = a_16;
  assign f_u_arrmul24_and16_17_b_17 = b_17;
  assign f_u_arrmul24_and16_17_y0 = f_u_arrmul24_and16_17_a_16 & f_u_arrmul24_and16_17_b_17;
  assign f_u_arrmul24_fa16_17_f_u_arrmul24_and16_17_y0 = f_u_arrmul24_and16_17_y0;
  assign f_u_arrmul24_fa16_17_f_u_arrmul24_fa17_16_y2 = f_u_arrmul24_fa17_16_y2;
  assign f_u_arrmul24_fa16_17_f_u_arrmul24_fa15_17_y4 = f_u_arrmul24_fa15_17_y4;
  assign f_u_arrmul24_fa16_17_y0 = f_u_arrmul24_fa16_17_f_u_arrmul24_and16_17_y0 ^ f_u_arrmul24_fa16_17_f_u_arrmul24_fa17_16_y2;
  assign f_u_arrmul24_fa16_17_y1 = f_u_arrmul24_fa16_17_f_u_arrmul24_and16_17_y0 & f_u_arrmul24_fa16_17_f_u_arrmul24_fa17_16_y2;
  assign f_u_arrmul24_fa16_17_y2 = f_u_arrmul24_fa16_17_y0 ^ f_u_arrmul24_fa16_17_f_u_arrmul24_fa15_17_y4;
  assign f_u_arrmul24_fa16_17_y3 = f_u_arrmul24_fa16_17_y0 & f_u_arrmul24_fa16_17_f_u_arrmul24_fa15_17_y4;
  assign f_u_arrmul24_fa16_17_y4 = f_u_arrmul24_fa16_17_y1 | f_u_arrmul24_fa16_17_y3;
  assign f_u_arrmul24_and17_17_a_17 = a_17;
  assign f_u_arrmul24_and17_17_b_17 = b_17;
  assign f_u_arrmul24_and17_17_y0 = f_u_arrmul24_and17_17_a_17 & f_u_arrmul24_and17_17_b_17;
  assign f_u_arrmul24_fa17_17_f_u_arrmul24_and17_17_y0 = f_u_arrmul24_and17_17_y0;
  assign f_u_arrmul24_fa17_17_f_u_arrmul24_fa18_16_y2 = f_u_arrmul24_fa18_16_y2;
  assign f_u_arrmul24_fa17_17_f_u_arrmul24_fa16_17_y4 = f_u_arrmul24_fa16_17_y4;
  assign f_u_arrmul24_fa17_17_y0 = f_u_arrmul24_fa17_17_f_u_arrmul24_and17_17_y0 ^ f_u_arrmul24_fa17_17_f_u_arrmul24_fa18_16_y2;
  assign f_u_arrmul24_fa17_17_y1 = f_u_arrmul24_fa17_17_f_u_arrmul24_and17_17_y0 & f_u_arrmul24_fa17_17_f_u_arrmul24_fa18_16_y2;
  assign f_u_arrmul24_fa17_17_y2 = f_u_arrmul24_fa17_17_y0 ^ f_u_arrmul24_fa17_17_f_u_arrmul24_fa16_17_y4;
  assign f_u_arrmul24_fa17_17_y3 = f_u_arrmul24_fa17_17_y0 & f_u_arrmul24_fa17_17_f_u_arrmul24_fa16_17_y4;
  assign f_u_arrmul24_fa17_17_y4 = f_u_arrmul24_fa17_17_y1 | f_u_arrmul24_fa17_17_y3;
  assign f_u_arrmul24_and18_17_a_18 = a_18;
  assign f_u_arrmul24_and18_17_b_17 = b_17;
  assign f_u_arrmul24_and18_17_y0 = f_u_arrmul24_and18_17_a_18 & f_u_arrmul24_and18_17_b_17;
  assign f_u_arrmul24_fa18_17_f_u_arrmul24_and18_17_y0 = f_u_arrmul24_and18_17_y0;
  assign f_u_arrmul24_fa18_17_f_u_arrmul24_fa19_16_y2 = f_u_arrmul24_fa19_16_y2;
  assign f_u_arrmul24_fa18_17_f_u_arrmul24_fa17_17_y4 = f_u_arrmul24_fa17_17_y4;
  assign f_u_arrmul24_fa18_17_y0 = f_u_arrmul24_fa18_17_f_u_arrmul24_and18_17_y0 ^ f_u_arrmul24_fa18_17_f_u_arrmul24_fa19_16_y2;
  assign f_u_arrmul24_fa18_17_y1 = f_u_arrmul24_fa18_17_f_u_arrmul24_and18_17_y0 & f_u_arrmul24_fa18_17_f_u_arrmul24_fa19_16_y2;
  assign f_u_arrmul24_fa18_17_y2 = f_u_arrmul24_fa18_17_y0 ^ f_u_arrmul24_fa18_17_f_u_arrmul24_fa17_17_y4;
  assign f_u_arrmul24_fa18_17_y3 = f_u_arrmul24_fa18_17_y0 & f_u_arrmul24_fa18_17_f_u_arrmul24_fa17_17_y4;
  assign f_u_arrmul24_fa18_17_y4 = f_u_arrmul24_fa18_17_y1 | f_u_arrmul24_fa18_17_y3;
  assign f_u_arrmul24_and19_17_a_19 = a_19;
  assign f_u_arrmul24_and19_17_b_17 = b_17;
  assign f_u_arrmul24_and19_17_y0 = f_u_arrmul24_and19_17_a_19 & f_u_arrmul24_and19_17_b_17;
  assign f_u_arrmul24_fa19_17_f_u_arrmul24_and19_17_y0 = f_u_arrmul24_and19_17_y0;
  assign f_u_arrmul24_fa19_17_f_u_arrmul24_fa20_16_y2 = f_u_arrmul24_fa20_16_y2;
  assign f_u_arrmul24_fa19_17_f_u_arrmul24_fa18_17_y4 = f_u_arrmul24_fa18_17_y4;
  assign f_u_arrmul24_fa19_17_y0 = f_u_arrmul24_fa19_17_f_u_arrmul24_and19_17_y0 ^ f_u_arrmul24_fa19_17_f_u_arrmul24_fa20_16_y2;
  assign f_u_arrmul24_fa19_17_y1 = f_u_arrmul24_fa19_17_f_u_arrmul24_and19_17_y0 & f_u_arrmul24_fa19_17_f_u_arrmul24_fa20_16_y2;
  assign f_u_arrmul24_fa19_17_y2 = f_u_arrmul24_fa19_17_y0 ^ f_u_arrmul24_fa19_17_f_u_arrmul24_fa18_17_y4;
  assign f_u_arrmul24_fa19_17_y3 = f_u_arrmul24_fa19_17_y0 & f_u_arrmul24_fa19_17_f_u_arrmul24_fa18_17_y4;
  assign f_u_arrmul24_fa19_17_y4 = f_u_arrmul24_fa19_17_y1 | f_u_arrmul24_fa19_17_y3;
  assign f_u_arrmul24_and20_17_a_20 = a_20;
  assign f_u_arrmul24_and20_17_b_17 = b_17;
  assign f_u_arrmul24_and20_17_y0 = f_u_arrmul24_and20_17_a_20 & f_u_arrmul24_and20_17_b_17;
  assign f_u_arrmul24_fa20_17_f_u_arrmul24_and20_17_y0 = f_u_arrmul24_and20_17_y0;
  assign f_u_arrmul24_fa20_17_f_u_arrmul24_fa21_16_y2 = f_u_arrmul24_fa21_16_y2;
  assign f_u_arrmul24_fa20_17_f_u_arrmul24_fa19_17_y4 = f_u_arrmul24_fa19_17_y4;
  assign f_u_arrmul24_fa20_17_y0 = f_u_arrmul24_fa20_17_f_u_arrmul24_and20_17_y0 ^ f_u_arrmul24_fa20_17_f_u_arrmul24_fa21_16_y2;
  assign f_u_arrmul24_fa20_17_y1 = f_u_arrmul24_fa20_17_f_u_arrmul24_and20_17_y0 & f_u_arrmul24_fa20_17_f_u_arrmul24_fa21_16_y2;
  assign f_u_arrmul24_fa20_17_y2 = f_u_arrmul24_fa20_17_y0 ^ f_u_arrmul24_fa20_17_f_u_arrmul24_fa19_17_y4;
  assign f_u_arrmul24_fa20_17_y3 = f_u_arrmul24_fa20_17_y0 & f_u_arrmul24_fa20_17_f_u_arrmul24_fa19_17_y4;
  assign f_u_arrmul24_fa20_17_y4 = f_u_arrmul24_fa20_17_y1 | f_u_arrmul24_fa20_17_y3;
  assign f_u_arrmul24_and21_17_a_21 = a_21;
  assign f_u_arrmul24_and21_17_b_17 = b_17;
  assign f_u_arrmul24_and21_17_y0 = f_u_arrmul24_and21_17_a_21 & f_u_arrmul24_and21_17_b_17;
  assign f_u_arrmul24_fa21_17_f_u_arrmul24_and21_17_y0 = f_u_arrmul24_and21_17_y0;
  assign f_u_arrmul24_fa21_17_f_u_arrmul24_fa22_16_y2 = f_u_arrmul24_fa22_16_y2;
  assign f_u_arrmul24_fa21_17_f_u_arrmul24_fa20_17_y4 = f_u_arrmul24_fa20_17_y4;
  assign f_u_arrmul24_fa21_17_y0 = f_u_arrmul24_fa21_17_f_u_arrmul24_and21_17_y0 ^ f_u_arrmul24_fa21_17_f_u_arrmul24_fa22_16_y2;
  assign f_u_arrmul24_fa21_17_y1 = f_u_arrmul24_fa21_17_f_u_arrmul24_and21_17_y0 & f_u_arrmul24_fa21_17_f_u_arrmul24_fa22_16_y2;
  assign f_u_arrmul24_fa21_17_y2 = f_u_arrmul24_fa21_17_y0 ^ f_u_arrmul24_fa21_17_f_u_arrmul24_fa20_17_y4;
  assign f_u_arrmul24_fa21_17_y3 = f_u_arrmul24_fa21_17_y0 & f_u_arrmul24_fa21_17_f_u_arrmul24_fa20_17_y4;
  assign f_u_arrmul24_fa21_17_y4 = f_u_arrmul24_fa21_17_y1 | f_u_arrmul24_fa21_17_y3;
  assign f_u_arrmul24_and22_17_a_22 = a_22;
  assign f_u_arrmul24_and22_17_b_17 = b_17;
  assign f_u_arrmul24_and22_17_y0 = f_u_arrmul24_and22_17_a_22 & f_u_arrmul24_and22_17_b_17;
  assign f_u_arrmul24_fa22_17_f_u_arrmul24_and22_17_y0 = f_u_arrmul24_and22_17_y0;
  assign f_u_arrmul24_fa22_17_f_u_arrmul24_fa23_16_y2 = f_u_arrmul24_fa23_16_y2;
  assign f_u_arrmul24_fa22_17_f_u_arrmul24_fa21_17_y4 = f_u_arrmul24_fa21_17_y4;
  assign f_u_arrmul24_fa22_17_y0 = f_u_arrmul24_fa22_17_f_u_arrmul24_and22_17_y0 ^ f_u_arrmul24_fa22_17_f_u_arrmul24_fa23_16_y2;
  assign f_u_arrmul24_fa22_17_y1 = f_u_arrmul24_fa22_17_f_u_arrmul24_and22_17_y0 & f_u_arrmul24_fa22_17_f_u_arrmul24_fa23_16_y2;
  assign f_u_arrmul24_fa22_17_y2 = f_u_arrmul24_fa22_17_y0 ^ f_u_arrmul24_fa22_17_f_u_arrmul24_fa21_17_y4;
  assign f_u_arrmul24_fa22_17_y3 = f_u_arrmul24_fa22_17_y0 & f_u_arrmul24_fa22_17_f_u_arrmul24_fa21_17_y4;
  assign f_u_arrmul24_fa22_17_y4 = f_u_arrmul24_fa22_17_y1 | f_u_arrmul24_fa22_17_y3;
  assign f_u_arrmul24_and23_17_a_23 = a_23;
  assign f_u_arrmul24_and23_17_b_17 = b_17;
  assign f_u_arrmul24_and23_17_y0 = f_u_arrmul24_and23_17_a_23 & f_u_arrmul24_and23_17_b_17;
  assign f_u_arrmul24_fa23_17_f_u_arrmul24_and23_17_y0 = f_u_arrmul24_and23_17_y0;
  assign f_u_arrmul24_fa23_17_f_u_arrmul24_fa23_16_y4 = f_u_arrmul24_fa23_16_y4;
  assign f_u_arrmul24_fa23_17_f_u_arrmul24_fa22_17_y4 = f_u_arrmul24_fa22_17_y4;
  assign f_u_arrmul24_fa23_17_y0 = f_u_arrmul24_fa23_17_f_u_arrmul24_and23_17_y0 ^ f_u_arrmul24_fa23_17_f_u_arrmul24_fa23_16_y4;
  assign f_u_arrmul24_fa23_17_y1 = f_u_arrmul24_fa23_17_f_u_arrmul24_and23_17_y0 & f_u_arrmul24_fa23_17_f_u_arrmul24_fa23_16_y4;
  assign f_u_arrmul24_fa23_17_y2 = f_u_arrmul24_fa23_17_y0 ^ f_u_arrmul24_fa23_17_f_u_arrmul24_fa22_17_y4;
  assign f_u_arrmul24_fa23_17_y3 = f_u_arrmul24_fa23_17_y0 & f_u_arrmul24_fa23_17_f_u_arrmul24_fa22_17_y4;
  assign f_u_arrmul24_fa23_17_y4 = f_u_arrmul24_fa23_17_y1 | f_u_arrmul24_fa23_17_y3;
  assign f_u_arrmul24_and0_18_a_0 = a_0;
  assign f_u_arrmul24_and0_18_b_18 = b_18;
  assign f_u_arrmul24_and0_18_y0 = f_u_arrmul24_and0_18_a_0 & f_u_arrmul24_and0_18_b_18;
  assign f_u_arrmul24_ha0_18_f_u_arrmul24_and0_18_y0 = f_u_arrmul24_and0_18_y0;
  assign f_u_arrmul24_ha0_18_f_u_arrmul24_fa1_17_y2 = f_u_arrmul24_fa1_17_y2;
  assign f_u_arrmul24_ha0_18_y0 = f_u_arrmul24_ha0_18_f_u_arrmul24_and0_18_y0 ^ f_u_arrmul24_ha0_18_f_u_arrmul24_fa1_17_y2;
  assign f_u_arrmul24_ha0_18_y1 = f_u_arrmul24_ha0_18_f_u_arrmul24_and0_18_y0 & f_u_arrmul24_ha0_18_f_u_arrmul24_fa1_17_y2;
  assign f_u_arrmul24_and1_18_a_1 = a_1;
  assign f_u_arrmul24_and1_18_b_18 = b_18;
  assign f_u_arrmul24_and1_18_y0 = f_u_arrmul24_and1_18_a_1 & f_u_arrmul24_and1_18_b_18;
  assign f_u_arrmul24_fa1_18_f_u_arrmul24_and1_18_y0 = f_u_arrmul24_and1_18_y0;
  assign f_u_arrmul24_fa1_18_f_u_arrmul24_fa2_17_y2 = f_u_arrmul24_fa2_17_y2;
  assign f_u_arrmul24_fa1_18_f_u_arrmul24_ha0_18_y1 = f_u_arrmul24_ha0_18_y1;
  assign f_u_arrmul24_fa1_18_y0 = f_u_arrmul24_fa1_18_f_u_arrmul24_and1_18_y0 ^ f_u_arrmul24_fa1_18_f_u_arrmul24_fa2_17_y2;
  assign f_u_arrmul24_fa1_18_y1 = f_u_arrmul24_fa1_18_f_u_arrmul24_and1_18_y0 & f_u_arrmul24_fa1_18_f_u_arrmul24_fa2_17_y2;
  assign f_u_arrmul24_fa1_18_y2 = f_u_arrmul24_fa1_18_y0 ^ f_u_arrmul24_fa1_18_f_u_arrmul24_ha0_18_y1;
  assign f_u_arrmul24_fa1_18_y3 = f_u_arrmul24_fa1_18_y0 & f_u_arrmul24_fa1_18_f_u_arrmul24_ha0_18_y1;
  assign f_u_arrmul24_fa1_18_y4 = f_u_arrmul24_fa1_18_y1 | f_u_arrmul24_fa1_18_y3;
  assign f_u_arrmul24_and2_18_a_2 = a_2;
  assign f_u_arrmul24_and2_18_b_18 = b_18;
  assign f_u_arrmul24_and2_18_y0 = f_u_arrmul24_and2_18_a_2 & f_u_arrmul24_and2_18_b_18;
  assign f_u_arrmul24_fa2_18_f_u_arrmul24_and2_18_y0 = f_u_arrmul24_and2_18_y0;
  assign f_u_arrmul24_fa2_18_f_u_arrmul24_fa3_17_y2 = f_u_arrmul24_fa3_17_y2;
  assign f_u_arrmul24_fa2_18_f_u_arrmul24_fa1_18_y4 = f_u_arrmul24_fa1_18_y4;
  assign f_u_arrmul24_fa2_18_y0 = f_u_arrmul24_fa2_18_f_u_arrmul24_and2_18_y0 ^ f_u_arrmul24_fa2_18_f_u_arrmul24_fa3_17_y2;
  assign f_u_arrmul24_fa2_18_y1 = f_u_arrmul24_fa2_18_f_u_arrmul24_and2_18_y0 & f_u_arrmul24_fa2_18_f_u_arrmul24_fa3_17_y2;
  assign f_u_arrmul24_fa2_18_y2 = f_u_arrmul24_fa2_18_y0 ^ f_u_arrmul24_fa2_18_f_u_arrmul24_fa1_18_y4;
  assign f_u_arrmul24_fa2_18_y3 = f_u_arrmul24_fa2_18_y0 & f_u_arrmul24_fa2_18_f_u_arrmul24_fa1_18_y4;
  assign f_u_arrmul24_fa2_18_y4 = f_u_arrmul24_fa2_18_y1 | f_u_arrmul24_fa2_18_y3;
  assign f_u_arrmul24_and3_18_a_3 = a_3;
  assign f_u_arrmul24_and3_18_b_18 = b_18;
  assign f_u_arrmul24_and3_18_y0 = f_u_arrmul24_and3_18_a_3 & f_u_arrmul24_and3_18_b_18;
  assign f_u_arrmul24_fa3_18_f_u_arrmul24_and3_18_y0 = f_u_arrmul24_and3_18_y0;
  assign f_u_arrmul24_fa3_18_f_u_arrmul24_fa4_17_y2 = f_u_arrmul24_fa4_17_y2;
  assign f_u_arrmul24_fa3_18_f_u_arrmul24_fa2_18_y4 = f_u_arrmul24_fa2_18_y4;
  assign f_u_arrmul24_fa3_18_y0 = f_u_arrmul24_fa3_18_f_u_arrmul24_and3_18_y0 ^ f_u_arrmul24_fa3_18_f_u_arrmul24_fa4_17_y2;
  assign f_u_arrmul24_fa3_18_y1 = f_u_arrmul24_fa3_18_f_u_arrmul24_and3_18_y0 & f_u_arrmul24_fa3_18_f_u_arrmul24_fa4_17_y2;
  assign f_u_arrmul24_fa3_18_y2 = f_u_arrmul24_fa3_18_y0 ^ f_u_arrmul24_fa3_18_f_u_arrmul24_fa2_18_y4;
  assign f_u_arrmul24_fa3_18_y3 = f_u_arrmul24_fa3_18_y0 & f_u_arrmul24_fa3_18_f_u_arrmul24_fa2_18_y4;
  assign f_u_arrmul24_fa3_18_y4 = f_u_arrmul24_fa3_18_y1 | f_u_arrmul24_fa3_18_y3;
  assign f_u_arrmul24_and4_18_a_4 = a_4;
  assign f_u_arrmul24_and4_18_b_18 = b_18;
  assign f_u_arrmul24_and4_18_y0 = f_u_arrmul24_and4_18_a_4 & f_u_arrmul24_and4_18_b_18;
  assign f_u_arrmul24_fa4_18_f_u_arrmul24_and4_18_y0 = f_u_arrmul24_and4_18_y0;
  assign f_u_arrmul24_fa4_18_f_u_arrmul24_fa5_17_y2 = f_u_arrmul24_fa5_17_y2;
  assign f_u_arrmul24_fa4_18_f_u_arrmul24_fa3_18_y4 = f_u_arrmul24_fa3_18_y4;
  assign f_u_arrmul24_fa4_18_y0 = f_u_arrmul24_fa4_18_f_u_arrmul24_and4_18_y0 ^ f_u_arrmul24_fa4_18_f_u_arrmul24_fa5_17_y2;
  assign f_u_arrmul24_fa4_18_y1 = f_u_arrmul24_fa4_18_f_u_arrmul24_and4_18_y0 & f_u_arrmul24_fa4_18_f_u_arrmul24_fa5_17_y2;
  assign f_u_arrmul24_fa4_18_y2 = f_u_arrmul24_fa4_18_y0 ^ f_u_arrmul24_fa4_18_f_u_arrmul24_fa3_18_y4;
  assign f_u_arrmul24_fa4_18_y3 = f_u_arrmul24_fa4_18_y0 & f_u_arrmul24_fa4_18_f_u_arrmul24_fa3_18_y4;
  assign f_u_arrmul24_fa4_18_y4 = f_u_arrmul24_fa4_18_y1 | f_u_arrmul24_fa4_18_y3;
  assign f_u_arrmul24_and5_18_a_5 = a_5;
  assign f_u_arrmul24_and5_18_b_18 = b_18;
  assign f_u_arrmul24_and5_18_y0 = f_u_arrmul24_and5_18_a_5 & f_u_arrmul24_and5_18_b_18;
  assign f_u_arrmul24_fa5_18_f_u_arrmul24_and5_18_y0 = f_u_arrmul24_and5_18_y0;
  assign f_u_arrmul24_fa5_18_f_u_arrmul24_fa6_17_y2 = f_u_arrmul24_fa6_17_y2;
  assign f_u_arrmul24_fa5_18_f_u_arrmul24_fa4_18_y4 = f_u_arrmul24_fa4_18_y4;
  assign f_u_arrmul24_fa5_18_y0 = f_u_arrmul24_fa5_18_f_u_arrmul24_and5_18_y0 ^ f_u_arrmul24_fa5_18_f_u_arrmul24_fa6_17_y2;
  assign f_u_arrmul24_fa5_18_y1 = f_u_arrmul24_fa5_18_f_u_arrmul24_and5_18_y0 & f_u_arrmul24_fa5_18_f_u_arrmul24_fa6_17_y2;
  assign f_u_arrmul24_fa5_18_y2 = f_u_arrmul24_fa5_18_y0 ^ f_u_arrmul24_fa5_18_f_u_arrmul24_fa4_18_y4;
  assign f_u_arrmul24_fa5_18_y3 = f_u_arrmul24_fa5_18_y0 & f_u_arrmul24_fa5_18_f_u_arrmul24_fa4_18_y4;
  assign f_u_arrmul24_fa5_18_y4 = f_u_arrmul24_fa5_18_y1 | f_u_arrmul24_fa5_18_y3;
  assign f_u_arrmul24_and6_18_a_6 = a_6;
  assign f_u_arrmul24_and6_18_b_18 = b_18;
  assign f_u_arrmul24_and6_18_y0 = f_u_arrmul24_and6_18_a_6 & f_u_arrmul24_and6_18_b_18;
  assign f_u_arrmul24_fa6_18_f_u_arrmul24_and6_18_y0 = f_u_arrmul24_and6_18_y0;
  assign f_u_arrmul24_fa6_18_f_u_arrmul24_fa7_17_y2 = f_u_arrmul24_fa7_17_y2;
  assign f_u_arrmul24_fa6_18_f_u_arrmul24_fa5_18_y4 = f_u_arrmul24_fa5_18_y4;
  assign f_u_arrmul24_fa6_18_y0 = f_u_arrmul24_fa6_18_f_u_arrmul24_and6_18_y0 ^ f_u_arrmul24_fa6_18_f_u_arrmul24_fa7_17_y2;
  assign f_u_arrmul24_fa6_18_y1 = f_u_arrmul24_fa6_18_f_u_arrmul24_and6_18_y0 & f_u_arrmul24_fa6_18_f_u_arrmul24_fa7_17_y2;
  assign f_u_arrmul24_fa6_18_y2 = f_u_arrmul24_fa6_18_y0 ^ f_u_arrmul24_fa6_18_f_u_arrmul24_fa5_18_y4;
  assign f_u_arrmul24_fa6_18_y3 = f_u_arrmul24_fa6_18_y0 & f_u_arrmul24_fa6_18_f_u_arrmul24_fa5_18_y4;
  assign f_u_arrmul24_fa6_18_y4 = f_u_arrmul24_fa6_18_y1 | f_u_arrmul24_fa6_18_y3;
  assign f_u_arrmul24_and7_18_a_7 = a_7;
  assign f_u_arrmul24_and7_18_b_18 = b_18;
  assign f_u_arrmul24_and7_18_y0 = f_u_arrmul24_and7_18_a_7 & f_u_arrmul24_and7_18_b_18;
  assign f_u_arrmul24_fa7_18_f_u_arrmul24_and7_18_y0 = f_u_arrmul24_and7_18_y0;
  assign f_u_arrmul24_fa7_18_f_u_arrmul24_fa8_17_y2 = f_u_arrmul24_fa8_17_y2;
  assign f_u_arrmul24_fa7_18_f_u_arrmul24_fa6_18_y4 = f_u_arrmul24_fa6_18_y4;
  assign f_u_arrmul24_fa7_18_y0 = f_u_arrmul24_fa7_18_f_u_arrmul24_and7_18_y0 ^ f_u_arrmul24_fa7_18_f_u_arrmul24_fa8_17_y2;
  assign f_u_arrmul24_fa7_18_y1 = f_u_arrmul24_fa7_18_f_u_arrmul24_and7_18_y0 & f_u_arrmul24_fa7_18_f_u_arrmul24_fa8_17_y2;
  assign f_u_arrmul24_fa7_18_y2 = f_u_arrmul24_fa7_18_y0 ^ f_u_arrmul24_fa7_18_f_u_arrmul24_fa6_18_y4;
  assign f_u_arrmul24_fa7_18_y3 = f_u_arrmul24_fa7_18_y0 & f_u_arrmul24_fa7_18_f_u_arrmul24_fa6_18_y4;
  assign f_u_arrmul24_fa7_18_y4 = f_u_arrmul24_fa7_18_y1 | f_u_arrmul24_fa7_18_y3;
  assign f_u_arrmul24_and8_18_a_8 = a_8;
  assign f_u_arrmul24_and8_18_b_18 = b_18;
  assign f_u_arrmul24_and8_18_y0 = f_u_arrmul24_and8_18_a_8 & f_u_arrmul24_and8_18_b_18;
  assign f_u_arrmul24_fa8_18_f_u_arrmul24_and8_18_y0 = f_u_arrmul24_and8_18_y0;
  assign f_u_arrmul24_fa8_18_f_u_arrmul24_fa9_17_y2 = f_u_arrmul24_fa9_17_y2;
  assign f_u_arrmul24_fa8_18_f_u_arrmul24_fa7_18_y4 = f_u_arrmul24_fa7_18_y4;
  assign f_u_arrmul24_fa8_18_y0 = f_u_arrmul24_fa8_18_f_u_arrmul24_and8_18_y0 ^ f_u_arrmul24_fa8_18_f_u_arrmul24_fa9_17_y2;
  assign f_u_arrmul24_fa8_18_y1 = f_u_arrmul24_fa8_18_f_u_arrmul24_and8_18_y0 & f_u_arrmul24_fa8_18_f_u_arrmul24_fa9_17_y2;
  assign f_u_arrmul24_fa8_18_y2 = f_u_arrmul24_fa8_18_y0 ^ f_u_arrmul24_fa8_18_f_u_arrmul24_fa7_18_y4;
  assign f_u_arrmul24_fa8_18_y3 = f_u_arrmul24_fa8_18_y0 & f_u_arrmul24_fa8_18_f_u_arrmul24_fa7_18_y4;
  assign f_u_arrmul24_fa8_18_y4 = f_u_arrmul24_fa8_18_y1 | f_u_arrmul24_fa8_18_y3;
  assign f_u_arrmul24_and9_18_a_9 = a_9;
  assign f_u_arrmul24_and9_18_b_18 = b_18;
  assign f_u_arrmul24_and9_18_y0 = f_u_arrmul24_and9_18_a_9 & f_u_arrmul24_and9_18_b_18;
  assign f_u_arrmul24_fa9_18_f_u_arrmul24_and9_18_y0 = f_u_arrmul24_and9_18_y0;
  assign f_u_arrmul24_fa9_18_f_u_arrmul24_fa10_17_y2 = f_u_arrmul24_fa10_17_y2;
  assign f_u_arrmul24_fa9_18_f_u_arrmul24_fa8_18_y4 = f_u_arrmul24_fa8_18_y4;
  assign f_u_arrmul24_fa9_18_y0 = f_u_arrmul24_fa9_18_f_u_arrmul24_and9_18_y0 ^ f_u_arrmul24_fa9_18_f_u_arrmul24_fa10_17_y2;
  assign f_u_arrmul24_fa9_18_y1 = f_u_arrmul24_fa9_18_f_u_arrmul24_and9_18_y0 & f_u_arrmul24_fa9_18_f_u_arrmul24_fa10_17_y2;
  assign f_u_arrmul24_fa9_18_y2 = f_u_arrmul24_fa9_18_y0 ^ f_u_arrmul24_fa9_18_f_u_arrmul24_fa8_18_y4;
  assign f_u_arrmul24_fa9_18_y3 = f_u_arrmul24_fa9_18_y0 & f_u_arrmul24_fa9_18_f_u_arrmul24_fa8_18_y4;
  assign f_u_arrmul24_fa9_18_y4 = f_u_arrmul24_fa9_18_y1 | f_u_arrmul24_fa9_18_y3;
  assign f_u_arrmul24_and10_18_a_10 = a_10;
  assign f_u_arrmul24_and10_18_b_18 = b_18;
  assign f_u_arrmul24_and10_18_y0 = f_u_arrmul24_and10_18_a_10 & f_u_arrmul24_and10_18_b_18;
  assign f_u_arrmul24_fa10_18_f_u_arrmul24_and10_18_y0 = f_u_arrmul24_and10_18_y0;
  assign f_u_arrmul24_fa10_18_f_u_arrmul24_fa11_17_y2 = f_u_arrmul24_fa11_17_y2;
  assign f_u_arrmul24_fa10_18_f_u_arrmul24_fa9_18_y4 = f_u_arrmul24_fa9_18_y4;
  assign f_u_arrmul24_fa10_18_y0 = f_u_arrmul24_fa10_18_f_u_arrmul24_and10_18_y0 ^ f_u_arrmul24_fa10_18_f_u_arrmul24_fa11_17_y2;
  assign f_u_arrmul24_fa10_18_y1 = f_u_arrmul24_fa10_18_f_u_arrmul24_and10_18_y0 & f_u_arrmul24_fa10_18_f_u_arrmul24_fa11_17_y2;
  assign f_u_arrmul24_fa10_18_y2 = f_u_arrmul24_fa10_18_y0 ^ f_u_arrmul24_fa10_18_f_u_arrmul24_fa9_18_y4;
  assign f_u_arrmul24_fa10_18_y3 = f_u_arrmul24_fa10_18_y0 & f_u_arrmul24_fa10_18_f_u_arrmul24_fa9_18_y4;
  assign f_u_arrmul24_fa10_18_y4 = f_u_arrmul24_fa10_18_y1 | f_u_arrmul24_fa10_18_y3;
  assign f_u_arrmul24_and11_18_a_11 = a_11;
  assign f_u_arrmul24_and11_18_b_18 = b_18;
  assign f_u_arrmul24_and11_18_y0 = f_u_arrmul24_and11_18_a_11 & f_u_arrmul24_and11_18_b_18;
  assign f_u_arrmul24_fa11_18_f_u_arrmul24_and11_18_y0 = f_u_arrmul24_and11_18_y0;
  assign f_u_arrmul24_fa11_18_f_u_arrmul24_fa12_17_y2 = f_u_arrmul24_fa12_17_y2;
  assign f_u_arrmul24_fa11_18_f_u_arrmul24_fa10_18_y4 = f_u_arrmul24_fa10_18_y4;
  assign f_u_arrmul24_fa11_18_y0 = f_u_arrmul24_fa11_18_f_u_arrmul24_and11_18_y0 ^ f_u_arrmul24_fa11_18_f_u_arrmul24_fa12_17_y2;
  assign f_u_arrmul24_fa11_18_y1 = f_u_arrmul24_fa11_18_f_u_arrmul24_and11_18_y0 & f_u_arrmul24_fa11_18_f_u_arrmul24_fa12_17_y2;
  assign f_u_arrmul24_fa11_18_y2 = f_u_arrmul24_fa11_18_y0 ^ f_u_arrmul24_fa11_18_f_u_arrmul24_fa10_18_y4;
  assign f_u_arrmul24_fa11_18_y3 = f_u_arrmul24_fa11_18_y0 & f_u_arrmul24_fa11_18_f_u_arrmul24_fa10_18_y4;
  assign f_u_arrmul24_fa11_18_y4 = f_u_arrmul24_fa11_18_y1 | f_u_arrmul24_fa11_18_y3;
  assign f_u_arrmul24_and12_18_a_12 = a_12;
  assign f_u_arrmul24_and12_18_b_18 = b_18;
  assign f_u_arrmul24_and12_18_y0 = f_u_arrmul24_and12_18_a_12 & f_u_arrmul24_and12_18_b_18;
  assign f_u_arrmul24_fa12_18_f_u_arrmul24_and12_18_y0 = f_u_arrmul24_and12_18_y0;
  assign f_u_arrmul24_fa12_18_f_u_arrmul24_fa13_17_y2 = f_u_arrmul24_fa13_17_y2;
  assign f_u_arrmul24_fa12_18_f_u_arrmul24_fa11_18_y4 = f_u_arrmul24_fa11_18_y4;
  assign f_u_arrmul24_fa12_18_y0 = f_u_arrmul24_fa12_18_f_u_arrmul24_and12_18_y0 ^ f_u_arrmul24_fa12_18_f_u_arrmul24_fa13_17_y2;
  assign f_u_arrmul24_fa12_18_y1 = f_u_arrmul24_fa12_18_f_u_arrmul24_and12_18_y0 & f_u_arrmul24_fa12_18_f_u_arrmul24_fa13_17_y2;
  assign f_u_arrmul24_fa12_18_y2 = f_u_arrmul24_fa12_18_y0 ^ f_u_arrmul24_fa12_18_f_u_arrmul24_fa11_18_y4;
  assign f_u_arrmul24_fa12_18_y3 = f_u_arrmul24_fa12_18_y0 & f_u_arrmul24_fa12_18_f_u_arrmul24_fa11_18_y4;
  assign f_u_arrmul24_fa12_18_y4 = f_u_arrmul24_fa12_18_y1 | f_u_arrmul24_fa12_18_y3;
  assign f_u_arrmul24_and13_18_a_13 = a_13;
  assign f_u_arrmul24_and13_18_b_18 = b_18;
  assign f_u_arrmul24_and13_18_y0 = f_u_arrmul24_and13_18_a_13 & f_u_arrmul24_and13_18_b_18;
  assign f_u_arrmul24_fa13_18_f_u_arrmul24_and13_18_y0 = f_u_arrmul24_and13_18_y0;
  assign f_u_arrmul24_fa13_18_f_u_arrmul24_fa14_17_y2 = f_u_arrmul24_fa14_17_y2;
  assign f_u_arrmul24_fa13_18_f_u_arrmul24_fa12_18_y4 = f_u_arrmul24_fa12_18_y4;
  assign f_u_arrmul24_fa13_18_y0 = f_u_arrmul24_fa13_18_f_u_arrmul24_and13_18_y0 ^ f_u_arrmul24_fa13_18_f_u_arrmul24_fa14_17_y2;
  assign f_u_arrmul24_fa13_18_y1 = f_u_arrmul24_fa13_18_f_u_arrmul24_and13_18_y0 & f_u_arrmul24_fa13_18_f_u_arrmul24_fa14_17_y2;
  assign f_u_arrmul24_fa13_18_y2 = f_u_arrmul24_fa13_18_y0 ^ f_u_arrmul24_fa13_18_f_u_arrmul24_fa12_18_y4;
  assign f_u_arrmul24_fa13_18_y3 = f_u_arrmul24_fa13_18_y0 & f_u_arrmul24_fa13_18_f_u_arrmul24_fa12_18_y4;
  assign f_u_arrmul24_fa13_18_y4 = f_u_arrmul24_fa13_18_y1 | f_u_arrmul24_fa13_18_y3;
  assign f_u_arrmul24_and14_18_a_14 = a_14;
  assign f_u_arrmul24_and14_18_b_18 = b_18;
  assign f_u_arrmul24_and14_18_y0 = f_u_arrmul24_and14_18_a_14 & f_u_arrmul24_and14_18_b_18;
  assign f_u_arrmul24_fa14_18_f_u_arrmul24_and14_18_y0 = f_u_arrmul24_and14_18_y0;
  assign f_u_arrmul24_fa14_18_f_u_arrmul24_fa15_17_y2 = f_u_arrmul24_fa15_17_y2;
  assign f_u_arrmul24_fa14_18_f_u_arrmul24_fa13_18_y4 = f_u_arrmul24_fa13_18_y4;
  assign f_u_arrmul24_fa14_18_y0 = f_u_arrmul24_fa14_18_f_u_arrmul24_and14_18_y0 ^ f_u_arrmul24_fa14_18_f_u_arrmul24_fa15_17_y2;
  assign f_u_arrmul24_fa14_18_y1 = f_u_arrmul24_fa14_18_f_u_arrmul24_and14_18_y0 & f_u_arrmul24_fa14_18_f_u_arrmul24_fa15_17_y2;
  assign f_u_arrmul24_fa14_18_y2 = f_u_arrmul24_fa14_18_y0 ^ f_u_arrmul24_fa14_18_f_u_arrmul24_fa13_18_y4;
  assign f_u_arrmul24_fa14_18_y3 = f_u_arrmul24_fa14_18_y0 & f_u_arrmul24_fa14_18_f_u_arrmul24_fa13_18_y4;
  assign f_u_arrmul24_fa14_18_y4 = f_u_arrmul24_fa14_18_y1 | f_u_arrmul24_fa14_18_y3;
  assign f_u_arrmul24_and15_18_a_15 = a_15;
  assign f_u_arrmul24_and15_18_b_18 = b_18;
  assign f_u_arrmul24_and15_18_y0 = f_u_arrmul24_and15_18_a_15 & f_u_arrmul24_and15_18_b_18;
  assign f_u_arrmul24_fa15_18_f_u_arrmul24_and15_18_y0 = f_u_arrmul24_and15_18_y0;
  assign f_u_arrmul24_fa15_18_f_u_arrmul24_fa16_17_y2 = f_u_arrmul24_fa16_17_y2;
  assign f_u_arrmul24_fa15_18_f_u_arrmul24_fa14_18_y4 = f_u_arrmul24_fa14_18_y4;
  assign f_u_arrmul24_fa15_18_y0 = f_u_arrmul24_fa15_18_f_u_arrmul24_and15_18_y0 ^ f_u_arrmul24_fa15_18_f_u_arrmul24_fa16_17_y2;
  assign f_u_arrmul24_fa15_18_y1 = f_u_arrmul24_fa15_18_f_u_arrmul24_and15_18_y0 & f_u_arrmul24_fa15_18_f_u_arrmul24_fa16_17_y2;
  assign f_u_arrmul24_fa15_18_y2 = f_u_arrmul24_fa15_18_y0 ^ f_u_arrmul24_fa15_18_f_u_arrmul24_fa14_18_y4;
  assign f_u_arrmul24_fa15_18_y3 = f_u_arrmul24_fa15_18_y0 & f_u_arrmul24_fa15_18_f_u_arrmul24_fa14_18_y4;
  assign f_u_arrmul24_fa15_18_y4 = f_u_arrmul24_fa15_18_y1 | f_u_arrmul24_fa15_18_y3;
  assign f_u_arrmul24_and16_18_a_16 = a_16;
  assign f_u_arrmul24_and16_18_b_18 = b_18;
  assign f_u_arrmul24_and16_18_y0 = f_u_arrmul24_and16_18_a_16 & f_u_arrmul24_and16_18_b_18;
  assign f_u_arrmul24_fa16_18_f_u_arrmul24_and16_18_y0 = f_u_arrmul24_and16_18_y0;
  assign f_u_arrmul24_fa16_18_f_u_arrmul24_fa17_17_y2 = f_u_arrmul24_fa17_17_y2;
  assign f_u_arrmul24_fa16_18_f_u_arrmul24_fa15_18_y4 = f_u_arrmul24_fa15_18_y4;
  assign f_u_arrmul24_fa16_18_y0 = f_u_arrmul24_fa16_18_f_u_arrmul24_and16_18_y0 ^ f_u_arrmul24_fa16_18_f_u_arrmul24_fa17_17_y2;
  assign f_u_arrmul24_fa16_18_y1 = f_u_arrmul24_fa16_18_f_u_arrmul24_and16_18_y0 & f_u_arrmul24_fa16_18_f_u_arrmul24_fa17_17_y2;
  assign f_u_arrmul24_fa16_18_y2 = f_u_arrmul24_fa16_18_y0 ^ f_u_arrmul24_fa16_18_f_u_arrmul24_fa15_18_y4;
  assign f_u_arrmul24_fa16_18_y3 = f_u_arrmul24_fa16_18_y0 & f_u_arrmul24_fa16_18_f_u_arrmul24_fa15_18_y4;
  assign f_u_arrmul24_fa16_18_y4 = f_u_arrmul24_fa16_18_y1 | f_u_arrmul24_fa16_18_y3;
  assign f_u_arrmul24_and17_18_a_17 = a_17;
  assign f_u_arrmul24_and17_18_b_18 = b_18;
  assign f_u_arrmul24_and17_18_y0 = f_u_arrmul24_and17_18_a_17 & f_u_arrmul24_and17_18_b_18;
  assign f_u_arrmul24_fa17_18_f_u_arrmul24_and17_18_y0 = f_u_arrmul24_and17_18_y0;
  assign f_u_arrmul24_fa17_18_f_u_arrmul24_fa18_17_y2 = f_u_arrmul24_fa18_17_y2;
  assign f_u_arrmul24_fa17_18_f_u_arrmul24_fa16_18_y4 = f_u_arrmul24_fa16_18_y4;
  assign f_u_arrmul24_fa17_18_y0 = f_u_arrmul24_fa17_18_f_u_arrmul24_and17_18_y0 ^ f_u_arrmul24_fa17_18_f_u_arrmul24_fa18_17_y2;
  assign f_u_arrmul24_fa17_18_y1 = f_u_arrmul24_fa17_18_f_u_arrmul24_and17_18_y0 & f_u_arrmul24_fa17_18_f_u_arrmul24_fa18_17_y2;
  assign f_u_arrmul24_fa17_18_y2 = f_u_arrmul24_fa17_18_y0 ^ f_u_arrmul24_fa17_18_f_u_arrmul24_fa16_18_y4;
  assign f_u_arrmul24_fa17_18_y3 = f_u_arrmul24_fa17_18_y0 & f_u_arrmul24_fa17_18_f_u_arrmul24_fa16_18_y4;
  assign f_u_arrmul24_fa17_18_y4 = f_u_arrmul24_fa17_18_y1 | f_u_arrmul24_fa17_18_y3;
  assign f_u_arrmul24_and18_18_a_18 = a_18;
  assign f_u_arrmul24_and18_18_b_18 = b_18;
  assign f_u_arrmul24_and18_18_y0 = f_u_arrmul24_and18_18_a_18 & f_u_arrmul24_and18_18_b_18;
  assign f_u_arrmul24_fa18_18_f_u_arrmul24_and18_18_y0 = f_u_arrmul24_and18_18_y0;
  assign f_u_arrmul24_fa18_18_f_u_arrmul24_fa19_17_y2 = f_u_arrmul24_fa19_17_y2;
  assign f_u_arrmul24_fa18_18_f_u_arrmul24_fa17_18_y4 = f_u_arrmul24_fa17_18_y4;
  assign f_u_arrmul24_fa18_18_y0 = f_u_arrmul24_fa18_18_f_u_arrmul24_and18_18_y0 ^ f_u_arrmul24_fa18_18_f_u_arrmul24_fa19_17_y2;
  assign f_u_arrmul24_fa18_18_y1 = f_u_arrmul24_fa18_18_f_u_arrmul24_and18_18_y0 & f_u_arrmul24_fa18_18_f_u_arrmul24_fa19_17_y2;
  assign f_u_arrmul24_fa18_18_y2 = f_u_arrmul24_fa18_18_y0 ^ f_u_arrmul24_fa18_18_f_u_arrmul24_fa17_18_y4;
  assign f_u_arrmul24_fa18_18_y3 = f_u_arrmul24_fa18_18_y0 & f_u_arrmul24_fa18_18_f_u_arrmul24_fa17_18_y4;
  assign f_u_arrmul24_fa18_18_y4 = f_u_arrmul24_fa18_18_y1 | f_u_arrmul24_fa18_18_y3;
  assign f_u_arrmul24_and19_18_a_19 = a_19;
  assign f_u_arrmul24_and19_18_b_18 = b_18;
  assign f_u_arrmul24_and19_18_y0 = f_u_arrmul24_and19_18_a_19 & f_u_arrmul24_and19_18_b_18;
  assign f_u_arrmul24_fa19_18_f_u_arrmul24_and19_18_y0 = f_u_arrmul24_and19_18_y0;
  assign f_u_arrmul24_fa19_18_f_u_arrmul24_fa20_17_y2 = f_u_arrmul24_fa20_17_y2;
  assign f_u_arrmul24_fa19_18_f_u_arrmul24_fa18_18_y4 = f_u_arrmul24_fa18_18_y4;
  assign f_u_arrmul24_fa19_18_y0 = f_u_arrmul24_fa19_18_f_u_arrmul24_and19_18_y0 ^ f_u_arrmul24_fa19_18_f_u_arrmul24_fa20_17_y2;
  assign f_u_arrmul24_fa19_18_y1 = f_u_arrmul24_fa19_18_f_u_arrmul24_and19_18_y0 & f_u_arrmul24_fa19_18_f_u_arrmul24_fa20_17_y2;
  assign f_u_arrmul24_fa19_18_y2 = f_u_arrmul24_fa19_18_y0 ^ f_u_arrmul24_fa19_18_f_u_arrmul24_fa18_18_y4;
  assign f_u_arrmul24_fa19_18_y3 = f_u_arrmul24_fa19_18_y0 & f_u_arrmul24_fa19_18_f_u_arrmul24_fa18_18_y4;
  assign f_u_arrmul24_fa19_18_y4 = f_u_arrmul24_fa19_18_y1 | f_u_arrmul24_fa19_18_y3;
  assign f_u_arrmul24_and20_18_a_20 = a_20;
  assign f_u_arrmul24_and20_18_b_18 = b_18;
  assign f_u_arrmul24_and20_18_y0 = f_u_arrmul24_and20_18_a_20 & f_u_arrmul24_and20_18_b_18;
  assign f_u_arrmul24_fa20_18_f_u_arrmul24_and20_18_y0 = f_u_arrmul24_and20_18_y0;
  assign f_u_arrmul24_fa20_18_f_u_arrmul24_fa21_17_y2 = f_u_arrmul24_fa21_17_y2;
  assign f_u_arrmul24_fa20_18_f_u_arrmul24_fa19_18_y4 = f_u_arrmul24_fa19_18_y4;
  assign f_u_arrmul24_fa20_18_y0 = f_u_arrmul24_fa20_18_f_u_arrmul24_and20_18_y0 ^ f_u_arrmul24_fa20_18_f_u_arrmul24_fa21_17_y2;
  assign f_u_arrmul24_fa20_18_y1 = f_u_arrmul24_fa20_18_f_u_arrmul24_and20_18_y0 & f_u_arrmul24_fa20_18_f_u_arrmul24_fa21_17_y2;
  assign f_u_arrmul24_fa20_18_y2 = f_u_arrmul24_fa20_18_y0 ^ f_u_arrmul24_fa20_18_f_u_arrmul24_fa19_18_y4;
  assign f_u_arrmul24_fa20_18_y3 = f_u_arrmul24_fa20_18_y0 & f_u_arrmul24_fa20_18_f_u_arrmul24_fa19_18_y4;
  assign f_u_arrmul24_fa20_18_y4 = f_u_arrmul24_fa20_18_y1 | f_u_arrmul24_fa20_18_y3;
  assign f_u_arrmul24_and21_18_a_21 = a_21;
  assign f_u_arrmul24_and21_18_b_18 = b_18;
  assign f_u_arrmul24_and21_18_y0 = f_u_arrmul24_and21_18_a_21 & f_u_arrmul24_and21_18_b_18;
  assign f_u_arrmul24_fa21_18_f_u_arrmul24_and21_18_y0 = f_u_arrmul24_and21_18_y0;
  assign f_u_arrmul24_fa21_18_f_u_arrmul24_fa22_17_y2 = f_u_arrmul24_fa22_17_y2;
  assign f_u_arrmul24_fa21_18_f_u_arrmul24_fa20_18_y4 = f_u_arrmul24_fa20_18_y4;
  assign f_u_arrmul24_fa21_18_y0 = f_u_arrmul24_fa21_18_f_u_arrmul24_and21_18_y0 ^ f_u_arrmul24_fa21_18_f_u_arrmul24_fa22_17_y2;
  assign f_u_arrmul24_fa21_18_y1 = f_u_arrmul24_fa21_18_f_u_arrmul24_and21_18_y0 & f_u_arrmul24_fa21_18_f_u_arrmul24_fa22_17_y2;
  assign f_u_arrmul24_fa21_18_y2 = f_u_arrmul24_fa21_18_y0 ^ f_u_arrmul24_fa21_18_f_u_arrmul24_fa20_18_y4;
  assign f_u_arrmul24_fa21_18_y3 = f_u_arrmul24_fa21_18_y0 & f_u_arrmul24_fa21_18_f_u_arrmul24_fa20_18_y4;
  assign f_u_arrmul24_fa21_18_y4 = f_u_arrmul24_fa21_18_y1 | f_u_arrmul24_fa21_18_y3;
  assign f_u_arrmul24_and22_18_a_22 = a_22;
  assign f_u_arrmul24_and22_18_b_18 = b_18;
  assign f_u_arrmul24_and22_18_y0 = f_u_arrmul24_and22_18_a_22 & f_u_arrmul24_and22_18_b_18;
  assign f_u_arrmul24_fa22_18_f_u_arrmul24_and22_18_y0 = f_u_arrmul24_and22_18_y0;
  assign f_u_arrmul24_fa22_18_f_u_arrmul24_fa23_17_y2 = f_u_arrmul24_fa23_17_y2;
  assign f_u_arrmul24_fa22_18_f_u_arrmul24_fa21_18_y4 = f_u_arrmul24_fa21_18_y4;
  assign f_u_arrmul24_fa22_18_y0 = f_u_arrmul24_fa22_18_f_u_arrmul24_and22_18_y0 ^ f_u_arrmul24_fa22_18_f_u_arrmul24_fa23_17_y2;
  assign f_u_arrmul24_fa22_18_y1 = f_u_arrmul24_fa22_18_f_u_arrmul24_and22_18_y0 & f_u_arrmul24_fa22_18_f_u_arrmul24_fa23_17_y2;
  assign f_u_arrmul24_fa22_18_y2 = f_u_arrmul24_fa22_18_y0 ^ f_u_arrmul24_fa22_18_f_u_arrmul24_fa21_18_y4;
  assign f_u_arrmul24_fa22_18_y3 = f_u_arrmul24_fa22_18_y0 & f_u_arrmul24_fa22_18_f_u_arrmul24_fa21_18_y4;
  assign f_u_arrmul24_fa22_18_y4 = f_u_arrmul24_fa22_18_y1 | f_u_arrmul24_fa22_18_y3;
  assign f_u_arrmul24_and23_18_a_23 = a_23;
  assign f_u_arrmul24_and23_18_b_18 = b_18;
  assign f_u_arrmul24_and23_18_y0 = f_u_arrmul24_and23_18_a_23 & f_u_arrmul24_and23_18_b_18;
  assign f_u_arrmul24_fa23_18_f_u_arrmul24_and23_18_y0 = f_u_arrmul24_and23_18_y0;
  assign f_u_arrmul24_fa23_18_f_u_arrmul24_fa23_17_y4 = f_u_arrmul24_fa23_17_y4;
  assign f_u_arrmul24_fa23_18_f_u_arrmul24_fa22_18_y4 = f_u_arrmul24_fa22_18_y4;
  assign f_u_arrmul24_fa23_18_y0 = f_u_arrmul24_fa23_18_f_u_arrmul24_and23_18_y0 ^ f_u_arrmul24_fa23_18_f_u_arrmul24_fa23_17_y4;
  assign f_u_arrmul24_fa23_18_y1 = f_u_arrmul24_fa23_18_f_u_arrmul24_and23_18_y0 & f_u_arrmul24_fa23_18_f_u_arrmul24_fa23_17_y4;
  assign f_u_arrmul24_fa23_18_y2 = f_u_arrmul24_fa23_18_y0 ^ f_u_arrmul24_fa23_18_f_u_arrmul24_fa22_18_y4;
  assign f_u_arrmul24_fa23_18_y3 = f_u_arrmul24_fa23_18_y0 & f_u_arrmul24_fa23_18_f_u_arrmul24_fa22_18_y4;
  assign f_u_arrmul24_fa23_18_y4 = f_u_arrmul24_fa23_18_y1 | f_u_arrmul24_fa23_18_y3;
  assign f_u_arrmul24_and0_19_a_0 = a_0;
  assign f_u_arrmul24_and0_19_b_19 = b_19;
  assign f_u_arrmul24_and0_19_y0 = f_u_arrmul24_and0_19_a_0 & f_u_arrmul24_and0_19_b_19;
  assign f_u_arrmul24_ha0_19_f_u_arrmul24_and0_19_y0 = f_u_arrmul24_and0_19_y0;
  assign f_u_arrmul24_ha0_19_f_u_arrmul24_fa1_18_y2 = f_u_arrmul24_fa1_18_y2;
  assign f_u_arrmul24_ha0_19_y0 = f_u_arrmul24_ha0_19_f_u_arrmul24_and0_19_y0 ^ f_u_arrmul24_ha0_19_f_u_arrmul24_fa1_18_y2;
  assign f_u_arrmul24_ha0_19_y1 = f_u_arrmul24_ha0_19_f_u_arrmul24_and0_19_y0 & f_u_arrmul24_ha0_19_f_u_arrmul24_fa1_18_y2;
  assign f_u_arrmul24_and1_19_a_1 = a_1;
  assign f_u_arrmul24_and1_19_b_19 = b_19;
  assign f_u_arrmul24_and1_19_y0 = f_u_arrmul24_and1_19_a_1 & f_u_arrmul24_and1_19_b_19;
  assign f_u_arrmul24_fa1_19_f_u_arrmul24_and1_19_y0 = f_u_arrmul24_and1_19_y0;
  assign f_u_arrmul24_fa1_19_f_u_arrmul24_fa2_18_y2 = f_u_arrmul24_fa2_18_y2;
  assign f_u_arrmul24_fa1_19_f_u_arrmul24_ha0_19_y1 = f_u_arrmul24_ha0_19_y1;
  assign f_u_arrmul24_fa1_19_y0 = f_u_arrmul24_fa1_19_f_u_arrmul24_and1_19_y0 ^ f_u_arrmul24_fa1_19_f_u_arrmul24_fa2_18_y2;
  assign f_u_arrmul24_fa1_19_y1 = f_u_arrmul24_fa1_19_f_u_arrmul24_and1_19_y0 & f_u_arrmul24_fa1_19_f_u_arrmul24_fa2_18_y2;
  assign f_u_arrmul24_fa1_19_y2 = f_u_arrmul24_fa1_19_y0 ^ f_u_arrmul24_fa1_19_f_u_arrmul24_ha0_19_y1;
  assign f_u_arrmul24_fa1_19_y3 = f_u_arrmul24_fa1_19_y0 & f_u_arrmul24_fa1_19_f_u_arrmul24_ha0_19_y1;
  assign f_u_arrmul24_fa1_19_y4 = f_u_arrmul24_fa1_19_y1 | f_u_arrmul24_fa1_19_y3;
  assign f_u_arrmul24_and2_19_a_2 = a_2;
  assign f_u_arrmul24_and2_19_b_19 = b_19;
  assign f_u_arrmul24_and2_19_y0 = f_u_arrmul24_and2_19_a_2 & f_u_arrmul24_and2_19_b_19;
  assign f_u_arrmul24_fa2_19_f_u_arrmul24_and2_19_y0 = f_u_arrmul24_and2_19_y0;
  assign f_u_arrmul24_fa2_19_f_u_arrmul24_fa3_18_y2 = f_u_arrmul24_fa3_18_y2;
  assign f_u_arrmul24_fa2_19_f_u_arrmul24_fa1_19_y4 = f_u_arrmul24_fa1_19_y4;
  assign f_u_arrmul24_fa2_19_y0 = f_u_arrmul24_fa2_19_f_u_arrmul24_and2_19_y0 ^ f_u_arrmul24_fa2_19_f_u_arrmul24_fa3_18_y2;
  assign f_u_arrmul24_fa2_19_y1 = f_u_arrmul24_fa2_19_f_u_arrmul24_and2_19_y0 & f_u_arrmul24_fa2_19_f_u_arrmul24_fa3_18_y2;
  assign f_u_arrmul24_fa2_19_y2 = f_u_arrmul24_fa2_19_y0 ^ f_u_arrmul24_fa2_19_f_u_arrmul24_fa1_19_y4;
  assign f_u_arrmul24_fa2_19_y3 = f_u_arrmul24_fa2_19_y0 & f_u_arrmul24_fa2_19_f_u_arrmul24_fa1_19_y4;
  assign f_u_arrmul24_fa2_19_y4 = f_u_arrmul24_fa2_19_y1 | f_u_arrmul24_fa2_19_y3;
  assign f_u_arrmul24_and3_19_a_3 = a_3;
  assign f_u_arrmul24_and3_19_b_19 = b_19;
  assign f_u_arrmul24_and3_19_y0 = f_u_arrmul24_and3_19_a_3 & f_u_arrmul24_and3_19_b_19;
  assign f_u_arrmul24_fa3_19_f_u_arrmul24_and3_19_y0 = f_u_arrmul24_and3_19_y0;
  assign f_u_arrmul24_fa3_19_f_u_arrmul24_fa4_18_y2 = f_u_arrmul24_fa4_18_y2;
  assign f_u_arrmul24_fa3_19_f_u_arrmul24_fa2_19_y4 = f_u_arrmul24_fa2_19_y4;
  assign f_u_arrmul24_fa3_19_y0 = f_u_arrmul24_fa3_19_f_u_arrmul24_and3_19_y0 ^ f_u_arrmul24_fa3_19_f_u_arrmul24_fa4_18_y2;
  assign f_u_arrmul24_fa3_19_y1 = f_u_arrmul24_fa3_19_f_u_arrmul24_and3_19_y0 & f_u_arrmul24_fa3_19_f_u_arrmul24_fa4_18_y2;
  assign f_u_arrmul24_fa3_19_y2 = f_u_arrmul24_fa3_19_y0 ^ f_u_arrmul24_fa3_19_f_u_arrmul24_fa2_19_y4;
  assign f_u_arrmul24_fa3_19_y3 = f_u_arrmul24_fa3_19_y0 & f_u_arrmul24_fa3_19_f_u_arrmul24_fa2_19_y4;
  assign f_u_arrmul24_fa3_19_y4 = f_u_arrmul24_fa3_19_y1 | f_u_arrmul24_fa3_19_y3;
  assign f_u_arrmul24_and4_19_a_4 = a_4;
  assign f_u_arrmul24_and4_19_b_19 = b_19;
  assign f_u_arrmul24_and4_19_y0 = f_u_arrmul24_and4_19_a_4 & f_u_arrmul24_and4_19_b_19;
  assign f_u_arrmul24_fa4_19_f_u_arrmul24_and4_19_y0 = f_u_arrmul24_and4_19_y0;
  assign f_u_arrmul24_fa4_19_f_u_arrmul24_fa5_18_y2 = f_u_arrmul24_fa5_18_y2;
  assign f_u_arrmul24_fa4_19_f_u_arrmul24_fa3_19_y4 = f_u_arrmul24_fa3_19_y4;
  assign f_u_arrmul24_fa4_19_y0 = f_u_arrmul24_fa4_19_f_u_arrmul24_and4_19_y0 ^ f_u_arrmul24_fa4_19_f_u_arrmul24_fa5_18_y2;
  assign f_u_arrmul24_fa4_19_y1 = f_u_arrmul24_fa4_19_f_u_arrmul24_and4_19_y0 & f_u_arrmul24_fa4_19_f_u_arrmul24_fa5_18_y2;
  assign f_u_arrmul24_fa4_19_y2 = f_u_arrmul24_fa4_19_y0 ^ f_u_arrmul24_fa4_19_f_u_arrmul24_fa3_19_y4;
  assign f_u_arrmul24_fa4_19_y3 = f_u_arrmul24_fa4_19_y0 & f_u_arrmul24_fa4_19_f_u_arrmul24_fa3_19_y4;
  assign f_u_arrmul24_fa4_19_y4 = f_u_arrmul24_fa4_19_y1 | f_u_arrmul24_fa4_19_y3;
  assign f_u_arrmul24_and5_19_a_5 = a_5;
  assign f_u_arrmul24_and5_19_b_19 = b_19;
  assign f_u_arrmul24_and5_19_y0 = f_u_arrmul24_and5_19_a_5 & f_u_arrmul24_and5_19_b_19;
  assign f_u_arrmul24_fa5_19_f_u_arrmul24_and5_19_y0 = f_u_arrmul24_and5_19_y0;
  assign f_u_arrmul24_fa5_19_f_u_arrmul24_fa6_18_y2 = f_u_arrmul24_fa6_18_y2;
  assign f_u_arrmul24_fa5_19_f_u_arrmul24_fa4_19_y4 = f_u_arrmul24_fa4_19_y4;
  assign f_u_arrmul24_fa5_19_y0 = f_u_arrmul24_fa5_19_f_u_arrmul24_and5_19_y0 ^ f_u_arrmul24_fa5_19_f_u_arrmul24_fa6_18_y2;
  assign f_u_arrmul24_fa5_19_y1 = f_u_arrmul24_fa5_19_f_u_arrmul24_and5_19_y0 & f_u_arrmul24_fa5_19_f_u_arrmul24_fa6_18_y2;
  assign f_u_arrmul24_fa5_19_y2 = f_u_arrmul24_fa5_19_y0 ^ f_u_arrmul24_fa5_19_f_u_arrmul24_fa4_19_y4;
  assign f_u_arrmul24_fa5_19_y3 = f_u_arrmul24_fa5_19_y0 & f_u_arrmul24_fa5_19_f_u_arrmul24_fa4_19_y4;
  assign f_u_arrmul24_fa5_19_y4 = f_u_arrmul24_fa5_19_y1 | f_u_arrmul24_fa5_19_y3;
  assign f_u_arrmul24_and6_19_a_6 = a_6;
  assign f_u_arrmul24_and6_19_b_19 = b_19;
  assign f_u_arrmul24_and6_19_y0 = f_u_arrmul24_and6_19_a_6 & f_u_arrmul24_and6_19_b_19;
  assign f_u_arrmul24_fa6_19_f_u_arrmul24_and6_19_y0 = f_u_arrmul24_and6_19_y0;
  assign f_u_arrmul24_fa6_19_f_u_arrmul24_fa7_18_y2 = f_u_arrmul24_fa7_18_y2;
  assign f_u_arrmul24_fa6_19_f_u_arrmul24_fa5_19_y4 = f_u_arrmul24_fa5_19_y4;
  assign f_u_arrmul24_fa6_19_y0 = f_u_arrmul24_fa6_19_f_u_arrmul24_and6_19_y0 ^ f_u_arrmul24_fa6_19_f_u_arrmul24_fa7_18_y2;
  assign f_u_arrmul24_fa6_19_y1 = f_u_arrmul24_fa6_19_f_u_arrmul24_and6_19_y0 & f_u_arrmul24_fa6_19_f_u_arrmul24_fa7_18_y2;
  assign f_u_arrmul24_fa6_19_y2 = f_u_arrmul24_fa6_19_y0 ^ f_u_arrmul24_fa6_19_f_u_arrmul24_fa5_19_y4;
  assign f_u_arrmul24_fa6_19_y3 = f_u_arrmul24_fa6_19_y0 & f_u_arrmul24_fa6_19_f_u_arrmul24_fa5_19_y4;
  assign f_u_arrmul24_fa6_19_y4 = f_u_arrmul24_fa6_19_y1 | f_u_arrmul24_fa6_19_y3;
  assign f_u_arrmul24_and7_19_a_7 = a_7;
  assign f_u_arrmul24_and7_19_b_19 = b_19;
  assign f_u_arrmul24_and7_19_y0 = f_u_arrmul24_and7_19_a_7 & f_u_arrmul24_and7_19_b_19;
  assign f_u_arrmul24_fa7_19_f_u_arrmul24_and7_19_y0 = f_u_arrmul24_and7_19_y0;
  assign f_u_arrmul24_fa7_19_f_u_arrmul24_fa8_18_y2 = f_u_arrmul24_fa8_18_y2;
  assign f_u_arrmul24_fa7_19_f_u_arrmul24_fa6_19_y4 = f_u_arrmul24_fa6_19_y4;
  assign f_u_arrmul24_fa7_19_y0 = f_u_arrmul24_fa7_19_f_u_arrmul24_and7_19_y0 ^ f_u_arrmul24_fa7_19_f_u_arrmul24_fa8_18_y2;
  assign f_u_arrmul24_fa7_19_y1 = f_u_arrmul24_fa7_19_f_u_arrmul24_and7_19_y0 & f_u_arrmul24_fa7_19_f_u_arrmul24_fa8_18_y2;
  assign f_u_arrmul24_fa7_19_y2 = f_u_arrmul24_fa7_19_y0 ^ f_u_arrmul24_fa7_19_f_u_arrmul24_fa6_19_y4;
  assign f_u_arrmul24_fa7_19_y3 = f_u_arrmul24_fa7_19_y0 & f_u_arrmul24_fa7_19_f_u_arrmul24_fa6_19_y4;
  assign f_u_arrmul24_fa7_19_y4 = f_u_arrmul24_fa7_19_y1 | f_u_arrmul24_fa7_19_y3;
  assign f_u_arrmul24_and8_19_a_8 = a_8;
  assign f_u_arrmul24_and8_19_b_19 = b_19;
  assign f_u_arrmul24_and8_19_y0 = f_u_arrmul24_and8_19_a_8 & f_u_arrmul24_and8_19_b_19;
  assign f_u_arrmul24_fa8_19_f_u_arrmul24_and8_19_y0 = f_u_arrmul24_and8_19_y0;
  assign f_u_arrmul24_fa8_19_f_u_arrmul24_fa9_18_y2 = f_u_arrmul24_fa9_18_y2;
  assign f_u_arrmul24_fa8_19_f_u_arrmul24_fa7_19_y4 = f_u_arrmul24_fa7_19_y4;
  assign f_u_arrmul24_fa8_19_y0 = f_u_arrmul24_fa8_19_f_u_arrmul24_and8_19_y0 ^ f_u_arrmul24_fa8_19_f_u_arrmul24_fa9_18_y2;
  assign f_u_arrmul24_fa8_19_y1 = f_u_arrmul24_fa8_19_f_u_arrmul24_and8_19_y0 & f_u_arrmul24_fa8_19_f_u_arrmul24_fa9_18_y2;
  assign f_u_arrmul24_fa8_19_y2 = f_u_arrmul24_fa8_19_y0 ^ f_u_arrmul24_fa8_19_f_u_arrmul24_fa7_19_y4;
  assign f_u_arrmul24_fa8_19_y3 = f_u_arrmul24_fa8_19_y0 & f_u_arrmul24_fa8_19_f_u_arrmul24_fa7_19_y4;
  assign f_u_arrmul24_fa8_19_y4 = f_u_arrmul24_fa8_19_y1 | f_u_arrmul24_fa8_19_y3;
  assign f_u_arrmul24_and9_19_a_9 = a_9;
  assign f_u_arrmul24_and9_19_b_19 = b_19;
  assign f_u_arrmul24_and9_19_y0 = f_u_arrmul24_and9_19_a_9 & f_u_arrmul24_and9_19_b_19;
  assign f_u_arrmul24_fa9_19_f_u_arrmul24_and9_19_y0 = f_u_arrmul24_and9_19_y0;
  assign f_u_arrmul24_fa9_19_f_u_arrmul24_fa10_18_y2 = f_u_arrmul24_fa10_18_y2;
  assign f_u_arrmul24_fa9_19_f_u_arrmul24_fa8_19_y4 = f_u_arrmul24_fa8_19_y4;
  assign f_u_arrmul24_fa9_19_y0 = f_u_arrmul24_fa9_19_f_u_arrmul24_and9_19_y0 ^ f_u_arrmul24_fa9_19_f_u_arrmul24_fa10_18_y2;
  assign f_u_arrmul24_fa9_19_y1 = f_u_arrmul24_fa9_19_f_u_arrmul24_and9_19_y0 & f_u_arrmul24_fa9_19_f_u_arrmul24_fa10_18_y2;
  assign f_u_arrmul24_fa9_19_y2 = f_u_arrmul24_fa9_19_y0 ^ f_u_arrmul24_fa9_19_f_u_arrmul24_fa8_19_y4;
  assign f_u_arrmul24_fa9_19_y3 = f_u_arrmul24_fa9_19_y0 & f_u_arrmul24_fa9_19_f_u_arrmul24_fa8_19_y4;
  assign f_u_arrmul24_fa9_19_y4 = f_u_arrmul24_fa9_19_y1 | f_u_arrmul24_fa9_19_y3;
  assign f_u_arrmul24_and10_19_a_10 = a_10;
  assign f_u_arrmul24_and10_19_b_19 = b_19;
  assign f_u_arrmul24_and10_19_y0 = f_u_arrmul24_and10_19_a_10 & f_u_arrmul24_and10_19_b_19;
  assign f_u_arrmul24_fa10_19_f_u_arrmul24_and10_19_y0 = f_u_arrmul24_and10_19_y0;
  assign f_u_arrmul24_fa10_19_f_u_arrmul24_fa11_18_y2 = f_u_arrmul24_fa11_18_y2;
  assign f_u_arrmul24_fa10_19_f_u_arrmul24_fa9_19_y4 = f_u_arrmul24_fa9_19_y4;
  assign f_u_arrmul24_fa10_19_y0 = f_u_arrmul24_fa10_19_f_u_arrmul24_and10_19_y0 ^ f_u_arrmul24_fa10_19_f_u_arrmul24_fa11_18_y2;
  assign f_u_arrmul24_fa10_19_y1 = f_u_arrmul24_fa10_19_f_u_arrmul24_and10_19_y0 & f_u_arrmul24_fa10_19_f_u_arrmul24_fa11_18_y2;
  assign f_u_arrmul24_fa10_19_y2 = f_u_arrmul24_fa10_19_y0 ^ f_u_arrmul24_fa10_19_f_u_arrmul24_fa9_19_y4;
  assign f_u_arrmul24_fa10_19_y3 = f_u_arrmul24_fa10_19_y0 & f_u_arrmul24_fa10_19_f_u_arrmul24_fa9_19_y4;
  assign f_u_arrmul24_fa10_19_y4 = f_u_arrmul24_fa10_19_y1 | f_u_arrmul24_fa10_19_y3;
  assign f_u_arrmul24_and11_19_a_11 = a_11;
  assign f_u_arrmul24_and11_19_b_19 = b_19;
  assign f_u_arrmul24_and11_19_y0 = f_u_arrmul24_and11_19_a_11 & f_u_arrmul24_and11_19_b_19;
  assign f_u_arrmul24_fa11_19_f_u_arrmul24_and11_19_y0 = f_u_arrmul24_and11_19_y0;
  assign f_u_arrmul24_fa11_19_f_u_arrmul24_fa12_18_y2 = f_u_arrmul24_fa12_18_y2;
  assign f_u_arrmul24_fa11_19_f_u_arrmul24_fa10_19_y4 = f_u_arrmul24_fa10_19_y4;
  assign f_u_arrmul24_fa11_19_y0 = f_u_arrmul24_fa11_19_f_u_arrmul24_and11_19_y0 ^ f_u_arrmul24_fa11_19_f_u_arrmul24_fa12_18_y2;
  assign f_u_arrmul24_fa11_19_y1 = f_u_arrmul24_fa11_19_f_u_arrmul24_and11_19_y0 & f_u_arrmul24_fa11_19_f_u_arrmul24_fa12_18_y2;
  assign f_u_arrmul24_fa11_19_y2 = f_u_arrmul24_fa11_19_y0 ^ f_u_arrmul24_fa11_19_f_u_arrmul24_fa10_19_y4;
  assign f_u_arrmul24_fa11_19_y3 = f_u_arrmul24_fa11_19_y0 & f_u_arrmul24_fa11_19_f_u_arrmul24_fa10_19_y4;
  assign f_u_arrmul24_fa11_19_y4 = f_u_arrmul24_fa11_19_y1 | f_u_arrmul24_fa11_19_y3;
  assign f_u_arrmul24_and12_19_a_12 = a_12;
  assign f_u_arrmul24_and12_19_b_19 = b_19;
  assign f_u_arrmul24_and12_19_y0 = f_u_arrmul24_and12_19_a_12 & f_u_arrmul24_and12_19_b_19;
  assign f_u_arrmul24_fa12_19_f_u_arrmul24_and12_19_y0 = f_u_arrmul24_and12_19_y0;
  assign f_u_arrmul24_fa12_19_f_u_arrmul24_fa13_18_y2 = f_u_arrmul24_fa13_18_y2;
  assign f_u_arrmul24_fa12_19_f_u_arrmul24_fa11_19_y4 = f_u_arrmul24_fa11_19_y4;
  assign f_u_arrmul24_fa12_19_y0 = f_u_arrmul24_fa12_19_f_u_arrmul24_and12_19_y0 ^ f_u_arrmul24_fa12_19_f_u_arrmul24_fa13_18_y2;
  assign f_u_arrmul24_fa12_19_y1 = f_u_arrmul24_fa12_19_f_u_arrmul24_and12_19_y0 & f_u_arrmul24_fa12_19_f_u_arrmul24_fa13_18_y2;
  assign f_u_arrmul24_fa12_19_y2 = f_u_arrmul24_fa12_19_y0 ^ f_u_arrmul24_fa12_19_f_u_arrmul24_fa11_19_y4;
  assign f_u_arrmul24_fa12_19_y3 = f_u_arrmul24_fa12_19_y0 & f_u_arrmul24_fa12_19_f_u_arrmul24_fa11_19_y4;
  assign f_u_arrmul24_fa12_19_y4 = f_u_arrmul24_fa12_19_y1 | f_u_arrmul24_fa12_19_y3;
  assign f_u_arrmul24_and13_19_a_13 = a_13;
  assign f_u_arrmul24_and13_19_b_19 = b_19;
  assign f_u_arrmul24_and13_19_y0 = f_u_arrmul24_and13_19_a_13 & f_u_arrmul24_and13_19_b_19;
  assign f_u_arrmul24_fa13_19_f_u_arrmul24_and13_19_y0 = f_u_arrmul24_and13_19_y0;
  assign f_u_arrmul24_fa13_19_f_u_arrmul24_fa14_18_y2 = f_u_arrmul24_fa14_18_y2;
  assign f_u_arrmul24_fa13_19_f_u_arrmul24_fa12_19_y4 = f_u_arrmul24_fa12_19_y4;
  assign f_u_arrmul24_fa13_19_y0 = f_u_arrmul24_fa13_19_f_u_arrmul24_and13_19_y0 ^ f_u_arrmul24_fa13_19_f_u_arrmul24_fa14_18_y2;
  assign f_u_arrmul24_fa13_19_y1 = f_u_arrmul24_fa13_19_f_u_arrmul24_and13_19_y0 & f_u_arrmul24_fa13_19_f_u_arrmul24_fa14_18_y2;
  assign f_u_arrmul24_fa13_19_y2 = f_u_arrmul24_fa13_19_y0 ^ f_u_arrmul24_fa13_19_f_u_arrmul24_fa12_19_y4;
  assign f_u_arrmul24_fa13_19_y3 = f_u_arrmul24_fa13_19_y0 & f_u_arrmul24_fa13_19_f_u_arrmul24_fa12_19_y4;
  assign f_u_arrmul24_fa13_19_y4 = f_u_arrmul24_fa13_19_y1 | f_u_arrmul24_fa13_19_y3;
  assign f_u_arrmul24_and14_19_a_14 = a_14;
  assign f_u_arrmul24_and14_19_b_19 = b_19;
  assign f_u_arrmul24_and14_19_y0 = f_u_arrmul24_and14_19_a_14 & f_u_arrmul24_and14_19_b_19;
  assign f_u_arrmul24_fa14_19_f_u_arrmul24_and14_19_y0 = f_u_arrmul24_and14_19_y0;
  assign f_u_arrmul24_fa14_19_f_u_arrmul24_fa15_18_y2 = f_u_arrmul24_fa15_18_y2;
  assign f_u_arrmul24_fa14_19_f_u_arrmul24_fa13_19_y4 = f_u_arrmul24_fa13_19_y4;
  assign f_u_arrmul24_fa14_19_y0 = f_u_arrmul24_fa14_19_f_u_arrmul24_and14_19_y0 ^ f_u_arrmul24_fa14_19_f_u_arrmul24_fa15_18_y2;
  assign f_u_arrmul24_fa14_19_y1 = f_u_arrmul24_fa14_19_f_u_arrmul24_and14_19_y0 & f_u_arrmul24_fa14_19_f_u_arrmul24_fa15_18_y2;
  assign f_u_arrmul24_fa14_19_y2 = f_u_arrmul24_fa14_19_y0 ^ f_u_arrmul24_fa14_19_f_u_arrmul24_fa13_19_y4;
  assign f_u_arrmul24_fa14_19_y3 = f_u_arrmul24_fa14_19_y0 & f_u_arrmul24_fa14_19_f_u_arrmul24_fa13_19_y4;
  assign f_u_arrmul24_fa14_19_y4 = f_u_arrmul24_fa14_19_y1 | f_u_arrmul24_fa14_19_y3;
  assign f_u_arrmul24_and15_19_a_15 = a_15;
  assign f_u_arrmul24_and15_19_b_19 = b_19;
  assign f_u_arrmul24_and15_19_y0 = f_u_arrmul24_and15_19_a_15 & f_u_arrmul24_and15_19_b_19;
  assign f_u_arrmul24_fa15_19_f_u_arrmul24_and15_19_y0 = f_u_arrmul24_and15_19_y0;
  assign f_u_arrmul24_fa15_19_f_u_arrmul24_fa16_18_y2 = f_u_arrmul24_fa16_18_y2;
  assign f_u_arrmul24_fa15_19_f_u_arrmul24_fa14_19_y4 = f_u_arrmul24_fa14_19_y4;
  assign f_u_arrmul24_fa15_19_y0 = f_u_arrmul24_fa15_19_f_u_arrmul24_and15_19_y0 ^ f_u_arrmul24_fa15_19_f_u_arrmul24_fa16_18_y2;
  assign f_u_arrmul24_fa15_19_y1 = f_u_arrmul24_fa15_19_f_u_arrmul24_and15_19_y0 & f_u_arrmul24_fa15_19_f_u_arrmul24_fa16_18_y2;
  assign f_u_arrmul24_fa15_19_y2 = f_u_arrmul24_fa15_19_y0 ^ f_u_arrmul24_fa15_19_f_u_arrmul24_fa14_19_y4;
  assign f_u_arrmul24_fa15_19_y3 = f_u_arrmul24_fa15_19_y0 & f_u_arrmul24_fa15_19_f_u_arrmul24_fa14_19_y4;
  assign f_u_arrmul24_fa15_19_y4 = f_u_arrmul24_fa15_19_y1 | f_u_arrmul24_fa15_19_y3;
  assign f_u_arrmul24_and16_19_a_16 = a_16;
  assign f_u_arrmul24_and16_19_b_19 = b_19;
  assign f_u_arrmul24_and16_19_y0 = f_u_arrmul24_and16_19_a_16 & f_u_arrmul24_and16_19_b_19;
  assign f_u_arrmul24_fa16_19_f_u_arrmul24_and16_19_y0 = f_u_arrmul24_and16_19_y0;
  assign f_u_arrmul24_fa16_19_f_u_arrmul24_fa17_18_y2 = f_u_arrmul24_fa17_18_y2;
  assign f_u_arrmul24_fa16_19_f_u_arrmul24_fa15_19_y4 = f_u_arrmul24_fa15_19_y4;
  assign f_u_arrmul24_fa16_19_y0 = f_u_arrmul24_fa16_19_f_u_arrmul24_and16_19_y0 ^ f_u_arrmul24_fa16_19_f_u_arrmul24_fa17_18_y2;
  assign f_u_arrmul24_fa16_19_y1 = f_u_arrmul24_fa16_19_f_u_arrmul24_and16_19_y0 & f_u_arrmul24_fa16_19_f_u_arrmul24_fa17_18_y2;
  assign f_u_arrmul24_fa16_19_y2 = f_u_arrmul24_fa16_19_y0 ^ f_u_arrmul24_fa16_19_f_u_arrmul24_fa15_19_y4;
  assign f_u_arrmul24_fa16_19_y3 = f_u_arrmul24_fa16_19_y0 & f_u_arrmul24_fa16_19_f_u_arrmul24_fa15_19_y4;
  assign f_u_arrmul24_fa16_19_y4 = f_u_arrmul24_fa16_19_y1 | f_u_arrmul24_fa16_19_y3;
  assign f_u_arrmul24_and17_19_a_17 = a_17;
  assign f_u_arrmul24_and17_19_b_19 = b_19;
  assign f_u_arrmul24_and17_19_y0 = f_u_arrmul24_and17_19_a_17 & f_u_arrmul24_and17_19_b_19;
  assign f_u_arrmul24_fa17_19_f_u_arrmul24_and17_19_y0 = f_u_arrmul24_and17_19_y0;
  assign f_u_arrmul24_fa17_19_f_u_arrmul24_fa18_18_y2 = f_u_arrmul24_fa18_18_y2;
  assign f_u_arrmul24_fa17_19_f_u_arrmul24_fa16_19_y4 = f_u_arrmul24_fa16_19_y4;
  assign f_u_arrmul24_fa17_19_y0 = f_u_arrmul24_fa17_19_f_u_arrmul24_and17_19_y0 ^ f_u_arrmul24_fa17_19_f_u_arrmul24_fa18_18_y2;
  assign f_u_arrmul24_fa17_19_y1 = f_u_arrmul24_fa17_19_f_u_arrmul24_and17_19_y0 & f_u_arrmul24_fa17_19_f_u_arrmul24_fa18_18_y2;
  assign f_u_arrmul24_fa17_19_y2 = f_u_arrmul24_fa17_19_y0 ^ f_u_arrmul24_fa17_19_f_u_arrmul24_fa16_19_y4;
  assign f_u_arrmul24_fa17_19_y3 = f_u_arrmul24_fa17_19_y0 & f_u_arrmul24_fa17_19_f_u_arrmul24_fa16_19_y4;
  assign f_u_arrmul24_fa17_19_y4 = f_u_arrmul24_fa17_19_y1 | f_u_arrmul24_fa17_19_y3;
  assign f_u_arrmul24_and18_19_a_18 = a_18;
  assign f_u_arrmul24_and18_19_b_19 = b_19;
  assign f_u_arrmul24_and18_19_y0 = f_u_arrmul24_and18_19_a_18 & f_u_arrmul24_and18_19_b_19;
  assign f_u_arrmul24_fa18_19_f_u_arrmul24_and18_19_y0 = f_u_arrmul24_and18_19_y0;
  assign f_u_arrmul24_fa18_19_f_u_arrmul24_fa19_18_y2 = f_u_arrmul24_fa19_18_y2;
  assign f_u_arrmul24_fa18_19_f_u_arrmul24_fa17_19_y4 = f_u_arrmul24_fa17_19_y4;
  assign f_u_arrmul24_fa18_19_y0 = f_u_arrmul24_fa18_19_f_u_arrmul24_and18_19_y0 ^ f_u_arrmul24_fa18_19_f_u_arrmul24_fa19_18_y2;
  assign f_u_arrmul24_fa18_19_y1 = f_u_arrmul24_fa18_19_f_u_arrmul24_and18_19_y0 & f_u_arrmul24_fa18_19_f_u_arrmul24_fa19_18_y2;
  assign f_u_arrmul24_fa18_19_y2 = f_u_arrmul24_fa18_19_y0 ^ f_u_arrmul24_fa18_19_f_u_arrmul24_fa17_19_y4;
  assign f_u_arrmul24_fa18_19_y3 = f_u_arrmul24_fa18_19_y0 & f_u_arrmul24_fa18_19_f_u_arrmul24_fa17_19_y4;
  assign f_u_arrmul24_fa18_19_y4 = f_u_arrmul24_fa18_19_y1 | f_u_arrmul24_fa18_19_y3;
  assign f_u_arrmul24_and19_19_a_19 = a_19;
  assign f_u_arrmul24_and19_19_b_19 = b_19;
  assign f_u_arrmul24_and19_19_y0 = f_u_arrmul24_and19_19_a_19 & f_u_arrmul24_and19_19_b_19;
  assign f_u_arrmul24_fa19_19_f_u_arrmul24_and19_19_y0 = f_u_arrmul24_and19_19_y0;
  assign f_u_arrmul24_fa19_19_f_u_arrmul24_fa20_18_y2 = f_u_arrmul24_fa20_18_y2;
  assign f_u_arrmul24_fa19_19_f_u_arrmul24_fa18_19_y4 = f_u_arrmul24_fa18_19_y4;
  assign f_u_arrmul24_fa19_19_y0 = f_u_arrmul24_fa19_19_f_u_arrmul24_and19_19_y0 ^ f_u_arrmul24_fa19_19_f_u_arrmul24_fa20_18_y2;
  assign f_u_arrmul24_fa19_19_y1 = f_u_arrmul24_fa19_19_f_u_arrmul24_and19_19_y0 & f_u_arrmul24_fa19_19_f_u_arrmul24_fa20_18_y2;
  assign f_u_arrmul24_fa19_19_y2 = f_u_arrmul24_fa19_19_y0 ^ f_u_arrmul24_fa19_19_f_u_arrmul24_fa18_19_y4;
  assign f_u_arrmul24_fa19_19_y3 = f_u_arrmul24_fa19_19_y0 & f_u_arrmul24_fa19_19_f_u_arrmul24_fa18_19_y4;
  assign f_u_arrmul24_fa19_19_y4 = f_u_arrmul24_fa19_19_y1 | f_u_arrmul24_fa19_19_y3;
  assign f_u_arrmul24_and20_19_a_20 = a_20;
  assign f_u_arrmul24_and20_19_b_19 = b_19;
  assign f_u_arrmul24_and20_19_y0 = f_u_arrmul24_and20_19_a_20 & f_u_arrmul24_and20_19_b_19;
  assign f_u_arrmul24_fa20_19_f_u_arrmul24_and20_19_y0 = f_u_arrmul24_and20_19_y0;
  assign f_u_arrmul24_fa20_19_f_u_arrmul24_fa21_18_y2 = f_u_arrmul24_fa21_18_y2;
  assign f_u_arrmul24_fa20_19_f_u_arrmul24_fa19_19_y4 = f_u_arrmul24_fa19_19_y4;
  assign f_u_arrmul24_fa20_19_y0 = f_u_arrmul24_fa20_19_f_u_arrmul24_and20_19_y0 ^ f_u_arrmul24_fa20_19_f_u_arrmul24_fa21_18_y2;
  assign f_u_arrmul24_fa20_19_y1 = f_u_arrmul24_fa20_19_f_u_arrmul24_and20_19_y0 & f_u_arrmul24_fa20_19_f_u_arrmul24_fa21_18_y2;
  assign f_u_arrmul24_fa20_19_y2 = f_u_arrmul24_fa20_19_y0 ^ f_u_arrmul24_fa20_19_f_u_arrmul24_fa19_19_y4;
  assign f_u_arrmul24_fa20_19_y3 = f_u_arrmul24_fa20_19_y0 & f_u_arrmul24_fa20_19_f_u_arrmul24_fa19_19_y4;
  assign f_u_arrmul24_fa20_19_y4 = f_u_arrmul24_fa20_19_y1 | f_u_arrmul24_fa20_19_y3;
  assign f_u_arrmul24_and21_19_a_21 = a_21;
  assign f_u_arrmul24_and21_19_b_19 = b_19;
  assign f_u_arrmul24_and21_19_y0 = f_u_arrmul24_and21_19_a_21 & f_u_arrmul24_and21_19_b_19;
  assign f_u_arrmul24_fa21_19_f_u_arrmul24_and21_19_y0 = f_u_arrmul24_and21_19_y0;
  assign f_u_arrmul24_fa21_19_f_u_arrmul24_fa22_18_y2 = f_u_arrmul24_fa22_18_y2;
  assign f_u_arrmul24_fa21_19_f_u_arrmul24_fa20_19_y4 = f_u_arrmul24_fa20_19_y4;
  assign f_u_arrmul24_fa21_19_y0 = f_u_arrmul24_fa21_19_f_u_arrmul24_and21_19_y0 ^ f_u_arrmul24_fa21_19_f_u_arrmul24_fa22_18_y2;
  assign f_u_arrmul24_fa21_19_y1 = f_u_arrmul24_fa21_19_f_u_arrmul24_and21_19_y0 & f_u_arrmul24_fa21_19_f_u_arrmul24_fa22_18_y2;
  assign f_u_arrmul24_fa21_19_y2 = f_u_arrmul24_fa21_19_y0 ^ f_u_arrmul24_fa21_19_f_u_arrmul24_fa20_19_y4;
  assign f_u_arrmul24_fa21_19_y3 = f_u_arrmul24_fa21_19_y0 & f_u_arrmul24_fa21_19_f_u_arrmul24_fa20_19_y4;
  assign f_u_arrmul24_fa21_19_y4 = f_u_arrmul24_fa21_19_y1 | f_u_arrmul24_fa21_19_y3;
  assign f_u_arrmul24_and22_19_a_22 = a_22;
  assign f_u_arrmul24_and22_19_b_19 = b_19;
  assign f_u_arrmul24_and22_19_y0 = f_u_arrmul24_and22_19_a_22 & f_u_arrmul24_and22_19_b_19;
  assign f_u_arrmul24_fa22_19_f_u_arrmul24_and22_19_y0 = f_u_arrmul24_and22_19_y0;
  assign f_u_arrmul24_fa22_19_f_u_arrmul24_fa23_18_y2 = f_u_arrmul24_fa23_18_y2;
  assign f_u_arrmul24_fa22_19_f_u_arrmul24_fa21_19_y4 = f_u_arrmul24_fa21_19_y4;
  assign f_u_arrmul24_fa22_19_y0 = f_u_arrmul24_fa22_19_f_u_arrmul24_and22_19_y0 ^ f_u_arrmul24_fa22_19_f_u_arrmul24_fa23_18_y2;
  assign f_u_arrmul24_fa22_19_y1 = f_u_arrmul24_fa22_19_f_u_arrmul24_and22_19_y0 & f_u_arrmul24_fa22_19_f_u_arrmul24_fa23_18_y2;
  assign f_u_arrmul24_fa22_19_y2 = f_u_arrmul24_fa22_19_y0 ^ f_u_arrmul24_fa22_19_f_u_arrmul24_fa21_19_y4;
  assign f_u_arrmul24_fa22_19_y3 = f_u_arrmul24_fa22_19_y0 & f_u_arrmul24_fa22_19_f_u_arrmul24_fa21_19_y4;
  assign f_u_arrmul24_fa22_19_y4 = f_u_arrmul24_fa22_19_y1 | f_u_arrmul24_fa22_19_y3;
  assign f_u_arrmul24_and23_19_a_23 = a_23;
  assign f_u_arrmul24_and23_19_b_19 = b_19;
  assign f_u_arrmul24_and23_19_y0 = f_u_arrmul24_and23_19_a_23 & f_u_arrmul24_and23_19_b_19;
  assign f_u_arrmul24_fa23_19_f_u_arrmul24_and23_19_y0 = f_u_arrmul24_and23_19_y0;
  assign f_u_arrmul24_fa23_19_f_u_arrmul24_fa23_18_y4 = f_u_arrmul24_fa23_18_y4;
  assign f_u_arrmul24_fa23_19_f_u_arrmul24_fa22_19_y4 = f_u_arrmul24_fa22_19_y4;
  assign f_u_arrmul24_fa23_19_y0 = f_u_arrmul24_fa23_19_f_u_arrmul24_and23_19_y0 ^ f_u_arrmul24_fa23_19_f_u_arrmul24_fa23_18_y4;
  assign f_u_arrmul24_fa23_19_y1 = f_u_arrmul24_fa23_19_f_u_arrmul24_and23_19_y0 & f_u_arrmul24_fa23_19_f_u_arrmul24_fa23_18_y4;
  assign f_u_arrmul24_fa23_19_y2 = f_u_arrmul24_fa23_19_y0 ^ f_u_arrmul24_fa23_19_f_u_arrmul24_fa22_19_y4;
  assign f_u_arrmul24_fa23_19_y3 = f_u_arrmul24_fa23_19_y0 & f_u_arrmul24_fa23_19_f_u_arrmul24_fa22_19_y4;
  assign f_u_arrmul24_fa23_19_y4 = f_u_arrmul24_fa23_19_y1 | f_u_arrmul24_fa23_19_y3;
  assign f_u_arrmul24_and0_20_a_0 = a_0;
  assign f_u_arrmul24_and0_20_b_20 = b_20;
  assign f_u_arrmul24_and0_20_y0 = f_u_arrmul24_and0_20_a_0 & f_u_arrmul24_and0_20_b_20;
  assign f_u_arrmul24_ha0_20_f_u_arrmul24_and0_20_y0 = f_u_arrmul24_and0_20_y0;
  assign f_u_arrmul24_ha0_20_f_u_arrmul24_fa1_19_y2 = f_u_arrmul24_fa1_19_y2;
  assign f_u_arrmul24_ha0_20_y0 = f_u_arrmul24_ha0_20_f_u_arrmul24_and0_20_y0 ^ f_u_arrmul24_ha0_20_f_u_arrmul24_fa1_19_y2;
  assign f_u_arrmul24_ha0_20_y1 = f_u_arrmul24_ha0_20_f_u_arrmul24_and0_20_y0 & f_u_arrmul24_ha0_20_f_u_arrmul24_fa1_19_y2;
  assign f_u_arrmul24_and1_20_a_1 = a_1;
  assign f_u_arrmul24_and1_20_b_20 = b_20;
  assign f_u_arrmul24_and1_20_y0 = f_u_arrmul24_and1_20_a_1 & f_u_arrmul24_and1_20_b_20;
  assign f_u_arrmul24_fa1_20_f_u_arrmul24_and1_20_y0 = f_u_arrmul24_and1_20_y0;
  assign f_u_arrmul24_fa1_20_f_u_arrmul24_fa2_19_y2 = f_u_arrmul24_fa2_19_y2;
  assign f_u_arrmul24_fa1_20_f_u_arrmul24_ha0_20_y1 = f_u_arrmul24_ha0_20_y1;
  assign f_u_arrmul24_fa1_20_y0 = f_u_arrmul24_fa1_20_f_u_arrmul24_and1_20_y0 ^ f_u_arrmul24_fa1_20_f_u_arrmul24_fa2_19_y2;
  assign f_u_arrmul24_fa1_20_y1 = f_u_arrmul24_fa1_20_f_u_arrmul24_and1_20_y0 & f_u_arrmul24_fa1_20_f_u_arrmul24_fa2_19_y2;
  assign f_u_arrmul24_fa1_20_y2 = f_u_arrmul24_fa1_20_y0 ^ f_u_arrmul24_fa1_20_f_u_arrmul24_ha0_20_y1;
  assign f_u_arrmul24_fa1_20_y3 = f_u_arrmul24_fa1_20_y0 & f_u_arrmul24_fa1_20_f_u_arrmul24_ha0_20_y1;
  assign f_u_arrmul24_fa1_20_y4 = f_u_arrmul24_fa1_20_y1 | f_u_arrmul24_fa1_20_y3;
  assign f_u_arrmul24_and2_20_a_2 = a_2;
  assign f_u_arrmul24_and2_20_b_20 = b_20;
  assign f_u_arrmul24_and2_20_y0 = f_u_arrmul24_and2_20_a_2 & f_u_arrmul24_and2_20_b_20;
  assign f_u_arrmul24_fa2_20_f_u_arrmul24_and2_20_y0 = f_u_arrmul24_and2_20_y0;
  assign f_u_arrmul24_fa2_20_f_u_arrmul24_fa3_19_y2 = f_u_arrmul24_fa3_19_y2;
  assign f_u_arrmul24_fa2_20_f_u_arrmul24_fa1_20_y4 = f_u_arrmul24_fa1_20_y4;
  assign f_u_arrmul24_fa2_20_y0 = f_u_arrmul24_fa2_20_f_u_arrmul24_and2_20_y0 ^ f_u_arrmul24_fa2_20_f_u_arrmul24_fa3_19_y2;
  assign f_u_arrmul24_fa2_20_y1 = f_u_arrmul24_fa2_20_f_u_arrmul24_and2_20_y0 & f_u_arrmul24_fa2_20_f_u_arrmul24_fa3_19_y2;
  assign f_u_arrmul24_fa2_20_y2 = f_u_arrmul24_fa2_20_y0 ^ f_u_arrmul24_fa2_20_f_u_arrmul24_fa1_20_y4;
  assign f_u_arrmul24_fa2_20_y3 = f_u_arrmul24_fa2_20_y0 & f_u_arrmul24_fa2_20_f_u_arrmul24_fa1_20_y4;
  assign f_u_arrmul24_fa2_20_y4 = f_u_arrmul24_fa2_20_y1 | f_u_arrmul24_fa2_20_y3;
  assign f_u_arrmul24_and3_20_a_3 = a_3;
  assign f_u_arrmul24_and3_20_b_20 = b_20;
  assign f_u_arrmul24_and3_20_y0 = f_u_arrmul24_and3_20_a_3 & f_u_arrmul24_and3_20_b_20;
  assign f_u_arrmul24_fa3_20_f_u_arrmul24_and3_20_y0 = f_u_arrmul24_and3_20_y0;
  assign f_u_arrmul24_fa3_20_f_u_arrmul24_fa4_19_y2 = f_u_arrmul24_fa4_19_y2;
  assign f_u_arrmul24_fa3_20_f_u_arrmul24_fa2_20_y4 = f_u_arrmul24_fa2_20_y4;
  assign f_u_arrmul24_fa3_20_y0 = f_u_arrmul24_fa3_20_f_u_arrmul24_and3_20_y0 ^ f_u_arrmul24_fa3_20_f_u_arrmul24_fa4_19_y2;
  assign f_u_arrmul24_fa3_20_y1 = f_u_arrmul24_fa3_20_f_u_arrmul24_and3_20_y0 & f_u_arrmul24_fa3_20_f_u_arrmul24_fa4_19_y2;
  assign f_u_arrmul24_fa3_20_y2 = f_u_arrmul24_fa3_20_y0 ^ f_u_arrmul24_fa3_20_f_u_arrmul24_fa2_20_y4;
  assign f_u_arrmul24_fa3_20_y3 = f_u_arrmul24_fa3_20_y0 & f_u_arrmul24_fa3_20_f_u_arrmul24_fa2_20_y4;
  assign f_u_arrmul24_fa3_20_y4 = f_u_arrmul24_fa3_20_y1 | f_u_arrmul24_fa3_20_y3;
  assign f_u_arrmul24_and4_20_a_4 = a_4;
  assign f_u_arrmul24_and4_20_b_20 = b_20;
  assign f_u_arrmul24_and4_20_y0 = f_u_arrmul24_and4_20_a_4 & f_u_arrmul24_and4_20_b_20;
  assign f_u_arrmul24_fa4_20_f_u_arrmul24_and4_20_y0 = f_u_arrmul24_and4_20_y0;
  assign f_u_arrmul24_fa4_20_f_u_arrmul24_fa5_19_y2 = f_u_arrmul24_fa5_19_y2;
  assign f_u_arrmul24_fa4_20_f_u_arrmul24_fa3_20_y4 = f_u_arrmul24_fa3_20_y4;
  assign f_u_arrmul24_fa4_20_y0 = f_u_arrmul24_fa4_20_f_u_arrmul24_and4_20_y0 ^ f_u_arrmul24_fa4_20_f_u_arrmul24_fa5_19_y2;
  assign f_u_arrmul24_fa4_20_y1 = f_u_arrmul24_fa4_20_f_u_arrmul24_and4_20_y0 & f_u_arrmul24_fa4_20_f_u_arrmul24_fa5_19_y2;
  assign f_u_arrmul24_fa4_20_y2 = f_u_arrmul24_fa4_20_y0 ^ f_u_arrmul24_fa4_20_f_u_arrmul24_fa3_20_y4;
  assign f_u_arrmul24_fa4_20_y3 = f_u_arrmul24_fa4_20_y0 & f_u_arrmul24_fa4_20_f_u_arrmul24_fa3_20_y4;
  assign f_u_arrmul24_fa4_20_y4 = f_u_arrmul24_fa4_20_y1 | f_u_arrmul24_fa4_20_y3;
  assign f_u_arrmul24_and5_20_a_5 = a_5;
  assign f_u_arrmul24_and5_20_b_20 = b_20;
  assign f_u_arrmul24_and5_20_y0 = f_u_arrmul24_and5_20_a_5 & f_u_arrmul24_and5_20_b_20;
  assign f_u_arrmul24_fa5_20_f_u_arrmul24_and5_20_y0 = f_u_arrmul24_and5_20_y0;
  assign f_u_arrmul24_fa5_20_f_u_arrmul24_fa6_19_y2 = f_u_arrmul24_fa6_19_y2;
  assign f_u_arrmul24_fa5_20_f_u_arrmul24_fa4_20_y4 = f_u_arrmul24_fa4_20_y4;
  assign f_u_arrmul24_fa5_20_y0 = f_u_arrmul24_fa5_20_f_u_arrmul24_and5_20_y0 ^ f_u_arrmul24_fa5_20_f_u_arrmul24_fa6_19_y2;
  assign f_u_arrmul24_fa5_20_y1 = f_u_arrmul24_fa5_20_f_u_arrmul24_and5_20_y0 & f_u_arrmul24_fa5_20_f_u_arrmul24_fa6_19_y2;
  assign f_u_arrmul24_fa5_20_y2 = f_u_arrmul24_fa5_20_y0 ^ f_u_arrmul24_fa5_20_f_u_arrmul24_fa4_20_y4;
  assign f_u_arrmul24_fa5_20_y3 = f_u_arrmul24_fa5_20_y0 & f_u_arrmul24_fa5_20_f_u_arrmul24_fa4_20_y4;
  assign f_u_arrmul24_fa5_20_y4 = f_u_arrmul24_fa5_20_y1 | f_u_arrmul24_fa5_20_y3;
  assign f_u_arrmul24_and6_20_a_6 = a_6;
  assign f_u_arrmul24_and6_20_b_20 = b_20;
  assign f_u_arrmul24_and6_20_y0 = f_u_arrmul24_and6_20_a_6 & f_u_arrmul24_and6_20_b_20;
  assign f_u_arrmul24_fa6_20_f_u_arrmul24_and6_20_y0 = f_u_arrmul24_and6_20_y0;
  assign f_u_arrmul24_fa6_20_f_u_arrmul24_fa7_19_y2 = f_u_arrmul24_fa7_19_y2;
  assign f_u_arrmul24_fa6_20_f_u_arrmul24_fa5_20_y4 = f_u_arrmul24_fa5_20_y4;
  assign f_u_arrmul24_fa6_20_y0 = f_u_arrmul24_fa6_20_f_u_arrmul24_and6_20_y0 ^ f_u_arrmul24_fa6_20_f_u_arrmul24_fa7_19_y2;
  assign f_u_arrmul24_fa6_20_y1 = f_u_arrmul24_fa6_20_f_u_arrmul24_and6_20_y0 & f_u_arrmul24_fa6_20_f_u_arrmul24_fa7_19_y2;
  assign f_u_arrmul24_fa6_20_y2 = f_u_arrmul24_fa6_20_y0 ^ f_u_arrmul24_fa6_20_f_u_arrmul24_fa5_20_y4;
  assign f_u_arrmul24_fa6_20_y3 = f_u_arrmul24_fa6_20_y0 & f_u_arrmul24_fa6_20_f_u_arrmul24_fa5_20_y4;
  assign f_u_arrmul24_fa6_20_y4 = f_u_arrmul24_fa6_20_y1 | f_u_arrmul24_fa6_20_y3;
  assign f_u_arrmul24_and7_20_a_7 = a_7;
  assign f_u_arrmul24_and7_20_b_20 = b_20;
  assign f_u_arrmul24_and7_20_y0 = f_u_arrmul24_and7_20_a_7 & f_u_arrmul24_and7_20_b_20;
  assign f_u_arrmul24_fa7_20_f_u_arrmul24_and7_20_y0 = f_u_arrmul24_and7_20_y0;
  assign f_u_arrmul24_fa7_20_f_u_arrmul24_fa8_19_y2 = f_u_arrmul24_fa8_19_y2;
  assign f_u_arrmul24_fa7_20_f_u_arrmul24_fa6_20_y4 = f_u_arrmul24_fa6_20_y4;
  assign f_u_arrmul24_fa7_20_y0 = f_u_arrmul24_fa7_20_f_u_arrmul24_and7_20_y0 ^ f_u_arrmul24_fa7_20_f_u_arrmul24_fa8_19_y2;
  assign f_u_arrmul24_fa7_20_y1 = f_u_arrmul24_fa7_20_f_u_arrmul24_and7_20_y0 & f_u_arrmul24_fa7_20_f_u_arrmul24_fa8_19_y2;
  assign f_u_arrmul24_fa7_20_y2 = f_u_arrmul24_fa7_20_y0 ^ f_u_arrmul24_fa7_20_f_u_arrmul24_fa6_20_y4;
  assign f_u_arrmul24_fa7_20_y3 = f_u_arrmul24_fa7_20_y0 & f_u_arrmul24_fa7_20_f_u_arrmul24_fa6_20_y4;
  assign f_u_arrmul24_fa7_20_y4 = f_u_arrmul24_fa7_20_y1 | f_u_arrmul24_fa7_20_y3;
  assign f_u_arrmul24_and8_20_a_8 = a_8;
  assign f_u_arrmul24_and8_20_b_20 = b_20;
  assign f_u_arrmul24_and8_20_y0 = f_u_arrmul24_and8_20_a_8 & f_u_arrmul24_and8_20_b_20;
  assign f_u_arrmul24_fa8_20_f_u_arrmul24_and8_20_y0 = f_u_arrmul24_and8_20_y0;
  assign f_u_arrmul24_fa8_20_f_u_arrmul24_fa9_19_y2 = f_u_arrmul24_fa9_19_y2;
  assign f_u_arrmul24_fa8_20_f_u_arrmul24_fa7_20_y4 = f_u_arrmul24_fa7_20_y4;
  assign f_u_arrmul24_fa8_20_y0 = f_u_arrmul24_fa8_20_f_u_arrmul24_and8_20_y0 ^ f_u_arrmul24_fa8_20_f_u_arrmul24_fa9_19_y2;
  assign f_u_arrmul24_fa8_20_y1 = f_u_arrmul24_fa8_20_f_u_arrmul24_and8_20_y0 & f_u_arrmul24_fa8_20_f_u_arrmul24_fa9_19_y2;
  assign f_u_arrmul24_fa8_20_y2 = f_u_arrmul24_fa8_20_y0 ^ f_u_arrmul24_fa8_20_f_u_arrmul24_fa7_20_y4;
  assign f_u_arrmul24_fa8_20_y3 = f_u_arrmul24_fa8_20_y0 & f_u_arrmul24_fa8_20_f_u_arrmul24_fa7_20_y4;
  assign f_u_arrmul24_fa8_20_y4 = f_u_arrmul24_fa8_20_y1 | f_u_arrmul24_fa8_20_y3;
  assign f_u_arrmul24_and9_20_a_9 = a_9;
  assign f_u_arrmul24_and9_20_b_20 = b_20;
  assign f_u_arrmul24_and9_20_y0 = f_u_arrmul24_and9_20_a_9 & f_u_arrmul24_and9_20_b_20;
  assign f_u_arrmul24_fa9_20_f_u_arrmul24_and9_20_y0 = f_u_arrmul24_and9_20_y0;
  assign f_u_arrmul24_fa9_20_f_u_arrmul24_fa10_19_y2 = f_u_arrmul24_fa10_19_y2;
  assign f_u_arrmul24_fa9_20_f_u_arrmul24_fa8_20_y4 = f_u_arrmul24_fa8_20_y4;
  assign f_u_arrmul24_fa9_20_y0 = f_u_arrmul24_fa9_20_f_u_arrmul24_and9_20_y0 ^ f_u_arrmul24_fa9_20_f_u_arrmul24_fa10_19_y2;
  assign f_u_arrmul24_fa9_20_y1 = f_u_arrmul24_fa9_20_f_u_arrmul24_and9_20_y0 & f_u_arrmul24_fa9_20_f_u_arrmul24_fa10_19_y2;
  assign f_u_arrmul24_fa9_20_y2 = f_u_arrmul24_fa9_20_y0 ^ f_u_arrmul24_fa9_20_f_u_arrmul24_fa8_20_y4;
  assign f_u_arrmul24_fa9_20_y3 = f_u_arrmul24_fa9_20_y0 & f_u_arrmul24_fa9_20_f_u_arrmul24_fa8_20_y4;
  assign f_u_arrmul24_fa9_20_y4 = f_u_arrmul24_fa9_20_y1 | f_u_arrmul24_fa9_20_y3;
  assign f_u_arrmul24_and10_20_a_10 = a_10;
  assign f_u_arrmul24_and10_20_b_20 = b_20;
  assign f_u_arrmul24_and10_20_y0 = f_u_arrmul24_and10_20_a_10 & f_u_arrmul24_and10_20_b_20;
  assign f_u_arrmul24_fa10_20_f_u_arrmul24_and10_20_y0 = f_u_arrmul24_and10_20_y0;
  assign f_u_arrmul24_fa10_20_f_u_arrmul24_fa11_19_y2 = f_u_arrmul24_fa11_19_y2;
  assign f_u_arrmul24_fa10_20_f_u_arrmul24_fa9_20_y4 = f_u_arrmul24_fa9_20_y4;
  assign f_u_arrmul24_fa10_20_y0 = f_u_arrmul24_fa10_20_f_u_arrmul24_and10_20_y0 ^ f_u_arrmul24_fa10_20_f_u_arrmul24_fa11_19_y2;
  assign f_u_arrmul24_fa10_20_y1 = f_u_arrmul24_fa10_20_f_u_arrmul24_and10_20_y0 & f_u_arrmul24_fa10_20_f_u_arrmul24_fa11_19_y2;
  assign f_u_arrmul24_fa10_20_y2 = f_u_arrmul24_fa10_20_y0 ^ f_u_arrmul24_fa10_20_f_u_arrmul24_fa9_20_y4;
  assign f_u_arrmul24_fa10_20_y3 = f_u_arrmul24_fa10_20_y0 & f_u_arrmul24_fa10_20_f_u_arrmul24_fa9_20_y4;
  assign f_u_arrmul24_fa10_20_y4 = f_u_arrmul24_fa10_20_y1 | f_u_arrmul24_fa10_20_y3;
  assign f_u_arrmul24_and11_20_a_11 = a_11;
  assign f_u_arrmul24_and11_20_b_20 = b_20;
  assign f_u_arrmul24_and11_20_y0 = f_u_arrmul24_and11_20_a_11 & f_u_arrmul24_and11_20_b_20;
  assign f_u_arrmul24_fa11_20_f_u_arrmul24_and11_20_y0 = f_u_arrmul24_and11_20_y0;
  assign f_u_arrmul24_fa11_20_f_u_arrmul24_fa12_19_y2 = f_u_arrmul24_fa12_19_y2;
  assign f_u_arrmul24_fa11_20_f_u_arrmul24_fa10_20_y4 = f_u_arrmul24_fa10_20_y4;
  assign f_u_arrmul24_fa11_20_y0 = f_u_arrmul24_fa11_20_f_u_arrmul24_and11_20_y0 ^ f_u_arrmul24_fa11_20_f_u_arrmul24_fa12_19_y2;
  assign f_u_arrmul24_fa11_20_y1 = f_u_arrmul24_fa11_20_f_u_arrmul24_and11_20_y0 & f_u_arrmul24_fa11_20_f_u_arrmul24_fa12_19_y2;
  assign f_u_arrmul24_fa11_20_y2 = f_u_arrmul24_fa11_20_y0 ^ f_u_arrmul24_fa11_20_f_u_arrmul24_fa10_20_y4;
  assign f_u_arrmul24_fa11_20_y3 = f_u_arrmul24_fa11_20_y0 & f_u_arrmul24_fa11_20_f_u_arrmul24_fa10_20_y4;
  assign f_u_arrmul24_fa11_20_y4 = f_u_arrmul24_fa11_20_y1 | f_u_arrmul24_fa11_20_y3;
  assign f_u_arrmul24_and12_20_a_12 = a_12;
  assign f_u_arrmul24_and12_20_b_20 = b_20;
  assign f_u_arrmul24_and12_20_y0 = f_u_arrmul24_and12_20_a_12 & f_u_arrmul24_and12_20_b_20;
  assign f_u_arrmul24_fa12_20_f_u_arrmul24_and12_20_y0 = f_u_arrmul24_and12_20_y0;
  assign f_u_arrmul24_fa12_20_f_u_arrmul24_fa13_19_y2 = f_u_arrmul24_fa13_19_y2;
  assign f_u_arrmul24_fa12_20_f_u_arrmul24_fa11_20_y4 = f_u_arrmul24_fa11_20_y4;
  assign f_u_arrmul24_fa12_20_y0 = f_u_arrmul24_fa12_20_f_u_arrmul24_and12_20_y0 ^ f_u_arrmul24_fa12_20_f_u_arrmul24_fa13_19_y2;
  assign f_u_arrmul24_fa12_20_y1 = f_u_arrmul24_fa12_20_f_u_arrmul24_and12_20_y0 & f_u_arrmul24_fa12_20_f_u_arrmul24_fa13_19_y2;
  assign f_u_arrmul24_fa12_20_y2 = f_u_arrmul24_fa12_20_y0 ^ f_u_arrmul24_fa12_20_f_u_arrmul24_fa11_20_y4;
  assign f_u_arrmul24_fa12_20_y3 = f_u_arrmul24_fa12_20_y0 & f_u_arrmul24_fa12_20_f_u_arrmul24_fa11_20_y4;
  assign f_u_arrmul24_fa12_20_y4 = f_u_arrmul24_fa12_20_y1 | f_u_arrmul24_fa12_20_y3;
  assign f_u_arrmul24_and13_20_a_13 = a_13;
  assign f_u_arrmul24_and13_20_b_20 = b_20;
  assign f_u_arrmul24_and13_20_y0 = f_u_arrmul24_and13_20_a_13 & f_u_arrmul24_and13_20_b_20;
  assign f_u_arrmul24_fa13_20_f_u_arrmul24_and13_20_y0 = f_u_arrmul24_and13_20_y0;
  assign f_u_arrmul24_fa13_20_f_u_arrmul24_fa14_19_y2 = f_u_arrmul24_fa14_19_y2;
  assign f_u_arrmul24_fa13_20_f_u_arrmul24_fa12_20_y4 = f_u_arrmul24_fa12_20_y4;
  assign f_u_arrmul24_fa13_20_y0 = f_u_arrmul24_fa13_20_f_u_arrmul24_and13_20_y0 ^ f_u_arrmul24_fa13_20_f_u_arrmul24_fa14_19_y2;
  assign f_u_arrmul24_fa13_20_y1 = f_u_arrmul24_fa13_20_f_u_arrmul24_and13_20_y0 & f_u_arrmul24_fa13_20_f_u_arrmul24_fa14_19_y2;
  assign f_u_arrmul24_fa13_20_y2 = f_u_arrmul24_fa13_20_y0 ^ f_u_arrmul24_fa13_20_f_u_arrmul24_fa12_20_y4;
  assign f_u_arrmul24_fa13_20_y3 = f_u_arrmul24_fa13_20_y0 & f_u_arrmul24_fa13_20_f_u_arrmul24_fa12_20_y4;
  assign f_u_arrmul24_fa13_20_y4 = f_u_arrmul24_fa13_20_y1 | f_u_arrmul24_fa13_20_y3;
  assign f_u_arrmul24_and14_20_a_14 = a_14;
  assign f_u_arrmul24_and14_20_b_20 = b_20;
  assign f_u_arrmul24_and14_20_y0 = f_u_arrmul24_and14_20_a_14 & f_u_arrmul24_and14_20_b_20;
  assign f_u_arrmul24_fa14_20_f_u_arrmul24_and14_20_y0 = f_u_arrmul24_and14_20_y0;
  assign f_u_arrmul24_fa14_20_f_u_arrmul24_fa15_19_y2 = f_u_arrmul24_fa15_19_y2;
  assign f_u_arrmul24_fa14_20_f_u_arrmul24_fa13_20_y4 = f_u_arrmul24_fa13_20_y4;
  assign f_u_arrmul24_fa14_20_y0 = f_u_arrmul24_fa14_20_f_u_arrmul24_and14_20_y0 ^ f_u_arrmul24_fa14_20_f_u_arrmul24_fa15_19_y2;
  assign f_u_arrmul24_fa14_20_y1 = f_u_arrmul24_fa14_20_f_u_arrmul24_and14_20_y0 & f_u_arrmul24_fa14_20_f_u_arrmul24_fa15_19_y2;
  assign f_u_arrmul24_fa14_20_y2 = f_u_arrmul24_fa14_20_y0 ^ f_u_arrmul24_fa14_20_f_u_arrmul24_fa13_20_y4;
  assign f_u_arrmul24_fa14_20_y3 = f_u_arrmul24_fa14_20_y0 & f_u_arrmul24_fa14_20_f_u_arrmul24_fa13_20_y4;
  assign f_u_arrmul24_fa14_20_y4 = f_u_arrmul24_fa14_20_y1 | f_u_arrmul24_fa14_20_y3;
  assign f_u_arrmul24_and15_20_a_15 = a_15;
  assign f_u_arrmul24_and15_20_b_20 = b_20;
  assign f_u_arrmul24_and15_20_y0 = f_u_arrmul24_and15_20_a_15 & f_u_arrmul24_and15_20_b_20;
  assign f_u_arrmul24_fa15_20_f_u_arrmul24_and15_20_y0 = f_u_arrmul24_and15_20_y0;
  assign f_u_arrmul24_fa15_20_f_u_arrmul24_fa16_19_y2 = f_u_arrmul24_fa16_19_y2;
  assign f_u_arrmul24_fa15_20_f_u_arrmul24_fa14_20_y4 = f_u_arrmul24_fa14_20_y4;
  assign f_u_arrmul24_fa15_20_y0 = f_u_arrmul24_fa15_20_f_u_arrmul24_and15_20_y0 ^ f_u_arrmul24_fa15_20_f_u_arrmul24_fa16_19_y2;
  assign f_u_arrmul24_fa15_20_y1 = f_u_arrmul24_fa15_20_f_u_arrmul24_and15_20_y0 & f_u_arrmul24_fa15_20_f_u_arrmul24_fa16_19_y2;
  assign f_u_arrmul24_fa15_20_y2 = f_u_arrmul24_fa15_20_y0 ^ f_u_arrmul24_fa15_20_f_u_arrmul24_fa14_20_y4;
  assign f_u_arrmul24_fa15_20_y3 = f_u_arrmul24_fa15_20_y0 & f_u_arrmul24_fa15_20_f_u_arrmul24_fa14_20_y4;
  assign f_u_arrmul24_fa15_20_y4 = f_u_arrmul24_fa15_20_y1 | f_u_arrmul24_fa15_20_y3;
  assign f_u_arrmul24_and16_20_a_16 = a_16;
  assign f_u_arrmul24_and16_20_b_20 = b_20;
  assign f_u_arrmul24_and16_20_y0 = f_u_arrmul24_and16_20_a_16 & f_u_arrmul24_and16_20_b_20;
  assign f_u_arrmul24_fa16_20_f_u_arrmul24_and16_20_y0 = f_u_arrmul24_and16_20_y0;
  assign f_u_arrmul24_fa16_20_f_u_arrmul24_fa17_19_y2 = f_u_arrmul24_fa17_19_y2;
  assign f_u_arrmul24_fa16_20_f_u_arrmul24_fa15_20_y4 = f_u_arrmul24_fa15_20_y4;
  assign f_u_arrmul24_fa16_20_y0 = f_u_arrmul24_fa16_20_f_u_arrmul24_and16_20_y0 ^ f_u_arrmul24_fa16_20_f_u_arrmul24_fa17_19_y2;
  assign f_u_arrmul24_fa16_20_y1 = f_u_arrmul24_fa16_20_f_u_arrmul24_and16_20_y0 & f_u_arrmul24_fa16_20_f_u_arrmul24_fa17_19_y2;
  assign f_u_arrmul24_fa16_20_y2 = f_u_arrmul24_fa16_20_y0 ^ f_u_arrmul24_fa16_20_f_u_arrmul24_fa15_20_y4;
  assign f_u_arrmul24_fa16_20_y3 = f_u_arrmul24_fa16_20_y0 & f_u_arrmul24_fa16_20_f_u_arrmul24_fa15_20_y4;
  assign f_u_arrmul24_fa16_20_y4 = f_u_arrmul24_fa16_20_y1 | f_u_arrmul24_fa16_20_y3;
  assign f_u_arrmul24_and17_20_a_17 = a_17;
  assign f_u_arrmul24_and17_20_b_20 = b_20;
  assign f_u_arrmul24_and17_20_y0 = f_u_arrmul24_and17_20_a_17 & f_u_arrmul24_and17_20_b_20;
  assign f_u_arrmul24_fa17_20_f_u_arrmul24_and17_20_y0 = f_u_arrmul24_and17_20_y0;
  assign f_u_arrmul24_fa17_20_f_u_arrmul24_fa18_19_y2 = f_u_arrmul24_fa18_19_y2;
  assign f_u_arrmul24_fa17_20_f_u_arrmul24_fa16_20_y4 = f_u_arrmul24_fa16_20_y4;
  assign f_u_arrmul24_fa17_20_y0 = f_u_arrmul24_fa17_20_f_u_arrmul24_and17_20_y0 ^ f_u_arrmul24_fa17_20_f_u_arrmul24_fa18_19_y2;
  assign f_u_arrmul24_fa17_20_y1 = f_u_arrmul24_fa17_20_f_u_arrmul24_and17_20_y0 & f_u_arrmul24_fa17_20_f_u_arrmul24_fa18_19_y2;
  assign f_u_arrmul24_fa17_20_y2 = f_u_arrmul24_fa17_20_y0 ^ f_u_arrmul24_fa17_20_f_u_arrmul24_fa16_20_y4;
  assign f_u_arrmul24_fa17_20_y3 = f_u_arrmul24_fa17_20_y0 & f_u_arrmul24_fa17_20_f_u_arrmul24_fa16_20_y4;
  assign f_u_arrmul24_fa17_20_y4 = f_u_arrmul24_fa17_20_y1 | f_u_arrmul24_fa17_20_y3;
  assign f_u_arrmul24_and18_20_a_18 = a_18;
  assign f_u_arrmul24_and18_20_b_20 = b_20;
  assign f_u_arrmul24_and18_20_y0 = f_u_arrmul24_and18_20_a_18 & f_u_arrmul24_and18_20_b_20;
  assign f_u_arrmul24_fa18_20_f_u_arrmul24_and18_20_y0 = f_u_arrmul24_and18_20_y0;
  assign f_u_arrmul24_fa18_20_f_u_arrmul24_fa19_19_y2 = f_u_arrmul24_fa19_19_y2;
  assign f_u_arrmul24_fa18_20_f_u_arrmul24_fa17_20_y4 = f_u_arrmul24_fa17_20_y4;
  assign f_u_arrmul24_fa18_20_y0 = f_u_arrmul24_fa18_20_f_u_arrmul24_and18_20_y0 ^ f_u_arrmul24_fa18_20_f_u_arrmul24_fa19_19_y2;
  assign f_u_arrmul24_fa18_20_y1 = f_u_arrmul24_fa18_20_f_u_arrmul24_and18_20_y0 & f_u_arrmul24_fa18_20_f_u_arrmul24_fa19_19_y2;
  assign f_u_arrmul24_fa18_20_y2 = f_u_arrmul24_fa18_20_y0 ^ f_u_arrmul24_fa18_20_f_u_arrmul24_fa17_20_y4;
  assign f_u_arrmul24_fa18_20_y3 = f_u_arrmul24_fa18_20_y0 & f_u_arrmul24_fa18_20_f_u_arrmul24_fa17_20_y4;
  assign f_u_arrmul24_fa18_20_y4 = f_u_arrmul24_fa18_20_y1 | f_u_arrmul24_fa18_20_y3;
  assign f_u_arrmul24_and19_20_a_19 = a_19;
  assign f_u_arrmul24_and19_20_b_20 = b_20;
  assign f_u_arrmul24_and19_20_y0 = f_u_arrmul24_and19_20_a_19 & f_u_arrmul24_and19_20_b_20;
  assign f_u_arrmul24_fa19_20_f_u_arrmul24_and19_20_y0 = f_u_arrmul24_and19_20_y0;
  assign f_u_arrmul24_fa19_20_f_u_arrmul24_fa20_19_y2 = f_u_arrmul24_fa20_19_y2;
  assign f_u_arrmul24_fa19_20_f_u_arrmul24_fa18_20_y4 = f_u_arrmul24_fa18_20_y4;
  assign f_u_arrmul24_fa19_20_y0 = f_u_arrmul24_fa19_20_f_u_arrmul24_and19_20_y0 ^ f_u_arrmul24_fa19_20_f_u_arrmul24_fa20_19_y2;
  assign f_u_arrmul24_fa19_20_y1 = f_u_arrmul24_fa19_20_f_u_arrmul24_and19_20_y0 & f_u_arrmul24_fa19_20_f_u_arrmul24_fa20_19_y2;
  assign f_u_arrmul24_fa19_20_y2 = f_u_arrmul24_fa19_20_y0 ^ f_u_arrmul24_fa19_20_f_u_arrmul24_fa18_20_y4;
  assign f_u_arrmul24_fa19_20_y3 = f_u_arrmul24_fa19_20_y0 & f_u_arrmul24_fa19_20_f_u_arrmul24_fa18_20_y4;
  assign f_u_arrmul24_fa19_20_y4 = f_u_arrmul24_fa19_20_y1 | f_u_arrmul24_fa19_20_y3;
  assign f_u_arrmul24_and20_20_a_20 = a_20;
  assign f_u_arrmul24_and20_20_b_20 = b_20;
  assign f_u_arrmul24_and20_20_y0 = f_u_arrmul24_and20_20_a_20 & f_u_arrmul24_and20_20_b_20;
  assign f_u_arrmul24_fa20_20_f_u_arrmul24_and20_20_y0 = f_u_arrmul24_and20_20_y0;
  assign f_u_arrmul24_fa20_20_f_u_arrmul24_fa21_19_y2 = f_u_arrmul24_fa21_19_y2;
  assign f_u_arrmul24_fa20_20_f_u_arrmul24_fa19_20_y4 = f_u_arrmul24_fa19_20_y4;
  assign f_u_arrmul24_fa20_20_y0 = f_u_arrmul24_fa20_20_f_u_arrmul24_and20_20_y0 ^ f_u_arrmul24_fa20_20_f_u_arrmul24_fa21_19_y2;
  assign f_u_arrmul24_fa20_20_y1 = f_u_arrmul24_fa20_20_f_u_arrmul24_and20_20_y0 & f_u_arrmul24_fa20_20_f_u_arrmul24_fa21_19_y2;
  assign f_u_arrmul24_fa20_20_y2 = f_u_arrmul24_fa20_20_y0 ^ f_u_arrmul24_fa20_20_f_u_arrmul24_fa19_20_y4;
  assign f_u_arrmul24_fa20_20_y3 = f_u_arrmul24_fa20_20_y0 & f_u_arrmul24_fa20_20_f_u_arrmul24_fa19_20_y4;
  assign f_u_arrmul24_fa20_20_y4 = f_u_arrmul24_fa20_20_y1 | f_u_arrmul24_fa20_20_y3;
  assign f_u_arrmul24_and21_20_a_21 = a_21;
  assign f_u_arrmul24_and21_20_b_20 = b_20;
  assign f_u_arrmul24_and21_20_y0 = f_u_arrmul24_and21_20_a_21 & f_u_arrmul24_and21_20_b_20;
  assign f_u_arrmul24_fa21_20_f_u_arrmul24_and21_20_y0 = f_u_arrmul24_and21_20_y0;
  assign f_u_arrmul24_fa21_20_f_u_arrmul24_fa22_19_y2 = f_u_arrmul24_fa22_19_y2;
  assign f_u_arrmul24_fa21_20_f_u_arrmul24_fa20_20_y4 = f_u_arrmul24_fa20_20_y4;
  assign f_u_arrmul24_fa21_20_y0 = f_u_arrmul24_fa21_20_f_u_arrmul24_and21_20_y0 ^ f_u_arrmul24_fa21_20_f_u_arrmul24_fa22_19_y2;
  assign f_u_arrmul24_fa21_20_y1 = f_u_arrmul24_fa21_20_f_u_arrmul24_and21_20_y0 & f_u_arrmul24_fa21_20_f_u_arrmul24_fa22_19_y2;
  assign f_u_arrmul24_fa21_20_y2 = f_u_arrmul24_fa21_20_y0 ^ f_u_arrmul24_fa21_20_f_u_arrmul24_fa20_20_y4;
  assign f_u_arrmul24_fa21_20_y3 = f_u_arrmul24_fa21_20_y0 & f_u_arrmul24_fa21_20_f_u_arrmul24_fa20_20_y4;
  assign f_u_arrmul24_fa21_20_y4 = f_u_arrmul24_fa21_20_y1 | f_u_arrmul24_fa21_20_y3;
  assign f_u_arrmul24_and22_20_a_22 = a_22;
  assign f_u_arrmul24_and22_20_b_20 = b_20;
  assign f_u_arrmul24_and22_20_y0 = f_u_arrmul24_and22_20_a_22 & f_u_arrmul24_and22_20_b_20;
  assign f_u_arrmul24_fa22_20_f_u_arrmul24_and22_20_y0 = f_u_arrmul24_and22_20_y0;
  assign f_u_arrmul24_fa22_20_f_u_arrmul24_fa23_19_y2 = f_u_arrmul24_fa23_19_y2;
  assign f_u_arrmul24_fa22_20_f_u_arrmul24_fa21_20_y4 = f_u_arrmul24_fa21_20_y4;
  assign f_u_arrmul24_fa22_20_y0 = f_u_arrmul24_fa22_20_f_u_arrmul24_and22_20_y0 ^ f_u_arrmul24_fa22_20_f_u_arrmul24_fa23_19_y2;
  assign f_u_arrmul24_fa22_20_y1 = f_u_arrmul24_fa22_20_f_u_arrmul24_and22_20_y0 & f_u_arrmul24_fa22_20_f_u_arrmul24_fa23_19_y2;
  assign f_u_arrmul24_fa22_20_y2 = f_u_arrmul24_fa22_20_y0 ^ f_u_arrmul24_fa22_20_f_u_arrmul24_fa21_20_y4;
  assign f_u_arrmul24_fa22_20_y3 = f_u_arrmul24_fa22_20_y0 & f_u_arrmul24_fa22_20_f_u_arrmul24_fa21_20_y4;
  assign f_u_arrmul24_fa22_20_y4 = f_u_arrmul24_fa22_20_y1 | f_u_arrmul24_fa22_20_y3;
  assign f_u_arrmul24_and23_20_a_23 = a_23;
  assign f_u_arrmul24_and23_20_b_20 = b_20;
  assign f_u_arrmul24_and23_20_y0 = f_u_arrmul24_and23_20_a_23 & f_u_arrmul24_and23_20_b_20;
  assign f_u_arrmul24_fa23_20_f_u_arrmul24_and23_20_y0 = f_u_arrmul24_and23_20_y0;
  assign f_u_arrmul24_fa23_20_f_u_arrmul24_fa23_19_y4 = f_u_arrmul24_fa23_19_y4;
  assign f_u_arrmul24_fa23_20_f_u_arrmul24_fa22_20_y4 = f_u_arrmul24_fa22_20_y4;
  assign f_u_arrmul24_fa23_20_y0 = f_u_arrmul24_fa23_20_f_u_arrmul24_and23_20_y0 ^ f_u_arrmul24_fa23_20_f_u_arrmul24_fa23_19_y4;
  assign f_u_arrmul24_fa23_20_y1 = f_u_arrmul24_fa23_20_f_u_arrmul24_and23_20_y0 & f_u_arrmul24_fa23_20_f_u_arrmul24_fa23_19_y4;
  assign f_u_arrmul24_fa23_20_y2 = f_u_arrmul24_fa23_20_y0 ^ f_u_arrmul24_fa23_20_f_u_arrmul24_fa22_20_y4;
  assign f_u_arrmul24_fa23_20_y3 = f_u_arrmul24_fa23_20_y0 & f_u_arrmul24_fa23_20_f_u_arrmul24_fa22_20_y4;
  assign f_u_arrmul24_fa23_20_y4 = f_u_arrmul24_fa23_20_y1 | f_u_arrmul24_fa23_20_y3;
  assign f_u_arrmul24_and0_21_a_0 = a_0;
  assign f_u_arrmul24_and0_21_b_21 = b_21;
  assign f_u_arrmul24_and0_21_y0 = f_u_arrmul24_and0_21_a_0 & f_u_arrmul24_and0_21_b_21;
  assign f_u_arrmul24_ha0_21_f_u_arrmul24_and0_21_y0 = f_u_arrmul24_and0_21_y0;
  assign f_u_arrmul24_ha0_21_f_u_arrmul24_fa1_20_y2 = f_u_arrmul24_fa1_20_y2;
  assign f_u_arrmul24_ha0_21_y0 = f_u_arrmul24_ha0_21_f_u_arrmul24_and0_21_y0 ^ f_u_arrmul24_ha0_21_f_u_arrmul24_fa1_20_y2;
  assign f_u_arrmul24_ha0_21_y1 = f_u_arrmul24_ha0_21_f_u_arrmul24_and0_21_y0 & f_u_arrmul24_ha0_21_f_u_arrmul24_fa1_20_y2;
  assign f_u_arrmul24_and1_21_a_1 = a_1;
  assign f_u_arrmul24_and1_21_b_21 = b_21;
  assign f_u_arrmul24_and1_21_y0 = f_u_arrmul24_and1_21_a_1 & f_u_arrmul24_and1_21_b_21;
  assign f_u_arrmul24_fa1_21_f_u_arrmul24_and1_21_y0 = f_u_arrmul24_and1_21_y0;
  assign f_u_arrmul24_fa1_21_f_u_arrmul24_fa2_20_y2 = f_u_arrmul24_fa2_20_y2;
  assign f_u_arrmul24_fa1_21_f_u_arrmul24_ha0_21_y1 = f_u_arrmul24_ha0_21_y1;
  assign f_u_arrmul24_fa1_21_y0 = f_u_arrmul24_fa1_21_f_u_arrmul24_and1_21_y0 ^ f_u_arrmul24_fa1_21_f_u_arrmul24_fa2_20_y2;
  assign f_u_arrmul24_fa1_21_y1 = f_u_arrmul24_fa1_21_f_u_arrmul24_and1_21_y0 & f_u_arrmul24_fa1_21_f_u_arrmul24_fa2_20_y2;
  assign f_u_arrmul24_fa1_21_y2 = f_u_arrmul24_fa1_21_y0 ^ f_u_arrmul24_fa1_21_f_u_arrmul24_ha0_21_y1;
  assign f_u_arrmul24_fa1_21_y3 = f_u_arrmul24_fa1_21_y0 & f_u_arrmul24_fa1_21_f_u_arrmul24_ha0_21_y1;
  assign f_u_arrmul24_fa1_21_y4 = f_u_arrmul24_fa1_21_y1 | f_u_arrmul24_fa1_21_y3;
  assign f_u_arrmul24_and2_21_a_2 = a_2;
  assign f_u_arrmul24_and2_21_b_21 = b_21;
  assign f_u_arrmul24_and2_21_y0 = f_u_arrmul24_and2_21_a_2 & f_u_arrmul24_and2_21_b_21;
  assign f_u_arrmul24_fa2_21_f_u_arrmul24_and2_21_y0 = f_u_arrmul24_and2_21_y0;
  assign f_u_arrmul24_fa2_21_f_u_arrmul24_fa3_20_y2 = f_u_arrmul24_fa3_20_y2;
  assign f_u_arrmul24_fa2_21_f_u_arrmul24_fa1_21_y4 = f_u_arrmul24_fa1_21_y4;
  assign f_u_arrmul24_fa2_21_y0 = f_u_arrmul24_fa2_21_f_u_arrmul24_and2_21_y0 ^ f_u_arrmul24_fa2_21_f_u_arrmul24_fa3_20_y2;
  assign f_u_arrmul24_fa2_21_y1 = f_u_arrmul24_fa2_21_f_u_arrmul24_and2_21_y0 & f_u_arrmul24_fa2_21_f_u_arrmul24_fa3_20_y2;
  assign f_u_arrmul24_fa2_21_y2 = f_u_arrmul24_fa2_21_y0 ^ f_u_arrmul24_fa2_21_f_u_arrmul24_fa1_21_y4;
  assign f_u_arrmul24_fa2_21_y3 = f_u_arrmul24_fa2_21_y0 & f_u_arrmul24_fa2_21_f_u_arrmul24_fa1_21_y4;
  assign f_u_arrmul24_fa2_21_y4 = f_u_arrmul24_fa2_21_y1 | f_u_arrmul24_fa2_21_y3;
  assign f_u_arrmul24_and3_21_a_3 = a_3;
  assign f_u_arrmul24_and3_21_b_21 = b_21;
  assign f_u_arrmul24_and3_21_y0 = f_u_arrmul24_and3_21_a_3 & f_u_arrmul24_and3_21_b_21;
  assign f_u_arrmul24_fa3_21_f_u_arrmul24_and3_21_y0 = f_u_arrmul24_and3_21_y0;
  assign f_u_arrmul24_fa3_21_f_u_arrmul24_fa4_20_y2 = f_u_arrmul24_fa4_20_y2;
  assign f_u_arrmul24_fa3_21_f_u_arrmul24_fa2_21_y4 = f_u_arrmul24_fa2_21_y4;
  assign f_u_arrmul24_fa3_21_y0 = f_u_arrmul24_fa3_21_f_u_arrmul24_and3_21_y0 ^ f_u_arrmul24_fa3_21_f_u_arrmul24_fa4_20_y2;
  assign f_u_arrmul24_fa3_21_y1 = f_u_arrmul24_fa3_21_f_u_arrmul24_and3_21_y0 & f_u_arrmul24_fa3_21_f_u_arrmul24_fa4_20_y2;
  assign f_u_arrmul24_fa3_21_y2 = f_u_arrmul24_fa3_21_y0 ^ f_u_arrmul24_fa3_21_f_u_arrmul24_fa2_21_y4;
  assign f_u_arrmul24_fa3_21_y3 = f_u_arrmul24_fa3_21_y0 & f_u_arrmul24_fa3_21_f_u_arrmul24_fa2_21_y4;
  assign f_u_arrmul24_fa3_21_y4 = f_u_arrmul24_fa3_21_y1 | f_u_arrmul24_fa3_21_y3;
  assign f_u_arrmul24_and4_21_a_4 = a_4;
  assign f_u_arrmul24_and4_21_b_21 = b_21;
  assign f_u_arrmul24_and4_21_y0 = f_u_arrmul24_and4_21_a_4 & f_u_arrmul24_and4_21_b_21;
  assign f_u_arrmul24_fa4_21_f_u_arrmul24_and4_21_y0 = f_u_arrmul24_and4_21_y0;
  assign f_u_arrmul24_fa4_21_f_u_arrmul24_fa5_20_y2 = f_u_arrmul24_fa5_20_y2;
  assign f_u_arrmul24_fa4_21_f_u_arrmul24_fa3_21_y4 = f_u_arrmul24_fa3_21_y4;
  assign f_u_arrmul24_fa4_21_y0 = f_u_arrmul24_fa4_21_f_u_arrmul24_and4_21_y0 ^ f_u_arrmul24_fa4_21_f_u_arrmul24_fa5_20_y2;
  assign f_u_arrmul24_fa4_21_y1 = f_u_arrmul24_fa4_21_f_u_arrmul24_and4_21_y0 & f_u_arrmul24_fa4_21_f_u_arrmul24_fa5_20_y2;
  assign f_u_arrmul24_fa4_21_y2 = f_u_arrmul24_fa4_21_y0 ^ f_u_arrmul24_fa4_21_f_u_arrmul24_fa3_21_y4;
  assign f_u_arrmul24_fa4_21_y3 = f_u_arrmul24_fa4_21_y0 & f_u_arrmul24_fa4_21_f_u_arrmul24_fa3_21_y4;
  assign f_u_arrmul24_fa4_21_y4 = f_u_arrmul24_fa4_21_y1 | f_u_arrmul24_fa4_21_y3;
  assign f_u_arrmul24_and5_21_a_5 = a_5;
  assign f_u_arrmul24_and5_21_b_21 = b_21;
  assign f_u_arrmul24_and5_21_y0 = f_u_arrmul24_and5_21_a_5 & f_u_arrmul24_and5_21_b_21;
  assign f_u_arrmul24_fa5_21_f_u_arrmul24_and5_21_y0 = f_u_arrmul24_and5_21_y0;
  assign f_u_arrmul24_fa5_21_f_u_arrmul24_fa6_20_y2 = f_u_arrmul24_fa6_20_y2;
  assign f_u_arrmul24_fa5_21_f_u_arrmul24_fa4_21_y4 = f_u_arrmul24_fa4_21_y4;
  assign f_u_arrmul24_fa5_21_y0 = f_u_arrmul24_fa5_21_f_u_arrmul24_and5_21_y0 ^ f_u_arrmul24_fa5_21_f_u_arrmul24_fa6_20_y2;
  assign f_u_arrmul24_fa5_21_y1 = f_u_arrmul24_fa5_21_f_u_arrmul24_and5_21_y0 & f_u_arrmul24_fa5_21_f_u_arrmul24_fa6_20_y2;
  assign f_u_arrmul24_fa5_21_y2 = f_u_arrmul24_fa5_21_y0 ^ f_u_arrmul24_fa5_21_f_u_arrmul24_fa4_21_y4;
  assign f_u_arrmul24_fa5_21_y3 = f_u_arrmul24_fa5_21_y0 & f_u_arrmul24_fa5_21_f_u_arrmul24_fa4_21_y4;
  assign f_u_arrmul24_fa5_21_y4 = f_u_arrmul24_fa5_21_y1 | f_u_arrmul24_fa5_21_y3;
  assign f_u_arrmul24_and6_21_a_6 = a_6;
  assign f_u_arrmul24_and6_21_b_21 = b_21;
  assign f_u_arrmul24_and6_21_y0 = f_u_arrmul24_and6_21_a_6 & f_u_arrmul24_and6_21_b_21;
  assign f_u_arrmul24_fa6_21_f_u_arrmul24_and6_21_y0 = f_u_arrmul24_and6_21_y0;
  assign f_u_arrmul24_fa6_21_f_u_arrmul24_fa7_20_y2 = f_u_arrmul24_fa7_20_y2;
  assign f_u_arrmul24_fa6_21_f_u_arrmul24_fa5_21_y4 = f_u_arrmul24_fa5_21_y4;
  assign f_u_arrmul24_fa6_21_y0 = f_u_arrmul24_fa6_21_f_u_arrmul24_and6_21_y0 ^ f_u_arrmul24_fa6_21_f_u_arrmul24_fa7_20_y2;
  assign f_u_arrmul24_fa6_21_y1 = f_u_arrmul24_fa6_21_f_u_arrmul24_and6_21_y0 & f_u_arrmul24_fa6_21_f_u_arrmul24_fa7_20_y2;
  assign f_u_arrmul24_fa6_21_y2 = f_u_arrmul24_fa6_21_y0 ^ f_u_arrmul24_fa6_21_f_u_arrmul24_fa5_21_y4;
  assign f_u_arrmul24_fa6_21_y3 = f_u_arrmul24_fa6_21_y0 & f_u_arrmul24_fa6_21_f_u_arrmul24_fa5_21_y4;
  assign f_u_arrmul24_fa6_21_y4 = f_u_arrmul24_fa6_21_y1 | f_u_arrmul24_fa6_21_y3;
  assign f_u_arrmul24_and7_21_a_7 = a_7;
  assign f_u_arrmul24_and7_21_b_21 = b_21;
  assign f_u_arrmul24_and7_21_y0 = f_u_arrmul24_and7_21_a_7 & f_u_arrmul24_and7_21_b_21;
  assign f_u_arrmul24_fa7_21_f_u_arrmul24_and7_21_y0 = f_u_arrmul24_and7_21_y0;
  assign f_u_arrmul24_fa7_21_f_u_arrmul24_fa8_20_y2 = f_u_arrmul24_fa8_20_y2;
  assign f_u_arrmul24_fa7_21_f_u_arrmul24_fa6_21_y4 = f_u_arrmul24_fa6_21_y4;
  assign f_u_arrmul24_fa7_21_y0 = f_u_arrmul24_fa7_21_f_u_arrmul24_and7_21_y0 ^ f_u_arrmul24_fa7_21_f_u_arrmul24_fa8_20_y2;
  assign f_u_arrmul24_fa7_21_y1 = f_u_arrmul24_fa7_21_f_u_arrmul24_and7_21_y0 & f_u_arrmul24_fa7_21_f_u_arrmul24_fa8_20_y2;
  assign f_u_arrmul24_fa7_21_y2 = f_u_arrmul24_fa7_21_y0 ^ f_u_arrmul24_fa7_21_f_u_arrmul24_fa6_21_y4;
  assign f_u_arrmul24_fa7_21_y3 = f_u_arrmul24_fa7_21_y0 & f_u_arrmul24_fa7_21_f_u_arrmul24_fa6_21_y4;
  assign f_u_arrmul24_fa7_21_y4 = f_u_arrmul24_fa7_21_y1 | f_u_arrmul24_fa7_21_y3;
  assign f_u_arrmul24_and8_21_a_8 = a_8;
  assign f_u_arrmul24_and8_21_b_21 = b_21;
  assign f_u_arrmul24_and8_21_y0 = f_u_arrmul24_and8_21_a_8 & f_u_arrmul24_and8_21_b_21;
  assign f_u_arrmul24_fa8_21_f_u_arrmul24_and8_21_y0 = f_u_arrmul24_and8_21_y0;
  assign f_u_arrmul24_fa8_21_f_u_arrmul24_fa9_20_y2 = f_u_arrmul24_fa9_20_y2;
  assign f_u_arrmul24_fa8_21_f_u_arrmul24_fa7_21_y4 = f_u_arrmul24_fa7_21_y4;
  assign f_u_arrmul24_fa8_21_y0 = f_u_arrmul24_fa8_21_f_u_arrmul24_and8_21_y0 ^ f_u_arrmul24_fa8_21_f_u_arrmul24_fa9_20_y2;
  assign f_u_arrmul24_fa8_21_y1 = f_u_arrmul24_fa8_21_f_u_arrmul24_and8_21_y0 & f_u_arrmul24_fa8_21_f_u_arrmul24_fa9_20_y2;
  assign f_u_arrmul24_fa8_21_y2 = f_u_arrmul24_fa8_21_y0 ^ f_u_arrmul24_fa8_21_f_u_arrmul24_fa7_21_y4;
  assign f_u_arrmul24_fa8_21_y3 = f_u_arrmul24_fa8_21_y0 & f_u_arrmul24_fa8_21_f_u_arrmul24_fa7_21_y4;
  assign f_u_arrmul24_fa8_21_y4 = f_u_arrmul24_fa8_21_y1 | f_u_arrmul24_fa8_21_y3;
  assign f_u_arrmul24_and9_21_a_9 = a_9;
  assign f_u_arrmul24_and9_21_b_21 = b_21;
  assign f_u_arrmul24_and9_21_y0 = f_u_arrmul24_and9_21_a_9 & f_u_arrmul24_and9_21_b_21;
  assign f_u_arrmul24_fa9_21_f_u_arrmul24_and9_21_y0 = f_u_arrmul24_and9_21_y0;
  assign f_u_arrmul24_fa9_21_f_u_arrmul24_fa10_20_y2 = f_u_arrmul24_fa10_20_y2;
  assign f_u_arrmul24_fa9_21_f_u_arrmul24_fa8_21_y4 = f_u_arrmul24_fa8_21_y4;
  assign f_u_arrmul24_fa9_21_y0 = f_u_arrmul24_fa9_21_f_u_arrmul24_and9_21_y0 ^ f_u_arrmul24_fa9_21_f_u_arrmul24_fa10_20_y2;
  assign f_u_arrmul24_fa9_21_y1 = f_u_arrmul24_fa9_21_f_u_arrmul24_and9_21_y0 & f_u_arrmul24_fa9_21_f_u_arrmul24_fa10_20_y2;
  assign f_u_arrmul24_fa9_21_y2 = f_u_arrmul24_fa9_21_y0 ^ f_u_arrmul24_fa9_21_f_u_arrmul24_fa8_21_y4;
  assign f_u_arrmul24_fa9_21_y3 = f_u_arrmul24_fa9_21_y0 & f_u_arrmul24_fa9_21_f_u_arrmul24_fa8_21_y4;
  assign f_u_arrmul24_fa9_21_y4 = f_u_arrmul24_fa9_21_y1 | f_u_arrmul24_fa9_21_y3;
  assign f_u_arrmul24_and10_21_a_10 = a_10;
  assign f_u_arrmul24_and10_21_b_21 = b_21;
  assign f_u_arrmul24_and10_21_y0 = f_u_arrmul24_and10_21_a_10 & f_u_arrmul24_and10_21_b_21;
  assign f_u_arrmul24_fa10_21_f_u_arrmul24_and10_21_y0 = f_u_arrmul24_and10_21_y0;
  assign f_u_arrmul24_fa10_21_f_u_arrmul24_fa11_20_y2 = f_u_arrmul24_fa11_20_y2;
  assign f_u_arrmul24_fa10_21_f_u_arrmul24_fa9_21_y4 = f_u_arrmul24_fa9_21_y4;
  assign f_u_arrmul24_fa10_21_y0 = f_u_arrmul24_fa10_21_f_u_arrmul24_and10_21_y0 ^ f_u_arrmul24_fa10_21_f_u_arrmul24_fa11_20_y2;
  assign f_u_arrmul24_fa10_21_y1 = f_u_arrmul24_fa10_21_f_u_arrmul24_and10_21_y0 & f_u_arrmul24_fa10_21_f_u_arrmul24_fa11_20_y2;
  assign f_u_arrmul24_fa10_21_y2 = f_u_arrmul24_fa10_21_y0 ^ f_u_arrmul24_fa10_21_f_u_arrmul24_fa9_21_y4;
  assign f_u_arrmul24_fa10_21_y3 = f_u_arrmul24_fa10_21_y0 & f_u_arrmul24_fa10_21_f_u_arrmul24_fa9_21_y4;
  assign f_u_arrmul24_fa10_21_y4 = f_u_arrmul24_fa10_21_y1 | f_u_arrmul24_fa10_21_y3;
  assign f_u_arrmul24_and11_21_a_11 = a_11;
  assign f_u_arrmul24_and11_21_b_21 = b_21;
  assign f_u_arrmul24_and11_21_y0 = f_u_arrmul24_and11_21_a_11 & f_u_arrmul24_and11_21_b_21;
  assign f_u_arrmul24_fa11_21_f_u_arrmul24_and11_21_y0 = f_u_arrmul24_and11_21_y0;
  assign f_u_arrmul24_fa11_21_f_u_arrmul24_fa12_20_y2 = f_u_arrmul24_fa12_20_y2;
  assign f_u_arrmul24_fa11_21_f_u_arrmul24_fa10_21_y4 = f_u_arrmul24_fa10_21_y4;
  assign f_u_arrmul24_fa11_21_y0 = f_u_arrmul24_fa11_21_f_u_arrmul24_and11_21_y0 ^ f_u_arrmul24_fa11_21_f_u_arrmul24_fa12_20_y2;
  assign f_u_arrmul24_fa11_21_y1 = f_u_arrmul24_fa11_21_f_u_arrmul24_and11_21_y0 & f_u_arrmul24_fa11_21_f_u_arrmul24_fa12_20_y2;
  assign f_u_arrmul24_fa11_21_y2 = f_u_arrmul24_fa11_21_y0 ^ f_u_arrmul24_fa11_21_f_u_arrmul24_fa10_21_y4;
  assign f_u_arrmul24_fa11_21_y3 = f_u_arrmul24_fa11_21_y0 & f_u_arrmul24_fa11_21_f_u_arrmul24_fa10_21_y4;
  assign f_u_arrmul24_fa11_21_y4 = f_u_arrmul24_fa11_21_y1 | f_u_arrmul24_fa11_21_y3;
  assign f_u_arrmul24_and12_21_a_12 = a_12;
  assign f_u_arrmul24_and12_21_b_21 = b_21;
  assign f_u_arrmul24_and12_21_y0 = f_u_arrmul24_and12_21_a_12 & f_u_arrmul24_and12_21_b_21;
  assign f_u_arrmul24_fa12_21_f_u_arrmul24_and12_21_y0 = f_u_arrmul24_and12_21_y0;
  assign f_u_arrmul24_fa12_21_f_u_arrmul24_fa13_20_y2 = f_u_arrmul24_fa13_20_y2;
  assign f_u_arrmul24_fa12_21_f_u_arrmul24_fa11_21_y4 = f_u_arrmul24_fa11_21_y4;
  assign f_u_arrmul24_fa12_21_y0 = f_u_arrmul24_fa12_21_f_u_arrmul24_and12_21_y0 ^ f_u_arrmul24_fa12_21_f_u_arrmul24_fa13_20_y2;
  assign f_u_arrmul24_fa12_21_y1 = f_u_arrmul24_fa12_21_f_u_arrmul24_and12_21_y0 & f_u_arrmul24_fa12_21_f_u_arrmul24_fa13_20_y2;
  assign f_u_arrmul24_fa12_21_y2 = f_u_arrmul24_fa12_21_y0 ^ f_u_arrmul24_fa12_21_f_u_arrmul24_fa11_21_y4;
  assign f_u_arrmul24_fa12_21_y3 = f_u_arrmul24_fa12_21_y0 & f_u_arrmul24_fa12_21_f_u_arrmul24_fa11_21_y4;
  assign f_u_arrmul24_fa12_21_y4 = f_u_arrmul24_fa12_21_y1 | f_u_arrmul24_fa12_21_y3;
  assign f_u_arrmul24_and13_21_a_13 = a_13;
  assign f_u_arrmul24_and13_21_b_21 = b_21;
  assign f_u_arrmul24_and13_21_y0 = f_u_arrmul24_and13_21_a_13 & f_u_arrmul24_and13_21_b_21;
  assign f_u_arrmul24_fa13_21_f_u_arrmul24_and13_21_y0 = f_u_arrmul24_and13_21_y0;
  assign f_u_arrmul24_fa13_21_f_u_arrmul24_fa14_20_y2 = f_u_arrmul24_fa14_20_y2;
  assign f_u_arrmul24_fa13_21_f_u_arrmul24_fa12_21_y4 = f_u_arrmul24_fa12_21_y4;
  assign f_u_arrmul24_fa13_21_y0 = f_u_arrmul24_fa13_21_f_u_arrmul24_and13_21_y0 ^ f_u_arrmul24_fa13_21_f_u_arrmul24_fa14_20_y2;
  assign f_u_arrmul24_fa13_21_y1 = f_u_arrmul24_fa13_21_f_u_arrmul24_and13_21_y0 & f_u_arrmul24_fa13_21_f_u_arrmul24_fa14_20_y2;
  assign f_u_arrmul24_fa13_21_y2 = f_u_arrmul24_fa13_21_y0 ^ f_u_arrmul24_fa13_21_f_u_arrmul24_fa12_21_y4;
  assign f_u_arrmul24_fa13_21_y3 = f_u_arrmul24_fa13_21_y0 & f_u_arrmul24_fa13_21_f_u_arrmul24_fa12_21_y4;
  assign f_u_arrmul24_fa13_21_y4 = f_u_arrmul24_fa13_21_y1 | f_u_arrmul24_fa13_21_y3;
  assign f_u_arrmul24_and14_21_a_14 = a_14;
  assign f_u_arrmul24_and14_21_b_21 = b_21;
  assign f_u_arrmul24_and14_21_y0 = f_u_arrmul24_and14_21_a_14 & f_u_arrmul24_and14_21_b_21;
  assign f_u_arrmul24_fa14_21_f_u_arrmul24_and14_21_y0 = f_u_arrmul24_and14_21_y0;
  assign f_u_arrmul24_fa14_21_f_u_arrmul24_fa15_20_y2 = f_u_arrmul24_fa15_20_y2;
  assign f_u_arrmul24_fa14_21_f_u_arrmul24_fa13_21_y4 = f_u_arrmul24_fa13_21_y4;
  assign f_u_arrmul24_fa14_21_y0 = f_u_arrmul24_fa14_21_f_u_arrmul24_and14_21_y0 ^ f_u_arrmul24_fa14_21_f_u_arrmul24_fa15_20_y2;
  assign f_u_arrmul24_fa14_21_y1 = f_u_arrmul24_fa14_21_f_u_arrmul24_and14_21_y0 & f_u_arrmul24_fa14_21_f_u_arrmul24_fa15_20_y2;
  assign f_u_arrmul24_fa14_21_y2 = f_u_arrmul24_fa14_21_y0 ^ f_u_arrmul24_fa14_21_f_u_arrmul24_fa13_21_y4;
  assign f_u_arrmul24_fa14_21_y3 = f_u_arrmul24_fa14_21_y0 & f_u_arrmul24_fa14_21_f_u_arrmul24_fa13_21_y4;
  assign f_u_arrmul24_fa14_21_y4 = f_u_arrmul24_fa14_21_y1 | f_u_arrmul24_fa14_21_y3;
  assign f_u_arrmul24_and15_21_a_15 = a_15;
  assign f_u_arrmul24_and15_21_b_21 = b_21;
  assign f_u_arrmul24_and15_21_y0 = f_u_arrmul24_and15_21_a_15 & f_u_arrmul24_and15_21_b_21;
  assign f_u_arrmul24_fa15_21_f_u_arrmul24_and15_21_y0 = f_u_arrmul24_and15_21_y0;
  assign f_u_arrmul24_fa15_21_f_u_arrmul24_fa16_20_y2 = f_u_arrmul24_fa16_20_y2;
  assign f_u_arrmul24_fa15_21_f_u_arrmul24_fa14_21_y4 = f_u_arrmul24_fa14_21_y4;
  assign f_u_arrmul24_fa15_21_y0 = f_u_arrmul24_fa15_21_f_u_arrmul24_and15_21_y0 ^ f_u_arrmul24_fa15_21_f_u_arrmul24_fa16_20_y2;
  assign f_u_arrmul24_fa15_21_y1 = f_u_arrmul24_fa15_21_f_u_arrmul24_and15_21_y0 & f_u_arrmul24_fa15_21_f_u_arrmul24_fa16_20_y2;
  assign f_u_arrmul24_fa15_21_y2 = f_u_arrmul24_fa15_21_y0 ^ f_u_arrmul24_fa15_21_f_u_arrmul24_fa14_21_y4;
  assign f_u_arrmul24_fa15_21_y3 = f_u_arrmul24_fa15_21_y0 & f_u_arrmul24_fa15_21_f_u_arrmul24_fa14_21_y4;
  assign f_u_arrmul24_fa15_21_y4 = f_u_arrmul24_fa15_21_y1 | f_u_arrmul24_fa15_21_y3;
  assign f_u_arrmul24_and16_21_a_16 = a_16;
  assign f_u_arrmul24_and16_21_b_21 = b_21;
  assign f_u_arrmul24_and16_21_y0 = f_u_arrmul24_and16_21_a_16 & f_u_arrmul24_and16_21_b_21;
  assign f_u_arrmul24_fa16_21_f_u_arrmul24_and16_21_y0 = f_u_arrmul24_and16_21_y0;
  assign f_u_arrmul24_fa16_21_f_u_arrmul24_fa17_20_y2 = f_u_arrmul24_fa17_20_y2;
  assign f_u_arrmul24_fa16_21_f_u_arrmul24_fa15_21_y4 = f_u_arrmul24_fa15_21_y4;
  assign f_u_arrmul24_fa16_21_y0 = f_u_arrmul24_fa16_21_f_u_arrmul24_and16_21_y0 ^ f_u_arrmul24_fa16_21_f_u_arrmul24_fa17_20_y2;
  assign f_u_arrmul24_fa16_21_y1 = f_u_arrmul24_fa16_21_f_u_arrmul24_and16_21_y0 & f_u_arrmul24_fa16_21_f_u_arrmul24_fa17_20_y2;
  assign f_u_arrmul24_fa16_21_y2 = f_u_arrmul24_fa16_21_y0 ^ f_u_arrmul24_fa16_21_f_u_arrmul24_fa15_21_y4;
  assign f_u_arrmul24_fa16_21_y3 = f_u_arrmul24_fa16_21_y0 & f_u_arrmul24_fa16_21_f_u_arrmul24_fa15_21_y4;
  assign f_u_arrmul24_fa16_21_y4 = f_u_arrmul24_fa16_21_y1 | f_u_arrmul24_fa16_21_y3;
  assign f_u_arrmul24_and17_21_a_17 = a_17;
  assign f_u_arrmul24_and17_21_b_21 = b_21;
  assign f_u_arrmul24_and17_21_y0 = f_u_arrmul24_and17_21_a_17 & f_u_arrmul24_and17_21_b_21;
  assign f_u_arrmul24_fa17_21_f_u_arrmul24_and17_21_y0 = f_u_arrmul24_and17_21_y0;
  assign f_u_arrmul24_fa17_21_f_u_arrmul24_fa18_20_y2 = f_u_arrmul24_fa18_20_y2;
  assign f_u_arrmul24_fa17_21_f_u_arrmul24_fa16_21_y4 = f_u_arrmul24_fa16_21_y4;
  assign f_u_arrmul24_fa17_21_y0 = f_u_arrmul24_fa17_21_f_u_arrmul24_and17_21_y0 ^ f_u_arrmul24_fa17_21_f_u_arrmul24_fa18_20_y2;
  assign f_u_arrmul24_fa17_21_y1 = f_u_arrmul24_fa17_21_f_u_arrmul24_and17_21_y0 & f_u_arrmul24_fa17_21_f_u_arrmul24_fa18_20_y2;
  assign f_u_arrmul24_fa17_21_y2 = f_u_arrmul24_fa17_21_y0 ^ f_u_arrmul24_fa17_21_f_u_arrmul24_fa16_21_y4;
  assign f_u_arrmul24_fa17_21_y3 = f_u_arrmul24_fa17_21_y0 & f_u_arrmul24_fa17_21_f_u_arrmul24_fa16_21_y4;
  assign f_u_arrmul24_fa17_21_y4 = f_u_arrmul24_fa17_21_y1 | f_u_arrmul24_fa17_21_y3;
  assign f_u_arrmul24_and18_21_a_18 = a_18;
  assign f_u_arrmul24_and18_21_b_21 = b_21;
  assign f_u_arrmul24_and18_21_y0 = f_u_arrmul24_and18_21_a_18 & f_u_arrmul24_and18_21_b_21;
  assign f_u_arrmul24_fa18_21_f_u_arrmul24_and18_21_y0 = f_u_arrmul24_and18_21_y0;
  assign f_u_arrmul24_fa18_21_f_u_arrmul24_fa19_20_y2 = f_u_arrmul24_fa19_20_y2;
  assign f_u_arrmul24_fa18_21_f_u_arrmul24_fa17_21_y4 = f_u_arrmul24_fa17_21_y4;
  assign f_u_arrmul24_fa18_21_y0 = f_u_arrmul24_fa18_21_f_u_arrmul24_and18_21_y0 ^ f_u_arrmul24_fa18_21_f_u_arrmul24_fa19_20_y2;
  assign f_u_arrmul24_fa18_21_y1 = f_u_arrmul24_fa18_21_f_u_arrmul24_and18_21_y0 & f_u_arrmul24_fa18_21_f_u_arrmul24_fa19_20_y2;
  assign f_u_arrmul24_fa18_21_y2 = f_u_arrmul24_fa18_21_y0 ^ f_u_arrmul24_fa18_21_f_u_arrmul24_fa17_21_y4;
  assign f_u_arrmul24_fa18_21_y3 = f_u_arrmul24_fa18_21_y0 & f_u_arrmul24_fa18_21_f_u_arrmul24_fa17_21_y4;
  assign f_u_arrmul24_fa18_21_y4 = f_u_arrmul24_fa18_21_y1 | f_u_arrmul24_fa18_21_y3;
  assign f_u_arrmul24_and19_21_a_19 = a_19;
  assign f_u_arrmul24_and19_21_b_21 = b_21;
  assign f_u_arrmul24_and19_21_y0 = f_u_arrmul24_and19_21_a_19 & f_u_arrmul24_and19_21_b_21;
  assign f_u_arrmul24_fa19_21_f_u_arrmul24_and19_21_y0 = f_u_arrmul24_and19_21_y0;
  assign f_u_arrmul24_fa19_21_f_u_arrmul24_fa20_20_y2 = f_u_arrmul24_fa20_20_y2;
  assign f_u_arrmul24_fa19_21_f_u_arrmul24_fa18_21_y4 = f_u_arrmul24_fa18_21_y4;
  assign f_u_arrmul24_fa19_21_y0 = f_u_arrmul24_fa19_21_f_u_arrmul24_and19_21_y0 ^ f_u_arrmul24_fa19_21_f_u_arrmul24_fa20_20_y2;
  assign f_u_arrmul24_fa19_21_y1 = f_u_arrmul24_fa19_21_f_u_arrmul24_and19_21_y0 & f_u_arrmul24_fa19_21_f_u_arrmul24_fa20_20_y2;
  assign f_u_arrmul24_fa19_21_y2 = f_u_arrmul24_fa19_21_y0 ^ f_u_arrmul24_fa19_21_f_u_arrmul24_fa18_21_y4;
  assign f_u_arrmul24_fa19_21_y3 = f_u_arrmul24_fa19_21_y0 & f_u_arrmul24_fa19_21_f_u_arrmul24_fa18_21_y4;
  assign f_u_arrmul24_fa19_21_y4 = f_u_arrmul24_fa19_21_y1 | f_u_arrmul24_fa19_21_y3;
  assign f_u_arrmul24_and20_21_a_20 = a_20;
  assign f_u_arrmul24_and20_21_b_21 = b_21;
  assign f_u_arrmul24_and20_21_y0 = f_u_arrmul24_and20_21_a_20 & f_u_arrmul24_and20_21_b_21;
  assign f_u_arrmul24_fa20_21_f_u_arrmul24_and20_21_y0 = f_u_arrmul24_and20_21_y0;
  assign f_u_arrmul24_fa20_21_f_u_arrmul24_fa21_20_y2 = f_u_arrmul24_fa21_20_y2;
  assign f_u_arrmul24_fa20_21_f_u_arrmul24_fa19_21_y4 = f_u_arrmul24_fa19_21_y4;
  assign f_u_arrmul24_fa20_21_y0 = f_u_arrmul24_fa20_21_f_u_arrmul24_and20_21_y0 ^ f_u_arrmul24_fa20_21_f_u_arrmul24_fa21_20_y2;
  assign f_u_arrmul24_fa20_21_y1 = f_u_arrmul24_fa20_21_f_u_arrmul24_and20_21_y0 & f_u_arrmul24_fa20_21_f_u_arrmul24_fa21_20_y2;
  assign f_u_arrmul24_fa20_21_y2 = f_u_arrmul24_fa20_21_y0 ^ f_u_arrmul24_fa20_21_f_u_arrmul24_fa19_21_y4;
  assign f_u_arrmul24_fa20_21_y3 = f_u_arrmul24_fa20_21_y0 & f_u_arrmul24_fa20_21_f_u_arrmul24_fa19_21_y4;
  assign f_u_arrmul24_fa20_21_y4 = f_u_arrmul24_fa20_21_y1 | f_u_arrmul24_fa20_21_y3;
  assign f_u_arrmul24_and21_21_a_21 = a_21;
  assign f_u_arrmul24_and21_21_b_21 = b_21;
  assign f_u_arrmul24_and21_21_y0 = f_u_arrmul24_and21_21_a_21 & f_u_arrmul24_and21_21_b_21;
  assign f_u_arrmul24_fa21_21_f_u_arrmul24_and21_21_y0 = f_u_arrmul24_and21_21_y0;
  assign f_u_arrmul24_fa21_21_f_u_arrmul24_fa22_20_y2 = f_u_arrmul24_fa22_20_y2;
  assign f_u_arrmul24_fa21_21_f_u_arrmul24_fa20_21_y4 = f_u_arrmul24_fa20_21_y4;
  assign f_u_arrmul24_fa21_21_y0 = f_u_arrmul24_fa21_21_f_u_arrmul24_and21_21_y0 ^ f_u_arrmul24_fa21_21_f_u_arrmul24_fa22_20_y2;
  assign f_u_arrmul24_fa21_21_y1 = f_u_arrmul24_fa21_21_f_u_arrmul24_and21_21_y0 & f_u_arrmul24_fa21_21_f_u_arrmul24_fa22_20_y2;
  assign f_u_arrmul24_fa21_21_y2 = f_u_arrmul24_fa21_21_y0 ^ f_u_arrmul24_fa21_21_f_u_arrmul24_fa20_21_y4;
  assign f_u_arrmul24_fa21_21_y3 = f_u_arrmul24_fa21_21_y0 & f_u_arrmul24_fa21_21_f_u_arrmul24_fa20_21_y4;
  assign f_u_arrmul24_fa21_21_y4 = f_u_arrmul24_fa21_21_y1 | f_u_arrmul24_fa21_21_y3;
  assign f_u_arrmul24_and22_21_a_22 = a_22;
  assign f_u_arrmul24_and22_21_b_21 = b_21;
  assign f_u_arrmul24_and22_21_y0 = f_u_arrmul24_and22_21_a_22 & f_u_arrmul24_and22_21_b_21;
  assign f_u_arrmul24_fa22_21_f_u_arrmul24_and22_21_y0 = f_u_arrmul24_and22_21_y0;
  assign f_u_arrmul24_fa22_21_f_u_arrmul24_fa23_20_y2 = f_u_arrmul24_fa23_20_y2;
  assign f_u_arrmul24_fa22_21_f_u_arrmul24_fa21_21_y4 = f_u_arrmul24_fa21_21_y4;
  assign f_u_arrmul24_fa22_21_y0 = f_u_arrmul24_fa22_21_f_u_arrmul24_and22_21_y0 ^ f_u_arrmul24_fa22_21_f_u_arrmul24_fa23_20_y2;
  assign f_u_arrmul24_fa22_21_y1 = f_u_arrmul24_fa22_21_f_u_arrmul24_and22_21_y0 & f_u_arrmul24_fa22_21_f_u_arrmul24_fa23_20_y2;
  assign f_u_arrmul24_fa22_21_y2 = f_u_arrmul24_fa22_21_y0 ^ f_u_arrmul24_fa22_21_f_u_arrmul24_fa21_21_y4;
  assign f_u_arrmul24_fa22_21_y3 = f_u_arrmul24_fa22_21_y0 & f_u_arrmul24_fa22_21_f_u_arrmul24_fa21_21_y4;
  assign f_u_arrmul24_fa22_21_y4 = f_u_arrmul24_fa22_21_y1 | f_u_arrmul24_fa22_21_y3;
  assign f_u_arrmul24_and23_21_a_23 = a_23;
  assign f_u_arrmul24_and23_21_b_21 = b_21;
  assign f_u_arrmul24_and23_21_y0 = f_u_arrmul24_and23_21_a_23 & f_u_arrmul24_and23_21_b_21;
  assign f_u_arrmul24_fa23_21_f_u_arrmul24_and23_21_y0 = f_u_arrmul24_and23_21_y0;
  assign f_u_arrmul24_fa23_21_f_u_arrmul24_fa23_20_y4 = f_u_arrmul24_fa23_20_y4;
  assign f_u_arrmul24_fa23_21_f_u_arrmul24_fa22_21_y4 = f_u_arrmul24_fa22_21_y4;
  assign f_u_arrmul24_fa23_21_y0 = f_u_arrmul24_fa23_21_f_u_arrmul24_and23_21_y0 ^ f_u_arrmul24_fa23_21_f_u_arrmul24_fa23_20_y4;
  assign f_u_arrmul24_fa23_21_y1 = f_u_arrmul24_fa23_21_f_u_arrmul24_and23_21_y0 & f_u_arrmul24_fa23_21_f_u_arrmul24_fa23_20_y4;
  assign f_u_arrmul24_fa23_21_y2 = f_u_arrmul24_fa23_21_y0 ^ f_u_arrmul24_fa23_21_f_u_arrmul24_fa22_21_y4;
  assign f_u_arrmul24_fa23_21_y3 = f_u_arrmul24_fa23_21_y0 & f_u_arrmul24_fa23_21_f_u_arrmul24_fa22_21_y4;
  assign f_u_arrmul24_fa23_21_y4 = f_u_arrmul24_fa23_21_y1 | f_u_arrmul24_fa23_21_y3;
  assign f_u_arrmul24_and0_22_a_0 = a_0;
  assign f_u_arrmul24_and0_22_b_22 = b_22;
  assign f_u_arrmul24_and0_22_y0 = f_u_arrmul24_and0_22_a_0 & f_u_arrmul24_and0_22_b_22;
  assign f_u_arrmul24_ha0_22_f_u_arrmul24_and0_22_y0 = f_u_arrmul24_and0_22_y0;
  assign f_u_arrmul24_ha0_22_f_u_arrmul24_fa1_21_y2 = f_u_arrmul24_fa1_21_y2;
  assign f_u_arrmul24_ha0_22_y0 = f_u_arrmul24_ha0_22_f_u_arrmul24_and0_22_y0 ^ f_u_arrmul24_ha0_22_f_u_arrmul24_fa1_21_y2;
  assign f_u_arrmul24_ha0_22_y1 = f_u_arrmul24_ha0_22_f_u_arrmul24_and0_22_y0 & f_u_arrmul24_ha0_22_f_u_arrmul24_fa1_21_y2;
  assign f_u_arrmul24_and1_22_a_1 = a_1;
  assign f_u_arrmul24_and1_22_b_22 = b_22;
  assign f_u_arrmul24_and1_22_y0 = f_u_arrmul24_and1_22_a_1 & f_u_arrmul24_and1_22_b_22;
  assign f_u_arrmul24_fa1_22_f_u_arrmul24_and1_22_y0 = f_u_arrmul24_and1_22_y0;
  assign f_u_arrmul24_fa1_22_f_u_arrmul24_fa2_21_y2 = f_u_arrmul24_fa2_21_y2;
  assign f_u_arrmul24_fa1_22_f_u_arrmul24_ha0_22_y1 = f_u_arrmul24_ha0_22_y1;
  assign f_u_arrmul24_fa1_22_y0 = f_u_arrmul24_fa1_22_f_u_arrmul24_and1_22_y0 ^ f_u_arrmul24_fa1_22_f_u_arrmul24_fa2_21_y2;
  assign f_u_arrmul24_fa1_22_y1 = f_u_arrmul24_fa1_22_f_u_arrmul24_and1_22_y0 & f_u_arrmul24_fa1_22_f_u_arrmul24_fa2_21_y2;
  assign f_u_arrmul24_fa1_22_y2 = f_u_arrmul24_fa1_22_y0 ^ f_u_arrmul24_fa1_22_f_u_arrmul24_ha0_22_y1;
  assign f_u_arrmul24_fa1_22_y3 = f_u_arrmul24_fa1_22_y0 & f_u_arrmul24_fa1_22_f_u_arrmul24_ha0_22_y1;
  assign f_u_arrmul24_fa1_22_y4 = f_u_arrmul24_fa1_22_y1 | f_u_arrmul24_fa1_22_y3;
  assign f_u_arrmul24_and2_22_a_2 = a_2;
  assign f_u_arrmul24_and2_22_b_22 = b_22;
  assign f_u_arrmul24_and2_22_y0 = f_u_arrmul24_and2_22_a_2 & f_u_arrmul24_and2_22_b_22;
  assign f_u_arrmul24_fa2_22_f_u_arrmul24_and2_22_y0 = f_u_arrmul24_and2_22_y0;
  assign f_u_arrmul24_fa2_22_f_u_arrmul24_fa3_21_y2 = f_u_arrmul24_fa3_21_y2;
  assign f_u_arrmul24_fa2_22_f_u_arrmul24_fa1_22_y4 = f_u_arrmul24_fa1_22_y4;
  assign f_u_arrmul24_fa2_22_y0 = f_u_arrmul24_fa2_22_f_u_arrmul24_and2_22_y0 ^ f_u_arrmul24_fa2_22_f_u_arrmul24_fa3_21_y2;
  assign f_u_arrmul24_fa2_22_y1 = f_u_arrmul24_fa2_22_f_u_arrmul24_and2_22_y0 & f_u_arrmul24_fa2_22_f_u_arrmul24_fa3_21_y2;
  assign f_u_arrmul24_fa2_22_y2 = f_u_arrmul24_fa2_22_y0 ^ f_u_arrmul24_fa2_22_f_u_arrmul24_fa1_22_y4;
  assign f_u_arrmul24_fa2_22_y3 = f_u_arrmul24_fa2_22_y0 & f_u_arrmul24_fa2_22_f_u_arrmul24_fa1_22_y4;
  assign f_u_arrmul24_fa2_22_y4 = f_u_arrmul24_fa2_22_y1 | f_u_arrmul24_fa2_22_y3;
  assign f_u_arrmul24_and3_22_a_3 = a_3;
  assign f_u_arrmul24_and3_22_b_22 = b_22;
  assign f_u_arrmul24_and3_22_y0 = f_u_arrmul24_and3_22_a_3 & f_u_arrmul24_and3_22_b_22;
  assign f_u_arrmul24_fa3_22_f_u_arrmul24_and3_22_y0 = f_u_arrmul24_and3_22_y0;
  assign f_u_arrmul24_fa3_22_f_u_arrmul24_fa4_21_y2 = f_u_arrmul24_fa4_21_y2;
  assign f_u_arrmul24_fa3_22_f_u_arrmul24_fa2_22_y4 = f_u_arrmul24_fa2_22_y4;
  assign f_u_arrmul24_fa3_22_y0 = f_u_arrmul24_fa3_22_f_u_arrmul24_and3_22_y0 ^ f_u_arrmul24_fa3_22_f_u_arrmul24_fa4_21_y2;
  assign f_u_arrmul24_fa3_22_y1 = f_u_arrmul24_fa3_22_f_u_arrmul24_and3_22_y0 & f_u_arrmul24_fa3_22_f_u_arrmul24_fa4_21_y2;
  assign f_u_arrmul24_fa3_22_y2 = f_u_arrmul24_fa3_22_y0 ^ f_u_arrmul24_fa3_22_f_u_arrmul24_fa2_22_y4;
  assign f_u_arrmul24_fa3_22_y3 = f_u_arrmul24_fa3_22_y0 & f_u_arrmul24_fa3_22_f_u_arrmul24_fa2_22_y4;
  assign f_u_arrmul24_fa3_22_y4 = f_u_arrmul24_fa3_22_y1 | f_u_arrmul24_fa3_22_y3;
  assign f_u_arrmul24_and4_22_a_4 = a_4;
  assign f_u_arrmul24_and4_22_b_22 = b_22;
  assign f_u_arrmul24_and4_22_y0 = f_u_arrmul24_and4_22_a_4 & f_u_arrmul24_and4_22_b_22;
  assign f_u_arrmul24_fa4_22_f_u_arrmul24_and4_22_y0 = f_u_arrmul24_and4_22_y0;
  assign f_u_arrmul24_fa4_22_f_u_arrmul24_fa5_21_y2 = f_u_arrmul24_fa5_21_y2;
  assign f_u_arrmul24_fa4_22_f_u_arrmul24_fa3_22_y4 = f_u_arrmul24_fa3_22_y4;
  assign f_u_arrmul24_fa4_22_y0 = f_u_arrmul24_fa4_22_f_u_arrmul24_and4_22_y0 ^ f_u_arrmul24_fa4_22_f_u_arrmul24_fa5_21_y2;
  assign f_u_arrmul24_fa4_22_y1 = f_u_arrmul24_fa4_22_f_u_arrmul24_and4_22_y0 & f_u_arrmul24_fa4_22_f_u_arrmul24_fa5_21_y2;
  assign f_u_arrmul24_fa4_22_y2 = f_u_arrmul24_fa4_22_y0 ^ f_u_arrmul24_fa4_22_f_u_arrmul24_fa3_22_y4;
  assign f_u_arrmul24_fa4_22_y3 = f_u_arrmul24_fa4_22_y0 & f_u_arrmul24_fa4_22_f_u_arrmul24_fa3_22_y4;
  assign f_u_arrmul24_fa4_22_y4 = f_u_arrmul24_fa4_22_y1 | f_u_arrmul24_fa4_22_y3;
  assign f_u_arrmul24_and5_22_a_5 = a_5;
  assign f_u_arrmul24_and5_22_b_22 = b_22;
  assign f_u_arrmul24_and5_22_y0 = f_u_arrmul24_and5_22_a_5 & f_u_arrmul24_and5_22_b_22;
  assign f_u_arrmul24_fa5_22_f_u_arrmul24_and5_22_y0 = f_u_arrmul24_and5_22_y0;
  assign f_u_arrmul24_fa5_22_f_u_arrmul24_fa6_21_y2 = f_u_arrmul24_fa6_21_y2;
  assign f_u_arrmul24_fa5_22_f_u_arrmul24_fa4_22_y4 = f_u_arrmul24_fa4_22_y4;
  assign f_u_arrmul24_fa5_22_y0 = f_u_arrmul24_fa5_22_f_u_arrmul24_and5_22_y0 ^ f_u_arrmul24_fa5_22_f_u_arrmul24_fa6_21_y2;
  assign f_u_arrmul24_fa5_22_y1 = f_u_arrmul24_fa5_22_f_u_arrmul24_and5_22_y0 & f_u_arrmul24_fa5_22_f_u_arrmul24_fa6_21_y2;
  assign f_u_arrmul24_fa5_22_y2 = f_u_arrmul24_fa5_22_y0 ^ f_u_arrmul24_fa5_22_f_u_arrmul24_fa4_22_y4;
  assign f_u_arrmul24_fa5_22_y3 = f_u_arrmul24_fa5_22_y0 & f_u_arrmul24_fa5_22_f_u_arrmul24_fa4_22_y4;
  assign f_u_arrmul24_fa5_22_y4 = f_u_arrmul24_fa5_22_y1 | f_u_arrmul24_fa5_22_y3;
  assign f_u_arrmul24_and6_22_a_6 = a_6;
  assign f_u_arrmul24_and6_22_b_22 = b_22;
  assign f_u_arrmul24_and6_22_y0 = f_u_arrmul24_and6_22_a_6 & f_u_arrmul24_and6_22_b_22;
  assign f_u_arrmul24_fa6_22_f_u_arrmul24_and6_22_y0 = f_u_arrmul24_and6_22_y0;
  assign f_u_arrmul24_fa6_22_f_u_arrmul24_fa7_21_y2 = f_u_arrmul24_fa7_21_y2;
  assign f_u_arrmul24_fa6_22_f_u_arrmul24_fa5_22_y4 = f_u_arrmul24_fa5_22_y4;
  assign f_u_arrmul24_fa6_22_y0 = f_u_arrmul24_fa6_22_f_u_arrmul24_and6_22_y0 ^ f_u_arrmul24_fa6_22_f_u_arrmul24_fa7_21_y2;
  assign f_u_arrmul24_fa6_22_y1 = f_u_arrmul24_fa6_22_f_u_arrmul24_and6_22_y0 & f_u_arrmul24_fa6_22_f_u_arrmul24_fa7_21_y2;
  assign f_u_arrmul24_fa6_22_y2 = f_u_arrmul24_fa6_22_y0 ^ f_u_arrmul24_fa6_22_f_u_arrmul24_fa5_22_y4;
  assign f_u_arrmul24_fa6_22_y3 = f_u_arrmul24_fa6_22_y0 & f_u_arrmul24_fa6_22_f_u_arrmul24_fa5_22_y4;
  assign f_u_arrmul24_fa6_22_y4 = f_u_arrmul24_fa6_22_y1 | f_u_arrmul24_fa6_22_y3;
  assign f_u_arrmul24_and7_22_a_7 = a_7;
  assign f_u_arrmul24_and7_22_b_22 = b_22;
  assign f_u_arrmul24_and7_22_y0 = f_u_arrmul24_and7_22_a_7 & f_u_arrmul24_and7_22_b_22;
  assign f_u_arrmul24_fa7_22_f_u_arrmul24_and7_22_y0 = f_u_arrmul24_and7_22_y0;
  assign f_u_arrmul24_fa7_22_f_u_arrmul24_fa8_21_y2 = f_u_arrmul24_fa8_21_y2;
  assign f_u_arrmul24_fa7_22_f_u_arrmul24_fa6_22_y4 = f_u_arrmul24_fa6_22_y4;
  assign f_u_arrmul24_fa7_22_y0 = f_u_arrmul24_fa7_22_f_u_arrmul24_and7_22_y0 ^ f_u_arrmul24_fa7_22_f_u_arrmul24_fa8_21_y2;
  assign f_u_arrmul24_fa7_22_y1 = f_u_arrmul24_fa7_22_f_u_arrmul24_and7_22_y0 & f_u_arrmul24_fa7_22_f_u_arrmul24_fa8_21_y2;
  assign f_u_arrmul24_fa7_22_y2 = f_u_arrmul24_fa7_22_y0 ^ f_u_arrmul24_fa7_22_f_u_arrmul24_fa6_22_y4;
  assign f_u_arrmul24_fa7_22_y3 = f_u_arrmul24_fa7_22_y0 & f_u_arrmul24_fa7_22_f_u_arrmul24_fa6_22_y4;
  assign f_u_arrmul24_fa7_22_y4 = f_u_arrmul24_fa7_22_y1 | f_u_arrmul24_fa7_22_y3;
  assign f_u_arrmul24_and8_22_a_8 = a_8;
  assign f_u_arrmul24_and8_22_b_22 = b_22;
  assign f_u_arrmul24_and8_22_y0 = f_u_arrmul24_and8_22_a_8 & f_u_arrmul24_and8_22_b_22;
  assign f_u_arrmul24_fa8_22_f_u_arrmul24_and8_22_y0 = f_u_arrmul24_and8_22_y0;
  assign f_u_arrmul24_fa8_22_f_u_arrmul24_fa9_21_y2 = f_u_arrmul24_fa9_21_y2;
  assign f_u_arrmul24_fa8_22_f_u_arrmul24_fa7_22_y4 = f_u_arrmul24_fa7_22_y4;
  assign f_u_arrmul24_fa8_22_y0 = f_u_arrmul24_fa8_22_f_u_arrmul24_and8_22_y0 ^ f_u_arrmul24_fa8_22_f_u_arrmul24_fa9_21_y2;
  assign f_u_arrmul24_fa8_22_y1 = f_u_arrmul24_fa8_22_f_u_arrmul24_and8_22_y0 & f_u_arrmul24_fa8_22_f_u_arrmul24_fa9_21_y2;
  assign f_u_arrmul24_fa8_22_y2 = f_u_arrmul24_fa8_22_y0 ^ f_u_arrmul24_fa8_22_f_u_arrmul24_fa7_22_y4;
  assign f_u_arrmul24_fa8_22_y3 = f_u_arrmul24_fa8_22_y0 & f_u_arrmul24_fa8_22_f_u_arrmul24_fa7_22_y4;
  assign f_u_arrmul24_fa8_22_y4 = f_u_arrmul24_fa8_22_y1 | f_u_arrmul24_fa8_22_y3;
  assign f_u_arrmul24_and9_22_a_9 = a_9;
  assign f_u_arrmul24_and9_22_b_22 = b_22;
  assign f_u_arrmul24_and9_22_y0 = f_u_arrmul24_and9_22_a_9 & f_u_arrmul24_and9_22_b_22;
  assign f_u_arrmul24_fa9_22_f_u_arrmul24_and9_22_y0 = f_u_arrmul24_and9_22_y0;
  assign f_u_arrmul24_fa9_22_f_u_arrmul24_fa10_21_y2 = f_u_arrmul24_fa10_21_y2;
  assign f_u_arrmul24_fa9_22_f_u_arrmul24_fa8_22_y4 = f_u_arrmul24_fa8_22_y4;
  assign f_u_arrmul24_fa9_22_y0 = f_u_arrmul24_fa9_22_f_u_arrmul24_and9_22_y0 ^ f_u_arrmul24_fa9_22_f_u_arrmul24_fa10_21_y2;
  assign f_u_arrmul24_fa9_22_y1 = f_u_arrmul24_fa9_22_f_u_arrmul24_and9_22_y0 & f_u_arrmul24_fa9_22_f_u_arrmul24_fa10_21_y2;
  assign f_u_arrmul24_fa9_22_y2 = f_u_arrmul24_fa9_22_y0 ^ f_u_arrmul24_fa9_22_f_u_arrmul24_fa8_22_y4;
  assign f_u_arrmul24_fa9_22_y3 = f_u_arrmul24_fa9_22_y0 & f_u_arrmul24_fa9_22_f_u_arrmul24_fa8_22_y4;
  assign f_u_arrmul24_fa9_22_y4 = f_u_arrmul24_fa9_22_y1 | f_u_arrmul24_fa9_22_y3;
  assign f_u_arrmul24_and10_22_a_10 = a_10;
  assign f_u_arrmul24_and10_22_b_22 = b_22;
  assign f_u_arrmul24_and10_22_y0 = f_u_arrmul24_and10_22_a_10 & f_u_arrmul24_and10_22_b_22;
  assign f_u_arrmul24_fa10_22_f_u_arrmul24_and10_22_y0 = f_u_arrmul24_and10_22_y0;
  assign f_u_arrmul24_fa10_22_f_u_arrmul24_fa11_21_y2 = f_u_arrmul24_fa11_21_y2;
  assign f_u_arrmul24_fa10_22_f_u_arrmul24_fa9_22_y4 = f_u_arrmul24_fa9_22_y4;
  assign f_u_arrmul24_fa10_22_y0 = f_u_arrmul24_fa10_22_f_u_arrmul24_and10_22_y0 ^ f_u_arrmul24_fa10_22_f_u_arrmul24_fa11_21_y2;
  assign f_u_arrmul24_fa10_22_y1 = f_u_arrmul24_fa10_22_f_u_arrmul24_and10_22_y0 & f_u_arrmul24_fa10_22_f_u_arrmul24_fa11_21_y2;
  assign f_u_arrmul24_fa10_22_y2 = f_u_arrmul24_fa10_22_y0 ^ f_u_arrmul24_fa10_22_f_u_arrmul24_fa9_22_y4;
  assign f_u_arrmul24_fa10_22_y3 = f_u_arrmul24_fa10_22_y0 & f_u_arrmul24_fa10_22_f_u_arrmul24_fa9_22_y4;
  assign f_u_arrmul24_fa10_22_y4 = f_u_arrmul24_fa10_22_y1 | f_u_arrmul24_fa10_22_y3;
  assign f_u_arrmul24_and11_22_a_11 = a_11;
  assign f_u_arrmul24_and11_22_b_22 = b_22;
  assign f_u_arrmul24_and11_22_y0 = f_u_arrmul24_and11_22_a_11 & f_u_arrmul24_and11_22_b_22;
  assign f_u_arrmul24_fa11_22_f_u_arrmul24_and11_22_y0 = f_u_arrmul24_and11_22_y0;
  assign f_u_arrmul24_fa11_22_f_u_arrmul24_fa12_21_y2 = f_u_arrmul24_fa12_21_y2;
  assign f_u_arrmul24_fa11_22_f_u_arrmul24_fa10_22_y4 = f_u_arrmul24_fa10_22_y4;
  assign f_u_arrmul24_fa11_22_y0 = f_u_arrmul24_fa11_22_f_u_arrmul24_and11_22_y0 ^ f_u_arrmul24_fa11_22_f_u_arrmul24_fa12_21_y2;
  assign f_u_arrmul24_fa11_22_y1 = f_u_arrmul24_fa11_22_f_u_arrmul24_and11_22_y0 & f_u_arrmul24_fa11_22_f_u_arrmul24_fa12_21_y2;
  assign f_u_arrmul24_fa11_22_y2 = f_u_arrmul24_fa11_22_y0 ^ f_u_arrmul24_fa11_22_f_u_arrmul24_fa10_22_y4;
  assign f_u_arrmul24_fa11_22_y3 = f_u_arrmul24_fa11_22_y0 & f_u_arrmul24_fa11_22_f_u_arrmul24_fa10_22_y4;
  assign f_u_arrmul24_fa11_22_y4 = f_u_arrmul24_fa11_22_y1 | f_u_arrmul24_fa11_22_y3;
  assign f_u_arrmul24_and12_22_a_12 = a_12;
  assign f_u_arrmul24_and12_22_b_22 = b_22;
  assign f_u_arrmul24_and12_22_y0 = f_u_arrmul24_and12_22_a_12 & f_u_arrmul24_and12_22_b_22;
  assign f_u_arrmul24_fa12_22_f_u_arrmul24_and12_22_y0 = f_u_arrmul24_and12_22_y0;
  assign f_u_arrmul24_fa12_22_f_u_arrmul24_fa13_21_y2 = f_u_arrmul24_fa13_21_y2;
  assign f_u_arrmul24_fa12_22_f_u_arrmul24_fa11_22_y4 = f_u_arrmul24_fa11_22_y4;
  assign f_u_arrmul24_fa12_22_y0 = f_u_arrmul24_fa12_22_f_u_arrmul24_and12_22_y0 ^ f_u_arrmul24_fa12_22_f_u_arrmul24_fa13_21_y2;
  assign f_u_arrmul24_fa12_22_y1 = f_u_arrmul24_fa12_22_f_u_arrmul24_and12_22_y0 & f_u_arrmul24_fa12_22_f_u_arrmul24_fa13_21_y2;
  assign f_u_arrmul24_fa12_22_y2 = f_u_arrmul24_fa12_22_y0 ^ f_u_arrmul24_fa12_22_f_u_arrmul24_fa11_22_y4;
  assign f_u_arrmul24_fa12_22_y3 = f_u_arrmul24_fa12_22_y0 & f_u_arrmul24_fa12_22_f_u_arrmul24_fa11_22_y4;
  assign f_u_arrmul24_fa12_22_y4 = f_u_arrmul24_fa12_22_y1 | f_u_arrmul24_fa12_22_y3;
  assign f_u_arrmul24_and13_22_a_13 = a_13;
  assign f_u_arrmul24_and13_22_b_22 = b_22;
  assign f_u_arrmul24_and13_22_y0 = f_u_arrmul24_and13_22_a_13 & f_u_arrmul24_and13_22_b_22;
  assign f_u_arrmul24_fa13_22_f_u_arrmul24_and13_22_y0 = f_u_arrmul24_and13_22_y0;
  assign f_u_arrmul24_fa13_22_f_u_arrmul24_fa14_21_y2 = f_u_arrmul24_fa14_21_y2;
  assign f_u_arrmul24_fa13_22_f_u_arrmul24_fa12_22_y4 = f_u_arrmul24_fa12_22_y4;
  assign f_u_arrmul24_fa13_22_y0 = f_u_arrmul24_fa13_22_f_u_arrmul24_and13_22_y0 ^ f_u_arrmul24_fa13_22_f_u_arrmul24_fa14_21_y2;
  assign f_u_arrmul24_fa13_22_y1 = f_u_arrmul24_fa13_22_f_u_arrmul24_and13_22_y0 & f_u_arrmul24_fa13_22_f_u_arrmul24_fa14_21_y2;
  assign f_u_arrmul24_fa13_22_y2 = f_u_arrmul24_fa13_22_y0 ^ f_u_arrmul24_fa13_22_f_u_arrmul24_fa12_22_y4;
  assign f_u_arrmul24_fa13_22_y3 = f_u_arrmul24_fa13_22_y0 & f_u_arrmul24_fa13_22_f_u_arrmul24_fa12_22_y4;
  assign f_u_arrmul24_fa13_22_y4 = f_u_arrmul24_fa13_22_y1 | f_u_arrmul24_fa13_22_y3;
  assign f_u_arrmul24_and14_22_a_14 = a_14;
  assign f_u_arrmul24_and14_22_b_22 = b_22;
  assign f_u_arrmul24_and14_22_y0 = f_u_arrmul24_and14_22_a_14 & f_u_arrmul24_and14_22_b_22;
  assign f_u_arrmul24_fa14_22_f_u_arrmul24_and14_22_y0 = f_u_arrmul24_and14_22_y0;
  assign f_u_arrmul24_fa14_22_f_u_arrmul24_fa15_21_y2 = f_u_arrmul24_fa15_21_y2;
  assign f_u_arrmul24_fa14_22_f_u_arrmul24_fa13_22_y4 = f_u_arrmul24_fa13_22_y4;
  assign f_u_arrmul24_fa14_22_y0 = f_u_arrmul24_fa14_22_f_u_arrmul24_and14_22_y0 ^ f_u_arrmul24_fa14_22_f_u_arrmul24_fa15_21_y2;
  assign f_u_arrmul24_fa14_22_y1 = f_u_arrmul24_fa14_22_f_u_arrmul24_and14_22_y0 & f_u_arrmul24_fa14_22_f_u_arrmul24_fa15_21_y2;
  assign f_u_arrmul24_fa14_22_y2 = f_u_arrmul24_fa14_22_y0 ^ f_u_arrmul24_fa14_22_f_u_arrmul24_fa13_22_y4;
  assign f_u_arrmul24_fa14_22_y3 = f_u_arrmul24_fa14_22_y0 & f_u_arrmul24_fa14_22_f_u_arrmul24_fa13_22_y4;
  assign f_u_arrmul24_fa14_22_y4 = f_u_arrmul24_fa14_22_y1 | f_u_arrmul24_fa14_22_y3;
  assign f_u_arrmul24_and15_22_a_15 = a_15;
  assign f_u_arrmul24_and15_22_b_22 = b_22;
  assign f_u_arrmul24_and15_22_y0 = f_u_arrmul24_and15_22_a_15 & f_u_arrmul24_and15_22_b_22;
  assign f_u_arrmul24_fa15_22_f_u_arrmul24_and15_22_y0 = f_u_arrmul24_and15_22_y0;
  assign f_u_arrmul24_fa15_22_f_u_arrmul24_fa16_21_y2 = f_u_arrmul24_fa16_21_y2;
  assign f_u_arrmul24_fa15_22_f_u_arrmul24_fa14_22_y4 = f_u_arrmul24_fa14_22_y4;
  assign f_u_arrmul24_fa15_22_y0 = f_u_arrmul24_fa15_22_f_u_arrmul24_and15_22_y0 ^ f_u_arrmul24_fa15_22_f_u_arrmul24_fa16_21_y2;
  assign f_u_arrmul24_fa15_22_y1 = f_u_arrmul24_fa15_22_f_u_arrmul24_and15_22_y0 & f_u_arrmul24_fa15_22_f_u_arrmul24_fa16_21_y2;
  assign f_u_arrmul24_fa15_22_y2 = f_u_arrmul24_fa15_22_y0 ^ f_u_arrmul24_fa15_22_f_u_arrmul24_fa14_22_y4;
  assign f_u_arrmul24_fa15_22_y3 = f_u_arrmul24_fa15_22_y0 & f_u_arrmul24_fa15_22_f_u_arrmul24_fa14_22_y4;
  assign f_u_arrmul24_fa15_22_y4 = f_u_arrmul24_fa15_22_y1 | f_u_arrmul24_fa15_22_y3;
  assign f_u_arrmul24_and16_22_a_16 = a_16;
  assign f_u_arrmul24_and16_22_b_22 = b_22;
  assign f_u_arrmul24_and16_22_y0 = f_u_arrmul24_and16_22_a_16 & f_u_arrmul24_and16_22_b_22;
  assign f_u_arrmul24_fa16_22_f_u_arrmul24_and16_22_y0 = f_u_arrmul24_and16_22_y0;
  assign f_u_arrmul24_fa16_22_f_u_arrmul24_fa17_21_y2 = f_u_arrmul24_fa17_21_y2;
  assign f_u_arrmul24_fa16_22_f_u_arrmul24_fa15_22_y4 = f_u_arrmul24_fa15_22_y4;
  assign f_u_arrmul24_fa16_22_y0 = f_u_arrmul24_fa16_22_f_u_arrmul24_and16_22_y0 ^ f_u_arrmul24_fa16_22_f_u_arrmul24_fa17_21_y2;
  assign f_u_arrmul24_fa16_22_y1 = f_u_arrmul24_fa16_22_f_u_arrmul24_and16_22_y0 & f_u_arrmul24_fa16_22_f_u_arrmul24_fa17_21_y2;
  assign f_u_arrmul24_fa16_22_y2 = f_u_arrmul24_fa16_22_y0 ^ f_u_arrmul24_fa16_22_f_u_arrmul24_fa15_22_y4;
  assign f_u_arrmul24_fa16_22_y3 = f_u_arrmul24_fa16_22_y0 & f_u_arrmul24_fa16_22_f_u_arrmul24_fa15_22_y4;
  assign f_u_arrmul24_fa16_22_y4 = f_u_arrmul24_fa16_22_y1 | f_u_arrmul24_fa16_22_y3;
  assign f_u_arrmul24_and17_22_a_17 = a_17;
  assign f_u_arrmul24_and17_22_b_22 = b_22;
  assign f_u_arrmul24_and17_22_y0 = f_u_arrmul24_and17_22_a_17 & f_u_arrmul24_and17_22_b_22;
  assign f_u_arrmul24_fa17_22_f_u_arrmul24_and17_22_y0 = f_u_arrmul24_and17_22_y0;
  assign f_u_arrmul24_fa17_22_f_u_arrmul24_fa18_21_y2 = f_u_arrmul24_fa18_21_y2;
  assign f_u_arrmul24_fa17_22_f_u_arrmul24_fa16_22_y4 = f_u_arrmul24_fa16_22_y4;
  assign f_u_arrmul24_fa17_22_y0 = f_u_arrmul24_fa17_22_f_u_arrmul24_and17_22_y0 ^ f_u_arrmul24_fa17_22_f_u_arrmul24_fa18_21_y2;
  assign f_u_arrmul24_fa17_22_y1 = f_u_arrmul24_fa17_22_f_u_arrmul24_and17_22_y0 & f_u_arrmul24_fa17_22_f_u_arrmul24_fa18_21_y2;
  assign f_u_arrmul24_fa17_22_y2 = f_u_arrmul24_fa17_22_y0 ^ f_u_arrmul24_fa17_22_f_u_arrmul24_fa16_22_y4;
  assign f_u_arrmul24_fa17_22_y3 = f_u_arrmul24_fa17_22_y0 & f_u_arrmul24_fa17_22_f_u_arrmul24_fa16_22_y4;
  assign f_u_arrmul24_fa17_22_y4 = f_u_arrmul24_fa17_22_y1 | f_u_arrmul24_fa17_22_y3;
  assign f_u_arrmul24_and18_22_a_18 = a_18;
  assign f_u_arrmul24_and18_22_b_22 = b_22;
  assign f_u_arrmul24_and18_22_y0 = f_u_arrmul24_and18_22_a_18 & f_u_arrmul24_and18_22_b_22;
  assign f_u_arrmul24_fa18_22_f_u_arrmul24_and18_22_y0 = f_u_arrmul24_and18_22_y0;
  assign f_u_arrmul24_fa18_22_f_u_arrmul24_fa19_21_y2 = f_u_arrmul24_fa19_21_y2;
  assign f_u_arrmul24_fa18_22_f_u_arrmul24_fa17_22_y4 = f_u_arrmul24_fa17_22_y4;
  assign f_u_arrmul24_fa18_22_y0 = f_u_arrmul24_fa18_22_f_u_arrmul24_and18_22_y0 ^ f_u_arrmul24_fa18_22_f_u_arrmul24_fa19_21_y2;
  assign f_u_arrmul24_fa18_22_y1 = f_u_arrmul24_fa18_22_f_u_arrmul24_and18_22_y0 & f_u_arrmul24_fa18_22_f_u_arrmul24_fa19_21_y2;
  assign f_u_arrmul24_fa18_22_y2 = f_u_arrmul24_fa18_22_y0 ^ f_u_arrmul24_fa18_22_f_u_arrmul24_fa17_22_y4;
  assign f_u_arrmul24_fa18_22_y3 = f_u_arrmul24_fa18_22_y0 & f_u_arrmul24_fa18_22_f_u_arrmul24_fa17_22_y4;
  assign f_u_arrmul24_fa18_22_y4 = f_u_arrmul24_fa18_22_y1 | f_u_arrmul24_fa18_22_y3;
  assign f_u_arrmul24_and19_22_a_19 = a_19;
  assign f_u_arrmul24_and19_22_b_22 = b_22;
  assign f_u_arrmul24_and19_22_y0 = f_u_arrmul24_and19_22_a_19 & f_u_arrmul24_and19_22_b_22;
  assign f_u_arrmul24_fa19_22_f_u_arrmul24_and19_22_y0 = f_u_arrmul24_and19_22_y0;
  assign f_u_arrmul24_fa19_22_f_u_arrmul24_fa20_21_y2 = f_u_arrmul24_fa20_21_y2;
  assign f_u_arrmul24_fa19_22_f_u_arrmul24_fa18_22_y4 = f_u_arrmul24_fa18_22_y4;
  assign f_u_arrmul24_fa19_22_y0 = f_u_arrmul24_fa19_22_f_u_arrmul24_and19_22_y0 ^ f_u_arrmul24_fa19_22_f_u_arrmul24_fa20_21_y2;
  assign f_u_arrmul24_fa19_22_y1 = f_u_arrmul24_fa19_22_f_u_arrmul24_and19_22_y0 & f_u_arrmul24_fa19_22_f_u_arrmul24_fa20_21_y2;
  assign f_u_arrmul24_fa19_22_y2 = f_u_arrmul24_fa19_22_y0 ^ f_u_arrmul24_fa19_22_f_u_arrmul24_fa18_22_y4;
  assign f_u_arrmul24_fa19_22_y3 = f_u_arrmul24_fa19_22_y0 & f_u_arrmul24_fa19_22_f_u_arrmul24_fa18_22_y4;
  assign f_u_arrmul24_fa19_22_y4 = f_u_arrmul24_fa19_22_y1 | f_u_arrmul24_fa19_22_y3;
  assign f_u_arrmul24_and20_22_a_20 = a_20;
  assign f_u_arrmul24_and20_22_b_22 = b_22;
  assign f_u_arrmul24_and20_22_y0 = f_u_arrmul24_and20_22_a_20 & f_u_arrmul24_and20_22_b_22;
  assign f_u_arrmul24_fa20_22_f_u_arrmul24_and20_22_y0 = f_u_arrmul24_and20_22_y0;
  assign f_u_arrmul24_fa20_22_f_u_arrmul24_fa21_21_y2 = f_u_arrmul24_fa21_21_y2;
  assign f_u_arrmul24_fa20_22_f_u_arrmul24_fa19_22_y4 = f_u_arrmul24_fa19_22_y4;
  assign f_u_arrmul24_fa20_22_y0 = f_u_arrmul24_fa20_22_f_u_arrmul24_and20_22_y0 ^ f_u_arrmul24_fa20_22_f_u_arrmul24_fa21_21_y2;
  assign f_u_arrmul24_fa20_22_y1 = f_u_arrmul24_fa20_22_f_u_arrmul24_and20_22_y0 & f_u_arrmul24_fa20_22_f_u_arrmul24_fa21_21_y2;
  assign f_u_arrmul24_fa20_22_y2 = f_u_arrmul24_fa20_22_y0 ^ f_u_arrmul24_fa20_22_f_u_arrmul24_fa19_22_y4;
  assign f_u_arrmul24_fa20_22_y3 = f_u_arrmul24_fa20_22_y0 & f_u_arrmul24_fa20_22_f_u_arrmul24_fa19_22_y4;
  assign f_u_arrmul24_fa20_22_y4 = f_u_arrmul24_fa20_22_y1 | f_u_arrmul24_fa20_22_y3;
  assign f_u_arrmul24_and21_22_a_21 = a_21;
  assign f_u_arrmul24_and21_22_b_22 = b_22;
  assign f_u_arrmul24_and21_22_y0 = f_u_arrmul24_and21_22_a_21 & f_u_arrmul24_and21_22_b_22;
  assign f_u_arrmul24_fa21_22_f_u_arrmul24_and21_22_y0 = f_u_arrmul24_and21_22_y0;
  assign f_u_arrmul24_fa21_22_f_u_arrmul24_fa22_21_y2 = f_u_arrmul24_fa22_21_y2;
  assign f_u_arrmul24_fa21_22_f_u_arrmul24_fa20_22_y4 = f_u_arrmul24_fa20_22_y4;
  assign f_u_arrmul24_fa21_22_y0 = f_u_arrmul24_fa21_22_f_u_arrmul24_and21_22_y0 ^ f_u_arrmul24_fa21_22_f_u_arrmul24_fa22_21_y2;
  assign f_u_arrmul24_fa21_22_y1 = f_u_arrmul24_fa21_22_f_u_arrmul24_and21_22_y0 & f_u_arrmul24_fa21_22_f_u_arrmul24_fa22_21_y2;
  assign f_u_arrmul24_fa21_22_y2 = f_u_arrmul24_fa21_22_y0 ^ f_u_arrmul24_fa21_22_f_u_arrmul24_fa20_22_y4;
  assign f_u_arrmul24_fa21_22_y3 = f_u_arrmul24_fa21_22_y0 & f_u_arrmul24_fa21_22_f_u_arrmul24_fa20_22_y4;
  assign f_u_arrmul24_fa21_22_y4 = f_u_arrmul24_fa21_22_y1 | f_u_arrmul24_fa21_22_y3;
  assign f_u_arrmul24_and22_22_a_22 = a_22;
  assign f_u_arrmul24_and22_22_b_22 = b_22;
  assign f_u_arrmul24_and22_22_y0 = f_u_arrmul24_and22_22_a_22 & f_u_arrmul24_and22_22_b_22;
  assign f_u_arrmul24_fa22_22_f_u_arrmul24_and22_22_y0 = f_u_arrmul24_and22_22_y0;
  assign f_u_arrmul24_fa22_22_f_u_arrmul24_fa23_21_y2 = f_u_arrmul24_fa23_21_y2;
  assign f_u_arrmul24_fa22_22_f_u_arrmul24_fa21_22_y4 = f_u_arrmul24_fa21_22_y4;
  assign f_u_arrmul24_fa22_22_y0 = f_u_arrmul24_fa22_22_f_u_arrmul24_and22_22_y0 ^ f_u_arrmul24_fa22_22_f_u_arrmul24_fa23_21_y2;
  assign f_u_arrmul24_fa22_22_y1 = f_u_arrmul24_fa22_22_f_u_arrmul24_and22_22_y0 & f_u_arrmul24_fa22_22_f_u_arrmul24_fa23_21_y2;
  assign f_u_arrmul24_fa22_22_y2 = f_u_arrmul24_fa22_22_y0 ^ f_u_arrmul24_fa22_22_f_u_arrmul24_fa21_22_y4;
  assign f_u_arrmul24_fa22_22_y3 = f_u_arrmul24_fa22_22_y0 & f_u_arrmul24_fa22_22_f_u_arrmul24_fa21_22_y4;
  assign f_u_arrmul24_fa22_22_y4 = f_u_arrmul24_fa22_22_y1 | f_u_arrmul24_fa22_22_y3;
  assign f_u_arrmul24_and23_22_a_23 = a_23;
  assign f_u_arrmul24_and23_22_b_22 = b_22;
  assign f_u_arrmul24_and23_22_y0 = f_u_arrmul24_and23_22_a_23 & f_u_arrmul24_and23_22_b_22;
  assign f_u_arrmul24_fa23_22_f_u_arrmul24_and23_22_y0 = f_u_arrmul24_and23_22_y0;
  assign f_u_arrmul24_fa23_22_f_u_arrmul24_fa23_21_y4 = f_u_arrmul24_fa23_21_y4;
  assign f_u_arrmul24_fa23_22_f_u_arrmul24_fa22_22_y4 = f_u_arrmul24_fa22_22_y4;
  assign f_u_arrmul24_fa23_22_y0 = f_u_arrmul24_fa23_22_f_u_arrmul24_and23_22_y0 ^ f_u_arrmul24_fa23_22_f_u_arrmul24_fa23_21_y4;
  assign f_u_arrmul24_fa23_22_y1 = f_u_arrmul24_fa23_22_f_u_arrmul24_and23_22_y0 & f_u_arrmul24_fa23_22_f_u_arrmul24_fa23_21_y4;
  assign f_u_arrmul24_fa23_22_y2 = f_u_arrmul24_fa23_22_y0 ^ f_u_arrmul24_fa23_22_f_u_arrmul24_fa22_22_y4;
  assign f_u_arrmul24_fa23_22_y3 = f_u_arrmul24_fa23_22_y0 & f_u_arrmul24_fa23_22_f_u_arrmul24_fa22_22_y4;
  assign f_u_arrmul24_fa23_22_y4 = f_u_arrmul24_fa23_22_y1 | f_u_arrmul24_fa23_22_y3;
  assign f_u_arrmul24_and0_23_a_0 = a_0;
  assign f_u_arrmul24_and0_23_b_23 = b_23;
  assign f_u_arrmul24_and0_23_y0 = f_u_arrmul24_and0_23_a_0 & f_u_arrmul24_and0_23_b_23;
  assign f_u_arrmul24_ha0_23_f_u_arrmul24_and0_23_y0 = f_u_arrmul24_and0_23_y0;
  assign f_u_arrmul24_ha0_23_f_u_arrmul24_fa1_22_y2 = f_u_arrmul24_fa1_22_y2;
  assign f_u_arrmul24_ha0_23_y0 = f_u_arrmul24_ha0_23_f_u_arrmul24_and0_23_y0 ^ f_u_arrmul24_ha0_23_f_u_arrmul24_fa1_22_y2;
  assign f_u_arrmul24_ha0_23_y1 = f_u_arrmul24_ha0_23_f_u_arrmul24_and0_23_y0 & f_u_arrmul24_ha0_23_f_u_arrmul24_fa1_22_y2;
  assign f_u_arrmul24_and1_23_a_1 = a_1;
  assign f_u_arrmul24_and1_23_b_23 = b_23;
  assign f_u_arrmul24_and1_23_y0 = f_u_arrmul24_and1_23_a_1 & f_u_arrmul24_and1_23_b_23;
  assign f_u_arrmul24_fa1_23_f_u_arrmul24_and1_23_y0 = f_u_arrmul24_and1_23_y0;
  assign f_u_arrmul24_fa1_23_f_u_arrmul24_fa2_22_y2 = f_u_arrmul24_fa2_22_y2;
  assign f_u_arrmul24_fa1_23_f_u_arrmul24_ha0_23_y1 = f_u_arrmul24_ha0_23_y1;
  assign f_u_arrmul24_fa1_23_y0 = f_u_arrmul24_fa1_23_f_u_arrmul24_and1_23_y0 ^ f_u_arrmul24_fa1_23_f_u_arrmul24_fa2_22_y2;
  assign f_u_arrmul24_fa1_23_y1 = f_u_arrmul24_fa1_23_f_u_arrmul24_and1_23_y0 & f_u_arrmul24_fa1_23_f_u_arrmul24_fa2_22_y2;
  assign f_u_arrmul24_fa1_23_y2 = f_u_arrmul24_fa1_23_y0 ^ f_u_arrmul24_fa1_23_f_u_arrmul24_ha0_23_y1;
  assign f_u_arrmul24_fa1_23_y3 = f_u_arrmul24_fa1_23_y0 & f_u_arrmul24_fa1_23_f_u_arrmul24_ha0_23_y1;
  assign f_u_arrmul24_fa1_23_y4 = f_u_arrmul24_fa1_23_y1 | f_u_arrmul24_fa1_23_y3;
  assign f_u_arrmul24_and2_23_a_2 = a_2;
  assign f_u_arrmul24_and2_23_b_23 = b_23;
  assign f_u_arrmul24_and2_23_y0 = f_u_arrmul24_and2_23_a_2 & f_u_arrmul24_and2_23_b_23;
  assign f_u_arrmul24_fa2_23_f_u_arrmul24_and2_23_y0 = f_u_arrmul24_and2_23_y0;
  assign f_u_arrmul24_fa2_23_f_u_arrmul24_fa3_22_y2 = f_u_arrmul24_fa3_22_y2;
  assign f_u_arrmul24_fa2_23_f_u_arrmul24_fa1_23_y4 = f_u_arrmul24_fa1_23_y4;
  assign f_u_arrmul24_fa2_23_y0 = f_u_arrmul24_fa2_23_f_u_arrmul24_and2_23_y0 ^ f_u_arrmul24_fa2_23_f_u_arrmul24_fa3_22_y2;
  assign f_u_arrmul24_fa2_23_y1 = f_u_arrmul24_fa2_23_f_u_arrmul24_and2_23_y0 & f_u_arrmul24_fa2_23_f_u_arrmul24_fa3_22_y2;
  assign f_u_arrmul24_fa2_23_y2 = f_u_arrmul24_fa2_23_y0 ^ f_u_arrmul24_fa2_23_f_u_arrmul24_fa1_23_y4;
  assign f_u_arrmul24_fa2_23_y3 = f_u_arrmul24_fa2_23_y0 & f_u_arrmul24_fa2_23_f_u_arrmul24_fa1_23_y4;
  assign f_u_arrmul24_fa2_23_y4 = f_u_arrmul24_fa2_23_y1 | f_u_arrmul24_fa2_23_y3;
  assign f_u_arrmul24_and3_23_a_3 = a_3;
  assign f_u_arrmul24_and3_23_b_23 = b_23;
  assign f_u_arrmul24_and3_23_y0 = f_u_arrmul24_and3_23_a_3 & f_u_arrmul24_and3_23_b_23;
  assign f_u_arrmul24_fa3_23_f_u_arrmul24_and3_23_y0 = f_u_arrmul24_and3_23_y0;
  assign f_u_arrmul24_fa3_23_f_u_arrmul24_fa4_22_y2 = f_u_arrmul24_fa4_22_y2;
  assign f_u_arrmul24_fa3_23_f_u_arrmul24_fa2_23_y4 = f_u_arrmul24_fa2_23_y4;
  assign f_u_arrmul24_fa3_23_y0 = f_u_arrmul24_fa3_23_f_u_arrmul24_and3_23_y0 ^ f_u_arrmul24_fa3_23_f_u_arrmul24_fa4_22_y2;
  assign f_u_arrmul24_fa3_23_y1 = f_u_arrmul24_fa3_23_f_u_arrmul24_and3_23_y0 & f_u_arrmul24_fa3_23_f_u_arrmul24_fa4_22_y2;
  assign f_u_arrmul24_fa3_23_y2 = f_u_arrmul24_fa3_23_y0 ^ f_u_arrmul24_fa3_23_f_u_arrmul24_fa2_23_y4;
  assign f_u_arrmul24_fa3_23_y3 = f_u_arrmul24_fa3_23_y0 & f_u_arrmul24_fa3_23_f_u_arrmul24_fa2_23_y4;
  assign f_u_arrmul24_fa3_23_y4 = f_u_arrmul24_fa3_23_y1 | f_u_arrmul24_fa3_23_y3;
  assign f_u_arrmul24_and4_23_a_4 = a_4;
  assign f_u_arrmul24_and4_23_b_23 = b_23;
  assign f_u_arrmul24_and4_23_y0 = f_u_arrmul24_and4_23_a_4 & f_u_arrmul24_and4_23_b_23;
  assign f_u_arrmul24_fa4_23_f_u_arrmul24_and4_23_y0 = f_u_arrmul24_and4_23_y0;
  assign f_u_arrmul24_fa4_23_f_u_arrmul24_fa5_22_y2 = f_u_arrmul24_fa5_22_y2;
  assign f_u_arrmul24_fa4_23_f_u_arrmul24_fa3_23_y4 = f_u_arrmul24_fa3_23_y4;
  assign f_u_arrmul24_fa4_23_y0 = f_u_arrmul24_fa4_23_f_u_arrmul24_and4_23_y0 ^ f_u_arrmul24_fa4_23_f_u_arrmul24_fa5_22_y2;
  assign f_u_arrmul24_fa4_23_y1 = f_u_arrmul24_fa4_23_f_u_arrmul24_and4_23_y0 & f_u_arrmul24_fa4_23_f_u_arrmul24_fa5_22_y2;
  assign f_u_arrmul24_fa4_23_y2 = f_u_arrmul24_fa4_23_y0 ^ f_u_arrmul24_fa4_23_f_u_arrmul24_fa3_23_y4;
  assign f_u_arrmul24_fa4_23_y3 = f_u_arrmul24_fa4_23_y0 & f_u_arrmul24_fa4_23_f_u_arrmul24_fa3_23_y4;
  assign f_u_arrmul24_fa4_23_y4 = f_u_arrmul24_fa4_23_y1 | f_u_arrmul24_fa4_23_y3;
  assign f_u_arrmul24_and5_23_a_5 = a_5;
  assign f_u_arrmul24_and5_23_b_23 = b_23;
  assign f_u_arrmul24_and5_23_y0 = f_u_arrmul24_and5_23_a_5 & f_u_arrmul24_and5_23_b_23;
  assign f_u_arrmul24_fa5_23_f_u_arrmul24_and5_23_y0 = f_u_arrmul24_and5_23_y0;
  assign f_u_arrmul24_fa5_23_f_u_arrmul24_fa6_22_y2 = f_u_arrmul24_fa6_22_y2;
  assign f_u_arrmul24_fa5_23_f_u_arrmul24_fa4_23_y4 = f_u_arrmul24_fa4_23_y4;
  assign f_u_arrmul24_fa5_23_y0 = f_u_arrmul24_fa5_23_f_u_arrmul24_and5_23_y0 ^ f_u_arrmul24_fa5_23_f_u_arrmul24_fa6_22_y2;
  assign f_u_arrmul24_fa5_23_y1 = f_u_arrmul24_fa5_23_f_u_arrmul24_and5_23_y0 & f_u_arrmul24_fa5_23_f_u_arrmul24_fa6_22_y2;
  assign f_u_arrmul24_fa5_23_y2 = f_u_arrmul24_fa5_23_y0 ^ f_u_arrmul24_fa5_23_f_u_arrmul24_fa4_23_y4;
  assign f_u_arrmul24_fa5_23_y3 = f_u_arrmul24_fa5_23_y0 & f_u_arrmul24_fa5_23_f_u_arrmul24_fa4_23_y4;
  assign f_u_arrmul24_fa5_23_y4 = f_u_arrmul24_fa5_23_y1 | f_u_arrmul24_fa5_23_y3;
  assign f_u_arrmul24_and6_23_a_6 = a_6;
  assign f_u_arrmul24_and6_23_b_23 = b_23;
  assign f_u_arrmul24_and6_23_y0 = f_u_arrmul24_and6_23_a_6 & f_u_arrmul24_and6_23_b_23;
  assign f_u_arrmul24_fa6_23_f_u_arrmul24_and6_23_y0 = f_u_arrmul24_and6_23_y0;
  assign f_u_arrmul24_fa6_23_f_u_arrmul24_fa7_22_y2 = f_u_arrmul24_fa7_22_y2;
  assign f_u_arrmul24_fa6_23_f_u_arrmul24_fa5_23_y4 = f_u_arrmul24_fa5_23_y4;
  assign f_u_arrmul24_fa6_23_y0 = f_u_arrmul24_fa6_23_f_u_arrmul24_and6_23_y0 ^ f_u_arrmul24_fa6_23_f_u_arrmul24_fa7_22_y2;
  assign f_u_arrmul24_fa6_23_y1 = f_u_arrmul24_fa6_23_f_u_arrmul24_and6_23_y0 & f_u_arrmul24_fa6_23_f_u_arrmul24_fa7_22_y2;
  assign f_u_arrmul24_fa6_23_y2 = f_u_arrmul24_fa6_23_y0 ^ f_u_arrmul24_fa6_23_f_u_arrmul24_fa5_23_y4;
  assign f_u_arrmul24_fa6_23_y3 = f_u_arrmul24_fa6_23_y0 & f_u_arrmul24_fa6_23_f_u_arrmul24_fa5_23_y4;
  assign f_u_arrmul24_fa6_23_y4 = f_u_arrmul24_fa6_23_y1 | f_u_arrmul24_fa6_23_y3;
  assign f_u_arrmul24_and7_23_a_7 = a_7;
  assign f_u_arrmul24_and7_23_b_23 = b_23;
  assign f_u_arrmul24_and7_23_y0 = f_u_arrmul24_and7_23_a_7 & f_u_arrmul24_and7_23_b_23;
  assign f_u_arrmul24_fa7_23_f_u_arrmul24_and7_23_y0 = f_u_arrmul24_and7_23_y0;
  assign f_u_arrmul24_fa7_23_f_u_arrmul24_fa8_22_y2 = f_u_arrmul24_fa8_22_y2;
  assign f_u_arrmul24_fa7_23_f_u_arrmul24_fa6_23_y4 = f_u_arrmul24_fa6_23_y4;
  assign f_u_arrmul24_fa7_23_y0 = f_u_arrmul24_fa7_23_f_u_arrmul24_and7_23_y0 ^ f_u_arrmul24_fa7_23_f_u_arrmul24_fa8_22_y2;
  assign f_u_arrmul24_fa7_23_y1 = f_u_arrmul24_fa7_23_f_u_arrmul24_and7_23_y0 & f_u_arrmul24_fa7_23_f_u_arrmul24_fa8_22_y2;
  assign f_u_arrmul24_fa7_23_y2 = f_u_arrmul24_fa7_23_y0 ^ f_u_arrmul24_fa7_23_f_u_arrmul24_fa6_23_y4;
  assign f_u_arrmul24_fa7_23_y3 = f_u_arrmul24_fa7_23_y0 & f_u_arrmul24_fa7_23_f_u_arrmul24_fa6_23_y4;
  assign f_u_arrmul24_fa7_23_y4 = f_u_arrmul24_fa7_23_y1 | f_u_arrmul24_fa7_23_y3;
  assign f_u_arrmul24_and8_23_a_8 = a_8;
  assign f_u_arrmul24_and8_23_b_23 = b_23;
  assign f_u_arrmul24_and8_23_y0 = f_u_arrmul24_and8_23_a_8 & f_u_arrmul24_and8_23_b_23;
  assign f_u_arrmul24_fa8_23_f_u_arrmul24_and8_23_y0 = f_u_arrmul24_and8_23_y0;
  assign f_u_arrmul24_fa8_23_f_u_arrmul24_fa9_22_y2 = f_u_arrmul24_fa9_22_y2;
  assign f_u_arrmul24_fa8_23_f_u_arrmul24_fa7_23_y4 = f_u_arrmul24_fa7_23_y4;
  assign f_u_arrmul24_fa8_23_y0 = f_u_arrmul24_fa8_23_f_u_arrmul24_and8_23_y0 ^ f_u_arrmul24_fa8_23_f_u_arrmul24_fa9_22_y2;
  assign f_u_arrmul24_fa8_23_y1 = f_u_arrmul24_fa8_23_f_u_arrmul24_and8_23_y0 & f_u_arrmul24_fa8_23_f_u_arrmul24_fa9_22_y2;
  assign f_u_arrmul24_fa8_23_y2 = f_u_arrmul24_fa8_23_y0 ^ f_u_arrmul24_fa8_23_f_u_arrmul24_fa7_23_y4;
  assign f_u_arrmul24_fa8_23_y3 = f_u_arrmul24_fa8_23_y0 & f_u_arrmul24_fa8_23_f_u_arrmul24_fa7_23_y4;
  assign f_u_arrmul24_fa8_23_y4 = f_u_arrmul24_fa8_23_y1 | f_u_arrmul24_fa8_23_y3;
  assign f_u_arrmul24_and9_23_a_9 = a_9;
  assign f_u_arrmul24_and9_23_b_23 = b_23;
  assign f_u_arrmul24_and9_23_y0 = f_u_arrmul24_and9_23_a_9 & f_u_arrmul24_and9_23_b_23;
  assign f_u_arrmul24_fa9_23_f_u_arrmul24_and9_23_y0 = f_u_arrmul24_and9_23_y0;
  assign f_u_arrmul24_fa9_23_f_u_arrmul24_fa10_22_y2 = f_u_arrmul24_fa10_22_y2;
  assign f_u_arrmul24_fa9_23_f_u_arrmul24_fa8_23_y4 = f_u_arrmul24_fa8_23_y4;
  assign f_u_arrmul24_fa9_23_y0 = f_u_arrmul24_fa9_23_f_u_arrmul24_and9_23_y0 ^ f_u_arrmul24_fa9_23_f_u_arrmul24_fa10_22_y2;
  assign f_u_arrmul24_fa9_23_y1 = f_u_arrmul24_fa9_23_f_u_arrmul24_and9_23_y0 & f_u_arrmul24_fa9_23_f_u_arrmul24_fa10_22_y2;
  assign f_u_arrmul24_fa9_23_y2 = f_u_arrmul24_fa9_23_y0 ^ f_u_arrmul24_fa9_23_f_u_arrmul24_fa8_23_y4;
  assign f_u_arrmul24_fa9_23_y3 = f_u_arrmul24_fa9_23_y0 & f_u_arrmul24_fa9_23_f_u_arrmul24_fa8_23_y4;
  assign f_u_arrmul24_fa9_23_y4 = f_u_arrmul24_fa9_23_y1 | f_u_arrmul24_fa9_23_y3;
  assign f_u_arrmul24_and10_23_a_10 = a_10;
  assign f_u_arrmul24_and10_23_b_23 = b_23;
  assign f_u_arrmul24_and10_23_y0 = f_u_arrmul24_and10_23_a_10 & f_u_arrmul24_and10_23_b_23;
  assign f_u_arrmul24_fa10_23_f_u_arrmul24_and10_23_y0 = f_u_arrmul24_and10_23_y0;
  assign f_u_arrmul24_fa10_23_f_u_arrmul24_fa11_22_y2 = f_u_arrmul24_fa11_22_y2;
  assign f_u_arrmul24_fa10_23_f_u_arrmul24_fa9_23_y4 = f_u_arrmul24_fa9_23_y4;
  assign f_u_arrmul24_fa10_23_y0 = f_u_arrmul24_fa10_23_f_u_arrmul24_and10_23_y0 ^ f_u_arrmul24_fa10_23_f_u_arrmul24_fa11_22_y2;
  assign f_u_arrmul24_fa10_23_y1 = f_u_arrmul24_fa10_23_f_u_arrmul24_and10_23_y0 & f_u_arrmul24_fa10_23_f_u_arrmul24_fa11_22_y2;
  assign f_u_arrmul24_fa10_23_y2 = f_u_arrmul24_fa10_23_y0 ^ f_u_arrmul24_fa10_23_f_u_arrmul24_fa9_23_y4;
  assign f_u_arrmul24_fa10_23_y3 = f_u_arrmul24_fa10_23_y0 & f_u_arrmul24_fa10_23_f_u_arrmul24_fa9_23_y4;
  assign f_u_arrmul24_fa10_23_y4 = f_u_arrmul24_fa10_23_y1 | f_u_arrmul24_fa10_23_y3;
  assign f_u_arrmul24_and11_23_a_11 = a_11;
  assign f_u_arrmul24_and11_23_b_23 = b_23;
  assign f_u_arrmul24_and11_23_y0 = f_u_arrmul24_and11_23_a_11 & f_u_arrmul24_and11_23_b_23;
  assign f_u_arrmul24_fa11_23_f_u_arrmul24_and11_23_y0 = f_u_arrmul24_and11_23_y0;
  assign f_u_arrmul24_fa11_23_f_u_arrmul24_fa12_22_y2 = f_u_arrmul24_fa12_22_y2;
  assign f_u_arrmul24_fa11_23_f_u_arrmul24_fa10_23_y4 = f_u_arrmul24_fa10_23_y4;
  assign f_u_arrmul24_fa11_23_y0 = f_u_arrmul24_fa11_23_f_u_arrmul24_and11_23_y0 ^ f_u_arrmul24_fa11_23_f_u_arrmul24_fa12_22_y2;
  assign f_u_arrmul24_fa11_23_y1 = f_u_arrmul24_fa11_23_f_u_arrmul24_and11_23_y0 & f_u_arrmul24_fa11_23_f_u_arrmul24_fa12_22_y2;
  assign f_u_arrmul24_fa11_23_y2 = f_u_arrmul24_fa11_23_y0 ^ f_u_arrmul24_fa11_23_f_u_arrmul24_fa10_23_y4;
  assign f_u_arrmul24_fa11_23_y3 = f_u_arrmul24_fa11_23_y0 & f_u_arrmul24_fa11_23_f_u_arrmul24_fa10_23_y4;
  assign f_u_arrmul24_fa11_23_y4 = f_u_arrmul24_fa11_23_y1 | f_u_arrmul24_fa11_23_y3;
  assign f_u_arrmul24_and12_23_a_12 = a_12;
  assign f_u_arrmul24_and12_23_b_23 = b_23;
  assign f_u_arrmul24_and12_23_y0 = f_u_arrmul24_and12_23_a_12 & f_u_arrmul24_and12_23_b_23;
  assign f_u_arrmul24_fa12_23_f_u_arrmul24_and12_23_y0 = f_u_arrmul24_and12_23_y0;
  assign f_u_arrmul24_fa12_23_f_u_arrmul24_fa13_22_y2 = f_u_arrmul24_fa13_22_y2;
  assign f_u_arrmul24_fa12_23_f_u_arrmul24_fa11_23_y4 = f_u_arrmul24_fa11_23_y4;
  assign f_u_arrmul24_fa12_23_y0 = f_u_arrmul24_fa12_23_f_u_arrmul24_and12_23_y0 ^ f_u_arrmul24_fa12_23_f_u_arrmul24_fa13_22_y2;
  assign f_u_arrmul24_fa12_23_y1 = f_u_arrmul24_fa12_23_f_u_arrmul24_and12_23_y0 & f_u_arrmul24_fa12_23_f_u_arrmul24_fa13_22_y2;
  assign f_u_arrmul24_fa12_23_y2 = f_u_arrmul24_fa12_23_y0 ^ f_u_arrmul24_fa12_23_f_u_arrmul24_fa11_23_y4;
  assign f_u_arrmul24_fa12_23_y3 = f_u_arrmul24_fa12_23_y0 & f_u_arrmul24_fa12_23_f_u_arrmul24_fa11_23_y4;
  assign f_u_arrmul24_fa12_23_y4 = f_u_arrmul24_fa12_23_y1 | f_u_arrmul24_fa12_23_y3;
  assign f_u_arrmul24_and13_23_a_13 = a_13;
  assign f_u_arrmul24_and13_23_b_23 = b_23;
  assign f_u_arrmul24_and13_23_y0 = f_u_arrmul24_and13_23_a_13 & f_u_arrmul24_and13_23_b_23;
  assign f_u_arrmul24_fa13_23_f_u_arrmul24_and13_23_y0 = f_u_arrmul24_and13_23_y0;
  assign f_u_arrmul24_fa13_23_f_u_arrmul24_fa14_22_y2 = f_u_arrmul24_fa14_22_y2;
  assign f_u_arrmul24_fa13_23_f_u_arrmul24_fa12_23_y4 = f_u_arrmul24_fa12_23_y4;
  assign f_u_arrmul24_fa13_23_y0 = f_u_arrmul24_fa13_23_f_u_arrmul24_and13_23_y0 ^ f_u_arrmul24_fa13_23_f_u_arrmul24_fa14_22_y2;
  assign f_u_arrmul24_fa13_23_y1 = f_u_arrmul24_fa13_23_f_u_arrmul24_and13_23_y0 & f_u_arrmul24_fa13_23_f_u_arrmul24_fa14_22_y2;
  assign f_u_arrmul24_fa13_23_y2 = f_u_arrmul24_fa13_23_y0 ^ f_u_arrmul24_fa13_23_f_u_arrmul24_fa12_23_y4;
  assign f_u_arrmul24_fa13_23_y3 = f_u_arrmul24_fa13_23_y0 & f_u_arrmul24_fa13_23_f_u_arrmul24_fa12_23_y4;
  assign f_u_arrmul24_fa13_23_y4 = f_u_arrmul24_fa13_23_y1 | f_u_arrmul24_fa13_23_y3;
  assign f_u_arrmul24_and14_23_a_14 = a_14;
  assign f_u_arrmul24_and14_23_b_23 = b_23;
  assign f_u_arrmul24_and14_23_y0 = f_u_arrmul24_and14_23_a_14 & f_u_arrmul24_and14_23_b_23;
  assign f_u_arrmul24_fa14_23_f_u_arrmul24_and14_23_y0 = f_u_arrmul24_and14_23_y0;
  assign f_u_arrmul24_fa14_23_f_u_arrmul24_fa15_22_y2 = f_u_arrmul24_fa15_22_y2;
  assign f_u_arrmul24_fa14_23_f_u_arrmul24_fa13_23_y4 = f_u_arrmul24_fa13_23_y4;
  assign f_u_arrmul24_fa14_23_y0 = f_u_arrmul24_fa14_23_f_u_arrmul24_and14_23_y0 ^ f_u_arrmul24_fa14_23_f_u_arrmul24_fa15_22_y2;
  assign f_u_arrmul24_fa14_23_y1 = f_u_arrmul24_fa14_23_f_u_arrmul24_and14_23_y0 & f_u_arrmul24_fa14_23_f_u_arrmul24_fa15_22_y2;
  assign f_u_arrmul24_fa14_23_y2 = f_u_arrmul24_fa14_23_y0 ^ f_u_arrmul24_fa14_23_f_u_arrmul24_fa13_23_y4;
  assign f_u_arrmul24_fa14_23_y3 = f_u_arrmul24_fa14_23_y0 & f_u_arrmul24_fa14_23_f_u_arrmul24_fa13_23_y4;
  assign f_u_arrmul24_fa14_23_y4 = f_u_arrmul24_fa14_23_y1 | f_u_arrmul24_fa14_23_y3;
  assign f_u_arrmul24_and15_23_a_15 = a_15;
  assign f_u_arrmul24_and15_23_b_23 = b_23;
  assign f_u_arrmul24_and15_23_y0 = f_u_arrmul24_and15_23_a_15 & f_u_arrmul24_and15_23_b_23;
  assign f_u_arrmul24_fa15_23_f_u_arrmul24_and15_23_y0 = f_u_arrmul24_and15_23_y0;
  assign f_u_arrmul24_fa15_23_f_u_arrmul24_fa16_22_y2 = f_u_arrmul24_fa16_22_y2;
  assign f_u_arrmul24_fa15_23_f_u_arrmul24_fa14_23_y4 = f_u_arrmul24_fa14_23_y4;
  assign f_u_arrmul24_fa15_23_y0 = f_u_arrmul24_fa15_23_f_u_arrmul24_and15_23_y0 ^ f_u_arrmul24_fa15_23_f_u_arrmul24_fa16_22_y2;
  assign f_u_arrmul24_fa15_23_y1 = f_u_arrmul24_fa15_23_f_u_arrmul24_and15_23_y0 & f_u_arrmul24_fa15_23_f_u_arrmul24_fa16_22_y2;
  assign f_u_arrmul24_fa15_23_y2 = f_u_arrmul24_fa15_23_y0 ^ f_u_arrmul24_fa15_23_f_u_arrmul24_fa14_23_y4;
  assign f_u_arrmul24_fa15_23_y3 = f_u_arrmul24_fa15_23_y0 & f_u_arrmul24_fa15_23_f_u_arrmul24_fa14_23_y4;
  assign f_u_arrmul24_fa15_23_y4 = f_u_arrmul24_fa15_23_y1 | f_u_arrmul24_fa15_23_y3;
  assign f_u_arrmul24_and16_23_a_16 = a_16;
  assign f_u_arrmul24_and16_23_b_23 = b_23;
  assign f_u_arrmul24_and16_23_y0 = f_u_arrmul24_and16_23_a_16 & f_u_arrmul24_and16_23_b_23;
  assign f_u_arrmul24_fa16_23_f_u_arrmul24_and16_23_y0 = f_u_arrmul24_and16_23_y0;
  assign f_u_arrmul24_fa16_23_f_u_arrmul24_fa17_22_y2 = f_u_arrmul24_fa17_22_y2;
  assign f_u_arrmul24_fa16_23_f_u_arrmul24_fa15_23_y4 = f_u_arrmul24_fa15_23_y4;
  assign f_u_arrmul24_fa16_23_y0 = f_u_arrmul24_fa16_23_f_u_arrmul24_and16_23_y0 ^ f_u_arrmul24_fa16_23_f_u_arrmul24_fa17_22_y2;
  assign f_u_arrmul24_fa16_23_y1 = f_u_arrmul24_fa16_23_f_u_arrmul24_and16_23_y0 & f_u_arrmul24_fa16_23_f_u_arrmul24_fa17_22_y2;
  assign f_u_arrmul24_fa16_23_y2 = f_u_arrmul24_fa16_23_y0 ^ f_u_arrmul24_fa16_23_f_u_arrmul24_fa15_23_y4;
  assign f_u_arrmul24_fa16_23_y3 = f_u_arrmul24_fa16_23_y0 & f_u_arrmul24_fa16_23_f_u_arrmul24_fa15_23_y4;
  assign f_u_arrmul24_fa16_23_y4 = f_u_arrmul24_fa16_23_y1 | f_u_arrmul24_fa16_23_y3;
  assign f_u_arrmul24_and17_23_a_17 = a_17;
  assign f_u_arrmul24_and17_23_b_23 = b_23;
  assign f_u_arrmul24_and17_23_y0 = f_u_arrmul24_and17_23_a_17 & f_u_arrmul24_and17_23_b_23;
  assign f_u_arrmul24_fa17_23_f_u_arrmul24_and17_23_y0 = f_u_arrmul24_and17_23_y0;
  assign f_u_arrmul24_fa17_23_f_u_arrmul24_fa18_22_y2 = f_u_arrmul24_fa18_22_y2;
  assign f_u_arrmul24_fa17_23_f_u_arrmul24_fa16_23_y4 = f_u_arrmul24_fa16_23_y4;
  assign f_u_arrmul24_fa17_23_y0 = f_u_arrmul24_fa17_23_f_u_arrmul24_and17_23_y0 ^ f_u_arrmul24_fa17_23_f_u_arrmul24_fa18_22_y2;
  assign f_u_arrmul24_fa17_23_y1 = f_u_arrmul24_fa17_23_f_u_arrmul24_and17_23_y0 & f_u_arrmul24_fa17_23_f_u_arrmul24_fa18_22_y2;
  assign f_u_arrmul24_fa17_23_y2 = f_u_arrmul24_fa17_23_y0 ^ f_u_arrmul24_fa17_23_f_u_arrmul24_fa16_23_y4;
  assign f_u_arrmul24_fa17_23_y3 = f_u_arrmul24_fa17_23_y0 & f_u_arrmul24_fa17_23_f_u_arrmul24_fa16_23_y4;
  assign f_u_arrmul24_fa17_23_y4 = f_u_arrmul24_fa17_23_y1 | f_u_arrmul24_fa17_23_y3;
  assign f_u_arrmul24_and18_23_a_18 = a_18;
  assign f_u_arrmul24_and18_23_b_23 = b_23;
  assign f_u_arrmul24_and18_23_y0 = f_u_arrmul24_and18_23_a_18 & f_u_arrmul24_and18_23_b_23;
  assign f_u_arrmul24_fa18_23_f_u_arrmul24_and18_23_y0 = f_u_arrmul24_and18_23_y0;
  assign f_u_arrmul24_fa18_23_f_u_arrmul24_fa19_22_y2 = f_u_arrmul24_fa19_22_y2;
  assign f_u_arrmul24_fa18_23_f_u_arrmul24_fa17_23_y4 = f_u_arrmul24_fa17_23_y4;
  assign f_u_arrmul24_fa18_23_y0 = f_u_arrmul24_fa18_23_f_u_arrmul24_and18_23_y0 ^ f_u_arrmul24_fa18_23_f_u_arrmul24_fa19_22_y2;
  assign f_u_arrmul24_fa18_23_y1 = f_u_arrmul24_fa18_23_f_u_arrmul24_and18_23_y0 & f_u_arrmul24_fa18_23_f_u_arrmul24_fa19_22_y2;
  assign f_u_arrmul24_fa18_23_y2 = f_u_arrmul24_fa18_23_y0 ^ f_u_arrmul24_fa18_23_f_u_arrmul24_fa17_23_y4;
  assign f_u_arrmul24_fa18_23_y3 = f_u_arrmul24_fa18_23_y0 & f_u_arrmul24_fa18_23_f_u_arrmul24_fa17_23_y4;
  assign f_u_arrmul24_fa18_23_y4 = f_u_arrmul24_fa18_23_y1 | f_u_arrmul24_fa18_23_y3;
  assign f_u_arrmul24_and19_23_a_19 = a_19;
  assign f_u_arrmul24_and19_23_b_23 = b_23;
  assign f_u_arrmul24_and19_23_y0 = f_u_arrmul24_and19_23_a_19 & f_u_arrmul24_and19_23_b_23;
  assign f_u_arrmul24_fa19_23_f_u_arrmul24_and19_23_y0 = f_u_arrmul24_and19_23_y0;
  assign f_u_arrmul24_fa19_23_f_u_arrmul24_fa20_22_y2 = f_u_arrmul24_fa20_22_y2;
  assign f_u_arrmul24_fa19_23_f_u_arrmul24_fa18_23_y4 = f_u_arrmul24_fa18_23_y4;
  assign f_u_arrmul24_fa19_23_y0 = f_u_arrmul24_fa19_23_f_u_arrmul24_and19_23_y0 ^ f_u_arrmul24_fa19_23_f_u_arrmul24_fa20_22_y2;
  assign f_u_arrmul24_fa19_23_y1 = f_u_arrmul24_fa19_23_f_u_arrmul24_and19_23_y0 & f_u_arrmul24_fa19_23_f_u_arrmul24_fa20_22_y2;
  assign f_u_arrmul24_fa19_23_y2 = f_u_arrmul24_fa19_23_y0 ^ f_u_arrmul24_fa19_23_f_u_arrmul24_fa18_23_y4;
  assign f_u_arrmul24_fa19_23_y3 = f_u_arrmul24_fa19_23_y0 & f_u_arrmul24_fa19_23_f_u_arrmul24_fa18_23_y4;
  assign f_u_arrmul24_fa19_23_y4 = f_u_arrmul24_fa19_23_y1 | f_u_arrmul24_fa19_23_y3;
  assign f_u_arrmul24_and20_23_a_20 = a_20;
  assign f_u_arrmul24_and20_23_b_23 = b_23;
  assign f_u_arrmul24_and20_23_y0 = f_u_arrmul24_and20_23_a_20 & f_u_arrmul24_and20_23_b_23;
  assign f_u_arrmul24_fa20_23_f_u_arrmul24_and20_23_y0 = f_u_arrmul24_and20_23_y0;
  assign f_u_arrmul24_fa20_23_f_u_arrmul24_fa21_22_y2 = f_u_arrmul24_fa21_22_y2;
  assign f_u_arrmul24_fa20_23_f_u_arrmul24_fa19_23_y4 = f_u_arrmul24_fa19_23_y4;
  assign f_u_arrmul24_fa20_23_y0 = f_u_arrmul24_fa20_23_f_u_arrmul24_and20_23_y0 ^ f_u_arrmul24_fa20_23_f_u_arrmul24_fa21_22_y2;
  assign f_u_arrmul24_fa20_23_y1 = f_u_arrmul24_fa20_23_f_u_arrmul24_and20_23_y0 & f_u_arrmul24_fa20_23_f_u_arrmul24_fa21_22_y2;
  assign f_u_arrmul24_fa20_23_y2 = f_u_arrmul24_fa20_23_y0 ^ f_u_arrmul24_fa20_23_f_u_arrmul24_fa19_23_y4;
  assign f_u_arrmul24_fa20_23_y3 = f_u_arrmul24_fa20_23_y0 & f_u_arrmul24_fa20_23_f_u_arrmul24_fa19_23_y4;
  assign f_u_arrmul24_fa20_23_y4 = f_u_arrmul24_fa20_23_y1 | f_u_arrmul24_fa20_23_y3;
  assign f_u_arrmul24_and21_23_a_21 = a_21;
  assign f_u_arrmul24_and21_23_b_23 = b_23;
  assign f_u_arrmul24_and21_23_y0 = f_u_arrmul24_and21_23_a_21 & f_u_arrmul24_and21_23_b_23;
  assign f_u_arrmul24_fa21_23_f_u_arrmul24_and21_23_y0 = f_u_arrmul24_and21_23_y0;
  assign f_u_arrmul24_fa21_23_f_u_arrmul24_fa22_22_y2 = f_u_arrmul24_fa22_22_y2;
  assign f_u_arrmul24_fa21_23_f_u_arrmul24_fa20_23_y4 = f_u_arrmul24_fa20_23_y4;
  assign f_u_arrmul24_fa21_23_y0 = f_u_arrmul24_fa21_23_f_u_arrmul24_and21_23_y0 ^ f_u_arrmul24_fa21_23_f_u_arrmul24_fa22_22_y2;
  assign f_u_arrmul24_fa21_23_y1 = f_u_arrmul24_fa21_23_f_u_arrmul24_and21_23_y0 & f_u_arrmul24_fa21_23_f_u_arrmul24_fa22_22_y2;
  assign f_u_arrmul24_fa21_23_y2 = f_u_arrmul24_fa21_23_y0 ^ f_u_arrmul24_fa21_23_f_u_arrmul24_fa20_23_y4;
  assign f_u_arrmul24_fa21_23_y3 = f_u_arrmul24_fa21_23_y0 & f_u_arrmul24_fa21_23_f_u_arrmul24_fa20_23_y4;
  assign f_u_arrmul24_fa21_23_y4 = f_u_arrmul24_fa21_23_y1 | f_u_arrmul24_fa21_23_y3;
  assign f_u_arrmul24_and22_23_a_22 = a_22;
  assign f_u_arrmul24_and22_23_b_23 = b_23;
  assign f_u_arrmul24_and22_23_y0 = f_u_arrmul24_and22_23_a_22 & f_u_arrmul24_and22_23_b_23;
  assign f_u_arrmul24_fa22_23_f_u_arrmul24_and22_23_y0 = f_u_arrmul24_and22_23_y0;
  assign f_u_arrmul24_fa22_23_f_u_arrmul24_fa23_22_y2 = f_u_arrmul24_fa23_22_y2;
  assign f_u_arrmul24_fa22_23_f_u_arrmul24_fa21_23_y4 = f_u_arrmul24_fa21_23_y4;
  assign f_u_arrmul24_fa22_23_y0 = f_u_arrmul24_fa22_23_f_u_arrmul24_and22_23_y0 ^ f_u_arrmul24_fa22_23_f_u_arrmul24_fa23_22_y2;
  assign f_u_arrmul24_fa22_23_y1 = f_u_arrmul24_fa22_23_f_u_arrmul24_and22_23_y0 & f_u_arrmul24_fa22_23_f_u_arrmul24_fa23_22_y2;
  assign f_u_arrmul24_fa22_23_y2 = f_u_arrmul24_fa22_23_y0 ^ f_u_arrmul24_fa22_23_f_u_arrmul24_fa21_23_y4;
  assign f_u_arrmul24_fa22_23_y3 = f_u_arrmul24_fa22_23_y0 & f_u_arrmul24_fa22_23_f_u_arrmul24_fa21_23_y4;
  assign f_u_arrmul24_fa22_23_y4 = f_u_arrmul24_fa22_23_y1 | f_u_arrmul24_fa22_23_y3;
  assign f_u_arrmul24_and23_23_a_23 = a_23;
  assign f_u_arrmul24_and23_23_b_23 = b_23;
  assign f_u_arrmul24_and23_23_y0 = f_u_arrmul24_and23_23_a_23 & f_u_arrmul24_and23_23_b_23;
  assign f_u_arrmul24_fa23_23_f_u_arrmul24_and23_23_y0 = f_u_arrmul24_and23_23_y0;
  assign f_u_arrmul24_fa23_23_f_u_arrmul24_fa23_22_y4 = f_u_arrmul24_fa23_22_y4;
  assign f_u_arrmul24_fa23_23_f_u_arrmul24_fa22_23_y4 = f_u_arrmul24_fa22_23_y4;
  assign f_u_arrmul24_fa23_23_y0 = f_u_arrmul24_fa23_23_f_u_arrmul24_and23_23_y0 ^ f_u_arrmul24_fa23_23_f_u_arrmul24_fa23_22_y4;
  assign f_u_arrmul24_fa23_23_y1 = f_u_arrmul24_fa23_23_f_u_arrmul24_and23_23_y0 & f_u_arrmul24_fa23_23_f_u_arrmul24_fa23_22_y4;
  assign f_u_arrmul24_fa23_23_y2 = f_u_arrmul24_fa23_23_y0 ^ f_u_arrmul24_fa23_23_f_u_arrmul24_fa22_23_y4;
  assign f_u_arrmul24_fa23_23_y3 = f_u_arrmul24_fa23_23_y0 & f_u_arrmul24_fa23_23_f_u_arrmul24_fa22_23_y4;
  assign f_u_arrmul24_fa23_23_y4 = f_u_arrmul24_fa23_23_y1 | f_u_arrmul24_fa23_23_y3;

  assign out[0] = f_u_arrmul24_and0_0_y0;
  assign out[1] = f_u_arrmul24_ha0_1_y0;
  assign out[2] = f_u_arrmul24_ha0_2_y0;
  assign out[3] = f_u_arrmul24_ha0_3_y0;
  assign out[4] = f_u_arrmul24_ha0_4_y0;
  assign out[5] = f_u_arrmul24_ha0_5_y0;
  assign out[6] = f_u_arrmul24_ha0_6_y0;
  assign out[7] = f_u_arrmul24_ha0_7_y0;
  assign out[8] = f_u_arrmul24_ha0_8_y0;
  assign out[9] = f_u_arrmul24_ha0_9_y0;
  assign out[10] = f_u_arrmul24_ha0_10_y0;
  assign out[11] = f_u_arrmul24_ha0_11_y0;
  assign out[12] = f_u_arrmul24_ha0_12_y0;
  assign out[13] = f_u_arrmul24_ha0_13_y0;
  assign out[14] = f_u_arrmul24_ha0_14_y0;
  assign out[15] = f_u_arrmul24_ha0_15_y0;
  assign out[16] = f_u_arrmul24_ha0_16_y0;
  assign out[17] = f_u_arrmul24_ha0_17_y0;
  assign out[18] = f_u_arrmul24_ha0_18_y0;
  assign out[19] = f_u_arrmul24_ha0_19_y0;
  assign out[20] = f_u_arrmul24_ha0_20_y0;
  assign out[21] = f_u_arrmul24_ha0_21_y0;
  assign out[22] = f_u_arrmul24_ha0_22_y0;
  assign out[23] = f_u_arrmul24_ha0_23_y0;
  assign out[24] = f_u_arrmul24_fa1_23_y2;
  assign out[25] = f_u_arrmul24_fa2_23_y2;
  assign out[26] = f_u_arrmul24_fa3_23_y2;
  assign out[27] = f_u_arrmul24_fa4_23_y2;
  assign out[28] = f_u_arrmul24_fa5_23_y2;
  assign out[29] = f_u_arrmul24_fa6_23_y2;
  assign out[30] = f_u_arrmul24_fa7_23_y2;
  assign out[31] = f_u_arrmul24_fa8_23_y2;
  assign out[32] = f_u_arrmul24_fa9_23_y2;
  assign out[33] = f_u_arrmul24_fa10_23_y2;
  assign out[34] = f_u_arrmul24_fa11_23_y2;
  assign out[35] = f_u_arrmul24_fa12_23_y2;
  assign out[36] = f_u_arrmul24_fa13_23_y2;
  assign out[37] = f_u_arrmul24_fa14_23_y2;
  assign out[38] = f_u_arrmul24_fa15_23_y2;
  assign out[39] = f_u_arrmul24_fa16_23_y2;
  assign out[40] = f_u_arrmul24_fa17_23_y2;
  assign out[41] = f_u_arrmul24_fa18_23_y2;
  assign out[42] = f_u_arrmul24_fa19_23_y2;
  assign out[43] = f_u_arrmul24_fa20_23_y2;
  assign out[44] = f_u_arrmul24_fa21_23_y2;
  assign out[45] = f_u_arrmul24_fa22_23_y2;
  assign out[46] = f_u_arrmul24_fa23_23_y2;
  assign out[47] = f_u_arrmul24_fa23_23_y4;
endmodule