module f_s_pg_rca24(input [23:0] a, input [23:0] b, output [24:0] f_s_pg_rca24_out);
  wire f_s_pg_rca24_pg_fa0_xor0;
  wire f_s_pg_rca24_pg_fa0_and0;
  wire f_s_pg_rca24_pg_fa1_xor0;
  wire f_s_pg_rca24_pg_fa1_and0;
  wire f_s_pg_rca24_pg_fa1_xor1;
  wire f_s_pg_rca24_and1;
  wire f_s_pg_rca24_or1;
  wire f_s_pg_rca24_pg_fa2_xor0;
  wire f_s_pg_rca24_pg_fa2_and0;
  wire f_s_pg_rca24_pg_fa2_xor1;
  wire f_s_pg_rca24_and2;
  wire f_s_pg_rca24_or2;
  wire f_s_pg_rca24_pg_fa3_xor0;
  wire f_s_pg_rca24_pg_fa3_and0;
  wire f_s_pg_rca24_pg_fa3_xor1;
  wire f_s_pg_rca24_and3;
  wire f_s_pg_rca24_or3;
  wire f_s_pg_rca24_pg_fa4_xor0;
  wire f_s_pg_rca24_pg_fa4_and0;
  wire f_s_pg_rca24_pg_fa4_xor1;
  wire f_s_pg_rca24_and4;
  wire f_s_pg_rca24_or4;
  wire f_s_pg_rca24_pg_fa5_xor0;
  wire f_s_pg_rca24_pg_fa5_and0;
  wire f_s_pg_rca24_pg_fa5_xor1;
  wire f_s_pg_rca24_and5;
  wire f_s_pg_rca24_or5;
  wire f_s_pg_rca24_pg_fa6_xor0;
  wire f_s_pg_rca24_pg_fa6_and0;
  wire f_s_pg_rca24_pg_fa6_xor1;
  wire f_s_pg_rca24_and6;
  wire f_s_pg_rca24_or6;
  wire f_s_pg_rca24_pg_fa7_xor0;
  wire f_s_pg_rca24_pg_fa7_and0;
  wire f_s_pg_rca24_pg_fa7_xor1;
  wire f_s_pg_rca24_and7;
  wire f_s_pg_rca24_or7;
  wire f_s_pg_rca24_pg_fa8_xor0;
  wire f_s_pg_rca24_pg_fa8_and0;
  wire f_s_pg_rca24_pg_fa8_xor1;
  wire f_s_pg_rca24_and8;
  wire f_s_pg_rca24_or8;
  wire f_s_pg_rca24_pg_fa9_xor0;
  wire f_s_pg_rca24_pg_fa9_and0;
  wire f_s_pg_rca24_pg_fa9_xor1;
  wire f_s_pg_rca24_and9;
  wire f_s_pg_rca24_or9;
  wire f_s_pg_rca24_pg_fa10_xor0;
  wire f_s_pg_rca24_pg_fa10_and0;
  wire f_s_pg_rca24_pg_fa10_xor1;
  wire f_s_pg_rca24_and10;
  wire f_s_pg_rca24_or10;
  wire f_s_pg_rca24_pg_fa11_xor0;
  wire f_s_pg_rca24_pg_fa11_and0;
  wire f_s_pg_rca24_pg_fa11_xor1;
  wire f_s_pg_rca24_and11;
  wire f_s_pg_rca24_or11;
  wire f_s_pg_rca24_pg_fa12_xor0;
  wire f_s_pg_rca24_pg_fa12_and0;
  wire f_s_pg_rca24_pg_fa12_xor1;
  wire f_s_pg_rca24_and12;
  wire f_s_pg_rca24_or12;
  wire f_s_pg_rca24_pg_fa13_xor0;
  wire f_s_pg_rca24_pg_fa13_and0;
  wire f_s_pg_rca24_pg_fa13_xor1;
  wire f_s_pg_rca24_and13;
  wire f_s_pg_rca24_or13;
  wire f_s_pg_rca24_pg_fa14_xor0;
  wire f_s_pg_rca24_pg_fa14_and0;
  wire f_s_pg_rca24_pg_fa14_xor1;
  wire f_s_pg_rca24_and14;
  wire f_s_pg_rca24_or14;
  wire f_s_pg_rca24_pg_fa15_xor0;
  wire f_s_pg_rca24_pg_fa15_and0;
  wire f_s_pg_rca24_pg_fa15_xor1;
  wire f_s_pg_rca24_and15;
  wire f_s_pg_rca24_or15;
  wire f_s_pg_rca24_pg_fa16_xor0;
  wire f_s_pg_rca24_pg_fa16_and0;
  wire f_s_pg_rca24_pg_fa16_xor1;
  wire f_s_pg_rca24_and16;
  wire f_s_pg_rca24_or16;
  wire f_s_pg_rca24_pg_fa17_xor0;
  wire f_s_pg_rca24_pg_fa17_and0;
  wire f_s_pg_rca24_pg_fa17_xor1;
  wire f_s_pg_rca24_and17;
  wire f_s_pg_rca24_or17;
  wire f_s_pg_rca24_pg_fa18_xor0;
  wire f_s_pg_rca24_pg_fa18_and0;
  wire f_s_pg_rca24_pg_fa18_xor1;
  wire f_s_pg_rca24_and18;
  wire f_s_pg_rca24_or18;
  wire f_s_pg_rca24_pg_fa19_xor0;
  wire f_s_pg_rca24_pg_fa19_and0;
  wire f_s_pg_rca24_pg_fa19_xor1;
  wire f_s_pg_rca24_and19;
  wire f_s_pg_rca24_or19;
  wire f_s_pg_rca24_pg_fa20_xor0;
  wire f_s_pg_rca24_pg_fa20_and0;
  wire f_s_pg_rca24_pg_fa20_xor1;
  wire f_s_pg_rca24_and20;
  wire f_s_pg_rca24_or20;
  wire f_s_pg_rca24_pg_fa21_xor0;
  wire f_s_pg_rca24_pg_fa21_and0;
  wire f_s_pg_rca24_pg_fa21_xor1;
  wire f_s_pg_rca24_and21;
  wire f_s_pg_rca24_or21;
  wire f_s_pg_rca24_pg_fa22_xor0;
  wire f_s_pg_rca24_pg_fa22_and0;
  wire f_s_pg_rca24_pg_fa22_xor1;
  wire f_s_pg_rca24_and22;
  wire f_s_pg_rca24_or22;
  wire f_s_pg_rca24_pg_fa23_xor0;
  wire f_s_pg_rca24_pg_fa23_and0;
  wire f_s_pg_rca24_pg_fa23_xor1;
  wire f_s_pg_rca24_and23;
  wire f_s_pg_rca24_or23;
  wire f_s_pg_rca24_xor0;
  wire f_s_pg_rca24_xor1;

  assign f_s_pg_rca24_pg_fa0_xor0 = a[0] ^ b[0];
  assign f_s_pg_rca24_pg_fa0_and0 = a[0] & b[0];
  assign f_s_pg_rca24_pg_fa1_xor0 = a[1] ^ b[1];
  assign f_s_pg_rca24_pg_fa1_and0 = a[1] & b[1];
  assign f_s_pg_rca24_pg_fa1_xor1 = f_s_pg_rca24_pg_fa1_xor0 ^ f_s_pg_rca24_pg_fa0_and0;
  assign f_s_pg_rca24_and1 = f_s_pg_rca24_pg_fa0_and0 & f_s_pg_rca24_pg_fa1_xor0;
  assign f_s_pg_rca24_or1 = f_s_pg_rca24_and1 | f_s_pg_rca24_pg_fa1_and0;
  assign f_s_pg_rca24_pg_fa2_xor0 = a[2] ^ b[2];
  assign f_s_pg_rca24_pg_fa2_and0 = a[2] & b[2];
  assign f_s_pg_rca24_pg_fa2_xor1 = f_s_pg_rca24_pg_fa2_xor0 ^ f_s_pg_rca24_or1;
  assign f_s_pg_rca24_and2 = f_s_pg_rca24_or1 & f_s_pg_rca24_pg_fa2_xor0;
  assign f_s_pg_rca24_or2 = f_s_pg_rca24_and2 | f_s_pg_rca24_pg_fa2_and0;
  assign f_s_pg_rca24_pg_fa3_xor0 = a[3] ^ b[3];
  assign f_s_pg_rca24_pg_fa3_and0 = a[3] & b[3];
  assign f_s_pg_rca24_pg_fa3_xor1 = f_s_pg_rca24_pg_fa3_xor0 ^ f_s_pg_rca24_or2;
  assign f_s_pg_rca24_and3 = f_s_pg_rca24_or2 & f_s_pg_rca24_pg_fa3_xor0;
  assign f_s_pg_rca24_or3 = f_s_pg_rca24_and3 | f_s_pg_rca24_pg_fa3_and0;
  assign f_s_pg_rca24_pg_fa4_xor0 = a[4] ^ b[4];
  assign f_s_pg_rca24_pg_fa4_and0 = a[4] & b[4];
  assign f_s_pg_rca24_pg_fa4_xor1 = f_s_pg_rca24_pg_fa4_xor0 ^ f_s_pg_rca24_or3;
  assign f_s_pg_rca24_and4 = f_s_pg_rca24_or3 & f_s_pg_rca24_pg_fa4_xor0;
  assign f_s_pg_rca24_or4 = f_s_pg_rca24_and4 | f_s_pg_rca24_pg_fa4_and0;
  assign f_s_pg_rca24_pg_fa5_xor0 = a[5] ^ b[5];
  assign f_s_pg_rca24_pg_fa5_and0 = a[5] & b[5];
  assign f_s_pg_rca24_pg_fa5_xor1 = f_s_pg_rca24_pg_fa5_xor0 ^ f_s_pg_rca24_or4;
  assign f_s_pg_rca24_and5 = f_s_pg_rca24_or4 & f_s_pg_rca24_pg_fa5_xor0;
  assign f_s_pg_rca24_or5 = f_s_pg_rca24_and5 | f_s_pg_rca24_pg_fa5_and0;
  assign f_s_pg_rca24_pg_fa6_xor0 = a[6] ^ b[6];
  assign f_s_pg_rca24_pg_fa6_and0 = a[6] & b[6];
  assign f_s_pg_rca24_pg_fa6_xor1 = f_s_pg_rca24_pg_fa6_xor0 ^ f_s_pg_rca24_or5;
  assign f_s_pg_rca24_and6 = f_s_pg_rca24_or5 & f_s_pg_rca24_pg_fa6_xor0;
  assign f_s_pg_rca24_or6 = f_s_pg_rca24_and6 | f_s_pg_rca24_pg_fa6_and0;
  assign f_s_pg_rca24_pg_fa7_xor0 = a[7] ^ b[7];
  assign f_s_pg_rca24_pg_fa7_and0 = a[7] & b[7];
  assign f_s_pg_rca24_pg_fa7_xor1 = f_s_pg_rca24_pg_fa7_xor0 ^ f_s_pg_rca24_or6;
  assign f_s_pg_rca24_and7 = f_s_pg_rca24_or6 & f_s_pg_rca24_pg_fa7_xor0;
  assign f_s_pg_rca24_or7 = f_s_pg_rca24_and7 | f_s_pg_rca24_pg_fa7_and0;
  assign f_s_pg_rca24_pg_fa8_xor0 = a[8] ^ b[8];
  assign f_s_pg_rca24_pg_fa8_and0 = a[8] & b[8];
  assign f_s_pg_rca24_pg_fa8_xor1 = f_s_pg_rca24_pg_fa8_xor0 ^ f_s_pg_rca24_or7;
  assign f_s_pg_rca24_and8 = f_s_pg_rca24_or7 & f_s_pg_rca24_pg_fa8_xor0;
  assign f_s_pg_rca24_or8 = f_s_pg_rca24_and8 | f_s_pg_rca24_pg_fa8_and0;
  assign f_s_pg_rca24_pg_fa9_xor0 = a[9] ^ b[9];
  assign f_s_pg_rca24_pg_fa9_and0 = a[9] & b[9];
  assign f_s_pg_rca24_pg_fa9_xor1 = f_s_pg_rca24_pg_fa9_xor0 ^ f_s_pg_rca24_or8;
  assign f_s_pg_rca24_and9 = f_s_pg_rca24_or8 & f_s_pg_rca24_pg_fa9_xor0;
  assign f_s_pg_rca24_or9 = f_s_pg_rca24_and9 | f_s_pg_rca24_pg_fa9_and0;
  assign f_s_pg_rca24_pg_fa10_xor0 = a[10] ^ b[10];
  assign f_s_pg_rca24_pg_fa10_and0 = a[10] & b[10];
  assign f_s_pg_rca24_pg_fa10_xor1 = f_s_pg_rca24_pg_fa10_xor0 ^ f_s_pg_rca24_or9;
  assign f_s_pg_rca24_and10 = f_s_pg_rca24_or9 & f_s_pg_rca24_pg_fa10_xor0;
  assign f_s_pg_rca24_or10 = f_s_pg_rca24_and10 | f_s_pg_rca24_pg_fa10_and0;
  assign f_s_pg_rca24_pg_fa11_xor0 = a[11] ^ b[11];
  assign f_s_pg_rca24_pg_fa11_and0 = a[11] & b[11];
  assign f_s_pg_rca24_pg_fa11_xor1 = f_s_pg_rca24_pg_fa11_xor0 ^ f_s_pg_rca24_or10;
  assign f_s_pg_rca24_and11 = f_s_pg_rca24_or10 & f_s_pg_rca24_pg_fa11_xor0;
  assign f_s_pg_rca24_or11 = f_s_pg_rca24_and11 | f_s_pg_rca24_pg_fa11_and0;
  assign f_s_pg_rca24_pg_fa12_xor0 = a[12] ^ b[12];
  assign f_s_pg_rca24_pg_fa12_and0 = a[12] & b[12];
  assign f_s_pg_rca24_pg_fa12_xor1 = f_s_pg_rca24_pg_fa12_xor0 ^ f_s_pg_rca24_or11;
  assign f_s_pg_rca24_and12 = f_s_pg_rca24_or11 & f_s_pg_rca24_pg_fa12_xor0;
  assign f_s_pg_rca24_or12 = f_s_pg_rca24_and12 | f_s_pg_rca24_pg_fa12_and0;
  assign f_s_pg_rca24_pg_fa13_xor0 = a[13] ^ b[13];
  assign f_s_pg_rca24_pg_fa13_and0 = a[13] & b[13];
  assign f_s_pg_rca24_pg_fa13_xor1 = f_s_pg_rca24_pg_fa13_xor0 ^ f_s_pg_rca24_or12;
  assign f_s_pg_rca24_and13 = f_s_pg_rca24_or12 & f_s_pg_rca24_pg_fa13_xor0;
  assign f_s_pg_rca24_or13 = f_s_pg_rca24_and13 | f_s_pg_rca24_pg_fa13_and0;
  assign f_s_pg_rca24_pg_fa14_xor0 = a[14] ^ b[14];
  assign f_s_pg_rca24_pg_fa14_and0 = a[14] & b[14];
  assign f_s_pg_rca24_pg_fa14_xor1 = f_s_pg_rca24_pg_fa14_xor0 ^ f_s_pg_rca24_or13;
  assign f_s_pg_rca24_and14 = f_s_pg_rca24_or13 & f_s_pg_rca24_pg_fa14_xor0;
  assign f_s_pg_rca24_or14 = f_s_pg_rca24_and14 | f_s_pg_rca24_pg_fa14_and0;
  assign f_s_pg_rca24_pg_fa15_xor0 = a[15] ^ b[15];
  assign f_s_pg_rca24_pg_fa15_and0 = a[15] & b[15];
  assign f_s_pg_rca24_pg_fa15_xor1 = f_s_pg_rca24_pg_fa15_xor0 ^ f_s_pg_rca24_or14;
  assign f_s_pg_rca24_and15 = f_s_pg_rca24_or14 & f_s_pg_rca24_pg_fa15_xor0;
  assign f_s_pg_rca24_or15 = f_s_pg_rca24_and15 | f_s_pg_rca24_pg_fa15_and0;
  assign f_s_pg_rca24_pg_fa16_xor0 = a[16] ^ b[16];
  assign f_s_pg_rca24_pg_fa16_and0 = a[16] & b[16];
  assign f_s_pg_rca24_pg_fa16_xor1 = f_s_pg_rca24_pg_fa16_xor0 ^ f_s_pg_rca24_or15;
  assign f_s_pg_rca24_and16 = f_s_pg_rca24_or15 & f_s_pg_rca24_pg_fa16_xor0;
  assign f_s_pg_rca24_or16 = f_s_pg_rca24_and16 | f_s_pg_rca24_pg_fa16_and0;
  assign f_s_pg_rca24_pg_fa17_xor0 = a[17] ^ b[17];
  assign f_s_pg_rca24_pg_fa17_and0 = a[17] & b[17];
  assign f_s_pg_rca24_pg_fa17_xor1 = f_s_pg_rca24_pg_fa17_xor0 ^ f_s_pg_rca24_or16;
  assign f_s_pg_rca24_and17 = f_s_pg_rca24_or16 & f_s_pg_rca24_pg_fa17_xor0;
  assign f_s_pg_rca24_or17 = f_s_pg_rca24_and17 | f_s_pg_rca24_pg_fa17_and0;
  assign f_s_pg_rca24_pg_fa18_xor0 = a[18] ^ b[18];
  assign f_s_pg_rca24_pg_fa18_and0 = a[18] & b[18];
  assign f_s_pg_rca24_pg_fa18_xor1 = f_s_pg_rca24_pg_fa18_xor0 ^ f_s_pg_rca24_or17;
  assign f_s_pg_rca24_and18 = f_s_pg_rca24_or17 & f_s_pg_rca24_pg_fa18_xor0;
  assign f_s_pg_rca24_or18 = f_s_pg_rca24_and18 | f_s_pg_rca24_pg_fa18_and0;
  assign f_s_pg_rca24_pg_fa19_xor0 = a[19] ^ b[19];
  assign f_s_pg_rca24_pg_fa19_and0 = a[19] & b[19];
  assign f_s_pg_rca24_pg_fa19_xor1 = f_s_pg_rca24_pg_fa19_xor0 ^ f_s_pg_rca24_or18;
  assign f_s_pg_rca24_and19 = f_s_pg_rca24_or18 & f_s_pg_rca24_pg_fa19_xor0;
  assign f_s_pg_rca24_or19 = f_s_pg_rca24_and19 | f_s_pg_rca24_pg_fa19_and0;
  assign f_s_pg_rca24_pg_fa20_xor0 = a[20] ^ b[20];
  assign f_s_pg_rca24_pg_fa20_and0 = a[20] & b[20];
  assign f_s_pg_rca24_pg_fa20_xor1 = f_s_pg_rca24_pg_fa20_xor0 ^ f_s_pg_rca24_or19;
  assign f_s_pg_rca24_and20 = f_s_pg_rca24_or19 & f_s_pg_rca24_pg_fa20_xor0;
  assign f_s_pg_rca24_or20 = f_s_pg_rca24_and20 | f_s_pg_rca24_pg_fa20_and0;
  assign f_s_pg_rca24_pg_fa21_xor0 = a[21] ^ b[21];
  assign f_s_pg_rca24_pg_fa21_and0 = a[21] & b[21];
  assign f_s_pg_rca24_pg_fa21_xor1 = f_s_pg_rca24_pg_fa21_xor0 ^ f_s_pg_rca24_or20;
  assign f_s_pg_rca24_and21 = f_s_pg_rca24_or20 & f_s_pg_rca24_pg_fa21_xor0;
  assign f_s_pg_rca24_or21 = f_s_pg_rca24_and21 | f_s_pg_rca24_pg_fa21_and0;
  assign f_s_pg_rca24_pg_fa22_xor0 = a[22] ^ b[22];
  assign f_s_pg_rca24_pg_fa22_and0 = a[22] & b[22];
  assign f_s_pg_rca24_pg_fa22_xor1 = f_s_pg_rca24_pg_fa22_xor0 ^ f_s_pg_rca24_or21;
  assign f_s_pg_rca24_and22 = f_s_pg_rca24_or21 & f_s_pg_rca24_pg_fa22_xor0;
  assign f_s_pg_rca24_or22 = f_s_pg_rca24_and22 | f_s_pg_rca24_pg_fa22_and0;
  assign f_s_pg_rca24_pg_fa23_xor0 = a[23] ^ b[23];
  assign f_s_pg_rca24_pg_fa23_and0 = a[23] & b[23];
  assign f_s_pg_rca24_pg_fa23_xor1 = f_s_pg_rca24_pg_fa23_xor0 ^ f_s_pg_rca24_or22;
  assign f_s_pg_rca24_and23 = f_s_pg_rca24_or22 & f_s_pg_rca24_pg_fa23_xor0;
  assign f_s_pg_rca24_or23 = f_s_pg_rca24_and23 | f_s_pg_rca24_pg_fa23_and0;
  assign f_s_pg_rca24_xor0 = a[23] ^ b[23];
  assign f_s_pg_rca24_xor1 = f_s_pg_rca24_xor0 ^ f_s_pg_rca24_or23;

  assign f_s_pg_rca24_out[0] = f_s_pg_rca24_pg_fa0_xor0;
  assign f_s_pg_rca24_out[1] = f_s_pg_rca24_pg_fa1_xor1;
  assign f_s_pg_rca24_out[2] = f_s_pg_rca24_pg_fa2_xor1;
  assign f_s_pg_rca24_out[3] = f_s_pg_rca24_pg_fa3_xor1;
  assign f_s_pg_rca24_out[4] = f_s_pg_rca24_pg_fa4_xor1;
  assign f_s_pg_rca24_out[5] = f_s_pg_rca24_pg_fa5_xor1;
  assign f_s_pg_rca24_out[6] = f_s_pg_rca24_pg_fa6_xor1;
  assign f_s_pg_rca24_out[7] = f_s_pg_rca24_pg_fa7_xor1;
  assign f_s_pg_rca24_out[8] = f_s_pg_rca24_pg_fa8_xor1;
  assign f_s_pg_rca24_out[9] = f_s_pg_rca24_pg_fa9_xor1;
  assign f_s_pg_rca24_out[10] = f_s_pg_rca24_pg_fa10_xor1;
  assign f_s_pg_rca24_out[11] = f_s_pg_rca24_pg_fa11_xor1;
  assign f_s_pg_rca24_out[12] = f_s_pg_rca24_pg_fa12_xor1;
  assign f_s_pg_rca24_out[13] = f_s_pg_rca24_pg_fa13_xor1;
  assign f_s_pg_rca24_out[14] = f_s_pg_rca24_pg_fa14_xor1;
  assign f_s_pg_rca24_out[15] = f_s_pg_rca24_pg_fa15_xor1;
  assign f_s_pg_rca24_out[16] = f_s_pg_rca24_pg_fa16_xor1;
  assign f_s_pg_rca24_out[17] = f_s_pg_rca24_pg_fa17_xor1;
  assign f_s_pg_rca24_out[18] = f_s_pg_rca24_pg_fa18_xor1;
  assign f_s_pg_rca24_out[19] = f_s_pg_rca24_pg_fa19_xor1;
  assign f_s_pg_rca24_out[20] = f_s_pg_rca24_pg_fa20_xor1;
  assign f_s_pg_rca24_out[21] = f_s_pg_rca24_pg_fa21_xor1;
  assign f_s_pg_rca24_out[22] = f_s_pg_rca24_pg_fa22_xor1;
  assign f_s_pg_rca24_out[23] = f_s_pg_rca24_pg_fa23_xor1;
  assign f_s_pg_rca24_out[24] = f_s_pg_rca24_xor1;
endmodule