module f_u_cska4(input [3:0] a, input [3:0] b, output [4:0] f_u_cska4_out);
  wire f_u_cska4_xor0;
  wire f_u_cska4_ha0_xor0;
  wire f_u_cska4_ha0_and0;
  wire f_u_cska4_xor1;
  wire f_u_cska4_fa0_xor0;
  wire f_u_cska4_fa0_and0;
  wire f_u_cska4_fa0_xor1;
  wire f_u_cska4_fa0_and1;
  wire f_u_cska4_fa0_or0;
  wire f_u_cska4_xor2;
  wire f_u_cska4_fa1_xor0;
  wire f_u_cska4_fa1_and0;
  wire f_u_cska4_fa1_xor1;
  wire f_u_cska4_fa1_and1;
  wire f_u_cska4_fa1_or0;
  wire f_u_cska4_xor3;
  wire f_u_cska4_fa2_xor0;
  wire f_u_cska4_fa2_and0;
  wire f_u_cska4_fa2_xor1;
  wire f_u_cska4_fa2_and1;
  wire f_u_cska4_fa2_or0;
  wire f_u_cska4_and_propagate00;
  wire f_u_cska4_and_propagate01;
  wire f_u_cska4_and_propagate02;
  wire f_u_cska4_mux2to10_not0;
  wire f_u_cska4_mux2to10_and1;

  assign f_u_cska4_xor0 = a[0] ^ b[0];
  assign f_u_cska4_ha0_xor0 = a[0] ^ b[0];
  assign f_u_cska4_ha0_and0 = a[0] & b[0];
  assign f_u_cska4_xor1 = a[1] ^ b[1];
  assign f_u_cska4_fa0_xor0 = a[1] ^ b[1];
  assign f_u_cska4_fa0_and0 = a[1] & b[1];
  assign f_u_cska4_fa0_xor1 = f_u_cska4_fa0_xor0 ^ f_u_cska4_ha0_and0;
  assign f_u_cska4_fa0_and1 = f_u_cska4_fa0_xor0 & f_u_cska4_ha0_and0;
  assign f_u_cska4_fa0_or0 = f_u_cska4_fa0_and0 | f_u_cska4_fa0_and1;
  assign f_u_cska4_xor2 = a[2] ^ b[2];
  assign f_u_cska4_fa1_xor0 = a[2] ^ b[2];
  assign f_u_cska4_fa1_and0 = a[2] & b[2];
  assign f_u_cska4_fa1_xor1 = f_u_cska4_fa1_xor0 ^ f_u_cska4_fa0_or0;
  assign f_u_cska4_fa1_and1 = f_u_cska4_fa1_xor0 & f_u_cska4_fa0_or0;
  assign f_u_cska4_fa1_or0 = f_u_cska4_fa1_and0 | f_u_cska4_fa1_and1;
  assign f_u_cska4_xor3 = a[3] ^ b[3];
  assign f_u_cska4_fa2_xor0 = a[3] ^ b[3];
  assign f_u_cska4_fa2_and0 = a[3] & b[3];
  assign f_u_cska4_fa2_xor1 = f_u_cska4_fa2_xor0 ^ f_u_cska4_fa1_or0;
  assign f_u_cska4_fa2_and1 = f_u_cska4_fa2_xor0 & f_u_cska4_fa1_or0;
  assign f_u_cska4_fa2_or0 = f_u_cska4_fa2_and0 | f_u_cska4_fa2_and1;
  assign f_u_cska4_and_propagate00 = f_u_cska4_xor0 & f_u_cska4_xor2;
  assign f_u_cska4_and_propagate01 = f_u_cska4_xor1 & f_u_cska4_xor3;
  assign f_u_cska4_and_propagate02 = f_u_cska4_and_propagate00 & f_u_cska4_and_propagate01;
  assign f_u_cska4_mux2to10_not0 = ~f_u_cska4_and_propagate02;
  assign f_u_cska4_mux2to10_and1 = f_u_cska4_fa2_or0 & f_u_cska4_mux2to10_not0;

  assign f_u_cska4_out[0] = f_u_cska4_ha0_xor0;
  assign f_u_cska4_out[1] = f_u_cska4_fa0_xor1;
  assign f_u_cska4_out[2] = f_u_cska4_fa1_xor1;
  assign f_u_cska4_out[3] = f_u_cska4_fa2_xor1;
  assign f_u_cska4_out[4] = f_u_cska4_mux2to10_and1;
endmodule