module f_u_cla8(input [7:0] a, input [7:0] b, output [8:0] f_u_cla8_out);
  wire f_u_cla8_pg_logic0_or0;
  wire f_u_cla8_pg_logic0_and0;
  wire f_u_cla8_pg_logic0_xor0;
  wire f_u_cla8_pg_logic1_or0;
  wire f_u_cla8_pg_logic1_and0;
  wire f_u_cla8_pg_logic1_xor0;
  wire f_u_cla8_xor1;
  wire f_u_cla8_and0;
  wire f_u_cla8_or0;
  wire f_u_cla8_pg_logic2_or0;
  wire f_u_cla8_pg_logic2_and0;
  wire f_u_cla8_pg_logic2_xor0;
  wire f_u_cla8_xor2;
  wire f_u_cla8_and1;
  wire f_u_cla8_and2;
  wire f_u_cla8_and3;
  wire f_u_cla8_and4;
  wire f_u_cla8_or1;
  wire f_u_cla8_or2;
  wire f_u_cla8_pg_logic3_or0;
  wire f_u_cla8_pg_logic3_and0;
  wire f_u_cla8_pg_logic3_xor0;
  wire f_u_cla8_xor3;
  wire f_u_cla8_and5;
  wire f_u_cla8_and6;
  wire f_u_cla8_and7;
  wire f_u_cla8_and8;
  wire f_u_cla8_and9;
  wire f_u_cla8_and10;
  wire f_u_cla8_and11;
  wire f_u_cla8_or3;
  wire f_u_cla8_or4;
  wire f_u_cla8_or5;
  wire f_u_cla8_pg_logic4_or0;
  wire f_u_cla8_pg_logic4_and0;
  wire f_u_cla8_pg_logic4_xor0;
  wire f_u_cla8_xor4;
  wire f_u_cla8_and12;
  wire f_u_cla8_or6;
  wire f_u_cla8_pg_logic5_or0;
  wire f_u_cla8_pg_logic5_and0;
  wire f_u_cla8_pg_logic5_xor0;
  wire f_u_cla8_xor5;
  wire f_u_cla8_and13;
  wire f_u_cla8_and14;
  wire f_u_cla8_and15;
  wire f_u_cla8_or7;
  wire f_u_cla8_or8;
  wire f_u_cla8_pg_logic6_or0;
  wire f_u_cla8_pg_logic6_and0;
  wire f_u_cla8_pg_logic6_xor0;
  wire f_u_cla8_xor6;
  wire f_u_cla8_and16;
  wire f_u_cla8_and17;
  wire f_u_cla8_and18;
  wire f_u_cla8_and19;
  wire f_u_cla8_and20;
  wire f_u_cla8_and21;
  wire f_u_cla8_or9;
  wire f_u_cla8_or10;
  wire f_u_cla8_or11;
  wire f_u_cla8_pg_logic7_or0;
  wire f_u_cla8_pg_logic7_and0;
  wire f_u_cla8_pg_logic7_xor0;
  wire f_u_cla8_xor7;
  wire f_u_cla8_and22;
  wire f_u_cla8_and23;
  wire f_u_cla8_and24;
  wire f_u_cla8_and25;
  wire f_u_cla8_and26;
  wire f_u_cla8_and27;
  wire f_u_cla8_and28;
  wire f_u_cla8_and29;
  wire f_u_cla8_and30;
  wire f_u_cla8_and31;
  wire f_u_cla8_or12;
  wire f_u_cla8_or13;
  wire f_u_cla8_or14;
  wire f_u_cla8_or15;

  assign f_u_cla8_pg_logic0_or0 = a[0] | b[0];
  assign f_u_cla8_pg_logic0_and0 = a[0] & b[0];
  assign f_u_cla8_pg_logic0_xor0 = a[0] ^ b[0];
  assign f_u_cla8_pg_logic1_or0 = a[1] | b[1];
  assign f_u_cla8_pg_logic1_and0 = a[1] & b[1];
  assign f_u_cla8_pg_logic1_xor0 = a[1] ^ b[1];
  assign f_u_cla8_xor1 = f_u_cla8_pg_logic1_xor0 ^ f_u_cla8_pg_logic0_and0;
  assign f_u_cla8_and0 = f_u_cla8_pg_logic0_and0 & f_u_cla8_pg_logic1_or0;
  assign f_u_cla8_or0 = f_u_cla8_pg_logic1_and0 | f_u_cla8_and0;
  assign f_u_cla8_pg_logic2_or0 = a[2] | b[2];
  assign f_u_cla8_pg_logic2_and0 = a[2] & b[2];
  assign f_u_cla8_pg_logic2_xor0 = a[2] ^ b[2];
  assign f_u_cla8_xor2 = f_u_cla8_pg_logic2_xor0 ^ f_u_cla8_or0;
  assign f_u_cla8_and1 = f_u_cla8_pg_logic2_or0 & f_u_cla8_pg_logic0_or0;
  assign f_u_cla8_and2 = f_u_cla8_pg_logic0_and0 & f_u_cla8_pg_logic2_or0;
  assign f_u_cla8_and3 = f_u_cla8_and2 & f_u_cla8_pg_logic1_or0;
  assign f_u_cla8_and4 = f_u_cla8_pg_logic1_and0 & f_u_cla8_pg_logic2_or0;
  assign f_u_cla8_or1 = f_u_cla8_and3 | f_u_cla8_and4;
  assign f_u_cla8_or2 = f_u_cla8_pg_logic2_and0 | f_u_cla8_or1;
  assign f_u_cla8_pg_logic3_or0 = a[3] | b[3];
  assign f_u_cla8_pg_logic3_and0 = a[3] & b[3];
  assign f_u_cla8_pg_logic3_xor0 = a[3] ^ b[3];
  assign f_u_cla8_xor3 = f_u_cla8_pg_logic3_xor0 ^ f_u_cla8_or2;
  assign f_u_cla8_and5 = f_u_cla8_pg_logic3_or0 & f_u_cla8_pg_logic1_or0;
  assign f_u_cla8_and6 = f_u_cla8_pg_logic0_and0 & f_u_cla8_pg_logic2_or0;
  assign f_u_cla8_and7 = f_u_cla8_pg_logic3_or0 & f_u_cla8_pg_logic1_or0;
  assign f_u_cla8_and8 = f_u_cla8_and6 & f_u_cla8_and7;
  assign f_u_cla8_and9 = f_u_cla8_pg_logic1_and0 & f_u_cla8_pg_logic3_or0;
  assign f_u_cla8_and10 = f_u_cla8_and9 & f_u_cla8_pg_logic2_or0;
  assign f_u_cla8_and11 = f_u_cla8_pg_logic2_and0 & f_u_cla8_pg_logic3_or0;
  assign f_u_cla8_or3 = f_u_cla8_and8 | f_u_cla8_and11;
  assign f_u_cla8_or4 = f_u_cla8_and10 | f_u_cla8_or3;
  assign f_u_cla8_or5 = f_u_cla8_pg_logic3_and0 | f_u_cla8_or4;
  assign f_u_cla8_pg_logic4_or0 = a[4] | b[4];
  assign f_u_cla8_pg_logic4_and0 = a[4] & b[4];
  assign f_u_cla8_pg_logic4_xor0 = a[4] ^ b[4];
  assign f_u_cla8_xor4 = f_u_cla8_pg_logic4_xor0 ^ f_u_cla8_or5;
  assign f_u_cla8_and12 = f_u_cla8_or5 & f_u_cla8_pg_logic4_or0;
  assign f_u_cla8_or6 = f_u_cla8_pg_logic4_and0 | f_u_cla8_and12;
  assign f_u_cla8_pg_logic5_or0 = a[5] | b[5];
  assign f_u_cla8_pg_logic5_and0 = a[5] & b[5];
  assign f_u_cla8_pg_logic5_xor0 = a[5] ^ b[5];
  assign f_u_cla8_xor5 = f_u_cla8_pg_logic5_xor0 ^ f_u_cla8_or6;
  assign f_u_cla8_and13 = f_u_cla8_or5 & f_u_cla8_pg_logic5_or0;
  assign f_u_cla8_and14 = f_u_cla8_and13 & f_u_cla8_pg_logic4_or0;
  assign f_u_cla8_and15 = f_u_cla8_pg_logic4_and0 & f_u_cla8_pg_logic5_or0;
  assign f_u_cla8_or7 = f_u_cla8_and14 | f_u_cla8_and15;
  assign f_u_cla8_or8 = f_u_cla8_pg_logic5_and0 | f_u_cla8_or7;
  assign f_u_cla8_pg_logic6_or0 = a[6] | b[6];
  assign f_u_cla8_pg_logic6_and0 = a[6] & b[6];
  assign f_u_cla8_pg_logic6_xor0 = a[6] ^ b[6];
  assign f_u_cla8_xor6 = f_u_cla8_pg_logic6_xor0 ^ f_u_cla8_or8;
  assign f_u_cla8_and16 = f_u_cla8_or5 & f_u_cla8_pg_logic5_or0;
  assign f_u_cla8_and17 = f_u_cla8_pg_logic6_or0 & f_u_cla8_pg_logic4_or0;
  assign f_u_cla8_and18 = f_u_cla8_and16 & f_u_cla8_and17;
  assign f_u_cla8_and19 = f_u_cla8_pg_logic4_and0 & f_u_cla8_pg_logic6_or0;
  assign f_u_cla8_and20 = f_u_cla8_and19 & f_u_cla8_pg_logic5_or0;
  assign f_u_cla8_and21 = f_u_cla8_pg_logic5_and0 & f_u_cla8_pg_logic6_or0;
  assign f_u_cla8_or9 = f_u_cla8_and18 | f_u_cla8_and20;
  assign f_u_cla8_or10 = f_u_cla8_or9 | f_u_cla8_and21;
  assign f_u_cla8_or11 = f_u_cla8_pg_logic6_and0 | f_u_cla8_or10;
  assign f_u_cla8_pg_logic7_or0 = a[7] | b[7];
  assign f_u_cla8_pg_logic7_and0 = a[7] & b[7];
  assign f_u_cla8_pg_logic7_xor0 = a[7] ^ b[7];
  assign f_u_cla8_xor7 = f_u_cla8_pg_logic7_xor0 ^ f_u_cla8_or11;
  assign f_u_cla8_and22 = f_u_cla8_or5 & f_u_cla8_pg_logic6_or0;
  assign f_u_cla8_and23 = f_u_cla8_pg_logic7_or0 & f_u_cla8_pg_logic5_or0;
  assign f_u_cla8_and24 = f_u_cla8_and22 & f_u_cla8_and23;
  assign f_u_cla8_and25 = f_u_cla8_and24 & f_u_cla8_pg_logic4_or0;
  assign f_u_cla8_and26 = f_u_cla8_pg_logic4_and0 & f_u_cla8_pg_logic6_or0;
  assign f_u_cla8_and27 = f_u_cla8_pg_logic7_or0 & f_u_cla8_pg_logic5_or0;
  assign f_u_cla8_and28 = f_u_cla8_and26 & f_u_cla8_and27;
  assign f_u_cla8_and29 = f_u_cla8_pg_logic5_and0 & f_u_cla8_pg_logic7_or0;
  assign f_u_cla8_and30 = f_u_cla8_and29 & f_u_cla8_pg_logic6_or0;
  assign f_u_cla8_and31 = f_u_cla8_pg_logic6_and0 & f_u_cla8_pg_logic7_or0;
  assign f_u_cla8_or12 = f_u_cla8_and25 | f_u_cla8_and30;
  assign f_u_cla8_or13 = f_u_cla8_and28 | f_u_cla8_and31;
  assign f_u_cla8_or14 = f_u_cla8_or12 | f_u_cla8_or13;
  assign f_u_cla8_or15 = f_u_cla8_pg_logic7_and0 | f_u_cla8_or14;

  assign f_u_cla8_out[0] = f_u_cla8_pg_logic0_xor0;
  assign f_u_cla8_out[1] = f_u_cla8_xor1;
  assign f_u_cla8_out[2] = f_u_cla8_xor2;
  assign f_u_cla8_out[3] = f_u_cla8_xor3;
  assign f_u_cla8_out[4] = f_u_cla8_xor4;
  assign f_u_cla8_out[5] = f_u_cla8_xor5;
  assign f_u_cla8_out[6] = f_u_cla8_xor6;
  assign f_u_cla8_out[7] = f_u_cla8_xor7;
  assign f_u_cla8_out[8] = f_u_cla8_or15;
endmodule