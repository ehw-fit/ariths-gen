module u_pg_rca16(input [15:0] a, input [15:0] b, output [16:0] u_pg_rca16_out);
  wire u_pg_rca16_pg_fa0_xor0;
  wire u_pg_rca16_pg_fa0_and0;
  wire u_pg_rca16_pg_fa1_xor0;
  wire u_pg_rca16_pg_fa1_and0;
  wire u_pg_rca16_pg_fa1_xor1;
  wire u_pg_rca16_and1;
  wire u_pg_rca16_or1;
  wire u_pg_rca16_pg_fa2_xor0;
  wire u_pg_rca16_pg_fa2_and0;
  wire u_pg_rca16_pg_fa2_xor1;
  wire u_pg_rca16_and2;
  wire u_pg_rca16_or2;
  wire u_pg_rca16_pg_fa3_xor0;
  wire u_pg_rca16_pg_fa3_and0;
  wire u_pg_rca16_pg_fa3_xor1;
  wire u_pg_rca16_and3;
  wire u_pg_rca16_or3;
  wire u_pg_rca16_pg_fa4_xor0;
  wire u_pg_rca16_pg_fa4_and0;
  wire u_pg_rca16_pg_fa4_xor1;
  wire u_pg_rca16_and4;
  wire u_pg_rca16_or4;
  wire u_pg_rca16_pg_fa5_xor0;
  wire u_pg_rca16_pg_fa5_and0;
  wire u_pg_rca16_pg_fa5_xor1;
  wire u_pg_rca16_and5;
  wire u_pg_rca16_or5;
  wire u_pg_rca16_pg_fa6_xor0;
  wire u_pg_rca16_pg_fa6_and0;
  wire u_pg_rca16_pg_fa6_xor1;
  wire u_pg_rca16_and6;
  wire u_pg_rca16_or6;
  wire u_pg_rca16_pg_fa7_xor0;
  wire u_pg_rca16_pg_fa7_and0;
  wire u_pg_rca16_pg_fa7_xor1;
  wire u_pg_rca16_and7;
  wire u_pg_rca16_or7;
  wire u_pg_rca16_pg_fa8_xor0;
  wire u_pg_rca16_pg_fa8_and0;
  wire u_pg_rca16_pg_fa8_xor1;
  wire u_pg_rca16_and8;
  wire u_pg_rca16_or8;
  wire u_pg_rca16_pg_fa9_xor0;
  wire u_pg_rca16_pg_fa9_and0;
  wire u_pg_rca16_pg_fa9_xor1;
  wire u_pg_rca16_and9;
  wire u_pg_rca16_or9;
  wire u_pg_rca16_pg_fa10_xor0;
  wire u_pg_rca16_pg_fa10_and0;
  wire u_pg_rca16_pg_fa10_xor1;
  wire u_pg_rca16_and10;
  wire u_pg_rca16_or10;
  wire u_pg_rca16_pg_fa11_xor0;
  wire u_pg_rca16_pg_fa11_and0;
  wire u_pg_rca16_pg_fa11_xor1;
  wire u_pg_rca16_and11;
  wire u_pg_rca16_or11;
  wire u_pg_rca16_pg_fa12_xor0;
  wire u_pg_rca16_pg_fa12_and0;
  wire u_pg_rca16_pg_fa12_xor1;
  wire u_pg_rca16_and12;
  wire u_pg_rca16_or12;
  wire u_pg_rca16_pg_fa13_xor0;
  wire u_pg_rca16_pg_fa13_and0;
  wire u_pg_rca16_pg_fa13_xor1;
  wire u_pg_rca16_and13;
  wire u_pg_rca16_or13;
  wire u_pg_rca16_pg_fa14_xor0;
  wire u_pg_rca16_pg_fa14_and0;
  wire u_pg_rca16_pg_fa14_xor1;
  wire u_pg_rca16_and14;
  wire u_pg_rca16_or14;
  wire u_pg_rca16_pg_fa15_xor0;
  wire u_pg_rca16_pg_fa15_and0;
  wire u_pg_rca16_pg_fa15_xor1;
  wire u_pg_rca16_and15;
  wire u_pg_rca16_or15;

  assign u_pg_rca16_pg_fa0_xor0 = a[0] ^ b[0];
  assign u_pg_rca16_pg_fa0_and0 = a[0] & b[0];
  assign u_pg_rca16_pg_fa1_xor0 = a[1] ^ b[1];
  assign u_pg_rca16_pg_fa1_and0 = a[1] & b[1];
  assign u_pg_rca16_pg_fa1_xor1 = u_pg_rca16_pg_fa1_xor0 ^ u_pg_rca16_pg_fa0_and0;
  assign u_pg_rca16_and1 = u_pg_rca16_pg_fa0_and0 & u_pg_rca16_pg_fa1_xor0;
  assign u_pg_rca16_or1 = u_pg_rca16_and1 | u_pg_rca16_pg_fa1_and0;
  assign u_pg_rca16_pg_fa2_xor0 = a[2] ^ b[2];
  assign u_pg_rca16_pg_fa2_and0 = a[2] & b[2];
  assign u_pg_rca16_pg_fa2_xor1 = u_pg_rca16_pg_fa2_xor0 ^ u_pg_rca16_or1;
  assign u_pg_rca16_and2 = u_pg_rca16_or1 & u_pg_rca16_pg_fa2_xor0;
  assign u_pg_rca16_or2 = u_pg_rca16_and2 | u_pg_rca16_pg_fa2_and0;
  assign u_pg_rca16_pg_fa3_xor0 = a[3] ^ b[3];
  assign u_pg_rca16_pg_fa3_and0 = a[3] & b[3];
  assign u_pg_rca16_pg_fa3_xor1 = u_pg_rca16_pg_fa3_xor0 ^ u_pg_rca16_or2;
  assign u_pg_rca16_and3 = u_pg_rca16_or2 & u_pg_rca16_pg_fa3_xor0;
  assign u_pg_rca16_or3 = u_pg_rca16_and3 | u_pg_rca16_pg_fa3_and0;
  assign u_pg_rca16_pg_fa4_xor0 = a[4] ^ b[4];
  assign u_pg_rca16_pg_fa4_and0 = a[4] & b[4];
  assign u_pg_rca16_pg_fa4_xor1 = u_pg_rca16_pg_fa4_xor0 ^ u_pg_rca16_or3;
  assign u_pg_rca16_and4 = u_pg_rca16_or3 & u_pg_rca16_pg_fa4_xor0;
  assign u_pg_rca16_or4 = u_pg_rca16_and4 | u_pg_rca16_pg_fa4_and0;
  assign u_pg_rca16_pg_fa5_xor0 = a[5] ^ b[5];
  assign u_pg_rca16_pg_fa5_and0 = a[5] & b[5];
  assign u_pg_rca16_pg_fa5_xor1 = u_pg_rca16_pg_fa5_xor0 ^ u_pg_rca16_or4;
  assign u_pg_rca16_and5 = u_pg_rca16_or4 & u_pg_rca16_pg_fa5_xor0;
  assign u_pg_rca16_or5 = u_pg_rca16_and5 | u_pg_rca16_pg_fa5_and0;
  assign u_pg_rca16_pg_fa6_xor0 = a[6] ^ b[6];
  assign u_pg_rca16_pg_fa6_and0 = a[6] & b[6];
  assign u_pg_rca16_pg_fa6_xor1 = u_pg_rca16_pg_fa6_xor0 ^ u_pg_rca16_or5;
  assign u_pg_rca16_and6 = u_pg_rca16_or5 & u_pg_rca16_pg_fa6_xor0;
  assign u_pg_rca16_or6 = u_pg_rca16_and6 | u_pg_rca16_pg_fa6_and0;
  assign u_pg_rca16_pg_fa7_xor0 = a[7] ^ b[7];
  assign u_pg_rca16_pg_fa7_and0 = a[7] & b[7];
  assign u_pg_rca16_pg_fa7_xor1 = u_pg_rca16_pg_fa7_xor0 ^ u_pg_rca16_or6;
  assign u_pg_rca16_and7 = u_pg_rca16_or6 & u_pg_rca16_pg_fa7_xor0;
  assign u_pg_rca16_or7 = u_pg_rca16_and7 | u_pg_rca16_pg_fa7_and0;
  assign u_pg_rca16_pg_fa8_xor0 = a[8] ^ b[8];
  assign u_pg_rca16_pg_fa8_and0 = a[8] & b[8];
  assign u_pg_rca16_pg_fa8_xor1 = u_pg_rca16_pg_fa8_xor0 ^ u_pg_rca16_or7;
  assign u_pg_rca16_and8 = u_pg_rca16_or7 & u_pg_rca16_pg_fa8_xor0;
  assign u_pg_rca16_or8 = u_pg_rca16_and8 | u_pg_rca16_pg_fa8_and0;
  assign u_pg_rca16_pg_fa9_xor0 = a[9] ^ b[9];
  assign u_pg_rca16_pg_fa9_and0 = a[9] & b[9];
  assign u_pg_rca16_pg_fa9_xor1 = u_pg_rca16_pg_fa9_xor0 ^ u_pg_rca16_or8;
  assign u_pg_rca16_and9 = u_pg_rca16_or8 & u_pg_rca16_pg_fa9_xor0;
  assign u_pg_rca16_or9 = u_pg_rca16_and9 | u_pg_rca16_pg_fa9_and0;
  assign u_pg_rca16_pg_fa10_xor0 = a[10] ^ b[10];
  assign u_pg_rca16_pg_fa10_and0 = a[10] & b[10];
  assign u_pg_rca16_pg_fa10_xor1 = u_pg_rca16_pg_fa10_xor0 ^ u_pg_rca16_or9;
  assign u_pg_rca16_and10 = u_pg_rca16_or9 & u_pg_rca16_pg_fa10_xor0;
  assign u_pg_rca16_or10 = u_pg_rca16_and10 | u_pg_rca16_pg_fa10_and0;
  assign u_pg_rca16_pg_fa11_xor0 = a[11] ^ b[11];
  assign u_pg_rca16_pg_fa11_and0 = a[11] & b[11];
  assign u_pg_rca16_pg_fa11_xor1 = u_pg_rca16_pg_fa11_xor0 ^ u_pg_rca16_or10;
  assign u_pg_rca16_and11 = u_pg_rca16_or10 & u_pg_rca16_pg_fa11_xor0;
  assign u_pg_rca16_or11 = u_pg_rca16_and11 | u_pg_rca16_pg_fa11_and0;
  assign u_pg_rca16_pg_fa12_xor0 = a[12] ^ b[12];
  assign u_pg_rca16_pg_fa12_and0 = a[12] & b[12];
  assign u_pg_rca16_pg_fa12_xor1 = u_pg_rca16_pg_fa12_xor0 ^ u_pg_rca16_or11;
  assign u_pg_rca16_and12 = u_pg_rca16_or11 & u_pg_rca16_pg_fa12_xor0;
  assign u_pg_rca16_or12 = u_pg_rca16_and12 | u_pg_rca16_pg_fa12_and0;
  assign u_pg_rca16_pg_fa13_xor0 = a[13] ^ b[13];
  assign u_pg_rca16_pg_fa13_and0 = a[13] & b[13];
  assign u_pg_rca16_pg_fa13_xor1 = u_pg_rca16_pg_fa13_xor0 ^ u_pg_rca16_or12;
  assign u_pg_rca16_and13 = u_pg_rca16_or12 & u_pg_rca16_pg_fa13_xor0;
  assign u_pg_rca16_or13 = u_pg_rca16_and13 | u_pg_rca16_pg_fa13_and0;
  assign u_pg_rca16_pg_fa14_xor0 = a[14] ^ b[14];
  assign u_pg_rca16_pg_fa14_and0 = a[14] & b[14];
  assign u_pg_rca16_pg_fa14_xor1 = u_pg_rca16_pg_fa14_xor0 ^ u_pg_rca16_or13;
  assign u_pg_rca16_and14 = u_pg_rca16_or13 & u_pg_rca16_pg_fa14_xor0;
  assign u_pg_rca16_or14 = u_pg_rca16_and14 | u_pg_rca16_pg_fa14_and0;
  assign u_pg_rca16_pg_fa15_xor0 = a[15] ^ b[15];
  assign u_pg_rca16_pg_fa15_and0 = a[15] & b[15];
  assign u_pg_rca16_pg_fa15_xor1 = u_pg_rca16_pg_fa15_xor0 ^ u_pg_rca16_or14;
  assign u_pg_rca16_and15 = u_pg_rca16_or14 & u_pg_rca16_pg_fa15_xor0;
  assign u_pg_rca16_or15 = u_pg_rca16_and15 | u_pg_rca16_pg_fa15_and0;

  assign u_pg_rca16_out[0] = u_pg_rca16_pg_fa0_xor0;
  assign u_pg_rca16_out[1] = u_pg_rca16_pg_fa1_xor1;
  assign u_pg_rca16_out[2] = u_pg_rca16_pg_fa2_xor1;
  assign u_pg_rca16_out[3] = u_pg_rca16_pg_fa3_xor1;
  assign u_pg_rca16_out[4] = u_pg_rca16_pg_fa4_xor1;
  assign u_pg_rca16_out[5] = u_pg_rca16_pg_fa5_xor1;
  assign u_pg_rca16_out[6] = u_pg_rca16_pg_fa6_xor1;
  assign u_pg_rca16_out[7] = u_pg_rca16_pg_fa7_xor1;
  assign u_pg_rca16_out[8] = u_pg_rca16_pg_fa8_xor1;
  assign u_pg_rca16_out[9] = u_pg_rca16_pg_fa9_xor1;
  assign u_pg_rca16_out[10] = u_pg_rca16_pg_fa10_xor1;
  assign u_pg_rca16_out[11] = u_pg_rca16_pg_fa11_xor1;
  assign u_pg_rca16_out[12] = u_pg_rca16_pg_fa12_xor1;
  assign u_pg_rca16_out[13] = u_pg_rca16_pg_fa13_xor1;
  assign u_pg_rca16_out[14] = u_pg_rca16_pg_fa14_xor1;
  assign u_pg_rca16_out[15] = u_pg_rca16_pg_fa15_xor1;
  assign u_pg_rca16_out[16] = u_pg_rca16_or15;
endmodule