module s_pg_rca32(input [31:0] a, input [31:0] b, output [32:0] s_pg_rca32_out);
  wire s_pg_rca32_pg_fa0_xor0;
  wire s_pg_rca32_pg_fa0_and0;
  wire s_pg_rca32_pg_fa1_xor0;
  wire s_pg_rca32_pg_fa1_and0;
  wire s_pg_rca32_pg_fa1_xor1;
  wire s_pg_rca32_and1;
  wire s_pg_rca32_or1;
  wire s_pg_rca32_pg_fa2_xor0;
  wire s_pg_rca32_pg_fa2_and0;
  wire s_pg_rca32_pg_fa2_xor1;
  wire s_pg_rca32_and2;
  wire s_pg_rca32_or2;
  wire s_pg_rca32_pg_fa3_xor0;
  wire s_pg_rca32_pg_fa3_and0;
  wire s_pg_rca32_pg_fa3_xor1;
  wire s_pg_rca32_and3;
  wire s_pg_rca32_or3;
  wire s_pg_rca32_pg_fa4_xor0;
  wire s_pg_rca32_pg_fa4_and0;
  wire s_pg_rca32_pg_fa4_xor1;
  wire s_pg_rca32_and4;
  wire s_pg_rca32_or4;
  wire s_pg_rca32_pg_fa5_xor0;
  wire s_pg_rca32_pg_fa5_and0;
  wire s_pg_rca32_pg_fa5_xor1;
  wire s_pg_rca32_and5;
  wire s_pg_rca32_or5;
  wire s_pg_rca32_pg_fa6_xor0;
  wire s_pg_rca32_pg_fa6_and0;
  wire s_pg_rca32_pg_fa6_xor1;
  wire s_pg_rca32_and6;
  wire s_pg_rca32_or6;
  wire s_pg_rca32_pg_fa7_xor0;
  wire s_pg_rca32_pg_fa7_and0;
  wire s_pg_rca32_pg_fa7_xor1;
  wire s_pg_rca32_and7;
  wire s_pg_rca32_or7;
  wire s_pg_rca32_pg_fa8_xor0;
  wire s_pg_rca32_pg_fa8_and0;
  wire s_pg_rca32_pg_fa8_xor1;
  wire s_pg_rca32_and8;
  wire s_pg_rca32_or8;
  wire s_pg_rca32_pg_fa9_xor0;
  wire s_pg_rca32_pg_fa9_and0;
  wire s_pg_rca32_pg_fa9_xor1;
  wire s_pg_rca32_and9;
  wire s_pg_rca32_or9;
  wire s_pg_rca32_pg_fa10_xor0;
  wire s_pg_rca32_pg_fa10_and0;
  wire s_pg_rca32_pg_fa10_xor1;
  wire s_pg_rca32_and10;
  wire s_pg_rca32_or10;
  wire s_pg_rca32_pg_fa11_xor0;
  wire s_pg_rca32_pg_fa11_and0;
  wire s_pg_rca32_pg_fa11_xor1;
  wire s_pg_rca32_and11;
  wire s_pg_rca32_or11;
  wire s_pg_rca32_pg_fa12_xor0;
  wire s_pg_rca32_pg_fa12_and0;
  wire s_pg_rca32_pg_fa12_xor1;
  wire s_pg_rca32_and12;
  wire s_pg_rca32_or12;
  wire s_pg_rca32_pg_fa13_xor0;
  wire s_pg_rca32_pg_fa13_and0;
  wire s_pg_rca32_pg_fa13_xor1;
  wire s_pg_rca32_and13;
  wire s_pg_rca32_or13;
  wire s_pg_rca32_pg_fa14_xor0;
  wire s_pg_rca32_pg_fa14_and0;
  wire s_pg_rca32_pg_fa14_xor1;
  wire s_pg_rca32_and14;
  wire s_pg_rca32_or14;
  wire s_pg_rca32_pg_fa15_xor0;
  wire s_pg_rca32_pg_fa15_and0;
  wire s_pg_rca32_pg_fa15_xor1;
  wire s_pg_rca32_and15;
  wire s_pg_rca32_or15;
  wire s_pg_rca32_pg_fa16_xor0;
  wire s_pg_rca32_pg_fa16_and0;
  wire s_pg_rca32_pg_fa16_xor1;
  wire s_pg_rca32_and16;
  wire s_pg_rca32_or16;
  wire s_pg_rca32_pg_fa17_xor0;
  wire s_pg_rca32_pg_fa17_and0;
  wire s_pg_rca32_pg_fa17_xor1;
  wire s_pg_rca32_and17;
  wire s_pg_rca32_or17;
  wire s_pg_rca32_pg_fa18_xor0;
  wire s_pg_rca32_pg_fa18_and0;
  wire s_pg_rca32_pg_fa18_xor1;
  wire s_pg_rca32_and18;
  wire s_pg_rca32_or18;
  wire s_pg_rca32_pg_fa19_xor0;
  wire s_pg_rca32_pg_fa19_and0;
  wire s_pg_rca32_pg_fa19_xor1;
  wire s_pg_rca32_and19;
  wire s_pg_rca32_or19;
  wire s_pg_rca32_pg_fa20_xor0;
  wire s_pg_rca32_pg_fa20_and0;
  wire s_pg_rca32_pg_fa20_xor1;
  wire s_pg_rca32_and20;
  wire s_pg_rca32_or20;
  wire s_pg_rca32_pg_fa21_xor0;
  wire s_pg_rca32_pg_fa21_and0;
  wire s_pg_rca32_pg_fa21_xor1;
  wire s_pg_rca32_and21;
  wire s_pg_rca32_or21;
  wire s_pg_rca32_pg_fa22_xor0;
  wire s_pg_rca32_pg_fa22_and0;
  wire s_pg_rca32_pg_fa22_xor1;
  wire s_pg_rca32_and22;
  wire s_pg_rca32_or22;
  wire s_pg_rca32_pg_fa23_xor0;
  wire s_pg_rca32_pg_fa23_and0;
  wire s_pg_rca32_pg_fa23_xor1;
  wire s_pg_rca32_and23;
  wire s_pg_rca32_or23;
  wire s_pg_rca32_pg_fa24_xor0;
  wire s_pg_rca32_pg_fa24_and0;
  wire s_pg_rca32_pg_fa24_xor1;
  wire s_pg_rca32_and24;
  wire s_pg_rca32_or24;
  wire s_pg_rca32_pg_fa25_xor0;
  wire s_pg_rca32_pg_fa25_and0;
  wire s_pg_rca32_pg_fa25_xor1;
  wire s_pg_rca32_and25;
  wire s_pg_rca32_or25;
  wire s_pg_rca32_pg_fa26_xor0;
  wire s_pg_rca32_pg_fa26_and0;
  wire s_pg_rca32_pg_fa26_xor1;
  wire s_pg_rca32_and26;
  wire s_pg_rca32_or26;
  wire s_pg_rca32_pg_fa27_xor0;
  wire s_pg_rca32_pg_fa27_and0;
  wire s_pg_rca32_pg_fa27_xor1;
  wire s_pg_rca32_and27;
  wire s_pg_rca32_or27;
  wire s_pg_rca32_pg_fa28_xor0;
  wire s_pg_rca32_pg_fa28_and0;
  wire s_pg_rca32_pg_fa28_xor1;
  wire s_pg_rca32_and28;
  wire s_pg_rca32_or28;
  wire s_pg_rca32_pg_fa29_xor0;
  wire s_pg_rca32_pg_fa29_and0;
  wire s_pg_rca32_pg_fa29_xor1;
  wire s_pg_rca32_and29;
  wire s_pg_rca32_or29;
  wire s_pg_rca32_pg_fa30_xor0;
  wire s_pg_rca32_pg_fa30_and0;
  wire s_pg_rca32_pg_fa30_xor1;
  wire s_pg_rca32_and30;
  wire s_pg_rca32_or30;
  wire s_pg_rca32_pg_fa31_xor0;
  wire s_pg_rca32_pg_fa31_and0;
  wire s_pg_rca32_pg_fa31_xor1;
  wire s_pg_rca32_and31;
  wire s_pg_rca32_or31;
  wire s_pg_rca32_xor0;
  wire s_pg_rca32_xor1;

  assign s_pg_rca32_pg_fa0_xor0 = a[0] ^ b[0];
  assign s_pg_rca32_pg_fa0_and0 = a[0] & b[0];
  assign s_pg_rca32_pg_fa1_xor0 = a[1] ^ b[1];
  assign s_pg_rca32_pg_fa1_and0 = a[1] & b[1];
  assign s_pg_rca32_pg_fa1_xor1 = s_pg_rca32_pg_fa1_xor0 ^ s_pg_rca32_pg_fa0_and0;
  assign s_pg_rca32_and1 = s_pg_rca32_pg_fa0_and0 & s_pg_rca32_pg_fa1_xor0;
  assign s_pg_rca32_or1 = s_pg_rca32_and1 | s_pg_rca32_pg_fa1_and0;
  assign s_pg_rca32_pg_fa2_xor0 = a[2] ^ b[2];
  assign s_pg_rca32_pg_fa2_and0 = a[2] & b[2];
  assign s_pg_rca32_pg_fa2_xor1 = s_pg_rca32_pg_fa2_xor0 ^ s_pg_rca32_or1;
  assign s_pg_rca32_and2 = s_pg_rca32_or1 & s_pg_rca32_pg_fa2_xor0;
  assign s_pg_rca32_or2 = s_pg_rca32_and2 | s_pg_rca32_pg_fa2_and0;
  assign s_pg_rca32_pg_fa3_xor0 = a[3] ^ b[3];
  assign s_pg_rca32_pg_fa3_and0 = a[3] & b[3];
  assign s_pg_rca32_pg_fa3_xor1 = s_pg_rca32_pg_fa3_xor0 ^ s_pg_rca32_or2;
  assign s_pg_rca32_and3 = s_pg_rca32_or2 & s_pg_rca32_pg_fa3_xor0;
  assign s_pg_rca32_or3 = s_pg_rca32_and3 | s_pg_rca32_pg_fa3_and0;
  assign s_pg_rca32_pg_fa4_xor0 = a[4] ^ b[4];
  assign s_pg_rca32_pg_fa4_and0 = a[4] & b[4];
  assign s_pg_rca32_pg_fa4_xor1 = s_pg_rca32_pg_fa4_xor0 ^ s_pg_rca32_or3;
  assign s_pg_rca32_and4 = s_pg_rca32_or3 & s_pg_rca32_pg_fa4_xor0;
  assign s_pg_rca32_or4 = s_pg_rca32_and4 | s_pg_rca32_pg_fa4_and0;
  assign s_pg_rca32_pg_fa5_xor0 = a[5] ^ b[5];
  assign s_pg_rca32_pg_fa5_and0 = a[5] & b[5];
  assign s_pg_rca32_pg_fa5_xor1 = s_pg_rca32_pg_fa5_xor0 ^ s_pg_rca32_or4;
  assign s_pg_rca32_and5 = s_pg_rca32_or4 & s_pg_rca32_pg_fa5_xor0;
  assign s_pg_rca32_or5 = s_pg_rca32_and5 | s_pg_rca32_pg_fa5_and0;
  assign s_pg_rca32_pg_fa6_xor0 = a[6] ^ b[6];
  assign s_pg_rca32_pg_fa6_and0 = a[6] & b[6];
  assign s_pg_rca32_pg_fa6_xor1 = s_pg_rca32_pg_fa6_xor0 ^ s_pg_rca32_or5;
  assign s_pg_rca32_and6 = s_pg_rca32_or5 & s_pg_rca32_pg_fa6_xor0;
  assign s_pg_rca32_or6 = s_pg_rca32_and6 | s_pg_rca32_pg_fa6_and0;
  assign s_pg_rca32_pg_fa7_xor0 = a[7] ^ b[7];
  assign s_pg_rca32_pg_fa7_and0 = a[7] & b[7];
  assign s_pg_rca32_pg_fa7_xor1 = s_pg_rca32_pg_fa7_xor0 ^ s_pg_rca32_or6;
  assign s_pg_rca32_and7 = s_pg_rca32_or6 & s_pg_rca32_pg_fa7_xor0;
  assign s_pg_rca32_or7 = s_pg_rca32_and7 | s_pg_rca32_pg_fa7_and0;
  assign s_pg_rca32_pg_fa8_xor0 = a[8] ^ b[8];
  assign s_pg_rca32_pg_fa8_and0 = a[8] & b[8];
  assign s_pg_rca32_pg_fa8_xor1 = s_pg_rca32_pg_fa8_xor0 ^ s_pg_rca32_or7;
  assign s_pg_rca32_and8 = s_pg_rca32_or7 & s_pg_rca32_pg_fa8_xor0;
  assign s_pg_rca32_or8 = s_pg_rca32_and8 | s_pg_rca32_pg_fa8_and0;
  assign s_pg_rca32_pg_fa9_xor0 = a[9] ^ b[9];
  assign s_pg_rca32_pg_fa9_and0 = a[9] & b[9];
  assign s_pg_rca32_pg_fa9_xor1 = s_pg_rca32_pg_fa9_xor0 ^ s_pg_rca32_or8;
  assign s_pg_rca32_and9 = s_pg_rca32_or8 & s_pg_rca32_pg_fa9_xor0;
  assign s_pg_rca32_or9 = s_pg_rca32_and9 | s_pg_rca32_pg_fa9_and0;
  assign s_pg_rca32_pg_fa10_xor0 = a[10] ^ b[10];
  assign s_pg_rca32_pg_fa10_and0 = a[10] & b[10];
  assign s_pg_rca32_pg_fa10_xor1 = s_pg_rca32_pg_fa10_xor0 ^ s_pg_rca32_or9;
  assign s_pg_rca32_and10 = s_pg_rca32_or9 & s_pg_rca32_pg_fa10_xor0;
  assign s_pg_rca32_or10 = s_pg_rca32_and10 | s_pg_rca32_pg_fa10_and0;
  assign s_pg_rca32_pg_fa11_xor0 = a[11] ^ b[11];
  assign s_pg_rca32_pg_fa11_and0 = a[11] & b[11];
  assign s_pg_rca32_pg_fa11_xor1 = s_pg_rca32_pg_fa11_xor0 ^ s_pg_rca32_or10;
  assign s_pg_rca32_and11 = s_pg_rca32_or10 & s_pg_rca32_pg_fa11_xor0;
  assign s_pg_rca32_or11 = s_pg_rca32_and11 | s_pg_rca32_pg_fa11_and0;
  assign s_pg_rca32_pg_fa12_xor0 = a[12] ^ b[12];
  assign s_pg_rca32_pg_fa12_and0 = a[12] & b[12];
  assign s_pg_rca32_pg_fa12_xor1 = s_pg_rca32_pg_fa12_xor0 ^ s_pg_rca32_or11;
  assign s_pg_rca32_and12 = s_pg_rca32_or11 & s_pg_rca32_pg_fa12_xor0;
  assign s_pg_rca32_or12 = s_pg_rca32_and12 | s_pg_rca32_pg_fa12_and0;
  assign s_pg_rca32_pg_fa13_xor0 = a[13] ^ b[13];
  assign s_pg_rca32_pg_fa13_and0 = a[13] & b[13];
  assign s_pg_rca32_pg_fa13_xor1 = s_pg_rca32_pg_fa13_xor0 ^ s_pg_rca32_or12;
  assign s_pg_rca32_and13 = s_pg_rca32_or12 & s_pg_rca32_pg_fa13_xor0;
  assign s_pg_rca32_or13 = s_pg_rca32_and13 | s_pg_rca32_pg_fa13_and0;
  assign s_pg_rca32_pg_fa14_xor0 = a[14] ^ b[14];
  assign s_pg_rca32_pg_fa14_and0 = a[14] & b[14];
  assign s_pg_rca32_pg_fa14_xor1 = s_pg_rca32_pg_fa14_xor0 ^ s_pg_rca32_or13;
  assign s_pg_rca32_and14 = s_pg_rca32_or13 & s_pg_rca32_pg_fa14_xor0;
  assign s_pg_rca32_or14 = s_pg_rca32_and14 | s_pg_rca32_pg_fa14_and0;
  assign s_pg_rca32_pg_fa15_xor0 = a[15] ^ b[15];
  assign s_pg_rca32_pg_fa15_and0 = a[15] & b[15];
  assign s_pg_rca32_pg_fa15_xor1 = s_pg_rca32_pg_fa15_xor0 ^ s_pg_rca32_or14;
  assign s_pg_rca32_and15 = s_pg_rca32_or14 & s_pg_rca32_pg_fa15_xor0;
  assign s_pg_rca32_or15 = s_pg_rca32_and15 | s_pg_rca32_pg_fa15_and0;
  assign s_pg_rca32_pg_fa16_xor0 = a[16] ^ b[16];
  assign s_pg_rca32_pg_fa16_and0 = a[16] & b[16];
  assign s_pg_rca32_pg_fa16_xor1 = s_pg_rca32_pg_fa16_xor0 ^ s_pg_rca32_or15;
  assign s_pg_rca32_and16 = s_pg_rca32_or15 & s_pg_rca32_pg_fa16_xor0;
  assign s_pg_rca32_or16 = s_pg_rca32_and16 | s_pg_rca32_pg_fa16_and0;
  assign s_pg_rca32_pg_fa17_xor0 = a[17] ^ b[17];
  assign s_pg_rca32_pg_fa17_and0 = a[17] & b[17];
  assign s_pg_rca32_pg_fa17_xor1 = s_pg_rca32_pg_fa17_xor0 ^ s_pg_rca32_or16;
  assign s_pg_rca32_and17 = s_pg_rca32_or16 & s_pg_rca32_pg_fa17_xor0;
  assign s_pg_rca32_or17 = s_pg_rca32_and17 | s_pg_rca32_pg_fa17_and0;
  assign s_pg_rca32_pg_fa18_xor0 = a[18] ^ b[18];
  assign s_pg_rca32_pg_fa18_and0 = a[18] & b[18];
  assign s_pg_rca32_pg_fa18_xor1 = s_pg_rca32_pg_fa18_xor0 ^ s_pg_rca32_or17;
  assign s_pg_rca32_and18 = s_pg_rca32_or17 & s_pg_rca32_pg_fa18_xor0;
  assign s_pg_rca32_or18 = s_pg_rca32_and18 | s_pg_rca32_pg_fa18_and0;
  assign s_pg_rca32_pg_fa19_xor0 = a[19] ^ b[19];
  assign s_pg_rca32_pg_fa19_and0 = a[19] & b[19];
  assign s_pg_rca32_pg_fa19_xor1 = s_pg_rca32_pg_fa19_xor0 ^ s_pg_rca32_or18;
  assign s_pg_rca32_and19 = s_pg_rca32_or18 & s_pg_rca32_pg_fa19_xor0;
  assign s_pg_rca32_or19 = s_pg_rca32_and19 | s_pg_rca32_pg_fa19_and0;
  assign s_pg_rca32_pg_fa20_xor0 = a[20] ^ b[20];
  assign s_pg_rca32_pg_fa20_and0 = a[20] & b[20];
  assign s_pg_rca32_pg_fa20_xor1 = s_pg_rca32_pg_fa20_xor0 ^ s_pg_rca32_or19;
  assign s_pg_rca32_and20 = s_pg_rca32_or19 & s_pg_rca32_pg_fa20_xor0;
  assign s_pg_rca32_or20 = s_pg_rca32_and20 | s_pg_rca32_pg_fa20_and0;
  assign s_pg_rca32_pg_fa21_xor0 = a[21] ^ b[21];
  assign s_pg_rca32_pg_fa21_and0 = a[21] & b[21];
  assign s_pg_rca32_pg_fa21_xor1 = s_pg_rca32_pg_fa21_xor0 ^ s_pg_rca32_or20;
  assign s_pg_rca32_and21 = s_pg_rca32_or20 & s_pg_rca32_pg_fa21_xor0;
  assign s_pg_rca32_or21 = s_pg_rca32_and21 | s_pg_rca32_pg_fa21_and0;
  assign s_pg_rca32_pg_fa22_xor0 = a[22] ^ b[22];
  assign s_pg_rca32_pg_fa22_and0 = a[22] & b[22];
  assign s_pg_rca32_pg_fa22_xor1 = s_pg_rca32_pg_fa22_xor0 ^ s_pg_rca32_or21;
  assign s_pg_rca32_and22 = s_pg_rca32_or21 & s_pg_rca32_pg_fa22_xor0;
  assign s_pg_rca32_or22 = s_pg_rca32_and22 | s_pg_rca32_pg_fa22_and0;
  assign s_pg_rca32_pg_fa23_xor0 = a[23] ^ b[23];
  assign s_pg_rca32_pg_fa23_and0 = a[23] & b[23];
  assign s_pg_rca32_pg_fa23_xor1 = s_pg_rca32_pg_fa23_xor0 ^ s_pg_rca32_or22;
  assign s_pg_rca32_and23 = s_pg_rca32_or22 & s_pg_rca32_pg_fa23_xor0;
  assign s_pg_rca32_or23 = s_pg_rca32_and23 | s_pg_rca32_pg_fa23_and0;
  assign s_pg_rca32_pg_fa24_xor0 = a[24] ^ b[24];
  assign s_pg_rca32_pg_fa24_and0 = a[24] & b[24];
  assign s_pg_rca32_pg_fa24_xor1 = s_pg_rca32_pg_fa24_xor0 ^ s_pg_rca32_or23;
  assign s_pg_rca32_and24 = s_pg_rca32_or23 & s_pg_rca32_pg_fa24_xor0;
  assign s_pg_rca32_or24 = s_pg_rca32_and24 | s_pg_rca32_pg_fa24_and0;
  assign s_pg_rca32_pg_fa25_xor0 = a[25] ^ b[25];
  assign s_pg_rca32_pg_fa25_and0 = a[25] & b[25];
  assign s_pg_rca32_pg_fa25_xor1 = s_pg_rca32_pg_fa25_xor0 ^ s_pg_rca32_or24;
  assign s_pg_rca32_and25 = s_pg_rca32_or24 & s_pg_rca32_pg_fa25_xor0;
  assign s_pg_rca32_or25 = s_pg_rca32_and25 | s_pg_rca32_pg_fa25_and0;
  assign s_pg_rca32_pg_fa26_xor0 = a[26] ^ b[26];
  assign s_pg_rca32_pg_fa26_and0 = a[26] & b[26];
  assign s_pg_rca32_pg_fa26_xor1 = s_pg_rca32_pg_fa26_xor0 ^ s_pg_rca32_or25;
  assign s_pg_rca32_and26 = s_pg_rca32_or25 & s_pg_rca32_pg_fa26_xor0;
  assign s_pg_rca32_or26 = s_pg_rca32_and26 | s_pg_rca32_pg_fa26_and0;
  assign s_pg_rca32_pg_fa27_xor0 = a[27] ^ b[27];
  assign s_pg_rca32_pg_fa27_and0 = a[27] & b[27];
  assign s_pg_rca32_pg_fa27_xor1 = s_pg_rca32_pg_fa27_xor0 ^ s_pg_rca32_or26;
  assign s_pg_rca32_and27 = s_pg_rca32_or26 & s_pg_rca32_pg_fa27_xor0;
  assign s_pg_rca32_or27 = s_pg_rca32_and27 | s_pg_rca32_pg_fa27_and0;
  assign s_pg_rca32_pg_fa28_xor0 = a[28] ^ b[28];
  assign s_pg_rca32_pg_fa28_and0 = a[28] & b[28];
  assign s_pg_rca32_pg_fa28_xor1 = s_pg_rca32_pg_fa28_xor0 ^ s_pg_rca32_or27;
  assign s_pg_rca32_and28 = s_pg_rca32_or27 & s_pg_rca32_pg_fa28_xor0;
  assign s_pg_rca32_or28 = s_pg_rca32_and28 | s_pg_rca32_pg_fa28_and0;
  assign s_pg_rca32_pg_fa29_xor0 = a[29] ^ b[29];
  assign s_pg_rca32_pg_fa29_and0 = a[29] & b[29];
  assign s_pg_rca32_pg_fa29_xor1 = s_pg_rca32_pg_fa29_xor0 ^ s_pg_rca32_or28;
  assign s_pg_rca32_and29 = s_pg_rca32_or28 & s_pg_rca32_pg_fa29_xor0;
  assign s_pg_rca32_or29 = s_pg_rca32_and29 | s_pg_rca32_pg_fa29_and0;
  assign s_pg_rca32_pg_fa30_xor0 = a[30] ^ b[30];
  assign s_pg_rca32_pg_fa30_and0 = a[30] & b[30];
  assign s_pg_rca32_pg_fa30_xor1 = s_pg_rca32_pg_fa30_xor0 ^ s_pg_rca32_or29;
  assign s_pg_rca32_and30 = s_pg_rca32_or29 & s_pg_rca32_pg_fa30_xor0;
  assign s_pg_rca32_or30 = s_pg_rca32_and30 | s_pg_rca32_pg_fa30_and0;
  assign s_pg_rca32_pg_fa31_xor0 = a[31] ^ b[31];
  assign s_pg_rca32_pg_fa31_and0 = a[31] & b[31];
  assign s_pg_rca32_pg_fa31_xor1 = s_pg_rca32_pg_fa31_xor0 ^ s_pg_rca32_or30;
  assign s_pg_rca32_and31 = s_pg_rca32_or30 & s_pg_rca32_pg_fa31_xor0;
  assign s_pg_rca32_or31 = s_pg_rca32_and31 | s_pg_rca32_pg_fa31_and0;
  assign s_pg_rca32_xor0 = a[31] ^ b[31];
  assign s_pg_rca32_xor1 = s_pg_rca32_xor0 ^ s_pg_rca32_or31;

  assign s_pg_rca32_out[0] = s_pg_rca32_pg_fa0_xor0;
  assign s_pg_rca32_out[1] = s_pg_rca32_pg_fa1_xor1;
  assign s_pg_rca32_out[2] = s_pg_rca32_pg_fa2_xor1;
  assign s_pg_rca32_out[3] = s_pg_rca32_pg_fa3_xor1;
  assign s_pg_rca32_out[4] = s_pg_rca32_pg_fa4_xor1;
  assign s_pg_rca32_out[5] = s_pg_rca32_pg_fa5_xor1;
  assign s_pg_rca32_out[6] = s_pg_rca32_pg_fa6_xor1;
  assign s_pg_rca32_out[7] = s_pg_rca32_pg_fa7_xor1;
  assign s_pg_rca32_out[8] = s_pg_rca32_pg_fa8_xor1;
  assign s_pg_rca32_out[9] = s_pg_rca32_pg_fa9_xor1;
  assign s_pg_rca32_out[10] = s_pg_rca32_pg_fa10_xor1;
  assign s_pg_rca32_out[11] = s_pg_rca32_pg_fa11_xor1;
  assign s_pg_rca32_out[12] = s_pg_rca32_pg_fa12_xor1;
  assign s_pg_rca32_out[13] = s_pg_rca32_pg_fa13_xor1;
  assign s_pg_rca32_out[14] = s_pg_rca32_pg_fa14_xor1;
  assign s_pg_rca32_out[15] = s_pg_rca32_pg_fa15_xor1;
  assign s_pg_rca32_out[16] = s_pg_rca32_pg_fa16_xor1;
  assign s_pg_rca32_out[17] = s_pg_rca32_pg_fa17_xor1;
  assign s_pg_rca32_out[18] = s_pg_rca32_pg_fa18_xor1;
  assign s_pg_rca32_out[19] = s_pg_rca32_pg_fa19_xor1;
  assign s_pg_rca32_out[20] = s_pg_rca32_pg_fa20_xor1;
  assign s_pg_rca32_out[21] = s_pg_rca32_pg_fa21_xor1;
  assign s_pg_rca32_out[22] = s_pg_rca32_pg_fa22_xor1;
  assign s_pg_rca32_out[23] = s_pg_rca32_pg_fa23_xor1;
  assign s_pg_rca32_out[24] = s_pg_rca32_pg_fa24_xor1;
  assign s_pg_rca32_out[25] = s_pg_rca32_pg_fa25_xor1;
  assign s_pg_rca32_out[26] = s_pg_rca32_pg_fa26_xor1;
  assign s_pg_rca32_out[27] = s_pg_rca32_pg_fa27_xor1;
  assign s_pg_rca32_out[28] = s_pg_rca32_pg_fa28_xor1;
  assign s_pg_rca32_out[29] = s_pg_rca32_pg_fa29_xor1;
  assign s_pg_rca32_out[30] = s_pg_rca32_pg_fa30_xor1;
  assign s_pg_rca32_out[31] = s_pg_rca32_pg_fa31_xor1;
  assign s_pg_rca32_out[32] = s_pg_rca32_xor1;
endmodule