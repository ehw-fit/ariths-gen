module u_CSAwallace_cska4(input [3:0] a, input [3:0] b, output [7:0] u_CSAwallace_cska4_out);
  wire u_CSAwallace_cska4_and_0_0;
  wire u_CSAwallace_cska4_and_1_0;
  wire u_CSAwallace_cska4_and_2_0;
  wire u_CSAwallace_cska4_and_3_0;
  wire u_CSAwallace_cska4_and_0_1;
  wire u_CSAwallace_cska4_and_1_1;
  wire u_CSAwallace_cska4_and_2_1;
  wire u_CSAwallace_cska4_and_3_1;
  wire u_CSAwallace_cska4_and_0_2;
  wire u_CSAwallace_cska4_and_1_2;
  wire u_CSAwallace_cska4_and_2_2;
  wire u_CSAwallace_cska4_and_3_2;
  wire u_CSAwallace_cska4_and_0_3;
  wire u_CSAwallace_cska4_and_1_3;
  wire u_CSAwallace_cska4_and_2_3;
  wire u_CSAwallace_cska4_and_3_3;
  wire u_CSAwallace_cska4_csa0_csa_component_fa1_xor0;
  wire u_CSAwallace_cska4_csa0_csa_component_fa1_and0;
  wire u_CSAwallace_cska4_csa0_csa_component_fa2_xor0;
  wire u_CSAwallace_cska4_csa0_csa_component_fa2_and0;
  wire u_CSAwallace_cska4_csa0_csa_component_fa2_xor1;
  wire u_CSAwallace_cska4_csa0_csa_component_fa2_and1;
  wire u_CSAwallace_cska4_csa0_csa_component_fa2_or0;
  wire u_CSAwallace_cska4_csa0_csa_component_fa3_xor0;
  wire u_CSAwallace_cska4_csa0_csa_component_fa3_and0;
  wire u_CSAwallace_cska4_csa0_csa_component_fa3_xor1;
  wire u_CSAwallace_cska4_csa0_csa_component_fa3_and1;
  wire u_CSAwallace_cska4_csa0_csa_component_fa3_or0;
  wire u_CSAwallace_cska4_csa0_csa_component_fa4_xor1;
  wire u_CSAwallace_cska4_csa0_csa_component_fa4_and1;
  wire u_CSAwallace_cska4_csa1_csa_component_fa2_xor0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa2_and0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa3_xor0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa3_and0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa3_xor1;
  wire u_CSAwallace_cska4_csa1_csa_component_fa3_and1;
  wire u_CSAwallace_cska4_csa1_csa_component_fa3_or0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa4_xor0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa4_and0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa4_xor1;
  wire u_CSAwallace_cska4_csa1_csa_component_fa4_and1;
  wire u_CSAwallace_cska4_csa1_csa_component_fa4_or0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa5_xor0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa5_and0;
  wire u_CSAwallace_cska4_csa1_csa_component_fa5_xor1;
  wire u_CSAwallace_cska4_csa1_csa_component_fa5_and1;
  wire u_CSAwallace_cska4_csa1_csa_component_fa5_or0;
  wire u_CSAwallace_cska4_u_cska8_xor3;
  wire u_CSAwallace_cska4_u_cska8_fa2_xor0;
  wire u_CSAwallace_cska4_u_cska8_fa2_and0;
  wire u_CSAwallace_cska4_u_cska8_and_propagate00;
  wire u_CSAwallace_cska4_u_cska8_and_propagate01;
  wire u_CSAwallace_cska4_u_cska8_and_propagate02;
  wire u_CSAwallace_cska4_u_cska8_mux2to10_not0;
  wire u_CSAwallace_cska4_u_cska8_mux2to10_and1;
  wire u_CSAwallace_cska4_u_cska8_xor4;
  wire u_CSAwallace_cska4_u_cska8_fa3_xor0;
  wire u_CSAwallace_cska4_u_cska8_fa3_and0;
  wire u_CSAwallace_cska4_u_cska8_fa3_xor1;
  wire u_CSAwallace_cska4_u_cska8_fa3_and1;
  wire u_CSAwallace_cska4_u_cska8_fa3_or0;
  wire u_CSAwallace_cska4_u_cska8_xor5;
  wire u_CSAwallace_cska4_u_cska8_fa4_xor0;
  wire u_CSAwallace_cska4_u_cska8_fa4_and0;
  wire u_CSAwallace_cska4_u_cska8_fa4_xor1;
  wire u_CSAwallace_cska4_u_cska8_fa4_and1;
  wire u_CSAwallace_cska4_u_cska8_fa4_or0;
  wire u_CSAwallace_cska4_u_cska8_xor6;
  wire u_CSAwallace_cska4_u_cska8_fa5_xor0;
  wire u_CSAwallace_cska4_u_cska8_fa5_and0;
  wire u_CSAwallace_cska4_u_cska8_fa5_xor1;
  wire u_CSAwallace_cska4_u_cska8_fa5_and1;
  wire u_CSAwallace_cska4_u_cska8_fa5_or0;
  wire u_CSAwallace_cska4_u_cska8_and_propagate13;

  assign u_CSAwallace_cska4_and_0_0 = a[0] & b[0];
  assign u_CSAwallace_cska4_and_1_0 = a[1] & b[0];
  assign u_CSAwallace_cska4_and_2_0 = a[2] & b[0];
  assign u_CSAwallace_cska4_and_3_0 = a[3] & b[0];
  assign u_CSAwallace_cska4_and_0_1 = a[0] & b[1];
  assign u_CSAwallace_cska4_and_1_1 = a[1] & b[1];
  assign u_CSAwallace_cska4_and_2_1 = a[2] & b[1];
  assign u_CSAwallace_cska4_and_3_1 = a[3] & b[1];
  assign u_CSAwallace_cska4_and_0_2 = a[0] & b[2];
  assign u_CSAwallace_cska4_and_1_2 = a[1] & b[2];
  assign u_CSAwallace_cska4_and_2_2 = a[2] & b[2];
  assign u_CSAwallace_cska4_and_3_2 = a[3] & b[2];
  assign u_CSAwallace_cska4_and_0_3 = a[0] & b[3];
  assign u_CSAwallace_cska4_and_1_3 = a[1] & b[3];
  assign u_CSAwallace_cska4_and_2_3 = a[2] & b[3];
  assign u_CSAwallace_cska4_and_3_3 = a[3] & b[3];
  assign u_CSAwallace_cska4_csa0_csa_component_fa1_xor0 = u_CSAwallace_cska4_and_1_0 ^ u_CSAwallace_cska4_and_0_1;
  assign u_CSAwallace_cska4_csa0_csa_component_fa1_and0 = u_CSAwallace_cska4_and_1_0 & u_CSAwallace_cska4_and_0_1;
  assign u_CSAwallace_cska4_csa0_csa_component_fa2_xor0 = u_CSAwallace_cska4_and_2_0 ^ u_CSAwallace_cska4_and_1_1;
  assign u_CSAwallace_cska4_csa0_csa_component_fa2_and0 = u_CSAwallace_cska4_and_2_0 & u_CSAwallace_cska4_and_1_1;
  assign u_CSAwallace_cska4_csa0_csa_component_fa2_xor1 = u_CSAwallace_cska4_csa0_csa_component_fa2_xor0 ^ u_CSAwallace_cska4_and_0_2;
  assign u_CSAwallace_cska4_csa0_csa_component_fa2_and1 = u_CSAwallace_cska4_csa0_csa_component_fa2_xor0 & u_CSAwallace_cska4_and_0_2;
  assign u_CSAwallace_cska4_csa0_csa_component_fa2_or0 = u_CSAwallace_cska4_csa0_csa_component_fa2_and0 | u_CSAwallace_cska4_csa0_csa_component_fa2_and1;
  assign u_CSAwallace_cska4_csa0_csa_component_fa3_xor0 = u_CSAwallace_cska4_and_3_0 ^ u_CSAwallace_cska4_and_2_1;
  assign u_CSAwallace_cska4_csa0_csa_component_fa3_and0 = u_CSAwallace_cska4_and_3_0 & u_CSAwallace_cska4_and_2_1;
  assign u_CSAwallace_cska4_csa0_csa_component_fa3_xor1 = u_CSAwallace_cska4_csa0_csa_component_fa3_xor0 ^ u_CSAwallace_cska4_and_1_2;
  assign u_CSAwallace_cska4_csa0_csa_component_fa3_and1 = u_CSAwallace_cska4_csa0_csa_component_fa3_xor0 & u_CSAwallace_cska4_and_1_2;
  assign u_CSAwallace_cska4_csa0_csa_component_fa3_or0 = u_CSAwallace_cska4_csa0_csa_component_fa3_and0 | u_CSAwallace_cska4_csa0_csa_component_fa3_and1;
  assign u_CSAwallace_cska4_csa0_csa_component_fa4_xor1 = u_CSAwallace_cska4_and_3_1 ^ u_CSAwallace_cska4_and_2_2;
  assign u_CSAwallace_cska4_csa0_csa_component_fa4_and1 = u_CSAwallace_cska4_and_3_1 & u_CSAwallace_cska4_and_2_2;
  assign u_CSAwallace_cska4_csa1_csa_component_fa2_xor0 = u_CSAwallace_cska4_csa0_csa_component_fa2_xor1 ^ u_CSAwallace_cska4_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_cska4_csa1_csa_component_fa2_and0 = u_CSAwallace_cska4_csa0_csa_component_fa2_xor1 & u_CSAwallace_cska4_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_cska4_csa1_csa_component_fa3_xor0 = u_CSAwallace_cska4_csa0_csa_component_fa3_xor1 ^ u_CSAwallace_cska4_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_cska4_csa1_csa_component_fa3_and0 = u_CSAwallace_cska4_csa0_csa_component_fa3_xor1 & u_CSAwallace_cska4_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_cska4_csa1_csa_component_fa3_xor1 = u_CSAwallace_cska4_csa1_csa_component_fa3_xor0 ^ u_CSAwallace_cska4_and_0_3;
  assign u_CSAwallace_cska4_csa1_csa_component_fa3_and1 = u_CSAwallace_cska4_csa1_csa_component_fa3_xor0 & u_CSAwallace_cska4_and_0_3;
  assign u_CSAwallace_cska4_csa1_csa_component_fa3_or0 = u_CSAwallace_cska4_csa1_csa_component_fa3_and0 | u_CSAwallace_cska4_csa1_csa_component_fa3_and1;
  assign u_CSAwallace_cska4_csa1_csa_component_fa4_xor0 = u_CSAwallace_cska4_csa0_csa_component_fa4_xor1 ^ u_CSAwallace_cska4_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_cska4_csa1_csa_component_fa4_and0 = u_CSAwallace_cska4_csa0_csa_component_fa4_xor1 & u_CSAwallace_cska4_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_cska4_csa1_csa_component_fa4_xor1 = u_CSAwallace_cska4_csa1_csa_component_fa4_xor0 ^ u_CSAwallace_cska4_and_1_3;
  assign u_CSAwallace_cska4_csa1_csa_component_fa4_and1 = u_CSAwallace_cska4_csa1_csa_component_fa4_xor0 & u_CSAwallace_cska4_and_1_3;
  assign u_CSAwallace_cska4_csa1_csa_component_fa4_or0 = u_CSAwallace_cska4_csa1_csa_component_fa4_and0 | u_CSAwallace_cska4_csa1_csa_component_fa4_and1;
  assign u_CSAwallace_cska4_csa1_csa_component_fa5_xor0 = u_CSAwallace_cska4_and_3_2 ^ u_CSAwallace_cska4_csa0_csa_component_fa4_and1;
  assign u_CSAwallace_cska4_csa1_csa_component_fa5_and0 = u_CSAwallace_cska4_and_3_2 & u_CSAwallace_cska4_csa0_csa_component_fa4_and1;
  assign u_CSAwallace_cska4_csa1_csa_component_fa5_xor1 = u_CSAwallace_cska4_csa1_csa_component_fa5_xor0 ^ u_CSAwallace_cska4_and_2_3;
  assign u_CSAwallace_cska4_csa1_csa_component_fa5_and1 = u_CSAwallace_cska4_csa1_csa_component_fa5_xor0 & u_CSAwallace_cska4_and_2_3;
  assign u_CSAwallace_cska4_csa1_csa_component_fa5_or0 = u_CSAwallace_cska4_csa1_csa_component_fa5_and0 | u_CSAwallace_cska4_csa1_csa_component_fa5_and1;
  assign u_CSAwallace_cska4_u_cska8_xor3 = u_CSAwallace_cska4_csa1_csa_component_fa3_xor1 ^ u_CSAwallace_cska4_csa1_csa_component_fa2_and0;
  assign u_CSAwallace_cska4_u_cska8_fa2_xor0 = u_CSAwallace_cska4_csa1_csa_component_fa3_xor1 ^ u_CSAwallace_cska4_csa1_csa_component_fa2_and0;
  assign u_CSAwallace_cska4_u_cska8_fa2_and0 = u_CSAwallace_cska4_csa1_csa_component_fa3_xor1 & u_CSAwallace_cska4_csa1_csa_component_fa2_and0;
  assign u_CSAwallace_cska4_u_cska8_and_propagate00 = u_CSAwallace_cska4_and_0_0 & u_CSAwallace_cska4_csa1_csa_component_fa2_xor0;
  assign u_CSAwallace_cska4_u_cska8_and_propagate01 = u_CSAwallace_cska4_csa0_csa_component_fa1_xor0 & u_CSAwallace_cska4_u_cska8_xor3;
  assign u_CSAwallace_cska4_u_cska8_and_propagate02 = u_CSAwallace_cska4_u_cska8_and_propagate00 & u_CSAwallace_cska4_u_cska8_and_propagate01;
  assign u_CSAwallace_cska4_u_cska8_mux2to10_not0 = ~u_CSAwallace_cska4_u_cska8_and_propagate02;
  assign u_CSAwallace_cska4_u_cska8_mux2to10_and1 = u_CSAwallace_cska4_u_cska8_fa2_and0 & u_CSAwallace_cska4_u_cska8_mux2to10_not0;
  assign u_CSAwallace_cska4_u_cska8_xor4 = u_CSAwallace_cska4_csa1_csa_component_fa4_xor1 ^ u_CSAwallace_cska4_csa1_csa_component_fa3_or0;
  assign u_CSAwallace_cska4_u_cska8_fa3_xor0 = u_CSAwallace_cska4_csa1_csa_component_fa4_xor1 ^ u_CSAwallace_cska4_csa1_csa_component_fa3_or0;
  assign u_CSAwallace_cska4_u_cska8_fa3_and0 = u_CSAwallace_cska4_csa1_csa_component_fa4_xor1 & u_CSAwallace_cska4_csa1_csa_component_fa3_or0;
  assign u_CSAwallace_cska4_u_cska8_fa3_xor1 = u_CSAwallace_cska4_u_cska8_fa3_xor0 ^ u_CSAwallace_cska4_u_cska8_mux2to10_and1;
  assign u_CSAwallace_cska4_u_cska8_fa3_and1 = u_CSAwallace_cska4_u_cska8_fa3_xor0 & u_CSAwallace_cska4_u_cska8_mux2to10_and1;
  assign u_CSAwallace_cska4_u_cska8_fa3_or0 = u_CSAwallace_cska4_u_cska8_fa3_and0 | u_CSAwallace_cska4_u_cska8_fa3_and1;
  assign u_CSAwallace_cska4_u_cska8_xor5 = u_CSAwallace_cska4_csa1_csa_component_fa5_xor1 ^ u_CSAwallace_cska4_csa1_csa_component_fa4_or0;
  assign u_CSAwallace_cska4_u_cska8_fa4_xor0 = u_CSAwallace_cska4_csa1_csa_component_fa5_xor1 ^ u_CSAwallace_cska4_csa1_csa_component_fa4_or0;
  assign u_CSAwallace_cska4_u_cska8_fa4_and0 = u_CSAwallace_cska4_csa1_csa_component_fa5_xor1 & u_CSAwallace_cska4_csa1_csa_component_fa4_or0;
  assign u_CSAwallace_cska4_u_cska8_fa4_xor1 = u_CSAwallace_cska4_u_cska8_fa4_xor0 ^ u_CSAwallace_cska4_u_cska8_fa3_or0;
  assign u_CSAwallace_cska4_u_cska8_fa4_and1 = u_CSAwallace_cska4_u_cska8_fa4_xor0 & u_CSAwallace_cska4_u_cska8_fa3_or0;
  assign u_CSAwallace_cska4_u_cska8_fa4_or0 = u_CSAwallace_cska4_u_cska8_fa4_and0 | u_CSAwallace_cska4_u_cska8_fa4_and1;
  assign u_CSAwallace_cska4_u_cska8_xor6 = u_CSAwallace_cska4_and_3_3 ^ u_CSAwallace_cska4_csa1_csa_component_fa5_or0;
  assign u_CSAwallace_cska4_u_cska8_fa5_xor0 = u_CSAwallace_cska4_and_3_3 ^ u_CSAwallace_cska4_csa1_csa_component_fa5_or0;
  assign u_CSAwallace_cska4_u_cska8_fa5_and0 = u_CSAwallace_cska4_and_3_3 & u_CSAwallace_cska4_csa1_csa_component_fa5_or0;
  assign u_CSAwallace_cska4_u_cska8_fa5_xor1 = u_CSAwallace_cska4_u_cska8_fa5_xor0 ^ u_CSAwallace_cska4_u_cska8_fa4_or0;
  assign u_CSAwallace_cska4_u_cska8_fa5_and1 = u_CSAwallace_cska4_u_cska8_fa5_xor0 & u_CSAwallace_cska4_u_cska8_fa4_or0;
  assign u_CSAwallace_cska4_u_cska8_fa5_or0 = u_CSAwallace_cska4_u_cska8_fa5_and0 | u_CSAwallace_cska4_u_cska8_fa5_and1;
  assign u_CSAwallace_cska4_u_cska8_and_propagate13 = u_CSAwallace_cska4_u_cska8_xor4 & u_CSAwallace_cska4_u_cska8_xor6;

  assign u_CSAwallace_cska4_out[0] = u_CSAwallace_cska4_and_0_0;
  assign u_CSAwallace_cska4_out[1] = u_CSAwallace_cska4_csa0_csa_component_fa1_xor0;
  assign u_CSAwallace_cska4_out[2] = u_CSAwallace_cska4_csa1_csa_component_fa2_xor0;
  assign u_CSAwallace_cska4_out[3] = u_CSAwallace_cska4_u_cska8_fa2_xor0;
  assign u_CSAwallace_cska4_out[4] = u_CSAwallace_cska4_u_cska8_fa3_xor1;
  assign u_CSAwallace_cska4_out[5] = u_CSAwallace_cska4_u_cska8_fa4_xor1;
  assign u_CSAwallace_cska4_out[6] = u_CSAwallace_cska4_u_cska8_fa5_xor1;
  assign u_CSAwallace_cska4_out[7] = u_CSAwallace_cska4_u_cska8_fa5_or0;
endmodule