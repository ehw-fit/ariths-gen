module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(.a(a[0]), .b(b[0]), .out(pg_logic_or0));
  and_gate and_gate_pg_logic_and0(.a(a[0]), .b(b[0]), .out(pg_logic_and0));
  xor_gate xor_gate_pg_logic_xor0(.a(a[0]), .b(b[0]), .out(pg_logic_xor0));
endmodule

module u_cla22(input [21:0] a, input [21:0] b, output [22:0] u_cla22_out);
  wire [0:0] u_cla22_pg_logic0_or0;
  wire [0:0] u_cla22_pg_logic0_and0;
  wire [0:0] u_cla22_pg_logic0_xor0;
  wire [0:0] u_cla22_pg_logic1_or0;
  wire [0:0] u_cla22_pg_logic1_and0;
  wire [0:0] u_cla22_pg_logic1_xor0;
  wire [0:0] u_cla22_xor1;
  wire [0:0] u_cla22_and0;
  wire [0:0] u_cla22_or0;
  wire [0:0] u_cla22_pg_logic2_or0;
  wire [0:0] u_cla22_pg_logic2_and0;
  wire [0:0] u_cla22_pg_logic2_xor0;
  wire [0:0] u_cla22_xor2;
  wire [0:0] u_cla22_and1;
  wire [0:0] u_cla22_and2;
  wire [0:0] u_cla22_and3;
  wire [0:0] u_cla22_and4;
  wire [0:0] u_cla22_or1;
  wire [0:0] u_cla22_or2;
  wire [0:0] u_cla22_pg_logic3_or0;
  wire [0:0] u_cla22_pg_logic3_and0;
  wire [0:0] u_cla22_pg_logic3_xor0;
  wire [0:0] u_cla22_xor3;
  wire [0:0] u_cla22_and5;
  wire [0:0] u_cla22_and6;
  wire [0:0] u_cla22_and7;
  wire [0:0] u_cla22_and8;
  wire [0:0] u_cla22_and9;
  wire [0:0] u_cla22_and10;
  wire [0:0] u_cla22_and11;
  wire [0:0] u_cla22_or3;
  wire [0:0] u_cla22_or4;
  wire [0:0] u_cla22_or5;
  wire [0:0] u_cla22_pg_logic4_or0;
  wire [0:0] u_cla22_pg_logic4_and0;
  wire [0:0] u_cla22_pg_logic4_xor0;
  wire [0:0] u_cla22_xor4;
  wire [0:0] u_cla22_and12;
  wire [0:0] u_cla22_or6;
  wire [0:0] u_cla22_pg_logic5_or0;
  wire [0:0] u_cla22_pg_logic5_and0;
  wire [0:0] u_cla22_pg_logic5_xor0;
  wire [0:0] u_cla22_xor5;
  wire [0:0] u_cla22_and13;
  wire [0:0] u_cla22_and14;
  wire [0:0] u_cla22_and15;
  wire [0:0] u_cla22_or7;
  wire [0:0] u_cla22_or8;
  wire [0:0] u_cla22_pg_logic6_or0;
  wire [0:0] u_cla22_pg_logic6_and0;
  wire [0:0] u_cla22_pg_logic6_xor0;
  wire [0:0] u_cla22_xor6;
  wire [0:0] u_cla22_and16;
  wire [0:0] u_cla22_and17;
  wire [0:0] u_cla22_and18;
  wire [0:0] u_cla22_and19;
  wire [0:0] u_cla22_and20;
  wire [0:0] u_cla22_and21;
  wire [0:0] u_cla22_or9;
  wire [0:0] u_cla22_or10;
  wire [0:0] u_cla22_or11;
  wire [0:0] u_cla22_pg_logic7_or0;
  wire [0:0] u_cla22_pg_logic7_and0;
  wire [0:0] u_cla22_pg_logic7_xor0;
  wire [0:0] u_cla22_xor7;
  wire [0:0] u_cla22_and22;
  wire [0:0] u_cla22_and23;
  wire [0:0] u_cla22_and24;
  wire [0:0] u_cla22_and25;
  wire [0:0] u_cla22_and26;
  wire [0:0] u_cla22_and27;
  wire [0:0] u_cla22_and28;
  wire [0:0] u_cla22_and29;
  wire [0:0] u_cla22_and30;
  wire [0:0] u_cla22_and31;
  wire [0:0] u_cla22_or12;
  wire [0:0] u_cla22_or13;
  wire [0:0] u_cla22_or14;
  wire [0:0] u_cla22_or15;
  wire [0:0] u_cla22_pg_logic8_or0;
  wire [0:0] u_cla22_pg_logic8_and0;
  wire [0:0] u_cla22_pg_logic8_xor0;
  wire [0:0] u_cla22_xor8;
  wire [0:0] u_cla22_and32;
  wire [0:0] u_cla22_or16;
  wire [0:0] u_cla22_pg_logic9_or0;
  wire [0:0] u_cla22_pg_logic9_and0;
  wire [0:0] u_cla22_pg_logic9_xor0;
  wire [0:0] u_cla22_xor9;
  wire [0:0] u_cla22_and33;
  wire [0:0] u_cla22_and34;
  wire [0:0] u_cla22_and35;
  wire [0:0] u_cla22_or17;
  wire [0:0] u_cla22_or18;
  wire [0:0] u_cla22_pg_logic10_or0;
  wire [0:0] u_cla22_pg_logic10_and0;
  wire [0:0] u_cla22_pg_logic10_xor0;
  wire [0:0] u_cla22_xor10;
  wire [0:0] u_cla22_and36;
  wire [0:0] u_cla22_and37;
  wire [0:0] u_cla22_and38;
  wire [0:0] u_cla22_and39;
  wire [0:0] u_cla22_and40;
  wire [0:0] u_cla22_and41;
  wire [0:0] u_cla22_or19;
  wire [0:0] u_cla22_or20;
  wire [0:0] u_cla22_or21;
  wire [0:0] u_cla22_pg_logic11_or0;
  wire [0:0] u_cla22_pg_logic11_and0;
  wire [0:0] u_cla22_pg_logic11_xor0;
  wire [0:0] u_cla22_xor11;
  wire [0:0] u_cla22_and42;
  wire [0:0] u_cla22_and43;
  wire [0:0] u_cla22_and44;
  wire [0:0] u_cla22_and45;
  wire [0:0] u_cla22_and46;
  wire [0:0] u_cla22_and47;
  wire [0:0] u_cla22_and48;
  wire [0:0] u_cla22_and49;
  wire [0:0] u_cla22_and50;
  wire [0:0] u_cla22_and51;
  wire [0:0] u_cla22_or22;
  wire [0:0] u_cla22_or23;
  wire [0:0] u_cla22_or24;
  wire [0:0] u_cla22_or25;
  wire [0:0] u_cla22_pg_logic12_or0;
  wire [0:0] u_cla22_pg_logic12_and0;
  wire [0:0] u_cla22_pg_logic12_xor0;
  wire [0:0] u_cla22_xor12;
  wire [0:0] u_cla22_and52;
  wire [0:0] u_cla22_or26;
  wire [0:0] u_cla22_pg_logic13_or0;
  wire [0:0] u_cla22_pg_logic13_and0;
  wire [0:0] u_cla22_pg_logic13_xor0;
  wire [0:0] u_cla22_xor13;
  wire [0:0] u_cla22_and53;
  wire [0:0] u_cla22_and54;
  wire [0:0] u_cla22_and55;
  wire [0:0] u_cla22_or27;
  wire [0:0] u_cla22_or28;
  wire [0:0] u_cla22_pg_logic14_or0;
  wire [0:0] u_cla22_pg_logic14_and0;
  wire [0:0] u_cla22_pg_logic14_xor0;
  wire [0:0] u_cla22_xor14;
  wire [0:0] u_cla22_and56;
  wire [0:0] u_cla22_and57;
  wire [0:0] u_cla22_and58;
  wire [0:0] u_cla22_and59;
  wire [0:0] u_cla22_and60;
  wire [0:0] u_cla22_and61;
  wire [0:0] u_cla22_or29;
  wire [0:0] u_cla22_or30;
  wire [0:0] u_cla22_or31;
  wire [0:0] u_cla22_pg_logic15_or0;
  wire [0:0] u_cla22_pg_logic15_and0;
  wire [0:0] u_cla22_pg_logic15_xor0;
  wire [0:0] u_cla22_xor15;
  wire [0:0] u_cla22_and62;
  wire [0:0] u_cla22_and63;
  wire [0:0] u_cla22_and64;
  wire [0:0] u_cla22_and65;
  wire [0:0] u_cla22_and66;
  wire [0:0] u_cla22_and67;
  wire [0:0] u_cla22_and68;
  wire [0:0] u_cla22_and69;
  wire [0:0] u_cla22_and70;
  wire [0:0] u_cla22_and71;
  wire [0:0] u_cla22_or32;
  wire [0:0] u_cla22_or33;
  wire [0:0] u_cla22_or34;
  wire [0:0] u_cla22_or35;
  wire [0:0] u_cla22_pg_logic16_or0;
  wire [0:0] u_cla22_pg_logic16_and0;
  wire [0:0] u_cla22_pg_logic16_xor0;
  wire [0:0] u_cla22_xor16;
  wire [0:0] u_cla22_and72;
  wire [0:0] u_cla22_or36;
  wire [0:0] u_cla22_pg_logic17_or0;
  wire [0:0] u_cla22_pg_logic17_and0;
  wire [0:0] u_cla22_pg_logic17_xor0;
  wire [0:0] u_cla22_xor17;
  wire [0:0] u_cla22_and73;
  wire [0:0] u_cla22_and74;
  wire [0:0] u_cla22_and75;
  wire [0:0] u_cla22_or37;
  wire [0:0] u_cla22_or38;
  wire [0:0] u_cla22_pg_logic18_or0;
  wire [0:0] u_cla22_pg_logic18_and0;
  wire [0:0] u_cla22_pg_logic18_xor0;
  wire [0:0] u_cla22_xor18;
  wire [0:0] u_cla22_and76;
  wire [0:0] u_cla22_and77;
  wire [0:0] u_cla22_and78;
  wire [0:0] u_cla22_and79;
  wire [0:0] u_cla22_and80;
  wire [0:0] u_cla22_and81;
  wire [0:0] u_cla22_or39;
  wire [0:0] u_cla22_or40;
  wire [0:0] u_cla22_or41;
  wire [0:0] u_cla22_pg_logic19_or0;
  wire [0:0] u_cla22_pg_logic19_and0;
  wire [0:0] u_cla22_pg_logic19_xor0;
  wire [0:0] u_cla22_xor19;
  wire [0:0] u_cla22_and82;
  wire [0:0] u_cla22_and83;
  wire [0:0] u_cla22_and84;
  wire [0:0] u_cla22_and85;
  wire [0:0] u_cla22_and86;
  wire [0:0] u_cla22_and87;
  wire [0:0] u_cla22_and88;
  wire [0:0] u_cla22_and89;
  wire [0:0] u_cla22_and90;
  wire [0:0] u_cla22_and91;
  wire [0:0] u_cla22_or42;
  wire [0:0] u_cla22_or43;
  wire [0:0] u_cla22_or44;
  wire [0:0] u_cla22_or45;
  wire [0:0] u_cla22_pg_logic20_or0;
  wire [0:0] u_cla22_pg_logic20_and0;
  wire [0:0] u_cla22_pg_logic20_xor0;
  wire [0:0] u_cla22_xor20;
  wire [0:0] u_cla22_and92;
  wire [0:0] u_cla22_or46;
  wire [0:0] u_cla22_pg_logic21_or0;
  wire [0:0] u_cla22_pg_logic21_and0;
  wire [0:0] u_cla22_pg_logic21_xor0;
  wire [0:0] u_cla22_xor21;
  wire [0:0] u_cla22_and93;
  wire [0:0] u_cla22_and94;
  wire [0:0] u_cla22_and95;
  wire [0:0] u_cla22_or47;
  wire [0:0] u_cla22_or48;

  pg_logic pg_logic_u_cla22_pg_logic0_out(.a(a[0]), .b(b[0]), .pg_logic_or0(u_cla22_pg_logic0_or0), .pg_logic_and0(u_cla22_pg_logic0_and0), .pg_logic_xor0(u_cla22_pg_logic0_xor0));
  pg_logic pg_logic_u_cla22_pg_logic1_out(.a(a[1]), .b(b[1]), .pg_logic_or0(u_cla22_pg_logic1_or0), .pg_logic_and0(u_cla22_pg_logic1_and0), .pg_logic_xor0(u_cla22_pg_logic1_xor0));
  xor_gate xor_gate_u_cla22_xor1(.a(u_cla22_pg_logic1_xor0[0]), .b(u_cla22_pg_logic0_and0[0]), .out(u_cla22_xor1));
  and_gate and_gate_u_cla22_and0(.a(u_cla22_pg_logic0_and0[0]), .b(u_cla22_pg_logic1_or0[0]), .out(u_cla22_and0));
  or_gate or_gate_u_cla22_or0(.a(u_cla22_pg_logic1_and0[0]), .b(u_cla22_and0[0]), .out(u_cla22_or0));
  pg_logic pg_logic_u_cla22_pg_logic2_out(.a(a[2]), .b(b[2]), .pg_logic_or0(u_cla22_pg_logic2_or0), .pg_logic_and0(u_cla22_pg_logic2_and0), .pg_logic_xor0(u_cla22_pg_logic2_xor0));
  xor_gate xor_gate_u_cla22_xor2(.a(u_cla22_pg_logic2_xor0[0]), .b(u_cla22_or0[0]), .out(u_cla22_xor2));
  and_gate and_gate_u_cla22_and1(.a(u_cla22_pg_logic2_or0[0]), .b(u_cla22_pg_logic0_or0[0]), .out(u_cla22_and1));
  and_gate and_gate_u_cla22_and2(.a(u_cla22_pg_logic0_and0[0]), .b(u_cla22_pg_logic2_or0[0]), .out(u_cla22_and2));
  and_gate and_gate_u_cla22_and3(.a(u_cla22_and2[0]), .b(u_cla22_pg_logic1_or0[0]), .out(u_cla22_and3));
  and_gate and_gate_u_cla22_and4(.a(u_cla22_pg_logic1_and0[0]), .b(u_cla22_pg_logic2_or0[0]), .out(u_cla22_and4));
  or_gate or_gate_u_cla22_or1(.a(u_cla22_and3[0]), .b(u_cla22_and4[0]), .out(u_cla22_or1));
  or_gate or_gate_u_cla22_or2(.a(u_cla22_pg_logic2_and0[0]), .b(u_cla22_or1[0]), .out(u_cla22_or2));
  pg_logic pg_logic_u_cla22_pg_logic3_out(.a(a[3]), .b(b[3]), .pg_logic_or0(u_cla22_pg_logic3_or0), .pg_logic_and0(u_cla22_pg_logic3_and0), .pg_logic_xor0(u_cla22_pg_logic3_xor0));
  xor_gate xor_gate_u_cla22_xor3(.a(u_cla22_pg_logic3_xor0[0]), .b(u_cla22_or2[0]), .out(u_cla22_xor3));
  and_gate and_gate_u_cla22_and5(.a(u_cla22_pg_logic3_or0[0]), .b(u_cla22_pg_logic1_or0[0]), .out(u_cla22_and5));
  and_gate and_gate_u_cla22_and6(.a(u_cla22_pg_logic0_and0[0]), .b(u_cla22_pg_logic2_or0[0]), .out(u_cla22_and6));
  and_gate and_gate_u_cla22_and7(.a(u_cla22_pg_logic3_or0[0]), .b(u_cla22_pg_logic1_or0[0]), .out(u_cla22_and7));
  and_gate and_gate_u_cla22_and8(.a(u_cla22_and6[0]), .b(u_cla22_and7[0]), .out(u_cla22_and8));
  and_gate and_gate_u_cla22_and9(.a(u_cla22_pg_logic1_and0[0]), .b(u_cla22_pg_logic3_or0[0]), .out(u_cla22_and9));
  and_gate and_gate_u_cla22_and10(.a(u_cla22_and9[0]), .b(u_cla22_pg_logic2_or0[0]), .out(u_cla22_and10));
  and_gate and_gate_u_cla22_and11(.a(u_cla22_pg_logic2_and0[0]), .b(u_cla22_pg_logic3_or0[0]), .out(u_cla22_and11));
  or_gate or_gate_u_cla22_or3(.a(u_cla22_and8[0]), .b(u_cla22_and11[0]), .out(u_cla22_or3));
  or_gate or_gate_u_cla22_or4(.a(u_cla22_and10[0]), .b(u_cla22_or3[0]), .out(u_cla22_or4));
  or_gate or_gate_u_cla22_or5(.a(u_cla22_pg_logic3_and0[0]), .b(u_cla22_or4[0]), .out(u_cla22_or5));
  pg_logic pg_logic_u_cla22_pg_logic4_out(.a(a[4]), .b(b[4]), .pg_logic_or0(u_cla22_pg_logic4_or0), .pg_logic_and0(u_cla22_pg_logic4_and0), .pg_logic_xor0(u_cla22_pg_logic4_xor0));
  xor_gate xor_gate_u_cla22_xor4(.a(u_cla22_pg_logic4_xor0[0]), .b(u_cla22_or5[0]), .out(u_cla22_xor4));
  and_gate and_gate_u_cla22_and12(.a(u_cla22_or5[0]), .b(u_cla22_pg_logic4_or0[0]), .out(u_cla22_and12));
  or_gate or_gate_u_cla22_or6(.a(u_cla22_pg_logic4_and0[0]), .b(u_cla22_and12[0]), .out(u_cla22_or6));
  pg_logic pg_logic_u_cla22_pg_logic5_out(.a(a[5]), .b(b[5]), .pg_logic_or0(u_cla22_pg_logic5_or0), .pg_logic_and0(u_cla22_pg_logic5_and0), .pg_logic_xor0(u_cla22_pg_logic5_xor0));
  xor_gate xor_gate_u_cla22_xor5(.a(u_cla22_pg_logic5_xor0[0]), .b(u_cla22_or6[0]), .out(u_cla22_xor5));
  and_gate and_gate_u_cla22_and13(.a(u_cla22_or5[0]), .b(u_cla22_pg_logic5_or0[0]), .out(u_cla22_and13));
  and_gate and_gate_u_cla22_and14(.a(u_cla22_and13[0]), .b(u_cla22_pg_logic4_or0[0]), .out(u_cla22_and14));
  and_gate and_gate_u_cla22_and15(.a(u_cla22_pg_logic4_and0[0]), .b(u_cla22_pg_logic5_or0[0]), .out(u_cla22_and15));
  or_gate or_gate_u_cla22_or7(.a(u_cla22_and14[0]), .b(u_cla22_and15[0]), .out(u_cla22_or7));
  or_gate or_gate_u_cla22_or8(.a(u_cla22_pg_logic5_and0[0]), .b(u_cla22_or7[0]), .out(u_cla22_or8));
  pg_logic pg_logic_u_cla22_pg_logic6_out(.a(a[6]), .b(b[6]), .pg_logic_or0(u_cla22_pg_logic6_or0), .pg_logic_and0(u_cla22_pg_logic6_and0), .pg_logic_xor0(u_cla22_pg_logic6_xor0));
  xor_gate xor_gate_u_cla22_xor6(.a(u_cla22_pg_logic6_xor0[0]), .b(u_cla22_or8[0]), .out(u_cla22_xor6));
  and_gate and_gate_u_cla22_and16(.a(u_cla22_or5[0]), .b(u_cla22_pg_logic5_or0[0]), .out(u_cla22_and16));
  and_gate and_gate_u_cla22_and17(.a(u_cla22_pg_logic6_or0[0]), .b(u_cla22_pg_logic4_or0[0]), .out(u_cla22_and17));
  and_gate and_gate_u_cla22_and18(.a(u_cla22_and16[0]), .b(u_cla22_and17[0]), .out(u_cla22_and18));
  and_gate and_gate_u_cla22_and19(.a(u_cla22_pg_logic4_and0[0]), .b(u_cla22_pg_logic6_or0[0]), .out(u_cla22_and19));
  and_gate and_gate_u_cla22_and20(.a(u_cla22_and19[0]), .b(u_cla22_pg_logic5_or0[0]), .out(u_cla22_and20));
  and_gate and_gate_u_cla22_and21(.a(u_cla22_pg_logic5_and0[0]), .b(u_cla22_pg_logic6_or0[0]), .out(u_cla22_and21));
  or_gate or_gate_u_cla22_or9(.a(u_cla22_and18[0]), .b(u_cla22_and20[0]), .out(u_cla22_or9));
  or_gate or_gate_u_cla22_or10(.a(u_cla22_or9[0]), .b(u_cla22_and21[0]), .out(u_cla22_or10));
  or_gate or_gate_u_cla22_or11(.a(u_cla22_pg_logic6_and0[0]), .b(u_cla22_or10[0]), .out(u_cla22_or11));
  pg_logic pg_logic_u_cla22_pg_logic7_out(.a(a[7]), .b(b[7]), .pg_logic_or0(u_cla22_pg_logic7_or0), .pg_logic_and0(u_cla22_pg_logic7_and0), .pg_logic_xor0(u_cla22_pg_logic7_xor0));
  xor_gate xor_gate_u_cla22_xor7(.a(u_cla22_pg_logic7_xor0[0]), .b(u_cla22_or11[0]), .out(u_cla22_xor7));
  and_gate and_gate_u_cla22_and22(.a(u_cla22_or5[0]), .b(u_cla22_pg_logic6_or0[0]), .out(u_cla22_and22));
  and_gate and_gate_u_cla22_and23(.a(u_cla22_pg_logic7_or0[0]), .b(u_cla22_pg_logic5_or0[0]), .out(u_cla22_and23));
  and_gate and_gate_u_cla22_and24(.a(u_cla22_and22[0]), .b(u_cla22_and23[0]), .out(u_cla22_and24));
  and_gate and_gate_u_cla22_and25(.a(u_cla22_and24[0]), .b(u_cla22_pg_logic4_or0[0]), .out(u_cla22_and25));
  and_gate and_gate_u_cla22_and26(.a(u_cla22_pg_logic4_and0[0]), .b(u_cla22_pg_logic6_or0[0]), .out(u_cla22_and26));
  and_gate and_gate_u_cla22_and27(.a(u_cla22_pg_logic7_or0[0]), .b(u_cla22_pg_logic5_or0[0]), .out(u_cla22_and27));
  and_gate and_gate_u_cla22_and28(.a(u_cla22_and26[0]), .b(u_cla22_and27[0]), .out(u_cla22_and28));
  and_gate and_gate_u_cla22_and29(.a(u_cla22_pg_logic5_and0[0]), .b(u_cla22_pg_logic7_or0[0]), .out(u_cla22_and29));
  and_gate and_gate_u_cla22_and30(.a(u_cla22_and29[0]), .b(u_cla22_pg_logic6_or0[0]), .out(u_cla22_and30));
  and_gate and_gate_u_cla22_and31(.a(u_cla22_pg_logic6_and0[0]), .b(u_cla22_pg_logic7_or0[0]), .out(u_cla22_and31));
  or_gate or_gate_u_cla22_or12(.a(u_cla22_and25[0]), .b(u_cla22_and30[0]), .out(u_cla22_or12));
  or_gate or_gate_u_cla22_or13(.a(u_cla22_and28[0]), .b(u_cla22_and31[0]), .out(u_cla22_or13));
  or_gate or_gate_u_cla22_or14(.a(u_cla22_or12[0]), .b(u_cla22_or13[0]), .out(u_cla22_or14));
  or_gate or_gate_u_cla22_or15(.a(u_cla22_pg_logic7_and0[0]), .b(u_cla22_or14[0]), .out(u_cla22_or15));
  pg_logic pg_logic_u_cla22_pg_logic8_out(.a(a[8]), .b(b[8]), .pg_logic_or0(u_cla22_pg_logic8_or0), .pg_logic_and0(u_cla22_pg_logic8_and0), .pg_logic_xor0(u_cla22_pg_logic8_xor0));
  xor_gate xor_gate_u_cla22_xor8(.a(u_cla22_pg_logic8_xor0[0]), .b(u_cla22_or15[0]), .out(u_cla22_xor8));
  and_gate and_gate_u_cla22_and32(.a(u_cla22_or15[0]), .b(u_cla22_pg_logic8_or0[0]), .out(u_cla22_and32));
  or_gate or_gate_u_cla22_or16(.a(u_cla22_pg_logic8_and0[0]), .b(u_cla22_and32[0]), .out(u_cla22_or16));
  pg_logic pg_logic_u_cla22_pg_logic9_out(.a(a[9]), .b(b[9]), .pg_logic_or0(u_cla22_pg_logic9_or0), .pg_logic_and0(u_cla22_pg_logic9_and0), .pg_logic_xor0(u_cla22_pg_logic9_xor0));
  xor_gate xor_gate_u_cla22_xor9(.a(u_cla22_pg_logic9_xor0[0]), .b(u_cla22_or16[0]), .out(u_cla22_xor9));
  and_gate and_gate_u_cla22_and33(.a(u_cla22_or15[0]), .b(u_cla22_pg_logic9_or0[0]), .out(u_cla22_and33));
  and_gate and_gate_u_cla22_and34(.a(u_cla22_and33[0]), .b(u_cla22_pg_logic8_or0[0]), .out(u_cla22_and34));
  and_gate and_gate_u_cla22_and35(.a(u_cla22_pg_logic8_and0[0]), .b(u_cla22_pg_logic9_or0[0]), .out(u_cla22_and35));
  or_gate or_gate_u_cla22_or17(.a(u_cla22_and34[0]), .b(u_cla22_and35[0]), .out(u_cla22_or17));
  or_gate or_gate_u_cla22_or18(.a(u_cla22_pg_logic9_and0[0]), .b(u_cla22_or17[0]), .out(u_cla22_or18));
  pg_logic pg_logic_u_cla22_pg_logic10_out(.a(a[10]), .b(b[10]), .pg_logic_or0(u_cla22_pg_logic10_or0), .pg_logic_and0(u_cla22_pg_logic10_and0), .pg_logic_xor0(u_cla22_pg_logic10_xor0));
  xor_gate xor_gate_u_cla22_xor10(.a(u_cla22_pg_logic10_xor0[0]), .b(u_cla22_or18[0]), .out(u_cla22_xor10));
  and_gate and_gate_u_cla22_and36(.a(u_cla22_or15[0]), .b(u_cla22_pg_logic9_or0[0]), .out(u_cla22_and36));
  and_gate and_gate_u_cla22_and37(.a(u_cla22_pg_logic10_or0[0]), .b(u_cla22_pg_logic8_or0[0]), .out(u_cla22_and37));
  and_gate and_gate_u_cla22_and38(.a(u_cla22_and36[0]), .b(u_cla22_and37[0]), .out(u_cla22_and38));
  and_gate and_gate_u_cla22_and39(.a(u_cla22_pg_logic8_and0[0]), .b(u_cla22_pg_logic10_or0[0]), .out(u_cla22_and39));
  and_gate and_gate_u_cla22_and40(.a(u_cla22_and39[0]), .b(u_cla22_pg_logic9_or0[0]), .out(u_cla22_and40));
  and_gate and_gate_u_cla22_and41(.a(u_cla22_pg_logic9_and0[0]), .b(u_cla22_pg_logic10_or0[0]), .out(u_cla22_and41));
  or_gate or_gate_u_cla22_or19(.a(u_cla22_and38[0]), .b(u_cla22_and40[0]), .out(u_cla22_or19));
  or_gate or_gate_u_cla22_or20(.a(u_cla22_or19[0]), .b(u_cla22_and41[0]), .out(u_cla22_or20));
  or_gate or_gate_u_cla22_or21(.a(u_cla22_pg_logic10_and0[0]), .b(u_cla22_or20[0]), .out(u_cla22_or21));
  pg_logic pg_logic_u_cla22_pg_logic11_out(.a(a[11]), .b(b[11]), .pg_logic_or0(u_cla22_pg_logic11_or0), .pg_logic_and0(u_cla22_pg_logic11_and0), .pg_logic_xor0(u_cla22_pg_logic11_xor0));
  xor_gate xor_gate_u_cla22_xor11(.a(u_cla22_pg_logic11_xor0[0]), .b(u_cla22_or21[0]), .out(u_cla22_xor11));
  and_gate and_gate_u_cla22_and42(.a(u_cla22_or15[0]), .b(u_cla22_pg_logic10_or0[0]), .out(u_cla22_and42));
  and_gate and_gate_u_cla22_and43(.a(u_cla22_pg_logic11_or0[0]), .b(u_cla22_pg_logic9_or0[0]), .out(u_cla22_and43));
  and_gate and_gate_u_cla22_and44(.a(u_cla22_and42[0]), .b(u_cla22_and43[0]), .out(u_cla22_and44));
  and_gate and_gate_u_cla22_and45(.a(u_cla22_and44[0]), .b(u_cla22_pg_logic8_or0[0]), .out(u_cla22_and45));
  and_gate and_gate_u_cla22_and46(.a(u_cla22_pg_logic8_and0[0]), .b(u_cla22_pg_logic10_or0[0]), .out(u_cla22_and46));
  and_gate and_gate_u_cla22_and47(.a(u_cla22_pg_logic11_or0[0]), .b(u_cla22_pg_logic9_or0[0]), .out(u_cla22_and47));
  and_gate and_gate_u_cla22_and48(.a(u_cla22_and46[0]), .b(u_cla22_and47[0]), .out(u_cla22_and48));
  and_gate and_gate_u_cla22_and49(.a(u_cla22_pg_logic9_and0[0]), .b(u_cla22_pg_logic11_or0[0]), .out(u_cla22_and49));
  and_gate and_gate_u_cla22_and50(.a(u_cla22_and49[0]), .b(u_cla22_pg_logic10_or0[0]), .out(u_cla22_and50));
  and_gate and_gate_u_cla22_and51(.a(u_cla22_pg_logic10_and0[0]), .b(u_cla22_pg_logic11_or0[0]), .out(u_cla22_and51));
  or_gate or_gate_u_cla22_or22(.a(u_cla22_and45[0]), .b(u_cla22_and50[0]), .out(u_cla22_or22));
  or_gate or_gate_u_cla22_or23(.a(u_cla22_and48[0]), .b(u_cla22_and51[0]), .out(u_cla22_or23));
  or_gate or_gate_u_cla22_or24(.a(u_cla22_or22[0]), .b(u_cla22_or23[0]), .out(u_cla22_or24));
  or_gate or_gate_u_cla22_or25(.a(u_cla22_pg_logic11_and0[0]), .b(u_cla22_or24[0]), .out(u_cla22_or25));
  pg_logic pg_logic_u_cla22_pg_logic12_out(.a(a[12]), .b(b[12]), .pg_logic_or0(u_cla22_pg_logic12_or0), .pg_logic_and0(u_cla22_pg_logic12_and0), .pg_logic_xor0(u_cla22_pg_logic12_xor0));
  xor_gate xor_gate_u_cla22_xor12(.a(u_cla22_pg_logic12_xor0[0]), .b(u_cla22_or25[0]), .out(u_cla22_xor12));
  and_gate and_gate_u_cla22_and52(.a(u_cla22_or25[0]), .b(u_cla22_pg_logic12_or0[0]), .out(u_cla22_and52));
  or_gate or_gate_u_cla22_or26(.a(u_cla22_pg_logic12_and0[0]), .b(u_cla22_and52[0]), .out(u_cla22_or26));
  pg_logic pg_logic_u_cla22_pg_logic13_out(.a(a[13]), .b(b[13]), .pg_logic_or0(u_cla22_pg_logic13_or0), .pg_logic_and0(u_cla22_pg_logic13_and0), .pg_logic_xor0(u_cla22_pg_logic13_xor0));
  xor_gate xor_gate_u_cla22_xor13(.a(u_cla22_pg_logic13_xor0[0]), .b(u_cla22_or26[0]), .out(u_cla22_xor13));
  and_gate and_gate_u_cla22_and53(.a(u_cla22_or25[0]), .b(u_cla22_pg_logic13_or0[0]), .out(u_cla22_and53));
  and_gate and_gate_u_cla22_and54(.a(u_cla22_and53[0]), .b(u_cla22_pg_logic12_or0[0]), .out(u_cla22_and54));
  and_gate and_gate_u_cla22_and55(.a(u_cla22_pg_logic12_and0[0]), .b(u_cla22_pg_logic13_or0[0]), .out(u_cla22_and55));
  or_gate or_gate_u_cla22_or27(.a(u_cla22_and54[0]), .b(u_cla22_and55[0]), .out(u_cla22_or27));
  or_gate or_gate_u_cla22_or28(.a(u_cla22_pg_logic13_and0[0]), .b(u_cla22_or27[0]), .out(u_cla22_or28));
  pg_logic pg_logic_u_cla22_pg_logic14_out(.a(a[14]), .b(b[14]), .pg_logic_or0(u_cla22_pg_logic14_or0), .pg_logic_and0(u_cla22_pg_logic14_and0), .pg_logic_xor0(u_cla22_pg_logic14_xor0));
  xor_gate xor_gate_u_cla22_xor14(.a(u_cla22_pg_logic14_xor0[0]), .b(u_cla22_or28[0]), .out(u_cla22_xor14));
  and_gate and_gate_u_cla22_and56(.a(u_cla22_or25[0]), .b(u_cla22_pg_logic13_or0[0]), .out(u_cla22_and56));
  and_gate and_gate_u_cla22_and57(.a(u_cla22_pg_logic14_or0[0]), .b(u_cla22_pg_logic12_or0[0]), .out(u_cla22_and57));
  and_gate and_gate_u_cla22_and58(.a(u_cla22_and56[0]), .b(u_cla22_and57[0]), .out(u_cla22_and58));
  and_gate and_gate_u_cla22_and59(.a(u_cla22_pg_logic12_and0[0]), .b(u_cla22_pg_logic14_or0[0]), .out(u_cla22_and59));
  and_gate and_gate_u_cla22_and60(.a(u_cla22_and59[0]), .b(u_cla22_pg_logic13_or0[0]), .out(u_cla22_and60));
  and_gate and_gate_u_cla22_and61(.a(u_cla22_pg_logic13_and0[0]), .b(u_cla22_pg_logic14_or0[0]), .out(u_cla22_and61));
  or_gate or_gate_u_cla22_or29(.a(u_cla22_and58[0]), .b(u_cla22_and60[0]), .out(u_cla22_or29));
  or_gate or_gate_u_cla22_or30(.a(u_cla22_or29[0]), .b(u_cla22_and61[0]), .out(u_cla22_or30));
  or_gate or_gate_u_cla22_or31(.a(u_cla22_pg_logic14_and0[0]), .b(u_cla22_or30[0]), .out(u_cla22_or31));
  pg_logic pg_logic_u_cla22_pg_logic15_out(.a(a[15]), .b(b[15]), .pg_logic_or0(u_cla22_pg_logic15_or0), .pg_logic_and0(u_cla22_pg_logic15_and0), .pg_logic_xor0(u_cla22_pg_logic15_xor0));
  xor_gate xor_gate_u_cla22_xor15(.a(u_cla22_pg_logic15_xor0[0]), .b(u_cla22_or31[0]), .out(u_cla22_xor15));
  and_gate and_gate_u_cla22_and62(.a(u_cla22_or25[0]), .b(u_cla22_pg_logic14_or0[0]), .out(u_cla22_and62));
  and_gate and_gate_u_cla22_and63(.a(u_cla22_pg_logic15_or0[0]), .b(u_cla22_pg_logic13_or0[0]), .out(u_cla22_and63));
  and_gate and_gate_u_cla22_and64(.a(u_cla22_and62[0]), .b(u_cla22_and63[0]), .out(u_cla22_and64));
  and_gate and_gate_u_cla22_and65(.a(u_cla22_and64[0]), .b(u_cla22_pg_logic12_or0[0]), .out(u_cla22_and65));
  and_gate and_gate_u_cla22_and66(.a(u_cla22_pg_logic12_and0[0]), .b(u_cla22_pg_logic14_or0[0]), .out(u_cla22_and66));
  and_gate and_gate_u_cla22_and67(.a(u_cla22_pg_logic15_or0[0]), .b(u_cla22_pg_logic13_or0[0]), .out(u_cla22_and67));
  and_gate and_gate_u_cla22_and68(.a(u_cla22_and66[0]), .b(u_cla22_and67[0]), .out(u_cla22_and68));
  and_gate and_gate_u_cla22_and69(.a(u_cla22_pg_logic13_and0[0]), .b(u_cla22_pg_logic15_or0[0]), .out(u_cla22_and69));
  and_gate and_gate_u_cla22_and70(.a(u_cla22_and69[0]), .b(u_cla22_pg_logic14_or0[0]), .out(u_cla22_and70));
  and_gate and_gate_u_cla22_and71(.a(u_cla22_pg_logic14_and0[0]), .b(u_cla22_pg_logic15_or0[0]), .out(u_cla22_and71));
  or_gate or_gate_u_cla22_or32(.a(u_cla22_and65[0]), .b(u_cla22_and70[0]), .out(u_cla22_or32));
  or_gate or_gate_u_cla22_or33(.a(u_cla22_and68[0]), .b(u_cla22_and71[0]), .out(u_cla22_or33));
  or_gate or_gate_u_cla22_or34(.a(u_cla22_or32[0]), .b(u_cla22_or33[0]), .out(u_cla22_or34));
  or_gate or_gate_u_cla22_or35(.a(u_cla22_pg_logic15_and0[0]), .b(u_cla22_or34[0]), .out(u_cla22_or35));
  pg_logic pg_logic_u_cla22_pg_logic16_out(.a(a[16]), .b(b[16]), .pg_logic_or0(u_cla22_pg_logic16_or0), .pg_logic_and0(u_cla22_pg_logic16_and0), .pg_logic_xor0(u_cla22_pg_logic16_xor0));
  xor_gate xor_gate_u_cla22_xor16(.a(u_cla22_pg_logic16_xor0[0]), .b(u_cla22_or35[0]), .out(u_cla22_xor16));
  and_gate and_gate_u_cla22_and72(.a(u_cla22_or35[0]), .b(u_cla22_pg_logic16_or0[0]), .out(u_cla22_and72));
  or_gate or_gate_u_cla22_or36(.a(u_cla22_pg_logic16_and0[0]), .b(u_cla22_and72[0]), .out(u_cla22_or36));
  pg_logic pg_logic_u_cla22_pg_logic17_out(.a(a[17]), .b(b[17]), .pg_logic_or0(u_cla22_pg_logic17_or0), .pg_logic_and0(u_cla22_pg_logic17_and0), .pg_logic_xor0(u_cla22_pg_logic17_xor0));
  xor_gate xor_gate_u_cla22_xor17(.a(u_cla22_pg_logic17_xor0[0]), .b(u_cla22_or36[0]), .out(u_cla22_xor17));
  and_gate and_gate_u_cla22_and73(.a(u_cla22_or35[0]), .b(u_cla22_pg_logic17_or0[0]), .out(u_cla22_and73));
  and_gate and_gate_u_cla22_and74(.a(u_cla22_and73[0]), .b(u_cla22_pg_logic16_or0[0]), .out(u_cla22_and74));
  and_gate and_gate_u_cla22_and75(.a(u_cla22_pg_logic16_and0[0]), .b(u_cla22_pg_logic17_or0[0]), .out(u_cla22_and75));
  or_gate or_gate_u_cla22_or37(.a(u_cla22_and74[0]), .b(u_cla22_and75[0]), .out(u_cla22_or37));
  or_gate or_gate_u_cla22_or38(.a(u_cla22_pg_logic17_and0[0]), .b(u_cla22_or37[0]), .out(u_cla22_or38));
  pg_logic pg_logic_u_cla22_pg_logic18_out(.a(a[18]), .b(b[18]), .pg_logic_or0(u_cla22_pg_logic18_or0), .pg_logic_and0(u_cla22_pg_logic18_and0), .pg_logic_xor0(u_cla22_pg_logic18_xor0));
  xor_gate xor_gate_u_cla22_xor18(.a(u_cla22_pg_logic18_xor0[0]), .b(u_cla22_or38[0]), .out(u_cla22_xor18));
  and_gate and_gate_u_cla22_and76(.a(u_cla22_or35[0]), .b(u_cla22_pg_logic17_or0[0]), .out(u_cla22_and76));
  and_gate and_gate_u_cla22_and77(.a(u_cla22_pg_logic18_or0[0]), .b(u_cla22_pg_logic16_or0[0]), .out(u_cla22_and77));
  and_gate and_gate_u_cla22_and78(.a(u_cla22_and76[0]), .b(u_cla22_and77[0]), .out(u_cla22_and78));
  and_gate and_gate_u_cla22_and79(.a(u_cla22_pg_logic16_and0[0]), .b(u_cla22_pg_logic18_or0[0]), .out(u_cla22_and79));
  and_gate and_gate_u_cla22_and80(.a(u_cla22_and79[0]), .b(u_cla22_pg_logic17_or0[0]), .out(u_cla22_and80));
  and_gate and_gate_u_cla22_and81(.a(u_cla22_pg_logic17_and0[0]), .b(u_cla22_pg_logic18_or0[0]), .out(u_cla22_and81));
  or_gate or_gate_u_cla22_or39(.a(u_cla22_and78[0]), .b(u_cla22_and80[0]), .out(u_cla22_or39));
  or_gate or_gate_u_cla22_or40(.a(u_cla22_or39[0]), .b(u_cla22_and81[0]), .out(u_cla22_or40));
  or_gate or_gate_u_cla22_or41(.a(u_cla22_pg_logic18_and0[0]), .b(u_cla22_or40[0]), .out(u_cla22_or41));
  pg_logic pg_logic_u_cla22_pg_logic19_out(.a(a[19]), .b(b[19]), .pg_logic_or0(u_cla22_pg_logic19_or0), .pg_logic_and0(u_cla22_pg_logic19_and0), .pg_logic_xor0(u_cla22_pg_logic19_xor0));
  xor_gate xor_gate_u_cla22_xor19(.a(u_cla22_pg_logic19_xor0[0]), .b(u_cla22_or41[0]), .out(u_cla22_xor19));
  and_gate and_gate_u_cla22_and82(.a(u_cla22_or35[0]), .b(u_cla22_pg_logic18_or0[0]), .out(u_cla22_and82));
  and_gate and_gate_u_cla22_and83(.a(u_cla22_pg_logic19_or0[0]), .b(u_cla22_pg_logic17_or0[0]), .out(u_cla22_and83));
  and_gate and_gate_u_cla22_and84(.a(u_cla22_and82[0]), .b(u_cla22_and83[0]), .out(u_cla22_and84));
  and_gate and_gate_u_cla22_and85(.a(u_cla22_and84[0]), .b(u_cla22_pg_logic16_or0[0]), .out(u_cla22_and85));
  and_gate and_gate_u_cla22_and86(.a(u_cla22_pg_logic16_and0[0]), .b(u_cla22_pg_logic18_or0[0]), .out(u_cla22_and86));
  and_gate and_gate_u_cla22_and87(.a(u_cla22_pg_logic19_or0[0]), .b(u_cla22_pg_logic17_or0[0]), .out(u_cla22_and87));
  and_gate and_gate_u_cla22_and88(.a(u_cla22_and86[0]), .b(u_cla22_and87[0]), .out(u_cla22_and88));
  and_gate and_gate_u_cla22_and89(.a(u_cla22_pg_logic17_and0[0]), .b(u_cla22_pg_logic19_or0[0]), .out(u_cla22_and89));
  and_gate and_gate_u_cla22_and90(.a(u_cla22_and89[0]), .b(u_cla22_pg_logic18_or0[0]), .out(u_cla22_and90));
  and_gate and_gate_u_cla22_and91(.a(u_cla22_pg_logic18_and0[0]), .b(u_cla22_pg_logic19_or0[0]), .out(u_cla22_and91));
  or_gate or_gate_u_cla22_or42(.a(u_cla22_and85[0]), .b(u_cla22_and90[0]), .out(u_cla22_or42));
  or_gate or_gate_u_cla22_or43(.a(u_cla22_and88[0]), .b(u_cla22_and91[0]), .out(u_cla22_or43));
  or_gate or_gate_u_cla22_or44(.a(u_cla22_or42[0]), .b(u_cla22_or43[0]), .out(u_cla22_or44));
  or_gate or_gate_u_cla22_or45(.a(u_cla22_pg_logic19_and0[0]), .b(u_cla22_or44[0]), .out(u_cla22_or45));
  pg_logic pg_logic_u_cla22_pg_logic20_out(.a(a[20]), .b(b[20]), .pg_logic_or0(u_cla22_pg_logic20_or0), .pg_logic_and0(u_cla22_pg_logic20_and0), .pg_logic_xor0(u_cla22_pg_logic20_xor0));
  xor_gate xor_gate_u_cla22_xor20(.a(u_cla22_pg_logic20_xor0[0]), .b(u_cla22_or45[0]), .out(u_cla22_xor20));
  and_gate and_gate_u_cla22_and92(.a(u_cla22_or45[0]), .b(u_cla22_pg_logic20_or0[0]), .out(u_cla22_and92));
  or_gate or_gate_u_cla22_or46(.a(u_cla22_pg_logic20_and0[0]), .b(u_cla22_and92[0]), .out(u_cla22_or46));
  pg_logic pg_logic_u_cla22_pg_logic21_out(.a(a[21]), .b(b[21]), .pg_logic_or0(u_cla22_pg_logic21_or0), .pg_logic_and0(u_cla22_pg_logic21_and0), .pg_logic_xor0(u_cla22_pg_logic21_xor0));
  xor_gate xor_gate_u_cla22_xor21(.a(u_cla22_pg_logic21_xor0[0]), .b(u_cla22_or46[0]), .out(u_cla22_xor21));
  and_gate and_gate_u_cla22_and93(.a(u_cla22_or45[0]), .b(u_cla22_pg_logic21_or0[0]), .out(u_cla22_and93));
  and_gate and_gate_u_cla22_and94(.a(u_cla22_and93[0]), .b(u_cla22_pg_logic20_or0[0]), .out(u_cla22_and94));
  and_gate and_gate_u_cla22_and95(.a(u_cla22_pg_logic20_and0[0]), .b(u_cla22_pg_logic21_or0[0]), .out(u_cla22_and95));
  or_gate or_gate_u_cla22_or47(.a(u_cla22_and94[0]), .b(u_cla22_and95[0]), .out(u_cla22_or47));
  or_gate or_gate_u_cla22_or48(.a(u_cla22_pg_logic21_and0[0]), .b(u_cla22_or47[0]), .out(u_cla22_or48));

  assign u_cla22_out[0] = u_cla22_pg_logic0_xor0[0];
  assign u_cla22_out[1] = u_cla22_xor1[0];
  assign u_cla22_out[2] = u_cla22_xor2[0];
  assign u_cla22_out[3] = u_cla22_xor3[0];
  assign u_cla22_out[4] = u_cla22_xor4[0];
  assign u_cla22_out[5] = u_cla22_xor5[0];
  assign u_cla22_out[6] = u_cla22_xor6[0];
  assign u_cla22_out[7] = u_cla22_xor7[0];
  assign u_cla22_out[8] = u_cla22_xor8[0];
  assign u_cla22_out[9] = u_cla22_xor9[0];
  assign u_cla22_out[10] = u_cla22_xor10[0];
  assign u_cla22_out[11] = u_cla22_xor11[0];
  assign u_cla22_out[12] = u_cla22_xor12[0];
  assign u_cla22_out[13] = u_cla22_xor13[0];
  assign u_cla22_out[14] = u_cla22_xor14[0];
  assign u_cla22_out[15] = u_cla22_xor15[0];
  assign u_cla22_out[16] = u_cla22_xor16[0];
  assign u_cla22_out[17] = u_cla22_xor17[0];
  assign u_cla22_out[18] = u_cla22_xor18[0];
  assign u_cla22_out[19] = u_cla22_xor19[0];
  assign u_cla22_out[20] = u_cla22_xor20[0];
  assign u_cla22_out[21] = u_cla22_xor21[0];
  assign u_cla22_out[22] = u_cla22_or48[0];
endmodule

module s_dadda_cla12(input [11:0] a, input [11:0] b, output [23:0] s_dadda_cla12_out);
  wire [0:0] s_dadda_cla12_and_9_0;
  wire [0:0] s_dadda_cla12_and_8_1;
  wire [0:0] s_dadda_cla12_ha0_xor0;
  wire [0:0] s_dadda_cla12_ha0_and0;
  wire [0:0] s_dadda_cla12_and_10_0;
  wire [0:0] s_dadda_cla12_and_9_1;
  wire [0:0] s_dadda_cla12_fa0_xor1;
  wire [0:0] s_dadda_cla12_fa0_or0;
  wire [0:0] s_dadda_cla12_and_8_2;
  wire [0:0] s_dadda_cla12_and_7_3;
  wire [0:0] s_dadda_cla12_ha1_xor0;
  wire [0:0] s_dadda_cla12_ha1_and0;
  wire [0:0] s_dadda_cla12_nand_11_0;
  wire [0:0] s_dadda_cla12_fa1_xor1;
  wire [0:0] s_dadda_cla12_fa1_or0;
  wire [0:0] s_dadda_cla12_and_10_1;
  wire [0:0] s_dadda_cla12_and_9_2;
  wire [0:0] s_dadda_cla12_and_8_3;
  wire [0:0] s_dadda_cla12_fa2_xor1;
  wire [0:0] s_dadda_cla12_fa2_or0;
  wire [0:0] s_dadda_cla12_and_7_4;
  wire [0:0] s_dadda_cla12_and_6_5;
  wire [0:0] s_dadda_cla12_ha2_xor0;
  wire [0:0] s_dadda_cla12_ha2_and0;
  wire [0:0] s_dadda_cla12_fa3_xor1;
  wire [0:0] s_dadda_cla12_fa3_or0;
  wire [0:0] s_dadda_cla12_nand_11_1;
  wire [0:0] s_dadda_cla12_and_10_2;
  wire [0:0] s_dadda_cla12_fa4_xor1;
  wire [0:0] s_dadda_cla12_fa4_or0;
  wire [0:0] s_dadda_cla12_and_9_3;
  wire [0:0] s_dadda_cla12_and_8_4;
  wire [0:0] s_dadda_cla12_and_7_5;
  wire [0:0] s_dadda_cla12_fa5_xor1;
  wire [0:0] s_dadda_cla12_fa5_or0;
  wire [0:0] s_dadda_cla12_fa6_xor1;
  wire [0:0] s_dadda_cla12_fa6_or0;
  wire [0:0] s_dadda_cla12_nand_11_2;
  wire [0:0] s_dadda_cla12_and_10_3;
  wire [0:0] s_dadda_cla12_and_9_4;
  wire [0:0] s_dadda_cla12_fa7_xor1;
  wire [0:0] s_dadda_cla12_fa7_or0;
  wire [0:0] s_dadda_cla12_nand_11_3;
  wire [0:0] s_dadda_cla12_fa8_xor1;
  wire [0:0] s_dadda_cla12_fa8_or0;
  wire [0:0] s_dadda_cla12_and_4_0;
  wire [0:0] s_dadda_cla12_and_3_1;
  wire [0:0] s_dadda_cla12_ha3_xor0;
  wire [0:0] s_dadda_cla12_ha3_and0;
  wire [0:0] s_dadda_cla12_and_5_0;
  wire [0:0] s_dadda_cla12_and_4_1;
  wire [0:0] s_dadda_cla12_fa9_xor1;
  wire [0:0] s_dadda_cla12_fa9_or0;
  wire [0:0] s_dadda_cla12_and_3_2;
  wire [0:0] s_dadda_cla12_and_2_3;
  wire [0:0] s_dadda_cla12_ha4_xor0;
  wire [0:0] s_dadda_cla12_ha4_and0;
  wire [0:0] s_dadda_cla12_and_6_0;
  wire [0:0] s_dadda_cla12_fa10_xor1;
  wire [0:0] s_dadda_cla12_fa10_or0;
  wire [0:0] s_dadda_cla12_and_5_1;
  wire [0:0] s_dadda_cla12_and_4_2;
  wire [0:0] s_dadda_cla12_and_3_3;
  wire [0:0] s_dadda_cla12_fa11_xor1;
  wire [0:0] s_dadda_cla12_fa11_or0;
  wire [0:0] s_dadda_cla12_and_2_4;
  wire [0:0] s_dadda_cla12_and_1_5;
  wire [0:0] s_dadda_cla12_ha5_xor0;
  wire [0:0] s_dadda_cla12_ha5_and0;
  wire [0:0] s_dadda_cla12_fa12_xor1;
  wire [0:0] s_dadda_cla12_fa12_or0;
  wire [0:0] s_dadda_cla12_and_7_0;
  wire [0:0] s_dadda_cla12_and_6_1;
  wire [0:0] s_dadda_cla12_and_5_2;
  wire [0:0] s_dadda_cla12_fa13_xor1;
  wire [0:0] s_dadda_cla12_fa13_or0;
  wire [0:0] s_dadda_cla12_and_4_3;
  wire [0:0] s_dadda_cla12_and_3_4;
  wire [0:0] s_dadda_cla12_and_2_5;
  wire [0:0] s_dadda_cla12_fa14_xor1;
  wire [0:0] s_dadda_cla12_fa14_or0;
  wire [0:0] s_dadda_cla12_and_1_6;
  wire [0:0] s_dadda_cla12_and_0_7;
  wire [0:0] s_dadda_cla12_ha6_xor0;
  wire [0:0] s_dadda_cla12_ha6_and0;
  wire [0:0] s_dadda_cla12_fa15_xor1;
  wire [0:0] s_dadda_cla12_fa15_or0;
  wire [0:0] s_dadda_cla12_and_8_0;
  wire [0:0] s_dadda_cla12_and_7_1;
  wire [0:0] s_dadda_cla12_fa16_xor1;
  wire [0:0] s_dadda_cla12_fa16_or0;
  wire [0:0] s_dadda_cla12_and_6_2;
  wire [0:0] s_dadda_cla12_and_5_3;
  wire [0:0] s_dadda_cla12_and_4_4;
  wire [0:0] s_dadda_cla12_fa17_xor1;
  wire [0:0] s_dadda_cla12_fa17_or0;
  wire [0:0] s_dadda_cla12_and_3_5;
  wire [0:0] s_dadda_cla12_and_2_6;
  wire [0:0] s_dadda_cla12_and_1_7;
  wire [0:0] s_dadda_cla12_fa18_xor1;
  wire [0:0] s_dadda_cla12_fa18_or0;
  wire [0:0] s_dadda_cla12_and_0_8;
  wire [0:0] s_dadda_cla12_ha7_xor0;
  wire [0:0] s_dadda_cla12_ha7_and0;
  wire [0:0] s_dadda_cla12_fa19_xor1;
  wire [0:0] s_dadda_cla12_fa19_or0;
  wire [0:0] s_dadda_cla12_and_7_2;
  wire [0:0] s_dadda_cla12_fa20_xor1;
  wire [0:0] s_dadda_cla12_fa20_or0;
  wire [0:0] s_dadda_cla12_and_6_3;
  wire [0:0] s_dadda_cla12_and_5_4;
  wire [0:0] s_dadda_cla12_and_4_5;
  wire [0:0] s_dadda_cla12_fa21_xor1;
  wire [0:0] s_dadda_cla12_fa21_or0;
  wire [0:0] s_dadda_cla12_and_3_6;
  wire [0:0] s_dadda_cla12_and_2_7;
  wire [0:0] s_dadda_cla12_and_1_8;
  wire [0:0] s_dadda_cla12_fa22_xor1;
  wire [0:0] s_dadda_cla12_fa22_or0;
  wire [0:0] s_dadda_cla12_and_0_9;
  wire [0:0] s_dadda_cla12_fa23_xor1;
  wire [0:0] s_dadda_cla12_fa23_or0;
  wire [0:0] s_dadda_cla12_fa24_xor1;
  wire [0:0] s_dadda_cla12_fa24_or0;
  wire [0:0] s_dadda_cla12_and_6_4;
  wire [0:0] s_dadda_cla12_fa25_xor1;
  wire [0:0] s_dadda_cla12_fa25_or0;
  wire [0:0] s_dadda_cla12_and_5_5;
  wire [0:0] s_dadda_cla12_and_4_6;
  wire [0:0] s_dadda_cla12_and_3_7;
  wire [0:0] s_dadda_cla12_fa26_xor1;
  wire [0:0] s_dadda_cla12_fa26_or0;
  wire [0:0] s_dadda_cla12_and_2_8;
  wire [0:0] s_dadda_cla12_and_1_9;
  wire [0:0] s_dadda_cla12_and_0_10;
  wire [0:0] s_dadda_cla12_fa27_xor1;
  wire [0:0] s_dadda_cla12_fa27_or0;
  wire [0:0] s_dadda_cla12_fa28_xor1;
  wire [0:0] s_dadda_cla12_fa28_or0;
  wire [0:0] s_dadda_cla12_fa29_xor1;
  wire [0:0] s_dadda_cla12_fa29_or0;
  wire [0:0] s_dadda_cla12_and_5_6;
  wire [0:0] s_dadda_cla12_fa30_xor1;
  wire [0:0] s_dadda_cla12_fa30_or0;
  wire [0:0] s_dadda_cla12_and_4_7;
  wire [0:0] s_dadda_cla12_and_3_8;
  wire [0:0] s_dadda_cla12_and_2_9;
  wire [0:0] s_dadda_cla12_fa31_xor1;
  wire [0:0] s_dadda_cla12_fa31_or0;
  wire [0:0] s_dadda_cla12_and_1_10;
  wire [0:0] s_dadda_cla12_nand_0_11;
  wire [0:0] s_dadda_cla12_fa32_xor1;
  wire [0:0] s_dadda_cla12_fa32_or0;
  wire [0:0] s_dadda_cla12_fa33_xor1;
  wire [0:0] s_dadda_cla12_fa33_or0;
  wire [0:0] s_dadda_cla12_fa34_xor1;
  wire [0:0] s_dadda_cla12_fa34_or0;
  wire [0:0] s_dadda_cla12_and_6_6;
  wire [0:0] s_dadda_cla12_fa35_xor1;
  wire [0:0] s_dadda_cla12_fa35_or0;
  wire [0:0] s_dadda_cla12_and_5_7;
  wire [0:0] s_dadda_cla12_and_4_8;
  wire [0:0] s_dadda_cla12_and_3_9;
  wire [0:0] s_dadda_cla12_fa36_xor1;
  wire [0:0] s_dadda_cla12_fa36_or0;
  wire [0:0] s_dadda_cla12_and_2_10;
  wire [0:0] s_dadda_cla12_nand_1_11;
  wire [0:0] s_dadda_cla12_fa37_xor1;
  wire [0:0] s_dadda_cla12_fa37_or0;
  wire [0:0] s_dadda_cla12_fa38_xor1;
  wire [0:0] s_dadda_cla12_fa38_or0;
  wire [0:0] s_dadda_cla12_fa39_xor1;
  wire [0:0] s_dadda_cla12_fa39_or0;
  wire [0:0] s_dadda_cla12_and_8_5;
  wire [0:0] s_dadda_cla12_fa40_xor1;
  wire [0:0] s_dadda_cla12_fa40_or0;
  wire [0:0] s_dadda_cla12_and_7_6;
  wire [0:0] s_dadda_cla12_and_6_7;
  wire [0:0] s_dadda_cla12_and_5_8;
  wire [0:0] s_dadda_cla12_fa41_xor1;
  wire [0:0] s_dadda_cla12_fa41_or0;
  wire [0:0] s_dadda_cla12_and_4_9;
  wire [0:0] s_dadda_cla12_and_3_10;
  wire [0:0] s_dadda_cla12_nand_2_11;
  wire [0:0] s_dadda_cla12_fa42_xor1;
  wire [0:0] s_dadda_cla12_fa42_or0;
  wire [0:0] s_dadda_cla12_fa43_xor1;
  wire [0:0] s_dadda_cla12_fa43_or0;
  wire [0:0] s_dadda_cla12_fa44_xor1;
  wire [0:0] s_dadda_cla12_fa44_or0;
  wire [0:0] s_dadda_cla12_and_10_4;
  wire [0:0] s_dadda_cla12_fa45_xor1;
  wire [0:0] s_dadda_cla12_fa45_or0;
  wire [0:0] s_dadda_cla12_and_9_5;
  wire [0:0] s_dadda_cla12_and_8_6;
  wire [0:0] s_dadda_cla12_and_7_7;
  wire [0:0] s_dadda_cla12_fa46_xor1;
  wire [0:0] s_dadda_cla12_fa46_or0;
  wire [0:0] s_dadda_cla12_and_6_8;
  wire [0:0] s_dadda_cla12_and_5_9;
  wire [0:0] s_dadda_cla12_and_4_10;
  wire [0:0] s_dadda_cla12_fa47_xor1;
  wire [0:0] s_dadda_cla12_fa47_or0;
  wire [0:0] s_dadda_cla12_nand_3_11;
  wire [0:0] s_dadda_cla12_fa48_xor1;
  wire [0:0] s_dadda_cla12_fa48_or0;
  wire [0:0] s_dadda_cla12_fa49_xor1;
  wire [0:0] s_dadda_cla12_fa49_or0;
  wire [0:0] s_dadda_cla12_fa50_xor1;
  wire [0:0] s_dadda_cla12_fa50_or0;
  wire [0:0] s_dadda_cla12_nand_11_4;
  wire [0:0] s_dadda_cla12_and_10_5;
  wire [0:0] s_dadda_cla12_and_9_6;
  wire [0:0] s_dadda_cla12_fa51_xor1;
  wire [0:0] s_dadda_cla12_fa51_or0;
  wire [0:0] s_dadda_cla12_and_8_7;
  wire [0:0] s_dadda_cla12_and_7_8;
  wire [0:0] s_dadda_cla12_and_6_9;
  wire [0:0] s_dadda_cla12_fa52_xor1;
  wire [0:0] s_dadda_cla12_fa52_or0;
  wire [0:0] s_dadda_cla12_and_5_10;
  wire [0:0] s_dadda_cla12_nand_4_11;
  wire [0:0] s_dadda_cla12_fa53_xor1;
  wire [0:0] s_dadda_cla12_fa53_or0;
  wire [0:0] s_dadda_cla12_fa54_xor1;
  wire [0:0] s_dadda_cla12_fa54_or0;
  wire [0:0] s_dadda_cla12_nand_11_5;
  wire [0:0] s_dadda_cla12_fa55_xor1;
  wire [0:0] s_dadda_cla12_fa55_or0;
  wire [0:0] s_dadda_cla12_and_10_6;
  wire [0:0] s_dadda_cla12_and_9_7;
  wire [0:0] s_dadda_cla12_and_8_8;
  wire [0:0] s_dadda_cla12_fa56_xor1;
  wire [0:0] s_dadda_cla12_fa56_or0;
  wire [0:0] s_dadda_cla12_and_7_9;
  wire [0:0] s_dadda_cla12_and_6_10;
  wire [0:0] s_dadda_cla12_nand_5_11;
  wire [0:0] s_dadda_cla12_fa57_xor1;
  wire [0:0] s_dadda_cla12_fa57_or0;
  wire [0:0] s_dadda_cla12_fa58_xor1;
  wire [0:0] s_dadda_cla12_fa58_or0;
  wire [0:0] s_dadda_cla12_nand_11_6;
  wire [0:0] s_dadda_cla12_and_10_7;
  wire [0:0] s_dadda_cla12_fa59_xor1;
  wire [0:0] s_dadda_cla12_fa59_or0;
  wire [0:0] s_dadda_cla12_and_9_8;
  wire [0:0] s_dadda_cla12_and_8_9;
  wire [0:0] s_dadda_cla12_and_7_10;
  wire [0:0] s_dadda_cla12_fa60_xor1;
  wire [0:0] s_dadda_cla12_fa60_or0;
  wire [0:0] s_dadda_cla12_fa61_xor1;
  wire [0:0] s_dadda_cla12_fa61_or0;
  wire [0:0] s_dadda_cla12_nand_11_7;
  wire [0:0] s_dadda_cla12_and_10_8;
  wire [0:0] s_dadda_cla12_and_9_9;
  wire [0:0] s_dadda_cla12_fa62_xor1;
  wire [0:0] s_dadda_cla12_fa62_or0;
  wire [0:0] s_dadda_cla12_nand_11_8;
  wire [0:0] s_dadda_cla12_fa63_xor1;
  wire [0:0] s_dadda_cla12_fa63_or0;
  wire [0:0] s_dadda_cla12_and_3_0;
  wire [0:0] s_dadda_cla12_and_2_1;
  wire [0:0] s_dadda_cla12_ha8_xor0;
  wire [0:0] s_dadda_cla12_ha8_and0;
  wire [0:0] s_dadda_cla12_and_2_2;
  wire [0:0] s_dadda_cla12_and_1_3;
  wire [0:0] s_dadda_cla12_fa64_xor1;
  wire [0:0] s_dadda_cla12_fa64_or0;
  wire [0:0] s_dadda_cla12_and_1_4;
  wire [0:0] s_dadda_cla12_and_0_5;
  wire [0:0] s_dadda_cla12_fa65_xor1;
  wire [0:0] s_dadda_cla12_fa65_or0;
  wire [0:0] s_dadda_cla12_and_0_6;
  wire [0:0] s_dadda_cla12_fa66_xor1;
  wire [0:0] s_dadda_cla12_fa66_or0;
  wire [0:0] s_dadda_cla12_fa67_xor1;
  wire [0:0] s_dadda_cla12_fa67_or0;
  wire [0:0] s_dadda_cla12_fa68_xor1;
  wire [0:0] s_dadda_cla12_fa68_or0;
  wire [0:0] s_dadda_cla12_fa69_xor1;
  wire [0:0] s_dadda_cla12_fa69_or0;
  wire [0:0] s_dadda_cla12_fa70_xor1;
  wire [0:0] s_dadda_cla12_fa70_or0;
  wire [0:0] s_dadda_cla12_fa71_xor1;
  wire [0:0] s_dadda_cla12_fa71_or0;
  wire [0:0] s_dadda_cla12_fa72_xor1;
  wire [0:0] s_dadda_cla12_fa72_or0;
  wire [0:0] s_dadda_cla12_fa73_xor1;
  wire [0:0] s_dadda_cla12_fa73_or0;
  wire [0:0] s_dadda_cla12_fa74_xor1;
  wire [0:0] s_dadda_cla12_fa74_or0;
  wire [0:0] s_dadda_cla12_fa75_xor1;
  wire [0:0] s_dadda_cla12_fa75_or0;
  wire [0:0] s_dadda_cla12_fa76_xor1;
  wire [0:0] s_dadda_cla12_fa76_or0;
  wire [0:0] s_dadda_cla12_nand_6_11;
  wire [0:0] s_dadda_cla12_fa77_xor1;
  wire [0:0] s_dadda_cla12_fa77_or0;
  wire [0:0] s_dadda_cla12_and_8_10;
  wire [0:0] s_dadda_cla12_nand_7_11;
  wire [0:0] s_dadda_cla12_fa78_xor1;
  wire [0:0] s_dadda_cla12_fa78_or0;
  wire [0:0] s_dadda_cla12_and_10_9;
  wire [0:0] s_dadda_cla12_and_9_10;
  wire [0:0] s_dadda_cla12_fa79_xor1;
  wire [0:0] s_dadda_cla12_fa79_or0;
  wire [0:0] s_dadda_cla12_nand_11_9;
  wire [0:0] s_dadda_cla12_fa80_xor1;
  wire [0:0] s_dadda_cla12_fa80_or0;
  wire [0:0] s_dadda_cla12_and_2_0;
  wire [0:0] s_dadda_cla12_and_1_1;
  wire [0:0] s_dadda_cla12_ha9_xor0;
  wire [0:0] s_dadda_cla12_ha9_and0;
  wire [0:0] s_dadda_cla12_and_1_2;
  wire [0:0] s_dadda_cla12_and_0_3;
  wire [0:0] s_dadda_cla12_fa81_xor1;
  wire [0:0] s_dadda_cla12_fa81_or0;
  wire [0:0] s_dadda_cla12_and_0_4;
  wire [0:0] s_dadda_cla12_fa82_xor1;
  wire [0:0] s_dadda_cla12_fa82_or0;
  wire [0:0] s_dadda_cla12_fa83_xor1;
  wire [0:0] s_dadda_cla12_fa83_or0;
  wire [0:0] s_dadda_cla12_fa84_xor1;
  wire [0:0] s_dadda_cla12_fa84_or0;
  wire [0:0] s_dadda_cla12_fa85_xor1;
  wire [0:0] s_dadda_cla12_fa85_or0;
  wire [0:0] s_dadda_cla12_fa86_xor1;
  wire [0:0] s_dadda_cla12_fa86_or0;
  wire [0:0] s_dadda_cla12_fa87_xor1;
  wire [0:0] s_dadda_cla12_fa87_or0;
  wire [0:0] s_dadda_cla12_fa88_xor1;
  wire [0:0] s_dadda_cla12_fa88_or0;
  wire [0:0] s_dadda_cla12_fa89_xor1;
  wire [0:0] s_dadda_cla12_fa89_or0;
  wire [0:0] s_dadda_cla12_fa90_xor1;
  wire [0:0] s_dadda_cla12_fa90_or0;
  wire [0:0] s_dadda_cla12_fa91_xor1;
  wire [0:0] s_dadda_cla12_fa91_or0;
  wire [0:0] s_dadda_cla12_fa92_xor1;
  wire [0:0] s_dadda_cla12_fa92_or0;
  wire [0:0] s_dadda_cla12_fa93_xor1;
  wire [0:0] s_dadda_cla12_fa93_or0;
  wire [0:0] s_dadda_cla12_fa94_xor1;
  wire [0:0] s_dadda_cla12_fa94_or0;
  wire [0:0] s_dadda_cla12_fa95_xor1;
  wire [0:0] s_dadda_cla12_fa95_or0;
  wire [0:0] s_dadda_cla12_fa96_xor1;
  wire [0:0] s_dadda_cla12_fa96_or0;
  wire [0:0] s_dadda_cla12_nand_8_11;
  wire [0:0] s_dadda_cla12_fa97_xor1;
  wire [0:0] s_dadda_cla12_fa97_or0;
  wire [0:0] s_dadda_cla12_and_10_10;
  wire [0:0] s_dadda_cla12_nand_9_11;
  wire [0:0] s_dadda_cla12_fa98_xor1;
  wire [0:0] s_dadda_cla12_fa98_or0;
  wire [0:0] s_dadda_cla12_nand_11_10;
  wire [0:0] s_dadda_cla12_fa99_xor1;
  wire [0:0] s_dadda_cla12_fa99_or0;
  wire [0:0] s_dadda_cla12_and_0_0;
  wire [0:0] s_dadda_cla12_and_1_0;
  wire [0:0] s_dadda_cla12_and_0_2;
  wire [0:0] s_dadda_cla12_nand_10_11;
  wire [0:0] s_dadda_cla12_and_0_1;
  wire [0:0] s_dadda_cla12_and_11_11;
  wire [21:0] s_dadda_cla12_u_cla22_a;
  wire [21:0] s_dadda_cla12_u_cla22_b;
  wire [22:0] s_dadda_cla12_u_cla22_out;
  wire [0:0] s_dadda_cla12_xor0;

  and_gate and_gate_s_dadda_cla12_and_9_0(.a(a[9]), .b(b[0]), .out(s_dadda_cla12_and_9_0));
  and_gate and_gate_s_dadda_cla12_and_8_1(.a(a[8]), .b(b[1]), .out(s_dadda_cla12_and_8_1));
  ha ha_s_dadda_cla12_ha0_out(.a(s_dadda_cla12_and_9_0[0]), .b(s_dadda_cla12_and_8_1[0]), .ha_xor0(s_dadda_cla12_ha0_xor0), .ha_and0(s_dadda_cla12_ha0_and0));
  and_gate and_gate_s_dadda_cla12_and_10_0(.a(a[10]), .b(b[0]), .out(s_dadda_cla12_and_10_0));
  and_gate and_gate_s_dadda_cla12_and_9_1(.a(a[9]), .b(b[1]), .out(s_dadda_cla12_and_9_1));
  fa fa_s_dadda_cla12_fa0_out(.a(s_dadda_cla12_ha0_and0[0]), .b(s_dadda_cla12_and_10_0[0]), .cin(s_dadda_cla12_and_9_1[0]), .fa_xor1(s_dadda_cla12_fa0_xor1), .fa_or0(s_dadda_cla12_fa0_or0));
  and_gate and_gate_s_dadda_cla12_and_8_2(.a(a[8]), .b(b[2]), .out(s_dadda_cla12_and_8_2));
  and_gate and_gate_s_dadda_cla12_and_7_3(.a(a[7]), .b(b[3]), .out(s_dadda_cla12_and_7_3));
  ha ha_s_dadda_cla12_ha1_out(.a(s_dadda_cla12_and_8_2[0]), .b(s_dadda_cla12_and_7_3[0]), .ha_xor0(s_dadda_cla12_ha1_xor0), .ha_and0(s_dadda_cla12_ha1_and0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_0(.a(a[11]), .b(b[0]), .out(s_dadda_cla12_nand_11_0));
  fa fa_s_dadda_cla12_fa1_out(.a(s_dadda_cla12_ha1_and0[0]), .b(s_dadda_cla12_fa0_or0[0]), .cin(s_dadda_cla12_nand_11_0[0]), .fa_xor1(s_dadda_cla12_fa1_xor1), .fa_or0(s_dadda_cla12_fa1_or0));
  and_gate and_gate_s_dadda_cla12_and_10_1(.a(a[10]), .b(b[1]), .out(s_dadda_cla12_and_10_1));
  and_gate and_gate_s_dadda_cla12_and_9_2(.a(a[9]), .b(b[2]), .out(s_dadda_cla12_and_9_2));
  and_gate and_gate_s_dadda_cla12_and_8_3(.a(a[8]), .b(b[3]), .out(s_dadda_cla12_and_8_3));
  fa fa_s_dadda_cla12_fa2_out(.a(s_dadda_cla12_and_10_1[0]), .b(s_dadda_cla12_and_9_2[0]), .cin(s_dadda_cla12_and_8_3[0]), .fa_xor1(s_dadda_cla12_fa2_xor1), .fa_or0(s_dadda_cla12_fa2_or0));
  and_gate and_gate_s_dadda_cla12_and_7_4(.a(a[7]), .b(b[4]), .out(s_dadda_cla12_and_7_4));
  and_gate and_gate_s_dadda_cla12_and_6_5(.a(a[6]), .b(b[5]), .out(s_dadda_cla12_and_6_5));
  ha ha_s_dadda_cla12_ha2_out(.a(s_dadda_cla12_and_7_4[0]), .b(s_dadda_cla12_and_6_5[0]), .ha_xor0(s_dadda_cla12_ha2_xor0), .ha_and0(s_dadda_cla12_ha2_and0));
  fa fa_s_dadda_cla12_fa3_out(.a(s_dadda_cla12_ha2_and0[0]), .b(s_dadda_cla12_fa2_or0[0]), .cin(s_dadda_cla12_fa1_or0[0]), .fa_xor1(s_dadda_cla12_fa3_xor1), .fa_or0(s_dadda_cla12_fa3_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_1(.a(a[11]), .b(b[1]), .out(s_dadda_cla12_nand_11_1));
  and_gate and_gate_s_dadda_cla12_and_10_2(.a(a[10]), .b(b[2]), .out(s_dadda_cla12_and_10_2));
  fa fa_s_dadda_cla12_fa4_out(.a(1'b1), .b(s_dadda_cla12_nand_11_1[0]), .cin(s_dadda_cla12_and_10_2[0]), .fa_xor1(s_dadda_cla12_fa4_xor1), .fa_or0(s_dadda_cla12_fa4_or0));
  and_gate and_gate_s_dadda_cla12_and_9_3(.a(a[9]), .b(b[3]), .out(s_dadda_cla12_and_9_3));
  and_gate and_gate_s_dadda_cla12_and_8_4(.a(a[8]), .b(b[4]), .out(s_dadda_cla12_and_8_4));
  and_gate and_gate_s_dadda_cla12_and_7_5(.a(a[7]), .b(b[5]), .out(s_dadda_cla12_and_7_5));
  fa fa_s_dadda_cla12_fa5_out(.a(s_dadda_cla12_and_9_3[0]), .b(s_dadda_cla12_and_8_4[0]), .cin(s_dadda_cla12_and_7_5[0]), .fa_xor1(s_dadda_cla12_fa5_xor1), .fa_or0(s_dadda_cla12_fa5_or0));
  fa fa_s_dadda_cla12_fa6_out(.a(s_dadda_cla12_fa5_or0[0]), .b(s_dadda_cla12_fa4_or0[0]), .cin(s_dadda_cla12_fa3_or0[0]), .fa_xor1(s_dadda_cla12_fa6_xor1), .fa_or0(s_dadda_cla12_fa6_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_2(.a(a[11]), .b(b[2]), .out(s_dadda_cla12_nand_11_2));
  and_gate and_gate_s_dadda_cla12_and_10_3(.a(a[10]), .b(b[3]), .out(s_dadda_cla12_and_10_3));
  and_gate and_gate_s_dadda_cla12_and_9_4(.a(a[9]), .b(b[4]), .out(s_dadda_cla12_and_9_4));
  fa fa_s_dadda_cla12_fa7_out(.a(s_dadda_cla12_nand_11_2[0]), .b(s_dadda_cla12_and_10_3[0]), .cin(s_dadda_cla12_and_9_4[0]), .fa_xor1(s_dadda_cla12_fa7_xor1), .fa_or0(s_dadda_cla12_fa7_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_3(.a(a[11]), .b(b[3]), .out(s_dadda_cla12_nand_11_3));
  fa fa_s_dadda_cla12_fa8_out(.a(s_dadda_cla12_fa7_or0[0]), .b(s_dadda_cla12_fa6_or0[0]), .cin(s_dadda_cla12_nand_11_3[0]), .fa_xor1(s_dadda_cla12_fa8_xor1), .fa_or0(s_dadda_cla12_fa8_or0));
  and_gate and_gate_s_dadda_cla12_and_4_0(.a(a[4]), .b(b[0]), .out(s_dadda_cla12_and_4_0));
  and_gate and_gate_s_dadda_cla12_and_3_1(.a(a[3]), .b(b[1]), .out(s_dadda_cla12_and_3_1));
  ha ha_s_dadda_cla12_ha3_out(.a(s_dadda_cla12_and_4_0[0]), .b(s_dadda_cla12_and_3_1[0]), .ha_xor0(s_dadda_cla12_ha3_xor0), .ha_and0(s_dadda_cla12_ha3_and0));
  and_gate and_gate_s_dadda_cla12_and_5_0(.a(a[5]), .b(b[0]), .out(s_dadda_cla12_and_5_0));
  and_gate and_gate_s_dadda_cla12_and_4_1(.a(a[4]), .b(b[1]), .out(s_dadda_cla12_and_4_1));
  fa fa_s_dadda_cla12_fa9_out(.a(s_dadda_cla12_ha3_and0[0]), .b(s_dadda_cla12_and_5_0[0]), .cin(s_dadda_cla12_and_4_1[0]), .fa_xor1(s_dadda_cla12_fa9_xor1), .fa_or0(s_dadda_cla12_fa9_or0));
  and_gate and_gate_s_dadda_cla12_and_3_2(.a(a[3]), .b(b[2]), .out(s_dadda_cla12_and_3_2));
  and_gate and_gate_s_dadda_cla12_and_2_3(.a(a[2]), .b(b[3]), .out(s_dadda_cla12_and_2_3));
  ha ha_s_dadda_cla12_ha4_out(.a(s_dadda_cla12_and_3_2[0]), .b(s_dadda_cla12_and_2_3[0]), .ha_xor0(s_dadda_cla12_ha4_xor0), .ha_and0(s_dadda_cla12_ha4_and0));
  and_gate and_gate_s_dadda_cla12_and_6_0(.a(a[6]), .b(b[0]), .out(s_dadda_cla12_and_6_0));
  fa fa_s_dadda_cla12_fa10_out(.a(s_dadda_cla12_ha4_and0[0]), .b(s_dadda_cla12_fa9_or0[0]), .cin(s_dadda_cla12_and_6_0[0]), .fa_xor1(s_dadda_cla12_fa10_xor1), .fa_or0(s_dadda_cla12_fa10_or0));
  and_gate and_gate_s_dadda_cla12_and_5_1(.a(a[5]), .b(b[1]), .out(s_dadda_cla12_and_5_1));
  and_gate and_gate_s_dadda_cla12_and_4_2(.a(a[4]), .b(b[2]), .out(s_dadda_cla12_and_4_2));
  and_gate and_gate_s_dadda_cla12_and_3_3(.a(a[3]), .b(b[3]), .out(s_dadda_cla12_and_3_3));
  fa fa_s_dadda_cla12_fa11_out(.a(s_dadda_cla12_and_5_1[0]), .b(s_dadda_cla12_and_4_2[0]), .cin(s_dadda_cla12_and_3_3[0]), .fa_xor1(s_dadda_cla12_fa11_xor1), .fa_or0(s_dadda_cla12_fa11_or0));
  and_gate and_gate_s_dadda_cla12_and_2_4(.a(a[2]), .b(b[4]), .out(s_dadda_cla12_and_2_4));
  and_gate and_gate_s_dadda_cla12_and_1_5(.a(a[1]), .b(b[5]), .out(s_dadda_cla12_and_1_5));
  ha ha_s_dadda_cla12_ha5_out(.a(s_dadda_cla12_and_2_4[0]), .b(s_dadda_cla12_and_1_5[0]), .ha_xor0(s_dadda_cla12_ha5_xor0), .ha_and0(s_dadda_cla12_ha5_and0));
  fa fa_s_dadda_cla12_fa12_out(.a(s_dadda_cla12_ha5_and0[0]), .b(s_dadda_cla12_fa11_or0[0]), .cin(s_dadda_cla12_fa10_or0[0]), .fa_xor1(s_dadda_cla12_fa12_xor1), .fa_or0(s_dadda_cla12_fa12_or0));
  and_gate and_gate_s_dadda_cla12_and_7_0(.a(a[7]), .b(b[0]), .out(s_dadda_cla12_and_7_0));
  and_gate and_gate_s_dadda_cla12_and_6_1(.a(a[6]), .b(b[1]), .out(s_dadda_cla12_and_6_1));
  and_gate and_gate_s_dadda_cla12_and_5_2(.a(a[5]), .b(b[2]), .out(s_dadda_cla12_and_5_2));
  fa fa_s_dadda_cla12_fa13_out(.a(s_dadda_cla12_and_7_0[0]), .b(s_dadda_cla12_and_6_1[0]), .cin(s_dadda_cla12_and_5_2[0]), .fa_xor1(s_dadda_cla12_fa13_xor1), .fa_or0(s_dadda_cla12_fa13_or0));
  and_gate and_gate_s_dadda_cla12_and_4_3(.a(a[4]), .b(b[3]), .out(s_dadda_cla12_and_4_3));
  and_gate and_gate_s_dadda_cla12_and_3_4(.a(a[3]), .b(b[4]), .out(s_dadda_cla12_and_3_4));
  and_gate and_gate_s_dadda_cla12_and_2_5(.a(a[2]), .b(b[5]), .out(s_dadda_cla12_and_2_5));
  fa fa_s_dadda_cla12_fa14_out(.a(s_dadda_cla12_and_4_3[0]), .b(s_dadda_cla12_and_3_4[0]), .cin(s_dadda_cla12_and_2_5[0]), .fa_xor1(s_dadda_cla12_fa14_xor1), .fa_or0(s_dadda_cla12_fa14_or0));
  and_gate and_gate_s_dadda_cla12_and_1_6(.a(a[1]), .b(b[6]), .out(s_dadda_cla12_and_1_6));
  and_gate and_gate_s_dadda_cla12_and_0_7(.a(a[0]), .b(b[7]), .out(s_dadda_cla12_and_0_7));
  ha ha_s_dadda_cla12_ha6_out(.a(s_dadda_cla12_and_1_6[0]), .b(s_dadda_cla12_and_0_7[0]), .ha_xor0(s_dadda_cla12_ha6_xor0), .ha_and0(s_dadda_cla12_ha6_and0));
  fa fa_s_dadda_cla12_fa15_out(.a(s_dadda_cla12_ha6_and0[0]), .b(s_dadda_cla12_fa14_or0[0]), .cin(s_dadda_cla12_fa13_or0[0]), .fa_xor1(s_dadda_cla12_fa15_xor1), .fa_or0(s_dadda_cla12_fa15_or0));
  and_gate and_gate_s_dadda_cla12_and_8_0(.a(a[8]), .b(b[0]), .out(s_dadda_cla12_and_8_0));
  and_gate and_gate_s_dadda_cla12_and_7_1(.a(a[7]), .b(b[1]), .out(s_dadda_cla12_and_7_1));
  fa fa_s_dadda_cla12_fa16_out(.a(s_dadda_cla12_fa12_or0[0]), .b(s_dadda_cla12_and_8_0[0]), .cin(s_dadda_cla12_and_7_1[0]), .fa_xor1(s_dadda_cla12_fa16_xor1), .fa_or0(s_dadda_cla12_fa16_or0));
  and_gate and_gate_s_dadda_cla12_and_6_2(.a(a[6]), .b(b[2]), .out(s_dadda_cla12_and_6_2));
  and_gate and_gate_s_dadda_cla12_and_5_3(.a(a[5]), .b(b[3]), .out(s_dadda_cla12_and_5_3));
  and_gate and_gate_s_dadda_cla12_and_4_4(.a(a[4]), .b(b[4]), .out(s_dadda_cla12_and_4_4));
  fa fa_s_dadda_cla12_fa17_out(.a(s_dadda_cla12_and_6_2[0]), .b(s_dadda_cla12_and_5_3[0]), .cin(s_dadda_cla12_and_4_4[0]), .fa_xor1(s_dadda_cla12_fa17_xor1), .fa_or0(s_dadda_cla12_fa17_or0));
  and_gate and_gate_s_dadda_cla12_and_3_5(.a(a[3]), .b(b[5]), .out(s_dadda_cla12_and_3_5));
  and_gate and_gate_s_dadda_cla12_and_2_6(.a(a[2]), .b(b[6]), .out(s_dadda_cla12_and_2_6));
  and_gate and_gate_s_dadda_cla12_and_1_7(.a(a[1]), .b(b[7]), .out(s_dadda_cla12_and_1_7));
  fa fa_s_dadda_cla12_fa18_out(.a(s_dadda_cla12_and_3_5[0]), .b(s_dadda_cla12_and_2_6[0]), .cin(s_dadda_cla12_and_1_7[0]), .fa_xor1(s_dadda_cla12_fa18_xor1), .fa_or0(s_dadda_cla12_fa18_or0));
  and_gate and_gate_s_dadda_cla12_and_0_8(.a(a[0]), .b(b[8]), .out(s_dadda_cla12_and_0_8));
  ha ha_s_dadda_cla12_ha7_out(.a(s_dadda_cla12_and_0_8[0]), .b(s_dadda_cla12_fa15_xor1[0]), .ha_xor0(s_dadda_cla12_ha7_xor0), .ha_and0(s_dadda_cla12_ha7_and0));
  fa fa_s_dadda_cla12_fa19_out(.a(s_dadda_cla12_ha7_and0[0]), .b(s_dadda_cla12_fa18_or0[0]), .cin(s_dadda_cla12_fa17_or0[0]), .fa_xor1(s_dadda_cla12_fa19_xor1), .fa_or0(s_dadda_cla12_fa19_or0));
  and_gate and_gate_s_dadda_cla12_and_7_2(.a(a[7]), .b(b[2]), .out(s_dadda_cla12_and_7_2));
  fa fa_s_dadda_cla12_fa20_out(.a(s_dadda_cla12_fa16_or0[0]), .b(s_dadda_cla12_fa15_or0[0]), .cin(s_dadda_cla12_and_7_2[0]), .fa_xor1(s_dadda_cla12_fa20_xor1), .fa_or0(s_dadda_cla12_fa20_or0));
  and_gate and_gate_s_dadda_cla12_and_6_3(.a(a[6]), .b(b[3]), .out(s_dadda_cla12_and_6_3));
  and_gate and_gate_s_dadda_cla12_and_5_4(.a(a[5]), .b(b[4]), .out(s_dadda_cla12_and_5_4));
  and_gate and_gate_s_dadda_cla12_and_4_5(.a(a[4]), .b(b[5]), .out(s_dadda_cla12_and_4_5));
  fa fa_s_dadda_cla12_fa21_out(.a(s_dadda_cla12_and_6_3[0]), .b(s_dadda_cla12_and_5_4[0]), .cin(s_dadda_cla12_and_4_5[0]), .fa_xor1(s_dadda_cla12_fa21_xor1), .fa_or0(s_dadda_cla12_fa21_or0));
  and_gate and_gate_s_dadda_cla12_and_3_6(.a(a[3]), .b(b[6]), .out(s_dadda_cla12_and_3_6));
  and_gate and_gate_s_dadda_cla12_and_2_7(.a(a[2]), .b(b[7]), .out(s_dadda_cla12_and_2_7));
  and_gate and_gate_s_dadda_cla12_and_1_8(.a(a[1]), .b(b[8]), .out(s_dadda_cla12_and_1_8));
  fa fa_s_dadda_cla12_fa22_out(.a(s_dadda_cla12_and_3_6[0]), .b(s_dadda_cla12_and_2_7[0]), .cin(s_dadda_cla12_and_1_8[0]), .fa_xor1(s_dadda_cla12_fa22_xor1), .fa_or0(s_dadda_cla12_fa22_or0));
  and_gate and_gate_s_dadda_cla12_and_0_9(.a(a[0]), .b(b[9]), .out(s_dadda_cla12_and_0_9));
  fa fa_s_dadda_cla12_fa23_out(.a(s_dadda_cla12_and_0_9[0]), .b(s_dadda_cla12_ha0_xor0[0]), .cin(s_dadda_cla12_fa19_xor1[0]), .fa_xor1(s_dadda_cla12_fa23_xor1), .fa_or0(s_dadda_cla12_fa23_or0));
  fa fa_s_dadda_cla12_fa24_out(.a(s_dadda_cla12_fa23_or0[0]), .b(s_dadda_cla12_fa22_or0[0]), .cin(s_dadda_cla12_fa21_or0[0]), .fa_xor1(s_dadda_cla12_fa24_xor1), .fa_or0(s_dadda_cla12_fa24_or0));
  and_gate and_gate_s_dadda_cla12_and_6_4(.a(a[6]), .b(b[4]), .out(s_dadda_cla12_and_6_4));
  fa fa_s_dadda_cla12_fa25_out(.a(s_dadda_cla12_fa20_or0[0]), .b(s_dadda_cla12_fa19_or0[0]), .cin(s_dadda_cla12_and_6_4[0]), .fa_xor1(s_dadda_cla12_fa25_xor1), .fa_or0(s_dadda_cla12_fa25_or0));
  and_gate and_gate_s_dadda_cla12_and_5_5(.a(a[5]), .b(b[5]), .out(s_dadda_cla12_and_5_5));
  and_gate and_gate_s_dadda_cla12_and_4_6(.a(a[4]), .b(b[6]), .out(s_dadda_cla12_and_4_6));
  and_gate and_gate_s_dadda_cla12_and_3_7(.a(a[3]), .b(b[7]), .out(s_dadda_cla12_and_3_7));
  fa fa_s_dadda_cla12_fa26_out(.a(s_dadda_cla12_and_5_5[0]), .b(s_dadda_cla12_and_4_6[0]), .cin(s_dadda_cla12_and_3_7[0]), .fa_xor1(s_dadda_cla12_fa26_xor1), .fa_or0(s_dadda_cla12_fa26_or0));
  and_gate and_gate_s_dadda_cla12_and_2_8(.a(a[2]), .b(b[8]), .out(s_dadda_cla12_and_2_8));
  and_gate and_gate_s_dadda_cla12_and_1_9(.a(a[1]), .b(b[9]), .out(s_dadda_cla12_and_1_9));
  and_gate and_gate_s_dadda_cla12_and_0_10(.a(a[0]), .b(b[10]), .out(s_dadda_cla12_and_0_10));
  fa fa_s_dadda_cla12_fa27_out(.a(s_dadda_cla12_and_2_8[0]), .b(s_dadda_cla12_and_1_9[0]), .cin(s_dadda_cla12_and_0_10[0]), .fa_xor1(s_dadda_cla12_fa27_xor1), .fa_or0(s_dadda_cla12_fa27_or0));
  fa fa_s_dadda_cla12_fa28_out(.a(s_dadda_cla12_fa0_xor1[0]), .b(s_dadda_cla12_ha1_xor0[0]), .cin(s_dadda_cla12_fa24_xor1[0]), .fa_xor1(s_dadda_cla12_fa28_xor1), .fa_or0(s_dadda_cla12_fa28_or0));
  fa fa_s_dadda_cla12_fa29_out(.a(s_dadda_cla12_fa28_or0[0]), .b(s_dadda_cla12_fa27_or0[0]), .cin(s_dadda_cla12_fa26_or0[0]), .fa_xor1(s_dadda_cla12_fa29_xor1), .fa_or0(s_dadda_cla12_fa29_or0));
  and_gate and_gate_s_dadda_cla12_and_5_6(.a(a[5]), .b(b[6]), .out(s_dadda_cla12_and_5_6));
  fa fa_s_dadda_cla12_fa30_out(.a(s_dadda_cla12_fa25_or0[0]), .b(s_dadda_cla12_fa24_or0[0]), .cin(s_dadda_cla12_and_5_6[0]), .fa_xor1(s_dadda_cla12_fa30_xor1), .fa_or0(s_dadda_cla12_fa30_or0));
  and_gate and_gate_s_dadda_cla12_and_4_7(.a(a[4]), .b(b[7]), .out(s_dadda_cla12_and_4_7));
  and_gate and_gate_s_dadda_cla12_and_3_8(.a(a[3]), .b(b[8]), .out(s_dadda_cla12_and_3_8));
  and_gate and_gate_s_dadda_cla12_and_2_9(.a(a[2]), .b(b[9]), .out(s_dadda_cla12_and_2_9));
  fa fa_s_dadda_cla12_fa31_out(.a(s_dadda_cla12_and_4_7[0]), .b(s_dadda_cla12_and_3_8[0]), .cin(s_dadda_cla12_and_2_9[0]), .fa_xor1(s_dadda_cla12_fa31_xor1), .fa_or0(s_dadda_cla12_fa31_or0));
  and_gate and_gate_s_dadda_cla12_and_1_10(.a(a[1]), .b(b[10]), .out(s_dadda_cla12_and_1_10));
  nand_gate nand_gate_s_dadda_cla12_nand_0_11(.a(a[0]), .b(b[11]), .out(s_dadda_cla12_nand_0_11));
  fa fa_s_dadda_cla12_fa32_out(.a(s_dadda_cla12_and_1_10[0]), .b(s_dadda_cla12_nand_0_11[0]), .cin(s_dadda_cla12_fa1_xor1[0]), .fa_xor1(s_dadda_cla12_fa32_xor1), .fa_or0(s_dadda_cla12_fa32_or0));
  fa fa_s_dadda_cla12_fa33_out(.a(s_dadda_cla12_fa2_xor1[0]), .b(s_dadda_cla12_ha2_xor0[0]), .cin(s_dadda_cla12_fa29_xor1[0]), .fa_xor1(s_dadda_cla12_fa33_xor1), .fa_or0(s_dadda_cla12_fa33_or0));
  fa fa_s_dadda_cla12_fa34_out(.a(s_dadda_cla12_fa33_or0[0]), .b(s_dadda_cla12_fa32_or0[0]), .cin(s_dadda_cla12_fa31_or0[0]), .fa_xor1(s_dadda_cla12_fa34_xor1), .fa_or0(s_dadda_cla12_fa34_or0));
  and_gate and_gate_s_dadda_cla12_and_6_6(.a(a[6]), .b(b[6]), .out(s_dadda_cla12_and_6_6));
  fa fa_s_dadda_cla12_fa35_out(.a(s_dadda_cla12_fa30_or0[0]), .b(s_dadda_cla12_fa29_or0[0]), .cin(s_dadda_cla12_and_6_6[0]), .fa_xor1(s_dadda_cla12_fa35_xor1), .fa_or0(s_dadda_cla12_fa35_or0));
  and_gate and_gate_s_dadda_cla12_and_5_7(.a(a[5]), .b(b[7]), .out(s_dadda_cla12_and_5_7));
  and_gate and_gate_s_dadda_cla12_and_4_8(.a(a[4]), .b(b[8]), .out(s_dadda_cla12_and_4_8));
  and_gate and_gate_s_dadda_cla12_and_3_9(.a(a[3]), .b(b[9]), .out(s_dadda_cla12_and_3_9));
  fa fa_s_dadda_cla12_fa36_out(.a(s_dadda_cla12_and_5_7[0]), .b(s_dadda_cla12_and_4_8[0]), .cin(s_dadda_cla12_and_3_9[0]), .fa_xor1(s_dadda_cla12_fa36_xor1), .fa_or0(s_dadda_cla12_fa36_or0));
  and_gate and_gate_s_dadda_cla12_and_2_10(.a(a[2]), .b(b[10]), .out(s_dadda_cla12_and_2_10));
  nand_gate nand_gate_s_dadda_cla12_nand_1_11(.a(a[1]), .b(b[11]), .out(s_dadda_cla12_nand_1_11));
  fa fa_s_dadda_cla12_fa37_out(.a(s_dadda_cla12_and_2_10[0]), .b(s_dadda_cla12_nand_1_11[0]), .cin(s_dadda_cla12_fa3_xor1[0]), .fa_xor1(s_dadda_cla12_fa37_xor1), .fa_or0(s_dadda_cla12_fa37_or0));
  fa fa_s_dadda_cla12_fa38_out(.a(s_dadda_cla12_fa4_xor1[0]), .b(s_dadda_cla12_fa5_xor1[0]), .cin(s_dadda_cla12_fa34_xor1[0]), .fa_xor1(s_dadda_cla12_fa38_xor1), .fa_or0(s_dadda_cla12_fa38_or0));
  fa fa_s_dadda_cla12_fa39_out(.a(s_dadda_cla12_fa38_or0[0]), .b(s_dadda_cla12_fa37_or0[0]), .cin(s_dadda_cla12_fa36_or0[0]), .fa_xor1(s_dadda_cla12_fa39_xor1), .fa_or0(s_dadda_cla12_fa39_or0));
  and_gate and_gate_s_dadda_cla12_and_8_5(.a(a[8]), .b(b[5]), .out(s_dadda_cla12_and_8_5));
  fa fa_s_dadda_cla12_fa40_out(.a(s_dadda_cla12_fa35_or0[0]), .b(s_dadda_cla12_fa34_or0[0]), .cin(s_dadda_cla12_and_8_5[0]), .fa_xor1(s_dadda_cla12_fa40_xor1), .fa_or0(s_dadda_cla12_fa40_or0));
  and_gate and_gate_s_dadda_cla12_and_7_6(.a(a[7]), .b(b[6]), .out(s_dadda_cla12_and_7_6));
  and_gate and_gate_s_dadda_cla12_and_6_7(.a(a[6]), .b(b[7]), .out(s_dadda_cla12_and_6_7));
  and_gate and_gate_s_dadda_cla12_and_5_8(.a(a[5]), .b(b[8]), .out(s_dadda_cla12_and_5_8));
  fa fa_s_dadda_cla12_fa41_out(.a(s_dadda_cla12_and_7_6[0]), .b(s_dadda_cla12_and_6_7[0]), .cin(s_dadda_cla12_and_5_8[0]), .fa_xor1(s_dadda_cla12_fa41_xor1), .fa_or0(s_dadda_cla12_fa41_or0));
  and_gate and_gate_s_dadda_cla12_and_4_9(.a(a[4]), .b(b[9]), .out(s_dadda_cla12_and_4_9));
  and_gate and_gate_s_dadda_cla12_and_3_10(.a(a[3]), .b(b[10]), .out(s_dadda_cla12_and_3_10));
  nand_gate nand_gate_s_dadda_cla12_nand_2_11(.a(a[2]), .b(b[11]), .out(s_dadda_cla12_nand_2_11));
  fa fa_s_dadda_cla12_fa42_out(.a(s_dadda_cla12_and_4_9[0]), .b(s_dadda_cla12_and_3_10[0]), .cin(s_dadda_cla12_nand_2_11[0]), .fa_xor1(s_dadda_cla12_fa42_xor1), .fa_or0(s_dadda_cla12_fa42_or0));
  fa fa_s_dadda_cla12_fa43_out(.a(s_dadda_cla12_fa6_xor1[0]), .b(s_dadda_cla12_fa7_xor1[0]), .cin(s_dadda_cla12_fa39_xor1[0]), .fa_xor1(s_dadda_cla12_fa43_xor1), .fa_or0(s_dadda_cla12_fa43_or0));
  fa fa_s_dadda_cla12_fa44_out(.a(s_dadda_cla12_fa43_or0[0]), .b(s_dadda_cla12_fa42_or0[0]), .cin(s_dadda_cla12_fa41_or0[0]), .fa_xor1(s_dadda_cla12_fa44_xor1), .fa_or0(s_dadda_cla12_fa44_or0));
  and_gate and_gate_s_dadda_cla12_and_10_4(.a(a[10]), .b(b[4]), .out(s_dadda_cla12_and_10_4));
  fa fa_s_dadda_cla12_fa45_out(.a(s_dadda_cla12_fa40_or0[0]), .b(s_dadda_cla12_fa39_or0[0]), .cin(s_dadda_cla12_and_10_4[0]), .fa_xor1(s_dadda_cla12_fa45_xor1), .fa_or0(s_dadda_cla12_fa45_or0));
  and_gate and_gate_s_dadda_cla12_and_9_5(.a(a[9]), .b(b[5]), .out(s_dadda_cla12_and_9_5));
  and_gate and_gate_s_dadda_cla12_and_8_6(.a(a[8]), .b(b[6]), .out(s_dadda_cla12_and_8_6));
  and_gate and_gate_s_dadda_cla12_and_7_7(.a(a[7]), .b(b[7]), .out(s_dadda_cla12_and_7_7));
  fa fa_s_dadda_cla12_fa46_out(.a(s_dadda_cla12_and_9_5[0]), .b(s_dadda_cla12_and_8_6[0]), .cin(s_dadda_cla12_and_7_7[0]), .fa_xor1(s_dadda_cla12_fa46_xor1), .fa_or0(s_dadda_cla12_fa46_or0));
  and_gate and_gate_s_dadda_cla12_and_6_8(.a(a[6]), .b(b[8]), .out(s_dadda_cla12_and_6_8));
  and_gate and_gate_s_dadda_cla12_and_5_9(.a(a[5]), .b(b[9]), .out(s_dadda_cla12_and_5_9));
  and_gate and_gate_s_dadda_cla12_and_4_10(.a(a[4]), .b(b[10]), .out(s_dadda_cla12_and_4_10));
  fa fa_s_dadda_cla12_fa47_out(.a(s_dadda_cla12_and_6_8[0]), .b(s_dadda_cla12_and_5_9[0]), .cin(s_dadda_cla12_and_4_10[0]), .fa_xor1(s_dadda_cla12_fa47_xor1), .fa_or0(s_dadda_cla12_fa47_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_3_11(.a(a[3]), .b(b[11]), .out(s_dadda_cla12_nand_3_11));
  fa fa_s_dadda_cla12_fa48_out(.a(s_dadda_cla12_nand_3_11[0]), .b(s_dadda_cla12_fa8_xor1[0]), .cin(s_dadda_cla12_fa44_xor1[0]), .fa_xor1(s_dadda_cla12_fa48_xor1), .fa_or0(s_dadda_cla12_fa48_or0));
  fa fa_s_dadda_cla12_fa49_out(.a(s_dadda_cla12_fa48_or0[0]), .b(s_dadda_cla12_fa47_or0[0]), .cin(s_dadda_cla12_fa46_or0[0]), .fa_xor1(s_dadda_cla12_fa49_xor1), .fa_or0(s_dadda_cla12_fa49_or0));
  fa fa_s_dadda_cla12_fa50_out(.a(s_dadda_cla12_fa45_or0[0]), .b(s_dadda_cla12_fa44_or0[0]), .cin(s_dadda_cla12_fa8_or0[0]), .fa_xor1(s_dadda_cla12_fa50_xor1), .fa_or0(s_dadda_cla12_fa50_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_4(.a(a[11]), .b(b[4]), .out(s_dadda_cla12_nand_11_4));
  and_gate and_gate_s_dadda_cla12_and_10_5(.a(a[10]), .b(b[5]), .out(s_dadda_cla12_and_10_5));
  and_gate and_gate_s_dadda_cla12_and_9_6(.a(a[9]), .b(b[6]), .out(s_dadda_cla12_and_9_6));
  fa fa_s_dadda_cla12_fa51_out(.a(s_dadda_cla12_nand_11_4[0]), .b(s_dadda_cla12_and_10_5[0]), .cin(s_dadda_cla12_and_9_6[0]), .fa_xor1(s_dadda_cla12_fa51_xor1), .fa_or0(s_dadda_cla12_fa51_or0));
  and_gate and_gate_s_dadda_cla12_and_8_7(.a(a[8]), .b(b[7]), .out(s_dadda_cla12_and_8_7));
  and_gate and_gate_s_dadda_cla12_and_7_8(.a(a[7]), .b(b[8]), .out(s_dadda_cla12_and_7_8));
  and_gate and_gate_s_dadda_cla12_and_6_9(.a(a[6]), .b(b[9]), .out(s_dadda_cla12_and_6_9));
  fa fa_s_dadda_cla12_fa52_out(.a(s_dadda_cla12_and_8_7[0]), .b(s_dadda_cla12_and_7_8[0]), .cin(s_dadda_cla12_and_6_9[0]), .fa_xor1(s_dadda_cla12_fa52_xor1), .fa_or0(s_dadda_cla12_fa52_or0));
  and_gate and_gate_s_dadda_cla12_and_5_10(.a(a[5]), .b(b[10]), .out(s_dadda_cla12_and_5_10));
  nand_gate nand_gate_s_dadda_cla12_nand_4_11(.a(a[4]), .b(b[11]), .out(s_dadda_cla12_nand_4_11));
  fa fa_s_dadda_cla12_fa53_out(.a(s_dadda_cla12_and_5_10[0]), .b(s_dadda_cla12_nand_4_11[0]), .cin(s_dadda_cla12_fa49_xor1[0]), .fa_xor1(s_dadda_cla12_fa53_xor1), .fa_or0(s_dadda_cla12_fa53_or0));
  fa fa_s_dadda_cla12_fa54_out(.a(s_dadda_cla12_fa53_or0[0]), .b(s_dadda_cla12_fa52_or0[0]), .cin(s_dadda_cla12_fa51_or0[0]), .fa_xor1(s_dadda_cla12_fa54_xor1), .fa_or0(s_dadda_cla12_fa54_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_5(.a(a[11]), .b(b[5]), .out(s_dadda_cla12_nand_11_5));
  fa fa_s_dadda_cla12_fa55_out(.a(s_dadda_cla12_fa50_or0[0]), .b(s_dadda_cla12_fa49_or0[0]), .cin(s_dadda_cla12_nand_11_5[0]), .fa_xor1(s_dadda_cla12_fa55_xor1), .fa_or0(s_dadda_cla12_fa55_or0));
  and_gate and_gate_s_dadda_cla12_and_10_6(.a(a[10]), .b(b[6]), .out(s_dadda_cla12_and_10_6));
  and_gate and_gate_s_dadda_cla12_and_9_7(.a(a[9]), .b(b[7]), .out(s_dadda_cla12_and_9_7));
  and_gate and_gate_s_dadda_cla12_and_8_8(.a(a[8]), .b(b[8]), .out(s_dadda_cla12_and_8_8));
  fa fa_s_dadda_cla12_fa56_out(.a(s_dadda_cla12_and_10_6[0]), .b(s_dadda_cla12_and_9_7[0]), .cin(s_dadda_cla12_and_8_8[0]), .fa_xor1(s_dadda_cla12_fa56_xor1), .fa_or0(s_dadda_cla12_fa56_or0));
  and_gate and_gate_s_dadda_cla12_and_7_9(.a(a[7]), .b(b[9]), .out(s_dadda_cla12_and_7_9));
  and_gate and_gate_s_dadda_cla12_and_6_10(.a(a[6]), .b(b[10]), .out(s_dadda_cla12_and_6_10));
  nand_gate nand_gate_s_dadda_cla12_nand_5_11(.a(a[5]), .b(b[11]), .out(s_dadda_cla12_nand_5_11));
  fa fa_s_dadda_cla12_fa57_out(.a(s_dadda_cla12_and_7_9[0]), .b(s_dadda_cla12_and_6_10[0]), .cin(s_dadda_cla12_nand_5_11[0]), .fa_xor1(s_dadda_cla12_fa57_xor1), .fa_or0(s_dadda_cla12_fa57_or0));
  fa fa_s_dadda_cla12_fa58_out(.a(s_dadda_cla12_fa57_or0[0]), .b(s_dadda_cla12_fa56_or0[0]), .cin(s_dadda_cla12_fa55_or0[0]), .fa_xor1(s_dadda_cla12_fa58_xor1), .fa_or0(s_dadda_cla12_fa58_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_6(.a(a[11]), .b(b[6]), .out(s_dadda_cla12_nand_11_6));
  and_gate and_gate_s_dadda_cla12_and_10_7(.a(a[10]), .b(b[7]), .out(s_dadda_cla12_and_10_7));
  fa fa_s_dadda_cla12_fa59_out(.a(s_dadda_cla12_fa54_or0[0]), .b(s_dadda_cla12_nand_11_6[0]), .cin(s_dadda_cla12_and_10_7[0]), .fa_xor1(s_dadda_cla12_fa59_xor1), .fa_or0(s_dadda_cla12_fa59_or0));
  and_gate and_gate_s_dadda_cla12_and_9_8(.a(a[9]), .b(b[8]), .out(s_dadda_cla12_and_9_8));
  and_gate and_gate_s_dadda_cla12_and_8_9(.a(a[8]), .b(b[9]), .out(s_dadda_cla12_and_8_9));
  and_gate and_gate_s_dadda_cla12_and_7_10(.a(a[7]), .b(b[10]), .out(s_dadda_cla12_and_7_10));
  fa fa_s_dadda_cla12_fa60_out(.a(s_dadda_cla12_and_9_8[0]), .b(s_dadda_cla12_and_8_9[0]), .cin(s_dadda_cla12_and_7_10[0]), .fa_xor1(s_dadda_cla12_fa60_xor1), .fa_or0(s_dadda_cla12_fa60_or0));
  fa fa_s_dadda_cla12_fa61_out(.a(s_dadda_cla12_fa60_or0[0]), .b(s_dadda_cla12_fa59_or0[0]), .cin(s_dadda_cla12_fa58_or0[0]), .fa_xor1(s_dadda_cla12_fa61_xor1), .fa_or0(s_dadda_cla12_fa61_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_7(.a(a[11]), .b(b[7]), .out(s_dadda_cla12_nand_11_7));
  and_gate and_gate_s_dadda_cla12_and_10_8(.a(a[10]), .b(b[8]), .out(s_dadda_cla12_and_10_8));
  and_gate and_gate_s_dadda_cla12_and_9_9(.a(a[9]), .b(b[9]), .out(s_dadda_cla12_and_9_9));
  fa fa_s_dadda_cla12_fa62_out(.a(s_dadda_cla12_nand_11_7[0]), .b(s_dadda_cla12_and_10_8[0]), .cin(s_dadda_cla12_and_9_9[0]), .fa_xor1(s_dadda_cla12_fa62_xor1), .fa_or0(s_dadda_cla12_fa62_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_8(.a(a[11]), .b(b[8]), .out(s_dadda_cla12_nand_11_8));
  fa fa_s_dadda_cla12_fa63_out(.a(s_dadda_cla12_fa62_or0[0]), .b(s_dadda_cla12_fa61_or0[0]), .cin(s_dadda_cla12_nand_11_8[0]), .fa_xor1(s_dadda_cla12_fa63_xor1), .fa_or0(s_dadda_cla12_fa63_or0));
  and_gate and_gate_s_dadda_cla12_and_3_0(.a(a[3]), .b(b[0]), .out(s_dadda_cla12_and_3_0));
  and_gate and_gate_s_dadda_cla12_and_2_1(.a(a[2]), .b(b[1]), .out(s_dadda_cla12_and_2_1));
  ha ha_s_dadda_cla12_ha8_out(.a(s_dadda_cla12_and_3_0[0]), .b(s_dadda_cla12_and_2_1[0]), .ha_xor0(s_dadda_cla12_ha8_xor0), .ha_and0(s_dadda_cla12_ha8_and0));
  and_gate and_gate_s_dadda_cla12_and_2_2(.a(a[2]), .b(b[2]), .out(s_dadda_cla12_and_2_2));
  and_gate and_gate_s_dadda_cla12_and_1_3(.a(a[1]), .b(b[3]), .out(s_dadda_cla12_and_1_3));
  fa fa_s_dadda_cla12_fa64_out(.a(s_dadda_cla12_ha8_and0[0]), .b(s_dadda_cla12_and_2_2[0]), .cin(s_dadda_cla12_and_1_3[0]), .fa_xor1(s_dadda_cla12_fa64_xor1), .fa_or0(s_dadda_cla12_fa64_or0));
  and_gate and_gate_s_dadda_cla12_and_1_4(.a(a[1]), .b(b[4]), .out(s_dadda_cla12_and_1_4));
  and_gate and_gate_s_dadda_cla12_and_0_5(.a(a[0]), .b(b[5]), .out(s_dadda_cla12_and_0_5));
  fa fa_s_dadda_cla12_fa65_out(.a(s_dadda_cla12_fa64_or0[0]), .b(s_dadda_cla12_and_1_4[0]), .cin(s_dadda_cla12_and_0_5[0]), .fa_xor1(s_dadda_cla12_fa65_xor1), .fa_or0(s_dadda_cla12_fa65_or0));
  and_gate and_gate_s_dadda_cla12_and_0_6(.a(a[0]), .b(b[6]), .out(s_dadda_cla12_and_0_6));
  fa fa_s_dadda_cla12_fa66_out(.a(s_dadda_cla12_fa65_or0[0]), .b(s_dadda_cla12_and_0_6[0]), .cin(s_dadda_cla12_fa10_xor1[0]), .fa_xor1(s_dadda_cla12_fa66_xor1), .fa_or0(s_dadda_cla12_fa66_or0));
  fa fa_s_dadda_cla12_fa67_out(.a(s_dadda_cla12_fa66_or0[0]), .b(s_dadda_cla12_fa12_xor1[0]), .cin(s_dadda_cla12_fa13_xor1[0]), .fa_xor1(s_dadda_cla12_fa67_xor1), .fa_or0(s_dadda_cla12_fa67_or0));
  fa fa_s_dadda_cla12_fa68_out(.a(s_dadda_cla12_fa67_or0[0]), .b(s_dadda_cla12_fa16_xor1[0]), .cin(s_dadda_cla12_fa17_xor1[0]), .fa_xor1(s_dadda_cla12_fa68_xor1), .fa_or0(s_dadda_cla12_fa68_or0));
  fa fa_s_dadda_cla12_fa69_out(.a(s_dadda_cla12_fa68_or0[0]), .b(s_dadda_cla12_fa20_xor1[0]), .cin(s_dadda_cla12_fa21_xor1[0]), .fa_xor1(s_dadda_cla12_fa69_xor1), .fa_or0(s_dadda_cla12_fa69_or0));
  fa fa_s_dadda_cla12_fa70_out(.a(s_dadda_cla12_fa69_or0[0]), .b(s_dadda_cla12_fa25_xor1[0]), .cin(s_dadda_cla12_fa26_xor1[0]), .fa_xor1(s_dadda_cla12_fa70_xor1), .fa_or0(s_dadda_cla12_fa70_or0));
  fa fa_s_dadda_cla12_fa71_out(.a(s_dadda_cla12_fa70_or0[0]), .b(s_dadda_cla12_fa30_xor1[0]), .cin(s_dadda_cla12_fa31_xor1[0]), .fa_xor1(s_dadda_cla12_fa71_xor1), .fa_or0(s_dadda_cla12_fa71_or0));
  fa fa_s_dadda_cla12_fa72_out(.a(s_dadda_cla12_fa71_or0[0]), .b(s_dadda_cla12_fa35_xor1[0]), .cin(s_dadda_cla12_fa36_xor1[0]), .fa_xor1(s_dadda_cla12_fa72_xor1), .fa_or0(s_dadda_cla12_fa72_or0));
  fa fa_s_dadda_cla12_fa73_out(.a(s_dadda_cla12_fa72_or0[0]), .b(s_dadda_cla12_fa40_xor1[0]), .cin(s_dadda_cla12_fa41_xor1[0]), .fa_xor1(s_dadda_cla12_fa73_xor1), .fa_or0(s_dadda_cla12_fa73_or0));
  fa fa_s_dadda_cla12_fa74_out(.a(s_dadda_cla12_fa73_or0[0]), .b(s_dadda_cla12_fa45_xor1[0]), .cin(s_dadda_cla12_fa46_xor1[0]), .fa_xor1(s_dadda_cla12_fa74_xor1), .fa_or0(s_dadda_cla12_fa74_or0));
  fa fa_s_dadda_cla12_fa75_out(.a(s_dadda_cla12_fa74_or0[0]), .b(s_dadda_cla12_fa50_xor1[0]), .cin(s_dadda_cla12_fa51_xor1[0]), .fa_xor1(s_dadda_cla12_fa75_xor1), .fa_or0(s_dadda_cla12_fa75_or0));
  fa fa_s_dadda_cla12_fa76_out(.a(s_dadda_cla12_fa75_or0[0]), .b(s_dadda_cla12_fa54_xor1[0]), .cin(s_dadda_cla12_fa55_xor1[0]), .fa_xor1(s_dadda_cla12_fa76_xor1), .fa_or0(s_dadda_cla12_fa76_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_6_11(.a(a[6]), .b(b[11]), .out(s_dadda_cla12_nand_6_11));
  fa fa_s_dadda_cla12_fa77_out(.a(s_dadda_cla12_fa76_or0[0]), .b(s_dadda_cla12_nand_6_11[0]), .cin(s_dadda_cla12_fa58_xor1[0]), .fa_xor1(s_dadda_cla12_fa77_xor1), .fa_or0(s_dadda_cla12_fa77_or0));
  and_gate and_gate_s_dadda_cla12_and_8_10(.a(a[8]), .b(b[10]), .out(s_dadda_cla12_and_8_10));
  nand_gate nand_gate_s_dadda_cla12_nand_7_11(.a(a[7]), .b(b[11]), .out(s_dadda_cla12_nand_7_11));
  fa fa_s_dadda_cla12_fa78_out(.a(s_dadda_cla12_fa77_or0[0]), .b(s_dadda_cla12_and_8_10[0]), .cin(s_dadda_cla12_nand_7_11[0]), .fa_xor1(s_dadda_cla12_fa78_xor1), .fa_or0(s_dadda_cla12_fa78_or0));
  and_gate and_gate_s_dadda_cla12_and_10_9(.a(a[10]), .b(b[9]), .out(s_dadda_cla12_and_10_9));
  and_gate and_gate_s_dadda_cla12_and_9_10(.a(a[9]), .b(b[10]), .out(s_dadda_cla12_and_9_10));
  fa fa_s_dadda_cla12_fa79_out(.a(s_dadda_cla12_fa78_or0[0]), .b(s_dadda_cla12_and_10_9[0]), .cin(s_dadda_cla12_and_9_10[0]), .fa_xor1(s_dadda_cla12_fa79_xor1), .fa_or0(s_dadda_cla12_fa79_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_9(.a(a[11]), .b(b[9]), .out(s_dadda_cla12_nand_11_9));
  fa fa_s_dadda_cla12_fa80_out(.a(s_dadda_cla12_fa79_or0[0]), .b(s_dadda_cla12_fa63_or0[0]), .cin(s_dadda_cla12_nand_11_9[0]), .fa_xor1(s_dadda_cla12_fa80_xor1), .fa_or0(s_dadda_cla12_fa80_or0));
  and_gate and_gate_s_dadda_cla12_and_2_0(.a(a[2]), .b(b[0]), .out(s_dadda_cla12_and_2_0));
  and_gate and_gate_s_dadda_cla12_and_1_1(.a(a[1]), .b(b[1]), .out(s_dadda_cla12_and_1_1));
  ha ha_s_dadda_cla12_ha9_out(.a(s_dadda_cla12_and_2_0[0]), .b(s_dadda_cla12_and_1_1[0]), .ha_xor0(s_dadda_cla12_ha9_xor0), .ha_and0(s_dadda_cla12_ha9_and0));
  and_gate and_gate_s_dadda_cla12_and_1_2(.a(a[1]), .b(b[2]), .out(s_dadda_cla12_and_1_2));
  and_gate and_gate_s_dadda_cla12_and_0_3(.a(a[0]), .b(b[3]), .out(s_dadda_cla12_and_0_3));
  fa fa_s_dadda_cla12_fa81_out(.a(s_dadda_cla12_ha9_and0[0]), .b(s_dadda_cla12_and_1_2[0]), .cin(s_dadda_cla12_and_0_3[0]), .fa_xor1(s_dadda_cla12_fa81_xor1), .fa_or0(s_dadda_cla12_fa81_or0));
  and_gate and_gate_s_dadda_cla12_and_0_4(.a(a[0]), .b(b[4]), .out(s_dadda_cla12_and_0_4));
  fa fa_s_dadda_cla12_fa82_out(.a(s_dadda_cla12_fa81_or0[0]), .b(s_dadda_cla12_and_0_4[0]), .cin(s_dadda_cla12_ha3_xor0[0]), .fa_xor1(s_dadda_cla12_fa82_xor1), .fa_or0(s_dadda_cla12_fa82_or0));
  fa fa_s_dadda_cla12_fa83_out(.a(s_dadda_cla12_fa82_or0[0]), .b(s_dadda_cla12_fa9_xor1[0]), .cin(s_dadda_cla12_ha4_xor0[0]), .fa_xor1(s_dadda_cla12_fa83_xor1), .fa_or0(s_dadda_cla12_fa83_or0));
  fa fa_s_dadda_cla12_fa84_out(.a(s_dadda_cla12_fa83_or0[0]), .b(s_dadda_cla12_fa11_xor1[0]), .cin(s_dadda_cla12_ha5_xor0[0]), .fa_xor1(s_dadda_cla12_fa84_xor1), .fa_or0(s_dadda_cla12_fa84_or0));
  fa fa_s_dadda_cla12_fa85_out(.a(s_dadda_cla12_fa84_or0[0]), .b(s_dadda_cla12_fa14_xor1[0]), .cin(s_dadda_cla12_ha6_xor0[0]), .fa_xor1(s_dadda_cla12_fa85_xor1), .fa_or0(s_dadda_cla12_fa85_or0));
  fa fa_s_dadda_cla12_fa86_out(.a(s_dadda_cla12_fa85_or0[0]), .b(s_dadda_cla12_fa18_xor1[0]), .cin(s_dadda_cla12_ha7_xor0[0]), .fa_xor1(s_dadda_cla12_fa86_xor1), .fa_or0(s_dadda_cla12_fa86_or0));
  fa fa_s_dadda_cla12_fa87_out(.a(s_dadda_cla12_fa86_or0[0]), .b(s_dadda_cla12_fa22_xor1[0]), .cin(s_dadda_cla12_fa23_xor1[0]), .fa_xor1(s_dadda_cla12_fa87_xor1), .fa_or0(s_dadda_cla12_fa87_or0));
  fa fa_s_dadda_cla12_fa88_out(.a(s_dadda_cla12_fa87_or0[0]), .b(s_dadda_cla12_fa27_xor1[0]), .cin(s_dadda_cla12_fa28_xor1[0]), .fa_xor1(s_dadda_cla12_fa88_xor1), .fa_or0(s_dadda_cla12_fa88_or0));
  fa fa_s_dadda_cla12_fa89_out(.a(s_dadda_cla12_fa88_or0[0]), .b(s_dadda_cla12_fa32_xor1[0]), .cin(s_dadda_cla12_fa33_xor1[0]), .fa_xor1(s_dadda_cla12_fa89_xor1), .fa_or0(s_dadda_cla12_fa89_or0));
  fa fa_s_dadda_cla12_fa90_out(.a(s_dadda_cla12_fa89_or0[0]), .b(s_dadda_cla12_fa37_xor1[0]), .cin(s_dadda_cla12_fa38_xor1[0]), .fa_xor1(s_dadda_cla12_fa90_xor1), .fa_or0(s_dadda_cla12_fa90_or0));
  fa fa_s_dadda_cla12_fa91_out(.a(s_dadda_cla12_fa90_or0[0]), .b(s_dadda_cla12_fa42_xor1[0]), .cin(s_dadda_cla12_fa43_xor1[0]), .fa_xor1(s_dadda_cla12_fa91_xor1), .fa_or0(s_dadda_cla12_fa91_or0));
  fa fa_s_dadda_cla12_fa92_out(.a(s_dadda_cla12_fa91_or0[0]), .b(s_dadda_cla12_fa47_xor1[0]), .cin(s_dadda_cla12_fa48_xor1[0]), .fa_xor1(s_dadda_cla12_fa92_xor1), .fa_or0(s_dadda_cla12_fa92_or0));
  fa fa_s_dadda_cla12_fa93_out(.a(s_dadda_cla12_fa92_or0[0]), .b(s_dadda_cla12_fa52_xor1[0]), .cin(s_dadda_cla12_fa53_xor1[0]), .fa_xor1(s_dadda_cla12_fa93_xor1), .fa_or0(s_dadda_cla12_fa93_or0));
  fa fa_s_dadda_cla12_fa94_out(.a(s_dadda_cla12_fa93_or0[0]), .b(s_dadda_cla12_fa56_xor1[0]), .cin(s_dadda_cla12_fa57_xor1[0]), .fa_xor1(s_dadda_cla12_fa94_xor1), .fa_or0(s_dadda_cla12_fa94_or0));
  fa fa_s_dadda_cla12_fa95_out(.a(s_dadda_cla12_fa94_or0[0]), .b(s_dadda_cla12_fa59_xor1[0]), .cin(s_dadda_cla12_fa60_xor1[0]), .fa_xor1(s_dadda_cla12_fa95_xor1), .fa_or0(s_dadda_cla12_fa95_or0));
  fa fa_s_dadda_cla12_fa96_out(.a(s_dadda_cla12_fa95_or0[0]), .b(s_dadda_cla12_fa61_xor1[0]), .cin(s_dadda_cla12_fa62_xor1[0]), .fa_xor1(s_dadda_cla12_fa96_xor1), .fa_or0(s_dadda_cla12_fa96_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_8_11(.a(a[8]), .b(b[11]), .out(s_dadda_cla12_nand_8_11));
  fa fa_s_dadda_cla12_fa97_out(.a(s_dadda_cla12_fa96_or0[0]), .b(s_dadda_cla12_nand_8_11[0]), .cin(s_dadda_cla12_fa63_xor1[0]), .fa_xor1(s_dadda_cla12_fa97_xor1), .fa_or0(s_dadda_cla12_fa97_or0));
  and_gate and_gate_s_dadda_cla12_and_10_10(.a(a[10]), .b(b[10]), .out(s_dadda_cla12_and_10_10));
  nand_gate nand_gate_s_dadda_cla12_nand_9_11(.a(a[9]), .b(b[11]), .out(s_dadda_cla12_nand_9_11));
  fa fa_s_dadda_cla12_fa98_out(.a(s_dadda_cla12_fa97_or0[0]), .b(s_dadda_cla12_and_10_10[0]), .cin(s_dadda_cla12_nand_9_11[0]), .fa_xor1(s_dadda_cla12_fa98_xor1), .fa_or0(s_dadda_cla12_fa98_or0));
  nand_gate nand_gate_s_dadda_cla12_nand_11_10(.a(a[11]), .b(b[10]), .out(s_dadda_cla12_nand_11_10));
  fa fa_s_dadda_cla12_fa99_out(.a(s_dadda_cla12_fa98_or0[0]), .b(s_dadda_cla12_fa80_or0[0]), .cin(s_dadda_cla12_nand_11_10[0]), .fa_xor1(s_dadda_cla12_fa99_xor1), .fa_or0(s_dadda_cla12_fa99_or0));
  and_gate and_gate_s_dadda_cla12_and_0_0(.a(a[0]), .b(b[0]), .out(s_dadda_cla12_and_0_0));
  and_gate and_gate_s_dadda_cla12_and_1_0(.a(a[1]), .b(b[0]), .out(s_dadda_cla12_and_1_0));
  and_gate and_gate_s_dadda_cla12_and_0_2(.a(a[0]), .b(b[2]), .out(s_dadda_cla12_and_0_2));
  nand_gate nand_gate_s_dadda_cla12_nand_10_11(.a(a[10]), .b(b[11]), .out(s_dadda_cla12_nand_10_11));
  and_gate and_gate_s_dadda_cla12_and_0_1(.a(a[0]), .b(b[1]), .out(s_dadda_cla12_and_0_1));
  and_gate and_gate_s_dadda_cla12_and_11_11(.a(a[11]), .b(b[11]), .out(s_dadda_cla12_and_11_11));
  assign s_dadda_cla12_u_cla22_a[0] = s_dadda_cla12_and_1_0[0];
  assign s_dadda_cla12_u_cla22_a[1] = s_dadda_cla12_and_0_2[0];
  assign s_dadda_cla12_u_cla22_a[2] = s_dadda_cla12_ha8_xor0[0];
  assign s_dadda_cla12_u_cla22_a[3] = s_dadda_cla12_fa64_xor1[0];
  assign s_dadda_cla12_u_cla22_a[4] = s_dadda_cla12_fa65_xor1[0];
  assign s_dadda_cla12_u_cla22_a[5] = s_dadda_cla12_fa66_xor1[0];
  assign s_dadda_cla12_u_cla22_a[6] = s_dadda_cla12_fa67_xor1[0];
  assign s_dadda_cla12_u_cla22_a[7] = s_dadda_cla12_fa68_xor1[0];
  assign s_dadda_cla12_u_cla22_a[8] = s_dadda_cla12_fa69_xor1[0];
  assign s_dadda_cla12_u_cla22_a[9] = s_dadda_cla12_fa70_xor1[0];
  assign s_dadda_cla12_u_cla22_a[10] = s_dadda_cla12_fa71_xor1[0];
  assign s_dadda_cla12_u_cla22_a[11] = s_dadda_cla12_fa72_xor1[0];
  assign s_dadda_cla12_u_cla22_a[12] = s_dadda_cla12_fa73_xor1[0];
  assign s_dadda_cla12_u_cla22_a[13] = s_dadda_cla12_fa74_xor1[0];
  assign s_dadda_cla12_u_cla22_a[14] = s_dadda_cla12_fa75_xor1[0];
  assign s_dadda_cla12_u_cla22_a[15] = s_dadda_cla12_fa76_xor1[0];
  assign s_dadda_cla12_u_cla22_a[16] = s_dadda_cla12_fa77_xor1[0];
  assign s_dadda_cla12_u_cla22_a[17] = s_dadda_cla12_fa78_xor1[0];
  assign s_dadda_cla12_u_cla22_a[18] = s_dadda_cla12_fa79_xor1[0];
  assign s_dadda_cla12_u_cla22_a[19] = s_dadda_cla12_fa80_xor1[0];
  assign s_dadda_cla12_u_cla22_a[20] = s_dadda_cla12_nand_10_11[0];
  assign s_dadda_cla12_u_cla22_a[21] = s_dadda_cla12_fa99_or0[0];
  assign s_dadda_cla12_u_cla22_b[0] = s_dadda_cla12_and_0_1[0];
  assign s_dadda_cla12_u_cla22_b[1] = s_dadda_cla12_ha9_xor0[0];
  assign s_dadda_cla12_u_cla22_b[2] = s_dadda_cla12_fa81_xor1[0];
  assign s_dadda_cla12_u_cla22_b[3] = s_dadda_cla12_fa82_xor1[0];
  assign s_dadda_cla12_u_cla22_b[4] = s_dadda_cla12_fa83_xor1[0];
  assign s_dadda_cla12_u_cla22_b[5] = s_dadda_cla12_fa84_xor1[0];
  assign s_dadda_cla12_u_cla22_b[6] = s_dadda_cla12_fa85_xor1[0];
  assign s_dadda_cla12_u_cla22_b[7] = s_dadda_cla12_fa86_xor1[0];
  assign s_dadda_cla12_u_cla22_b[8] = s_dadda_cla12_fa87_xor1[0];
  assign s_dadda_cla12_u_cla22_b[9] = s_dadda_cla12_fa88_xor1[0];
  assign s_dadda_cla12_u_cla22_b[10] = s_dadda_cla12_fa89_xor1[0];
  assign s_dadda_cla12_u_cla22_b[11] = s_dadda_cla12_fa90_xor1[0];
  assign s_dadda_cla12_u_cla22_b[12] = s_dadda_cla12_fa91_xor1[0];
  assign s_dadda_cla12_u_cla22_b[13] = s_dadda_cla12_fa92_xor1[0];
  assign s_dadda_cla12_u_cla22_b[14] = s_dadda_cla12_fa93_xor1[0];
  assign s_dadda_cla12_u_cla22_b[15] = s_dadda_cla12_fa94_xor1[0];
  assign s_dadda_cla12_u_cla22_b[16] = s_dadda_cla12_fa95_xor1[0];
  assign s_dadda_cla12_u_cla22_b[17] = s_dadda_cla12_fa96_xor1[0];
  assign s_dadda_cla12_u_cla22_b[18] = s_dadda_cla12_fa97_xor1[0];
  assign s_dadda_cla12_u_cla22_b[19] = s_dadda_cla12_fa98_xor1[0];
  assign s_dadda_cla12_u_cla22_b[20] = s_dadda_cla12_fa99_xor1[0];
  assign s_dadda_cla12_u_cla22_b[21] = s_dadda_cla12_and_11_11[0];
  u_cla22 u_cla22_s_dadda_cla12_u_cla22_out(.a(s_dadda_cla12_u_cla22_a), .b(s_dadda_cla12_u_cla22_b), .u_cla22_out(s_dadda_cla12_u_cla22_out));
  not_gate not_gate_s_dadda_cla12_xor0(.a(s_dadda_cla12_u_cla22_out[22]), .out(s_dadda_cla12_xor0));

  assign s_dadda_cla12_out[0] = s_dadda_cla12_and_0_0[0];
  assign s_dadda_cla12_out[1] = s_dadda_cla12_u_cla22_out[0];
  assign s_dadda_cla12_out[2] = s_dadda_cla12_u_cla22_out[1];
  assign s_dadda_cla12_out[3] = s_dadda_cla12_u_cla22_out[2];
  assign s_dadda_cla12_out[4] = s_dadda_cla12_u_cla22_out[3];
  assign s_dadda_cla12_out[5] = s_dadda_cla12_u_cla22_out[4];
  assign s_dadda_cla12_out[6] = s_dadda_cla12_u_cla22_out[5];
  assign s_dadda_cla12_out[7] = s_dadda_cla12_u_cla22_out[6];
  assign s_dadda_cla12_out[8] = s_dadda_cla12_u_cla22_out[7];
  assign s_dadda_cla12_out[9] = s_dadda_cla12_u_cla22_out[8];
  assign s_dadda_cla12_out[10] = s_dadda_cla12_u_cla22_out[9];
  assign s_dadda_cla12_out[11] = s_dadda_cla12_u_cla22_out[10];
  assign s_dadda_cla12_out[12] = s_dadda_cla12_u_cla22_out[11];
  assign s_dadda_cla12_out[13] = s_dadda_cla12_u_cla22_out[12];
  assign s_dadda_cla12_out[14] = s_dadda_cla12_u_cla22_out[13];
  assign s_dadda_cla12_out[15] = s_dadda_cla12_u_cla22_out[14];
  assign s_dadda_cla12_out[16] = s_dadda_cla12_u_cla22_out[15];
  assign s_dadda_cla12_out[17] = s_dadda_cla12_u_cla22_out[16];
  assign s_dadda_cla12_out[18] = s_dadda_cla12_u_cla22_out[17];
  assign s_dadda_cla12_out[19] = s_dadda_cla12_u_cla22_out[18];
  assign s_dadda_cla12_out[20] = s_dadda_cla12_u_cla22_out[19];
  assign s_dadda_cla12_out[21] = s_dadda_cla12_u_cla22_out[20];
  assign s_dadda_cla12_out[22] = s_dadda_cla12_u_cla22_out[21];
  assign s_dadda_cla12_out[23] = s_dadda_cla12_xor0[0];
endmodule