module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(.a(a[0]), .b(b[0]), .out(pg_logic_or0));
  and_gate and_gate_pg_logic_and0(.a(a[0]), .b(b[0]), .out(pg_logic_and0));
  xor_gate xor_gate_pg_logic_xor0(.a(a[0]), .b(b[0]), .out(pg_logic_xor0));
endmodule

module u_cla32(input [31:0] a, input [31:0] b, output [32:0] u_cla32_out);
  wire [0:0] u_cla32_pg_logic0_or0;
  wire [0:0] u_cla32_pg_logic0_and0;
  wire [0:0] u_cla32_pg_logic0_xor0;
  wire [0:0] u_cla32_pg_logic1_or0;
  wire [0:0] u_cla32_pg_logic1_and0;
  wire [0:0] u_cla32_pg_logic1_xor0;
  wire [0:0] u_cla32_xor1;
  wire [0:0] u_cla32_and0;
  wire [0:0] u_cla32_or0;
  wire [0:0] u_cla32_pg_logic2_or0;
  wire [0:0] u_cla32_pg_logic2_and0;
  wire [0:0] u_cla32_pg_logic2_xor0;
  wire [0:0] u_cla32_xor2;
  wire [0:0] u_cla32_and1;
  wire [0:0] u_cla32_and2;
  wire [0:0] u_cla32_and3;
  wire [0:0] u_cla32_and4;
  wire [0:0] u_cla32_or1;
  wire [0:0] u_cla32_or2;
  wire [0:0] u_cla32_pg_logic3_or0;
  wire [0:0] u_cla32_pg_logic3_and0;
  wire [0:0] u_cla32_pg_logic3_xor0;
  wire [0:0] u_cla32_xor3;
  wire [0:0] u_cla32_and5;
  wire [0:0] u_cla32_and6;
  wire [0:0] u_cla32_and7;
  wire [0:0] u_cla32_and8;
  wire [0:0] u_cla32_and9;
  wire [0:0] u_cla32_and10;
  wire [0:0] u_cla32_and11;
  wire [0:0] u_cla32_or3;
  wire [0:0] u_cla32_or4;
  wire [0:0] u_cla32_or5;
  wire [0:0] u_cla32_pg_logic4_or0;
  wire [0:0] u_cla32_pg_logic4_and0;
  wire [0:0] u_cla32_pg_logic4_xor0;
  wire [0:0] u_cla32_xor4;
  wire [0:0] u_cla32_and12;
  wire [0:0] u_cla32_or6;
  wire [0:0] u_cla32_pg_logic5_or0;
  wire [0:0] u_cla32_pg_logic5_and0;
  wire [0:0] u_cla32_pg_logic5_xor0;
  wire [0:0] u_cla32_xor5;
  wire [0:0] u_cla32_and13;
  wire [0:0] u_cla32_and14;
  wire [0:0] u_cla32_and15;
  wire [0:0] u_cla32_or7;
  wire [0:0] u_cla32_or8;
  wire [0:0] u_cla32_pg_logic6_or0;
  wire [0:0] u_cla32_pg_logic6_and0;
  wire [0:0] u_cla32_pg_logic6_xor0;
  wire [0:0] u_cla32_xor6;
  wire [0:0] u_cla32_and16;
  wire [0:0] u_cla32_and17;
  wire [0:0] u_cla32_and18;
  wire [0:0] u_cla32_and19;
  wire [0:0] u_cla32_and20;
  wire [0:0] u_cla32_and21;
  wire [0:0] u_cla32_or9;
  wire [0:0] u_cla32_or10;
  wire [0:0] u_cla32_or11;
  wire [0:0] u_cla32_pg_logic7_or0;
  wire [0:0] u_cla32_pg_logic7_and0;
  wire [0:0] u_cla32_pg_logic7_xor0;
  wire [0:0] u_cla32_xor7;
  wire [0:0] u_cla32_and22;
  wire [0:0] u_cla32_and23;
  wire [0:0] u_cla32_and24;
  wire [0:0] u_cla32_and25;
  wire [0:0] u_cla32_and26;
  wire [0:0] u_cla32_and27;
  wire [0:0] u_cla32_and28;
  wire [0:0] u_cla32_and29;
  wire [0:0] u_cla32_and30;
  wire [0:0] u_cla32_and31;
  wire [0:0] u_cla32_or12;
  wire [0:0] u_cla32_or13;
  wire [0:0] u_cla32_or14;
  wire [0:0] u_cla32_or15;
  wire [0:0] u_cla32_pg_logic8_or0;
  wire [0:0] u_cla32_pg_logic8_and0;
  wire [0:0] u_cla32_pg_logic8_xor0;
  wire [0:0] u_cla32_xor8;
  wire [0:0] u_cla32_and32;
  wire [0:0] u_cla32_or16;
  wire [0:0] u_cla32_pg_logic9_or0;
  wire [0:0] u_cla32_pg_logic9_and0;
  wire [0:0] u_cla32_pg_logic9_xor0;
  wire [0:0] u_cla32_xor9;
  wire [0:0] u_cla32_and33;
  wire [0:0] u_cla32_and34;
  wire [0:0] u_cla32_and35;
  wire [0:0] u_cla32_or17;
  wire [0:0] u_cla32_or18;
  wire [0:0] u_cla32_pg_logic10_or0;
  wire [0:0] u_cla32_pg_logic10_and0;
  wire [0:0] u_cla32_pg_logic10_xor0;
  wire [0:0] u_cla32_xor10;
  wire [0:0] u_cla32_and36;
  wire [0:0] u_cla32_and37;
  wire [0:0] u_cla32_and38;
  wire [0:0] u_cla32_and39;
  wire [0:0] u_cla32_and40;
  wire [0:0] u_cla32_and41;
  wire [0:0] u_cla32_or19;
  wire [0:0] u_cla32_or20;
  wire [0:0] u_cla32_or21;
  wire [0:0] u_cla32_pg_logic11_or0;
  wire [0:0] u_cla32_pg_logic11_and0;
  wire [0:0] u_cla32_pg_logic11_xor0;
  wire [0:0] u_cla32_xor11;
  wire [0:0] u_cla32_and42;
  wire [0:0] u_cla32_and43;
  wire [0:0] u_cla32_and44;
  wire [0:0] u_cla32_and45;
  wire [0:0] u_cla32_and46;
  wire [0:0] u_cla32_and47;
  wire [0:0] u_cla32_and48;
  wire [0:0] u_cla32_and49;
  wire [0:0] u_cla32_and50;
  wire [0:0] u_cla32_and51;
  wire [0:0] u_cla32_or22;
  wire [0:0] u_cla32_or23;
  wire [0:0] u_cla32_or24;
  wire [0:0] u_cla32_or25;
  wire [0:0] u_cla32_pg_logic12_or0;
  wire [0:0] u_cla32_pg_logic12_and0;
  wire [0:0] u_cla32_pg_logic12_xor0;
  wire [0:0] u_cla32_xor12;
  wire [0:0] u_cla32_and52;
  wire [0:0] u_cla32_or26;
  wire [0:0] u_cla32_pg_logic13_or0;
  wire [0:0] u_cla32_pg_logic13_and0;
  wire [0:0] u_cla32_pg_logic13_xor0;
  wire [0:0] u_cla32_xor13;
  wire [0:0] u_cla32_and53;
  wire [0:0] u_cla32_and54;
  wire [0:0] u_cla32_and55;
  wire [0:0] u_cla32_or27;
  wire [0:0] u_cla32_or28;
  wire [0:0] u_cla32_pg_logic14_or0;
  wire [0:0] u_cla32_pg_logic14_and0;
  wire [0:0] u_cla32_pg_logic14_xor0;
  wire [0:0] u_cla32_xor14;
  wire [0:0] u_cla32_and56;
  wire [0:0] u_cla32_and57;
  wire [0:0] u_cla32_and58;
  wire [0:0] u_cla32_and59;
  wire [0:0] u_cla32_and60;
  wire [0:0] u_cla32_and61;
  wire [0:0] u_cla32_or29;
  wire [0:0] u_cla32_or30;
  wire [0:0] u_cla32_or31;
  wire [0:0] u_cla32_pg_logic15_or0;
  wire [0:0] u_cla32_pg_logic15_and0;
  wire [0:0] u_cla32_pg_logic15_xor0;
  wire [0:0] u_cla32_xor15;
  wire [0:0] u_cla32_and62;
  wire [0:0] u_cla32_and63;
  wire [0:0] u_cla32_and64;
  wire [0:0] u_cla32_and65;
  wire [0:0] u_cla32_and66;
  wire [0:0] u_cla32_and67;
  wire [0:0] u_cla32_and68;
  wire [0:0] u_cla32_and69;
  wire [0:0] u_cla32_and70;
  wire [0:0] u_cla32_and71;
  wire [0:0] u_cla32_or32;
  wire [0:0] u_cla32_or33;
  wire [0:0] u_cla32_or34;
  wire [0:0] u_cla32_or35;
  wire [0:0] u_cla32_pg_logic16_or0;
  wire [0:0] u_cla32_pg_logic16_and0;
  wire [0:0] u_cla32_pg_logic16_xor0;
  wire [0:0] u_cla32_xor16;
  wire [0:0] u_cla32_and72;
  wire [0:0] u_cla32_or36;
  wire [0:0] u_cla32_pg_logic17_or0;
  wire [0:0] u_cla32_pg_logic17_and0;
  wire [0:0] u_cla32_pg_logic17_xor0;
  wire [0:0] u_cla32_xor17;
  wire [0:0] u_cla32_and73;
  wire [0:0] u_cla32_and74;
  wire [0:0] u_cla32_and75;
  wire [0:0] u_cla32_or37;
  wire [0:0] u_cla32_or38;
  wire [0:0] u_cla32_pg_logic18_or0;
  wire [0:0] u_cla32_pg_logic18_and0;
  wire [0:0] u_cla32_pg_logic18_xor0;
  wire [0:0] u_cla32_xor18;
  wire [0:0] u_cla32_and76;
  wire [0:0] u_cla32_and77;
  wire [0:0] u_cla32_and78;
  wire [0:0] u_cla32_and79;
  wire [0:0] u_cla32_and80;
  wire [0:0] u_cla32_and81;
  wire [0:0] u_cla32_or39;
  wire [0:0] u_cla32_or40;
  wire [0:0] u_cla32_or41;
  wire [0:0] u_cla32_pg_logic19_or0;
  wire [0:0] u_cla32_pg_logic19_and0;
  wire [0:0] u_cla32_pg_logic19_xor0;
  wire [0:0] u_cla32_xor19;
  wire [0:0] u_cla32_and82;
  wire [0:0] u_cla32_and83;
  wire [0:0] u_cla32_and84;
  wire [0:0] u_cla32_and85;
  wire [0:0] u_cla32_and86;
  wire [0:0] u_cla32_and87;
  wire [0:0] u_cla32_and88;
  wire [0:0] u_cla32_and89;
  wire [0:0] u_cla32_and90;
  wire [0:0] u_cla32_and91;
  wire [0:0] u_cla32_or42;
  wire [0:0] u_cla32_or43;
  wire [0:0] u_cla32_or44;
  wire [0:0] u_cla32_or45;
  wire [0:0] u_cla32_pg_logic20_or0;
  wire [0:0] u_cla32_pg_logic20_and0;
  wire [0:0] u_cla32_pg_logic20_xor0;
  wire [0:0] u_cla32_xor20;
  wire [0:0] u_cla32_and92;
  wire [0:0] u_cla32_or46;
  wire [0:0] u_cla32_pg_logic21_or0;
  wire [0:0] u_cla32_pg_logic21_and0;
  wire [0:0] u_cla32_pg_logic21_xor0;
  wire [0:0] u_cla32_xor21;
  wire [0:0] u_cla32_and93;
  wire [0:0] u_cla32_and94;
  wire [0:0] u_cla32_and95;
  wire [0:0] u_cla32_or47;
  wire [0:0] u_cla32_or48;
  wire [0:0] u_cla32_pg_logic22_or0;
  wire [0:0] u_cla32_pg_logic22_and0;
  wire [0:0] u_cla32_pg_logic22_xor0;
  wire [0:0] u_cla32_xor22;
  wire [0:0] u_cla32_and96;
  wire [0:0] u_cla32_and97;
  wire [0:0] u_cla32_and98;
  wire [0:0] u_cla32_and99;
  wire [0:0] u_cla32_and100;
  wire [0:0] u_cla32_and101;
  wire [0:0] u_cla32_or49;
  wire [0:0] u_cla32_or50;
  wire [0:0] u_cla32_or51;
  wire [0:0] u_cla32_pg_logic23_or0;
  wire [0:0] u_cla32_pg_logic23_and0;
  wire [0:0] u_cla32_pg_logic23_xor0;
  wire [0:0] u_cla32_xor23;
  wire [0:0] u_cla32_and102;
  wire [0:0] u_cla32_and103;
  wire [0:0] u_cla32_and104;
  wire [0:0] u_cla32_and105;
  wire [0:0] u_cla32_and106;
  wire [0:0] u_cla32_and107;
  wire [0:0] u_cla32_and108;
  wire [0:0] u_cla32_and109;
  wire [0:0] u_cla32_and110;
  wire [0:0] u_cla32_and111;
  wire [0:0] u_cla32_or52;
  wire [0:0] u_cla32_or53;
  wire [0:0] u_cla32_or54;
  wire [0:0] u_cla32_or55;
  wire [0:0] u_cla32_pg_logic24_or0;
  wire [0:0] u_cla32_pg_logic24_and0;
  wire [0:0] u_cla32_pg_logic24_xor0;
  wire [0:0] u_cla32_xor24;
  wire [0:0] u_cla32_and112;
  wire [0:0] u_cla32_or56;
  wire [0:0] u_cla32_pg_logic25_or0;
  wire [0:0] u_cla32_pg_logic25_and0;
  wire [0:0] u_cla32_pg_logic25_xor0;
  wire [0:0] u_cla32_xor25;
  wire [0:0] u_cla32_and113;
  wire [0:0] u_cla32_and114;
  wire [0:0] u_cla32_and115;
  wire [0:0] u_cla32_or57;
  wire [0:0] u_cla32_or58;
  wire [0:0] u_cla32_pg_logic26_or0;
  wire [0:0] u_cla32_pg_logic26_and0;
  wire [0:0] u_cla32_pg_logic26_xor0;
  wire [0:0] u_cla32_xor26;
  wire [0:0] u_cla32_and116;
  wire [0:0] u_cla32_and117;
  wire [0:0] u_cla32_and118;
  wire [0:0] u_cla32_and119;
  wire [0:0] u_cla32_and120;
  wire [0:0] u_cla32_and121;
  wire [0:0] u_cla32_or59;
  wire [0:0] u_cla32_or60;
  wire [0:0] u_cla32_or61;
  wire [0:0] u_cla32_pg_logic27_or0;
  wire [0:0] u_cla32_pg_logic27_and0;
  wire [0:0] u_cla32_pg_logic27_xor0;
  wire [0:0] u_cla32_xor27;
  wire [0:0] u_cla32_and122;
  wire [0:0] u_cla32_and123;
  wire [0:0] u_cla32_and124;
  wire [0:0] u_cla32_and125;
  wire [0:0] u_cla32_and126;
  wire [0:0] u_cla32_and127;
  wire [0:0] u_cla32_and128;
  wire [0:0] u_cla32_and129;
  wire [0:0] u_cla32_and130;
  wire [0:0] u_cla32_and131;
  wire [0:0] u_cla32_or62;
  wire [0:0] u_cla32_or63;
  wire [0:0] u_cla32_or64;
  wire [0:0] u_cla32_or65;
  wire [0:0] u_cla32_pg_logic28_or0;
  wire [0:0] u_cla32_pg_logic28_and0;
  wire [0:0] u_cla32_pg_logic28_xor0;
  wire [0:0] u_cla32_xor28;
  wire [0:0] u_cla32_and132;
  wire [0:0] u_cla32_or66;
  wire [0:0] u_cla32_pg_logic29_or0;
  wire [0:0] u_cla32_pg_logic29_and0;
  wire [0:0] u_cla32_pg_logic29_xor0;
  wire [0:0] u_cla32_xor29;
  wire [0:0] u_cla32_and133;
  wire [0:0] u_cla32_and134;
  wire [0:0] u_cla32_and135;
  wire [0:0] u_cla32_or67;
  wire [0:0] u_cla32_or68;
  wire [0:0] u_cla32_pg_logic30_or0;
  wire [0:0] u_cla32_pg_logic30_and0;
  wire [0:0] u_cla32_pg_logic30_xor0;
  wire [0:0] u_cla32_xor30;
  wire [0:0] u_cla32_and136;
  wire [0:0] u_cla32_and137;
  wire [0:0] u_cla32_and138;
  wire [0:0] u_cla32_and139;
  wire [0:0] u_cla32_and140;
  wire [0:0] u_cla32_and141;
  wire [0:0] u_cla32_or69;
  wire [0:0] u_cla32_or70;
  wire [0:0] u_cla32_or71;
  wire [0:0] u_cla32_pg_logic31_or0;
  wire [0:0] u_cla32_pg_logic31_and0;
  wire [0:0] u_cla32_pg_logic31_xor0;
  wire [0:0] u_cla32_xor31;
  wire [0:0] u_cla32_and142;
  wire [0:0] u_cla32_and143;
  wire [0:0] u_cla32_and144;
  wire [0:0] u_cla32_and145;
  wire [0:0] u_cla32_and146;
  wire [0:0] u_cla32_and147;
  wire [0:0] u_cla32_and148;
  wire [0:0] u_cla32_and149;
  wire [0:0] u_cla32_and150;
  wire [0:0] u_cla32_and151;
  wire [0:0] u_cla32_or72;
  wire [0:0] u_cla32_or73;
  wire [0:0] u_cla32_or74;
  wire [0:0] u_cla32_or75;

  pg_logic pg_logic_u_cla32_pg_logic0_out(.a(a[0]), .b(b[0]), .pg_logic_or0(u_cla32_pg_logic0_or0), .pg_logic_and0(u_cla32_pg_logic0_and0), .pg_logic_xor0(u_cla32_pg_logic0_xor0));
  pg_logic pg_logic_u_cla32_pg_logic1_out(.a(a[1]), .b(b[1]), .pg_logic_or0(u_cla32_pg_logic1_or0), .pg_logic_and0(u_cla32_pg_logic1_and0), .pg_logic_xor0(u_cla32_pg_logic1_xor0));
  xor_gate xor_gate_u_cla32_xor1(.a(u_cla32_pg_logic1_xor0[0]), .b(u_cla32_pg_logic0_and0[0]), .out(u_cla32_xor1));
  and_gate and_gate_u_cla32_and0(.a(u_cla32_pg_logic0_and0[0]), .b(u_cla32_pg_logic1_or0[0]), .out(u_cla32_and0));
  or_gate or_gate_u_cla32_or0(.a(u_cla32_pg_logic1_and0[0]), .b(u_cla32_and0[0]), .out(u_cla32_or0));
  pg_logic pg_logic_u_cla32_pg_logic2_out(.a(a[2]), .b(b[2]), .pg_logic_or0(u_cla32_pg_logic2_or0), .pg_logic_and0(u_cla32_pg_logic2_and0), .pg_logic_xor0(u_cla32_pg_logic2_xor0));
  xor_gate xor_gate_u_cla32_xor2(.a(u_cla32_pg_logic2_xor0[0]), .b(u_cla32_or0[0]), .out(u_cla32_xor2));
  and_gate and_gate_u_cla32_and1(.a(u_cla32_pg_logic2_or0[0]), .b(u_cla32_pg_logic0_or0[0]), .out(u_cla32_and1));
  and_gate and_gate_u_cla32_and2(.a(u_cla32_pg_logic0_and0[0]), .b(u_cla32_pg_logic2_or0[0]), .out(u_cla32_and2));
  and_gate and_gate_u_cla32_and3(.a(u_cla32_and2[0]), .b(u_cla32_pg_logic1_or0[0]), .out(u_cla32_and3));
  and_gate and_gate_u_cla32_and4(.a(u_cla32_pg_logic1_and0[0]), .b(u_cla32_pg_logic2_or0[0]), .out(u_cla32_and4));
  or_gate or_gate_u_cla32_or1(.a(u_cla32_and3[0]), .b(u_cla32_and4[0]), .out(u_cla32_or1));
  or_gate or_gate_u_cla32_or2(.a(u_cla32_pg_logic2_and0[0]), .b(u_cla32_or1[0]), .out(u_cla32_or2));
  pg_logic pg_logic_u_cla32_pg_logic3_out(.a(a[3]), .b(b[3]), .pg_logic_or0(u_cla32_pg_logic3_or0), .pg_logic_and0(u_cla32_pg_logic3_and0), .pg_logic_xor0(u_cla32_pg_logic3_xor0));
  xor_gate xor_gate_u_cla32_xor3(.a(u_cla32_pg_logic3_xor0[0]), .b(u_cla32_or2[0]), .out(u_cla32_xor3));
  and_gate and_gate_u_cla32_and5(.a(u_cla32_pg_logic3_or0[0]), .b(u_cla32_pg_logic1_or0[0]), .out(u_cla32_and5));
  and_gate and_gate_u_cla32_and6(.a(u_cla32_pg_logic0_and0[0]), .b(u_cla32_pg_logic2_or0[0]), .out(u_cla32_and6));
  and_gate and_gate_u_cla32_and7(.a(u_cla32_pg_logic3_or0[0]), .b(u_cla32_pg_logic1_or0[0]), .out(u_cla32_and7));
  and_gate and_gate_u_cla32_and8(.a(u_cla32_and6[0]), .b(u_cla32_and7[0]), .out(u_cla32_and8));
  and_gate and_gate_u_cla32_and9(.a(u_cla32_pg_logic1_and0[0]), .b(u_cla32_pg_logic3_or0[0]), .out(u_cla32_and9));
  and_gate and_gate_u_cla32_and10(.a(u_cla32_and9[0]), .b(u_cla32_pg_logic2_or0[0]), .out(u_cla32_and10));
  and_gate and_gate_u_cla32_and11(.a(u_cla32_pg_logic2_and0[0]), .b(u_cla32_pg_logic3_or0[0]), .out(u_cla32_and11));
  or_gate or_gate_u_cla32_or3(.a(u_cla32_and8[0]), .b(u_cla32_and11[0]), .out(u_cla32_or3));
  or_gate or_gate_u_cla32_or4(.a(u_cla32_and10[0]), .b(u_cla32_or3[0]), .out(u_cla32_or4));
  or_gate or_gate_u_cla32_or5(.a(u_cla32_pg_logic3_and0[0]), .b(u_cla32_or4[0]), .out(u_cla32_or5));
  pg_logic pg_logic_u_cla32_pg_logic4_out(.a(a[4]), .b(b[4]), .pg_logic_or0(u_cla32_pg_logic4_or0), .pg_logic_and0(u_cla32_pg_logic4_and0), .pg_logic_xor0(u_cla32_pg_logic4_xor0));
  xor_gate xor_gate_u_cla32_xor4(.a(u_cla32_pg_logic4_xor0[0]), .b(u_cla32_or5[0]), .out(u_cla32_xor4));
  and_gate and_gate_u_cla32_and12(.a(u_cla32_or5[0]), .b(u_cla32_pg_logic4_or0[0]), .out(u_cla32_and12));
  or_gate or_gate_u_cla32_or6(.a(u_cla32_pg_logic4_and0[0]), .b(u_cla32_and12[0]), .out(u_cla32_or6));
  pg_logic pg_logic_u_cla32_pg_logic5_out(.a(a[5]), .b(b[5]), .pg_logic_or0(u_cla32_pg_logic5_or0), .pg_logic_and0(u_cla32_pg_logic5_and0), .pg_logic_xor0(u_cla32_pg_logic5_xor0));
  xor_gate xor_gate_u_cla32_xor5(.a(u_cla32_pg_logic5_xor0[0]), .b(u_cla32_or6[0]), .out(u_cla32_xor5));
  and_gate and_gate_u_cla32_and13(.a(u_cla32_or5[0]), .b(u_cla32_pg_logic5_or0[0]), .out(u_cla32_and13));
  and_gate and_gate_u_cla32_and14(.a(u_cla32_and13[0]), .b(u_cla32_pg_logic4_or0[0]), .out(u_cla32_and14));
  and_gate and_gate_u_cla32_and15(.a(u_cla32_pg_logic4_and0[0]), .b(u_cla32_pg_logic5_or0[0]), .out(u_cla32_and15));
  or_gate or_gate_u_cla32_or7(.a(u_cla32_and14[0]), .b(u_cla32_and15[0]), .out(u_cla32_or7));
  or_gate or_gate_u_cla32_or8(.a(u_cla32_pg_logic5_and0[0]), .b(u_cla32_or7[0]), .out(u_cla32_or8));
  pg_logic pg_logic_u_cla32_pg_logic6_out(.a(a[6]), .b(b[6]), .pg_logic_or0(u_cla32_pg_logic6_or0), .pg_logic_and0(u_cla32_pg_logic6_and0), .pg_logic_xor0(u_cla32_pg_logic6_xor0));
  xor_gate xor_gate_u_cla32_xor6(.a(u_cla32_pg_logic6_xor0[0]), .b(u_cla32_or8[0]), .out(u_cla32_xor6));
  and_gate and_gate_u_cla32_and16(.a(u_cla32_or5[0]), .b(u_cla32_pg_logic5_or0[0]), .out(u_cla32_and16));
  and_gate and_gate_u_cla32_and17(.a(u_cla32_pg_logic6_or0[0]), .b(u_cla32_pg_logic4_or0[0]), .out(u_cla32_and17));
  and_gate and_gate_u_cla32_and18(.a(u_cla32_and16[0]), .b(u_cla32_and17[0]), .out(u_cla32_and18));
  and_gate and_gate_u_cla32_and19(.a(u_cla32_pg_logic4_and0[0]), .b(u_cla32_pg_logic6_or0[0]), .out(u_cla32_and19));
  and_gate and_gate_u_cla32_and20(.a(u_cla32_and19[0]), .b(u_cla32_pg_logic5_or0[0]), .out(u_cla32_and20));
  and_gate and_gate_u_cla32_and21(.a(u_cla32_pg_logic5_and0[0]), .b(u_cla32_pg_logic6_or0[0]), .out(u_cla32_and21));
  or_gate or_gate_u_cla32_or9(.a(u_cla32_and18[0]), .b(u_cla32_and20[0]), .out(u_cla32_or9));
  or_gate or_gate_u_cla32_or10(.a(u_cla32_or9[0]), .b(u_cla32_and21[0]), .out(u_cla32_or10));
  or_gate or_gate_u_cla32_or11(.a(u_cla32_pg_logic6_and0[0]), .b(u_cla32_or10[0]), .out(u_cla32_or11));
  pg_logic pg_logic_u_cla32_pg_logic7_out(.a(a[7]), .b(b[7]), .pg_logic_or0(u_cla32_pg_logic7_or0), .pg_logic_and0(u_cla32_pg_logic7_and0), .pg_logic_xor0(u_cla32_pg_logic7_xor0));
  xor_gate xor_gate_u_cla32_xor7(.a(u_cla32_pg_logic7_xor0[0]), .b(u_cla32_or11[0]), .out(u_cla32_xor7));
  and_gate and_gate_u_cla32_and22(.a(u_cla32_or5[0]), .b(u_cla32_pg_logic6_or0[0]), .out(u_cla32_and22));
  and_gate and_gate_u_cla32_and23(.a(u_cla32_pg_logic7_or0[0]), .b(u_cla32_pg_logic5_or0[0]), .out(u_cla32_and23));
  and_gate and_gate_u_cla32_and24(.a(u_cla32_and22[0]), .b(u_cla32_and23[0]), .out(u_cla32_and24));
  and_gate and_gate_u_cla32_and25(.a(u_cla32_and24[0]), .b(u_cla32_pg_logic4_or0[0]), .out(u_cla32_and25));
  and_gate and_gate_u_cla32_and26(.a(u_cla32_pg_logic4_and0[0]), .b(u_cla32_pg_logic6_or0[0]), .out(u_cla32_and26));
  and_gate and_gate_u_cla32_and27(.a(u_cla32_pg_logic7_or0[0]), .b(u_cla32_pg_logic5_or0[0]), .out(u_cla32_and27));
  and_gate and_gate_u_cla32_and28(.a(u_cla32_and26[0]), .b(u_cla32_and27[0]), .out(u_cla32_and28));
  and_gate and_gate_u_cla32_and29(.a(u_cla32_pg_logic5_and0[0]), .b(u_cla32_pg_logic7_or0[0]), .out(u_cla32_and29));
  and_gate and_gate_u_cla32_and30(.a(u_cla32_and29[0]), .b(u_cla32_pg_logic6_or0[0]), .out(u_cla32_and30));
  and_gate and_gate_u_cla32_and31(.a(u_cla32_pg_logic6_and0[0]), .b(u_cla32_pg_logic7_or0[0]), .out(u_cla32_and31));
  or_gate or_gate_u_cla32_or12(.a(u_cla32_and25[0]), .b(u_cla32_and30[0]), .out(u_cla32_or12));
  or_gate or_gate_u_cla32_or13(.a(u_cla32_and28[0]), .b(u_cla32_and31[0]), .out(u_cla32_or13));
  or_gate or_gate_u_cla32_or14(.a(u_cla32_or12[0]), .b(u_cla32_or13[0]), .out(u_cla32_or14));
  or_gate or_gate_u_cla32_or15(.a(u_cla32_pg_logic7_and0[0]), .b(u_cla32_or14[0]), .out(u_cla32_or15));
  pg_logic pg_logic_u_cla32_pg_logic8_out(.a(a[8]), .b(b[8]), .pg_logic_or0(u_cla32_pg_logic8_or0), .pg_logic_and0(u_cla32_pg_logic8_and0), .pg_logic_xor0(u_cla32_pg_logic8_xor0));
  xor_gate xor_gate_u_cla32_xor8(.a(u_cla32_pg_logic8_xor0[0]), .b(u_cla32_or15[0]), .out(u_cla32_xor8));
  and_gate and_gate_u_cla32_and32(.a(u_cla32_or15[0]), .b(u_cla32_pg_logic8_or0[0]), .out(u_cla32_and32));
  or_gate or_gate_u_cla32_or16(.a(u_cla32_pg_logic8_and0[0]), .b(u_cla32_and32[0]), .out(u_cla32_or16));
  pg_logic pg_logic_u_cla32_pg_logic9_out(.a(a[9]), .b(b[9]), .pg_logic_or0(u_cla32_pg_logic9_or0), .pg_logic_and0(u_cla32_pg_logic9_and0), .pg_logic_xor0(u_cla32_pg_logic9_xor0));
  xor_gate xor_gate_u_cla32_xor9(.a(u_cla32_pg_logic9_xor0[0]), .b(u_cla32_or16[0]), .out(u_cla32_xor9));
  and_gate and_gate_u_cla32_and33(.a(u_cla32_or15[0]), .b(u_cla32_pg_logic9_or0[0]), .out(u_cla32_and33));
  and_gate and_gate_u_cla32_and34(.a(u_cla32_and33[0]), .b(u_cla32_pg_logic8_or0[0]), .out(u_cla32_and34));
  and_gate and_gate_u_cla32_and35(.a(u_cla32_pg_logic8_and0[0]), .b(u_cla32_pg_logic9_or0[0]), .out(u_cla32_and35));
  or_gate or_gate_u_cla32_or17(.a(u_cla32_and34[0]), .b(u_cla32_and35[0]), .out(u_cla32_or17));
  or_gate or_gate_u_cla32_or18(.a(u_cla32_pg_logic9_and0[0]), .b(u_cla32_or17[0]), .out(u_cla32_or18));
  pg_logic pg_logic_u_cla32_pg_logic10_out(.a(a[10]), .b(b[10]), .pg_logic_or0(u_cla32_pg_logic10_or0), .pg_logic_and0(u_cla32_pg_logic10_and0), .pg_logic_xor0(u_cla32_pg_logic10_xor0));
  xor_gate xor_gate_u_cla32_xor10(.a(u_cla32_pg_logic10_xor0[0]), .b(u_cla32_or18[0]), .out(u_cla32_xor10));
  and_gate and_gate_u_cla32_and36(.a(u_cla32_or15[0]), .b(u_cla32_pg_logic9_or0[0]), .out(u_cla32_and36));
  and_gate and_gate_u_cla32_and37(.a(u_cla32_pg_logic10_or0[0]), .b(u_cla32_pg_logic8_or0[0]), .out(u_cla32_and37));
  and_gate and_gate_u_cla32_and38(.a(u_cla32_and36[0]), .b(u_cla32_and37[0]), .out(u_cla32_and38));
  and_gate and_gate_u_cla32_and39(.a(u_cla32_pg_logic8_and0[0]), .b(u_cla32_pg_logic10_or0[0]), .out(u_cla32_and39));
  and_gate and_gate_u_cla32_and40(.a(u_cla32_and39[0]), .b(u_cla32_pg_logic9_or0[0]), .out(u_cla32_and40));
  and_gate and_gate_u_cla32_and41(.a(u_cla32_pg_logic9_and0[0]), .b(u_cla32_pg_logic10_or0[0]), .out(u_cla32_and41));
  or_gate or_gate_u_cla32_or19(.a(u_cla32_and38[0]), .b(u_cla32_and40[0]), .out(u_cla32_or19));
  or_gate or_gate_u_cla32_or20(.a(u_cla32_or19[0]), .b(u_cla32_and41[0]), .out(u_cla32_or20));
  or_gate or_gate_u_cla32_or21(.a(u_cla32_pg_logic10_and0[0]), .b(u_cla32_or20[0]), .out(u_cla32_or21));
  pg_logic pg_logic_u_cla32_pg_logic11_out(.a(a[11]), .b(b[11]), .pg_logic_or0(u_cla32_pg_logic11_or0), .pg_logic_and0(u_cla32_pg_logic11_and0), .pg_logic_xor0(u_cla32_pg_logic11_xor0));
  xor_gate xor_gate_u_cla32_xor11(.a(u_cla32_pg_logic11_xor0[0]), .b(u_cla32_or21[0]), .out(u_cla32_xor11));
  and_gate and_gate_u_cla32_and42(.a(u_cla32_or15[0]), .b(u_cla32_pg_logic10_or0[0]), .out(u_cla32_and42));
  and_gate and_gate_u_cla32_and43(.a(u_cla32_pg_logic11_or0[0]), .b(u_cla32_pg_logic9_or0[0]), .out(u_cla32_and43));
  and_gate and_gate_u_cla32_and44(.a(u_cla32_and42[0]), .b(u_cla32_and43[0]), .out(u_cla32_and44));
  and_gate and_gate_u_cla32_and45(.a(u_cla32_and44[0]), .b(u_cla32_pg_logic8_or0[0]), .out(u_cla32_and45));
  and_gate and_gate_u_cla32_and46(.a(u_cla32_pg_logic8_and0[0]), .b(u_cla32_pg_logic10_or0[0]), .out(u_cla32_and46));
  and_gate and_gate_u_cla32_and47(.a(u_cla32_pg_logic11_or0[0]), .b(u_cla32_pg_logic9_or0[0]), .out(u_cla32_and47));
  and_gate and_gate_u_cla32_and48(.a(u_cla32_and46[0]), .b(u_cla32_and47[0]), .out(u_cla32_and48));
  and_gate and_gate_u_cla32_and49(.a(u_cla32_pg_logic9_and0[0]), .b(u_cla32_pg_logic11_or0[0]), .out(u_cla32_and49));
  and_gate and_gate_u_cla32_and50(.a(u_cla32_and49[0]), .b(u_cla32_pg_logic10_or0[0]), .out(u_cla32_and50));
  and_gate and_gate_u_cla32_and51(.a(u_cla32_pg_logic10_and0[0]), .b(u_cla32_pg_logic11_or0[0]), .out(u_cla32_and51));
  or_gate or_gate_u_cla32_or22(.a(u_cla32_and45[0]), .b(u_cla32_and50[0]), .out(u_cla32_or22));
  or_gate or_gate_u_cla32_or23(.a(u_cla32_and48[0]), .b(u_cla32_and51[0]), .out(u_cla32_or23));
  or_gate or_gate_u_cla32_or24(.a(u_cla32_or22[0]), .b(u_cla32_or23[0]), .out(u_cla32_or24));
  or_gate or_gate_u_cla32_or25(.a(u_cla32_pg_logic11_and0[0]), .b(u_cla32_or24[0]), .out(u_cla32_or25));
  pg_logic pg_logic_u_cla32_pg_logic12_out(.a(a[12]), .b(b[12]), .pg_logic_or0(u_cla32_pg_logic12_or0), .pg_logic_and0(u_cla32_pg_logic12_and0), .pg_logic_xor0(u_cla32_pg_logic12_xor0));
  xor_gate xor_gate_u_cla32_xor12(.a(u_cla32_pg_logic12_xor0[0]), .b(u_cla32_or25[0]), .out(u_cla32_xor12));
  and_gate and_gate_u_cla32_and52(.a(u_cla32_or25[0]), .b(u_cla32_pg_logic12_or0[0]), .out(u_cla32_and52));
  or_gate or_gate_u_cla32_or26(.a(u_cla32_pg_logic12_and0[0]), .b(u_cla32_and52[0]), .out(u_cla32_or26));
  pg_logic pg_logic_u_cla32_pg_logic13_out(.a(a[13]), .b(b[13]), .pg_logic_or0(u_cla32_pg_logic13_or0), .pg_logic_and0(u_cla32_pg_logic13_and0), .pg_logic_xor0(u_cla32_pg_logic13_xor0));
  xor_gate xor_gate_u_cla32_xor13(.a(u_cla32_pg_logic13_xor0[0]), .b(u_cla32_or26[0]), .out(u_cla32_xor13));
  and_gate and_gate_u_cla32_and53(.a(u_cla32_or25[0]), .b(u_cla32_pg_logic13_or0[0]), .out(u_cla32_and53));
  and_gate and_gate_u_cla32_and54(.a(u_cla32_and53[0]), .b(u_cla32_pg_logic12_or0[0]), .out(u_cla32_and54));
  and_gate and_gate_u_cla32_and55(.a(u_cla32_pg_logic12_and0[0]), .b(u_cla32_pg_logic13_or0[0]), .out(u_cla32_and55));
  or_gate or_gate_u_cla32_or27(.a(u_cla32_and54[0]), .b(u_cla32_and55[0]), .out(u_cla32_or27));
  or_gate or_gate_u_cla32_or28(.a(u_cla32_pg_logic13_and0[0]), .b(u_cla32_or27[0]), .out(u_cla32_or28));
  pg_logic pg_logic_u_cla32_pg_logic14_out(.a(a[14]), .b(b[14]), .pg_logic_or0(u_cla32_pg_logic14_or0), .pg_logic_and0(u_cla32_pg_logic14_and0), .pg_logic_xor0(u_cla32_pg_logic14_xor0));
  xor_gate xor_gate_u_cla32_xor14(.a(u_cla32_pg_logic14_xor0[0]), .b(u_cla32_or28[0]), .out(u_cla32_xor14));
  and_gate and_gate_u_cla32_and56(.a(u_cla32_or25[0]), .b(u_cla32_pg_logic13_or0[0]), .out(u_cla32_and56));
  and_gate and_gate_u_cla32_and57(.a(u_cla32_pg_logic14_or0[0]), .b(u_cla32_pg_logic12_or0[0]), .out(u_cla32_and57));
  and_gate and_gate_u_cla32_and58(.a(u_cla32_and56[0]), .b(u_cla32_and57[0]), .out(u_cla32_and58));
  and_gate and_gate_u_cla32_and59(.a(u_cla32_pg_logic12_and0[0]), .b(u_cla32_pg_logic14_or0[0]), .out(u_cla32_and59));
  and_gate and_gate_u_cla32_and60(.a(u_cla32_and59[0]), .b(u_cla32_pg_logic13_or0[0]), .out(u_cla32_and60));
  and_gate and_gate_u_cla32_and61(.a(u_cla32_pg_logic13_and0[0]), .b(u_cla32_pg_logic14_or0[0]), .out(u_cla32_and61));
  or_gate or_gate_u_cla32_or29(.a(u_cla32_and58[0]), .b(u_cla32_and60[0]), .out(u_cla32_or29));
  or_gate or_gate_u_cla32_or30(.a(u_cla32_or29[0]), .b(u_cla32_and61[0]), .out(u_cla32_or30));
  or_gate or_gate_u_cla32_or31(.a(u_cla32_pg_logic14_and0[0]), .b(u_cla32_or30[0]), .out(u_cla32_or31));
  pg_logic pg_logic_u_cla32_pg_logic15_out(.a(a[15]), .b(b[15]), .pg_logic_or0(u_cla32_pg_logic15_or0), .pg_logic_and0(u_cla32_pg_logic15_and0), .pg_logic_xor0(u_cla32_pg_logic15_xor0));
  xor_gate xor_gate_u_cla32_xor15(.a(u_cla32_pg_logic15_xor0[0]), .b(u_cla32_or31[0]), .out(u_cla32_xor15));
  and_gate and_gate_u_cla32_and62(.a(u_cla32_or25[0]), .b(u_cla32_pg_logic14_or0[0]), .out(u_cla32_and62));
  and_gate and_gate_u_cla32_and63(.a(u_cla32_pg_logic15_or0[0]), .b(u_cla32_pg_logic13_or0[0]), .out(u_cla32_and63));
  and_gate and_gate_u_cla32_and64(.a(u_cla32_and62[0]), .b(u_cla32_and63[0]), .out(u_cla32_and64));
  and_gate and_gate_u_cla32_and65(.a(u_cla32_and64[0]), .b(u_cla32_pg_logic12_or0[0]), .out(u_cla32_and65));
  and_gate and_gate_u_cla32_and66(.a(u_cla32_pg_logic12_and0[0]), .b(u_cla32_pg_logic14_or0[0]), .out(u_cla32_and66));
  and_gate and_gate_u_cla32_and67(.a(u_cla32_pg_logic15_or0[0]), .b(u_cla32_pg_logic13_or0[0]), .out(u_cla32_and67));
  and_gate and_gate_u_cla32_and68(.a(u_cla32_and66[0]), .b(u_cla32_and67[0]), .out(u_cla32_and68));
  and_gate and_gate_u_cla32_and69(.a(u_cla32_pg_logic13_and0[0]), .b(u_cla32_pg_logic15_or0[0]), .out(u_cla32_and69));
  and_gate and_gate_u_cla32_and70(.a(u_cla32_and69[0]), .b(u_cla32_pg_logic14_or0[0]), .out(u_cla32_and70));
  and_gate and_gate_u_cla32_and71(.a(u_cla32_pg_logic14_and0[0]), .b(u_cla32_pg_logic15_or0[0]), .out(u_cla32_and71));
  or_gate or_gate_u_cla32_or32(.a(u_cla32_and65[0]), .b(u_cla32_and70[0]), .out(u_cla32_or32));
  or_gate or_gate_u_cla32_or33(.a(u_cla32_and68[0]), .b(u_cla32_and71[0]), .out(u_cla32_or33));
  or_gate or_gate_u_cla32_or34(.a(u_cla32_or32[0]), .b(u_cla32_or33[0]), .out(u_cla32_or34));
  or_gate or_gate_u_cla32_or35(.a(u_cla32_pg_logic15_and0[0]), .b(u_cla32_or34[0]), .out(u_cla32_or35));
  pg_logic pg_logic_u_cla32_pg_logic16_out(.a(a[16]), .b(b[16]), .pg_logic_or0(u_cla32_pg_logic16_or0), .pg_logic_and0(u_cla32_pg_logic16_and0), .pg_logic_xor0(u_cla32_pg_logic16_xor0));
  xor_gate xor_gate_u_cla32_xor16(.a(u_cla32_pg_logic16_xor0[0]), .b(u_cla32_or35[0]), .out(u_cla32_xor16));
  and_gate and_gate_u_cla32_and72(.a(u_cla32_or35[0]), .b(u_cla32_pg_logic16_or0[0]), .out(u_cla32_and72));
  or_gate or_gate_u_cla32_or36(.a(u_cla32_pg_logic16_and0[0]), .b(u_cla32_and72[0]), .out(u_cla32_or36));
  pg_logic pg_logic_u_cla32_pg_logic17_out(.a(a[17]), .b(b[17]), .pg_logic_or0(u_cla32_pg_logic17_or0), .pg_logic_and0(u_cla32_pg_logic17_and0), .pg_logic_xor0(u_cla32_pg_logic17_xor0));
  xor_gate xor_gate_u_cla32_xor17(.a(u_cla32_pg_logic17_xor0[0]), .b(u_cla32_or36[0]), .out(u_cla32_xor17));
  and_gate and_gate_u_cla32_and73(.a(u_cla32_or35[0]), .b(u_cla32_pg_logic17_or0[0]), .out(u_cla32_and73));
  and_gate and_gate_u_cla32_and74(.a(u_cla32_and73[0]), .b(u_cla32_pg_logic16_or0[0]), .out(u_cla32_and74));
  and_gate and_gate_u_cla32_and75(.a(u_cla32_pg_logic16_and0[0]), .b(u_cla32_pg_logic17_or0[0]), .out(u_cla32_and75));
  or_gate or_gate_u_cla32_or37(.a(u_cla32_and74[0]), .b(u_cla32_and75[0]), .out(u_cla32_or37));
  or_gate or_gate_u_cla32_or38(.a(u_cla32_pg_logic17_and0[0]), .b(u_cla32_or37[0]), .out(u_cla32_or38));
  pg_logic pg_logic_u_cla32_pg_logic18_out(.a(a[18]), .b(b[18]), .pg_logic_or0(u_cla32_pg_logic18_or0), .pg_logic_and0(u_cla32_pg_logic18_and0), .pg_logic_xor0(u_cla32_pg_logic18_xor0));
  xor_gate xor_gate_u_cla32_xor18(.a(u_cla32_pg_logic18_xor0[0]), .b(u_cla32_or38[0]), .out(u_cla32_xor18));
  and_gate and_gate_u_cla32_and76(.a(u_cla32_or35[0]), .b(u_cla32_pg_logic17_or0[0]), .out(u_cla32_and76));
  and_gate and_gate_u_cla32_and77(.a(u_cla32_pg_logic18_or0[0]), .b(u_cla32_pg_logic16_or0[0]), .out(u_cla32_and77));
  and_gate and_gate_u_cla32_and78(.a(u_cla32_and76[0]), .b(u_cla32_and77[0]), .out(u_cla32_and78));
  and_gate and_gate_u_cla32_and79(.a(u_cla32_pg_logic16_and0[0]), .b(u_cla32_pg_logic18_or0[0]), .out(u_cla32_and79));
  and_gate and_gate_u_cla32_and80(.a(u_cla32_and79[0]), .b(u_cla32_pg_logic17_or0[0]), .out(u_cla32_and80));
  and_gate and_gate_u_cla32_and81(.a(u_cla32_pg_logic17_and0[0]), .b(u_cla32_pg_logic18_or0[0]), .out(u_cla32_and81));
  or_gate or_gate_u_cla32_or39(.a(u_cla32_and78[0]), .b(u_cla32_and80[0]), .out(u_cla32_or39));
  or_gate or_gate_u_cla32_or40(.a(u_cla32_or39[0]), .b(u_cla32_and81[0]), .out(u_cla32_or40));
  or_gate or_gate_u_cla32_or41(.a(u_cla32_pg_logic18_and0[0]), .b(u_cla32_or40[0]), .out(u_cla32_or41));
  pg_logic pg_logic_u_cla32_pg_logic19_out(.a(a[19]), .b(b[19]), .pg_logic_or0(u_cla32_pg_logic19_or0), .pg_logic_and0(u_cla32_pg_logic19_and0), .pg_logic_xor0(u_cla32_pg_logic19_xor0));
  xor_gate xor_gate_u_cla32_xor19(.a(u_cla32_pg_logic19_xor0[0]), .b(u_cla32_or41[0]), .out(u_cla32_xor19));
  and_gate and_gate_u_cla32_and82(.a(u_cla32_or35[0]), .b(u_cla32_pg_logic18_or0[0]), .out(u_cla32_and82));
  and_gate and_gate_u_cla32_and83(.a(u_cla32_pg_logic19_or0[0]), .b(u_cla32_pg_logic17_or0[0]), .out(u_cla32_and83));
  and_gate and_gate_u_cla32_and84(.a(u_cla32_and82[0]), .b(u_cla32_and83[0]), .out(u_cla32_and84));
  and_gate and_gate_u_cla32_and85(.a(u_cla32_and84[0]), .b(u_cla32_pg_logic16_or0[0]), .out(u_cla32_and85));
  and_gate and_gate_u_cla32_and86(.a(u_cla32_pg_logic16_and0[0]), .b(u_cla32_pg_logic18_or0[0]), .out(u_cla32_and86));
  and_gate and_gate_u_cla32_and87(.a(u_cla32_pg_logic19_or0[0]), .b(u_cla32_pg_logic17_or0[0]), .out(u_cla32_and87));
  and_gate and_gate_u_cla32_and88(.a(u_cla32_and86[0]), .b(u_cla32_and87[0]), .out(u_cla32_and88));
  and_gate and_gate_u_cla32_and89(.a(u_cla32_pg_logic17_and0[0]), .b(u_cla32_pg_logic19_or0[0]), .out(u_cla32_and89));
  and_gate and_gate_u_cla32_and90(.a(u_cla32_and89[0]), .b(u_cla32_pg_logic18_or0[0]), .out(u_cla32_and90));
  and_gate and_gate_u_cla32_and91(.a(u_cla32_pg_logic18_and0[0]), .b(u_cla32_pg_logic19_or0[0]), .out(u_cla32_and91));
  or_gate or_gate_u_cla32_or42(.a(u_cla32_and85[0]), .b(u_cla32_and90[0]), .out(u_cla32_or42));
  or_gate or_gate_u_cla32_or43(.a(u_cla32_and88[0]), .b(u_cla32_and91[0]), .out(u_cla32_or43));
  or_gate or_gate_u_cla32_or44(.a(u_cla32_or42[0]), .b(u_cla32_or43[0]), .out(u_cla32_or44));
  or_gate or_gate_u_cla32_or45(.a(u_cla32_pg_logic19_and0[0]), .b(u_cla32_or44[0]), .out(u_cla32_or45));
  pg_logic pg_logic_u_cla32_pg_logic20_out(.a(a[20]), .b(b[20]), .pg_logic_or0(u_cla32_pg_logic20_or0), .pg_logic_and0(u_cla32_pg_logic20_and0), .pg_logic_xor0(u_cla32_pg_logic20_xor0));
  xor_gate xor_gate_u_cla32_xor20(.a(u_cla32_pg_logic20_xor0[0]), .b(u_cla32_or45[0]), .out(u_cla32_xor20));
  and_gate and_gate_u_cla32_and92(.a(u_cla32_or45[0]), .b(u_cla32_pg_logic20_or0[0]), .out(u_cla32_and92));
  or_gate or_gate_u_cla32_or46(.a(u_cla32_pg_logic20_and0[0]), .b(u_cla32_and92[0]), .out(u_cla32_or46));
  pg_logic pg_logic_u_cla32_pg_logic21_out(.a(a[21]), .b(b[21]), .pg_logic_or0(u_cla32_pg_logic21_or0), .pg_logic_and0(u_cla32_pg_logic21_and0), .pg_logic_xor0(u_cla32_pg_logic21_xor0));
  xor_gate xor_gate_u_cla32_xor21(.a(u_cla32_pg_logic21_xor0[0]), .b(u_cla32_or46[0]), .out(u_cla32_xor21));
  and_gate and_gate_u_cla32_and93(.a(u_cla32_or45[0]), .b(u_cla32_pg_logic21_or0[0]), .out(u_cla32_and93));
  and_gate and_gate_u_cla32_and94(.a(u_cla32_and93[0]), .b(u_cla32_pg_logic20_or0[0]), .out(u_cla32_and94));
  and_gate and_gate_u_cla32_and95(.a(u_cla32_pg_logic20_and0[0]), .b(u_cla32_pg_logic21_or0[0]), .out(u_cla32_and95));
  or_gate or_gate_u_cla32_or47(.a(u_cla32_and94[0]), .b(u_cla32_and95[0]), .out(u_cla32_or47));
  or_gate or_gate_u_cla32_or48(.a(u_cla32_pg_logic21_and0[0]), .b(u_cla32_or47[0]), .out(u_cla32_or48));
  pg_logic pg_logic_u_cla32_pg_logic22_out(.a(a[22]), .b(b[22]), .pg_logic_or0(u_cla32_pg_logic22_or0), .pg_logic_and0(u_cla32_pg_logic22_and0), .pg_logic_xor0(u_cla32_pg_logic22_xor0));
  xor_gate xor_gate_u_cla32_xor22(.a(u_cla32_pg_logic22_xor0[0]), .b(u_cla32_or48[0]), .out(u_cla32_xor22));
  and_gate and_gate_u_cla32_and96(.a(u_cla32_or45[0]), .b(u_cla32_pg_logic21_or0[0]), .out(u_cla32_and96));
  and_gate and_gate_u_cla32_and97(.a(u_cla32_pg_logic22_or0[0]), .b(u_cla32_pg_logic20_or0[0]), .out(u_cla32_and97));
  and_gate and_gate_u_cla32_and98(.a(u_cla32_and96[0]), .b(u_cla32_and97[0]), .out(u_cla32_and98));
  and_gate and_gate_u_cla32_and99(.a(u_cla32_pg_logic20_and0[0]), .b(u_cla32_pg_logic22_or0[0]), .out(u_cla32_and99));
  and_gate and_gate_u_cla32_and100(.a(u_cla32_and99[0]), .b(u_cla32_pg_logic21_or0[0]), .out(u_cla32_and100));
  and_gate and_gate_u_cla32_and101(.a(u_cla32_pg_logic21_and0[0]), .b(u_cla32_pg_logic22_or0[0]), .out(u_cla32_and101));
  or_gate or_gate_u_cla32_or49(.a(u_cla32_and98[0]), .b(u_cla32_and100[0]), .out(u_cla32_or49));
  or_gate or_gate_u_cla32_or50(.a(u_cla32_or49[0]), .b(u_cla32_and101[0]), .out(u_cla32_or50));
  or_gate or_gate_u_cla32_or51(.a(u_cla32_pg_logic22_and0[0]), .b(u_cla32_or50[0]), .out(u_cla32_or51));
  pg_logic pg_logic_u_cla32_pg_logic23_out(.a(a[23]), .b(b[23]), .pg_logic_or0(u_cla32_pg_logic23_or0), .pg_logic_and0(u_cla32_pg_logic23_and0), .pg_logic_xor0(u_cla32_pg_logic23_xor0));
  xor_gate xor_gate_u_cla32_xor23(.a(u_cla32_pg_logic23_xor0[0]), .b(u_cla32_or51[0]), .out(u_cla32_xor23));
  and_gate and_gate_u_cla32_and102(.a(u_cla32_or45[0]), .b(u_cla32_pg_logic22_or0[0]), .out(u_cla32_and102));
  and_gate and_gate_u_cla32_and103(.a(u_cla32_pg_logic23_or0[0]), .b(u_cla32_pg_logic21_or0[0]), .out(u_cla32_and103));
  and_gate and_gate_u_cla32_and104(.a(u_cla32_and102[0]), .b(u_cla32_and103[0]), .out(u_cla32_and104));
  and_gate and_gate_u_cla32_and105(.a(u_cla32_and104[0]), .b(u_cla32_pg_logic20_or0[0]), .out(u_cla32_and105));
  and_gate and_gate_u_cla32_and106(.a(u_cla32_pg_logic20_and0[0]), .b(u_cla32_pg_logic22_or0[0]), .out(u_cla32_and106));
  and_gate and_gate_u_cla32_and107(.a(u_cla32_pg_logic23_or0[0]), .b(u_cla32_pg_logic21_or0[0]), .out(u_cla32_and107));
  and_gate and_gate_u_cla32_and108(.a(u_cla32_and106[0]), .b(u_cla32_and107[0]), .out(u_cla32_and108));
  and_gate and_gate_u_cla32_and109(.a(u_cla32_pg_logic21_and0[0]), .b(u_cla32_pg_logic23_or0[0]), .out(u_cla32_and109));
  and_gate and_gate_u_cla32_and110(.a(u_cla32_and109[0]), .b(u_cla32_pg_logic22_or0[0]), .out(u_cla32_and110));
  and_gate and_gate_u_cla32_and111(.a(u_cla32_pg_logic22_and0[0]), .b(u_cla32_pg_logic23_or0[0]), .out(u_cla32_and111));
  or_gate or_gate_u_cla32_or52(.a(u_cla32_and105[0]), .b(u_cla32_and110[0]), .out(u_cla32_or52));
  or_gate or_gate_u_cla32_or53(.a(u_cla32_and108[0]), .b(u_cla32_and111[0]), .out(u_cla32_or53));
  or_gate or_gate_u_cla32_or54(.a(u_cla32_or52[0]), .b(u_cla32_or53[0]), .out(u_cla32_or54));
  or_gate or_gate_u_cla32_or55(.a(u_cla32_pg_logic23_and0[0]), .b(u_cla32_or54[0]), .out(u_cla32_or55));
  pg_logic pg_logic_u_cla32_pg_logic24_out(.a(a[24]), .b(b[24]), .pg_logic_or0(u_cla32_pg_logic24_or0), .pg_logic_and0(u_cla32_pg_logic24_and0), .pg_logic_xor0(u_cla32_pg_logic24_xor0));
  xor_gate xor_gate_u_cla32_xor24(.a(u_cla32_pg_logic24_xor0[0]), .b(u_cla32_or55[0]), .out(u_cla32_xor24));
  and_gate and_gate_u_cla32_and112(.a(u_cla32_or55[0]), .b(u_cla32_pg_logic24_or0[0]), .out(u_cla32_and112));
  or_gate or_gate_u_cla32_or56(.a(u_cla32_pg_logic24_and0[0]), .b(u_cla32_and112[0]), .out(u_cla32_or56));
  pg_logic pg_logic_u_cla32_pg_logic25_out(.a(a[25]), .b(b[25]), .pg_logic_or0(u_cla32_pg_logic25_or0), .pg_logic_and0(u_cla32_pg_logic25_and0), .pg_logic_xor0(u_cla32_pg_logic25_xor0));
  xor_gate xor_gate_u_cla32_xor25(.a(u_cla32_pg_logic25_xor0[0]), .b(u_cla32_or56[0]), .out(u_cla32_xor25));
  and_gate and_gate_u_cla32_and113(.a(u_cla32_or55[0]), .b(u_cla32_pg_logic25_or0[0]), .out(u_cla32_and113));
  and_gate and_gate_u_cla32_and114(.a(u_cla32_and113[0]), .b(u_cla32_pg_logic24_or0[0]), .out(u_cla32_and114));
  and_gate and_gate_u_cla32_and115(.a(u_cla32_pg_logic24_and0[0]), .b(u_cla32_pg_logic25_or0[0]), .out(u_cla32_and115));
  or_gate or_gate_u_cla32_or57(.a(u_cla32_and114[0]), .b(u_cla32_and115[0]), .out(u_cla32_or57));
  or_gate or_gate_u_cla32_or58(.a(u_cla32_pg_logic25_and0[0]), .b(u_cla32_or57[0]), .out(u_cla32_or58));
  pg_logic pg_logic_u_cla32_pg_logic26_out(.a(a[26]), .b(b[26]), .pg_logic_or0(u_cla32_pg_logic26_or0), .pg_logic_and0(u_cla32_pg_logic26_and0), .pg_logic_xor0(u_cla32_pg_logic26_xor0));
  xor_gate xor_gate_u_cla32_xor26(.a(u_cla32_pg_logic26_xor0[0]), .b(u_cla32_or58[0]), .out(u_cla32_xor26));
  and_gate and_gate_u_cla32_and116(.a(u_cla32_or55[0]), .b(u_cla32_pg_logic25_or0[0]), .out(u_cla32_and116));
  and_gate and_gate_u_cla32_and117(.a(u_cla32_pg_logic26_or0[0]), .b(u_cla32_pg_logic24_or0[0]), .out(u_cla32_and117));
  and_gate and_gate_u_cla32_and118(.a(u_cla32_and116[0]), .b(u_cla32_and117[0]), .out(u_cla32_and118));
  and_gate and_gate_u_cla32_and119(.a(u_cla32_pg_logic24_and0[0]), .b(u_cla32_pg_logic26_or0[0]), .out(u_cla32_and119));
  and_gate and_gate_u_cla32_and120(.a(u_cla32_and119[0]), .b(u_cla32_pg_logic25_or0[0]), .out(u_cla32_and120));
  and_gate and_gate_u_cla32_and121(.a(u_cla32_pg_logic25_and0[0]), .b(u_cla32_pg_logic26_or0[0]), .out(u_cla32_and121));
  or_gate or_gate_u_cla32_or59(.a(u_cla32_and118[0]), .b(u_cla32_and120[0]), .out(u_cla32_or59));
  or_gate or_gate_u_cla32_or60(.a(u_cla32_or59[0]), .b(u_cla32_and121[0]), .out(u_cla32_or60));
  or_gate or_gate_u_cla32_or61(.a(u_cla32_pg_logic26_and0[0]), .b(u_cla32_or60[0]), .out(u_cla32_or61));
  pg_logic pg_logic_u_cla32_pg_logic27_out(.a(a[27]), .b(b[27]), .pg_logic_or0(u_cla32_pg_logic27_or0), .pg_logic_and0(u_cla32_pg_logic27_and0), .pg_logic_xor0(u_cla32_pg_logic27_xor0));
  xor_gate xor_gate_u_cla32_xor27(.a(u_cla32_pg_logic27_xor0[0]), .b(u_cla32_or61[0]), .out(u_cla32_xor27));
  and_gate and_gate_u_cla32_and122(.a(u_cla32_or55[0]), .b(u_cla32_pg_logic26_or0[0]), .out(u_cla32_and122));
  and_gate and_gate_u_cla32_and123(.a(u_cla32_pg_logic27_or0[0]), .b(u_cla32_pg_logic25_or0[0]), .out(u_cla32_and123));
  and_gate and_gate_u_cla32_and124(.a(u_cla32_and122[0]), .b(u_cla32_and123[0]), .out(u_cla32_and124));
  and_gate and_gate_u_cla32_and125(.a(u_cla32_and124[0]), .b(u_cla32_pg_logic24_or0[0]), .out(u_cla32_and125));
  and_gate and_gate_u_cla32_and126(.a(u_cla32_pg_logic24_and0[0]), .b(u_cla32_pg_logic26_or0[0]), .out(u_cla32_and126));
  and_gate and_gate_u_cla32_and127(.a(u_cla32_pg_logic27_or0[0]), .b(u_cla32_pg_logic25_or0[0]), .out(u_cla32_and127));
  and_gate and_gate_u_cla32_and128(.a(u_cla32_and126[0]), .b(u_cla32_and127[0]), .out(u_cla32_and128));
  and_gate and_gate_u_cla32_and129(.a(u_cla32_pg_logic25_and0[0]), .b(u_cla32_pg_logic27_or0[0]), .out(u_cla32_and129));
  and_gate and_gate_u_cla32_and130(.a(u_cla32_and129[0]), .b(u_cla32_pg_logic26_or0[0]), .out(u_cla32_and130));
  and_gate and_gate_u_cla32_and131(.a(u_cla32_pg_logic26_and0[0]), .b(u_cla32_pg_logic27_or0[0]), .out(u_cla32_and131));
  or_gate or_gate_u_cla32_or62(.a(u_cla32_and125[0]), .b(u_cla32_and130[0]), .out(u_cla32_or62));
  or_gate or_gate_u_cla32_or63(.a(u_cla32_and128[0]), .b(u_cla32_and131[0]), .out(u_cla32_or63));
  or_gate or_gate_u_cla32_or64(.a(u_cla32_or62[0]), .b(u_cla32_or63[0]), .out(u_cla32_or64));
  or_gate or_gate_u_cla32_or65(.a(u_cla32_pg_logic27_and0[0]), .b(u_cla32_or64[0]), .out(u_cla32_or65));
  pg_logic pg_logic_u_cla32_pg_logic28_out(.a(a[28]), .b(b[28]), .pg_logic_or0(u_cla32_pg_logic28_or0), .pg_logic_and0(u_cla32_pg_logic28_and0), .pg_logic_xor0(u_cla32_pg_logic28_xor0));
  xor_gate xor_gate_u_cla32_xor28(.a(u_cla32_pg_logic28_xor0[0]), .b(u_cla32_or65[0]), .out(u_cla32_xor28));
  and_gate and_gate_u_cla32_and132(.a(u_cla32_or65[0]), .b(u_cla32_pg_logic28_or0[0]), .out(u_cla32_and132));
  or_gate or_gate_u_cla32_or66(.a(u_cla32_pg_logic28_and0[0]), .b(u_cla32_and132[0]), .out(u_cla32_or66));
  pg_logic pg_logic_u_cla32_pg_logic29_out(.a(a[29]), .b(b[29]), .pg_logic_or0(u_cla32_pg_logic29_or0), .pg_logic_and0(u_cla32_pg_logic29_and0), .pg_logic_xor0(u_cla32_pg_logic29_xor0));
  xor_gate xor_gate_u_cla32_xor29(.a(u_cla32_pg_logic29_xor0[0]), .b(u_cla32_or66[0]), .out(u_cla32_xor29));
  and_gate and_gate_u_cla32_and133(.a(u_cla32_or65[0]), .b(u_cla32_pg_logic29_or0[0]), .out(u_cla32_and133));
  and_gate and_gate_u_cla32_and134(.a(u_cla32_and133[0]), .b(u_cla32_pg_logic28_or0[0]), .out(u_cla32_and134));
  and_gate and_gate_u_cla32_and135(.a(u_cla32_pg_logic28_and0[0]), .b(u_cla32_pg_logic29_or0[0]), .out(u_cla32_and135));
  or_gate or_gate_u_cla32_or67(.a(u_cla32_and134[0]), .b(u_cla32_and135[0]), .out(u_cla32_or67));
  or_gate or_gate_u_cla32_or68(.a(u_cla32_pg_logic29_and0[0]), .b(u_cla32_or67[0]), .out(u_cla32_or68));
  pg_logic pg_logic_u_cla32_pg_logic30_out(.a(a[30]), .b(b[30]), .pg_logic_or0(u_cla32_pg_logic30_or0), .pg_logic_and0(u_cla32_pg_logic30_and0), .pg_logic_xor0(u_cla32_pg_logic30_xor0));
  xor_gate xor_gate_u_cla32_xor30(.a(u_cla32_pg_logic30_xor0[0]), .b(u_cla32_or68[0]), .out(u_cla32_xor30));
  and_gate and_gate_u_cla32_and136(.a(u_cla32_or65[0]), .b(u_cla32_pg_logic29_or0[0]), .out(u_cla32_and136));
  and_gate and_gate_u_cla32_and137(.a(u_cla32_pg_logic30_or0[0]), .b(u_cla32_pg_logic28_or0[0]), .out(u_cla32_and137));
  and_gate and_gate_u_cla32_and138(.a(u_cla32_and136[0]), .b(u_cla32_and137[0]), .out(u_cla32_and138));
  and_gate and_gate_u_cla32_and139(.a(u_cla32_pg_logic28_and0[0]), .b(u_cla32_pg_logic30_or0[0]), .out(u_cla32_and139));
  and_gate and_gate_u_cla32_and140(.a(u_cla32_and139[0]), .b(u_cla32_pg_logic29_or0[0]), .out(u_cla32_and140));
  and_gate and_gate_u_cla32_and141(.a(u_cla32_pg_logic29_and0[0]), .b(u_cla32_pg_logic30_or0[0]), .out(u_cla32_and141));
  or_gate or_gate_u_cla32_or69(.a(u_cla32_and138[0]), .b(u_cla32_and140[0]), .out(u_cla32_or69));
  or_gate or_gate_u_cla32_or70(.a(u_cla32_or69[0]), .b(u_cla32_and141[0]), .out(u_cla32_or70));
  or_gate or_gate_u_cla32_or71(.a(u_cla32_pg_logic30_and0[0]), .b(u_cla32_or70[0]), .out(u_cla32_or71));
  pg_logic pg_logic_u_cla32_pg_logic31_out(.a(a[31]), .b(b[31]), .pg_logic_or0(u_cla32_pg_logic31_or0), .pg_logic_and0(u_cla32_pg_logic31_and0), .pg_logic_xor0(u_cla32_pg_logic31_xor0));
  xor_gate xor_gate_u_cla32_xor31(.a(u_cla32_pg_logic31_xor0[0]), .b(u_cla32_or71[0]), .out(u_cla32_xor31));
  and_gate and_gate_u_cla32_and142(.a(u_cla32_or65[0]), .b(u_cla32_pg_logic30_or0[0]), .out(u_cla32_and142));
  and_gate and_gate_u_cla32_and143(.a(u_cla32_pg_logic31_or0[0]), .b(u_cla32_pg_logic29_or0[0]), .out(u_cla32_and143));
  and_gate and_gate_u_cla32_and144(.a(u_cla32_and142[0]), .b(u_cla32_and143[0]), .out(u_cla32_and144));
  and_gate and_gate_u_cla32_and145(.a(u_cla32_and144[0]), .b(u_cla32_pg_logic28_or0[0]), .out(u_cla32_and145));
  and_gate and_gate_u_cla32_and146(.a(u_cla32_pg_logic28_and0[0]), .b(u_cla32_pg_logic30_or0[0]), .out(u_cla32_and146));
  and_gate and_gate_u_cla32_and147(.a(u_cla32_pg_logic31_or0[0]), .b(u_cla32_pg_logic29_or0[0]), .out(u_cla32_and147));
  and_gate and_gate_u_cla32_and148(.a(u_cla32_and146[0]), .b(u_cla32_and147[0]), .out(u_cla32_and148));
  and_gate and_gate_u_cla32_and149(.a(u_cla32_pg_logic29_and0[0]), .b(u_cla32_pg_logic31_or0[0]), .out(u_cla32_and149));
  and_gate and_gate_u_cla32_and150(.a(u_cla32_and149[0]), .b(u_cla32_pg_logic30_or0[0]), .out(u_cla32_and150));
  and_gate and_gate_u_cla32_and151(.a(u_cla32_pg_logic30_and0[0]), .b(u_cla32_pg_logic31_or0[0]), .out(u_cla32_and151));
  or_gate or_gate_u_cla32_or72(.a(u_cla32_and145[0]), .b(u_cla32_and150[0]), .out(u_cla32_or72));
  or_gate or_gate_u_cla32_or73(.a(u_cla32_and148[0]), .b(u_cla32_and151[0]), .out(u_cla32_or73));
  or_gate or_gate_u_cla32_or74(.a(u_cla32_or72[0]), .b(u_cla32_or73[0]), .out(u_cla32_or74));
  or_gate or_gate_u_cla32_or75(.a(u_cla32_pg_logic31_and0[0]), .b(u_cla32_or74[0]), .out(u_cla32_or75));

  assign u_cla32_out[0] = u_cla32_pg_logic0_xor0[0];
  assign u_cla32_out[1] = u_cla32_xor1[0];
  assign u_cla32_out[2] = u_cla32_xor2[0];
  assign u_cla32_out[3] = u_cla32_xor3[0];
  assign u_cla32_out[4] = u_cla32_xor4[0];
  assign u_cla32_out[5] = u_cla32_xor5[0];
  assign u_cla32_out[6] = u_cla32_xor6[0];
  assign u_cla32_out[7] = u_cla32_xor7[0];
  assign u_cla32_out[8] = u_cla32_xor8[0];
  assign u_cla32_out[9] = u_cla32_xor9[0];
  assign u_cla32_out[10] = u_cla32_xor10[0];
  assign u_cla32_out[11] = u_cla32_xor11[0];
  assign u_cla32_out[12] = u_cla32_xor12[0];
  assign u_cla32_out[13] = u_cla32_xor13[0];
  assign u_cla32_out[14] = u_cla32_xor14[0];
  assign u_cla32_out[15] = u_cla32_xor15[0];
  assign u_cla32_out[16] = u_cla32_xor16[0];
  assign u_cla32_out[17] = u_cla32_xor17[0];
  assign u_cla32_out[18] = u_cla32_xor18[0];
  assign u_cla32_out[19] = u_cla32_xor19[0];
  assign u_cla32_out[20] = u_cla32_xor20[0];
  assign u_cla32_out[21] = u_cla32_xor21[0];
  assign u_cla32_out[22] = u_cla32_xor22[0];
  assign u_cla32_out[23] = u_cla32_xor23[0];
  assign u_cla32_out[24] = u_cla32_xor24[0];
  assign u_cla32_out[25] = u_cla32_xor25[0];
  assign u_cla32_out[26] = u_cla32_xor26[0];
  assign u_cla32_out[27] = u_cla32_xor27[0];
  assign u_cla32_out[28] = u_cla32_xor28[0];
  assign u_cla32_out[29] = u_cla32_xor29[0];
  assign u_cla32_out[30] = u_cla32_xor30[0];
  assign u_cla32_out[31] = u_cla32_xor31[0];
  assign u_cla32_out[32] = u_cla32_or75[0];
endmodule

module u_csamul_cla32(input [31:0] a, input [31:0] b, output [63:0] u_csamul_cla32_out);
  wire [0:0] u_csamul_cla32_and0_0;
  wire [0:0] u_csamul_cla32_and1_0;
  wire [0:0] u_csamul_cla32_and2_0;
  wire [0:0] u_csamul_cla32_and3_0;
  wire [0:0] u_csamul_cla32_and4_0;
  wire [0:0] u_csamul_cla32_and5_0;
  wire [0:0] u_csamul_cla32_and6_0;
  wire [0:0] u_csamul_cla32_and7_0;
  wire [0:0] u_csamul_cla32_and8_0;
  wire [0:0] u_csamul_cla32_and9_0;
  wire [0:0] u_csamul_cla32_and10_0;
  wire [0:0] u_csamul_cla32_and11_0;
  wire [0:0] u_csamul_cla32_and12_0;
  wire [0:0] u_csamul_cla32_and13_0;
  wire [0:0] u_csamul_cla32_and14_0;
  wire [0:0] u_csamul_cla32_and15_0;
  wire [0:0] u_csamul_cla32_and16_0;
  wire [0:0] u_csamul_cla32_and17_0;
  wire [0:0] u_csamul_cla32_and18_0;
  wire [0:0] u_csamul_cla32_and19_0;
  wire [0:0] u_csamul_cla32_and20_0;
  wire [0:0] u_csamul_cla32_and21_0;
  wire [0:0] u_csamul_cla32_and22_0;
  wire [0:0] u_csamul_cla32_and23_0;
  wire [0:0] u_csamul_cla32_and24_0;
  wire [0:0] u_csamul_cla32_and25_0;
  wire [0:0] u_csamul_cla32_and26_0;
  wire [0:0] u_csamul_cla32_and27_0;
  wire [0:0] u_csamul_cla32_and28_0;
  wire [0:0] u_csamul_cla32_and29_0;
  wire [0:0] u_csamul_cla32_and30_0;
  wire [0:0] u_csamul_cla32_and31_0;
  wire [0:0] u_csamul_cla32_and0_1;
  wire [0:0] u_csamul_cla32_ha0_1_xor0;
  wire [0:0] u_csamul_cla32_ha0_1_and0;
  wire [0:0] u_csamul_cla32_and1_1;
  wire [0:0] u_csamul_cla32_ha1_1_xor0;
  wire [0:0] u_csamul_cla32_ha1_1_and0;
  wire [0:0] u_csamul_cla32_and2_1;
  wire [0:0] u_csamul_cla32_ha2_1_xor0;
  wire [0:0] u_csamul_cla32_ha2_1_and0;
  wire [0:0] u_csamul_cla32_and3_1;
  wire [0:0] u_csamul_cla32_ha3_1_xor0;
  wire [0:0] u_csamul_cla32_ha3_1_and0;
  wire [0:0] u_csamul_cla32_and4_1;
  wire [0:0] u_csamul_cla32_ha4_1_xor0;
  wire [0:0] u_csamul_cla32_ha4_1_and0;
  wire [0:0] u_csamul_cla32_and5_1;
  wire [0:0] u_csamul_cla32_ha5_1_xor0;
  wire [0:0] u_csamul_cla32_ha5_1_and0;
  wire [0:0] u_csamul_cla32_and6_1;
  wire [0:0] u_csamul_cla32_ha6_1_xor0;
  wire [0:0] u_csamul_cla32_ha6_1_and0;
  wire [0:0] u_csamul_cla32_and7_1;
  wire [0:0] u_csamul_cla32_ha7_1_xor0;
  wire [0:0] u_csamul_cla32_ha7_1_and0;
  wire [0:0] u_csamul_cla32_and8_1;
  wire [0:0] u_csamul_cla32_ha8_1_xor0;
  wire [0:0] u_csamul_cla32_ha8_1_and0;
  wire [0:0] u_csamul_cla32_and9_1;
  wire [0:0] u_csamul_cla32_ha9_1_xor0;
  wire [0:0] u_csamul_cla32_ha9_1_and0;
  wire [0:0] u_csamul_cla32_and10_1;
  wire [0:0] u_csamul_cla32_ha10_1_xor0;
  wire [0:0] u_csamul_cla32_ha10_1_and0;
  wire [0:0] u_csamul_cla32_and11_1;
  wire [0:0] u_csamul_cla32_ha11_1_xor0;
  wire [0:0] u_csamul_cla32_ha11_1_and0;
  wire [0:0] u_csamul_cla32_and12_1;
  wire [0:0] u_csamul_cla32_ha12_1_xor0;
  wire [0:0] u_csamul_cla32_ha12_1_and0;
  wire [0:0] u_csamul_cla32_and13_1;
  wire [0:0] u_csamul_cla32_ha13_1_xor0;
  wire [0:0] u_csamul_cla32_ha13_1_and0;
  wire [0:0] u_csamul_cla32_and14_1;
  wire [0:0] u_csamul_cla32_ha14_1_xor0;
  wire [0:0] u_csamul_cla32_ha14_1_and0;
  wire [0:0] u_csamul_cla32_and15_1;
  wire [0:0] u_csamul_cla32_ha15_1_xor0;
  wire [0:0] u_csamul_cla32_ha15_1_and0;
  wire [0:0] u_csamul_cla32_and16_1;
  wire [0:0] u_csamul_cla32_ha16_1_xor0;
  wire [0:0] u_csamul_cla32_ha16_1_and0;
  wire [0:0] u_csamul_cla32_and17_1;
  wire [0:0] u_csamul_cla32_ha17_1_xor0;
  wire [0:0] u_csamul_cla32_ha17_1_and0;
  wire [0:0] u_csamul_cla32_and18_1;
  wire [0:0] u_csamul_cla32_ha18_1_xor0;
  wire [0:0] u_csamul_cla32_ha18_1_and0;
  wire [0:0] u_csamul_cla32_and19_1;
  wire [0:0] u_csamul_cla32_ha19_1_xor0;
  wire [0:0] u_csamul_cla32_ha19_1_and0;
  wire [0:0] u_csamul_cla32_and20_1;
  wire [0:0] u_csamul_cla32_ha20_1_xor0;
  wire [0:0] u_csamul_cla32_ha20_1_and0;
  wire [0:0] u_csamul_cla32_and21_1;
  wire [0:0] u_csamul_cla32_ha21_1_xor0;
  wire [0:0] u_csamul_cla32_ha21_1_and0;
  wire [0:0] u_csamul_cla32_and22_1;
  wire [0:0] u_csamul_cla32_ha22_1_xor0;
  wire [0:0] u_csamul_cla32_ha22_1_and0;
  wire [0:0] u_csamul_cla32_and23_1;
  wire [0:0] u_csamul_cla32_ha23_1_xor0;
  wire [0:0] u_csamul_cla32_ha23_1_and0;
  wire [0:0] u_csamul_cla32_and24_1;
  wire [0:0] u_csamul_cla32_ha24_1_xor0;
  wire [0:0] u_csamul_cla32_ha24_1_and0;
  wire [0:0] u_csamul_cla32_and25_1;
  wire [0:0] u_csamul_cla32_ha25_1_xor0;
  wire [0:0] u_csamul_cla32_ha25_1_and0;
  wire [0:0] u_csamul_cla32_and26_1;
  wire [0:0] u_csamul_cla32_ha26_1_xor0;
  wire [0:0] u_csamul_cla32_ha26_1_and0;
  wire [0:0] u_csamul_cla32_and27_1;
  wire [0:0] u_csamul_cla32_ha27_1_xor0;
  wire [0:0] u_csamul_cla32_ha27_1_and0;
  wire [0:0] u_csamul_cla32_and28_1;
  wire [0:0] u_csamul_cla32_ha28_1_xor0;
  wire [0:0] u_csamul_cla32_ha28_1_and0;
  wire [0:0] u_csamul_cla32_and29_1;
  wire [0:0] u_csamul_cla32_ha29_1_xor0;
  wire [0:0] u_csamul_cla32_ha29_1_and0;
  wire [0:0] u_csamul_cla32_and30_1;
  wire [0:0] u_csamul_cla32_ha30_1_xor0;
  wire [0:0] u_csamul_cla32_ha30_1_and0;
  wire [0:0] u_csamul_cla32_and31_1;
  wire [0:0] u_csamul_cla32_and0_2;
  wire [0:0] u_csamul_cla32_fa0_2_xor1;
  wire [0:0] u_csamul_cla32_fa0_2_or0;
  wire [0:0] u_csamul_cla32_and1_2;
  wire [0:0] u_csamul_cla32_fa1_2_xor1;
  wire [0:0] u_csamul_cla32_fa1_2_or0;
  wire [0:0] u_csamul_cla32_and2_2;
  wire [0:0] u_csamul_cla32_fa2_2_xor1;
  wire [0:0] u_csamul_cla32_fa2_2_or0;
  wire [0:0] u_csamul_cla32_and3_2;
  wire [0:0] u_csamul_cla32_fa3_2_xor1;
  wire [0:0] u_csamul_cla32_fa3_2_or0;
  wire [0:0] u_csamul_cla32_and4_2;
  wire [0:0] u_csamul_cla32_fa4_2_xor1;
  wire [0:0] u_csamul_cla32_fa4_2_or0;
  wire [0:0] u_csamul_cla32_and5_2;
  wire [0:0] u_csamul_cla32_fa5_2_xor1;
  wire [0:0] u_csamul_cla32_fa5_2_or0;
  wire [0:0] u_csamul_cla32_and6_2;
  wire [0:0] u_csamul_cla32_fa6_2_xor1;
  wire [0:0] u_csamul_cla32_fa6_2_or0;
  wire [0:0] u_csamul_cla32_and7_2;
  wire [0:0] u_csamul_cla32_fa7_2_xor1;
  wire [0:0] u_csamul_cla32_fa7_2_or0;
  wire [0:0] u_csamul_cla32_and8_2;
  wire [0:0] u_csamul_cla32_fa8_2_xor1;
  wire [0:0] u_csamul_cla32_fa8_2_or0;
  wire [0:0] u_csamul_cla32_and9_2;
  wire [0:0] u_csamul_cla32_fa9_2_xor1;
  wire [0:0] u_csamul_cla32_fa9_2_or0;
  wire [0:0] u_csamul_cla32_and10_2;
  wire [0:0] u_csamul_cla32_fa10_2_xor1;
  wire [0:0] u_csamul_cla32_fa10_2_or0;
  wire [0:0] u_csamul_cla32_and11_2;
  wire [0:0] u_csamul_cla32_fa11_2_xor1;
  wire [0:0] u_csamul_cla32_fa11_2_or0;
  wire [0:0] u_csamul_cla32_and12_2;
  wire [0:0] u_csamul_cla32_fa12_2_xor1;
  wire [0:0] u_csamul_cla32_fa12_2_or0;
  wire [0:0] u_csamul_cla32_and13_2;
  wire [0:0] u_csamul_cla32_fa13_2_xor1;
  wire [0:0] u_csamul_cla32_fa13_2_or0;
  wire [0:0] u_csamul_cla32_and14_2;
  wire [0:0] u_csamul_cla32_fa14_2_xor1;
  wire [0:0] u_csamul_cla32_fa14_2_or0;
  wire [0:0] u_csamul_cla32_and15_2;
  wire [0:0] u_csamul_cla32_fa15_2_xor1;
  wire [0:0] u_csamul_cla32_fa15_2_or0;
  wire [0:0] u_csamul_cla32_and16_2;
  wire [0:0] u_csamul_cla32_fa16_2_xor1;
  wire [0:0] u_csamul_cla32_fa16_2_or0;
  wire [0:0] u_csamul_cla32_and17_2;
  wire [0:0] u_csamul_cla32_fa17_2_xor1;
  wire [0:0] u_csamul_cla32_fa17_2_or0;
  wire [0:0] u_csamul_cla32_and18_2;
  wire [0:0] u_csamul_cla32_fa18_2_xor1;
  wire [0:0] u_csamul_cla32_fa18_2_or0;
  wire [0:0] u_csamul_cla32_and19_2;
  wire [0:0] u_csamul_cla32_fa19_2_xor1;
  wire [0:0] u_csamul_cla32_fa19_2_or0;
  wire [0:0] u_csamul_cla32_and20_2;
  wire [0:0] u_csamul_cla32_fa20_2_xor1;
  wire [0:0] u_csamul_cla32_fa20_2_or0;
  wire [0:0] u_csamul_cla32_and21_2;
  wire [0:0] u_csamul_cla32_fa21_2_xor1;
  wire [0:0] u_csamul_cla32_fa21_2_or0;
  wire [0:0] u_csamul_cla32_and22_2;
  wire [0:0] u_csamul_cla32_fa22_2_xor1;
  wire [0:0] u_csamul_cla32_fa22_2_or0;
  wire [0:0] u_csamul_cla32_and23_2;
  wire [0:0] u_csamul_cla32_fa23_2_xor1;
  wire [0:0] u_csamul_cla32_fa23_2_or0;
  wire [0:0] u_csamul_cla32_and24_2;
  wire [0:0] u_csamul_cla32_fa24_2_xor1;
  wire [0:0] u_csamul_cla32_fa24_2_or0;
  wire [0:0] u_csamul_cla32_and25_2;
  wire [0:0] u_csamul_cla32_fa25_2_xor1;
  wire [0:0] u_csamul_cla32_fa25_2_or0;
  wire [0:0] u_csamul_cla32_and26_2;
  wire [0:0] u_csamul_cla32_fa26_2_xor1;
  wire [0:0] u_csamul_cla32_fa26_2_or0;
  wire [0:0] u_csamul_cla32_and27_2;
  wire [0:0] u_csamul_cla32_fa27_2_xor1;
  wire [0:0] u_csamul_cla32_fa27_2_or0;
  wire [0:0] u_csamul_cla32_and28_2;
  wire [0:0] u_csamul_cla32_fa28_2_xor1;
  wire [0:0] u_csamul_cla32_fa28_2_or0;
  wire [0:0] u_csamul_cla32_and29_2;
  wire [0:0] u_csamul_cla32_fa29_2_xor1;
  wire [0:0] u_csamul_cla32_fa29_2_or0;
  wire [0:0] u_csamul_cla32_and30_2;
  wire [0:0] u_csamul_cla32_fa30_2_xor1;
  wire [0:0] u_csamul_cla32_fa30_2_or0;
  wire [0:0] u_csamul_cla32_and31_2;
  wire [0:0] u_csamul_cla32_and0_3;
  wire [0:0] u_csamul_cla32_fa0_3_xor1;
  wire [0:0] u_csamul_cla32_fa0_3_or0;
  wire [0:0] u_csamul_cla32_and1_3;
  wire [0:0] u_csamul_cla32_fa1_3_xor1;
  wire [0:0] u_csamul_cla32_fa1_3_or0;
  wire [0:0] u_csamul_cla32_and2_3;
  wire [0:0] u_csamul_cla32_fa2_3_xor1;
  wire [0:0] u_csamul_cla32_fa2_3_or0;
  wire [0:0] u_csamul_cla32_and3_3;
  wire [0:0] u_csamul_cla32_fa3_3_xor1;
  wire [0:0] u_csamul_cla32_fa3_3_or0;
  wire [0:0] u_csamul_cla32_and4_3;
  wire [0:0] u_csamul_cla32_fa4_3_xor1;
  wire [0:0] u_csamul_cla32_fa4_3_or0;
  wire [0:0] u_csamul_cla32_and5_3;
  wire [0:0] u_csamul_cla32_fa5_3_xor1;
  wire [0:0] u_csamul_cla32_fa5_3_or0;
  wire [0:0] u_csamul_cla32_and6_3;
  wire [0:0] u_csamul_cla32_fa6_3_xor1;
  wire [0:0] u_csamul_cla32_fa6_3_or0;
  wire [0:0] u_csamul_cla32_and7_3;
  wire [0:0] u_csamul_cla32_fa7_3_xor1;
  wire [0:0] u_csamul_cla32_fa7_3_or0;
  wire [0:0] u_csamul_cla32_and8_3;
  wire [0:0] u_csamul_cla32_fa8_3_xor1;
  wire [0:0] u_csamul_cla32_fa8_3_or0;
  wire [0:0] u_csamul_cla32_and9_3;
  wire [0:0] u_csamul_cla32_fa9_3_xor1;
  wire [0:0] u_csamul_cla32_fa9_3_or0;
  wire [0:0] u_csamul_cla32_and10_3;
  wire [0:0] u_csamul_cla32_fa10_3_xor1;
  wire [0:0] u_csamul_cla32_fa10_3_or0;
  wire [0:0] u_csamul_cla32_and11_3;
  wire [0:0] u_csamul_cla32_fa11_3_xor1;
  wire [0:0] u_csamul_cla32_fa11_3_or0;
  wire [0:0] u_csamul_cla32_and12_3;
  wire [0:0] u_csamul_cla32_fa12_3_xor1;
  wire [0:0] u_csamul_cla32_fa12_3_or0;
  wire [0:0] u_csamul_cla32_and13_3;
  wire [0:0] u_csamul_cla32_fa13_3_xor1;
  wire [0:0] u_csamul_cla32_fa13_3_or0;
  wire [0:0] u_csamul_cla32_and14_3;
  wire [0:0] u_csamul_cla32_fa14_3_xor1;
  wire [0:0] u_csamul_cla32_fa14_3_or0;
  wire [0:0] u_csamul_cla32_and15_3;
  wire [0:0] u_csamul_cla32_fa15_3_xor1;
  wire [0:0] u_csamul_cla32_fa15_3_or0;
  wire [0:0] u_csamul_cla32_and16_3;
  wire [0:0] u_csamul_cla32_fa16_3_xor1;
  wire [0:0] u_csamul_cla32_fa16_3_or0;
  wire [0:0] u_csamul_cla32_and17_3;
  wire [0:0] u_csamul_cla32_fa17_3_xor1;
  wire [0:0] u_csamul_cla32_fa17_3_or0;
  wire [0:0] u_csamul_cla32_and18_3;
  wire [0:0] u_csamul_cla32_fa18_3_xor1;
  wire [0:0] u_csamul_cla32_fa18_3_or0;
  wire [0:0] u_csamul_cla32_and19_3;
  wire [0:0] u_csamul_cla32_fa19_3_xor1;
  wire [0:0] u_csamul_cla32_fa19_3_or0;
  wire [0:0] u_csamul_cla32_and20_3;
  wire [0:0] u_csamul_cla32_fa20_3_xor1;
  wire [0:0] u_csamul_cla32_fa20_3_or0;
  wire [0:0] u_csamul_cla32_and21_3;
  wire [0:0] u_csamul_cla32_fa21_3_xor1;
  wire [0:0] u_csamul_cla32_fa21_3_or0;
  wire [0:0] u_csamul_cla32_and22_3;
  wire [0:0] u_csamul_cla32_fa22_3_xor1;
  wire [0:0] u_csamul_cla32_fa22_3_or0;
  wire [0:0] u_csamul_cla32_and23_3;
  wire [0:0] u_csamul_cla32_fa23_3_xor1;
  wire [0:0] u_csamul_cla32_fa23_3_or0;
  wire [0:0] u_csamul_cla32_and24_3;
  wire [0:0] u_csamul_cla32_fa24_3_xor1;
  wire [0:0] u_csamul_cla32_fa24_3_or0;
  wire [0:0] u_csamul_cla32_and25_3;
  wire [0:0] u_csamul_cla32_fa25_3_xor1;
  wire [0:0] u_csamul_cla32_fa25_3_or0;
  wire [0:0] u_csamul_cla32_and26_3;
  wire [0:0] u_csamul_cla32_fa26_3_xor1;
  wire [0:0] u_csamul_cla32_fa26_3_or0;
  wire [0:0] u_csamul_cla32_and27_3;
  wire [0:0] u_csamul_cla32_fa27_3_xor1;
  wire [0:0] u_csamul_cla32_fa27_3_or0;
  wire [0:0] u_csamul_cla32_and28_3;
  wire [0:0] u_csamul_cla32_fa28_3_xor1;
  wire [0:0] u_csamul_cla32_fa28_3_or0;
  wire [0:0] u_csamul_cla32_and29_3;
  wire [0:0] u_csamul_cla32_fa29_3_xor1;
  wire [0:0] u_csamul_cla32_fa29_3_or0;
  wire [0:0] u_csamul_cla32_and30_3;
  wire [0:0] u_csamul_cla32_fa30_3_xor1;
  wire [0:0] u_csamul_cla32_fa30_3_or0;
  wire [0:0] u_csamul_cla32_and31_3;
  wire [0:0] u_csamul_cla32_and0_4;
  wire [0:0] u_csamul_cla32_fa0_4_xor1;
  wire [0:0] u_csamul_cla32_fa0_4_or0;
  wire [0:0] u_csamul_cla32_and1_4;
  wire [0:0] u_csamul_cla32_fa1_4_xor1;
  wire [0:0] u_csamul_cla32_fa1_4_or0;
  wire [0:0] u_csamul_cla32_and2_4;
  wire [0:0] u_csamul_cla32_fa2_4_xor1;
  wire [0:0] u_csamul_cla32_fa2_4_or0;
  wire [0:0] u_csamul_cla32_and3_4;
  wire [0:0] u_csamul_cla32_fa3_4_xor1;
  wire [0:0] u_csamul_cla32_fa3_4_or0;
  wire [0:0] u_csamul_cla32_and4_4;
  wire [0:0] u_csamul_cla32_fa4_4_xor1;
  wire [0:0] u_csamul_cla32_fa4_4_or0;
  wire [0:0] u_csamul_cla32_and5_4;
  wire [0:0] u_csamul_cla32_fa5_4_xor1;
  wire [0:0] u_csamul_cla32_fa5_4_or0;
  wire [0:0] u_csamul_cla32_and6_4;
  wire [0:0] u_csamul_cla32_fa6_4_xor1;
  wire [0:0] u_csamul_cla32_fa6_4_or0;
  wire [0:0] u_csamul_cla32_and7_4;
  wire [0:0] u_csamul_cla32_fa7_4_xor1;
  wire [0:0] u_csamul_cla32_fa7_4_or0;
  wire [0:0] u_csamul_cla32_and8_4;
  wire [0:0] u_csamul_cla32_fa8_4_xor1;
  wire [0:0] u_csamul_cla32_fa8_4_or0;
  wire [0:0] u_csamul_cla32_and9_4;
  wire [0:0] u_csamul_cla32_fa9_4_xor1;
  wire [0:0] u_csamul_cla32_fa9_4_or0;
  wire [0:0] u_csamul_cla32_and10_4;
  wire [0:0] u_csamul_cla32_fa10_4_xor1;
  wire [0:0] u_csamul_cla32_fa10_4_or0;
  wire [0:0] u_csamul_cla32_and11_4;
  wire [0:0] u_csamul_cla32_fa11_4_xor1;
  wire [0:0] u_csamul_cla32_fa11_4_or0;
  wire [0:0] u_csamul_cla32_and12_4;
  wire [0:0] u_csamul_cla32_fa12_4_xor1;
  wire [0:0] u_csamul_cla32_fa12_4_or0;
  wire [0:0] u_csamul_cla32_and13_4;
  wire [0:0] u_csamul_cla32_fa13_4_xor1;
  wire [0:0] u_csamul_cla32_fa13_4_or0;
  wire [0:0] u_csamul_cla32_and14_4;
  wire [0:0] u_csamul_cla32_fa14_4_xor1;
  wire [0:0] u_csamul_cla32_fa14_4_or0;
  wire [0:0] u_csamul_cla32_and15_4;
  wire [0:0] u_csamul_cla32_fa15_4_xor1;
  wire [0:0] u_csamul_cla32_fa15_4_or0;
  wire [0:0] u_csamul_cla32_and16_4;
  wire [0:0] u_csamul_cla32_fa16_4_xor1;
  wire [0:0] u_csamul_cla32_fa16_4_or0;
  wire [0:0] u_csamul_cla32_and17_4;
  wire [0:0] u_csamul_cla32_fa17_4_xor1;
  wire [0:0] u_csamul_cla32_fa17_4_or0;
  wire [0:0] u_csamul_cla32_and18_4;
  wire [0:0] u_csamul_cla32_fa18_4_xor1;
  wire [0:0] u_csamul_cla32_fa18_4_or0;
  wire [0:0] u_csamul_cla32_and19_4;
  wire [0:0] u_csamul_cla32_fa19_4_xor1;
  wire [0:0] u_csamul_cla32_fa19_4_or0;
  wire [0:0] u_csamul_cla32_and20_4;
  wire [0:0] u_csamul_cla32_fa20_4_xor1;
  wire [0:0] u_csamul_cla32_fa20_4_or0;
  wire [0:0] u_csamul_cla32_and21_4;
  wire [0:0] u_csamul_cla32_fa21_4_xor1;
  wire [0:0] u_csamul_cla32_fa21_4_or0;
  wire [0:0] u_csamul_cla32_and22_4;
  wire [0:0] u_csamul_cla32_fa22_4_xor1;
  wire [0:0] u_csamul_cla32_fa22_4_or0;
  wire [0:0] u_csamul_cla32_and23_4;
  wire [0:0] u_csamul_cla32_fa23_4_xor1;
  wire [0:0] u_csamul_cla32_fa23_4_or0;
  wire [0:0] u_csamul_cla32_and24_4;
  wire [0:0] u_csamul_cla32_fa24_4_xor1;
  wire [0:0] u_csamul_cla32_fa24_4_or0;
  wire [0:0] u_csamul_cla32_and25_4;
  wire [0:0] u_csamul_cla32_fa25_4_xor1;
  wire [0:0] u_csamul_cla32_fa25_4_or0;
  wire [0:0] u_csamul_cla32_and26_4;
  wire [0:0] u_csamul_cla32_fa26_4_xor1;
  wire [0:0] u_csamul_cla32_fa26_4_or0;
  wire [0:0] u_csamul_cla32_and27_4;
  wire [0:0] u_csamul_cla32_fa27_4_xor1;
  wire [0:0] u_csamul_cla32_fa27_4_or0;
  wire [0:0] u_csamul_cla32_and28_4;
  wire [0:0] u_csamul_cla32_fa28_4_xor1;
  wire [0:0] u_csamul_cla32_fa28_4_or0;
  wire [0:0] u_csamul_cla32_and29_4;
  wire [0:0] u_csamul_cla32_fa29_4_xor1;
  wire [0:0] u_csamul_cla32_fa29_4_or0;
  wire [0:0] u_csamul_cla32_and30_4;
  wire [0:0] u_csamul_cla32_fa30_4_xor1;
  wire [0:0] u_csamul_cla32_fa30_4_or0;
  wire [0:0] u_csamul_cla32_and31_4;
  wire [0:0] u_csamul_cla32_and0_5;
  wire [0:0] u_csamul_cla32_fa0_5_xor1;
  wire [0:0] u_csamul_cla32_fa0_5_or0;
  wire [0:0] u_csamul_cla32_and1_5;
  wire [0:0] u_csamul_cla32_fa1_5_xor1;
  wire [0:0] u_csamul_cla32_fa1_5_or0;
  wire [0:0] u_csamul_cla32_and2_5;
  wire [0:0] u_csamul_cla32_fa2_5_xor1;
  wire [0:0] u_csamul_cla32_fa2_5_or0;
  wire [0:0] u_csamul_cla32_and3_5;
  wire [0:0] u_csamul_cla32_fa3_5_xor1;
  wire [0:0] u_csamul_cla32_fa3_5_or0;
  wire [0:0] u_csamul_cla32_and4_5;
  wire [0:0] u_csamul_cla32_fa4_5_xor1;
  wire [0:0] u_csamul_cla32_fa4_5_or0;
  wire [0:0] u_csamul_cla32_and5_5;
  wire [0:0] u_csamul_cla32_fa5_5_xor1;
  wire [0:0] u_csamul_cla32_fa5_5_or0;
  wire [0:0] u_csamul_cla32_and6_5;
  wire [0:0] u_csamul_cla32_fa6_5_xor1;
  wire [0:0] u_csamul_cla32_fa6_5_or0;
  wire [0:0] u_csamul_cla32_and7_5;
  wire [0:0] u_csamul_cla32_fa7_5_xor1;
  wire [0:0] u_csamul_cla32_fa7_5_or0;
  wire [0:0] u_csamul_cla32_and8_5;
  wire [0:0] u_csamul_cla32_fa8_5_xor1;
  wire [0:0] u_csamul_cla32_fa8_5_or0;
  wire [0:0] u_csamul_cla32_and9_5;
  wire [0:0] u_csamul_cla32_fa9_5_xor1;
  wire [0:0] u_csamul_cla32_fa9_5_or0;
  wire [0:0] u_csamul_cla32_and10_5;
  wire [0:0] u_csamul_cla32_fa10_5_xor1;
  wire [0:0] u_csamul_cla32_fa10_5_or0;
  wire [0:0] u_csamul_cla32_and11_5;
  wire [0:0] u_csamul_cla32_fa11_5_xor1;
  wire [0:0] u_csamul_cla32_fa11_5_or0;
  wire [0:0] u_csamul_cla32_and12_5;
  wire [0:0] u_csamul_cla32_fa12_5_xor1;
  wire [0:0] u_csamul_cla32_fa12_5_or0;
  wire [0:0] u_csamul_cla32_and13_5;
  wire [0:0] u_csamul_cla32_fa13_5_xor1;
  wire [0:0] u_csamul_cla32_fa13_5_or0;
  wire [0:0] u_csamul_cla32_and14_5;
  wire [0:0] u_csamul_cla32_fa14_5_xor1;
  wire [0:0] u_csamul_cla32_fa14_5_or0;
  wire [0:0] u_csamul_cla32_and15_5;
  wire [0:0] u_csamul_cla32_fa15_5_xor1;
  wire [0:0] u_csamul_cla32_fa15_5_or0;
  wire [0:0] u_csamul_cla32_and16_5;
  wire [0:0] u_csamul_cla32_fa16_5_xor1;
  wire [0:0] u_csamul_cla32_fa16_5_or0;
  wire [0:0] u_csamul_cla32_and17_5;
  wire [0:0] u_csamul_cla32_fa17_5_xor1;
  wire [0:0] u_csamul_cla32_fa17_5_or0;
  wire [0:0] u_csamul_cla32_and18_5;
  wire [0:0] u_csamul_cla32_fa18_5_xor1;
  wire [0:0] u_csamul_cla32_fa18_5_or0;
  wire [0:0] u_csamul_cla32_and19_5;
  wire [0:0] u_csamul_cla32_fa19_5_xor1;
  wire [0:0] u_csamul_cla32_fa19_5_or0;
  wire [0:0] u_csamul_cla32_and20_5;
  wire [0:0] u_csamul_cla32_fa20_5_xor1;
  wire [0:0] u_csamul_cla32_fa20_5_or0;
  wire [0:0] u_csamul_cla32_and21_5;
  wire [0:0] u_csamul_cla32_fa21_5_xor1;
  wire [0:0] u_csamul_cla32_fa21_5_or0;
  wire [0:0] u_csamul_cla32_and22_5;
  wire [0:0] u_csamul_cla32_fa22_5_xor1;
  wire [0:0] u_csamul_cla32_fa22_5_or0;
  wire [0:0] u_csamul_cla32_and23_5;
  wire [0:0] u_csamul_cla32_fa23_5_xor1;
  wire [0:0] u_csamul_cla32_fa23_5_or0;
  wire [0:0] u_csamul_cla32_and24_5;
  wire [0:0] u_csamul_cla32_fa24_5_xor1;
  wire [0:0] u_csamul_cla32_fa24_5_or0;
  wire [0:0] u_csamul_cla32_and25_5;
  wire [0:0] u_csamul_cla32_fa25_5_xor1;
  wire [0:0] u_csamul_cla32_fa25_5_or0;
  wire [0:0] u_csamul_cla32_and26_5;
  wire [0:0] u_csamul_cla32_fa26_5_xor1;
  wire [0:0] u_csamul_cla32_fa26_5_or0;
  wire [0:0] u_csamul_cla32_and27_5;
  wire [0:0] u_csamul_cla32_fa27_5_xor1;
  wire [0:0] u_csamul_cla32_fa27_5_or0;
  wire [0:0] u_csamul_cla32_and28_5;
  wire [0:0] u_csamul_cla32_fa28_5_xor1;
  wire [0:0] u_csamul_cla32_fa28_5_or0;
  wire [0:0] u_csamul_cla32_and29_5;
  wire [0:0] u_csamul_cla32_fa29_5_xor1;
  wire [0:0] u_csamul_cla32_fa29_5_or0;
  wire [0:0] u_csamul_cla32_and30_5;
  wire [0:0] u_csamul_cla32_fa30_5_xor1;
  wire [0:0] u_csamul_cla32_fa30_5_or0;
  wire [0:0] u_csamul_cla32_and31_5;
  wire [0:0] u_csamul_cla32_and0_6;
  wire [0:0] u_csamul_cla32_fa0_6_xor1;
  wire [0:0] u_csamul_cla32_fa0_6_or0;
  wire [0:0] u_csamul_cla32_and1_6;
  wire [0:0] u_csamul_cla32_fa1_6_xor1;
  wire [0:0] u_csamul_cla32_fa1_6_or0;
  wire [0:0] u_csamul_cla32_and2_6;
  wire [0:0] u_csamul_cla32_fa2_6_xor1;
  wire [0:0] u_csamul_cla32_fa2_6_or0;
  wire [0:0] u_csamul_cla32_and3_6;
  wire [0:0] u_csamul_cla32_fa3_6_xor1;
  wire [0:0] u_csamul_cla32_fa3_6_or0;
  wire [0:0] u_csamul_cla32_and4_6;
  wire [0:0] u_csamul_cla32_fa4_6_xor1;
  wire [0:0] u_csamul_cla32_fa4_6_or0;
  wire [0:0] u_csamul_cla32_and5_6;
  wire [0:0] u_csamul_cla32_fa5_6_xor1;
  wire [0:0] u_csamul_cla32_fa5_6_or0;
  wire [0:0] u_csamul_cla32_and6_6;
  wire [0:0] u_csamul_cla32_fa6_6_xor1;
  wire [0:0] u_csamul_cla32_fa6_6_or0;
  wire [0:0] u_csamul_cla32_and7_6;
  wire [0:0] u_csamul_cla32_fa7_6_xor1;
  wire [0:0] u_csamul_cla32_fa7_6_or0;
  wire [0:0] u_csamul_cla32_and8_6;
  wire [0:0] u_csamul_cla32_fa8_6_xor1;
  wire [0:0] u_csamul_cla32_fa8_6_or0;
  wire [0:0] u_csamul_cla32_and9_6;
  wire [0:0] u_csamul_cla32_fa9_6_xor1;
  wire [0:0] u_csamul_cla32_fa9_6_or0;
  wire [0:0] u_csamul_cla32_and10_6;
  wire [0:0] u_csamul_cla32_fa10_6_xor1;
  wire [0:0] u_csamul_cla32_fa10_6_or0;
  wire [0:0] u_csamul_cla32_and11_6;
  wire [0:0] u_csamul_cla32_fa11_6_xor1;
  wire [0:0] u_csamul_cla32_fa11_6_or0;
  wire [0:0] u_csamul_cla32_and12_6;
  wire [0:0] u_csamul_cla32_fa12_6_xor1;
  wire [0:0] u_csamul_cla32_fa12_6_or0;
  wire [0:0] u_csamul_cla32_and13_6;
  wire [0:0] u_csamul_cla32_fa13_6_xor1;
  wire [0:0] u_csamul_cla32_fa13_6_or0;
  wire [0:0] u_csamul_cla32_and14_6;
  wire [0:0] u_csamul_cla32_fa14_6_xor1;
  wire [0:0] u_csamul_cla32_fa14_6_or0;
  wire [0:0] u_csamul_cla32_and15_6;
  wire [0:0] u_csamul_cla32_fa15_6_xor1;
  wire [0:0] u_csamul_cla32_fa15_6_or0;
  wire [0:0] u_csamul_cla32_and16_6;
  wire [0:0] u_csamul_cla32_fa16_6_xor1;
  wire [0:0] u_csamul_cla32_fa16_6_or0;
  wire [0:0] u_csamul_cla32_and17_6;
  wire [0:0] u_csamul_cla32_fa17_6_xor1;
  wire [0:0] u_csamul_cla32_fa17_6_or0;
  wire [0:0] u_csamul_cla32_and18_6;
  wire [0:0] u_csamul_cla32_fa18_6_xor1;
  wire [0:0] u_csamul_cla32_fa18_6_or0;
  wire [0:0] u_csamul_cla32_and19_6;
  wire [0:0] u_csamul_cla32_fa19_6_xor1;
  wire [0:0] u_csamul_cla32_fa19_6_or0;
  wire [0:0] u_csamul_cla32_and20_6;
  wire [0:0] u_csamul_cla32_fa20_6_xor1;
  wire [0:0] u_csamul_cla32_fa20_6_or0;
  wire [0:0] u_csamul_cla32_and21_6;
  wire [0:0] u_csamul_cla32_fa21_6_xor1;
  wire [0:0] u_csamul_cla32_fa21_6_or0;
  wire [0:0] u_csamul_cla32_and22_6;
  wire [0:0] u_csamul_cla32_fa22_6_xor1;
  wire [0:0] u_csamul_cla32_fa22_6_or0;
  wire [0:0] u_csamul_cla32_and23_6;
  wire [0:0] u_csamul_cla32_fa23_6_xor1;
  wire [0:0] u_csamul_cla32_fa23_6_or0;
  wire [0:0] u_csamul_cla32_and24_6;
  wire [0:0] u_csamul_cla32_fa24_6_xor1;
  wire [0:0] u_csamul_cla32_fa24_6_or0;
  wire [0:0] u_csamul_cla32_and25_6;
  wire [0:0] u_csamul_cla32_fa25_6_xor1;
  wire [0:0] u_csamul_cla32_fa25_6_or0;
  wire [0:0] u_csamul_cla32_and26_6;
  wire [0:0] u_csamul_cla32_fa26_6_xor1;
  wire [0:0] u_csamul_cla32_fa26_6_or0;
  wire [0:0] u_csamul_cla32_and27_6;
  wire [0:0] u_csamul_cla32_fa27_6_xor1;
  wire [0:0] u_csamul_cla32_fa27_6_or0;
  wire [0:0] u_csamul_cla32_and28_6;
  wire [0:0] u_csamul_cla32_fa28_6_xor1;
  wire [0:0] u_csamul_cla32_fa28_6_or0;
  wire [0:0] u_csamul_cla32_and29_6;
  wire [0:0] u_csamul_cla32_fa29_6_xor1;
  wire [0:0] u_csamul_cla32_fa29_6_or0;
  wire [0:0] u_csamul_cla32_and30_6;
  wire [0:0] u_csamul_cla32_fa30_6_xor1;
  wire [0:0] u_csamul_cla32_fa30_6_or0;
  wire [0:0] u_csamul_cla32_and31_6;
  wire [0:0] u_csamul_cla32_and0_7;
  wire [0:0] u_csamul_cla32_fa0_7_xor1;
  wire [0:0] u_csamul_cla32_fa0_7_or0;
  wire [0:0] u_csamul_cla32_and1_7;
  wire [0:0] u_csamul_cla32_fa1_7_xor1;
  wire [0:0] u_csamul_cla32_fa1_7_or0;
  wire [0:0] u_csamul_cla32_and2_7;
  wire [0:0] u_csamul_cla32_fa2_7_xor1;
  wire [0:0] u_csamul_cla32_fa2_7_or0;
  wire [0:0] u_csamul_cla32_and3_7;
  wire [0:0] u_csamul_cla32_fa3_7_xor1;
  wire [0:0] u_csamul_cla32_fa3_7_or0;
  wire [0:0] u_csamul_cla32_and4_7;
  wire [0:0] u_csamul_cla32_fa4_7_xor1;
  wire [0:0] u_csamul_cla32_fa4_7_or0;
  wire [0:0] u_csamul_cla32_and5_7;
  wire [0:0] u_csamul_cla32_fa5_7_xor1;
  wire [0:0] u_csamul_cla32_fa5_7_or0;
  wire [0:0] u_csamul_cla32_and6_7;
  wire [0:0] u_csamul_cla32_fa6_7_xor1;
  wire [0:0] u_csamul_cla32_fa6_7_or0;
  wire [0:0] u_csamul_cla32_and7_7;
  wire [0:0] u_csamul_cla32_fa7_7_xor1;
  wire [0:0] u_csamul_cla32_fa7_7_or0;
  wire [0:0] u_csamul_cla32_and8_7;
  wire [0:0] u_csamul_cla32_fa8_7_xor1;
  wire [0:0] u_csamul_cla32_fa8_7_or0;
  wire [0:0] u_csamul_cla32_and9_7;
  wire [0:0] u_csamul_cla32_fa9_7_xor1;
  wire [0:0] u_csamul_cla32_fa9_7_or0;
  wire [0:0] u_csamul_cla32_and10_7;
  wire [0:0] u_csamul_cla32_fa10_7_xor1;
  wire [0:0] u_csamul_cla32_fa10_7_or0;
  wire [0:0] u_csamul_cla32_and11_7;
  wire [0:0] u_csamul_cla32_fa11_7_xor1;
  wire [0:0] u_csamul_cla32_fa11_7_or0;
  wire [0:0] u_csamul_cla32_and12_7;
  wire [0:0] u_csamul_cla32_fa12_7_xor1;
  wire [0:0] u_csamul_cla32_fa12_7_or0;
  wire [0:0] u_csamul_cla32_and13_7;
  wire [0:0] u_csamul_cla32_fa13_7_xor1;
  wire [0:0] u_csamul_cla32_fa13_7_or0;
  wire [0:0] u_csamul_cla32_and14_7;
  wire [0:0] u_csamul_cla32_fa14_7_xor1;
  wire [0:0] u_csamul_cla32_fa14_7_or0;
  wire [0:0] u_csamul_cla32_and15_7;
  wire [0:0] u_csamul_cla32_fa15_7_xor1;
  wire [0:0] u_csamul_cla32_fa15_7_or0;
  wire [0:0] u_csamul_cla32_and16_7;
  wire [0:0] u_csamul_cla32_fa16_7_xor1;
  wire [0:0] u_csamul_cla32_fa16_7_or0;
  wire [0:0] u_csamul_cla32_and17_7;
  wire [0:0] u_csamul_cla32_fa17_7_xor1;
  wire [0:0] u_csamul_cla32_fa17_7_or0;
  wire [0:0] u_csamul_cla32_and18_7;
  wire [0:0] u_csamul_cla32_fa18_7_xor1;
  wire [0:0] u_csamul_cla32_fa18_7_or0;
  wire [0:0] u_csamul_cla32_and19_7;
  wire [0:0] u_csamul_cla32_fa19_7_xor1;
  wire [0:0] u_csamul_cla32_fa19_7_or0;
  wire [0:0] u_csamul_cla32_and20_7;
  wire [0:0] u_csamul_cla32_fa20_7_xor1;
  wire [0:0] u_csamul_cla32_fa20_7_or0;
  wire [0:0] u_csamul_cla32_and21_7;
  wire [0:0] u_csamul_cla32_fa21_7_xor1;
  wire [0:0] u_csamul_cla32_fa21_7_or0;
  wire [0:0] u_csamul_cla32_and22_7;
  wire [0:0] u_csamul_cla32_fa22_7_xor1;
  wire [0:0] u_csamul_cla32_fa22_7_or0;
  wire [0:0] u_csamul_cla32_and23_7;
  wire [0:0] u_csamul_cla32_fa23_7_xor1;
  wire [0:0] u_csamul_cla32_fa23_7_or0;
  wire [0:0] u_csamul_cla32_and24_7;
  wire [0:0] u_csamul_cla32_fa24_7_xor1;
  wire [0:0] u_csamul_cla32_fa24_7_or0;
  wire [0:0] u_csamul_cla32_and25_7;
  wire [0:0] u_csamul_cla32_fa25_7_xor1;
  wire [0:0] u_csamul_cla32_fa25_7_or0;
  wire [0:0] u_csamul_cla32_and26_7;
  wire [0:0] u_csamul_cla32_fa26_7_xor1;
  wire [0:0] u_csamul_cla32_fa26_7_or0;
  wire [0:0] u_csamul_cla32_and27_7;
  wire [0:0] u_csamul_cla32_fa27_7_xor1;
  wire [0:0] u_csamul_cla32_fa27_7_or0;
  wire [0:0] u_csamul_cla32_and28_7;
  wire [0:0] u_csamul_cla32_fa28_7_xor1;
  wire [0:0] u_csamul_cla32_fa28_7_or0;
  wire [0:0] u_csamul_cla32_and29_7;
  wire [0:0] u_csamul_cla32_fa29_7_xor1;
  wire [0:0] u_csamul_cla32_fa29_7_or0;
  wire [0:0] u_csamul_cla32_and30_7;
  wire [0:0] u_csamul_cla32_fa30_7_xor1;
  wire [0:0] u_csamul_cla32_fa30_7_or0;
  wire [0:0] u_csamul_cla32_and31_7;
  wire [0:0] u_csamul_cla32_and0_8;
  wire [0:0] u_csamul_cla32_fa0_8_xor1;
  wire [0:0] u_csamul_cla32_fa0_8_or0;
  wire [0:0] u_csamul_cla32_and1_8;
  wire [0:0] u_csamul_cla32_fa1_8_xor1;
  wire [0:0] u_csamul_cla32_fa1_8_or0;
  wire [0:0] u_csamul_cla32_and2_8;
  wire [0:0] u_csamul_cla32_fa2_8_xor1;
  wire [0:0] u_csamul_cla32_fa2_8_or0;
  wire [0:0] u_csamul_cla32_and3_8;
  wire [0:0] u_csamul_cla32_fa3_8_xor1;
  wire [0:0] u_csamul_cla32_fa3_8_or0;
  wire [0:0] u_csamul_cla32_and4_8;
  wire [0:0] u_csamul_cla32_fa4_8_xor1;
  wire [0:0] u_csamul_cla32_fa4_8_or0;
  wire [0:0] u_csamul_cla32_and5_8;
  wire [0:0] u_csamul_cla32_fa5_8_xor1;
  wire [0:0] u_csamul_cla32_fa5_8_or0;
  wire [0:0] u_csamul_cla32_and6_8;
  wire [0:0] u_csamul_cla32_fa6_8_xor1;
  wire [0:0] u_csamul_cla32_fa6_8_or0;
  wire [0:0] u_csamul_cla32_and7_8;
  wire [0:0] u_csamul_cla32_fa7_8_xor1;
  wire [0:0] u_csamul_cla32_fa7_8_or0;
  wire [0:0] u_csamul_cla32_and8_8;
  wire [0:0] u_csamul_cla32_fa8_8_xor1;
  wire [0:0] u_csamul_cla32_fa8_8_or0;
  wire [0:0] u_csamul_cla32_and9_8;
  wire [0:0] u_csamul_cla32_fa9_8_xor1;
  wire [0:0] u_csamul_cla32_fa9_8_or0;
  wire [0:0] u_csamul_cla32_and10_8;
  wire [0:0] u_csamul_cla32_fa10_8_xor1;
  wire [0:0] u_csamul_cla32_fa10_8_or0;
  wire [0:0] u_csamul_cla32_and11_8;
  wire [0:0] u_csamul_cla32_fa11_8_xor1;
  wire [0:0] u_csamul_cla32_fa11_8_or0;
  wire [0:0] u_csamul_cla32_and12_8;
  wire [0:0] u_csamul_cla32_fa12_8_xor1;
  wire [0:0] u_csamul_cla32_fa12_8_or0;
  wire [0:0] u_csamul_cla32_and13_8;
  wire [0:0] u_csamul_cla32_fa13_8_xor1;
  wire [0:0] u_csamul_cla32_fa13_8_or0;
  wire [0:0] u_csamul_cla32_and14_8;
  wire [0:0] u_csamul_cla32_fa14_8_xor1;
  wire [0:0] u_csamul_cla32_fa14_8_or0;
  wire [0:0] u_csamul_cla32_and15_8;
  wire [0:0] u_csamul_cla32_fa15_8_xor1;
  wire [0:0] u_csamul_cla32_fa15_8_or0;
  wire [0:0] u_csamul_cla32_and16_8;
  wire [0:0] u_csamul_cla32_fa16_8_xor1;
  wire [0:0] u_csamul_cla32_fa16_8_or0;
  wire [0:0] u_csamul_cla32_and17_8;
  wire [0:0] u_csamul_cla32_fa17_8_xor1;
  wire [0:0] u_csamul_cla32_fa17_8_or0;
  wire [0:0] u_csamul_cla32_and18_8;
  wire [0:0] u_csamul_cla32_fa18_8_xor1;
  wire [0:0] u_csamul_cla32_fa18_8_or0;
  wire [0:0] u_csamul_cla32_and19_8;
  wire [0:0] u_csamul_cla32_fa19_8_xor1;
  wire [0:0] u_csamul_cla32_fa19_8_or0;
  wire [0:0] u_csamul_cla32_and20_8;
  wire [0:0] u_csamul_cla32_fa20_8_xor1;
  wire [0:0] u_csamul_cla32_fa20_8_or0;
  wire [0:0] u_csamul_cla32_and21_8;
  wire [0:0] u_csamul_cla32_fa21_8_xor1;
  wire [0:0] u_csamul_cla32_fa21_8_or0;
  wire [0:0] u_csamul_cla32_and22_8;
  wire [0:0] u_csamul_cla32_fa22_8_xor1;
  wire [0:0] u_csamul_cla32_fa22_8_or0;
  wire [0:0] u_csamul_cla32_and23_8;
  wire [0:0] u_csamul_cla32_fa23_8_xor1;
  wire [0:0] u_csamul_cla32_fa23_8_or0;
  wire [0:0] u_csamul_cla32_and24_8;
  wire [0:0] u_csamul_cla32_fa24_8_xor1;
  wire [0:0] u_csamul_cla32_fa24_8_or0;
  wire [0:0] u_csamul_cla32_and25_8;
  wire [0:0] u_csamul_cla32_fa25_8_xor1;
  wire [0:0] u_csamul_cla32_fa25_8_or0;
  wire [0:0] u_csamul_cla32_and26_8;
  wire [0:0] u_csamul_cla32_fa26_8_xor1;
  wire [0:0] u_csamul_cla32_fa26_8_or0;
  wire [0:0] u_csamul_cla32_and27_8;
  wire [0:0] u_csamul_cla32_fa27_8_xor1;
  wire [0:0] u_csamul_cla32_fa27_8_or0;
  wire [0:0] u_csamul_cla32_and28_8;
  wire [0:0] u_csamul_cla32_fa28_8_xor1;
  wire [0:0] u_csamul_cla32_fa28_8_or0;
  wire [0:0] u_csamul_cla32_and29_8;
  wire [0:0] u_csamul_cla32_fa29_8_xor1;
  wire [0:0] u_csamul_cla32_fa29_8_or0;
  wire [0:0] u_csamul_cla32_and30_8;
  wire [0:0] u_csamul_cla32_fa30_8_xor1;
  wire [0:0] u_csamul_cla32_fa30_8_or0;
  wire [0:0] u_csamul_cla32_and31_8;
  wire [0:0] u_csamul_cla32_and0_9;
  wire [0:0] u_csamul_cla32_fa0_9_xor1;
  wire [0:0] u_csamul_cla32_fa0_9_or0;
  wire [0:0] u_csamul_cla32_and1_9;
  wire [0:0] u_csamul_cla32_fa1_9_xor1;
  wire [0:0] u_csamul_cla32_fa1_9_or0;
  wire [0:0] u_csamul_cla32_and2_9;
  wire [0:0] u_csamul_cla32_fa2_9_xor1;
  wire [0:0] u_csamul_cla32_fa2_9_or0;
  wire [0:0] u_csamul_cla32_and3_9;
  wire [0:0] u_csamul_cla32_fa3_9_xor1;
  wire [0:0] u_csamul_cla32_fa3_9_or0;
  wire [0:0] u_csamul_cla32_and4_9;
  wire [0:0] u_csamul_cla32_fa4_9_xor1;
  wire [0:0] u_csamul_cla32_fa4_9_or0;
  wire [0:0] u_csamul_cla32_and5_9;
  wire [0:0] u_csamul_cla32_fa5_9_xor1;
  wire [0:0] u_csamul_cla32_fa5_9_or0;
  wire [0:0] u_csamul_cla32_and6_9;
  wire [0:0] u_csamul_cla32_fa6_9_xor1;
  wire [0:0] u_csamul_cla32_fa6_9_or0;
  wire [0:0] u_csamul_cla32_and7_9;
  wire [0:0] u_csamul_cla32_fa7_9_xor1;
  wire [0:0] u_csamul_cla32_fa7_9_or0;
  wire [0:0] u_csamul_cla32_and8_9;
  wire [0:0] u_csamul_cla32_fa8_9_xor1;
  wire [0:0] u_csamul_cla32_fa8_9_or0;
  wire [0:0] u_csamul_cla32_and9_9;
  wire [0:0] u_csamul_cla32_fa9_9_xor1;
  wire [0:0] u_csamul_cla32_fa9_9_or0;
  wire [0:0] u_csamul_cla32_and10_9;
  wire [0:0] u_csamul_cla32_fa10_9_xor1;
  wire [0:0] u_csamul_cla32_fa10_9_or0;
  wire [0:0] u_csamul_cla32_and11_9;
  wire [0:0] u_csamul_cla32_fa11_9_xor1;
  wire [0:0] u_csamul_cla32_fa11_9_or0;
  wire [0:0] u_csamul_cla32_and12_9;
  wire [0:0] u_csamul_cla32_fa12_9_xor1;
  wire [0:0] u_csamul_cla32_fa12_9_or0;
  wire [0:0] u_csamul_cla32_and13_9;
  wire [0:0] u_csamul_cla32_fa13_9_xor1;
  wire [0:0] u_csamul_cla32_fa13_9_or0;
  wire [0:0] u_csamul_cla32_and14_9;
  wire [0:0] u_csamul_cla32_fa14_9_xor1;
  wire [0:0] u_csamul_cla32_fa14_9_or0;
  wire [0:0] u_csamul_cla32_and15_9;
  wire [0:0] u_csamul_cla32_fa15_9_xor1;
  wire [0:0] u_csamul_cla32_fa15_9_or0;
  wire [0:0] u_csamul_cla32_and16_9;
  wire [0:0] u_csamul_cla32_fa16_9_xor1;
  wire [0:0] u_csamul_cla32_fa16_9_or0;
  wire [0:0] u_csamul_cla32_and17_9;
  wire [0:0] u_csamul_cla32_fa17_9_xor1;
  wire [0:0] u_csamul_cla32_fa17_9_or0;
  wire [0:0] u_csamul_cla32_and18_9;
  wire [0:0] u_csamul_cla32_fa18_9_xor1;
  wire [0:0] u_csamul_cla32_fa18_9_or0;
  wire [0:0] u_csamul_cla32_and19_9;
  wire [0:0] u_csamul_cla32_fa19_9_xor1;
  wire [0:0] u_csamul_cla32_fa19_9_or0;
  wire [0:0] u_csamul_cla32_and20_9;
  wire [0:0] u_csamul_cla32_fa20_9_xor1;
  wire [0:0] u_csamul_cla32_fa20_9_or0;
  wire [0:0] u_csamul_cla32_and21_9;
  wire [0:0] u_csamul_cla32_fa21_9_xor1;
  wire [0:0] u_csamul_cla32_fa21_9_or0;
  wire [0:0] u_csamul_cla32_and22_9;
  wire [0:0] u_csamul_cla32_fa22_9_xor1;
  wire [0:0] u_csamul_cla32_fa22_9_or0;
  wire [0:0] u_csamul_cla32_and23_9;
  wire [0:0] u_csamul_cla32_fa23_9_xor1;
  wire [0:0] u_csamul_cla32_fa23_9_or0;
  wire [0:0] u_csamul_cla32_and24_9;
  wire [0:0] u_csamul_cla32_fa24_9_xor1;
  wire [0:0] u_csamul_cla32_fa24_9_or0;
  wire [0:0] u_csamul_cla32_and25_9;
  wire [0:0] u_csamul_cla32_fa25_9_xor1;
  wire [0:0] u_csamul_cla32_fa25_9_or0;
  wire [0:0] u_csamul_cla32_and26_9;
  wire [0:0] u_csamul_cla32_fa26_9_xor1;
  wire [0:0] u_csamul_cla32_fa26_9_or0;
  wire [0:0] u_csamul_cla32_and27_9;
  wire [0:0] u_csamul_cla32_fa27_9_xor1;
  wire [0:0] u_csamul_cla32_fa27_9_or0;
  wire [0:0] u_csamul_cla32_and28_9;
  wire [0:0] u_csamul_cla32_fa28_9_xor1;
  wire [0:0] u_csamul_cla32_fa28_9_or0;
  wire [0:0] u_csamul_cla32_and29_9;
  wire [0:0] u_csamul_cla32_fa29_9_xor1;
  wire [0:0] u_csamul_cla32_fa29_9_or0;
  wire [0:0] u_csamul_cla32_and30_9;
  wire [0:0] u_csamul_cla32_fa30_9_xor1;
  wire [0:0] u_csamul_cla32_fa30_9_or0;
  wire [0:0] u_csamul_cla32_and31_9;
  wire [0:0] u_csamul_cla32_and0_10;
  wire [0:0] u_csamul_cla32_fa0_10_xor1;
  wire [0:0] u_csamul_cla32_fa0_10_or0;
  wire [0:0] u_csamul_cla32_and1_10;
  wire [0:0] u_csamul_cla32_fa1_10_xor1;
  wire [0:0] u_csamul_cla32_fa1_10_or0;
  wire [0:0] u_csamul_cla32_and2_10;
  wire [0:0] u_csamul_cla32_fa2_10_xor1;
  wire [0:0] u_csamul_cla32_fa2_10_or0;
  wire [0:0] u_csamul_cla32_and3_10;
  wire [0:0] u_csamul_cla32_fa3_10_xor1;
  wire [0:0] u_csamul_cla32_fa3_10_or0;
  wire [0:0] u_csamul_cla32_and4_10;
  wire [0:0] u_csamul_cla32_fa4_10_xor1;
  wire [0:0] u_csamul_cla32_fa4_10_or0;
  wire [0:0] u_csamul_cla32_and5_10;
  wire [0:0] u_csamul_cla32_fa5_10_xor1;
  wire [0:0] u_csamul_cla32_fa5_10_or0;
  wire [0:0] u_csamul_cla32_and6_10;
  wire [0:0] u_csamul_cla32_fa6_10_xor1;
  wire [0:0] u_csamul_cla32_fa6_10_or0;
  wire [0:0] u_csamul_cla32_and7_10;
  wire [0:0] u_csamul_cla32_fa7_10_xor1;
  wire [0:0] u_csamul_cla32_fa7_10_or0;
  wire [0:0] u_csamul_cla32_and8_10;
  wire [0:0] u_csamul_cla32_fa8_10_xor1;
  wire [0:0] u_csamul_cla32_fa8_10_or0;
  wire [0:0] u_csamul_cla32_and9_10;
  wire [0:0] u_csamul_cla32_fa9_10_xor1;
  wire [0:0] u_csamul_cla32_fa9_10_or0;
  wire [0:0] u_csamul_cla32_and10_10;
  wire [0:0] u_csamul_cla32_fa10_10_xor1;
  wire [0:0] u_csamul_cla32_fa10_10_or0;
  wire [0:0] u_csamul_cla32_and11_10;
  wire [0:0] u_csamul_cla32_fa11_10_xor1;
  wire [0:0] u_csamul_cla32_fa11_10_or0;
  wire [0:0] u_csamul_cla32_and12_10;
  wire [0:0] u_csamul_cla32_fa12_10_xor1;
  wire [0:0] u_csamul_cla32_fa12_10_or0;
  wire [0:0] u_csamul_cla32_and13_10;
  wire [0:0] u_csamul_cla32_fa13_10_xor1;
  wire [0:0] u_csamul_cla32_fa13_10_or0;
  wire [0:0] u_csamul_cla32_and14_10;
  wire [0:0] u_csamul_cla32_fa14_10_xor1;
  wire [0:0] u_csamul_cla32_fa14_10_or0;
  wire [0:0] u_csamul_cla32_and15_10;
  wire [0:0] u_csamul_cla32_fa15_10_xor1;
  wire [0:0] u_csamul_cla32_fa15_10_or0;
  wire [0:0] u_csamul_cla32_and16_10;
  wire [0:0] u_csamul_cla32_fa16_10_xor1;
  wire [0:0] u_csamul_cla32_fa16_10_or0;
  wire [0:0] u_csamul_cla32_and17_10;
  wire [0:0] u_csamul_cla32_fa17_10_xor1;
  wire [0:0] u_csamul_cla32_fa17_10_or0;
  wire [0:0] u_csamul_cla32_and18_10;
  wire [0:0] u_csamul_cla32_fa18_10_xor1;
  wire [0:0] u_csamul_cla32_fa18_10_or0;
  wire [0:0] u_csamul_cla32_and19_10;
  wire [0:0] u_csamul_cla32_fa19_10_xor1;
  wire [0:0] u_csamul_cla32_fa19_10_or0;
  wire [0:0] u_csamul_cla32_and20_10;
  wire [0:0] u_csamul_cla32_fa20_10_xor1;
  wire [0:0] u_csamul_cla32_fa20_10_or0;
  wire [0:0] u_csamul_cla32_and21_10;
  wire [0:0] u_csamul_cla32_fa21_10_xor1;
  wire [0:0] u_csamul_cla32_fa21_10_or0;
  wire [0:0] u_csamul_cla32_and22_10;
  wire [0:0] u_csamul_cla32_fa22_10_xor1;
  wire [0:0] u_csamul_cla32_fa22_10_or0;
  wire [0:0] u_csamul_cla32_and23_10;
  wire [0:0] u_csamul_cla32_fa23_10_xor1;
  wire [0:0] u_csamul_cla32_fa23_10_or0;
  wire [0:0] u_csamul_cla32_and24_10;
  wire [0:0] u_csamul_cla32_fa24_10_xor1;
  wire [0:0] u_csamul_cla32_fa24_10_or0;
  wire [0:0] u_csamul_cla32_and25_10;
  wire [0:0] u_csamul_cla32_fa25_10_xor1;
  wire [0:0] u_csamul_cla32_fa25_10_or0;
  wire [0:0] u_csamul_cla32_and26_10;
  wire [0:0] u_csamul_cla32_fa26_10_xor1;
  wire [0:0] u_csamul_cla32_fa26_10_or0;
  wire [0:0] u_csamul_cla32_and27_10;
  wire [0:0] u_csamul_cla32_fa27_10_xor1;
  wire [0:0] u_csamul_cla32_fa27_10_or0;
  wire [0:0] u_csamul_cla32_and28_10;
  wire [0:0] u_csamul_cla32_fa28_10_xor1;
  wire [0:0] u_csamul_cla32_fa28_10_or0;
  wire [0:0] u_csamul_cla32_and29_10;
  wire [0:0] u_csamul_cla32_fa29_10_xor1;
  wire [0:0] u_csamul_cla32_fa29_10_or0;
  wire [0:0] u_csamul_cla32_and30_10;
  wire [0:0] u_csamul_cla32_fa30_10_xor1;
  wire [0:0] u_csamul_cla32_fa30_10_or0;
  wire [0:0] u_csamul_cla32_and31_10;
  wire [0:0] u_csamul_cla32_and0_11;
  wire [0:0] u_csamul_cla32_fa0_11_xor1;
  wire [0:0] u_csamul_cla32_fa0_11_or0;
  wire [0:0] u_csamul_cla32_and1_11;
  wire [0:0] u_csamul_cla32_fa1_11_xor1;
  wire [0:0] u_csamul_cla32_fa1_11_or0;
  wire [0:0] u_csamul_cla32_and2_11;
  wire [0:0] u_csamul_cla32_fa2_11_xor1;
  wire [0:0] u_csamul_cla32_fa2_11_or0;
  wire [0:0] u_csamul_cla32_and3_11;
  wire [0:0] u_csamul_cla32_fa3_11_xor1;
  wire [0:0] u_csamul_cla32_fa3_11_or0;
  wire [0:0] u_csamul_cla32_and4_11;
  wire [0:0] u_csamul_cla32_fa4_11_xor1;
  wire [0:0] u_csamul_cla32_fa4_11_or0;
  wire [0:0] u_csamul_cla32_and5_11;
  wire [0:0] u_csamul_cla32_fa5_11_xor1;
  wire [0:0] u_csamul_cla32_fa5_11_or0;
  wire [0:0] u_csamul_cla32_and6_11;
  wire [0:0] u_csamul_cla32_fa6_11_xor1;
  wire [0:0] u_csamul_cla32_fa6_11_or0;
  wire [0:0] u_csamul_cla32_and7_11;
  wire [0:0] u_csamul_cla32_fa7_11_xor1;
  wire [0:0] u_csamul_cla32_fa7_11_or0;
  wire [0:0] u_csamul_cla32_and8_11;
  wire [0:0] u_csamul_cla32_fa8_11_xor1;
  wire [0:0] u_csamul_cla32_fa8_11_or0;
  wire [0:0] u_csamul_cla32_and9_11;
  wire [0:0] u_csamul_cla32_fa9_11_xor1;
  wire [0:0] u_csamul_cla32_fa9_11_or0;
  wire [0:0] u_csamul_cla32_and10_11;
  wire [0:0] u_csamul_cla32_fa10_11_xor1;
  wire [0:0] u_csamul_cla32_fa10_11_or0;
  wire [0:0] u_csamul_cla32_and11_11;
  wire [0:0] u_csamul_cla32_fa11_11_xor1;
  wire [0:0] u_csamul_cla32_fa11_11_or0;
  wire [0:0] u_csamul_cla32_and12_11;
  wire [0:0] u_csamul_cla32_fa12_11_xor1;
  wire [0:0] u_csamul_cla32_fa12_11_or0;
  wire [0:0] u_csamul_cla32_and13_11;
  wire [0:0] u_csamul_cla32_fa13_11_xor1;
  wire [0:0] u_csamul_cla32_fa13_11_or0;
  wire [0:0] u_csamul_cla32_and14_11;
  wire [0:0] u_csamul_cla32_fa14_11_xor1;
  wire [0:0] u_csamul_cla32_fa14_11_or0;
  wire [0:0] u_csamul_cla32_and15_11;
  wire [0:0] u_csamul_cla32_fa15_11_xor1;
  wire [0:0] u_csamul_cla32_fa15_11_or0;
  wire [0:0] u_csamul_cla32_and16_11;
  wire [0:0] u_csamul_cla32_fa16_11_xor1;
  wire [0:0] u_csamul_cla32_fa16_11_or0;
  wire [0:0] u_csamul_cla32_and17_11;
  wire [0:0] u_csamul_cla32_fa17_11_xor1;
  wire [0:0] u_csamul_cla32_fa17_11_or0;
  wire [0:0] u_csamul_cla32_and18_11;
  wire [0:0] u_csamul_cla32_fa18_11_xor1;
  wire [0:0] u_csamul_cla32_fa18_11_or0;
  wire [0:0] u_csamul_cla32_and19_11;
  wire [0:0] u_csamul_cla32_fa19_11_xor1;
  wire [0:0] u_csamul_cla32_fa19_11_or0;
  wire [0:0] u_csamul_cla32_and20_11;
  wire [0:0] u_csamul_cla32_fa20_11_xor1;
  wire [0:0] u_csamul_cla32_fa20_11_or0;
  wire [0:0] u_csamul_cla32_and21_11;
  wire [0:0] u_csamul_cla32_fa21_11_xor1;
  wire [0:0] u_csamul_cla32_fa21_11_or0;
  wire [0:0] u_csamul_cla32_and22_11;
  wire [0:0] u_csamul_cla32_fa22_11_xor1;
  wire [0:0] u_csamul_cla32_fa22_11_or0;
  wire [0:0] u_csamul_cla32_and23_11;
  wire [0:0] u_csamul_cla32_fa23_11_xor1;
  wire [0:0] u_csamul_cla32_fa23_11_or0;
  wire [0:0] u_csamul_cla32_and24_11;
  wire [0:0] u_csamul_cla32_fa24_11_xor1;
  wire [0:0] u_csamul_cla32_fa24_11_or0;
  wire [0:0] u_csamul_cla32_and25_11;
  wire [0:0] u_csamul_cla32_fa25_11_xor1;
  wire [0:0] u_csamul_cla32_fa25_11_or0;
  wire [0:0] u_csamul_cla32_and26_11;
  wire [0:0] u_csamul_cla32_fa26_11_xor1;
  wire [0:0] u_csamul_cla32_fa26_11_or0;
  wire [0:0] u_csamul_cla32_and27_11;
  wire [0:0] u_csamul_cla32_fa27_11_xor1;
  wire [0:0] u_csamul_cla32_fa27_11_or0;
  wire [0:0] u_csamul_cla32_and28_11;
  wire [0:0] u_csamul_cla32_fa28_11_xor1;
  wire [0:0] u_csamul_cla32_fa28_11_or0;
  wire [0:0] u_csamul_cla32_and29_11;
  wire [0:0] u_csamul_cla32_fa29_11_xor1;
  wire [0:0] u_csamul_cla32_fa29_11_or0;
  wire [0:0] u_csamul_cla32_and30_11;
  wire [0:0] u_csamul_cla32_fa30_11_xor1;
  wire [0:0] u_csamul_cla32_fa30_11_or0;
  wire [0:0] u_csamul_cla32_and31_11;
  wire [0:0] u_csamul_cla32_and0_12;
  wire [0:0] u_csamul_cla32_fa0_12_xor1;
  wire [0:0] u_csamul_cla32_fa0_12_or0;
  wire [0:0] u_csamul_cla32_and1_12;
  wire [0:0] u_csamul_cla32_fa1_12_xor1;
  wire [0:0] u_csamul_cla32_fa1_12_or0;
  wire [0:0] u_csamul_cla32_and2_12;
  wire [0:0] u_csamul_cla32_fa2_12_xor1;
  wire [0:0] u_csamul_cla32_fa2_12_or0;
  wire [0:0] u_csamul_cla32_and3_12;
  wire [0:0] u_csamul_cla32_fa3_12_xor1;
  wire [0:0] u_csamul_cla32_fa3_12_or0;
  wire [0:0] u_csamul_cla32_and4_12;
  wire [0:0] u_csamul_cla32_fa4_12_xor1;
  wire [0:0] u_csamul_cla32_fa4_12_or0;
  wire [0:0] u_csamul_cla32_and5_12;
  wire [0:0] u_csamul_cla32_fa5_12_xor1;
  wire [0:0] u_csamul_cla32_fa5_12_or0;
  wire [0:0] u_csamul_cla32_and6_12;
  wire [0:0] u_csamul_cla32_fa6_12_xor1;
  wire [0:0] u_csamul_cla32_fa6_12_or0;
  wire [0:0] u_csamul_cla32_and7_12;
  wire [0:0] u_csamul_cla32_fa7_12_xor1;
  wire [0:0] u_csamul_cla32_fa7_12_or0;
  wire [0:0] u_csamul_cla32_and8_12;
  wire [0:0] u_csamul_cla32_fa8_12_xor1;
  wire [0:0] u_csamul_cla32_fa8_12_or0;
  wire [0:0] u_csamul_cla32_and9_12;
  wire [0:0] u_csamul_cla32_fa9_12_xor1;
  wire [0:0] u_csamul_cla32_fa9_12_or0;
  wire [0:0] u_csamul_cla32_and10_12;
  wire [0:0] u_csamul_cla32_fa10_12_xor1;
  wire [0:0] u_csamul_cla32_fa10_12_or0;
  wire [0:0] u_csamul_cla32_and11_12;
  wire [0:0] u_csamul_cla32_fa11_12_xor1;
  wire [0:0] u_csamul_cla32_fa11_12_or0;
  wire [0:0] u_csamul_cla32_and12_12;
  wire [0:0] u_csamul_cla32_fa12_12_xor1;
  wire [0:0] u_csamul_cla32_fa12_12_or0;
  wire [0:0] u_csamul_cla32_and13_12;
  wire [0:0] u_csamul_cla32_fa13_12_xor1;
  wire [0:0] u_csamul_cla32_fa13_12_or0;
  wire [0:0] u_csamul_cla32_and14_12;
  wire [0:0] u_csamul_cla32_fa14_12_xor1;
  wire [0:0] u_csamul_cla32_fa14_12_or0;
  wire [0:0] u_csamul_cla32_and15_12;
  wire [0:0] u_csamul_cla32_fa15_12_xor1;
  wire [0:0] u_csamul_cla32_fa15_12_or0;
  wire [0:0] u_csamul_cla32_and16_12;
  wire [0:0] u_csamul_cla32_fa16_12_xor1;
  wire [0:0] u_csamul_cla32_fa16_12_or0;
  wire [0:0] u_csamul_cla32_and17_12;
  wire [0:0] u_csamul_cla32_fa17_12_xor1;
  wire [0:0] u_csamul_cla32_fa17_12_or0;
  wire [0:0] u_csamul_cla32_and18_12;
  wire [0:0] u_csamul_cla32_fa18_12_xor1;
  wire [0:0] u_csamul_cla32_fa18_12_or0;
  wire [0:0] u_csamul_cla32_and19_12;
  wire [0:0] u_csamul_cla32_fa19_12_xor1;
  wire [0:0] u_csamul_cla32_fa19_12_or0;
  wire [0:0] u_csamul_cla32_and20_12;
  wire [0:0] u_csamul_cla32_fa20_12_xor1;
  wire [0:0] u_csamul_cla32_fa20_12_or0;
  wire [0:0] u_csamul_cla32_and21_12;
  wire [0:0] u_csamul_cla32_fa21_12_xor1;
  wire [0:0] u_csamul_cla32_fa21_12_or0;
  wire [0:0] u_csamul_cla32_and22_12;
  wire [0:0] u_csamul_cla32_fa22_12_xor1;
  wire [0:0] u_csamul_cla32_fa22_12_or0;
  wire [0:0] u_csamul_cla32_and23_12;
  wire [0:0] u_csamul_cla32_fa23_12_xor1;
  wire [0:0] u_csamul_cla32_fa23_12_or0;
  wire [0:0] u_csamul_cla32_and24_12;
  wire [0:0] u_csamul_cla32_fa24_12_xor1;
  wire [0:0] u_csamul_cla32_fa24_12_or0;
  wire [0:0] u_csamul_cla32_and25_12;
  wire [0:0] u_csamul_cla32_fa25_12_xor1;
  wire [0:0] u_csamul_cla32_fa25_12_or0;
  wire [0:0] u_csamul_cla32_and26_12;
  wire [0:0] u_csamul_cla32_fa26_12_xor1;
  wire [0:0] u_csamul_cla32_fa26_12_or0;
  wire [0:0] u_csamul_cla32_and27_12;
  wire [0:0] u_csamul_cla32_fa27_12_xor1;
  wire [0:0] u_csamul_cla32_fa27_12_or0;
  wire [0:0] u_csamul_cla32_and28_12;
  wire [0:0] u_csamul_cla32_fa28_12_xor1;
  wire [0:0] u_csamul_cla32_fa28_12_or0;
  wire [0:0] u_csamul_cla32_and29_12;
  wire [0:0] u_csamul_cla32_fa29_12_xor1;
  wire [0:0] u_csamul_cla32_fa29_12_or0;
  wire [0:0] u_csamul_cla32_and30_12;
  wire [0:0] u_csamul_cla32_fa30_12_xor1;
  wire [0:0] u_csamul_cla32_fa30_12_or0;
  wire [0:0] u_csamul_cla32_and31_12;
  wire [0:0] u_csamul_cla32_and0_13;
  wire [0:0] u_csamul_cla32_fa0_13_xor1;
  wire [0:0] u_csamul_cla32_fa0_13_or0;
  wire [0:0] u_csamul_cla32_and1_13;
  wire [0:0] u_csamul_cla32_fa1_13_xor1;
  wire [0:0] u_csamul_cla32_fa1_13_or0;
  wire [0:0] u_csamul_cla32_and2_13;
  wire [0:0] u_csamul_cla32_fa2_13_xor1;
  wire [0:0] u_csamul_cla32_fa2_13_or0;
  wire [0:0] u_csamul_cla32_and3_13;
  wire [0:0] u_csamul_cla32_fa3_13_xor1;
  wire [0:0] u_csamul_cla32_fa3_13_or0;
  wire [0:0] u_csamul_cla32_and4_13;
  wire [0:0] u_csamul_cla32_fa4_13_xor1;
  wire [0:0] u_csamul_cla32_fa4_13_or0;
  wire [0:0] u_csamul_cla32_and5_13;
  wire [0:0] u_csamul_cla32_fa5_13_xor1;
  wire [0:0] u_csamul_cla32_fa5_13_or0;
  wire [0:0] u_csamul_cla32_and6_13;
  wire [0:0] u_csamul_cla32_fa6_13_xor1;
  wire [0:0] u_csamul_cla32_fa6_13_or0;
  wire [0:0] u_csamul_cla32_and7_13;
  wire [0:0] u_csamul_cla32_fa7_13_xor1;
  wire [0:0] u_csamul_cla32_fa7_13_or0;
  wire [0:0] u_csamul_cla32_and8_13;
  wire [0:0] u_csamul_cla32_fa8_13_xor1;
  wire [0:0] u_csamul_cla32_fa8_13_or0;
  wire [0:0] u_csamul_cla32_and9_13;
  wire [0:0] u_csamul_cla32_fa9_13_xor1;
  wire [0:0] u_csamul_cla32_fa9_13_or0;
  wire [0:0] u_csamul_cla32_and10_13;
  wire [0:0] u_csamul_cla32_fa10_13_xor1;
  wire [0:0] u_csamul_cla32_fa10_13_or0;
  wire [0:0] u_csamul_cla32_and11_13;
  wire [0:0] u_csamul_cla32_fa11_13_xor1;
  wire [0:0] u_csamul_cla32_fa11_13_or0;
  wire [0:0] u_csamul_cla32_and12_13;
  wire [0:0] u_csamul_cla32_fa12_13_xor1;
  wire [0:0] u_csamul_cla32_fa12_13_or0;
  wire [0:0] u_csamul_cla32_and13_13;
  wire [0:0] u_csamul_cla32_fa13_13_xor1;
  wire [0:0] u_csamul_cla32_fa13_13_or0;
  wire [0:0] u_csamul_cla32_and14_13;
  wire [0:0] u_csamul_cla32_fa14_13_xor1;
  wire [0:0] u_csamul_cla32_fa14_13_or0;
  wire [0:0] u_csamul_cla32_and15_13;
  wire [0:0] u_csamul_cla32_fa15_13_xor1;
  wire [0:0] u_csamul_cla32_fa15_13_or0;
  wire [0:0] u_csamul_cla32_and16_13;
  wire [0:0] u_csamul_cla32_fa16_13_xor1;
  wire [0:0] u_csamul_cla32_fa16_13_or0;
  wire [0:0] u_csamul_cla32_and17_13;
  wire [0:0] u_csamul_cla32_fa17_13_xor1;
  wire [0:0] u_csamul_cla32_fa17_13_or0;
  wire [0:0] u_csamul_cla32_and18_13;
  wire [0:0] u_csamul_cla32_fa18_13_xor1;
  wire [0:0] u_csamul_cla32_fa18_13_or0;
  wire [0:0] u_csamul_cla32_and19_13;
  wire [0:0] u_csamul_cla32_fa19_13_xor1;
  wire [0:0] u_csamul_cla32_fa19_13_or0;
  wire [0:0] u_csamul_cla32_and20_13;
  wire [0:0] u_csamul_cla32_fa20_13_xor1;
  wire [0:0] u_csamul_cla32_fa20_13_or0;
  wire [0:0] u_csamul_cla32_and21_13;
  wire [0:0] u_csamul_cla32_fa21_13_xor1;
  wire [0:0] u_csamul_cla32_fa21_13_or0;
  wire [0:0] u_csamul_cla32_and22_13;
  wire [0:0] u_csamul_cla32_fa22_13_xor1;
  wire [0:0] u_csamul_cla32_fa22_13_or0;
  wire [0:0] u_csamul_cla32_and23_13;
  wire [0:0] u_csamul_cla32_fa23_13_xor1;
  wire [0:0] u_csamul_cla32_fa23_13_or0;
  wire [0:0] u_csamul_cla32_and24_13;
  wire [0:0] u_csamul_cla32_fa24_13_xor1;
  wire [0:0] u_csamul_cla32_fa24_13_or0;
  wire [0:0] u_csamul_cla32_and25_13;
  wire [0:0] u_csamul_cla32_fa25_13_xor1;
  wire [0:0] u_csamul_cla32_fa25_13_or0;
  wire [0:0] u_csamul_cla32_and26_13;
  wire [0:0] u_csamul_cla32_fa26_13_xor1;
  wire [0:0] u_csamul_cla32_fa26_13_or0;
  wire [0:0] u_csamul_cla32_and27_13;
  wire [0:0] u_csamul_cla32_fa27_13_xor1;
  wire [0:0] u_csamul_cla32_fa27_13_or0;
  wire [0:0] u_csamul_cla32_and28_13;
  wire [0:0] u_csamul_cla32_fa28_13_xor1;
  wire [0:0] u_csamul_cla32_fa28_13_or0;
  wire [0:0] u_csamul_cla32_and29_13;
  wire [0:0] u_csamul_cla32_fa29_13_xor1;
  wire [0:0] u_csamul_cla32_fa29_13_or0;
  wire [0:0] u_csamul_cla32_and30_13;
  wire [0:0] u_csamul_cla32_fa30_13_xor1;
  wire [0:0] u_csamul_cla32_fa30_13_or0;
  wire [0:0] u_csamul_cla32_and31_13;
  wire [0:0] u_csamul_cla32_and0_14;
  wire [0:0] u_csamul_cla32_fa0_14_xor1;
  wire [0:0] u_csamul_cla32_fa0_14_or0;
  wire [0:0] u_csamul_cla32_and1_14;
  wire [0:0] u_csamul_cla32_fa1_14_xor1;
  wire [0:0] u_csamul_cla32_fa1_14_or0;
  wire [0:0] u_csamul_cla32_and2_14;
  wire [0:0] u_csamul_cla32_fa2_14_xor1;
  wire [0:0] u_csamul_cla32_fa2_14_or0;
  wire [0:0] u_csamul_cla32_and3_14;
  wire [0:0] u_csamul_cla32_fa3_14_xor1;
  wire [0:0] u_csamul_cla32_fa3_14_or0;
  wire [0:0] u_csamul_cla32_and4_14;
  wire [0:0] u_csamul_cla32_fa4_14_xor1;
  wire [0:0] u_csamul_cla32_fa4_14_or0;
  wire [0:0] u_csamul_cla32_and5_14;
  wire [0:0] u_csamul_cla32_fa5_14_xor1;
  wire [0:0] u_csamul_cla32_fa5_14_or0;
  wire [0:0] u_csamul_cla32_and6_14;
  wire [0:0] u_csamul_cla32_fa6_14_xor1;
  wire [0:0] u_csamul_cla32_fa6_14_or0;
  wire [0:0] u_csamul_cla32_and7_14;
  wire [0:0] u_csamul_cla32_fa7_14_xor1;
  wire [0:0] u_csamul_cla32_fa7_14_or0;
  wire [0:0] u_csamul_cla32_and8_14;
  wire [0:0] u_csamul_cla32_fa8_14_xor1;
  wire [0:0] u_csamul_cla32_fa8_14_or0;
  wire [0:0] u_csamul_cla32_and9_14;
  wire [0:0] u_csamul_cla32_fa9_14_xor1;
  wire [0:0] u_csamul_cla32_fa9_14_or0;
  wire [0:0] u_csamul_cla32_and10_14;
  wire [0:0] u_csamul_cla32_fa10_14_xor1;
  wire [0:0] u_csamul_cla32_fa10_14_or0;
  wire [0:0] u_csamul_cla32_and11_14;
  wire [0:0] u_csamul_cla32_fa11_14_xor1;
  wire [0:0] u_csamul_cla32_fa11_14_or0;
  wire [0:0] u_csamul_cla32_and12_14;
  wire [0:0] u_csamul_cla32_fa12_14_xor1;
  wire [0:0] u_csamul_cla32_fa12_14_or0;
  wire [0:0] u_csamul_cla32_and13_14;
  wire [0:0] u_csamul_cla32_fa13_14_xor1;
  wire [0:0] u_csamul_cla32_fa13_14_or0;
  wire [0:0] u_csamul_cla32_and14_14;
  wire [0:0] u_csamul_cla32_fa14_14_xor1;
  wire [0:0] u_csamul_cla32_fa14_14_or0;
  wire [0:0] u_csamul_cla32_and15_14;
  wire [0:0] u_csamul_cla32_fa15_14_xor1;
  wire [0:0] u_csamul_cla32_fa15_14_or0;
  wire [0:0] u_csamul_cla32_and16_14;
  wire [0:0] u_csamul_cla32_fa16_14_xor1;
  wire [0:0] u_csamul_cla32_fa16_14_or0;
  wire [0:0] u_csamul_cla32_and17_14;
  wire [0:0] u_csamul_cla32_fa17_14_xor1;
  wire [0:0] u_csamul_cla32_fa17_14_or0;
  wire [0:0] u_csamul_cla32_and18_14;
  wire [0:0] u_csamul_cla32_fa18_14_xor1;
  wire [0:0] u_csamul_cla32_fa18_14_or0;
  wire [0:0] u_csamul_cla32_and19_14;
  wire [0:0] u_csamul_cla32_fa19_14_xor1;
  wire [0:0] u_csamul_cla32_fa19_14_or0;
  wire [0:0] u_csamul_cla32_and20_14;
  wire [0:0] u_csamul_cla32_fa20_14_xor1;
  wire [0:0] u_csamul_cla32_fa20_14_or0;
  wire [0:0] u_csamul_cla32_and21_14;
  wire [0:0] u_csamul_cla32_fa21_14_xor1;
  wire [0:0] u_csamul_cla32_fa21_14_or0;
  wire [0:0] u_csamul_cla32_and22_14;
  wire [0:0] u_csamul_cla32_fa22_14_xor1;
  wire [0:0] u_csamul_cla32_fa22_14_or0;
  wire [0:0] u_csamul_cla32_and23_14;
  wire [0:0] u_csamul_cla32_fa23_14_xor1;
  wire [0:0] u_csamul_cla32_fa23_14_or0;
  wire [0:0] u_csamul_cla32_and24_14;
  wire [0:0] u_csamul_cla32_fa24_14_xor1;
  wire [0:0] u_csamul_cla32_fa24_14_or0;
  wire [0:0] u_csamul_cla32_and25_14;
  wire [0:0] u_csamul_cla32_fa25_14_xor1;
  wire [0:0] u_csamul_cla32_fa25_14_or0;
  wire [0:0] u_csamul_cla32_and26_14;
  wire [0:0] u_csamul_cla32_fa26_14_xor1;
  wire [0:0] u_csamul_cla32_fa26_14_or0;
  wire [0:0] u_csamul_cla32_and27_14;
  wire [0:0] u_csamul_cla32_fa27_14_xor1;
  wire [0:0] u_csamul_cla32_fa27_14_or0;
  wire [0:0] u_csamul_cla32_and28_14;
  wire [0:0] u_csamul_cla32_fa28_14_xor1;
  wire [0:0] u_csamul_cla32_fa28_14_or0;
  wire [0:0] u_csamul_cla32_and29_14;
  wire [0:0] u_csamul_cla32_fa29_14_xor1;
  wire [0:0] u_csamul_cla32_fa29_14_or0;
  wire [0:0] u_csamul_cla32_and30_14;
  wire [0:0] u_csamul_cla32_fa30_14_xor1;
  wire [0:0] u_csamul_cla32_fa30_14_or0;
  wire [0:0] u_csamul_cla32_and31_14;
  wire [0:0] u_csamul_cla32_and0_15;
  wire [0:0] u_csamul_cla32_fa0_15_xor1;
  wire [0:0] u_csamul_cla32_fa0_15_or0;
  wire [0:0] u_csamul_cla32_and1_15;
  wire [0:0] u_csamul_cla32_fa1_15_xor1;
  wire [0:0] u_csamul_cla32_fa1_15_or0;
  wire [0:0] u_csamul_cla32_and2_15;
  wire [0:0] u_csamul_cla32_fa2_15_xor1;
  wire [0:0] u_csamul_cla32_fa2_15_or0;
  wire [0:0] u_csamul_cla32_and3_15;
  wire [0:0] u_csamul_cla32_fa3_15_xor1;
  wire [0:0] u_csamul_cla32_fa3_15_or0;
  wire [0:0] u_csamul_cla32_and4_15;
  wire [0:0] u_csamul_cla32_fa4_15_xor1;
  wire [0:0] u_csamul_cla32_fa4_15_or0;
  wire [0:0] u_csamul_cla32_and5_15;
  wire [0:0] u_csamul_cla32_fa5_15_xor1;
  wire [0:0] u_csamul_cla32_fa5_15_or0;
  wire [0:0] u_csamul_cla32_and6_15;
  wire [0:0] u_csamul_cla32_fa6_15_xor1;
  wire [0:0] u_csamul_cla32_fa6_15_or0;
  wire [0:0] u_csamul_cla32_and7_15;
  wire [0:0] u_csamul_cla32_fa7_15_xor1;
  wire [0:0] u_csamul_cla32_fa7_15_or0;
  wire [0:0] u_csamul_cla32_and8_15;
  wire [0:0] u_csamul_cla32_fa8_15_xor1;
  wire [0:0] u_csamul_cla32_fa8_15_or0;
  wire [0:0] u_csamul_cla32_and9_15;
  wire [0:0] u_csamul_cla32_fa9_15_xor1;
  wire [0:0] u_csamul_cla32_fa9_15_or0;
  wire [0:0] u_csamul_cla32_and10_15;
  wire [0:0] u_csamul_cla32_fa10_15_xor1;
  wire [0:0] u_csamul_cla32_fa10_15_or0;
  wire [0:0] u_csamul_cla32_and11_15;
  wire [0:0] u_csamul_cla32_fa11_15_xor1;
  wire [0:0] u_csamul_cla32_fa11_15_or0;
  wire [0:0] u_csamul_cla32_and12_15;
  wire [0:0] u_csamul_cla32_fa12_15_xor1;
  wire [0:0] u_csamul_cla32_fa12_15_or0;
  wire [0:0] u_csamul_cla32_and13_15;
  wire [0:0] u_csamul_cla32_fa13_15_xor1;
  wire [0:0] u_csamul_cla32_fa13_15_or0;
  wire [0:0] u_csamul_cla32_and14_15;
  wire [0:0] u_csamul_cla32_fa14_15_xor1;
  wire [0:0] u_csamul_cla32_fa14_15_or0;
  wire [0:0] u_csamul_cla32_and15_15;
  wire [0:0] u_csamul_cla32_fa15_15_xor1;
  wire [0:0] u_csamul_cla32_fa15_15_or0;
  wire [0:0] u_csamul_cla32_and16_15;
  wire [0:0] u_csamul_cla32_fa16_15_xor1;
  wire [0:0] u_csamul_cla32_fa16_15_or0;
  wire [0:0] u_csamul_cla32_and17_15;
  wire [0:0] u_csamul_cla32_fa17_15_xor1;
  wire [0:0] u_csamul_cla32_fa17_15_or0;
  wire [0:0] u_csamul_cla32_and18_15;
  wire [0:0] u_csamul_cla32_fa18_15_xor1;
  wire [0:0] u_csamul_cla32_fa18_15_or0;
  wire [0:0] u_csamul_cla32_and19_15;
  wire [0:0] u_csamul_cla32_fa19_15_xor1;
  wire [0:0] u_csamul_cla32_fa19_15_or0;
  wire [0:0] u_csamul_cla32_and20_15;
  wire [0:0] u_csamul_cla32_fa20_15_xor1;
  wire [0:0] u_csamul_cla32_fa20_15_or0;
  wire [0:0] u_csamul_cla32_and21_15;
  wire [0:0] u_csamul_cla32_fa21_15_xor1;
  wire [0:0] u_csamul_cla32_fa21_15_or0;
  wire [0:0] u_csamul_cla32_and22_15;
  wire [0:0] u_csamul_cla32_fa22_15_xor1;
  wire [0:0] u_csamul_cla32_fa22_15_or0;
  wire [0:0] u_csamul_cla32_and23_15;
  wire [0:0] u_csamul_cla32_fa23_15_xor1;
  wire [0:0] u_csamul_cla32_fa23_15_or0;
  wire [0:0] u_csamul_cla32_and24_15;
  wire [0:0] u_csamul_cla32_fa24_15_xor1;
  wire [0:0] u_csamul_cla32_fa24_15_or0;
  wire [0:0] u_csamul_cla32_and25_15;
  wire [0:0] u_csamul_cla32_fa25_15_xor1;
  wire [0:0] u_csamul_cla32_fa25_15_or0;
  wire [0:0] u_csamul_cla32_and26_15;
  wire [0:0] u_csamul_cla32_fa26_15_xor1;
  wire [0:0] u_csamul_cla32_fa26_15_or0;
  wire [0:0] u_csamul_cla32_and27_15;
  wire [0:0] u_csamul_cla32_fa27_15_xor1;
  wire [0:0] u_csamul_cla32_fa27_15_or0;
  wire [0:0] u_csamul_cla32_and28_15;
  wire [0:0] u_csamul_cla32_fa28_15_xor1;
  wire [0:0] u_csamul_cla32_fa28_15_or0;
  wire [0:0] u_csamul_cla32_and29_15;
  wire [0:0] u_csamul_cla32_fa29_15_xor1;
  wire [0:0] u_csamul_cla32_fa29_15_or0;
  wire [0:0] u_csamul_cla32_and30_15;
  wire [0:0] u_csamul_cla32_fa30_15_xor1;
  wire [0:0] u_csamul_cla32_fa30_15_or0;
  wire [0:0] u_csamul_cla32_and31_15;
  wire [0:0] u_csamul_cla32_and0_16;
  wire [0:0] u_csamul_cla32_fa0_16_xor1;
  wire [0:0] u_csamul_cla32_fa0_16_or0;
  wire [0:0] u_csamul_cla32_and1_16;
  wire [0:0] u_csamul_cla32_fa1_16_xor1;
  wire [0:0] u_csamul_cla32_fa1_16_or0;
  wire [0:0] u_csamul_cla32_and2_16;
  wire [0:0] u_csamul_cla32_fa2_16_xor1;
  wire [0:0] u_csamul_cla32_fa2_16_or0;
  wire [0:0] u_csamul_cla32_and3_16;
  wire [0:0] u_csamul_cla32_fa3_16_xor1;
  wire [0:0] u_csamul_cla32_fa3_16_or0;
  wire [0:0] u_csamul_cla32_and4_16;
  wire [0:0] u_csamul_cla32_fa4_16_xor1;
  wire [0:0] u_csamul_cla32_fa4_16_or0;
  wire [0:0] u_csamul_cla32_and5_16;
  wire [0:0] u_csamul_cla32_fa5_16_xor1;
  wire [0:0] u_csamul_cla32_fa5_16_or0;
  wire [0:0] u_csamul_cla32_and6_16;
  wire [0:0] u_csamul_cla32_fa6_16_xor1;
  wire [0:0] u_csamul_cla32_fa6_16_or0;
  wire [0:0] u_csamul_cla32_and7_16;
  wire [0:0] u_csamul_cla32_fa7_16_xor1;
  wire [0:0] u_csamul_cla32_fa7_16_or0;
  wire [0:0] u_csamul_cla32_and8_16;
  wire [0:0] u_csamul_cla32_fa8_16_xor1;
  wire [0:0] u_csamul_cla32_fa8_16_or0;
  wire [0:0] u_csamul_cla32_and9_16;
  wire [0:0] u_csamul_cla32_fa9_16_xor1;
  wire [0:0] u_csamul_cla32_fa9_16_or0;
  wire [0:0] u_csamul_cla32_and10_16;
  wire [0:0] u_csamul_cla32_fa10_16_xor1;
  wire [0:0] u_csamul_cla32_fa10_16_or0;
  wire [0:0] u_csamul_cla32_and11_16;
  wire [0:0] u_csamul_cla32_fa11_16_xor1;
  wire [0:0] u_csamul_cla32_fa11_16_or0;
  wire [0:0] u_csamul_cla32_and12_16;
  wire [0:0] u_csamul_cla32_fa12_16_xor1;
  wire [0:0] u_csamul_cla32_fa12_16_or0;
  wire [0:0] u_csamul_cla32_and13_16;
  wire [0:0] u_csamul_cla32_fa13_16_xor1;
  wire [0:0] u_csamul_cla32_fa13_16_or0;
  wire [0:0] u_csamul_cla32_and14_16;
  wire [0:0] u_csamul_cla32_fa14_16_xor1;
  wire [0:0] u_csamul_cla32_fa14_16_or0;
  wire [0:0] u_csamul_cla32_and15_16;
  wire [0:0] u_csamul_cla32_fa15_16_xor1;
  wire [0:0] u_csamul_cla32_fa15_16_or0;
  wire [0:0] u_csamul_cla32_and16_16;
  wire [0:0] u_csamul_cla32_fa16_16_xor1;
  wire [0:0] u_csamul_cla32_fa16_16_or0;
  wire [0:0] u_csamul_cla32_and17_16;
  wire [0:0] u_csamul_cla32_fa17_16_xor1;
  wire [0:0] u_csamul_cla32_fa17_16_or0;
  wire [0:0] u_csamul_cla32_and18_16;
  wire [0:0] u_csamul_cla32_fa18_16_xor1;
  wire [0:0] u_csamul_cla32_fa18_16_or0;
  wire [0:0] u_csamul_cla32_and19_16;
  wire [0:0] u_csamul_cla32_fa19_16_xor1;
  wire [0:0] u_csamul_cla32_fa19_16_or0;
  wire [0:0] u_csamul_cla32_and20_16;
  wire [0:0] u_csamul_cla32_fa20_16_xor1;
  wire [0:0] u_csamul_cla32_fa20_16_or0;
  wire [0:0] u_csamul_cla32_and21_16;
  wire [0:0] u_csamul_cla32_fa21_16_xor1;
  wire [0:0] u_csamul_cla32_fa21_16_or0;
  wire [0:0] u_csamul_cla32_and22_16;
  wire [0:0] u_csamul_cla32_fa22_16_xor1;
  wire [0:0] u_csamul_cla32_fa22_16_or0;
  wire [0:0] u_csamul_cla32_and23_16;
  wire [0:0] u_csamul_cla32_fa23_16_xor1;
  wire [0:0] u_csamul_cla32_fa23_16_or0;
  wire [0:0] u_csamul_cla32_and24_16;
  wire [0:0] u_csamul_cla32_fa24_16_xor1;
  wire [0:0] u_csamul_cla32_fa24_16_or0;
  wire [0:0] u_csamul_cla32_and25_16;
  wire [0:0] u_csamul_cla32_fa25_16_xor1;
  wire [0:0] u_csamul_cla32_fa25_16_or0;
  wire [0:0] u_csamul_cla32_and26_16;
  wire [0:0] u_csamul_cla32_fa26_16_xor1;
  wire [0:0] u_csamul_cla32_fa26_16_or0;
  wire [0:0] u_csamul_cla32_and27_16;
  wire [0:0] u_csamul_cla32_fa27_16_xor1;
  wire [0:0] u_csamul_cla32_fa27_16_or0;
  wire [0:0] u_csamul_cla32_and28_16;
  wire [0:0] u_csamul_cla32_fa28_16_xor1;
  wire [0:0] u_csamul_cla32_fa28_16_or0;
  wire [0:0] u_csamul_cla32_and29_16;
  wire [0:0] u_csamul_cla32_fa29_16_xor1;
  wire [0:0] u_csamul_cla32_fa29_16_or0;
  wire [0:0] u_csamul_cla32_and30_16;
  wire [0:0] u_csamul_cla32_fa30_16_xor1;
  wire [0:0] u_csamul_cla32_fa30_16_or0;
  wire [0:0] u_csamul_cla32_and31_16;
  wire [0:0] u_csamul_cla32_and0_17;
  wire [0:0] u_csamul_cla32_fa0_17_xor1;
  wire [0:0] u_csamul_cla32_fa0_17_or0;
  wire [0:0] u_csamul_cla32_and1_17;
  wire [0:0] u_csamul_cla32_fa1_17_xor1;
  wire [0:0] u_csamul_cla32_fa1_17_or0;
  wire [0:0] u_csamul_cla32_and2_17;
  wire [0:0] u_csamul_cla32_fa2_17_xor1;
  wire [0:0] u_csamul_cla32_fa2_17_or0;
  wire [0:0] u_csamul_cla32_and3_17;
  wire [0:0] u_csamul_cla32_fa3_17_xor1;
  wire [0:0] u_csamul_cla32_fa3_17_or0;
  wire [0:0] u_csamul_cla32_and4_17;
  wire [0:0] u_csamul_cla32_fa4_17_xor1;
  wire [0:0] u_csamul_cla32_fa4_17_or0;
  wire [0:0] u_csamul_cla32_and5_17;
  wire [0:0] u_csamul_cla32_fa5_17_xor1;
  wire [0:0] u_csamul_cla32_fa5_17_or0;
  wire [0:0] u_csamul_cla32_and6_17;
  wire [0:0] u_csamul_cla32_fa6_17_xor1;
  wire [0:0] u_csamul_cla32_fa6_17_or0;
  wire [0:0] u_csamul_cla32_and7_17;
  wire [0:0] u_csamul_cla32_fa7_17_xor1;
  wire [0:0] u_csamul_cla32_fa7_17_or0;
  wire [0:0] u_csamul_cla32_and8_17;
  wire [0:0] u_csamul_cla32_fa8_17_xor1;
  wire [0:0] u_csamul_cla32_fa8_17_or0;
  wire [0:0] u_csamul_cla32_and9_17;
  wire [0:0] u_csamul_cla32_fa9_17_xor1;
  wire [0:0] u_csamul_cla32_fa9_17_or0;
  wire [0:0] u_csamul_cla32_and10_17;
  wire [0:0] u_csamul_cla32_fa10_17_xor1;
  wire [0:0] u_csamul_cla32_fa10_17_or0;
  wire [0:0] u_csamul_cla32_and11_17;
  wire [0:0] u_csamul_cla32_fa11_17_xor1;
  wire [0:0] u_csamul_cla32_fa11_17_or0;
  wire [0:0] u_csamul_cla32_and12_17;
  wire [0:0] u_csamul_cla32_fa12_17_xor1;
  wire [0:0] u_csamul_cla32_fa12_17_or0;
  wire [0:0] u_csamul_cla32_and13_17;
  wire [0:0] u_csamul_cla32_fa13_17_xor1;
  wire [0:0] u_csamul_cla32_fa13_17_or0;
  wire [0:0] u_csamul_cla32_and14_17;
  wire [0:0] u_csamul_cla32_fa14_17_xor1;
  wire [0:0] u_csamul_cla32_fa14_17_or0;
  wire [0:0] u_csamul_cla32_and15_17;
  wire [0:0] u_csamul_cla32_fa15_17_xor1;
  wire [0:0] u_csamul_cla32_fa15_17_or0;
  wire [0:0] u_csamul_cla32_and16_17;
  wire [0:0] u_csamul_cla32_fa16_17_xor1;
  wire [0:0] u_csamul_cla32_fa16_17_or0;
  wire [0:0] u_csamul_cla32_and17_17;
  wire [0:0] u_csamul_cla32_fa17_17_xor1;
  wire [0:0] u_csamul_cla32_fa17_17_or0;
  wire [0:0] u_csamul_cla32_and18_17;
  wire [0:0] u_csamul_cla32_fa18_17_xor1;
  wire [0:0] u_csamul_cla32_fa18_17_or0;
  wire [0:0] u_csamul_cla32_and19_17;
  wire [0:0] u_csamul_cla32_fa19_17_xor1;
  wire [0:0] u_csamul_cla32_fa19_17_or0;
  wire [0:0] u_csamul_cla32_and20_17;
  wire [0:0] u_csamul_cla32_fa20_17_xor1;
  wire [0:0] u_csamul_cla32_fa20_17_or0;
  wire [0:0] u_csamul_cla32_and21_17;
  wire [0:0] u_csamul_cla32_fa21_17_xor1;
  wire [0:0] u_csamul_cla32_fa21_17_or0;
  wire [0:0] u_csamul_cla32_and22_17;
  wire [0:0] u_csamul_cla32_fa22_17_xor1;
  wire [0:0] u_csamul_cla32_fa22_17_or0;
  wire [0:0] u_csamul_cla32_and23_17;
  wire [0:0] u_csamul_cla32_fa23_17_xor1;
  wire [0:0] u_csamul_cla32_fa23_17_or0;
  wire [0:0] u_csamul_cla32_and24_17;
  wire [0:0] u_csamul_cla32_fa24_17_xor1;
  wire [0:0] u_csamul_cla32_fa24_17_or0;
  wire [0:0] u_csamul_cla32_and25_17;
  wire [0:0] u_csamul_cla32_fa25_17_xor1;
  wire [0:0] u_csamul_cla32_fa25_17_or0;
  wire [0:0] u_csamul_cla32_and26_17;
  wire [0:0] u_csamul_cla32_fa26_17_xor1;
  wire [0:0] u_csamul_cla32_fa26_17_or0;
  wire [0:0] u_csamul_cla32_and27_17;
  wire [0:0] u_csamul_cla32_fa27_17_xor1;
  wire [0:0] u_csamul_cla32_fa27_17_or0;
  wire [0:0] u_csamul_cla32_and28_17;
  wire [0:0] u_csamul_cla32_fa28_17_xor1;
  wire [0:0] u_csamul_cla32_fa28_17_or0;
  wire [0:0] u_csamul_cla32_and29_17;
  wire [0:0] u_csamul_cla32_fa29_17_xor1;
  wire [0:0] u_csamul_cla32_fa29_17_or0;
  wire [0:0] u_csamul_cla32_and30_17;
  wire [0:0] u_csamul_cla32_fa30_17_xor1;
  wire [0:0] u_csamul_cla32_fa30_17_or0;
  wire [0:0] u_csamul_cla32_and31_17;
  wire [0:0] u_csamul_cla32_and0_18;
  wire [0:0] u_csamul_cla32_fa0_18_xor1;
  wire [0:0] u_csamul_cla32_fa0_18_or0;
  wire [0:0] u_csamul_cla32_and1_18;
  wire [0:0] u_csamul_cla32_fa1_18_xor1;
  wire [0:0] u_csamul_cla32_fa1_18_or0;
  wire [0:0] u_csamul_cla32_and2_18;
  wire [0:0] u_csamul_cla32_fa2_18_xor1;
  wire [0:0] u_csamul_cla32_fa2_18_or0;
  wire [0:0] u_csamul_cla32_and3_18;
  wire [0:0] u_csamul_cla32_fa3_18_xor1;
  wire [0:0] u_csamul_cla32_fa3_18_or0;
  wire [0:0] u_csamul_cla32_and4_18;
  wire [0:0] u_csamul_cla32_fa4_18_xor1;
  wire [0:0] u_csamul_cla32_fa4_18_or0;
  wire [0:0] u_csamul_cla32_and5_18;
  wire [0:0] u_csamul_cla32_fa5_18_xor1;
  wire [0:0] u_csamul_cla32_fa5_18_or0;
  wire [0:0] u_csamul_cla32_and6_18;
  wire [0:0] u_csamul_cla32_fa6_18_xor1;
  wire [0:0] u_csamul_cla32_fa6_18_or0;
  wire [0:0] u_csamul_cla32_and7_18;
  wire [0:0] u_csamul_cla32_fa7_18_xor1;
  wire [0:0] u_csamul_cla32_fa7_18_or0;
  wire [0:0] u_csamul_cla32_and8_18;
  wire [0:0] u_csamul_cla32_fa8_18_xor1;
  wire [0:0] u_csamul_cla32_fa8_18_or0;
  wire [0:0] u_csamul_cla32_and9_18;
  wire [0:0] u_csamul_cla32_fa9_18_xor1;
  wire [0:0] u_csamul_cla32_fa9_18_or0;
  wire [0:0] u_csamul_cla32_and10_18;
  wire [0:0] u_csamul_cla32_fa10_18_xor1;
  wire [0:0] u_csamul_cla32_fa10_18_or0;
  wire [0:0] u_csamul_cla32_and11_18;
  wire [0:0] u_csamul_cla32_fa11_18_xor1;
  wire [0:0] u_csamul_cla32_fa11_18_or0;
  wire [0:0] u_csamul_cla32_and12_18;
  wire [0:0] u_csamul_cla32_fa12_18_xor1;
  wire [0:0] u_csamul_cla32_fa12_18_or0;
  wire [0:0] u_csamul_cla32_and13_18;
  wire [0:0] u_csamul_cla32_fa13_18_xor1;
  wire [0:0] u_csamul_cla32_fa13_18_or0;
  wire [0:0] u_csamul_cla32_and14_18;
  wire [0:0] u_csamul_cla32_fa14_18_xor1;
  wire [0:0] u_csamul_cla32_fa14_18_or0;
  wire [0:0] u_csamul_cla32_and15_18;
  wire [0:0] u_csamul_cla32_fa15_18_xor1;
  wire [0:0] u_csamul_cla32_fa15_18_or0;
  wire [0:0] u_csamul_cla32_and16_18;
  wire [0:0] u_csamul_cla32_fa16_18_xor1;
  wire [0:0] u_csamul_cla32_fa16_18_or0;
  wire [0:0] u_csamul_cla32_and17_18;
  wire [0:0] u_csamul_cla32_fa17_18_xor1;
  wire [0:0] u_csamul_cla32_fa17_18_or0;
  wire [0:0] u_csamul_cla32_and18_18;
  wire [0:0] u_csamul_cla32_fa18_18_xor1;
  wire [0:0] u_csamul_cla32_fa18_18_or0;
  wire [0:0] u_csamul_cla32_and19_18;
  wire [0:0] u_csamul_cla32_fa19_18_xor1;
  wire [0:0] u_csamul_cla32_fa19_18_or0;
  wire [0:0] u_csamul_cla32_and20_18;
  wire [0:0] u_csamul_cla32_fa20_18_xor1;
  wire [0:0] u_csamul_cla32_fa20_18_or0;
  wire [0:0] u_csamul_cla32_and21_18;
  wire [0:0] u_csamul_cla32_fa21_18_xor1;
  wire [0:0] u_csamul_cla32_fa21_18_or0;
  wire [0:0] u_csamul_cla32_and22_18;
  wire [0:0] u_csamul_cla32_fa22_18_xor1;
  wire [0:0] u_csamul_cla32_fa22_18_or0;
  wire [0:0] u_csamul_cla32_and23_18;
  wire [0:0] u_csamul_cla32_fa23_18_xor1;
  wire [0:0] u_csamul_cla32_fa23_18_or0;
  wire [0:0] u_csamul_cla32_and24_18;
  wire [0:0] u_csamul_cla32_fa24_18_xor1;
  wire [0:0] u_csamul_cla32_fa24_18_or0;
  wire [0:0] u_csamul_cla32_and25_18;
  wire [0:0] u_csamul_cla32_fa25_18_xor1;
  wire [0:0] u_csamul_cla32_fa25_18_or0;
  wire [0:0] u_csamul_cla32_and26_18;
  wire [0:0] u_csamul_cla32_fa26_18_xor1;
  wire [0:0] u_csamul_cla32_fa26_18_or0;
  wire [0:0] u_csamul_cla32_and27_18;
  wire [0:0] u_csamul_cla32_fa27_18_xor1;
  wire [0:0] u_csamul_cla32_fa27_18_or0;
  wire [0:0] u_csamul_cla32_and28_18;
  wire [0:0] u_csamul_cla32_fa28_18_xor1;
  wire [0:0] u_csamul_cla32_fa28_18_or0;
  wire [0:0] u_csamul_cla32_and29_18;
  wire [0:0] u_csamul_cla32_fa29_18_xor1;
  wire [0:0] u_csamul_cla32_fa29_18_or0;
  wire [0:0] u_csamul_cla32_and30_18;
  wire [0:0] u_csamul_cla32_fa30_18_xor1;
  wire [0:0] u_csamul_cla32_fa30_18_or0;
  wire [0:0] u_csamul_cla32_and31_18;
  wire [0:0] u_csamul_cla32_and0_19;
  wire [0:0] u_csamul_cla32_fa0_19_xor1;
  wire [0:0] u_csamul_cla32_fa0_19_or0;
  wire [0:0] u_csamul_cla32_and1_19;
  wire [0:0] u_csamul_cla32_fa1_19_xor1;
  wire [0:0] u_csamul_cla32_fa1_19_or0;
  wire [0:0] u_csamul_cla32_and2_19;
  wire [0:0] u_csamul_cla32_fa2_19_xor1;
  wire [0:0] u_csamul_cla32_fa2_19_or0;
  wire [0:0] u_csamul_cla32_and3_19;
  wire [0:0] u_csamul_cla32_fa3_19_xor1;
  wire [0:0] u_csamul_cla32_fa3_19_or0;
  wire [0:0] u_csamul_cla32_and4_19;
  wire [0:0] u_csamul_cla32_fa4_19_xor1;
  wire [0:0] u_csamul_cla32_fa4_19_or0;
  wire [0:0] u_csamul_cla32_and5_19;
  wire [0:0] u_csamul_cla32_fa5_19_xor1;
  wire [0:0] u_csamul_cla32_fa5_19_or0;
  wire [0:0] u_csamul_cla32_and6_19;
  wire [0:0] u_csamul_cla32_fa6_19_xor1;
  wire [0:0] u_csamul_cla32_fa6_19_or0;
  wire [0:0] u_csamul_cla32_and7_19;
  wire [0:0] u_csamul_cla32_fa7_19_xor1;
  wire [0:0] u_csamul_cla32_fa7_19_or0;
  wire [0:0] u_csamul_cla32_and8_19;
  wire [0:0] u_csamul_cla32_fa8_19_xor1;
  wire [0:0] u_csamul_cla32_fa8_19_or0;
  wire [0:0] u_csamul_cla32_and9_19;
  wire [0:0] u_csamul_cla32_fa9_19_xor1;
  wire [0:0] u_csamul_cla32_fa9_19_or0;
  wire [0:0] u_csamul_cla32_and10_19;
  wire [0:0] u_csamul_cla32_fa10_19_xor1;
  wire [0:0] u_csamul_cla32_fa10_19_or0;
  wire [0:0] u_csamul_cla32_and11_19;
  wire [0:0] u_csamul_cla32_fa11_19_xor1;
  wire [0:0] u_csamul_cla32_fa11_19_or0;
  wire [0:0] u_csamul_cla32_and12_19;
  wire [0:0] u_csamul_cla32_fa12_19_xor1;
  wire [0:0] u_csamul_cla32_fa12_19_or0;
  wire [0:0] u_csamul_cla32_and13_19;
  wire [0:0] u_csamul_cla32_fa13_19_xor1;
  wire [0:0] u_csamul_cla32_fa13_19_or0;
  wire [0:0] u_csamul_cla32_and14_19;
  wire [0:0] u_csamul_cla32_fa14_19_xor1;
  wire [0:0] u_csamul_cla32_fa14_19_or0;
  wire [0:0] u_csamul_cla32_and15_19;
  wire [0:0] u_csamul_cla32_fa15_19_xor1;
  wire [0:0] u_csamul_cla32_fa15_19_or0;
  wire [0:0] u_csamul_cla32_and16_19;
  wire [0:0] u_csamul_cla32_fa16_19_xor1;
  wire [0:0] u_csamul_cla32_fa16_19_or0;
  wire [0:0] u_csamul_cla32_and17_19;
  wire [0:0] u_csamul_cla32_fa17_19_xor1;
  wire [0:0] u_csamul_cla32_fa17_19_or0;
  wire [0:0] u_csamul_cla32_and18_19;
  wire [0:0] u_csamul_cla32_fa18_19_xor1;
  wire [0:0] u_csamul_cla32_fa18_19_or0;
  wire [0:0] u_csamul_cla32_and19_19;
  wire [0:0] u_csamul_cla32_fa19_19_xor1;
  wire [0:0] u_csamul_cla32_fa19_19_or0;
  wire [0:0] u_csamul_cla32_and20_19;
  wire [0:0] u_csamul_cla32_fa20_19_xor1;
  wire [0:0] u_csamul_cla32_fa20_19_or0;
  wire [0:0] u_csamul_cla32_and21_19;
  wire [0:0] u_csamul_cla32_fa21_19_xor1;
  wire [0:0] u_csamul_cla32_fa21_19_or0;
  wire [0:0] u_csamul_cla32_and22_19;
  wire [0:0] u_csamul_cla32_fa22_19_xor1;
  wire [0:0] u_csamul_cla32_fa22_19_or0;
  wire [0:0] u_csamul_cla32_and23_19;
  wire [0:0] u_csamul_cla32_fa23_19_xor1;
  wire [0:0] u_csamul_cla32_fa23_19_or0;
  wire [0:0] u_csamul_cla32_and24_19;
  wire [0:0] u_csamul_cla32_fa24_19_xor1;
  wire [0:0] u_csamul_cla32_fa24_19_or0;
  wire [0:0] u_csamul_cla32_and25_19;
  wire [0:0] u_csamul_cla32_fa25_19_xor1;
  wire [0:0] u_csamul_cla32_fa25_19_or0;
  wire [0:0] u_csamul_cla32_and26_19;
  wire [0:0] u_csamul_cla32_fa26_19_xor1;
  wire [0:0] u_csamul_cla32_fa26_19_or0;
  wire [0:0] u_csamul_cla32_and27_19;
  wire [0:0] u_csamul_cla32_fa27_19_xor1;
  wire [0:0] u_csamul_cla32_fa27_19_or0;
  wire [0:0] u_csamul_cla32_and28_19;
  wire [0:0] u_csamul_cla32_fa28_19_xor1;
  wire [0:0] u_csamul_cla32_fa28_19_or0;
  wire [0:0] u_csamul_cla32_and29_19;
  wire [0:0] u_csamul_cla32_fa29_19_xor1;
  wire [0:0] u_csamul_cla32_fa29_19_or0;
  wire [0:0] u_csamul_cla32_and30_19;
  wire [0:0] u_csamul_cla32_fa30_19_xor1;
  wire [0:0] u_csamul_cla32_fa30_19_or0;
  wire [0:0] u_csamul_cla32_and31_19;
  wire [0:0] u_csamul_cla32_and0_20;
  wire [0:0] u_csamul_cla32_fa0_20_xor1;
  wire [0:0] u_csamul_cla32_fa0_20_or0;
  wire [0:0] u_csamul_cla32_and1_20;
  wire [0:0] u_csamul_cla32_fa1_20_xor1;
  wire [0:0] u_csamul_cla32_fa1_20_or0;
  wire [0:0] u_csamul_cla32_and2_20;
  wire [0:0] u_csamul_cla32_fa2_20_xor1;
  wire [0:0] u_csamul_cla32_fa2_20_or0;
  wire [0:0] u_csamul_cla32_and3_20;
  wire [0:0] u_csamul_cla32_fa3_20_xor1;
  wire [0:0] u_csamul_cla32_fa3_20_or0;
  wire [0:0] u_csamul_cla32_and4_20;
  wire [0:0] u_csamul_cla32_fa4_20_xor1;
  wire [0:0] u_csamul_cla32_fa4_20_or0;
  wire [0:0] u_csamul_cla32_and5_20;
  wire [0:0] u_csamul_cla32_fa5_20_xor1;
  wire [0:0] u_csamul_cla32_fa5_20_or0;
  wire [0:0] u_csamul_cla32_and6_20;
  wire [0:0] u_csamul_cla32_fa6_20_xor1;
  wire [0:0] u_csamul_cla32_fa6_20_or0;
  wire [0:0] u_csamul_cla32_and7_20;
  wire [0:0] u_csamul_cla32_fa7_20_xor1;
  wire [0:0] u_csamul_cla32_fa7_20_or0;
  wire [0:0] u_csamul_cla32_and8_20;
  wire [0:0] u_csamul_cla32_fa8_20_xor1;
  wire [0:0] u_csamul_cla32_fa8_20_or0;
  wire [0:0] u_csamul_cla32_and9_20;
  wire [0:0] u_csamul_cla32_fa9_20_xor1;
  wire [0:0] u_csamul_cla32_fa9_20_or0;
  wire [0:0] u_csamul_cla32_and10_20;
  wire [0:0] u_csamul_cla32_fa10_20_xor1;
  wire [0:0] u_csamul_cla32_fa10_20_or0;
  wire [0:0] u_csamul_cla32_and11_20;
  wire [0:0] u_csamul_cla32_fa11_20_xor1;
  wire [0:0] u_csamul_cla32_fa11_20_or0;
  wire [0:0] u_csamul_cla32_and12_20;
  wire [0:0] u_csamul_cla32_fa12_20_xor1;
  wire [0:0] u_csamul_cla32_fa12_20_or0;
  wire [0:0] u_csamul_cla32_and13_20;
  wire [0:0] u_csamul_cla32_fa13_20_xor1;
  wire [0:0] u_csamul_cla32_fa13_20_or0;
  wire [0:0] u_csamul_cla32_and14_20;
  wire [0:0] u_csamul_cla32_fa14_20_xor1;
  wire [0:0] u_csamul_cla32_fa14_20_or0;
  wire [0:0] u_csamul_cla32_and15_20;
  wire [0:0] u_csamul_cla32_fa15_20_xor1;
  wire [0:0] u_csamul_cla32_fa15_20_or0;
  wire [0:0] u_csamul_cla32_and16_20;
  wire [0:0] u_csamul_cla32_fa16_20_xor1;
  wire [0:0] u_csamul_cla32_fa16_20_or0;
  wire [0:0] u_csamul_cla32_and17_20;
  wire [0:0] u_csamul_cla32_fa17_20_xor1;
  wire [0:0] u_csamul_cla32_fa17_20_or0;
  wire [0:0] u_csamul_cla32_and18_20;
  wire [0:0] u_csamul_cla32_fa18_20_xor1;
  wire [0:0] u_csamul_cla32_fa18_20_or0;
  wire [0:0] u_csamul_cla32_and19_20;
  wire [0:0] u_csamul_cla32_fa19_20_xor1;
  wire [0:0] u_csamul_cla32_fa19_20_or0;
  wire [0:0] u_csamul_cla32_and20_20;
  wire [0:0] u_csamul_cla32_fa20_20_xor1;
  wire [0:0] u_csamul_cla32_fa20_20_or0;
  wire [0:0] u_csamul_cla32_and21_20;
  wire [0:0] u_csamul_cla32_fa21_20_xor1;
  wire [0:0] u_csamul_cla32_fa21_20_or0;
  wire [0:0] u_csamul_cla32_and22_20;
  wire [0:0] u_csamul_cla32_fa22_20_xor1;
  wire [0:0] u_csamul_cla32_fa22_20_or0;
  wire [0:0] u_csamul_cla32_and23_20;
  wire [0:0] u_csamul_cla32_fa23_20_xor1;
  wire [0:0] u_csamul_cla32_fa23_20_or0;
  wire [0:0] u_csamul_cla32_and24_20;
  wire [0:0] u_csamul_cla32_fa24_20_xor1;
  wire [0:0] u_csamul_cla32_fa24_20_or0;
  wire [0:0] u_csamul_cla32_and25_20;
  wire [0:0] u_csamul_cla32_fa25_20_xor1;
  wire [0:0] u_csamul_cla32_fa25_20_or0;
  wire [0:0] u_csamul_cla32_and26_20;
  wire [0:0] u_csamul_cla32_fa26_20_xor1;
  wire [0:0] u_csamul_cla32_fa26_20_or0;
  wire [0:0] u_csamul_cla32_and27_20;
  wire [0:0] u_csamul_cla32_fa27_20_xor1;
  wire [0:0] u_csamul_cla32_fa27_20_or0;
  wire [0:0] u_csamul_cla32_and28_20;
  wire [0:0] u_csamul_cla32_fa28_20_xor1;
  wire [0:0] u_csamul_cla32_fa28_20_or0;
  wire [0:0] u_csamul_cla32_and29_20;
  wire [0:0] u_csamul_cla32_fa29_20_xor1;
  wire [0:0] u_csamul_cla32_fa29_20_or0;
  wire [0:0] u_csamul_cla32_and30_20;
  wire [0:0] u_csamul_cla32_fa30_20_xor1;
  wire [0:0] u_csamul_cla32_fa30_20_or0;
  wire [0:0] u_csamul_cla32_and31_20;
  wire [0:0] u_csamul_cla32_and0_21;
  wire [0:0] u_csamul_cla32_fa0_21_xor1;
  wire [0:0] u_csamul_cla32_fa0_21_or0;
  wire [0:0] u_csamul_cla32_and1_21;
  wire [0:0] u_csamul_cla32_fa1_21_xor1;
  wire [0:0] u_csamul_cla32_fa1_21_or0;
  wire [0:0] u_csamul_cla32_and2_21;
  wire [0:0] u_csamul_cla32_fa2_21_xor1;
  wire [0:0] u_csamul_cla32_fa2_21_or0;
  wire [0:0] u_csamul_cla32_and3_21;
  wire [0:0] u_csamul_cla32_fa3_21_xor1;
  wire [0:0] u_csamul_cla32_fa3_21_or0;
  wire [0:0] u_csamul_cla32_and4_21;
  wire [0:0] u_csamul_cla32_fa4_21_xor1;
  wire [0:0] u_csamul_cla32_fa4_21_or0;
  wire [0:0] u_csamul_cla32_and5_21;
  wire [0:0] u_csamul_cla32_fa5_21_xor1;
  wire [0:0] u_csamul_cla32_fa5_21_or0;
  wire [0:0] u_csamul_cla32_and6_21;
  wire [0:0] u_csamul_cla32_fa6_21_xor1;
  wire [0:0] u_csamul_cla32_fa6_21_or0;
  wire [0:0] u_csamul_cla32_and7_21;
  wire [0:0] u_csamul_cla32_fa7_21_xor1;
  wire [0:0] u_csamul_cla32_fa7_21_or0;
  wire [0:0] u_csamul_cla32_and8_21;
  wire [0:0] u_csamul_cla32_fa8_21_xor1;
  wire [0:0] u_csamul_cla32_fa8_21_or0;
  wire [0:0] u_csamul_cla32_and9_21;
  wire [0:0] u_csamul_cla32_fa9_21_xor1;
  wire [0:0] u_csamul_cla32_fa9_21_or0;
  wire [0:0] u_csamul_cla32_and10_21;
  wire [0:0] u_csamul_cla32_fa10_21_xor1;
  wire [0:0] u_csamul_cla32_fa10_21_or0;
  wire [0:0] u_csamul_cla32_and11_21;
  wire [0:0] u_csamul_cla32_fa11_21_xor1;
  wire [0:0] u_csamul_cla32_fa11_21_or0;
  wire [0:0] u_csamul_cla32_and12_21;
  wire [0:0] u_csamul_cla32_fa12_21_xor1;
  wire [0:0] u_csamul_cla32_fa12_21_or0;
  wire [0:0] u_csamul_cla32_and13_21;
  wire [0:0] u_csamul_cla32_fa13_21_xor1;
  wire [0:0] u_csamul_cla32_fa13_21_or0;
  wire [0:0] u_csamul_cla32_and14_21;
  wire [0:0] u_csamul_cla32_fa14_21_xor1;
  wire [0:0] u_csamul_cla32_fa14_21_or0;
  wire [0:0] u_csamul_cla32_and15_21;
  wire [0:0] u_csamul_cla32_fa15_21_xor1;
  wire [0:0] u_csamul_cla32_fa15_21_or0;
  wire [0:0] u_csamul_cla32_and16_21;
  wire [0:0] u_csamul_cla32_fa16_21_xor1;
  wire [0:0] u_csamul_cla32_fa16_21_or0;
  wire [0:0] u_csamul_cla32_and17_21;
  wire [0:0] u_csamul_cla32_fa17_21_xor1;
  wire [0:0] u_csamul_cla32_fa17_21_or0;
  wire [0:0] u_csamul_cla32_and18_21;
  wire [0:0] u_csamul_cla32_fa18_21_xor1;
  wire [0:0] u_csamul_cla32_fa18_21_or0;
  wire [0:0] u_csamul_cla32_and19_21;
  wire [0:0] u_csamul_cla32_fa19_21_xor1;
  wire [0:0] u_csamul_cla32_fa19_21_or0;
  wire [0:0] u_csamul_cla32_and20_21;
  wire [0:0] u_csamul_cla32_fa20_21_xor1;
  wire [0:0] u_csamul_cla32_fa20_21_or0;
  wire [0:0] u_csamul_cla32_and21_21;
  wire [0:0] u_csamul_cla32_fa21_21_xor1;
  wire [0:0] u_csamul_cla32_fa21_21_or0;
  wire [0:0] u_csamul_cla32_and22_21;
  wire [0:0] u_csamul_cla32_fa22_21_xor1;
  wire [0:0] u_csamul_cla32_fa22_21_or0;
  wire [0:0] u_csamul_cla32_and23_21;
  wire [0:0] u_csamul_cla32_fa23_21_xor1;
  wire [0:0] u_csamul_cla32_fa23_21_or0;
  wire [0:0] u_csamul_cla32_and24_21;
  wire [0:0] u_csamul_cla32_fa24_21_xor1;
  wire [0:0] u_csamul_cla32_fa24_21_or0;
  wire [0:0] u_csamul_cla32_and25_21;
  wire [0:0] u_csamul_cla32_fa25_21_xor1;
  wire [0:0] u_csamul_cla32_fa25_21_or0;
  wire [0:0] u_csamul_cla32_and26_21;
  wire [0:0] u_csamul_cla32_fa26_21_xor1;
  wire [0:0] u_csamul_cla32_fa26_21_or0;
  wire [0:0] u_csamul_cla32_and27_21;
  wire [0:0] u_csamul_cla32_fa27_21_xor1;
  wire [0:0] u_csamul_cla32_fa27_21_or0;
  wire [0:0] u_csamul_cla32_and28_21;
  wire [0:0] u_csamul_cla32_fa28_21_xor1;
  wire [0:0] u_csamul_cla32_fa28_21_or0;
  wire [0:0] u_csamul_cla32_and29_21;
  wire [0:0] u_csamul_cla32_fa29_21_xor1;
  wire [0:0] u_csamul_cla32_fa29_21_or0;
  wire [0:0] u_csamul_cla32_and30_21;
  wire [0:0] u_csamul_cla32_fa30_21_xor1;
  wire [0:0] u_csamul_cla32_fa30_21_or0;
  wire [0:0] u_csamul_cla32_and31_21;
  wire [0:0] u_csamul_cla32_and0_22;
  wire [0:0] u_csamul_cla32_fa0_22_xor1;
  wire [0:0] u_csamul_cla32_fa0_22_or0;
  wire [0:0] u_csamul_cla32_and1_22;
  wire [0:0] u_csamul_cla32_fa1_22_xor1;
  wire [0:0] u_csamul_cla32_fa1_22_or0;
  wire [0:0] u_csamul_cla32_and2_22;
  wire [0:0] u_csamul_cla32_fa2_22_xor1;
  wire [0:0] u_csamul_cla32_fa2_22_or0;
  wire [0:0] u_csamul_cla32_and3_22;
  wire [0:0] u_csamul_cla32_fa3_22_xor1;
  wire [0:0] u_csamul_cla32_fa3_22_or0;
  wire [0:0] u_csamul_cla32_and4_22;
  wire [0:0] u_csamul_cla32_fa4_22_xor1;
  wire [0:0] u_csamul_cla32_fa4_22_or0;
  wire [0:0] u_csamul_cla32_and5_22;
  wire [0:0] u_csamul_cla32_fa5_22_xor1;
  wire [0:0] u_csamul_cla32_fa5_22_or0;
  wire [0:0] u_csamul_cla32_and6_22;
  wire [0:0] u_csamul_cla32_fa6_22_xor1;
  wire [0:0] u_csamul_cla32_fa6_22_or0;
  wire [0:0] u_csamul_cla32_and7_22;
  wire [0:0] u_csamul_cla32_fa7_22_xor1;
  wire [0:0] u_csamul_cla32_fa7_22_or0;
  wire [0:0] u_csamul_cla32_and8_22;
  wire [0:0] u_csamul_cla32_fa8_22_xor1;
  wire [0:0] u_csamul_cla32_fa8_22_or0;
  wire [0:0] u_csamul_cla32_and9_22;
  wire [0:0] u_csamul_cla32_fa9_22_xor1;
  wire [0:0] u_csamul_cla32_fa9_22_or0;
  wire [0:0] u_csamul_cla32_and10_22;
  wire [0:0] u_csamul_cla32_fa10_22_xor1;
  wire [0:0] u_csamul_cla32_fa10_22_or0;
  wire [0:0] u_csamul_cla32_and11_22;
  wire [0:0] u_csamul_cla32_fa11_22_xor1;
  wire [0:0] u_csamul_cla32_fa11_22_or0;
  wire [0:0] u_csamul_cla32_and12_22;
  wire [0:0] u_csamul_cla32_fa12_22_xor1;
  wire [0:0] u_csamul_cla32_fa12_22_or0;
  wire [0:0] u_csamul_cla32_and13_22;
  wire [0:0] u_csamul_cla32_fa13_22_xor1;
  wire [0:0] u_csamul_cla32_fa13_22_or0;
  wire [0:0] u_csamul_cla32_and14_22;
  wire [0:0] u_csamul_cla32_fa14_22_xor1;
  wire [0:0] u_csamul_cla32_fa14_22_or0;
  wire [0:0] u_csamul_cla32_and15_22;
  wire [0:0] u_csamul_cla32_fa15_22_xor1;
  wire [0:0] u_csamul_cla32_fa15_22_or0;
  wire [0:0] u_csamul_cla32_and16_22;
  wire [0:0] u_csamul_cla32_fa16_22_xor1;
  wire [0:0] u_csamul_cla32_fa16_22_or0;
  wire [0:0] u_csamul_cla32_and17_22;
  wire [0:0] u_csamul_cla32_fa17_22_xor1;
  wire [0:0] u_csamul_cla32_fa17_22_or0;
  wire [0:0] u_csamul_cla32_and18_22;
  wire [0:0] u_csamul_cla32_fa18_22_xor1;
  wire [0:0] u_csamul_cla32_fa18_22_or0;
  wire [0:0] u_csamul_cla32_and19_22;
  wire [0:0] u_csamul_cla32_fa19_22_xor1;
  wire [0:0] u_csamul_cla32_fa19_22_or0;
  wire [0:0] u_csamul_cla32_and20_22;
  wire [0:0] u_csamul_cla32_fa20_22_xor1;
  wire [0:0] u_csamul_cla32_fa20_22_or0;
  wire [0:0] u_csamul_cla32_and21_22;
  wire [0:0] u_csamul_cla32_fa21_22_xor1;
  wire [0:0] u_csamul_cla32_fa21_22_or0;
  wire [0:0] u_csamul_cla32_and22_22;
  wire [0:0] u_csamul_cla32_fa22_22_xor1;
  wire [0:0] u_csamul_cla32_fa22_22_or0;
  wire [0:0] u_csamul_cla32_and23_22;
  wire [0:0] u_csamul_cla32_fa23_22_xor1;
  wire [0:0] u_csamul_cla32_fa23_22_or0;
  wire [0:0] u_csamul_cla32_and24_22;
  wire [0:0] u_csamul_cla32_fa24_22_xor1;
  wire [0:0] u_csamul_cla32_fa24_22_or0;
  wire [0:0] u_csamul_cla32_and25_22;
  wire [0:0] u_csamul_cla32_fa25_22_xor1;
  wire [0:0] u_csamul_cla32_fa25_22_or0;
  wire [0:0] u_csamul_cla32_and26_22;
  wire [0:0] u_csamul_cla32_fa26_22_xor1;
  wire [0:0] u_csamul_cla32_fa26_22_or0;
  wire [0:0] u_csamul_cla32_and27_22;
  wire [0:0] u_csamul_cla32_fa27_22_xor1;
  wire [0:0] u_csamul_cla32_fa27_22_or0;
  wire [0:0] u_csamul_cla32_and28_22;
  wire [0:0] u_csamul_cla32_fa28_22_xor1;
  wire [0:0] u_csamul_cla32_fa28_22_or0;
  wire [0:0] u_csamul_cla32_and29_22;
  wire [0:0] u_csamul_cla32_fa29_22_xor1;
  wire [0:0] u_csamul_cla32_fa29_22_or0;
  wire [0:0] u_csamul_cla32_and30_22;
  wire [0:0] u_csamul_cla32_fa30_22_xor1;
  wire [0:0] u_csamul_cla32_fa30_22_or0;
  wire [0:0] u_csamul_cla32_and31_22;
  wire [0:0] u_csamul_cla32_and0_23;
  wire [0:0] u_csamul_cla32_fa0_23_xor1;
  wire [0:0] u_csamul_cla32_fa0_23_or0;
  wire [0:0] u_csamul_cla32_and1_23;
  wire [0:0] u_csamul_cla32_fa1_23_xor1;
  wire [0:0] u_csamul_cla32_fa1_23_or0;
  wire [0:0] u_csamul_cla32_and2_23;
  wire [0:0] u_csamul_cla32_fa2_23_xor1;
  wire [0:0] u_csamul_cla32_fa2_23_or0;
  wire [0:0] u_csamul_cla32_and3_23;
  wire [0:0] u_csamul_cla32_fa3_23_xor1;
  wire [0:0] u_csamul_cla32_fa3_23_or0;
  wire [0:0] u_csamul_cla32_and4_23;
  wire [0:0] u_csamul_cla32_fa4_23_xor1;
  wire [0:0] u_csamul_cla32_fa4_23_or0;
  wire [0:0] u_csamul_cla32_and5_23;
  wire [0:0] u_csamul_cla32_fa5_23_xor1;
  wire [0:0] u_csamul_cla32_fa5_23_or0;
  wire [0:0] u_csamul_cla32_and6_23;
  wire [0:0] u_csamul_cla32_fa6_23_xor1;
  wire [0:0] u_csamul_cla32_fa6_23_or0;
  wire [0:0] u_csamul_cla32_and7_23;
  wire [0:0] u_csamul_cla32_fa7_23_xor1;
  wire [0:0] u_csamul_cla32_fa7_23_or0;
  wire [0:0] u_csamul_cla32_and8_23;
  wire [0:0] u_csamul_cla32_fa8_23_xor1;
  wire [0:0] u_csamul_cla32_fa8_23_or0;
  wire [0:0] u_csamul_cla32_and9_23;
  wire [0:0] u_csamul_cla32_fa9_23_xor1;
  wire [0:0] u_csamul_cla32_fa9_23_or0;
  wire [0:0] u_csamul_cla32_and10_23;
  wire [0:0] u_csamul_cla32_fa10_23_xor1;
  wire [0:0] u_csamul_cla32_fa10_23_or0;
  wire [0:0] u_csamul_cla32_and11_23;
  wire [0:0] u_csamul_cla32_fa11_23_xor1;
  wire [0:0] u_csamul_cla32_fa11_23_or0;
  wire [0:0] u_csamul_cla32_and12_23;
  wire [0:0] u_csamul_cla32_fa12_23_xor1;
  wire [0:0] u_csamul_cla32_fa12_23_or0;
  wire [0:0] u_csamul_cla32_and13_23;
  wire [0:0] u_csamul_cla32_fa13_23_xor1;
  wire [0:0] u_csamul_cla32_fa13_23_or0;
  wire [0:0] u_csamul_cla32_and14_23;
  wire [0:0] u_csamul_cla32_fa14_23_xor1;
  wire [0:0] u_csamul_cla32_fa14_23_or0;
  wire [0:0] u_csamul_cla32_and15_23;
  wire [0:0] u_csamul_cla32_fa15_23_xor1;
  wire [0:0] u_csamul_cla32_fa15_23_or0;
  wire [0:0] u_csamul_cla32_and16_23;
  wire [0:0] u_csamul_cla32_fa16_23_xor1;
  wire [0:0] u_csamul_cla32_fa16_23_or0;
  wire [0:0] u_csamul_cla32_and17_23;
  wire [0:0] u_csamul_cla32_fa17_23_xor1;
  wire [0:0] u_csamul_cla32_fa17_23_or0;
  wire [0:0] u_csamul_cla32_and18_23;
  wire [0:0] u_csamul_cla32_fa18_23_xor1;
  wire [0:0] u_csamul_cla32_fa18_23_or0;
  wire [0:0] u_csamul_cla32_and19_23;
  wire [0:0] u_csamul_cla32_fa19_23_xor1;
  wire [0:0] u_csamul_cla32_fa19_23_or0;
  wire [0:0] u_csamul_cla32_and20_23;
  wire [0:0] u_csamul_cla32_fa20_23_xor1;
  wire [0:0] u_csamul_cla32_fa20_23_or0;
  wire [0:0] u_csamul_cla32_and21_23;
  wire [0:0] u_csamul_cla32_fa21_23_xor1;
  wire [0:0] u_csamul_cla32_fa21_23_or0;
  wire [0:0] u_csamul_cla32_and22_23;
  wire [0:0] u_csamul_cla32_fa22_23_xor1;
  wire [0:0] u_csamul_cla32_fa22_23_or0;
  wire [0:0] u_csamul_cla32_and23_23;
  wire [0:0] u_csamul_cla32_fa23_23_xor1;
  wire [0:0] u_csamul_cla32_fa23_23_or0;
  wire [0:0] u_csamul_cla32_and24_23;
  wire [0:0] u_csamul_cla32_fa24_23_xor1;
  wire [0:0] u_csamul_cla32_fa24_23_or0;
  wire [0:0] u_csamul_cla32_and25_23;
  wire [0:0] u_csamul_cla32_fa25_23_xor1;
  wire [0:0] u_csamul_cla32_fa25_23_or0;
  wire [0:0] u_csamul_cla32_and26_23;
  wire [0:0] u_csamul_cla32_fa26_23_xor1;
  wire [0:0] u_csamul_cla32_fa26_23_or0;
  wire [0:0] u_csamul_cla32_and27_23;
  wire [0:0] u_csamul_cla32_fa27_23_xor1;
  wire [0:0] u_csamul_cla32_fa27_23_or0;
  wire [0:0] u_csamul_cla32_and28_23;
  wire [0:0] u_csamul_cla32_fa28_23_xor1;
  wire [0:0] u_csamul_cla32_fa28_23_or0;
  wire [0:0] u_csamul_cla32_and29_23;
  wire [0:0] u_csamul_cla32_fa29_23_xor1;
  wire [0:0] u_csamul_cla32_fa29_23_or0;
  wire [0:0] u_csamul_cla32_and30_23;
  wire [0:0] u_csamul_cla32_fa30_23_xor1;
  wire [0:0] u_csamul_cla32_fa30_23_or0;
  wire [0:0] u_csamul_cla32_and31_23;
  wire [0:0] u_csamul_cla32_and0_24;
  wire [0:0] u_csamul_cla32_fa0_24_xor1;
  wire [0:0] u_csamul_cla32_fa0_24_or0;
  wire [0:0] u_csamul_cla32_and1_24;
  wire [0:0] u_csamul_cla32_fa1_24_xor1;
  wire [0:0] u_csamul_cla32_fa1_24_or0;
  wire [0:0] u_csamul_cla32_and2_24;
  wire [0:0] u_csamul_cla32_fa2_24_xor1;
  wire [0:0] u_csamul_cla32_fa2_24_or0;
  wire [0:0] u_csamul_cla32_and3_24;
  wire [0:0] u_csamul_cla32_fa3_24_xor1;
  wire [0:0] u_csamul_cla32_fa3_24_or0;
  wire [0:0] u_csamul_cla32_and4_24;
  wire [0:0] u_csamul_cla32_fa4_24_xor1;
  wire [0:0] u_csamul_cla32_fa4_24_or0;
  wire [0:0] u_csamul_cla32_and5_24;
  wire [0:0] u_csamul_cla32_fa5_24_xor1;
  wire [0:0] u_csamul_cla32_fa5_24_or0;
  wire [0:0] u_csamul_cla32_and6_24;
  wire [0:0] u_csamul_cla32_fa6_24_xor1;
  wire [0:0] u_csamul_cla32_fa6_24_or0;
  wire [0:0] u_csamul_cla32_and7_24;
  wire [0:0] u_csamul_cla32_fa7_24_xor1;
  wire [0:0] u_csamul_cla32_fa7_24_or0;
  wire [0:0] u_csamul_cla32_and8_24;
  wire [0:0] u_csamul_cla32_fa8_24_xor1;
  wire [0:0] u_csamul_cla32_fa8_24_or0;
  wire [0:0] u_csamul_cla32_and9_24;
  wire [0:0] u_csamul_cla32_fa9_24_xor1;
  wire [0:0] u_csamul_cla32_fa9_24_or0;
  wire [0:0] u_csamul_cla32_and10_24;
  wire [0:0] u_csamul_cla32_fa10_24_xor1;
  wire [0:0] u_csamul_cla32_fa10_24_or0;
  wire [0:0] u_csamul_cla32_and11_24;
  wire [0:0] u_csamul_cla32_fa11_24_xor1;
  wire [0:0] u_csamul_cla32_fa11_24_or0;
  wire [0:0] u_csamul_cla32_and12_24;
  wire [0:0] u_csamul_cla32_fa12_24_xor1;
  wire [0:0] u_csamul_cla32_fa12_24_or0;
  wire [0:0] u_csamul_cla32_and13_24;
  wire [0:0] u_csamul_cla32_fa13_24_xor1;
  wire [0:0] u_csamul_cla32_fa13_24_or0;
  wire [0:0] u_csamul_cla32_and14_24;
  wire [0:0] u_csamul_cla32_fa14_24_xor1;
  wire [0:0] u_csamul_cla32_fa14_24_or0;
  wire [0:0] u_csamul_cla32_and15_24;
  wire [0:0] u_csamul_cla32_fa15_24_xor1;
  wire [0:0] u_csamul_cla32_fa15_24_or0;
  wire [0:0] u_csamul_cla32_and16_24;
  wire [0:0] u_csamul_cla32_fa16_24_xor1;
  wire [0:0] u_csamul_cla32_fa16_24_or0;
  wire [0:0] u_csamul_cla32_and17_24;
  wire [0:0] u_csamul_cla32_fa17_24_xor1;
  wire [0:0] u_csamul_cla32_fa17_24_or0;
  wire [0:0] u_csamul_cla32_and18_24;
  wire [0:0] u_csamul_cla32_fa18_24_xor1;
  wire [0:0] u_csamul_cla32_fa18_24_or0;
  wire [0:0] u_csamul_cla32_and19_24;
  wire [0:0] u_csamul_cla32_fa19_24_xor1;
  wire [0:0] u_csamul_cla32_fa19_24_or0;
  wire [0:0] u_csamul_cla32_and20_24;
  wire [0:0] u_csamul_cla32_fa20_24_xor1;
  wire [0:0] u_csamul_cla32_fa20_24_or0;
  wire [0:0] u_csamul_cla32_and21_24;
  wire [0:0] u_csamul_cla32_fa21_24_xor1;
  wire [0:0] u_csamul_cla32_fa21_24_or0;
  wire [0:0] u_csamul_cla32_and22_24;
  wire [0:0] u_csamul_cla32_fa22_24_xor1;
  wire [0:0] u_csamul_cla32_fa22_24_or0;
  wire [0:0] u_csamul_cla32_and23_24;
  wire [0:0] u_csamul_cla32_fa23_24_xor1;
  wire [0:0] u_csamul_cla32_fa23_24_or0;
  wire [0:0] u_csamul_cla32_and24_24;
  wire [0:0] u_csamul_cla32_fa24_24_xor1;
  wire [0:0] u_csamul_cla32_fa24_24_or0;
  wire [0:0] u_csamul_cla32_and25_24;
  wire [0:0] u_csamul_cla32_fa25_24_xor1;
  wire [0:0] u_csamul_cla32_fa25_24_or0;
  wire [0:0] u_csamul_cla32_and26_24;
  wire [0:0] u_csamul_cla32_fa26_24_xor1;
  wire [0:0] u_csamul_cla32_fa26_24_or0;
  wire [0:0] u_csamul_cla32_and27_24;
  wire [0:0] u_csamul_cla32_fa27_24_xor1;
  wire [0:0] u_csamul_cla32_fa27_24_or0;
  wire [0:0] u_csamul_cla32_and28_24;
  wire [0:0] u_csamul_cla32_fa28_24_xor1;
  wire [0:0] u_csamul_cla32_fa28_24_or0;
  wire [0:0] u_csamul_cla32_and29_24;
  wire [0:0] u_csamul_cla32_fa29_24_xor1;
  wire [0:0] u_csamul_cla32_fa29_24_or0;
  wire [0:0] u_csamul_cla32_and30_24;
  wire [0:0] u_csamul_cla32_fa30_24_xor1;
  wire [0:0] u_csamul_cla32_fa30_24_or0;
  wire [0:0] u_csamul_cla32_and31_24;
  wire [0:0] u_csamul_cla32_and0_25;
  wire [0:0] u_csamul_cla32_fa0_25_xor1;
  wire [0:0] u_csamul_cla32_fa0_25_or0;
  wire [0:0] u_csamul_cla32_and1_25;
  wire [0:0] u_csamul_cla32_fa1_25_xor1;
  wire [0:0] u_csamul_cla32_fa1_25_or0;
  wire [0:0] u_csamul_cla32_and2_25;
  wire [0:0] u_csamul_cla32_fa2_25_xor1;
  wire [0:0] u_csamul_cla32_fa2_25_or0;
  wire [0:0] u_csamul_cla32_and3_25;
  wire [0:0] u_csamul_cla32_fa3_25_xor1;
  wire [0:0] u_csamul_cla32_fa3_25_or0;
  wire [0:0] u_csamul_cla32_and4_25;
  wire [0:0] u_csamul_cla32_fa4_25_xor1;
  wire [0:0] u_csamul_cla32_fa4_25_or0;
  wire [0:0] u_csamul_cla32_and5_25;
  wire [0:0] u_csamul_cla32_fa5_25_xor1;
  wire [0:0] u_csamul_cla32_fa5_25_or0;
  wire [0:0] u_csamul_cla32_and6_25;
  wire [0:0] u_csamul_cla32_fa6_25_xor1;
  wire [0:0] u_csamul_cla32_fa6_25_or0;
  wire [0:0] u_csamul_cla32_and7_25;
  wire [0:0] u_csamul_cla32_fa7_25_xor1;
  wire [0:0] u_csamul_cla32_fa7_25_or0;
  wire [0:0] u_csamul_cla32_and8_25;
  wire [0:0] u_csamul_cla32_fa8_25_xor1;
  wire [0:0] u_csamul_cla32_fa8_25_or0;
  wire [0:0] u_csamul_cla32_and9_25;
  wire [0:0] u_csamul_cla32_fa9_25_xor1;
  wire [0:0] u_csamul_cla32_fa9_25_or0;
  wire [0:0] u_csamul_cla32_and10_25;
  wire [0:0] u_csamul_cla32_fa10_25_xor1;
  wire [0:0] u_csamul_cla32_fa10_25_or0;
  wire [0:0] u_csamul_cla32_and11_25;
  wire [0:0] u_csamul_cla32_fa11_25_xor1;
  wire [0:0] u_csamul_cla32_fa11_25_or0;
  wire [0:0] u_csamul_cla32_and12_25;
  wire [0:0] u_csamul_cla32_fa12_25_xor1;
  wire [0:0] u_csamul_cla32_fa12_25_or0;
  wire [0:0] u_csamul_cla32_and13_25;
  wire [0:0] u_csamul_cla32_fa13_25_xor1;
  wire [0:0] u_csamul_cla32_fa13_25_or0;
  wire [0:0] u_csamul_cla32_and14_25;
  wire [0:0] u_csamul_cla32_fa14_25_xor1;
  wire [0:0] u_csamul_cla32_fa14_25_or0;
  wire [0:0] u_csamul_cla32_and15_25;
  wire [0:0] u_csamul_cla32_fa15_25_xor1;
  wire [0:0] u_csamul_cla32_fa15_25_or0;
  wire [0:0] u_csamul_cla32_and16_25;
  wire [0:0] u_csamul_cla32_fa16_25_xor1;
  wire [0:0] u_csamul_cla32_fa16_25_or0;
  wire [0:0] u_csamul_cla32_and17_25;
  wire [0:0] u_csamul_cla32_fa17_25_xor1;
  wire [0:0] u_csamul_cla32_fa17_25_or0;
  wire [0:0] u_csamul_cla32_and18_25;
  wire [0:0] u_csamul_cla32_fa18_25_xor1;
  wire [0:0] u_csamul_cla32_fa18_25_or0;
  wire [0:0] u_csamul_cla32_and19_25;
  wire [0:0] u_csamul_cla32_fa19_25_xor1;
  wire [0:0] u_csamul_cla32_fa19_25_or0;
  wire [0:0] u_csamul_cla32_and20_25;
  wire [0:0] u_csamul_cla32_fa20_25_xor1;
  wire [0:0] u_csamul_cla32_fa20_25_or0;
  wire [0:0] u_csamul_cla32_and21_25;
  wire [0:0] u_csamul_cla32_fa21_25_xor1;
  wire [0:0] u_csamul_cla32_fa21_25_or0;
  wire [0:0] u_csamul_cla32_and22_25;
  wire [0:0] u_csamul_cla32_fa22_25_xor1;
  wire [0:0] u_csamul_cla32_fa22_25_or0;
  wire [0:0] u_csamul_cla32_and23_25;
  wire [0:0] u_csamul_cla32_fa23_25_xor1;
  wire [0:0] u_csamul_cla32_fa23_25_or0;
  wire [0:0] u_csamul_cla32_and24_25;
  wire [0:0] u_csamul_cla32_fa24_25_xor1;
  wire [0:0] u_csamul_cla32_fa24_25_or0;
  wire [0:0] u_csamul_cla32_and25_25;
  wire [0:0] u_csamul_cla32_fa25_25_xor1;
  wire [0:0] u_csamul_cla32_fa25_25_or0;
  wire [0:0] u_csamul_cla32_and26_25;
  wire [0:0] u_csamul_cla32_fa26_25_xor1;
  wire [0:0] u_csamul_cla32_fa26_25_or0;
  wire [0:0] u_csamul_cla32_and27_25;
  wire [0:0] u_csamul_cla32_fa27_25_xor1;
  wire [0:0] u_csamul_cla32_fa27_25_or0;
  wire [0:0] u_csamul_cla32_and28_25;
  wire [0:0] u_csamul_cla32_fa28_25_xor1;
  wire [0:0] u_csamul_cla32_fa28_25_or0;
  wire [0:0] u_csamul_cla32_and29_25;
  wire [0:0] u_csamul_cla32_fa29_25_xor1;
  wire [0:0] u_csamul_cla32_fa29_25_or0;
  wire [0:0] u_csamul_cla32_and30_25;
  wire [0:0] u_csamul_cla32_fa30_25_xor1;
  wire [0:0] u_csamul_cla32_fa30_25_or0;
  wire [0:0] u_csamul_cla32_and31_25;
  wire [0:0] u_csamul_cla32_and0_26;
  wire [0:0] u_csamul_cla32_fa0_26_xor1;
  wire [0:0] u_csamul_cla32_fa0_26_or0;
  wire [0:0] u_csamul_cla32_and1_26;
  wire [0:0] u_csamul_cla32_fa1_26_xor1;
  wire [0:0] u_csamul_cla32_fa1_26_or0;
  wire [0:0] u_csamul_cla32_and2_26;
  wire [0:0] u_csamul_cla32_fa2_26_xor1;
  wire [0:0] u_csamul_cla32_fa2_26_or0;
  wire [0:0] u_csamul_cla32_and3_26;
  wire [0:0] u_csamul_cla32_fa3_26_xor1;
  wire [0:0] u_csamul_cla32_fa3_26_or0;
  wire [0:0] u_csamul_cla32_and4_26;
  wire [0:0] u_csamul_cla32_fa4_26_xor1;
  wire [0:0] u_csamul_cla32_fa4_26_or0;
  wire [0:0] u_csamul_cla32_and5_26;
  wire [0:0] u_csamul_cla32_fa5_26_xor1;
  wire [0:0] u_csamul_cla32_fa5_26_or0;
  wire [0:0] u_csamul_cla32_and6_26;
  wire [0:0] u_csamul_cla32_fa6_26_xor1;
  wire [0:0] u_csamul_cla32_fa6_26_or0;
  wire [0:0] u_csamul_cla32_and7_26;
  wire [0:0] u_csamul_cla32_fa7_26_xor1;
  wire [0:0] u_csamul_cla32_fa7_26_or0;
  wire [0:0] u_csamul_cla32_and8_26;
  wire [0:0] u_csamul_cla32_fa8_26_xor1;
  wire [0:0] u_csamul_cla32_fa8_26_or0;
  wire [0:0] u_csamul_cla32_and9_26;
  wire [0:0] u_csamul_cla32_fa9_26_xor1;
  wire [0:0] u_csamul_cla32_fa9_26_or0;
  wire [0:0] u_csamul_cla32_and10_26;
  wire [0:0] u_csamul_cla32_fa10_26_xor1;
  wire [0:0] u_csamul_cla32_fa10_26_or0;
  wire [0:0] u_csamul_cla32_and11_26;
  wire [0:0] u_csamul_cla32_fa11_26_xor1;
  wire [0:0] u_csamul_cla32_fa11_26_or0;
  wire [0:0] u_csamul_cla32_and12_26;
  wire [0:0] u_csamul_cla32_fa12_26_xor1;
  wire [0:0] u_csamul_cla32_fa12_26_or0;
  wire [0:0] u_csamul_cla32_and13_26;
  wire [0:0] u_csamul_cla32_fa13_26_xor1;
  wire [0:0] u_csamul_cla32_fa13_26_or0;
  wire [0:0] u_csamul_cla32_and14_26;
  wire [0:0] u_csamul_cla32_fa14_26_xor1;
  wire [0:0] u_csamul_cla32_fa14_26_or0;
  wire [0:0] u_csamul_cla32_and15_26;
  wire [0:0] u_csamul_cla32_fa15_26_xor1;
  wire [0:0] u_csamul_cla32_fa15_26_or0;
  wire [0:0] u_csamul_cla32_and16_26;
  wire [0:0] u_csamul_cla32_fa16_26_xor1;
  wire [0:0] u_csamul_cla32_fa16_26_or0;
  wire [0:0] u_csamul_cla32_and17_26;
  wire [0:0] u_csamul_cla32_fa17_26_xor1;
  wire [0:0] u_csamul_cla32_fa17_26_or0;
  wire [0:0] u_csamul_cla32_and18_26;
  wire [0:0] u_csamul_cla32_fa18_26_xor1;
  wire [0:0] u_csamul_cla32_fa18_26_or0;
  wire [0:0] u_csamul_cla32_and19_26;
  wire [0:0] u_csamul_cla32_fa19_26_xor1;
  wire [0:0] u_csamul_cla32_fa19_26_or0;
  wire [0:0] u_csamul_cla32_and20_26;
  wire [0:0] u_csamul_cla32_fa20_26_xor1;
  wire [0:0] u_csamul_cla32_fa20_26_or0;
  wire [0:0] u_csamul_cla32_and21_26;
  wire [0:0] u_csamul_cla32_fa21_26_xor1;
  wire [0:0] u_csamul_cla32_fa21_26_or0;
  wire [0:0] u_csamul_cla32_and22_26;
  wire [0:0] u_csamul_cla32_fa22_26_xor1;
  wire [0:0] u_csamul_cla32_fa22_26_or0;
  wire [0:0] u_csamul_cla32_and23_26;
  wire [0:0] u_csamul_cla32_fa23_26_xor1;
  wire [0:0] u_csamul_cla32_fa23_26_or0;
  wire [0:0] u_csamul_cla32_and24_26;
  wire [0:0] u_csamul_cla32_fa24_26_xor1;
  wire [0:0] u_csamul_cla32_fa24_26_or0;
  wire [0:0] u_csamul_cla32_and25_26;
  wire [0:0] u_csamul_cla32_fa25_26_xor1;
  wire [0:0] u_csamul_cla32_fa25_26_or0;
  wire [0:0] u_csamul_cla32_and26_26;
  wire [0:0] u_csamul_cla32_fa26_26_xor1;
  wire [0:0] u_csamul_cla32_fa26_26_or0;
  wire [0:0] u_csamul_cla32_and27_26;
  wire [0:0] u_csamul_cla32_fa27_26_xor1;
  wire [0:0] u_csamul_cla32_fa27_26_or0;
  wire [0:0] u_csamul_cla32_and28_26;
  wire [0:0] u_csamul_cla32_fa28_26_xor1;
  wire [0:0] u_csamul_cla32_fa28_26_or0;
  wire [0:0] u_csamul_cla32_and29_26;
  wire [0:0] u_csamul_cla32_fa29_26_xor1;
  wire [0:0] u_csamul_cla32_fa29_26_or0;
  wire [0:0] u_csamul_cla32_and30_26;
  wire [0:0] u_csamul_cla32_fa30_26_xor1;
  wire [0:0] u_csamul_cla32_fa30_26_or0;
  wire [0:0] u_csamul_cla32_and31_26;
  wire [0:0] u_csamul_cla32_and0_27;
  wire [0:0] u_csamul_cla32_fa0_27_xor1;
  wire [0:0] u_csamul_cla32_fa0_27_or0;
  wire [0:0] u_csamul_cla32_and1_27;
  wire [0:0] u_csamul_cla32_fa1_27_xor1;
  wire [0:0] u_csamul_cla32_fa1_27_or0;
  wire [0:0] u_csamul_cla32_and2_27;
  wire [0:0] u_csamul_cla32_fa2_27_xor1;
  wire [0:0] u_csamul_cla32_fa2_27_or0;
  wire [0:0] u_csamul_cla32_and3_27;
  wire [0:0] u_csamul_cla32_fa3_27_xor1;
  wire [0:0] u_csamul_cla32_fa3_27_or0;
  wire [0:0] u_csamul_cla32_and4_27;
  wire [0:0] u_csamul_cla32_fa4_27_xor1;
  wire [0:0] u_csamul_cla32_fa4_27_or0;
  wire [0:0] u_csamul_cla32_and5_27;
  wire [0:0] u_csamul_cla32_fa5_27_xor1;
  wire [0:0] u_csamul_cla32_fa5_27_or0;
  wire [0:0] u_csamul_cla32_and6_27;
  wire [0:0] u_csamul_cla32_fa6_27_xor1;
  wire [0:0] u_csamul_cla32_fa6_27_or0;
  wire [0:0] u_csamul_cla32_and7_27;
  wire [0:0] u_csamul_cla32_fa7_27_xor1;
  wire [0:0] u_csamul_cla32_fa7_27_or0;
  wire [0:0] u_csamul_cla32_and8_27;
  wire [0:0] u_csamul_cla32_fa8_27_xor1;
  wire [0:0] u_csamul_cla32_fa8_27_or0;
  wire [0:0] u_csamul_cla32_and9_27;
  wire [0:0] u_csamul_cla32_fa9_27_xor1;
  wire [0:0] u_csamul_cla32_fa9_27_or0;
  wire [0:0] u_csamul_cla32_and10_27;
  wire [0:0] u_csamul_cla32_fa10_27_xor1;
  wire [0:0] u_csamul_cla32_fa10_27_or0;
  wire [0:0] u_csamul_cla32_and11_27;
  wire [0:0] u_csamul_cla32_fa11_27_xor1;
  wire [0:0] u_csamul_cla32_fa11_27_or0;
  wire [0:0] u_csamul_cla32_and12_27;
  wire [0:0] u_csamul_cla32_fa12_27_xor1;
  wire [0:0] u_csamul_cla32_fa12_27_or0;
  wire [0:0] u_csamul_cla32_and13_27;
  wire [0:0] u_csamul_cla32_fa13_27_xor1;
  wire [0:0] u_csamul_cla32_fa13_27_or0;
  wire [0:0] u_csamul_cla32_and14_27;
  wire [0:0] u_csamul_cla32_fa14_27_xor1;
  wire [0:0] u_csamul_cla32_fa14_27_or0;
  wire [0:0] u_csamul_cla32_and15_27;
  wire [0:0] u_csamul_cla32_fa15_27_xor1;
  wire [0:0] u_csamul_cla32_fa15_27_or0;
  wire [0:0] u_csamul_cla32_and16_27;
  wire [0:0] u_csamul_cla32_fa16_27_xor1;
  wire [0:0] u_csamul_cla32_fa16_27_or0;
  wire [0:0] u_csamul_cla32_and17_27;
  wire [0:0] u_csamul_cla32_fa17_27_xor1;
  wire [0:0] u_csamul_cla32_fa17_27_or0;
  wire [0:0] u_csamul_cla32_and18_27;
  wire [0:0] u_csamul_cla32_fa18_27_xor1;
  wire [0:0] u_csamul_cla32_fa18_27_or0;
  wire [0:0] u_csamul_cla32_and19_27;
  wire [0:0] u_csamul_cla32_fa19_27_xor1;
  wire [0:0] u_csamul_cla32_fa19_27_or0;
  wire [0:0] u_csamul_cla32_and20_27;
  wire [0:0] u_csamul_cla32_fa20_27_xor1;
  wire [0:0] u_csamul_cla32_fa20_27_or0;
  wire [0:0] u_csamul_cla32_and21_27;
  wire [0:0] u_csamul_cla32_fa21_27_xor1;
  wire [0:0] u_csamul_cla32_fa21_27_or0;
  wire [0:0] u_csamul_cla32_and22_27;
  wire [0:0] u_csamul_cla32_fa22_27_xor1;
  wire [0:0] u_csamul_cla32_fa22_27_or0;
  wire [0:0] u_csamul_cla32_and23_27;
  wire [0:0] u_csamul_cla32_fa23_27_xor1;
  wire [0:0] u_csamul_cla32_fa23_27_or0;
  wire [0:0] u_csamul_cla32_and24_27;
  wire [0:0] u_csamul_cla32_fa24_27_xor1;
  wire [0:0] u_csamul_cla32_fa24_27_or0;
  wire [0:0] u_csamul_cla32_and25_27;
  wire [0:0] u_csamul_cla32_fa25_27_xor1;
  wire [0:0] u_csamul_cla32_fa25_27_or0;
  wire [0:0] u_csamul_cla32_and26_27;
  wire [0:0] u_csamul_cla32_fa26_27_xor1;
  wire [0:0] u_csamul_cla32_fa26_27_or0;
  wire [0:0] u_csamul_cla32_and27_27;
  wire [0:0] u_csamul_cla32_fa27_27_xor1;
  wire [0:0] u_csamul_cla32_fa27_27_or0;
  wire [0:0] u_csamul_cla32_and28_27;
  wire [0:0] u_csamul_cla32_fa28_27_xor1;
  wire [0:0] u_csamul_cla32_fa28_27_or0;
  wire [0:0] u_csamul_cla32_and29_27;
  wire [0:0] u_csamul_cla32_fa29_27_xor1;
  wire [0:0] u_csamul_cla32_fa29_27_or0;
  wire [0:0] u_csamul_cla32_and30_27;
  wire [0:0] u_csamul_cla32_fa30_27_xor1;
  wire [0:0] u_csamul_cla32_fa30_27_or0;
  wire [0:0] u_csamul_cla32_and31_27;
  wire [0:0] u_csamul_cla32_and0_28;
  wire [0:0] u_csamul_cla32_fa0_28_xor1;
  wire [0:0] u_csamul_cla32_fa0_28_or0;
  wire [0:0] u_csamul_cla32_and1_28;
  wire [0:0] u_csamul_cla32_fa1_28_xor1;
  wire [0:0] u_csamul_cla32_fa1_28_or0;
  wire [0:0] u_csamul_cla32_and2_28;
  wire [0:0] u_csamul_cla32_fa2_28_xor1;
  wire [0:0] u_csamul_cla32_fa2_28_or0;
  wire [0:0] u_csamul_cla32_and3_28;
  wire [0:0] u_csamul_cla32_fa3_28_xor1;
  wire [0:0] u_csamul_cla32_fa3_28_or0;
  wire [0:0] u_csamul_cla32_and4_28;
  wire [0:0] u_csamul_cla32_fa4_28_xor1;
  wire [0:0] u_csamul_cla32_fa4_28_or0;
  wire [0:0] u_csamul_cla32_and5_28;
  wire [0:0] u_csamul_cla32_fa5_28_xor1;
  wire [0:0] u_csamul_cla32_fa5_28_or0;
  wire [0:0] u_csamul_cla32_and6_28;
  wire [0:0] u_csamul_cla32_fa6_28_xor1;
  wire [0:0] u_csamul_cla32_fa6_28_or0;
  wire [0:0] u_csamul_cla32_and7_28;
  wire [0:0] u_csamul_cla32_fa7_28_xor1;
  wire [0:0] u_csamul_cla32_fa7_28_or0;
  wire [0:0] u_csamul_cla32_and8_28;
  wire [0:0] u_csamul_cla32_fa8_28_xor1;
  wire [0:0] u_csamul_cla32_fa8_28_or0;
  wire [0:0] u_csamul_cla32_and9_28;
  wire [0:0] u_csamul_cla32_fa9_28_xor1;
  wire [0:0] u_csamul_cla32_fa9_28_or0;
  wire [0:0] u_csamul_cla32_and10_28;
  wire [0:0] u_csamul_cla32_fa10_28_xor1;
  wire [0:0] u_csamul_cla32_fa10_28_or0;
  wire [0:0] u_csamul_cla32_and11_28;
  wire [0:0] u_csamul_cla32_fa11_28_xor1;
  wire [0:0] u_csamul_cla32_fa11_28_or0;
  wire [0:0] u_csamul_cla32_and12_28;
  wire [0:0] u_csamul_cla32_fa12_28_xor1;
  wire [0:0] u_csamul_cla32_fa12_28_or0;
  wire [0:0] u_csamul_cla32_and13_28;
  wire [0:0] u_csamul_cla32_fa13_28_xor1;
  wire [0:0] u_csamul_cla32_fa13_28_or0;
  wire [0:0] u_csamul_cla32_and14_28;
  wire [0:0] u_csamul_cla32_fa14_28_xor1;
  wire [0:0] u_csamul_cla32_fa14_28_or0;
  wire [0:0] u_csamul_cla32_and15_28;
  wire [0:0] u_csamul_cla32_fa15_28_xor1;
  wire [0:0] u_csamul_cla32_fa15_28_or0;
  wire [0:0] u_csamul_cla32_and16_28;
  wire [0:0] u_csamul_cla32_fa16_28_xor1;
  wire [0:0] u_csamul_cla32_fa16_28_or0;
  wire [0:0] u_csamul_cla32_and17_28;
  wire [0:0] u_csamul_cla32_fa17_28_xor1;
  wire [0:0] u_csamul_cla32_fa17_28_or0;
  wire [0:0] u_csamul_cla32_and18_28;
  wire [0:0] u_csamul_cla32_fa18_28_xor1;
  wire [0:0] u_csamul_cla32_fa18_28_or0;
  wire [0:0] u_csamul_cla32_and19_28;
  wire [0:0] u_csamul_cla32_fa19_28_xor1;
  wire [0:0] u_csamul_cla32_fa19_28_or0;
  wire [0:0] u_csamul_cla32_and20_28;
  wire [0:0] u_csamul_cla32_fa20_28_xor1;
  wire [0:0] u_csamul_cla32_fa20_28_or0;
  wire [0:0] u_csamul_cla32_and21_28;
  wire [0:0] u_csamul_cla32_fa21_28_xor1;
  wire [0:0] u_csamul_cla32_fa21_28_or0;
  wire [0:0] u_csamul_cla32_and22_28;
  wire [0:0] u_csamul_cla32_fa22_28_xor1;
  wire [0:0] u_csamul_cla32_fa22_28_or0;
  wire [0:0] u_csamul_cla32_and23_28;
  wire [0:0] u_csamul_cla32_fa23_28_xor1;
  wire [0:0] u_csamul_cla32_fa23_28_or0;
  wire [0:0] u_csamul_cla32_and24_28;
  wire [0:0] u_csamul_cla32_fa24_28_xor1;
  wire [0:0] u_csamul_cla32_fa24_28_or0;
  wire [0:0] u_csamul_cla32_and25_28;
  wire [0:0] u_csamul_cla32_fa25_28_xor1;
  wire [0:0] u_csamul_cla32_fa25_28_or0;
  wire [0:0] u_csamul_cla32_and26_28;
  wire [0:0] u_csamul_cla32_fa26_28_xor1;
  wire [0:0] u_csamul_cla32_fa26_28_or0;
  wire [0:0] u_csamul_cla32_and27_28;
  wire [0:0] u_csamul_cla32_fa27_28_xor1;
  wire [0:0] u_csamul_cla32_fa27_28_or0;
  wire [0:0] u_csamul_cla32_and28_28;
  wire [0:0] u_csamul_cla32_fa28_28_xor1;
  wire [0:0] u_csamul_cla32_fa28_28_or0;
  wire [0:0] u_csamul_cla32_and29_28;
  wire [0:0] u_csamul_cla32_fa29_28_xor1;
  wire [0:0] u_csamul_cla32_fa29_28_or0;
  wire [0:0] u_csamul_cla32_and30_28;
  wire [0:0] u_csamul_cla32_fa30_28_xor1;
  wire [0:0] u_csamul_cla32_fa30_28_or0;
  wire [0:0] u_csamul_cla32_and31_28;
  wire [0:0] u_csamul_cla32_and0_29;
  wire [0:0] u_csamul_cla32_fa0_29_xor1;
  wire [0:0] u_csamul_cla32_fa0_29_or0;
  wire [0:0] u_csamul_cla32_and1_29;
  wire [0:0] u_csamul_cla32_fa1_29_xor1;
  wire [0:0] u_csamul_cla32_fa1_29_or0;
  wire [0:0] u_csamul_cla32_and2_29;
  wire [0:0] u_csamul_cla32_fa2_29_xor1;
  wire [0:0] u_csamul_cla32_fa2_29_or0;
  wire [0:0] u_csamul_cla32_and3_29;
  wire [0:0] u_csamul_cla32_fa3_29_xor1;
  wire [0:0] u_csamul_cla32_fa3_29_or0;
  wire [0:0] u_csamul_cla32_and4_29;
  wire [0:0] u_csamul_cla32_fa4_29_xor1;
  wire [0:0] u_csamul_cla32_fa4_29_or0;
  wire [0:0] u_csamul_cla32_and5_29;
  wire [0:0] u_csamul_cla32_fa5_29_xor1;
  wire [0:0] u_csamul_cla32_fa5_29_or0;
  wire [0:0] u_csamul_cla32_and6_29;
  wire [0:0] u_csamul_cla32_fa6_29_xor1;
  wire [0:0] u_csamul_cla32_fa6_29_or0;
  wire [0:0] u_csamul_cla32_and7_29;
  wire [0:0] u_csamul_cla32_fa7_29_xor1;
  wire [0:0] u_csamul_cla32_fa7_29_or0;
  wire [0:0] u_csamul_cla32_and8_29;
  wire [0:0] u_csamul_cla32_fa8_29_xor1;
  wire [0:0] u_csamul_cla32_fa8_29_or0;
  wire [0:0] u_csamul_cla32_and9_29;
  wire [0:0] u_csamul_cla32_fa9_29_xor1;
  wire [0:0] u_csamul_cla32_fa9_29_or0;
  wire [0:0] u_csamul_cla32_and10_29;
  wire [0:0] u_csamul_cla32_fa10_29_xor1;
  wire [0:0] u_csamul_cla32_fa10_29_or0;
  wire [0:0] u_csamul_cla32_and11_29;
  wire [0:0] u_csamul_cla32_fa11_29_xor1;
  wire [0:0] u_csamul_cla32_fa11_29_or0;
  wire [0:0] u_csamul_cla32_and12_29;
  wire [0:0] u_csamul_cla32_fa12_29_xor1;
  wire [0:0] u_csamul_cla32_fa12_29_or0;
  wire [0:0] u_csamul_cla32_and13_29;
  wire [0:0] u_csamul_cla32_fa13_29_xor1;
  wire [0:0] u_csamul_cla32_fa13_29_or0;
  wire [0:0] u_csamul_cla32_and14_29;
  wire [0:0] u_csamul_cla32_fa14_29_xor1;
  wire [0:0] u_csamul_cla32_fa14_29_or0;
  wire [0:0] u_csamul_cla32_and15_29;
  wire [0:0] u_csamul_cla32_fa15_29_xor1;
  wire [0:0] u_csamul_cla32_fa15_29_or0;
  wire [0:0] u_csamul_cla32_and16_29;
  wire [0:0] u_csamul_cla32_fa16_29_xor1;
  wire [0:0] u_csamul_cla32_fa16_29_or0;
  wire [0:0] u_csamul_cla32_and17_29;
  wire [0:0] u_csamul_cla32_fa17_29_xor1;
  wire [0:0] u_csamul_cla32_fa17_29_or0;
  wire [0:0] u_csamul_cla32_and18_29;
  wire [0:0] u_csamul_cla32_fa18_29_xor1;
  wire [0:0] u_csamul_cla32_fa18_29_or0;
  wire [0:0] u_csamul_cla32_and19_29;
  wire [0:0] u_csamul_cla32_fa19_29_xor1;
  wire [0:0] u_csamul_cla32_fa19_29_or0;
  wire [0:0] u_csamul_cla32_and20_29;
  wire [0:0] u_csamul_cla32_fa20_29_xor1;
  wire [0:0] u_csamul_cla32_fa20_29_or0;
  wire [0:0] u_csamul_cla32_and21_29;
  wire [0:0] u_csamul_cla32_fa21_29_xor1;
  wire [0:0] u_csamul_cla32_fa21_29_or0;
  wire [0:0] u_csamul_cla32_and22_29;
  wire [0:0] u_csamul_cla32_fa22_29_xor1;
  wire [0:0] u_csamul_cla32_fa22_29_or0;
  wire [0:0] u_csamul_cla32_and23_29;
  wire [0:0] u_csamul_cla32_fa23_29_xor1;
  wire [0:0] u_csamul_cla32_fa23_29_or0;
  wire [0:0] u_csamul_cla32_and24_29;
  wire [0:0] u_csamul_cla32_fa24_29_xor1;
  wire [0:0] u_csamul_cla32_fa24_29_or0;
  wire [0:0] u_csamul_cla32_and25_29;
  wire [0:0] u_csamul_cla32_fa25_29_xor1;
  wire [0:0] u_csamul_cla32_fa25_29_or0;
  wire [0:0] u_csamul_cla32_and26_29;
  wire [0:0] u_csamul_cla32_fa26_29_xor1;
  wire [0:0] u_csamul_cla32_fa26_29_or0;
  wire [0:0] u_csamul_cla32_and27_29;
  wire [0:0] u_csamul_cla32_fa27_29_xor1;
  wire [0:0] u_csamul_cla32_fa27_29_or0;
  wire [0:0] u_csamul_cla32_and28_29;
  wire [0:0] u_csamul_cla32_fa28_29_xor1;
  wire [0:0] u_csamul_cla32_fa28_29_or0;
  wire [0:0] u_csamul_cla32_and29_29;
  wire [0:0] u_csamul_cla32_fa29_29_xor1;
  wire [0:0] u_csamul_cla32_fa29_29_or0;
  wire [0:0] u_csamul_cla32_and30_29;
  wire [0:0] u_csamul_cla32_fa30_29_xor1;
  wire [0:0] u_csamul_cla32_fa30_29_or0;
  wire [0:0] u_csamul_cla32_and31_29;
  wire [0:0] u_csamul_cla32_and0_30;
  wire [0:0] u_csamul_cla32_fa0_30_xor1;
  wire [0:0] u_csamul_cla32_fa0_30_or0;
  wire [0:0] u_csamul_cla32_and1_30;
  wire [0:0] u_csamul_cla32_fa1_30_xor1;
  wire [0:0] u_csamul_cla32_fa1_30_or0;
  wire [0:0] u_csamul_cla32_and2_30;
  wire [0:0] u_csamul_cla32_fa2_30_xor1;
  wire [0:0] u_csamul_cla32_fa2_30_or0;
  wire [0:0] u_csamul_cla32_and3_30;
  wire [0:0] u_csamul_cla32_fa3_30_xor1;
  wire [0:0] u_csamul_cla32_fa3_30_or0;
  wire [0:0] u_csamul_cla32_and4_30;
  wire [0:0] u_csamul_cla32_fa4_30_xor1;
  wire [0:0] u_csamul_cla32_fa4_30_or0;
  wire [0:0] u_csamul_cla32_and5_30;
  wire [0:0] u_csamul_cla32_fa5_30_xor1;
  wire [0:0] u_csamul_cla32_fa5_30_or0;
  wire [0:0] u_csamul_cla32_and6_30;
  wire [0:0] u_csamul_cla32_fa6_30_xor1;
  wire [0:0] u_csamul_cla32_fa6_30_or0;
  wire [0:0] u_csamul_cla32_and7_30;
  wire [0:0] u_csamul_cla32_fa7_30_xor1;
  wire [0:0] u_csamul_cla32_fa7_30_or0;
  wire [0:0] u_csamul_cla32_and8_30;
  wire [0:0] u_csamul_cla32_fa8_30_xor1;
  wire [0:0] u_csamul_cla32_fa8_30_or0;
  wire [0:0] u_csamul_cla32_and9_30;
  wire [0:0] u_csamul_cla32_fa9_30_xor1;
  wire [0:0] u_csamul_cla32_fa9_30_or0;
  wire [0:0] u_csamul_cla32_and10_30;
  wire [0:0] u_csamul_cla32_fa10_30_xor1;
  wire [0:0] u_csamul_cla32_fa10_30_or0;
  wire [0:0] u_csamul_cla32_and11_30;
  wire [0:0] u_csamul_cla32_fa11_30_xor1;
  wire [0:0] u_csamul_cla32_fa11_30_or0;
  wire [0:0] u_csamul_cla32_and12_30;
  wire [0:0] u_csamul_cla32_fa12_30_xor1;
  wire [0:0] u_csamul_cla32_fa12_30_or0;
  wire [0:0] u_csamul_cla32_and13_30;
  wire [0:0] u_csamul_cla32_fa13_30_xor1;
  wire [0:0] u_csamul_cla32_fa13_30_or0;
  wire [0:0] u_csamul_cla32_and14_30;
  wire [0:0] u_csamul_cla32_fa14_30_xor1;
  wire [0:0] u_csamul_cla32_fa14_30_or0;
  wire [0:0] u_csamul_cla32_and15_30;
  wire [0:0] u_csamul_cla32_fa15_30_xor1;
  wire [0:0] u_csamul_cla32_fa15_30_or0;
  wire [0:0] u_csamul_cla32_and16_30;
  wire [0:0] u_csamul_cla32_fa16_30_xor1;
  wire [0:0] u_csamul_cla32_fa16_30_or0;
  wire [0:0] u_csamul_cla32_and17_30;
  wire [0:0] u_csamul_cla32_fa17_30_xor1;
  wire [0:0] u_csamul_cla32_fa17_30_or0;
  wire [0:0] u_csamul_cla32_and18_30;
  wire [0:0] u_csamul_cla32_fa18_30_xor1;
  wire [0:0] u_csamul_cla32_fa18_30_or0;
  wire [0:0] u_csamul_cla32_and19_30;
  wire [0:0] u_csamul_cla32_fa19_30_xor1;
  wire [0:0] u_csamul_cla32_fa19_30_or0;
  wire [0:0] u_csamul_cla32_and20_30;
  wire [0:0] u_csamul_cla32_fa20_30_xor1;
  wire [0:0] u_csamul_cla32_fa20_30_or0;
  wire [0:0] u_csamul_cla32_and21_30;
  wire [0:0] u_csamul_cla32_fa21_30_xor1;
  wire [0:0] u_csamul_cla32_fa21_30_or0;
  wire [0:0] u_csamul_cla32_and22_30;
  wire [0:0] u_csamul_cla32_fa22_30_xor1;
  wire [0:0] u_csamul_cla32_fa22_30_or0;
  wire [0:0] u_csamul_cla32_and23_30;
  wire [0:0] u_csamul_cla32_fa23_30_xor1;
  wire [0:0] u_csamul_cla32_fa23_30_or0;
  wire [0:0] u_csamul_cla32_and24_30;
  wire [0:0] u_csamul_cla32_fa24_30_xor1;
  wire [0:0] u_csamul_cla32_fa24_30_or0;
  wire [0:0] u_csamul_cla32_and25_30;
  wire [0:0] u_csamul_cla32_fa25_30_xor1;
  wire [0:0] u_csamul_cla32_fa25_30_or0;
  wire [0:0] u_csamul_cla32_and26_30;
  wire [0:0] u_csamul_cla32_fa26_30_xor1;
  wire [0:0] u_csamul_cla32_fa26_30_or0;
  wire [0:0] u_csamul_cla32_and27_30;
  wire [0:0] u_csamul_cla32_fa27_30_xor1;
  wire [0:0] u_csamul_cla32_fa27_30_or0;
  wire [0:0] u_csamul_cla32_and28_30;
  wire [0:0] u_csamul_cla32_fa28_30_xor1;
  wire [0:0] u_csamul_cla32_fa28_30_or0;
  wire [0:0] u_csamul_cla32_and29_30;
  wire [0:0] u_csamul_cla32_fa29_30_xor1;
  wire [0:0] u_csamul_cla32_fa29_30_or0;
  wire [0:0] u_csamul_cla32_and30_30;
  wire [0:0] u_csamul_cla32_fa30_30_xor1;
  wire [0:0] u_csamul_cla32_fa30_30_or0;
  wire [0:0] u_csamul_cla32_and31_30;
  wire [0:0] u_csamul_cla32_and0_31;
  wire [0:0] u_csamul_cla32_fa0_31_xor1;
  wire [0:0] u_csamul_cla32_fa0_31_or0;
  wire [0:0] u_csamul_cla32_and1_31;
  wire [0:0] u_csamul_cla32_fa1_31_xor1;
  wire [0:0] u_csamul_cla32_fa1_31_or0;
  wire [0:0] u_csamul_cla32_and2_31;
  wire [0:0] u_csamul_cla32_fa2_31_xor1;
  wire [0:0] u_csamul_cla32_fa2_31_or0;
  wire [0:0] u_csamul_cla32_and3_31;
  wire [0:0] u_csamul_cla32_fa3_31_xor1;
  wire [0:0] u_csamul_cla32_fa3_31_or0;
  wire [0:0] u_csamul_cla32_and4_31;
  wire [0:0] u_csamul_cla32_fa4_31_xor1;
  wire [0:0] u_csamul_cla32_fa4_31_or0;
  wire [0:0] u_csamul_cla32_and5_31;
  wire [0:0] u_csamul_cla32_fa5_31_xor1;
  wire [0:0] u_csamul_cla32_fa5_31_or0;
  wire [0:0] u_csamul_cla32_and6_31;
  wire [0:0] u_csamul_cla32_fa6_31_xor1;
  wire [0:0] u_csamul_cla32_fa6_31_or0;
  wire [0:0] u_csamul_cla32_and7_31;
  wire [0:0] u_csamul_cla32_fa7_31_xor1;
  wire [0:0] u_csamul_cla32_fa7_31_or0;
  wire [0:0] u_csamul_cla32_and8_31;
  wire [0:0] u_csamul_cla32_fa8_31_xor1;
  wire [0:0] u_csamul_cla32_fa8_31_or0;
  wire [0:0] u_csamul_cla32_and9_31;
  wire [0:0] u_csamul_cla32_fa9_31_xor1;
  wire [0:0] u_csamul_cla32_fa9_31_or0;
  wire [0:0] u_csamul_cla32_and10_31;
  wire [0:0] u_csamul_cla32_fa10_31_xor1;
  wire [0:0] u_csamul_cla32_fa10_31_or0;
  wire [0:0] u_csamul_cla32_and11_31;
  wire [0:0] u_csamul_cla32_fa11_31_xor1;
  wire [0:0] u_csamul_cla32_fa11_31_or0;
  wire [0:0] u_csamul_cla32_and12_31;
  wire [0:0] u_csamul_cla32_fa12_31_xor1;
  wire [0:0] u_csamul_cla32_fa12_31_or0;
  wire [0:0] u_csamul_cla32_and13_31;
  wire [0:0] u_csamul_cla32_fa13_31_xor1;
  wire [0:0] u_csamul_cla32_fa13_31_or0;
  wire [0:0] u_csamul_cla32_and14_31;
  wire [0:0] u_csamul_cla32_fa14_31_xor1;
  wire [0:0] u_csamul_cla32_fa14_31_or0;
  wire [0:0] u_csamul_cla32_and15_31;
  wire [0:0] u_csamul_cla32_fa15_31_xor1;
  wire [0:0] u_csamul_cla32_fa15_31_or0;
  wire [0:0] u_csamul_cla32_and16_31;
  wire [0:0] u_csamul_cla32_fa16_31_xor1;
  wire [0:0] u_csamul_cla32_fa16_31_or0;
  wire [0:0] u_csamul_cla32_and17_31;
  wire [0:0] u_csamul_cla32_fa17_31_xor1;
  wire [0:0] u_csamul_cla32_fa17_31_or0;
  wire [0:0] u_csamul_cla32_and18_31;
  wire [0:0] u_csamul_cla32_fa18_31_xor1;
  wire [0:0] u_csamul_cla32_fa18_31_or0;
  wire [0:0] u_csamul_cla32_and19_31;
  wire [0:0] u_csamul_cla32_fa19_31_xor1;
  wire [0:0] u_csamul_cla32_fa19_31_or0;
  wire [0:0] u_csamul_cla32_and20_31;
  wire [0:0] u_csamul_cla32_fa20_31_xor1;
  wire [0:0] u_csamul_cla32_fa20_31_or0;
  wire [0:0] u_csamul_cla32_and21_31;
  wire [0:0] u_csamul_cla32_fa21_31_xor1;
  wire [0:0] u_csamul_cla32_fa21_31_or0;
  wire [0:0] u_csamul_cla32_and22_31;
  wire [0:0] u_csamul_cla32_fa22_31_xor1;
  wire [0:0] u_csamul_cla32_fa22_31_or0;
  wire [0:0] u_csamul_cla32_and23_31;
  wire [0:0] u_csamul_cla32_fa23_31_xor1;
  wire [0:0] u_csamul_cla32_fa23_31_or0;
  wire [0:0] u_csamul_cla32_and24_31;
  wire [0:0] u_csamul_cla32_fa24_31_xor1;
  wire [0:0] u_csamul_cla32_fa24_31_or0;
  wire [0:0] u_csamul_cla32_and25_31;
  wire [0:0] u_csamul_cla32_fa25_31_xor1;
  wire [0:0] u_csamul_cla32_fa25_31_or0;
  wire [0:0] u_csamul_cla32_and26_31;
  wire [0:0] u_csamul_cla32_fa26_31_xor1;
  wire [0:0] u_csamul_cla32_fa26_31_or0;
  wire [0:0] u_csamul_cla32_and27_31;
  wire [0:0] u_csamul_cla32_fa27_31_xor1;
  wire [0:0] u_csamul_cla32_fa27_31_or0;
  wire [0:0] u_csamul_cla32_and28_31;
  wire [0:0] u_csamul_cla32_fa28_31_xor1;
  wire [0:0] u_csamul_cla32_fa28_31_or0;
  wire [0:0] u_csamul_cla32_and29_31;
  wire [0:0] u_csamul_cla32_fa29_31_xor1;
  wire [0:0] u_csamul_cla32_fa29_31_or0;
  wire [0:0] u_csamul_cla32_and30_31;
  wire [0:0] u_csamul_cla32_fa30_31_xor1;
  wire [0:0] u_csamul_cla32_fa30_31_or0;
  wire [0:0] u_csamul_cla32_and31_31;
  wire [31:0] u_csamul_cla32_u_cla32_a;
  wire [31:0] u_csamul_cla32_u_cla32_b;
  wire [32:0] u_csamul_cla32_u_cla32_out;

  and_gate and_gate_u_csamul_cla32_and0_0(.a(a[0]), .b(b[0]), .out(u_csamul_cla32_and0_0));
  and_gate and_gate_u_csamul_cla32_and1_0(.a(a[1]), .b(b[0]), .out(u_csamul_cla32_and1_0));
  and_gate and_gate_u_csamul_cla32_and2_0(.a(a[2]), .b(b[0]), .out(u_csamul_cla32_and2_0));
  and_gate and_gate_u_csamul_cla32_and3_0(.a(a[3]), .b(b[0]), .out(u_csamul_cla32_and3_0));
  and_gate and_gate_u_csamul_cla32_and4_0(.a(a[4]), .b(b[0]), .out(u_csamul_cla32_and4_0));
  and_gate and_gate_u_csamul_cla32_and5_0(.a(a[5]), .b(b[0]), .out(u_csamul_cla32_and5_0));
  and_gate and_gate_u_csamul_cla32_and6_0(.a(a[6]), .b(b[0]), .out(u_csamul_cla32_and6_0));
  and_gate and_gate_u_csamul_cla32_and7_0(.a(a[7]), .b(b[0]), .out(u_csamul_cla32_and7_0));
  and_gate and_gate_u_csamul_cla32_and8_0(.a(a[8]), .b(b[0]), .out(u_csamul_cla32_and8_0));
  and_gate and_gate_u_csamul_cla32_and9_0(.a(a[9]), .b(b[0]), .out(u_csamul_cla32_and9_0));
  and_gate and_gate_u_csamul_cla32_and10_0(.a(a[10]), .b(b[0]), .out(u_csamul_cla32_and10_0));
  and_gate and_gate_u_csamul_cla32_and11_0(.a(a[11]), .b(b[0]), .out(u_csamul_cla32_and11_0));
  and_gate and_gate_u_csamul_cla32_and12_0(.a(a[12]), .b(b[0]), .out(u_csamul_cla32_and12_0));
  and_gate and_gate_u_csamul_cla32_and13_0(.a(a[13]), .b(b[0]), .out(u_csamul_cla32_and13_0));
  and_gate and_gate_u_csamul_cla32_and14_0(.a(a[14]), .b(b[0]), .out(u_csamul_cla32_and14_0));
  and_gate and_gate_u_csamul_cla32_and15_0(.a(a[15]), .b(b[0]), .out(u_csamul_cla32_and15_0));
  and_gate and_gate_u_csamul_cla32_and16_0(.a(a[16]), .b(b[0]), .out(u_csamul_cla32_and16_0));
  and_gate and_gate_u_csamul_cla32_and17_0(.a(a[17]), .b(b[0]), .out(u_csamul_cla32_and17_0));
  and_gate and_gate_u_csamul_cla32_and18_0(.a(a[18]), .b(b[0]), .out(u_csamul_cla32_and18_0));
  and_gate and_gate_u_csamul_cla32_and19_0(.a(a[19]), .b(b[0]), .out(u_csamul_cla32_and19_0));
  and_gate and_gate_u_csamul_cla32_and20_0(.a(a[20]), .b(b[0]), .out(u_csamul_cla32_and20_0));
  and_gate and_gate_u_csamul_cla32_and21_0(.a(a[21]), .b(b[0]), .out(u_csamul_cla32_and21_0));
  and_gate and_gate_u_csamul_cla32_and22_0(.a(a[22]), .b(b[0]), .out(u_csamul_cla32_and22_0));
  and_gate and_gate_u_csamul_cla32_and23_0(.a(a[23]), .b(b[0]), .out(u_csamul_cla32_and23_0));
  and_gate and_gate_u_csamul_cla32_and24_0(.a(a[24]), .b(b[0]), .out(u_csamul_cla32_and24_0));
  and_gate and_gate_u_csamul_cla32_and25_0(.a(a[25]), .b(b[0]), .out(u_csamul_cla32_and25_0));
  and_gate and_gate_u_csamul_cla32_and26_0(.a(a[26]), .b(b[0]), .out(u_csamul_cla32_and26_0));
  and_gate and_gate_u_csamul_cla32_and27_0(.a(a[27]), .b(b[0]), .out(u_csamul_cla32_and27_0));
  and_gate and_gate_u_csamul_cla32_and28_0(.a(a[28]), .b(b[0]), .out(u_csamul_cla32_and28_0));
  and_gate and_gate_u_csamul_cla32_and29_0(.a(a[29]), .b(b[0]), .out(u_csamul_cla32_and29_0));
  and_gate and_gate_u_csamul_cla32_and30_0(.a(a[30]), .b(b[0]), .out(u_csamul_cla32_and30_0));
  and_gate and_gate_u_csamul_cla32_and31_0(.a(a[31]), .b(b[0]), .out(u_csamul_cla32_and31_0));
  and_gate and_gate_u_csamul_cla32_and0_1(.a(a[0]), .b(b[1]), .out(u_csamul_cla32_and0_1));
  ha ha_u_csamul_cla32_ha0_1_out(.a(u_csamul_cla32_and0_1[0]), .b(u_csamul_cla32_and1_0[0]), .ha_xor0(u_csamul_cla32_ha0_1_xor0), .ha_and0(u_csamul_cla32_ha0_1_and0));
  and_gate and_gate_u_csamul_cla32_and1_1(.a(a[1]), .b(b[1]), .out(u_csamul_cla32_and1_1));
  ha ha_u_csamul_cla32_ha1_1_out(.a(u_csamul_cla32_and1_1[0]), .b(u_csamul_cla32_and2_0[0]), .ha_xor0(u_csamul_cla32_ha1_1_xor0), .ha_and0(u_csamul_cla32_ha1_1_and0));
  and_gate and_gate_u_csamul_cla32_and2_1(.a(a[2]), .b(b[1]), .out(u_csamul_cla32_and2_1));
  ha ha_u_csamul_cla32_ha2_1_out(.a(u_csamul_cla32_and2_1[0]), .b(u_csamul_cla32_and3_0[0]), .ha_xor0(u_csamul_cla32_ha2_1_xor0), .ha_and0(u_csamul_cla32_ha2_1_and0));
  and_gate and_gate_u_csamul_cla32_and3_1(.a(a[3]), .b(b[1]), .out(u_csamul_cla32_and3_1));
  ha ha_u_csamul_cla32_ha3_1_out(.a(u_csamul_cla32_and3_1[0]), .b(u_csamul_cla32_and4_0[0]), .ha_xor0(u_csamul_cla32_ha3_1_xor0), .ha_and0(u_csamul_cla32_ha3_1_and0));
  and_gate and_gate_u_csamul_cla32_and4_1(.a(a[4]), .b(b[1]), .out(u_csamul_cla32_and4_1));
  ha ha_u_csamul_cla32_ha4_1_out(.a(u_csamul_cla32_and4_1[0]), .b(u_csamul_cla32_and5_0[0]), .ha_xor0(u_csamul_cla32_ha4_1_xor0), .ha_and0(u_csamul_cla32_ha4_1_and0));
  and_gate and_gate_u_csamul_cla32_and5_1(.a(a[5]), .b(b[1]), .out(u_csamul_cla32_and5_1));
  ha ha_u_csamul_cla32_ha5_1_out(.a(u_csamul_cla32_and5_1[0]), .b(u_csamul_cla32_and6_0[0]), .ha_xor0(u_csamul_cla32_ha5_1_xor0), .ha_and0(u_csamul_cla32_ha5_1_and0));
  and_gate and_gate_u_csamul_cla32_and6_1(.a(a[6]), .b(b[1]), .out(u_csamul_cla32_and6_1));
  ha ha_u_csamul_cla32_ha6_1_out(.a(u_csamul_cla32_and6_1[0]), .b(u_csamul_cla32_and7_0[0]), .ha_xor0(u_csamul_cla32_ha6_1_xor0), .ha_and0(u_csamul_cla32_ha6_1_and0));
  and_gate and_gate_u_csamul_cla32_and7_1(.a(a[7]), .b(b[1]), .out(u_csamul_cla32_and7_1));
  ha ha_u_csamul_cla32_ha7_1_out(.a(u_csamul_cla32_and7_1[0]), .b(u_csamul_cla32_and8_0[0]), .ha_xor0(u_csamul_cla32_ha7_1_xor0), .ha_and0(u_csamul_cla32_ha7_1_and0));
  and_gate and_gate_u_csamul_cla32_and8_1(.a(a[8]), .b(b[1]), .out(u_csamul_cla32_and8_1));
  ha ha_u_csamul_cla32_ha8_1_out(.a(u_csamul_cla32_and8_1[0]), .b(u_csamul_cla32_and9_0[0]), .ha_xor0(u_csamul_cla32_ha8_1_xor0), .ha_and0(u_csamul_cla32_ha8_1_and0));
  and_gate and_gate_u_csamul_cla32_and9_1(.a(a[9]), .b(b[1]), .out(u_csamul_cla32_and9_1));
  ha ha_u_csamul_cla32_ha9_1_out(.a(u_csamul_cla32_and9_1[0]), .b(u_csamul_cla32_and10_0[0]), .ha_xor0(u_csamul_cla32_ha9_1_xor0), .ha_and0(u_csamul_cla32_ha9_1_and0));
  and_gate and_gate_u_csamul_cla32_and10_1(.a(a[10]), .b(b[1]), .out(u_csamul_cla32_and10_1));
  ha ha_u_csamul_cla32_ha10_1_out(.a(u_csamul_cla32_and10_1[0]), .b(u_csamul_cla32_and11_0[0]), .ha_xor0(u_csamul_cla32_ha10_1_xor0), .ha_and0(u_csamul_cla32_ha10_1_and0));
  and_gate and_gate_u_csamul_cla32_and11_1(.a(a[11]), .b(b[1]), .out(u_csamul_cla32_and11_1));
  ha ha_u_csamul_cla32_ha11_1_out(.a(u_csamul_cla32_and11_1[0]), .b(u_csamul_cla32_and12_0[0]), .ha_xor0(u_csamul_cla32_ha11_1_xor0), .ha_and0(u_csamul_cla32_ha11_1_and0));
  and_gate and_gate_u_csamul_cla32_and12_1(.a(a[12]), .b(b[1]), .out(u_csamul_cla32_and12_1));
  ha ha_u_csamul_cla32_ha12_1_out(.a(u_csamul_cla32_and12_1[0]), .b(u_csamul_cla32_and13_0[0]), .ha_xor0(u_csamul_cla32_ha12_1_xor0), .ha_and0(u_csamul_cla32_ha12_1_and0));
  and_gate and_gate_u_csamul_cla32_and13_1(.a(a[13]), .b(b[1]), .out(u_csamul_cla32_and13_1));
  ha ha_u_csamul_cla32_ha13_1_out(.a(u_csamul_cla32_and13_1[0]), .b(u_csamul_cla32_and14_0[0]), .ha_xor0(u_csamul_cla32_ha13_1_xor0), .ha_and0(u_csamul_cla32_ha13_1_and0));
  and_gate and_gate_u_csamul_cla32_and14_1(.a(a[14]), .b(b[1]), .out(u_csamul_cla32_and14_1));
  ha ha_u_csamul_cla32_ha14_1_out(.a(u_csamul_cla32_and14_1[0]), .b(u_csamul_cla32_and15_0[0]), .ha_xor0(u_csamul_cla32_ha14_1_xor0), .ha_and0(u_csamul_cla32_ha14_1_and0));
  and_gate and_gate_u_csamul_cla32_and15_1(.a(a[15]), .b(b[1]), .out(u_csamul_cla32_and15_1));
  ha ha_u_csamul_cla32_ha15_1_out(.a(u_csamul_cla32_and15_1[0]), .b(u_csamul_cla32_and16_0[0]), .ha_xor0(u_csamul_cla32_ha15_1_xor0), .ha_and0(u_csamul_cla32_ha15_1_and0));
  and_gate and_gate_u_csamul_cla32_and16_1(.a(a[16]), .b(b[1]), .out(u_csamul_cla32_and16_1));
  ha ha_u_csamul_cla32_ha16_1_out(.a(u_csamul_cla32_and16_1[0]), .b(u_csamul_cla32_and17_0[0]), .ha_xor0(u_csamul_cla32_ha16_1_xor0), .ha_and0(u_csamul_cla32_ha16_1_and0));
  and_gate and_gate_u_csamul_cla32_and17_1(.a(a[17]), .b(b[1]), .out(u_csamul_cla32_and17_1));
  ha ha_u_csamul_cla32_ha17_1_out(.a(u_csamul_cla32_and17_1[0]), .b(u_csamul_cla32_and18_0[0]), .ha_xor0(u_csamul_cla32_ha17_1_xor0), .ha_and0(u_csamul_cla32_ha17_1_and0));
  and_gate and_gate_u_csamul_cla32_and18_1(.a(a[18]), .b(b[1]), .out(u_csamul_cla32_and18_1));
  ha ha_u_csamul_cla32_ha18_1_out(.a(u_csamul_cla32_and18_1[0]), .b(u_csamul_cla32_and19_0[0]), .ha_xor0(u_csamul_cla32_ha18_1_xor0), .ha_and0(u_csamul_cla32_ha18_1_and0));
  and_gate and_gate_u_csamul_cla32_and19_1(.a(a[19]), .b(b[1]), .out(u_csamul_cla32_and19_1));
  ha ha_u_csamul_cla32_ha19_1_out(.a(u_csamul_cla32_and19_1[0]), .b(u_csamul_cla32_and20_0[0]), .ha_xor0(u_csamul_cla32_ha19_1_xor0), .ha_and0(u_csamul_cla32_ha19_1_and0));
  and_gate and_gate_u_csamul_cla32_and20_1(.a(a[20]), .b(b[1]), .out(u_csamul_cla32_and20_1));
  ha ha_u_csamul_cla32_ha20_1_out(.a(u_csamul_cla32_and20_1[0]), .b(u_csamul_cla32_and21_0[0]), .ha_xor0(u_csamul_cla32_ha20_1_xor0), .ha_and0(u_csamul_cla32_ha20_1_and0));
  and_gate and_gate_u_csamul_cla32_and21_1(.a(a[21]), .b(b[1]), .out(u_csamul_cla32_and21_1));
  ha ha_u_csamul_cla32_ha21_1_out(.a(u_csamul_cla32_and21_1[0]), .b(u_csamul_cla32_and22_0[0]), .ha_xor0(u_csamul_cla32_ha21_1_xor0), .ha_and0(u_csamul_cla32_ha21_1_and0));
  and_gate and_gate_u_csamul_cla32_and22_1(.a(a[22]), .b(b[1]), .out(u_csamul_cla32_and22_1));
  ha ha_u_csamul_cla32_ha22_1_out(.a(u_csamul_cla32_and22_1[0]), .b(u_csamul_cla32_and23_0[0]), .ha_xor0(u_csamul_cla32_ha22_1_xor0), .ha_and0(u_csamul_cla32_ha22_1_and0));
  and_gate and_gate_u_csamul_cla32_and23_1(.a(a[23]), .b(b[1]), .out(u_csamul_cla32_and23_1));
  ha ha_u_csamul_cla32_ha23_1_out(.a(u_csamul_cla32_and23_1[0]), .b(u_csamul_cla32_and24_0[0]), .ha_xor0(u_csamul_cla32_ha23_1_xor0), .ha_and0(u_csamul_cla32_ha23_1_and0));
  and_gate and_gate_u_csamul_cla32_and24_1(.a(a[24]), .b(b[1]), .out(u_csamul_cla32_and24_1));
  ha ha_u_csamul_cla32_ha24_1_out(.a(u_csamul_cla32_and24_1[0]), .b(u_csamul_cla32_and25_0[0]), .ha_xor0(u_csamul_cla32_ha24_1_xor0), .ha_and0(u_csamul_cla32_ha24_1_and0));
  and_gate and_gate_u_csamul_cla32_and25_1(.a(a[25]), .b(b[1]), .out(u_csamul_cla32_and25_1));
  ha ha_u_csamul_cla32_ha25_1_out(.a(u_csamul_cla32_and25_1[0]), .b(u_csamul_cla32_and26_0[0]), .ha_xor0(u_csamul_cla32_ha25_1_xor0), .ha_and0(u_csamul_cla32_ha25_1_and0));
  and_gate and_gate_u_csamul_cla32_and26_1(.a(a[26]), .b(b[1]), .out(u_csamul_cla32_and26_1));
  ha ha_u_csamul_cla32_ha26_1_out(.a(u_csamul_cla32_and26_1[0]), .b(u_csamul_cla32_and27_0[0]), .ha_xor0(u_csamul_cla32_ha26_1_xor0), .ha_and0(u_csamul_cla32_ha26_1_and0));
  and_gate and_gate_u_csamul_cla32_and27_1(.a(a[27]), .b(b[1]), .out(u_csamul_cla32_and27_1));
  ha ha_u_csamul_cla32_ha27_1_out(.a(u_csamul_cla32_and27_1[0]), .b(u_csamul_cla32_and28_0[0]), .ha_xor0(u_csamul_cla32_ha27_1_xor0), .ha_and0(u_csamul_cla32_ha27_1_and0));
  and_gate and_gate_u_csamul_cla32_and28_1(.a(a[28]), .b(b[1]), .out(u_csamul_cla32_and28_1));
  ha ha_u_csamul_cla32_ha28_1_out(.a(u_csamul_cla32_and28_1[0]), .b(u_csamul_cla32_and29_0[0]), .ha_xor0(u_csamul_cla32_ha28_1_xor0), .ha_and0(u_csamul_cla32_ha28_1_and0));
  and_gate and_gate_u_csamul_cla32_and29_1(.a(a[29]), .b(b[1]), .out(u_csamul_cla32_and29_1));
  ha ha_u_csamul_cla32_ha29_1_out(.a(u_csamul_cla32_and29_1[0]), .b(u_csamul_cla32_and30_0[0]), .ha_xor0(u_csamul_cla32_ha29_1_xor0), .ha_and0(u_csamul_cla32_ha29_1_and0));
  and_gate and_gate_u_csamul_cla32_and30_1(.a(a[30]), .b(b[1]), .out(u_csamul_cla32_and30_1));
  ha ha_u_csamul_cla32_ha30_1_out(.a(u_csamul_cla32_and30_1[0]), .b(u_csamul_cla32_and31_0[0]), .ha_xor0(u_csamul_cla32_ha30_1_xor0), .ha_and0(u_csamul_cla32_ha30_1_and0));
  and_gate and_gate_u_csamul_cla32_and31_1(.a(a[31]), .b(b[1]), .out(u_csamul_cla32_and31_1));
  and_gate and_gate_u_csamul_cla32_and0_2(.a(a[0]), .b(b[2]), .out(u_csamul_cla32_and0_2));
  fa fa_u_csamul_cla32_fa0_2_out(.a(u_csamul_cla32_and0_2[0]), .b(u_csamul_cla32_ha1_1_xor0[0]), .cin(u_csamul_cla32_ha0_1_and0[0]), .fa_xor1(u_csamul_cla32_fa0_2_xor1), .fa_or0(u_csamul_cla32_fa0_2_or0));
  and_gate and_gate_u_csamul_cla32_and1_2(.a(a[1]), .b(b[2]), .out(u_csamul_cla32_and1_2));
  fa fa_u_csamul_cla32_fa1_2_out(.a(u_csamul_cla32_and1_2[0]), .b(u_csamul_cla32_ha2_1_xor0[0]), .cin(u_csamul_cla32_ha1_1_and0[0]), .fa_xor1(u_csamul_cla32_fa1_2_xor1), .fa_or0(u_csamul_cla32_fa1_2_or0));
  and_gate and_gate_u_csamul_cla32_and2_2(.a(a[2]), .b(b[2]), .out(u_csamul_cla32_and2_2));
  fa fa_u_csamul_cla32_fa2_2_out(.a(u_csamul_cla32_and2_2[0]), .b(u_csamul_cla32_ha3_1_xor0[0]), .cin(u_csamul_cla32_ha2_1_and0[0]), .fa_xor1(u_csamul_cla32_fa2_2_xor1), .fa_or0(u_csamul_cla32_fa2_2_or0));
  and_gate and_gate_u_csamul_cla32_and3_2(.a(a[3]), .b(b[2]), .out(u_csamul_cla32_and3_2));
  fa fa_u_csamul_cla32_fa3_2_out(.a(u_csamul_cla32_and3_2[0]), .b(u_csamul_cla32_ha4_1_xor0[0]), .cin(u_csamul_cla32_ha3_1_and0[0]), .fa_xor1(u_csamul_cla32_fa3_2_xor1), .fa_or0(u_csamul_cla32_fa3_2_or0));
  and_gate and_gate_u_csamul_cla32_and4_2(.a(a[4]), .b(b[2]), .out(u_csamul_cla32_and4_2));
  fa fa_u_csamul_cla32_fa4_2_out(.a(u_csamul_cla32_and4_2[0]), .b(u_csamul_cla32_ha5_1_xor0[0]), .cin(u_csamul_cla32_ha4_1_and0[0]), .fa_xor1(u_csamul_cla32_fa4_2_xor1), .fa_or0(u_csamul_cla32_fa4_2_or0));
  and_gate and_gate_u_csamul_cla32_and5_2(.a(a[5]), .b(b[2]), .out(u_csamul_cla32_and5_2));
  fa fa_u_csamul_cla32_fa5_2_out(.a(u_csamul_cla32_and5_2[0]), .b(u_csamul_cla32_ha6_1_xor0[0]), .cin(u_csamul_cla32_ha5_1_and0[0]), .fa_xor1(u_csamul_cla32_fa5_2_xor1), .fa_or0(u_csamul_cla32_fa5_2_or0));
  and_gate and_gate_u_csamul_cla32_and6_2(.a(a[6]), .b(b[2]), .out(u_csamul_cla32_and6_2));
  fa fa_u_csamul_cla32_fa6_2_out(.a(u_csamul_cla32_and6_2[0]), .b(u_csamul_cla32_ha7_1_xor0[0]), .cin(u_csamul_cla32_ha6_1_and0[0]), .fa_xor1(u_csamul_cla32_fa6_2_xor1), .fa_or0(u_csamul_cla32_fa6_2_or0));
  and_gate and_gate_u_csamul_cla32_and7_2(.a(a[7]), .b(b[2]), .out(u_csamul_cla32_and7_2));
  fa fa_u_csamul_cla32_fa7_2_out(.a(u_csamul_cla32_and7_2[0]), .b(u_csamul_cla32_ha8_1_xor0[0]), .cin(u_csamul_cla32_ha7_1_and0[0]), .fa_xor1(u_csamul_cla32_fa7_2_xor1), .fa_or0(u_csamul_cla32_fa7_2_or0));
  and_gate and_gate_u_csamul_cla32_and8_2(.a(a[8]), .b(b[2]), .out(u_csamul_cla32_and8_2));
  fa fa_u_csamul_cla32_fa8_2_out(.a(u_csamul_cla32_and8_2[0]), .b(u_csamul_cla32_ha9_1_xor0[0]), .cin(u_csamul_cla32_ha8_1_and0[0]), .fa_xor1(u_csamul_cla32_fa8_2_xor1), .fa_or0(u_csamul_cla32_fa8_2_or0));
  and_gate and_gate_u_csamul_cla32_and9_2(.a(a[9]), .b(b[2]), .out(u_csamul_cla32_and9_2));
  fa fa_u_csamul_cla32_fa9_2_out(.a(u_csamul_cla32_and9_2[0]), .b(u_csamul_cla32_ha10_1_xor0[0]), .cin(u_csamul_cla32_ha9_1_and0[0]), .fa_xor1(u_csamul_cla32_fa9_2_xor1), .fa_or0(u_csamul_cla32_fa9_2_or0));
  and_gate and_gate_u_csamul_cla32_and10_2(.a(a[10]), .b(b[2]), .out(u_csamul_cla32_and10_2));
  fa fa_u_csamul_cla32_fa10_2_out(.a(u_csamul_cla32_and10_2[0]), .b(u_csamul_cla32_ha11_1_xor0[0]), .cin(u_csamul_cla32_ha10_1_and0[0]), .fa_xor1(u_csamul_cla32_fa10_2_xor1), .fa_or0(u_csamul_cla32_fa10_2_or0));
  and_gate and_gate_u_csamul_cla32_and11_2(.a(a[11]), .b(b[2]), .out(u_csamul_cla32_and11_2));
  fa fa_u_csamul_cla32_fa11_2_out(.a(u_csamul_cla32_and11_2[0]), .b(u_csamul_cla32_ha12_1_xor0[0]), .cin(u_csamul_cla32_ha11_1_and0[0]), .fa_xor1(u_csamul_cla32_fa11_2_xor1), .fa_or0(u_csamul_cla32_fa11_2_or0));
  and_gate and_gate_u_csamul_cla32_and12_2(.a(a[12]), .b(b[2]), .out(u_csamul_cla32_and12_2));
  fa fa_u_csamul_cla32_fa12_2_out(.a(u_csamul_cla32_and12_2[0]), .b(u_csamul_cla32_ha13_1_xor0[0]), .cin(u_csamul_cla32_ha12_1_and0[0]), .fa_xor1(u_csamul_cla32_fa12_2_xor1), .fa_or0(u_csamul_cla32_fa12_2_or0));
  and_gate and_gate_u_csamul_cla32_and13_2(.a(a[13]), .b(b[2]), .out(u_csamul_cla32_and13_2));
  fa fa_u_csamul_cla32_fa13_2_out(.a(u_csamul_cla32_and13_2[0]), .b(u_csamul_cla32_ha14_1_xor0[0]), .cin(u_csamul_cla32_ha13_1_and0[0]), .fa_xor1(u_csamul_cla32_fa13_2_xor1), .fa_or0(u_csamul_cla32_fa13_2_or0));
  and_gate and_gate_u_csamul_cla32_and14_2(.a(a[14]), .b(b[2]), .out(u_csamul_cla32_and14_2));
  fa fa_u_csamul_cla32_fa14_2_out(.a(u_csamul_cla32_and14_2[0]), .b(u_csamul_cla32_ha15_1_xor0[0]), .cin(u_csamul_cla32_ha14_1_and0[0]), .fa_xor1(u_csamul_cla32_fa14_2_xor1), .fa_or0(u_csamul_cla32_fa14_2_or0));
  and_gate and_gate_u_csamul_cla32_and15_2(.a(a[15]), .b(b[2]), .out(u_csamul_cla32_and15_2));
  fa fa_u_csamul_cla32_fa15_2_out(.a(u_csamul_cla32_and15_2[0]), .b(u_csamul_cla32_ha16_1_xor0[0]), .cin(u_csamul_cla32_ha15_1_and0[0]), .fa_xor1(u_csamul_cla32_fa15_2_xor1), .fa_or0(u_csamul_cla32_fa15_2_or0));
  and_gate and_gate_u_csamul_cla32_and16_2(.a(a[16]), .b(b[2]), .out(u_csamul_cla32_and16_2));
  fa fa_u_csamul_cla32_fa16_2_out(.a(u_csamul_cla32_and16_2[0]), .b(u_csamul_cla32_ha17_1_xor0[0]), .cin(u_csamul_cla32_ha16_1_and0[0]), .fa_xor1(u_csamul_cla32_fa16_2_xor1), .fa_or0(u_csamul_cla32_fa16_2_or0));
  and_gate and_gate_u_csamul_cla32_and17_2(.a(a[17]), .b(b[2]), .out(u_csamul_cla32_and17_2));
  fa fa_u_csamul_cla32_fa17_2_out(.a(u_csamul_cla32_and17_2[0]), .b(u_csamul_cla32_ha18_1_xor0[0]), .cin(u_csamul_cla32_ha17_1_and0[0]), .fa_xor1(u_csamul_cla32_fa17_2_xor1), .fa_or0(u_csamul_cla32_fa17_2_or0));
  and_gate and_gate_u_csamul_cla32_and18_2(.a(a[18]), .b(b[2]), .out(u_csamul_cla32_and18_2));
  fa fa_u_csamul_cla32_fa18_2_out(.a(u_csamul_cla32_and18_2[0]), .b(u_csamul_cla32_ha19_1_xor0[0]), .cin(u_csamul_cla32_ha18_1_and0[0]), .fa_xor1(u_csamul_cla32_fa18_2_xor1), .fa_or0(u_csamul_cla32_fa18_2_or0));
  and_gate and_gate_u_csamul_cla32_and19_2(.a(a[19]), .b(b[2]), .out(u_csamul_cla32_and19_2));
  fa fa_u_csamul_cla32_fa19_2_out(.a(u_csamul_cla32_and19_2[0]), .b(u_csamul_cla32_ha20_1_xor0[0]), .cin(u_csamul_cla32_ha19_1_and0[0]), .fa_xor1(u_csamul_cla32_fa19_2_xor1), .fa_or0(u_csamul_cla32_fa19_2_or0));
  and_gate and_gate_u_csamul_cla32_and20_2(.a(a[20]), .b(b[2]), .out(u_csamul_cla32_and20_2));
  fa fa_u_csamul_cla32_fa20_2_out(.a(u_csamul_cla32_and20_2[0]), .b(u_csamul_cla32_ha21_1_xor0[0]), .cin(u_csamul_cla32_ha20_1_and0[0]), .fa_xor1(u_csamul_cla32_fa20_2_xor1), .fa_or0(u_csamul_cla32_fa20_2_or0));
  and_gate and_gate_u_csamul_cla32_and21_2(.a(a[21]), .b(b[2]), .out(u_csamul_cla32_and21_2));
  fa fa_u_csamul_cla32_fa21_2_out(.a(u_csamul_cla32_and21_2[0]), .b(u_csamul_cla32_ha22_1_xor0[0]), .cin(u_csamul_cla32_ha21_1_and0[0]), .fa_xor1(u_csamul_cla32_fa21_2_xor1), .fa_or0(u_csamul_cla32_fa21_2_or0));
  and_gate and_gate_u_csamul_cla32_and22_2(.a(a[22]), .b(b[2]), .out(u_csamul_cla32_and22_2));
  fa fa_u_csamul_cla32_fa22_2_out(.a(u_csamul_cla32_and22_2[0]), .b(u_csamul_cla32_ha23_1_xor0[0]), .cin(u_csamul_cla32_ha22_1_and0[0]), .fa_xor1(u_csamul_cla32_fa22_2_xor1), .fa_or0(u_csamul_cla32_fa22_2_or0));
  and_gate and_gate_u_csamul_cla32_and23_2(.a(a[23]), .b(b[2]), .out(u_csamul_cla32_and23_2));
  fa fa_u_csamul_cla32_fa23_2_out(.a(u_csamul_cla32_and23_2[0]), .b(u_csamul_cla32_ha24_1_xor0[0]), .cin(u_csamul_cla32_ha23_1_and0[0]), .fa_xor1(u_csamul_cla32_fa23_2_xor1), .fa_or0(u_csamul_cla32_fa23_2_or0));
  and_gate and_gate_u_csamul_cla32_and24_2(.a(a[24]), .b(b[2]), .out(u_csamul_cla32_and24_2));
  fa fa_u_csamul_cla32_fa24_2_out(.a(u_csamul_cla32_and24_2[0]), .b(u_csamul_cla32_ha25_1_xor0[0]), .cin(u_csamul_cla32_ha24_1_and0[0]), .fa_xor1(u_csamul_cla32_fa24_2_xor1), .fa_or0(u_csamul_cla32_fa24_2_or0));
  and_gate and_gate_u_csamul_cla32_and25_2(.a(a[25]), .b(b[2]), .out(u_csamul_cla32_and25_2));
  fa fa_u_csamul_cla32_fa25_2_out(.a(u_csamul_cla32_and25_2[0]), .b(u_csamul_cla32_ha26_1_xor0[0]), .cin(u_csamul_cla32_ha25_1_and0[0]), .fa_xor1(u_csamul_cla32_fa25_2_xor1), .fa_or0(u_csamul_cla32_fa25_2_or0));
  and_gate and_gate_u_csamul_cla32_and26_2(.a(a[26]), .b(b[2]), .out(u_csamul_cla32_and26_2));
  fa fa_u_csamul_cla32_fa26_2_out(.a(u_csamul_cla32_and26_2[0]), .b(u_csamul_cla32_ha27_1_xor0[0]), .cin(u_csamul_cla32_ha26_1_and0[0]), .fa_xor1(u_csamul_cla32_fa26_2_xor1), .fa_or0(u_csamul_cla32_fa26_2_or0));
  and_gate and_gate_u_csamul_cla32_and27_2(.a(a[27]), .b(b[2]), .out(u_csamul_cla32_and27_2));
  fa fa_u_csamul_cla32_fa27_2_out(.a(u_csamul_cla32_and27_2[0]), .b(u_csamul_cla32_ha28_1_xor0[0]), .cin(u_csamul_cla32_ha27_1_and0[0]), .fa_xor1(u_csamul_cla32_fa27_2_xor1), .fa_or0(u_csamul_cla32_fa27_2_or0));
  and_gate and_gate_u_csamul_cla32_and28_2(.a(a[28]), .b(b[2]), .out(u_csamul_cla32_and28_2));
  fa fa_u_csamul_cla32_fa28_2_out(.a(u_csamul_cla32_and28_2[0]), .b(u_csamul_cla32_ha29_1_xor0[0]), .cin(u_csamul_cla32_ha28_1_and0[0]), .fa_xor1(u_csamul_cla32_fa28_2_xor1), .fa_or0(u_csamul_cla32_fa28_2_or0));
  and_gate and_gate_u_csamul_cla32_and29_2(.a(a[29]), .b(b[2]), .out(u_csamul_cla32_and29_2));
  fa fa_u_csamul_cla32_fa29_2_out(.a(u_csamul_cla32_and29_2[0]), .b(u_csamul_cla32_ha30_1_xor0[0]), .cin(u_csamul_cla32_ha29_1_and0[0]), .fa_xor1(u_csamul_cla32_fa29_2_xor1), .fa_or0(u_csamul_cla32_fa29_2_or0));
  and_gate and_gate_u_csamul_cla32_and30_2(.a(a[30]), .b(b[2]), .out(u_csamul_cla32_and30_2));
  fa fa_u_csamul_cla32_fa30_2_out(.a(u_csamul_cla32_and30_2[0]), .b(u_csamul_cla32_and31_1[0]), .cin(u_csamul_cla32_ha30_1_and0[0]), .fa_xor1(u_csamul_cla32_fa30_2_xor1), .fa_or0(u_csamul_cla32_fa30_2_or0));
  and_gate and_gate_u_csamul_cla32_and31_2(.a(a[31]), .b(b[2]), .out(u_csamul_cla32_and31_2));
  and_gate and_gate_u_csamul_cla32_and0_3(.a(a[0]), .b(b[3]), .out(u_csamul_cla32_and0_3));
  fa fa_u_csamul_cla32_fa0_3_out(.a(u_csamul_cla32_and0_3[0]), .b(u_csamul_cla32_fa1_2_xor1[0]), .cin(u_csamul_cla32_fa0_2_or0[0]), .fa_xor1(u_csamul_cla32_fa0_3_xor1), .fa_or0(u_csamul_cla32_fa0_3_or0));
  and_gate and_gate_u_csamul_cla32_and1_3(.a(a[1]), .b(b[3]), .out(u_csamul_cla32_and1_3));
  fa fa_u_csamul_cla32_fa1_3_out(.a(u_csamul_cla32_and1_3[0]), .b(u_csamul_cla32_fa2_2_xor1[0]), .cin(u_csamul_cla32_fa1_2_or0[0]), .fa_xor1(u_csamul_cla32_fa1_3_xor1), .fa_or0(u_csamul_cla32_fa1_3_or0));
  and_gate and_gate_u_csamul_cla32_and2_3(.a(a[2]), .b(b[3]), .out(u_csamul_cla32_and2_3));
  fa fa_u_csamul_cla32_fa2_3_out(.a(u_csamul_cla32_and2_3[0]), .b(u_csamul_cla32_fa3_2_xor1[0]), .cin(u_csamul_cla32_fa2_2_or0[0]), .fa_xor1(u_csamul_cla32_fa2_3_xor1), .fa_or0(u_csamul_cla32_fa2_3_or0));
  and_gate and_gate_u_csamul_cla32_and3_3(.a(a[3]), .b(b[3]), .out(u_csamul_cla32_and3_3));
  fa fa_u_csamul_cla32_fa3_3_out(.a(u_csamul_cla32_and3_3[0]), .b(u_csamul_cla32_fa4_2_xor1[0]), .cin(u_csamul_cla32_fa3_2_or0[0]), .fa_xor1(u_csamul_cla32_fa3_3_xor1), .fa_or0(u_csamul_cla32_fa3_3_or0));
  and_gate and_gate_u_csamul_cla32_and4_3(.a(a[4]), .b(b[3]), .out(u_csamul_cla32_and4_3));
  fa fa_u_csamul_cla32_fa4_3_out(.a(u_csamul_cla32_and4_3[0]), .b(u_csamul_cla32_fa5_2_xor1[0]), .cin(u_csamul_cla32_fa4_2_or0[0]), .fa_xor1(u_csamul_cla32_fa4_3_xor1), .fa_or0(u_csamul_cla32_fa4_3_or0));
  and_gate and_gate_u_csamul_cla32_and5_3(.a(a[5]), .b(b[3]), .out(u_csamul_cla32_and5_3));
  fa fa_u_csamul_cla32_fa5_3_out(.a(u_csamul_cla32_and5_3[0]), .b(u_csamul_cla32_fa6_2_xor1[0]), .cin(u_csamul_cla32_fa5_2_or0[0]), .fa_xor1(u_csamul_cla32_fa5_3_xor1), .fa_or0(u_csamul_cla32_fa5_3_or0));
  and_gate and_gate_u_csamul_cla32_and6_3(.a(a[6]), .b(b[3]), .out(u_csamul_cla32_and6_3));
  fa fa_u_csamul_cla32_fa6_3_out(.a(u_csamul_cla32_and6_3[0]), .b(u_csamul_cla32_fa7_2_xor1[0]), .cin(u_csamul_cla32_fa6_2_or0[0]), .fa_xor1(u_csamul_cla32_fa6_3_xor1), .fa_or0(u_csamul_cla32_fa6_3_or0));
  and_gate and_gate_u_csamul_cla32_and7_3(.a(a[7]), .b(b[3]), .out(u_csamul_cla32_and7_3));
  fa fa_u_csamul_cla32_fa7_3_out(.a(u_csamul_cla32_and7_3[0]), .b(u_csamul_cla32_fa8_2_xor1[0]), .cin(u_csamul_cla32_fa7_2_or0[0]), .fa_xor1(u_csamul_cla32_fa7_3_xor1), .fa_or0(u_csamul_cla32_fa7_3_or0));
  and_gate and_gate_u_csamul_cla32_and8_3(.a(a[8]), .b(b[3]), .out(u_csamul_cla32_and8_3));
  fa fa_u_csamul_cla32_fa8_3_out(.a(u_csamul_cla32_and8_3[0]), .b(u_csamul_cla32_fa9_2_xor1[0]), .cin(u_csamul_cla32_fa8_2_or0[0]), .fa_xor1(u_csamul_cla32_fa8_3_xor1), .fa_or0(u_csamul_cla32_fa8_3_or0));
  and_gate and_gate_u_csamul_cla32_and9_3(.a(a[9]), .b(b[3]), .out(u_csamul_cla32_and9_3));
  fa fa_u_csamul_cla32_fa9_3_out(.a(u_csamul_cla32_and9_3[0]), .b(u_csamul_cla32_fa10_2_xor1[0]), .cin(u_csamul_cla32_fa9_2_or0[0]), .fa_xor1(u_csamul_cla32_fa9_3_xor1), .fa_or0(u_csamul_cla32_fa9_3_or0));
  and_gate and_gate_u_csamul_cla32_and10_3(.a(a[10]), .b(b[3]), .out(u_csamul_cla32_and10_3));
  fa fa_u_csamul_cla32_fa10_3_out(.a(u_csamul_cla32_and10_3[0]), .b(u_csamul_cla32_fa11_2_xor1[0]), .cin(u_csamul_cla32_fa10_2_or0[0]), .fa_xor1(u_csamul_cla32_fa10_3_xor1), .fa_or0(u_csamul_cla32_fa10_3_or0));
  and_gate and_gate_u_csamul_cla32_and11_3(.a(a[11]), .b(b[3]), .out(u_csamul_cla32_and11_3));
  fa fa_u_csamul_cla32_fa11_3_out(.a(u_csamul_cla32_and11_3[0]), .b(u_csamul_cla32_fa12_2_xor1[0]), .cin(u_csamul_cla32_fa11_2_or0[0]), .fa_xor1(u_csamul_cla32_fa11_3_xor1), .fa_or0(u_csamul_cla32_fa11_3_or0));
  and_gate and_gate_u_csamul_cla32_and12_3(.a(a[12]), .b(b[3]), .out(u_csamul_cla32_and12_3));
  fa fa_u_csamul_cla32_fa12_3_out(.a(u_csamul_cla32_and12_3[0]), .b(u_csamul_cla32_fa13_2_xor1[0]), .cin(u_csamul_cla32_fa12_2_or0[0]), .fa_xor1(u_csamul_cla32_fa12_3_xor1), .fa_or0(u_csamul_cla32_fa12_3_or0));
  and_gate and_gate_u_csamul_cla32_and13_3(.a(a[13]), .b(b[3]), .out(u_csamul_cla32_and13_3));
  fa fa_u_csamul_cla32_fa13_3_out(.a(u_csamul_cla32_and13_3[0]), .b(u_csamul_cla32_fa14_2_xor1[0]), .cin(u_csamul_cla32_fa13_2_or0[0]), .fa_xor1(u_csamul_cla32_fa13_3_xor1), .fa_or0(u_csamul_cla32_fa13_3_or0));
  and_gate and_gate_u_csamul_cla32_and14_3(.a(a[14]), .b(b[3]), .out(u_csamul_cla32_and14_3));
  fa fa_u_csamul_cla32_fa14_3_out(.a(u_csamul_cla32_and14_3[0]), .b(u_csamul_cla32_fa15_2_xor1[0]), .cin(u_csamul_cla32_fa14_2_or0[0]), .fa_xor1(u_csamul_cla32_fa14_3_xor1), .fa_or0(u_csamul_cla32_fa14_3_or0));
  and_gate and_gate_u_csamul_cla32_and15_3(.a(a[15]), .b(b[3]), .out(u_csamul_cla32_and15_3));
  fa fa_u_csamul_cla32_fa15_3_out(.a(u_csamul_cla32_and15_3[0]), .b(u_csamul_cla32_fa16_2_xor1[0]), .cin(u_csamul_cla32_fa15_2_or0[0]), .fa_xor1(u_csamul_cla32_fa15_3_xor1), .fa_or0(u_csamul_cla32_fa15_3_or0));
  and_gate and_gate_u_csamul_cla32_and16_3(.a(a[16]), .b(b[3]), .out(u_csamul_cla32_and16_3));
  fa fa_u_csamul_cla32_fa16_3_out(.a(u_csamul_cla32_and16_3[0]), .b(u_csamul_cla32_fa17_2_xor1[0]), .cin(u_csamul_cla32_fa16_2_or0[0]), .fa_xor1(u_csamul_cla32_fa16_3_xor1), .fa_or0(u_csamul_cla32_fa16_3_or0));
  and_gate and_gate_u_csamul_cla32_and17_3(.a(a[17]), .b(b[3]), .out(u_csamul_cla32_and17_3));
  fa fa_u_csamul_cla32_fa17_3_out(.a(u_csamul_cla32_and17_3[0]), .b(u_csamul_cla32_fa18_2_xor1[0]), .cin(u_csamul_cla32_fa17_2_or0[0]), .fa_xor1(u_csamul_cla32_fa17_3_xor1), .fa_or0(u_csamul_cla32_fa17_3_or0));
  and_gate and_gate_u_csamul_cla32_and18_3(.a(a[18]), .b(b[3]), .out(u_csamul_cla32_and18_3));
  fa fa_u_csamul_cla32_fa18_3_out(.a(u_csamul_cla32_and18_3[0]), .b(u_csamul_cla32_fa19_2_xor1[0]), .cin(u_csamul_cla32_fa18_2_or0[0]), .fa_xor1(u_csamul_cla32_fa18_3_xor1), .fa_or0(u_csamul_cla32_fa18_3_or0));
  and_gate and_gate_u_csamul_cla32_and19_3(.a(a[19]), .b(b[3]), .out(u_csamul_cla32_and19_3));
  fa fa_u_csamul_cla32_fa19_3_out(.a(u_csamul_cla32_and19_3[0]), .b(u_csamul_cla32_fa20_2_xor1[0]), .cin(u_csamul_cla32_fa19_2_or0[0]), .fa_xor1(u_csamul_cla32_fa19_3_xor1), .fa_or0(u_csamul_cla32_fa19_3_or0));
  and_gate and_gate_u_csamul_cla32_and20_3(.a(a[20]), .b(b[3]), .out(u_csamul_cla32_and20_3));
  fa fa_u_csamul_cla32_fa20_3_out(.a(u_csamul_cla32_and20_3[0]), .b(u_csamul_cla32_fa21_2_xor1[0]), .cin(u_csamul_cla32_fa20_2_or0[0]), .fa_xor1(u_csamul_cla32_fa20_3_xor1), .fa_or0(u_csamul_cla32_fa20_3_or0));
  and_gate and_gate_u_csamul_cla32_and21_3(.a(a[21]), .b(b[3]), .out(u_csamul_cla32_and21_3));
  fa fa_u_csamul_cla32_fa21_3_out(.a(u_csamul_cla32_and21_3[0]), .b(u_csamul_cla32_fa22_2_xor1[0]), .cin(u_csamul_cla32_fa21_2_or0[0]), .fa_xor1(u_csamul_cla32_fa21_3_xor1), .fa_or0(u_csamul_cla32_fa21_3_or0));
  and_gate and_gate_u_csamul_cla32_and22_3(.a(a[22]), .b(b[3]), .out(u_csamul_cla32_and22_3));
  fa fa_u_csamul_cla32_fa22_3_out(.a(u_csamul_cla32_and22_3[0]), .b(u_csamul_cla32_fa23_2_xor1[0]), .cin(u_csamul_cla32_fa22_2_or0[0]), .fa_xor1(u_csamul_cla32_fa22_3_xor1), .fa_or0(u_csamul_cla32_fa22_3_or0));
  and_gate and_gate_u_csamul_cla32_and23_3(.a(a[23]), .b(b[3]), .out(u_csamul_cla32_and23_3));
  fa fa_u_csamul_cla32_fa23_3_out(.a(u_csamul_cla32_and23_3[0]), .b(u_csamul_cla32_fa24_2_xor1[0]), .cin(u_csamul_cla32_fa23_2_or0[0]), .fa_xor1(u_csamul_cla32_fa23_3_xor1), .fa_or0(u_csamul_cla32_fa23_3_or0));
  and_gate and_gate_u_csamul_cla32_and24_3(.a(a[24]), .b(b[3]), .out(u_csamul_cla32_and24_3));
  fa fa_u_csamul_cla32_fa24_3_out(.a(u_csamul_cla32_and24_3[0]), .b(u_csamul_cla32_fa25_2_xor1[0]), .cin(u_csamul_cla32_fa24_2_or0[0]), .fa_xor1(u_csamul_cla32_fa24_3_xor1), .fa_or0(u_csamul_cla32_fa24_3_or0));
  and_gate and_gate_u_csamul_cla32_and25_3(.a(a[25]), .b(b[3]), .out(u_csamul_cla32_and25_3));
  fa fa_u_csamul_cla32_fa25_3_out(.a(u_csamul_cla32_and25_3[0]), .b(u_csamul_cla32_fa26_2_xor1[0]), .cin(u_csamul_cla32_fa25_2_or0[0]), .fa_xor1(u_csamul_cla32_fa25_3_xor1), .fa_or0(u_csamul_cla32_fa25_3_or0));
  and_gate and_gate_u_csamul_cla32_and26_3(.a(a[26]), .b(b[3]), .out(u_csamul_cla32_and26_3));
  fa fa_u_csamul_cla32_fa26_3_out(.a(u_csamul_cla32_and26_3[0]), .b(u_csamul_cla32_fa27_2_xor1[0]), .cin(u_csamul_cla32_fa26_2_or0[0]), .fa_xor1(u_csamul_cla32_fa26_3_xor1), .fa_or0(u_csamul_cla32_fa26_3_or0));
  and_gate and_gate_u_csamul_cla32_and27_3(.a(a[27]), .b(b[3]), .out(u_csamul_cla32_and27_3));
  fa fa_u_csamul_cla32_fa27_3_out(.a(u_csamul_cla32_and27_3[0]), .b(u_csamul_cla32_fa28_2_xor1[0]), .cin(u_csamul_cla32_fa27_2_or0[0]), .fa_xor1(u_csamul_cla32_fa27_3_xor1), .fa_or0(u_csamul_cla32_fa27_3_or0));
  and_gate and_gate_u_csamul_cla32_and28_3(.a(a[28]), .b(b[3]), .out(u_csamul_cla32_and28_3));
  fa fa_u_csamul_cla32_fa28_3_out(.a(u_csamul_cla32_and28_3[0]), .b(u_csamul_cla32_fa29_2_xor1[0]), .cin(u_csamul_cla32_fa28_2_or0[0]), .fa_xor1(u_csamul_cla32_fa28_3_xor1), .fa_or0(u_csamul_cla32_fa28_3_or0));
  and_gate and_gate_u_csamul_cla32_and29_3(.a(a[29]), .b(b[3]), .out(u_csamul_cla32_and29_3));
  fa fa_u_csamul_cla32_fa29_3_out(.a(u_csamul_cla32_and29_3[0]), .b(u_csamul_cla32_fa30_2_xor1[0]), .cin(u_csamul_cla32_fa29_2_or0[0]), .fa_xor1(u_csamul_cla32_fa29_3_xor1), .fa_or0(u_csamul_cla32_fa29_3_or0));
  and_gate and_gate_u_csamul_cla32_and30_3(.a(a[30]), .b(b[3]), .out(u_csamul_cla32_and30_3));
  fa fa_u_csamul_cla32_fa30_3_out(.a(u_csamul_cla32_and30_3[0]), .b(u_csamul_cla32_and31_2[0]), .cin(u_csamul_cla32_fa30_2_or0[0]), .fa_xor1(u_csamul_cla32_fa30_3_xor1), .fa_or0(u_csamul_cla32_fa30_3_or0));
  and_gate and_gate_u_csamul_cla32_and31_3(.a(a[31]), .b(b[3]), .out(u_csamul_cla32_and31_3));
  and_gate and_gate_u_csamul_cla32_and0_4(.a(a[0]), .b(b[4]), .out(u_csamul_cla32_and0_4));
  fa fa_u_csamul_cla32_fa0_4_out(.a(u_csamul_cla32_and0_4[0]), .b(u_csamul_cla32_fa1_3_xor1[0]), .cin(u_csamul_cla32_fa0_3_or0[0]), .fa_xor1(u_csamul_cla32_fa0_4_xor1), .fa_or0(u_csamul_cla32_fa0_4_or0));
  and_gate and_gate_u_csamul_cla32_and1_4(.a(a[1]), .b(b[4]), .out(u_csamul_cla32_and1_4));
  fa fa_u_csamul_cla32_fa1_4_out(.a(u_csamul_cla32_and1_4[0]), .b(u_csamul_cla32_fa2_3_xor1[0]), .cin(u_csamul_cla32_fa1_3_or0[0]), .fa_xor1(u_csamul_cla32_fa1_4_xor1), .fa_or0(u_csamul_cla32_fa1_4_or0));
  and_gate and_gate_u_csamul_cla32_and2_4(.a(a[2]), .b(b[4]), .out(u_csamul_cla32_and2_4));
  fa fa_u_csamul_cla32_fa2_4_out(.a(u_csamul_cla32_and2_4[0]), .b(u_csamul_cla32_fa3_3_xor1[0]), .cin(u_csamul_cla32_fa2_3_or0[0]), .fa_xor1(u_csamul_cla32_fa2_4_xor1), .fa_or0(u_csamul_cla32_fa2_4_or0));
  and_gate and_gate_u_csamul_cla32_and3_4(.a(a[3]), .b(b[4]), .out(u_csamul_cla32_and3_4));
  fa fa_u_csamul_cla32_fa3_4_out(.a(u_csamul_cla32_and3_4[0]), .b(u_csamul_cla32_fa4_3_xor1[0]), .cin(u_csamul_cla32_fa3_3_or0[0]), .fa_xor1(u_csamul_cla32_fa3_4_xor1), .fa_or0(u_csamul_cla32_fa3_4_or0));
  and_gate and_gate_u_csamul_cla32_and4_4(.a(a[4]), .b(b[4]), .out(u_csamul_cla32_and4_4));
  fa fa_u_csamul_cla32_fa4_4_out(.a(u_csamul_cla32_and4_4[0]), .b(u_csamul_cla32_fa5_3_xor1[0]), .cin(u_csamul_cla32_fa4_3_or0[0]), .fa_xor1(u_csamul_cla32_fa4_4_xor1), .fa_or0(u_csamul_cla32_fa4_4_or0));
  and_gate and_gate_u_csamul_cla32_and5_4(.a(a[5]), .b(b[4]), .out(u_csamul_cla32_and5_4));
  fa fa_u_csamul_cla32_fa5_4_out(.a(u_csamul_cla32_and5_4[0]), .b(u_csamul_cla32_fa6_3_xor1[0]), .cin(u_csamul_cla32_fa5_3_or0[0]), .fa_xor1(u_csamul_cla32_fa5_4_xor1), .fa_or0(u_csamul_cla32_fa5_4_or0));
  and_gate and_gate_u_csamul_cla32_and6_4(.a(a[6]), .b(b[4]), .out(u_csamul_cla32_and6_4));
  fa fa_u_csamul_cla32_fa6_4_out(.a(u_csamul_cla32_and6_4[0]), .b(u_csamul_cla32_fa7_3_xor1[0]), .cin(u_csamul_cla32_fa6_3_or0[0]), .fa_xor1(u_csamul_cla32_fa6_4_xor1), .fa_or0(u_csamul_cla32_fa6_4_or0));
  and_gate and_gate_u_csamul_cla32_and7_4(.a(a[7]), .b(b[4]), .out(u_csamul_cla32_and7_4));
  fa fa_u_csamul_cla32_fa7_4_out(.a(u_csamul_cla32_and7_4[0]), .b(u_csamul_cla32_fa8_3_xor1[0]), .cin(u_csamul_cla32_fa7_3_or0[0]), .fa_xor1(u_csamul_cla32_fa7_4_xor1), .fa_or0(u_csamul_cla32_fa7_4_or0));
  and_gate and_gate_u_csamul_cla32_and8_4(.a(a[8]), .b(b[4]), .out(u_csamul_cla32_and8_4));
  fa fa_u_csamul_cla32_fa8_4_out(.a(u_csamul_cla32_and8_4[0]), .b(u_csamul_cla32_fa9_3_xor1[0]), .cin(u_csamul_cla32_fa8_3_or0[0]), .fa_xor1(u_csamul_cla32_fa8_4_xor1), .fa_or0(u_csamul_cla32_fa8_4_or0));
  and_gate and_gate_u_csamul_cla32_and9_4(.a(a[9]), .b(b[4]), .out(u_csamul_cla32_and9_4));
  fa fa_u_csamul_cla32_fa9_4_out(.a(u_csamul_cla32_and9_4[0]), .b(u_csamul_cla32_fa10_3_xor1[0]), .cin(u_csamul_cla32_fa9_3_or0[0]), .fa_xor1(u_csamul_cla32_fa9_4_xor1), .fa_or0(u_csamul_cla32_fa9_4_or0));
  and_gate and_gate_u_csamul_cla32_and10_4(.a(a[10]), .b(b[4]), .out(u_csamul_cla32_and10_4));
  fa fa_u_csamul_cla32_fa10_4_out(.a(u_csamul_cla32_and10_4[0]), .b(u_csamul_cla32_fa11_3_xor1[0]), .cin(u_csamul_cla32_fa10_3_or0[0]), .fa_xor1(u_csamul_cla32_fa10_4_xor1), .fa_or0(u_csamul_cla32_fa10_4_or0));
  and_gate and_gate_u_csamul_cla32_and11_4(.a(a[11]), .b(b[4]), .out(u_csamul_cla32_and11_4));
  fa fa_u_csamul_cla32_fa11_4_out(.a(u_csamul_cla32_and11_4[0]), .b(u_csamul_cla32_fa12_3_xor1[0]), .cin(u_csamul_cla32_fa11_3_or0[0]), .fa_xor1(u_csamul_cla32_fa11_4_xor1), .fa_or0(u_csamul_cla32_fa11_4_or0));
  and_gate and_gate_u_csamul_cla32_and12_4(.a(a[12]), .b(b[4]), .out(u_csamul_cla32_and12_4));
  fa fa_u_csamul_cla32_fa12_4_out(.a(u_csamul_cla32_and12_4[0]), .b(u_csamul_cla32_fa13_3_xor1[0]), .cin(u_csamul_cla32_fa12_3_or0[0]), .fa_xor1(u_csamul_cla32_fa12_4_xor1), .fa_or0(u_csamul_cla32_fa12_4_or0));
  and_gate and_gate_u_csamul_cla32_and13_4(.a(a[13]), .b(b[4]), .out(u_csamul_cla32_and13_4));
  fa fa_u_csamul_cla32_fa13_4_out(.a(u_csamul_cla32_and13_4[0]), .b(u_csamul_cla32_fa14_3_xor1[0]), .cin(u_csamul_cla32_fa13_3_or0[0]), .fa_xor1(u_csamul_cla32_fa13_4_xor1), .fa_or0(u_csamul_cla32_fa13_4_or0));
  and_gate and_gate_u_csamul_cla32_and14_4(.a(a[14]), .b(b[4]), .out(u_csamul_cla32_and14_4));
  fa fa_u_csamul_cla32_fa14_4_out(.a(u_csamul_cla32_and14_4[0]), .b(u_csamul_cla32_fa15_3_xor1[0]), .cin(u_csamul_cla32_fa14_3_or0[0]), .fa_xor1(u_csamul_cla32_fa14_4_xor1), .fa_or0(u_csamul_cla32_fa14_4_or0));
  and_gate and_gate_u_csamul_cla32_and15_4(.a(a[15]), .b(b[4]), .out(u_csamul_cla32_and15_4));
  fa fa_u_csamul_cla32_fa15_4_out(.a(u_csamul_cla32_and15_4[0]), .b(u_csamul_cla32_fa16_3_xor1[0]), .cin(u_csamul_cla32_fa15_3_or0[0]), .fa_xor1(u_csamul_cla32_fa15_4_xor1), .fa_or0(u_csamul_cla32_fa15_4_or0));
  and_gate and_gate_u_csamul_cla32_and16_4(.a(a[16]), .b(b[4]), .out(u_csamul_cla32_and16_4));
  fa fa_u_csamul_cla32_fa16_4_out(.a(u_csamul_cla32_and16_4[0]), .b(u_csamul_cla32_fa17_3_xor1[0]), .cin(u_csamul_cla32_fa16_3_or0[0]), .fa_xor1(u_csamul_cla32_fa16_4_xor1), .fa_or0(u_csamul_cla32_fa16_4_or0));
  and_gate and_gate_u_csamul_cla32_and17_4(.a(a[17]), .b(b[4]), .out(u_csamul_cla32_and17_4));
  fa fa_u_csamul_cla32_fa17_4_out(.a(u_csamul_cla32_and17_4[0]), .b(u_csamul_cla32_fa18_3_xor1[0]), .cin(u_csamul_cla32_fa17_3_or0[0]), .fa_xor1(u_csamul_cla32_fa17_4_xor1), .fa_or0(u_csamul_cla32_fa17_4_or0));
  and_gate and_gate_u_csamul_cla32_and18_4(.a(a[18]), .b(b[4]), .out(u_csamul_cla32_and18_4));
  fa fa_u_csamul_cla32_fa18_4_out(.a(u_csamul_cla32_and18_4[0]), .b(u_csamul_cla32_fa19_3_xor1[0]), .cin(u_csamul_cla32_fa18_3_or0[0]), .fa_xor1(u_csamul_cla32_fa18_4_xor1), .fa_or0(u_csamul_cla32_fa18_4_or0));
  and_gate and_gate_u_csamul_cla32_and19_4(.a(a[19]), .b(b[4]), .out(u_csamul_cla32_and19_4));
  fa fa_u_csamul_cla32_fa19_4_out(.a(u_csamul_cla32_and19_4[0]), .b(u_csamul_cla32_fa20_3_xor1[0]), .cin(u_csamul_cla32_fa19_3_or0[0]), .fa_xor1(u_csamul_cla32_fa19_4_xor1), .fa_or0(u_csamul_cla32_fa19_4_or0));
  and_gate and_gate_u_csamul_cla32_and20_4(.a(a[20]), .b(b[4]), .out(u_csamul_cla32_and20_4));
  fa fa_u_csamul_cla32_fa20_4_out(.a(u_csamul_cla32_and20_4[0]), .b(u_csamul_cla32_fa21_3_xor1[0]), .cin(u_csamul_cla32_fa20_3_or0[0]), .fa_xor1(u_csamul_cla32_fa20_4_xor1), .fa_or0(u_csamul_cla32_fa20_4_or0));
  and_gate and_gate_u_csamul_cla32_and21_4(.a(a[21]), .b(b[4]), .out(u_csamul_cla32_and21_4));
  fa fa_u_csamul_cla32_fa21_4_out(.a(u_csamul_cla32_and21_4[0]), .b(u_csamul_cla32_fa22_3_xor1[0]), .cin(u_csamul_cla32_fa21_3_or0[0]), .fa_xor1(u_csamul_cla32_fa21_4_xor1), .fa_or0(u_csamul_cla32_fa21_4_or0));
  and_gate and_gate_u_csamul_cla32_and22_4(.a(a[22]), .b(b[4]), .out(u_csamul_cla32_and22_4));
  fa fa_u_csamul_cla32_fa22_4_out(.a(u_csamul_cla32_and22_4[0]), .b(u_csamul_cla32_fa23_3_xor1[0]), .cin(u_csamul_cla32_fa22_3_or0[0]), .fa_xor1(u_csamul_cla32_fa22_4_xor1), .fa_or0(u_csamul_cla32_fa22_4_or0));
  and_gate and_gate_u_csamul_cla32_and23_4(.a(a[23]), .b(b[4]), .out(u_csamul_cla32_and23_4));
  fa fa_u_csamul_cla32_fa23_4_out(.a(u_csamul_cla32_and23_4[0]), .b(u_csamul_cla32_fa24_3_xor1[0]), .cin(u_csamul_cla32_fa23_3_or0[0]), .fa_xor1(u_csamul_cla32_fa23_4_xor1), .fa_or0(u_csamul_cla32_fa23_4_or0));
  and_gate and_gate_u_csamul_cla32_and24_4(.a(a[24]), .b(b[4]), .out(u_csamul_cla32_and24_4));
  fa fa_u_csamul_cla32_fa24_4_out(.a(u_csamul_cla32_and24_4[0]), .b(u_csamul_cla32_fa25_3_xor1[0]), .cin(u_csamul_cla32_fa24_3_or0[0]), .fa_xor1(u_csamul_cla32_fa24_4_xor1), .fa_or0(u_csamul_cla32_fa24_4_or0));
  and_gate and_gate_u_csamul_cla32_and25_4(.a(a[25]), .b(b[4]), .out(u_csamul_cla32_and25_4));
  fa fa_u_csamul_cla32_fa25_4_out(.a(u_csamul_cla32_and25_4[0]), .b(u_csamul_cla32_fa26_3_xor1[0]), .cin(u_csamul_cla32_fa25_3_or0[0]), .fa_xor1(u_csamul_cla32_fa25_4_xor1), .fa_or0(u_csamul_cla32_fa25_4_or0));
  and_gate and_gate_u_csamul_cla32_and26_4(.a(a[26]), .b(b[4]), .out(u_csamul_cla32_and26_4));
  fa fa_u_csamul_cla32_fa26_4_out(.a(u_csamul_cla32_and26_4[0]), .b(u_csamul_cla32_fa27_3_xor1[0]), .cin(u_csamul_cla32_fa26_3_or0[0]), .fa_xor1(u_csamul_cla32_fa26_4_xor1), .fa_or0(u_csamul_cla32_fa26_4_or0));
  and_gate and_gate_u_csamul_cla32_and27_4(.a(a[27]), .b(b[4]), .out(u_csamul_cla32_and27_4));
  fa fa_u_csamul_cla32_fa27_4_out(.a(u_csamul_cla32_and27_4[0]), .b(u_csamul_cla32_fa28_3_xor1[0]), .cin(u_csamul_cla32_fa27_3_or0[0]), .fa_xor1(u_csamul_cla32_fa27_4_xor1), .fa_or0(u_csamul_cla32_fa27_4_or0));
  and_gate and_gate_u_csamul_cla32_and28_4(.a(a[28]), .b(b[4]), .out(u_csamul_cla32_and28_4));
  fa fa_u_csamul_cla32_fa28_4_out(.a(u_csamul_cla32_and28_4[0]), .b(u_csamul_cla32_fa29_3_xor1[0]), .cin(u_csamul_cla32_fa28_3_or0[0]), .fa_xor1(u_csamul_cla32_fa28_4_xor1), .fa_or0(u_csamul_cla32_fa28_4_or0));
  and_gate and_gate_u_csamul_cla32_and29_4(.a(a[29]), .b(b[4]), .out(u_csamul_cla32_and29_4));
  fa fa_u_csamul_cla32_fa29_4_out(.a(u_csamul_cla32_and29_4[0]), .b(u_csamul_cla32_fa30_3_xor1[0]), .cin(u_csamul_cla32_fa29_3_or0[0]), .fa_xor1(u_csamul_cla32_fa29_4_xor1), .fa_or0(u_csamul_cla32_fa29_4_or0));
  and_gate and_gate_u_csamul_cla32_and30_4(.a(a[30]), .b(b[4]), .out(u_csamul_cla32_and30_4));
  fa fa_u_csamul_cla32_fa30_4_out(.a(u_csamul_cla32_and30_4[0]), .b(u_csamul_cla32_and31_3[0]), .cin(u_csamul_cla32_fa30_3_or0[0]), .fa_xor1(u_csamul_cla32_fa30_4_xor1), .fa_or0(u_csamul_cla32_fa30_4_or0));
  and_gate and_gate_u_csamul_cla32_and31_4(.a(a[31]), .b(b[4]), .out(u_csamul_cla32_and31_4));
  and_gate and_gate_u_csamul_cla32_and0_5(.a(a[0]), .b(b[5]), .out(u_csamul_cla32_and0_5));
  fa fa_u_csamul_cla32_fa0_5_out(.a(u_csamul_cla32_and0_5[0]), .b(u_csamul_cla32_fa1_4_xor1[0]), .cin(u_csamul_cla32_fa0_4_or0[0]), .fa_xor1(u_csamul_cla32_fa0_5_xor1), .fa_or0(u_csamul_cla32_fa0_5_or0));
  and_gate and_gate_u_csamul_cla32_and1_5(.a(a[1]), .b(b[5]), .out(u_csamul_cla32_and1_5));
  fa fa_u_csamul_cla32_fa1_5_out(.a(u_csamul_cla32_and1_5[0]), .b(u_csamul_cla32_fa2_4_xor1[0]), .cin(u_csamul_cla32_fa1_4_or0[0]), .fa_xor1(u_csamul_cla32_fa1_5_xor1), .fa_or0(u_csamul_cla32_fa1_5_or0));
  and_gate and_gate_u_csamul_cla32_and2_5(.a(a[2]), .b(b[5]), .out(u_csamul_cla32_and2_5));
  fa fa_u_csamul_cla32_fa2_5_out(.a(u_csamul_cla32_and2_5[0]), .b(u_csamul_cla32_fa3_4_xor1[0]), .cin(u_csamul_cla32_fa2_4_or0[0]), .fa_xor1(u_csamul_cla32_fa2_5_xor1), .fa_or0(u_csamul_cla32_fa2_5_or0));
  and_gate and_gate_u_csamul_cla32_and3_5(.a(a[3]), .b(b[5]), .out(u_csamul_cla32_and3_5));
  fa fa_u_csamul_cla32_fa3_5_out(.a(u_csamul_cla32_and3_5[0]), .b(u_csamul_cla32_fa4_4_xor1[0]), .cin(u_csamul_cla32_fa3_4_or0[0]), .fa_xor1(u_csamul_cla32_fa3_5_xor1), .fa_or0(u_csamul_cla32_fa3_5_or0));
  and_gate and_gate_u_csamul_cla32_and4_5(.a(a[4]), .b(b[5]), .out(u_csamul_cla32_and4_5));
  fa fa_u_csamul_cla32_fa4_5_out(.a(u_csamul_cla32_and4_5[0]), .b(u_csamul_cla32_fa5_4_xor1[0]), .cin(u_csamul_cla32_fa4_4_or0[0]), .fa_xor1(u_csamul_cla32_fa4_5_xor1), .fa_or0(u_csamul_cla32_fa4_5_or0));
  and_gate and_gate_u_csamul_cla32_and5_5(.a(a[5]), .b(b[5]), .out(u_csamul_cla32_and5_5));
  fa fa_u_csamul_cla32_fa5_5_out(.a(u_csamul_cla32_and5_5[0]), .b(u_csamul_cla32_fa6_4_xor1[0]), .cin(u_csamul_cla32_fa5_4_or0[0]), .fa_xor1(u_csamul_cla32_fa5_5_xor1), .fa_or0(u_csamul_cla32_fa5_5_or0));
  and_gate and_gate_u_csamul_cla32_and6_5(.a(a[6]), .b(b[5]), .out(u_csamul_cla32_and6_5));
  fa fa_u_csamul_cla32_fa6_5_out(.a(u_csamul_cla32_and6_5[0]), .b(u_csamul_cla32_fa7_4_xor1[0]), .cin(u_csamul_cla32_fa6_4_or0[0]), .fa_xor1(u_csamul_cla32_fa6_5_xor1), .fa_or0(u_csamul_cla32_fa6_5_or0));
  and_gate and_gate_u_csamul_cla32_and7_5(.a(a[7]), .b(b[5]), .out(u_csamul_cla32_and7_5));
  fa fa_u_csamul_cla32_fa7_5_out(.a(u_csamul_cla32_and7_5[0]), .b(u_csamul_cla32_fa8_4_xor1[0]), .cin(u_csamul_cla32_fa7_4_or0[0]), .fa_xor1(u_csamul_cla32_fa7_5_xor1), .fa_or0(u_csamul_cla32_fa7_5_or0));
  and_gate and_gate_u_csamul_cla32_and8_5(.a(a[8]), .b(b[5]), .out(u_csamul_cla32_and8_5));
  fa fa_u_csamul_cla32_fa8_5_out(.a(u_csamul_cla32_and8_5[0]), .b(u_csamul_cla32_fa9_4_xor1[0]), .cin(u_csamul_cla32_fa8_4_or0[0]), .fa_xor1(u_csamul_cla32_fa8_5_xor1), .fa_or0(u_csamul_cla32_fa8_5_or0));
  and_gate and_gate_u_csamul_cla32_and9_5(.a(a[9]), .b(b[5]), .out(u_csamul_cla32_and9_5));
  fa fa_u_csamul_cla32_fa9_5_out(.a(u_csamul_cla32_and9_5[0]), .b(u_csamul_cla32_fa10_4_xor1[0]), .cin(u_csamul_cla32_fa9_4_or0[0]), .fa_xor1(u_csamul_cla32_fa9_5_xor1), .fa_or0(u_csamul_cla32_fa9_5_or0));
  and_gate and_gate_u_csamul_cla32_and10_5(.a(a[10]), .b(b[5]), .out(u_csamul_cla32_and10_5));
  fa fa_u_csamul_cla32_fa10_5_out(.a(u_csamul_cla32_and10_5[0]), .b(u_csamul_cla32_fa11_4_xor1[0]), .cin(u_csamul_cla32_fa10_4_or0[0]), .fa_xor1(u_csamul_cla32_fa10_5_xor1), .fa_or0(u_csamul_cla32_fa10_5_or0));
  and_gate and_gate_u_csamul_cla32_and11_5(.a(a[11]), .b(b[5]), .out(u_csamul_cla32_and11_5));
  fa fa_u_csamul_cla32_fa11_5_out(.a(u_csamul_cla32_and11_5[0]), .b(u_csamul_cla32_fa12_4_xor1[0]), .cin(u_csamul_cla32_fa11_4_or0[0]), .fa_xor1(u_csamul_cla32_fa11_5_xor1), .fa_or0(u_csamul_cla32_fa11_5_or0));
  and_gate and_gate_u_csamul_cla32_and12_5(.a(a[12]), .b(b[5]), .out(u_csamul_cla32_and12_5));
  fa fa_u_csamul_cla32_fa12_5_out(.a(u_csamul_cla32_and12_5[0]), .b(u_csamul_cla32_fa13_4_xor1[0]), .cin(u_csamul_cla32_fa12_4_or0[0]), .fa_xor1(u_csamul_cla32_fa12_5_xor1), .fa_or0(u_csamul_cla32_fa12_5_or0));
  and_gate and_gate_u_csamul_cla32_and13_5(.a(a[13]), .b(b[5]), .out(u_csamul_cla32_and13_5));
  fa fa_u_csamul_cla32_fa13_5_out(.a(u_csamul_cla32_and13_5[0]), .b(u_csamul_cla32_fa14_4_xor1[0]), .cin(u_csamul_cla32_fa13_4_or0[0]), .fa_xor1(u_csamul_cla32_fa13_5_xor1), .fa_or0(u_csamul_cla32_fa13_5_or0));
  and_gate and_gate_u_csamul_cla32_and14_5(.a(a[14]), .b(b[5]), .out(u_csamul_cla32_and14_5));
  fa fa_u_csamul_cla32_fa14_5_out(.a(u_csamul_cla32_and14_5[0]), .b(u_csamul_cla32_fa15_4_xor1[0]), .cin(u_csamul_cla32_fa14_4_or0[0]), .fa_xor1(u_csamul_cla32_fa14_5_xor1), .fa_or0(u_csamul_cla32_fa14_5_or0));
  and_gate and_gate_u_csamul_cla32_and15_5(.a(a[15]), .b(b[5]), .out(u_csamul_cla32_and15_5));
  fa fa_u_csamul_cla32_fa15_5_out(.a(u_csamul_cla32_and15_5[0]), .b(u_csamul_cla32_fa16_4_xor1[0]), .cin(u_csamul_cla32_fa15_4_or0[0]), .fa_xor1(u_csamul_cla32_fa15_5_xor1), .fa_or0(u_csamul_cla32_fa15_5_or0));
  and_gate and_gate_u_csamul_cla32_and16_5(.a(a[16]), .b(b[5]), .out(u_csamul_cla32_and16_5));
  fa fa_u_csamul_cla32_fa16_5_out(.a(u_csamul_cla32_and16_5[0]), .b(u_csamul_cla32_fa17_4_xor1[0]), .cin(u_csamul_cla32_fa16_4_or0[0]), .fa_xor1(u_csamul_cla32_fa16_5_xor1), .fa_or0(u_csamul_cla32_fa16_5_or0));
  and_gate and_gate_u_csamul_cla32_and17_5(.a(a[17]), .b(b[5]), .out(u_csamul_cla32_and17_5));
  fa fa_u_csamul_cla32_fa17_5_out(.a(u_csamul_cla32_and17_5[0]), .b(u_csamul_cla32_fa18_4_xor1[0]), .cin(u_csamul_cla32_fa17_4_or0[0]), .fa_xor1(u_csamul_cla32_fa17_5_xor1), .fa_or0(u_csamul_cla32_fa17_5_or0));
  and_gate and_gate_u_csamul_cla32_and18_5(.a(a[18]), .b(b[5]), .out(u_csamul_cla32_and18_5));
  fa fa_u_csamul_cla32_fa18_5_out(.a(u_csamul_cla32_and18_5[0]), .b(u_csamul_cla32_fa19_4_xor1[0]), .cin(u_csamul_cla32_fa18_4_or0[0]), .fa_xor1(u_csamul_cla32_fa18_5_xor1), .fa_or0(u_csamul_cla32_fa18_5_or0));
  and_gate and_gate_u_csamul_cla32_and19_5(.a(a[19]), .b(b[5]), .out(u_csamul_cla32_and19_5));
  fa fa_u_csamul_cla32_fa19_5_out(.a(u_csamul_cla32_and19_5[0]), .b(u_csamul_cla32_fa20_4_xor1[0]), .cin(u_csamul_cla32_fa19_4_or0[0]), .fa_xor1(u_csamul_cla32_fa19_5_xor1), .fa_or0(u_csamul_cla32_fa19_5_or0));
  and_gate and_gate_u_csamul_cla32_and20_5(.a(a[20]), .b(b[5]), .out(u_csamul_cla32_and20_5));
  fa fa_u_csamul_cla32_fa20_5_out(.a(u_csamul_cla32_and20_5[0]), .b(u_csamul_cla32_fa21_4_xor1[0]), .cin(u_csamul_cla32_fa20_4_or0[0]), .fa_xor1(u_csamul_cla32_fa20_5_xor1), .fa_or0(u_csamul_cla32_fa20_5_or0));
  and_gate and_gate_u_csamul_cla32_and21_5(.a(a[21]), .b(b[5]), .out(u_csamul_cla32_and21_5));
  fa fa_u_csamul_cla32_fa21_5_out(.a(u_csamul_cla32_and21_5[0]), .b(u_csamul_cla32_fa22_4_xor1[0]), .cin(u_csamul_cla32_fa21_4_or0[0]), .fa_xor1(u_csamul_cla32_fa21_5_xor1), .fa_or0(u_csamul_cla32_fa21_5_or0));
  and_gate and_gate_u_csamul_cla32_and22_5(.a(a[22]), .b(b[5]), .out(u_csamul_cla32_and22_5));
  fa fa_u_csamul_cla32_fa22_5_out(.a(u_csamul_cla32_and22_5[0]), .b(u_csamul_cla32_fa23_4_xor1[0]), .cin(u_csamul_cla32_fa22_4_or0[0]), .fa_xor1(u_csamul_cla32_fa22_5_xor1), .fa_or0(u_csamul_cla32_fa22_5_or0));
  and_gate and_gate_u_csamul_cla32_and23_5(.a(a[23]), .b(b[5]), .out(u_csamul_cla32_and23_5));
  fa fa_u_csamul_cla32_fa23_5_out(.a(u_csamul_cla32_and23_5[0]), .b(u_csamul_cla32_fa24_4_xor1[0]), .cin(u_csamul_cla32_fa23_4_or0[0]), .fa_xor1(u_csamul_cla32_fa23_5_xor1), .fa_or0(u_csamul_cla32_fa23_5_or0));
  and_gate and_gate_u_csamul_cla32_and24_5(.a(a[24]), .b(b[5]), .out(u_csamul_cla32_and24_5));
  fa fa_u_csamul_cla32_fa24_5_out(.a(u_csamul_cla32_and24_5[0]), .b(u_csamul_cla32_fa25_4_xor1[0]), .cin(u_csamul_cla32_fa24_4_or0[0]), .fa_xor1(u_csamul_cla32_fa24_5_xor1), .fa_or0(u_csamul_cla32_fa24_5_or0));
  and_gate and_gate_u_csamul_cla32_and25_5(.a(a[25]), .b(b[5]), .out(u_csamul_cla32_and25_5));
  fa fa_u_csamul_cla32_fa25_5_out(.a(u_csamul_cla32_and25_5[0]), .b(u_csamul_cla32_fa26_4_xor1[0]), .cin(u_csamul_cla32_fa25_4_or0[0]), .fa_xor1(u_csamul_cla32_fa25_5_xor1), .fa_or0(u_csamul_cla32_fa25_5_or0));
  and_gate and_gate_u_csamul_cla32_and26_5(.a(a[26]), .b(b[5]), .out(u_csamul_cla32_and26_5));
  fa fa_u_csamul_cla32_fa26_5_out(.a(u_csamul_cla32_and26_5[0]), .b(u_csamul_cla32_fa27_4_xor1[0]), .cin(u_csamul_cla32_fa26_4_or0[0]), .fa_xor1(u_csamul_cla32_fa26_5_xor1), .fa_or0(u_csamul_cla32_fa26_5_or0));
  and_gate and_gate_u_csamul_cla32_and27_5(.a(a[27]), .b(b[5]), .out(u_csamul_cla32_and27_5));
  fa fa_u_csamul_cla32_fa27_5_out(.a(u_csamul_cla32_and27_5[0]), .b(u_csamul_cla32_fa28_4_xor1[0]), .cin(u_csamul_cla32_fa27_4_or0[0]), .fa_xor1(u_csamul_cla32_fa27_5_xor1), .fa_or0(u_csamul_cla32_fa27_5_or0));
  and_gate and_gate_u_csamul_cla32_and28_5(.a(a[28]), .b(b[5]), .out(u_csamul_cla32_and28_5));
  fa fa_u_csamul_cla32_fa28_5_out(.a(u_csamul_cla32_and28_5[0]), .b(u_csamul_cla32_fa29_4_xor1[0]), .cin(u_csamul_cla32_fa28_4_or0[0]), .fa_xor1(u_csamul_cla32_fa28_5_xor1), .fa_or0(u_csamul_cla32_fa28_5_or0));
  and_gate and_gate_u_csamul_cla32_and29_5(.a(a[29]), .b(b[5]), .out(u_csamul_cla32_and29_5));
  fa fa_u_csamul_cla32_fa29_5_out(.a(u_csamul_cla32_and29_5[0]), .b(u_csamul_cla32_fa30_4_xor1[0]), .cin(u_csamul_cla32_fa29_4_or0[0]), .fa_xor1(u_csamul_cla32_fa29_5_xor1), .fa_or0(u_csamul_cla32_fa29_5_or0));
  and_gate and_gate_u_csamul_cla32_and30_5(.a(a[30]), .b(b[5]), .out(u_csamul_cla32_and30_5));
  fa fa_u_csamul_cla32_fa30_5_out(.a(u_csamul_cla32_and30_5[0]), .b(u_csamul_cla32_and31_4[0]), .cin(u_csamul_cla32_fa30_4_or0[0]), .fa_xor1(u_csamul_cla32_fa30_5_xor1), .fa_or0(u_csamul_cla32_fa30_5_or0));
  and_gate and_gate_u_csamul_cla32_and31_5(.a(a[31]), .b(b[5]), .out(u_csamul_cla32_and31_5));
  and_gate and_gate_u_csamul_cla32_and0_6(.a(a[0]), .b(b[6]), .out(u_csamul_cla32_and0_6));
  fa fa_u_csamul_cla32_fa0_6_out(.a(u_csamul_cla32_and0_6[0]), .b(u_csamul_cla32_fa1_5_xor1[0]), .cin(u_csamul_cla32_fa0_5_or0[0]), .fa_xor1(u_csamul_cla32_fa0_6_xor1), .fa_or0(u_csamul_cla32_fa0_6_or0));
  and_gate and_gate_u_csamul_cla32_and1_6(.a(a[1]), .b(b[6]), .out(u_csamul_cla32_and1_6));
  fa fa_u_csamul_cla32_fa1_6_out(.a(u_csamul_cla32_and1_6[0]), .b(u_csamul_cla32_fa2_5_xor1[0]), .cin(u_csamul_cla32_fa1_5_or0[0]), .fa_xor1(u_csamul_cla32_fa1_6_xor1), .fa_or0(u_csamul_cla32_fa1_6_or0));
  and_gate and_gate_u_csamul_cla32_and2_6(.a(a[2]), .b(b[6]), .out(u_csamul_cla32_and2_6));
  fa fa_u_csamul_cla32_fa2_6_out(.a(u_csamul_cla32_and2_6[0]), .b(u_csamul_cla32_fa3_5_xor1[0]), .cin(u_csamul_cla32_fa2_5_or0[0]), .fa_xor1(u_csamul_cla32_fa2_6_xor1), .fa_or0(u_csamul_cla32_fa2_6_or0));
  and_gate and_gate_u_csamul_cla32_and3_6(.a(a[3]), .b(b[6]), .out(u_csamul_cla32_and3_6));
  fa fa_u_csamul_cla32_fa3_6_out(.a(u_csamul_cla32_and3_6[0]), .b(u_csamul_cla32_fa4_5_xor1[0]), .cin(u_csamul_cla32_fa3_5_or0[0]), .fa_xor1(u_csamul_cla32_fa3_6_xor1), .fa_or0(u_csamul_cla32_fa3_6_or0));
  and_gate and_gate_u_csamul_cla32_and4_6(.a(a[4]), .b(b[6]), .out(u_csamul_cla32_and4_6));
  fa fa_u_csamul_cla32_fa4_6_out(.a(u_csamul_cla32_and4_6[0]), .b(u_csamul_cla32_fa5_5_xor1[0]), .cin(u_csamul_cla32_fa4_5_or0[0]), .fa_xor1(u_csamul_cla32_fa4_6_xor1), .fa_or0(u_csamul_cla32_fa4_6_or0));
  and_gate and_gate_u_csamul_cla32_and5_6(.a(a[5]), .b(b[6]), .out(u_csamul_cla32_and5_6));
  fa fa_u_csamul_cla32_fa5_6_out(.a(u_csamul_cla32_and5_6[0]), .b(u_csamul_cla32_fa6_5_xor1[0]), .cin(u_csamul_cla32_fa5_5_or0[0]), .fa_xor1(u_csamul_cla32_fa5_6_xor1), .fa_or0(u_csamul_cla32_fa5_6_or0));
  and_gate and_gate_u_csamul_cla32_and6_6(.a(a[6]), .b(b[6]), .out(u_csamul_cla32_and6_6));
  fa fa_u_csamul_cla32_fa6_6_out(.a(u_csamul_cla32_and6_6[0]), .b(u_csamul_cla32_fa7_5_xor1[0]), .cin(u_csamul_cla32_fa6_5_or0[0]), .fa_xor1(u_csamul_cla32_fa6_6_xor1), .fa_or0(u_csamul_cla32_fa6_6_or0));
  and_gate and_gate_u_csamul_cla32_and7_6(.a(a[7]), .b(b[6]), .out(u_csamul_cla32_and7_6));
  fa fa_u_csamul_cla32_fa7_6_out(.a(u_csamul_cla32_and7_6[0]), .b(u_csamul_cla32_fa8_5_xor1[0]), .cin(u_csamul_cla32_fa7_5_or0[0]), .fa_xor1(u_csamul_cla32_fa7_6_xor1), .fa_or0(u_csamul_cla32_fa7_6_or0));
  and_gate and_gate_u_csamul_cla32_and8_6(.a(a[8]), .b(b[6]), .out(u_csamul_cla32_and8_6));
  fa fa_u_csamul_cla32_fa8_6_out(.a(u_csamul_cla32_and8_6[0]), .b(u_csamul_cla32_fa9_5_xor1[0]), .cin(u_csamul_cla32_fa8_5_or0[0]), .fa_xor1(u_csamul_cla32_fa8_6_xor1), .fa_or0(u_csamul_cla32_fa8_6_or0));
  and_gate and_gate_u_csamul_cla32_and9_6(.a(a[9]), .b(b[6]), .out(u_csamul_cla32_and9_6));
  fa fa_u_csamul_cla32_fa9_6_out(.a(u_csamul_cla32_and9_6[0]), .b(u_csamul_cla32_fa10_5_xor1[0]), .cin(u_csamul_cla32_fa9_5_or0[0]), .fa_xor1(u_csamul_cla32_fa9_6_xor1), .fa_or0(u_csamul_cla32_fa9_6_or0));
  and_gate and_gate_u_csamul_cla32_and10_6(.a(a[10]), .b(b[6]), .out(u_csamul_cla32_and10_6));
  fa fa_u_csamul_cla32_fa10_6_out(.a(u_csamul_cla32_and10_6[0]), .b(u_csamul_cla32_fa11_5_xor1[0]), .cin(u_csamul_cla32_fa10_5_or0[0]), .fa_xor1(u_csamul_cla32_fa10_6_xor1), .fa_or0(u_csamul_cla32_fa10_6_or0));
  and_gate and_gate_u_csamul_cla32_and11_6(.a(a[11]), .b(b[6]), .out(u_csamul_cla32_and11_6));
  fa fa_u_csamul_cla32_fa11_6_out(.a(u_csamul_cla32_and11_6[0]), .b(u_csamul_cla32_fa12_5_xor1[0]), .cin(u_csamul_cla32_fa11_5_or0[0]), .fa_xor1(u_csamul_cla32_fa11_6_xor1), .fa_or0(u_csamul_cla32_fa11_6_or0));
  and_gate and_gate_u_csamul_cla32_and12_6(.a(a[12]), .b(b[6]), .out(u_csamul_cla32_and12_6));
  fa fa_u_csamul_cla32_fa12_6_out(.a(u_csamul_cla32_and12_6[0]), .b(u_csamul_cla32_fa13_5_xor1[0]), .cin(u_csamul_cla32_fa12_5_or0[0]), .fa_xor1(u_csamul_cla32_fa12_6_xor1), .fa_or0(u_csamul_cla32_fa12_6_or0));
  and_gate and_gate_u_csamul_cla32_and13_6(.a(a[13]), .b(b[6]), .out(u_csamul_cla32_and13_6));
  fa fa_u_csamul_cla32_fa13_6_out(.a(u_csamul_cla32_and13_6[0]), .b(u_csamul_cla32_fa14_5_xor1[0]), .cin(u_csamul_cla32_fa13_5_or0[0]), .fa_xor1(u_csamul_cla32_fa13_6_xor1), .fa_or0(u_csamul_cla32_fa13_6_or0));
  and_gate and_gate_u_csamul_cla32_and14_6(.a(a[14]), .b(b[6]), .out(u_csamul_cla32_and14_6));
  fa fa_u_csamul_cla32_fa14_6_out(.a(u_csamul_cla32_and14_6[0]), .b(u_csamul_cla32_fa15_5_xor1[0]), .cin(u_csamul_cla32_fa14_5_or0[0]), .fa_xor1(u_csamul_cla32_fa14_6_xor1), .fa_or0(u_csamul_cla32_fa14_6_or0));
  and_gate and_gate_u_csamul_cla32_and15_6(.a(a[15]), .b(b[6]), .out(u_csamul_cla32_and15_6));
  fa fa_u_csamul_cla32_fa15_6_out(.a(u_csamul_cla32_and15_6[0]), .b(u_csamul_cla32_fa16_5_xor1[0]), .cin(u_csamul_cla32_fa15_5_or0[0]), .fa_xor1(u_csamul_cla32_fa15_6_xor1), .fa_or0(u_csamul_cla32_fa15_6_or0));
  and_gate and_gate_u_csamul_cla32_and16_6(.a(a[16]), .b(b[6]), .out(u_csamul_cla32_and16_6));
  fa fa_u_csamul_cla32_fa16_6_out(.a(u_csamul_cla32_and16_6[0]), .b(u_csamul_cla32_fa17_5_xor1[0]), .cin(u_csamul_cla32_fa16_5_or0[0]), .fa_xor1(u_csamul_cla32_fa16_6_xor1), .fa_or0(u_csamul_cla32_fa16_6_or0));
  and_gate and_gate_u_csamul_cla32_and17_6(.a(a[17]), .b(b[6]), .out(u_csamul_cla32_and17_6));
  fa fa_u_csamul_cla32_fa17_6_out(.a(u_csamul_cla32_and17_6[0]), .b(u_csamul_cla32_fa18_5_xor1[0]), .cin(u_csamul_cla32_fa17_5_or0[0]), .fa_xor1(u_csamul_cla32_fa17_6_xor1), .fa_or0(u_csamul_cla32_fa17_6_or0));
  and_gate and_gate_u_csamul_cla32_and18_6(.a(a[18]), .b(b[6]), .out(u_csamul_cla32_and18_6));
  fa fa_u_csamul_cla32_fa18_6_out(.a(u_csamul_cla32_and18_6[0]), .b(u_csamul_cla32_fa19_5_xor1[0]), .cin(u_csamul_cla32_fa18_5_or0[0]), .fa_xor1(u_csamul_cla32_fa18_6_xor1), .fa_or0(u_csamul_cla32_fa18_6_or0));
  and_gate and_gate_u_csamul_cla32_and19_6(.a(a[19]), .b(b[6]), .out(u_csamul_cla32_and19_6));
  fa fa_u_csamul_cla32_fa19_6_out(.a(u_csamul_cla32_and19_6[0]), .b(u_csamul_cla32_fa20_5_xor1[0]), .cin(u_csamul_cla32_fa19_5_or0[0]), .fa_xor1(u_csamul_cla32_fa19_6_xor1), .fa_or0(u_csamul_cla32_fa19_6_or0));
  and_gate and_gate_u_csamul_cla32_and20_6(.a(a[20]), .b(b[6]), .out(u_csamul_cla32_and20_6));
  fa fa_u_csamul_cla32_fa20_6_out(.a(u_csamul_cla32_and20_6[0]), .b(u_csamul_cla32_fa21_5_xor1[0]), .cin(u_csamul_cla32_fa20_5_or0[0]), .fa_xor1(u_csamul_cla32_fa20_6_xor1), .fa_or0(u_csamul_cla32_fa20_6_or0));
  and_gate and_gate_u_csamul_cla32_and21_6(.a(a[21]), .b(b[6]), .out(u_csamul_cla32_and21_6));
  fa fa_u_csamul_cla32_fa21_6_out(.a(u_csamul_cla32_and21_6[0]), .b(u_csamul_cla32_fa22_5_xor1[0]), .cin(u_csamul_cla32_fa21_5_or0[0]), .fa_xor1(u_csamul_cla32_fa21_6_xor1), .fa_or0(u_csamul_cla32_fa21_6_or0));
  and_gate and_gate_u_csamul_cla32_and22_6(.a(a[22]), .b(b[6]), .out(u_csamul_cla32_and22_6));
  fa fa_u_csamul_cla32_fa22_6_out(.a(u_csamul_cla32_and22_6[0]), .b(u_csamul_cla32_fa23_5_xor1[0]), .cin(u_csamul_cla32_fa22_5_or0[0]), .fa_xor1(u_csamul_cla32_fa22_6_xor1), .fa_or0(u_csamul_cla32_fa22_6_or0));
  and_gate and_gate_u_csamul_cla32_and23_6(.a(a[23]), .b(b[6]), .out(u_csamul_cla32_and23_6));
  fa fa_u_csamul_cla32_fa23_6_out(.a(u_csamul_cla32_and23_6[0]), .b(u_csamul_cla32_fa24_5_xor1[0]), .cin(u_csamul_cla32_fa23_5_or0[0]), .fa_xor1(u_csamul_cla32_fa23_6_xor1), .fa_or0(u_csamul_cla32_fa23_6_or0));
  and_gate and_gate_u_csamul_cla32_and24_6(.a(a[24]), .b(b[6]), .out(u_csamul_cla32_and24_6));
  fa fa_u_csamul_cla32_fa24_6_out(.a(u_csamul_cla32_and24_6[0]), .b(u_csamul_cla32_fa25_5_xor1[0]), .cin(u_csamul_cla32_fa24_5_or0[0]), .fa_xor1(u_csamul_cla32_fa24_6_xor1), .fa_or0(u_csamul_cla32_fa24_6_or0));
  and_gate and_gate_u_csamul_cla32_and25_6(.a(a[25]), .b(b[6]), .out(u_csamul_cla32_and25_6));
  fa fa_u_csamul_cla32_fa25_6_out(.a(u_csamul_cla32_and25_6[0]), .b(u_csamul_cla32_fa26_5_xor1[0]), .cin(u_csamul_cla32_fa25_5_or0[0]), .fa_xor1(u_csamul_cla32_fa25_6_xor1), .fa_or0(u_csamul_cla32_fa25_6_or0));
  and_gate and_gate_u_csamul_cla32_and26_6(.a(a[26]), .b(b[6]), .out(u_csamul_cla32_and26_6));
  fa fa_u_csamul_cla32_fa26_6_out(.a(u_csamul_cla32_and26_6[0]), .b(u_csamul_cla32_fa27_5_xor1[0]), .cin(u_csamul_cla32_fa26_5_or0[0]), .fa_xor1(u_csamul_cla32_fa26_6_xor1), .fa_or0(u_csamul_cla32_fa26_6_or0));
  and_gate and_gate_u_csamul_cla32_and27_6(.a(a[27]), .b(b[6]), .out(u_csamul_cla32_and27_6));
  fa fa_u_csamul_cla32_fa27_6_out(.a(u_csamul_cla32_and27_6[0]), .b(u_csamul_cla32_fa28_5_xor1[0]), .cin(u_csamul_cla32_fa27_5_or0[0]), .fa_xor1(u_csamul_cla32_fa27_6_xor1), .fa_or0(u_csamul_cla32_fa27_6_or0));
  and_gate and_gate_u_csamul_cla32_and28_6(.a(a[28]), .b(b[6]), .out(u_csamul_cla32_and28_6));
  fa fa_u_csamul_cla32_fa28_6_out(.a(u_csamul_cla32_and28_6[0]), .b(u_csamul_cla32_fa29_5_xor1[0]), .cin(u_csamul_cla32_fa28_5_or0[0]), .fa_xor1(u_csamul_cla32_fa28_6_xor1), .fa_or0(u_csamul_cla32_fa28_6_or0));
  and_gate and_gate_u_csamul_cla32_and29_6(.a(a[29]), .b(b[6]), .out(u_csamul_cla32_and29_6));
  fa fa_u_csamul_cla32_fa29_6_out(.a(u_csamul_cla32_and29_6[0]), .b(u_csamul_cla32_fa30_5_xor1[0]), .cin(u_csamul_cla32_fa29_5_or0[0]), .fa_xor1(u_csamul_cla32_fa29_6_xor1), .fa_or0(u_csamul_cla32_fa29_6_or0));
  and_gate and_gate_u_csamul_cla32_and30_6(.a(a[30]), .b(b[6]), .out(u_csamul_cla32_and30_6));
  fa fa_u_csamul_cla32_fa30_6_out(.a(u_csamul_cla32_and30_6[0]), .b(u_csamul_cla32_and31_5[0]), .cin(u_csamul_cla32_fa30_5_or0[0]), .fa_xor1(u_csamul_cla32_fa30_6_xor1), .fa_or0(u_csamul_cla32_fa30_6_or0));
  and_gate and_gate_u_csamul_cla32_and31_6(.a(a[31]), .b(b[6]), .out(u_csamul_cla32_and31_6));
  and_gate and_gate_u_csamul_cla32_and0_7(.a(a[0]), .b(b[7]), .out(u_csamul_cla32_and0_7));
  fa fa_u_csamul_cla32_fa0_7_out(.a(u_csamul_cla32_and0_7[0]), .b(u_csamul_cla32_fa1_6_xor1[0]), .cin(u_csamul_cla32_fa0_6_or0[0]), .fa_xor1(u_csamul_cla32_fa0_7_xor1), .fa_or0(u_csamul_cla32_fa0_7_or0));
  and_gate and_gate_u_csamul_cla32_and1_7(.a(a[1]), .b(b[7]), .out(u_csamul_cla32_and1_7));
  fa fa_u_csamul_cla32_fa1_7_out(.a(u_csamul_cla32_and1_7[0]), .b(u_csamul_cla32_fa2_6_xor1[0]), .cin(u_csamul_cla32_fa1_6_or0[0]), .fa_xor1(u_csamul_cla32_fa1_7_xor1), .fa_or0(u_csamul_cla32_fa1_7_or0));
  and_gate and_gate_u_csamul_cla32_and2_7(.a(a[2]), .b(b[7]), .out(u_csamul_cla32_and2_7));
  fa fa_u_csamul_cla32_fa2_7_out(.a(u_csamul_cla32_and2_7[0]), .b(u_csamul_cla32_fa3_6_xor1[0]), .cin(u_csamul_cla32_fa2_6_or0[0]), .fa_xor1(u_csamul_cla32_fa2_7_xor1), .fa_or0(u_csamul_cla32_fa2_7_or0));
  and_gate and_gate_u_csamul_cla32_and3_7(.a(a[3]), .b(b[7]), .out(u_csamul_cla32_and3_7));
  fa fa_u_csamul_cla32_fa3_7_out(.a(u_csamul_cla32_and3_7[0]), .b(u_csamul_cla32_fa4_6_xor1[0]), .cin(u_csamul_cla32_fa3_6_or0[0]), .fa_xor1(u_csamul_cla32_fa3_7_xor1), .fa_or0(u_csamul_cla32_fa3_7_or0));
  and_gate and_gate_u_csamul_cla32_and4_7(.a(a[4]), .b(b[7]), .out(u_csamul_cla32_and4_7));
  fa fa_u_csamul_cla32_fa4_7_out(.a(u_csamul_cla32_and4_7[0]), .b(u_csamul_cla32_fa5_6_xor1[0]), .cin(u_csamul_cla32_fa4_6_or0[0]), .fa_xor1(u_csamul_cla32_fa4_7_xor1), .fa_or0(u_csamul_cla32_fa4_7_or0));
  and_gate and_gate_u_csamul_cla32_and5_7(.a(a[5]), .b(b[7]), .out(u_csamul_cla32_and5_7));
  fa fa_u_csamul_cla32_fa5_7_out(.a(u_csamul_cla32_and5_7[0]), .b(u_csamul_cla32_fa6_6_xor1[0]), .cin(u_csamul_cla32_fa5_6_or0[0]), .fa_xor1(u_csamul_cla32_fa5_7_xor1), .fa_or0(u_csamul_cla32_fa5_7_or0));
  and_gate and_gate_u_csamul_cla32_and6_7(.a(a[6]), .b(b[7]), .out(u_csamul_cla32_and6_7));
  fa fa_u_csamul_cla32_fa6_7_out(.a(u_csamul_cla32_and6_7[0]), .b(u_csamul_cla32_fa7_6_xor1[0]), .cin(u_csamul_cla32_fa6_6_or0[0]), .fa_xor1(u_csamul_cla32_fa6_7_xor1), .fa_or0(u_csamul_cla32_fa6_7_or0));
  and_gate and_gate_u_csamul_cla32_and7_7(.a(a[7]), .b(b[7]), .out(u_csamul_cla32_and7_7));
  fa fa_u_csamul_cla32_fa7_7_out(.a(u_csamul_cla32_and7_7[0]), .b(u_csamul_cla32_fa8_6_xor1[0]), .cin(u_csamul_cla32_fa7_6_or0[0]), .fa_xor1(u_csamul_cla32_fa7_7_xor1), .fa_or0(u_csamul_cla32_fa7_7_or0));
  and_gate and_gate_u_csamul_cla32_and8_7(.a(a[8]), .b(b[7]), .out(u_csamul_cla32_and8_7));
  fa fa_u_csamul_cla32_fa8_7_out(.a(u_csamul_cla32_and8_7[0]), .b(u_csamul_cla32_fa9_6_xor1[0]), .cin(u_csamul_cla32_fa8_6_or0[0]), .fa_xor1(u_csamul_cla32_fa8_7_xor1), .fa_or0(u_csamul_cla32_fa8_7_or0));
  and_gate and_gate_u_csamul_cla32_and9_7(.a(a[9]), .b(b[7]), .out(u_csamul_cla32_and9_7));
  fa fa_u_csamul_cla32_fa9_7_out(.a(u_csamul_cla32_and9_7[0]), .b(u_csamul_cla32_fa10_6_xor1[0]), .cin(u_csamul_cla32_fa9_6_or0[0]), .fa_xor1(u_csamul_cla32_fa9_7_xor1), .fa_or0(u_csamul_cla32_fa9_7_or0));
  and_gate and_gate_u_csamul_cla32_and10_7(.a(a[10]), .b(b[7]), .out(u_csamul_cla32_and10_7));
  fa fa_u_csamul_cla32_fa10_7_out(.a(u_csamul_cla32_and10_7[0]), .b(u_csamul_cla32_fa11_6_xor1[0]), .cin(u_csamul_cla32_fa10_6_or0[0]), .fa_xor1(u_csamul_cla32_fa10_7_xor1), .fa_or0(u_csamul_cla32_fa10_7_or0));
  and_gate and_gate_u_csamul_cla32_and11_7(.a(a[11]), .b(b[7]), .out(u_csamul_cla32_and11_7));
  fa fa_u_csamul_cla32_fa11_7_out(.a(u_csamul_cla32_and11_7[0]), .b(u_csamul_cla32_fa12_6_xor1[0]), .cin(u_csamul_cla32_fa11_6_or0[0]), .fa_xor1(u_csamul_cla32_fa11_7_xor1), .fa_or0(u_csamul_cla32_fa11_7_or0));
  and_gate and_gate_u_csamul_cla32_and12_7(.a(a[12]), .b(b[7]), .out(u_csamul_cla32_and12_7));
  fa fa_u_csamul_cla32_fa12_7_out(.a(u_csamul_cla32_and12_7[0]), .b(u_csamul_cla32_fa13_6_xor1[0]), .cin(u_csamul_cla32_fa12_6_or0[0]), .fa_xor1(u_csamul_cla32_fa12_7_xor1), .fa_or0(u_csamul_cla32_fa12_7_or0));
  and_gate and_gate_u_csamul_cla32_and13_7(.a(a[13]), .b(b[7]), .out(u_csamul_cla32_and13_7));
  fa fa_u_csamul_cla32_fa13_7_out(.a(u_csamul_cla32_and13_7[0]), .b(u_csamul_cla32_fa14_6_xor1[0]), .cin(u_csamul_cla32_fa13_6_or0[0]), .fa_xor1(u_csamul_cla32_fa13_7_xor1), .fa_or0(u_csamul_cla32_fa13_7_or0));
  and_gate and_gate_u_csamul_cla32_and14_7(.a(a[14]), .b(b[7]), .out(u_csamul_cla32_and14_7));
  fa fa_u_csamul_cla32_fa14_7_out(.a(u_csamul_cla32_and14_7[0]), .b(u_csamul_cla32_fa15_6_xor1[0]), .cin(u_csamul_cla32_fa14_6_or0[0]), .fa_xor1(u_csamul_cla32_fa14_7_xor1), .fa_or0(u_csamul_cla32_fa14_7_or0));
  and_gate and_gate_u_csamul_cla32_and15_7(.a(a[15]), .b(b[7]), .out(u_csamul_cla32_and15_7));
  fa fa_u_csamul_cla32_fa15_7_out(.a(u_csamul_cla32_and15_7[0]), .b(u_csamul_cla32_fa16_6_xor1[0]), .cin(u_csamul_cla32_fa15_6_or0[0]), .fa_xor1(u_csamul_cla32_fa15_7_xor1), .fa_or0(u_csamul_cla32_fa15_7_or0));
  and_gate and_gate_u_csamul_cla32_and16_7(.a(a[16]), .b(b[7]), .out(u_csamul_cla32_and16_7));
  fa fa_u_csamul_cla32_fa16_7_out(.a(u_csamul_cla32_and16_7[0]), .b(u_csamul_cla32_fa17_6_xor1[0]), .cin(u_csamul_cla32_fa16_6_or0[0]), .fa_xor1(u_csamul_cla32_fa16_7_xor1), .fa_or0(u_csamul_cla32_fa16_7_or0));
  and_gate and_gate_u_csamul_cla32_and17_7(.a(a[17]), .b(b[7]), .out(u_csamul_cla32_and17_7));
  fa fa_u_csamul_cla32_fa17_7_out(.a(u_csamul_cla32_and17_7[0]), .b(u_csamul_cla32_fa18_6_xor1[0]), .cin(u_csamul_cla32_fa17_6_or0[0]), .fa_xor1(u_csamul_cla32_fa17_7_xor1), .fa_or0(u_csamul_cla32_fa17_7_or0));
  and_gate and_gate_u_csamul_cla32_and18_7(.a(a[18]), .b(b[7]), .out(u_csamul_cla32_and18_7));
  fa fa_u_csamul_cla32_fa18_7_out(.a(u_csamul_cla32_and18_7[0]), .b(u_csamul_cla32_fa19_6_xor1[0]), .cin(u_csamul_cla32_fa18_6_or0[0]), .fa_xor1(u_csamul_cla32_fa18_7_xor1), .fa_or0(u_csamul_cla32_fa18_7_or0));
  and_gate and_gate_u_csamul_cla32_and19_7(.a(a[19]), .b(b[7]), .out(u_csamul_cla32_and19_7));
  fa fa_u_csamul_cla32_fa19_7_out(.a(u_csamul_cla32_and19_7[0]), .b(u_csamul_cla32_fa20_6_xor1[0]), .cin(u_csamul_cla32_fa19_6_or0[0]), .fa_xor1(u_csamul_cla32_fa19_7_xor1), .fa_or0(u_csamul_cla32_fa19_7_or0));
  and_gate and_gate_u_csamul_cla32_and20_7(.a(a[20]), .b(b[7]), .out(u_csamul_cla32_and20_7));
  fa fa_u_csamul_cla32_fa20_7_out(.a(u_csamul_cla32_and20_7[0]), .b(u_csamul_cla32_fa21_6_xor1[0]), .cin(u_csamul_cla32_fa20_6_or0[0]), .fa_xor1(u_csamul_cla32_fa20_7_xor1), .fa_or0(u_csamul_cla32_fa20_7_or0));
  and_gate and_gate_u_csamul_cla32_and21_7(.a(a[21]), .b(b[7]), .out(u_csamul_cla32_and21_7));
  fa fa_u_csamul_cla32_fa21_7_out(.a(u_csamul_cla32_and21_7[0]), .b(u_csamul_cla32_fa22_6_xor1[0]), .cin(u_csamul_cla32_fa21_6_or0[0]), .fa_xor1(u_csamul_cla32_fa21_7_xor1), .fa_or0(u_csamul_cla32_fa21_7_or0));
  and_gate and_gate_u_csamul_cla32_and22_7(.a(a[22]), .b(b[7]), .out(u_csamul_cla32_and22_7));
  fa fa_u_csamul_cla32_fa22_7_out(.a(u_csamul_cla32_and22_7[0]), .b(u_csamul_cla32_fa23_6_xor1[0]), .cin(u_csamul_cla32_fa22_6_or0[0]), .fa_xor1(u_csamul_cla32_fa22_7_xor1), .fa_or0(u_csamul_cla32_fa22_7_or0));
  and_gate and_gate_u_csamul_cla32_and23_7(.a(a[23]), .b(b[7]), .out(u_csamul_cla32_and23_7));
  fa fa_u_csamul_cla32_fa23_7_out(.a(u_csamul_cla32_and23_7[0]), .b(u_csamul_cla32_fa24_6_xor1[0]), .cin(u_csamul_cla32_fa23_6_or0[0]), .fa_xor1(u_csamul_cla32_fa23_7_xor1), .fa_or0(u_csamul_cla32_fa23_7_or0));
  and_gate and_gate_u_csamul_cla32_and24_7(.a(a[24]), .b(b[7]), .out(u_csamul_cla32_and24_7));
  fa fa_u_csamul_cla32_fa24_7_out(.a(u_csamul_cla32_and24_7[0]), .b(u_csamul_cla32_fa25_6_xor1[0]), .cin(u_csamul_cla32_fa24_6_or0[0]), .fa_xor1(u_csamul_cla32_fa24_7_xor1), .fa_or0(u_csamul_cla32_fa24_7_or0));
  and_gate and_gate_u_csamul_cla32_and25_7(.a(a[25]), .b(b[7]), .out(u_csamul_cla32_and25_7));
  fa fa_u_csamul_cla32_fa25_7_out(.a(u_csamul_cla32_and25_7[0]), .b(u_csamul_cla32_fa26_6_xor1[0]), .cin(u_csamul_cla32_fa25_6_or0[0]), .fa_xor1(u_csamul_cla32_fa25_7_xor1), .fa_or0(u_csamul_cla32_fa25_7_or0));
  and_gate and_gate_u_csamul_cla32_and26_7(.a(a[26]), .b(b[7]), .out(u_csamul_cla32_and26_7));
  fa fa_u_csamul_cla32_fa26_7_out(.a(u_csamul_cla32_and26_7[0]), .b(u_csamul_cla32_fa27_6_xor1[0]), .cin(u_csamul_cla32_fa26_6_or0[0]), .fa_xor1(u_csamul_cla32_fa26_7_xor1), .fa_or0(u_csamul_cla32_fa26_7_or0));
  and_gate and_gate_u_csamul_cla32_and27_7(.a(a[27]), .b(b[7]), .out(u_csamul_cla32_and27_7));
  fa fa_u_csamul_cla32_fa27_7_out(.a(u_csamul_cla32_and27_7[0]), .b(u_csamul_cla32_fa28_6_xor1[0]), .cin(u_csamul_cla32_fa27_6_or0[0]), .fa_xor1(u_csamul_cla32_fa27_7_xor1), .fa_or0(u_csamul_cla32_fa27_7_or0));
  and_gate and_gate_u_csamul_cla32_and28_7(.a(a[28]), .b(b[7]), .out(u_csamul_cla32_and28_7));
  fa fa_u_csamul_cla32_fa28_7_out(.a(u_csamul_cla32_and28_7[0]), .b(u_csamul_cla32_fa29_6_xor1[0]), .cin(u_csamul_cla32_fa28_6_or0[0]), .fa_xor1(u_csamul_cla32_fa28_7_xor1), .fa_or0(u_csamul_cla32_fa28_7_or0));
  and_gate and_gate_u_csamul_cla32_and29_7(.a(a[29]), .b(b[7]), .out(u_csamul_cla32_and29_7));
  fa fa_u_csamul_cla32_fa29_7_out(.a(u_csamul_cla32_and29_7[0]), .b(u_csamul_cla32_fa30_6_xor1[0]), .cin(u_csamul_cla32_fa29_6_or0[0]), .fa_xor1(u_csamul_cla32_fa29_7_xor1), .fa_or0(u_csamul_cla32_fa29_7_or0));
  and_gate and_gate_u_csamul_cla32_and30_7(.a(a[30]), .b(b[7]), .out(u_csamul_cla32_and30_7));
  fa fa_u_csamul_cla32_fa30_7_out(.a(u_csamul_cla32_and30_7[0]), .b(u_csamul_cla32_and31_6[0]), .cin(u_csamul_cla32_fa30_6_or0[0]), .fa_xor1(u_csamul_cla32_fa30_7_xor1), .fa_or0(u_csamul_cla32_fa30_7_or0));
  and_gate and_gate_u_csamul_cla32_and31_7(.a(a[31]), .b(b[7]), .out(u_csamul_cla32_and31_7));
  and_gate and_gate_u_csamul_cla32_and0_8(.a(a[0]), .b(b[8]), .out(u_csamul_cla32_and0_8));
  fa fa_u_csamul_cla32_fa0_8_out(.a(u_csamul_cla32_and0_8[0]), .b(u_csamul_cla32_fa1_7_xor1[0]), .cin(u_csamul_cla32_fa0_7_or0[0]), .fa_xor1(u_csamul_cla32_fa0_8_xor1), .fa_or0(u_csamul_cla32_fa0_8_or0));
  and_gate and_gate_u_csamul_cla32_and1_8(.a(a[1]), .b(b[8]), .out(u_csamul_cla32_and1_8));
  fa fa_u_csamul_cla32_fa1_8_out(.a(u_csamul_cla32_and1_8[0]), .b(u_csamul_cla32_fa2_7_xor1[0]), .cin(u_csamul_cla32_fa1_7_or0[0]), .fa_xor1(u_csamul_cla32_fa1_8_xor1), .fa_or0(u_csamul_cla32_fa1_8_or0));
  and_gate and_gate_u_csamul_cla32_and2_8(.a(a[2]), .b(b[8]), .out(u_csamul_cla32_and2_8));
  fa fa_u_csamul_cla32_fa2_8_out(.a(u_csamul_cla32_and2_8[0]), .b(u_csamul_cla32_fa3_7_xor1[0]), .cin(u_csamul_cla32_fa2_7_or0[0]), .fa_xor1(u_csamul_cla32_fa2_8_xor1), .fa_or0(u_csamul_cla32_fa2_8_or0));
  and_gate and_gate_u_csamul_cla32_and3_8(.a(a[3]), .b(b[8]), .out(u_csamul_cla32_and3_8));
  fa fa_u_csamul_cla32_fa3_8_out(.a(u_csamul_cla32_and3_8[0]), .b(u_csamul_cla32_fa4_7_xor1[0]), .cin(u_csamul_cla32_fa3_7_or0[0]), .fa_xor1(u_csamul_cla32_fa3_8_xor1), .fa_or0(u_csamul_cla32_fa3_8_or0));
  and_gate and_gate_u_csamul_cla32_and4_8(.a(a[4]), .b(b[8]), .out(u_csamul_cla32_and4_8));
  fa fa_u_csamul_cla32_fa4_8_out(.a(u_csamul_cla32_and4_8[0]), .b(u_csamul_cla32_fa5_7_xor1[0]), .cin(u_csamul_cla32_fa4_7_or0[0]), .fa_xor1(u_csamul_cla32_fa4_8_xor1), .fa_or0(u_csamul_cla32_fa4_8_or0));
  and_gate and_gate_u_csamul_cla32_and5_8(.a(a[5]), .b(b[8]), .out(u_csamul_cla32_and5_8));
  fa fa_u_csamul_cla32_fa5_8_out(.a(u_csamul_cla32_and5_8[0]), .b(u_csamul_cla32_fa6_7_xor1[0]), .cin(u_csamul_cla32_fa5_7_or0[0]), .fa_xor1(u_csamul_cla32_fa5_8_xor1), .fa_or0(u_csamul_cla32_fa5_8_or0));
  and_gate and_gate_u_csamul_cla32_and6_8(.a(a[6]), .b(b[8]), .out(u_csamul_cla32_and6_8));
  fa fa_u_csamul_cla32_fa6_8_out(.a(u_csamul_cla32_and6_8[0]), .b(u_csamul_cla32_fa7_7_xor1[0]), .cin(u_csamul_cla32_fa6_7_or0[0]), .fa_xor1(u_csamul_cla32_fa6_8_xor1), .fa_or0(u_csamul_cla32_fa6_8_or0));
  and_gate and_gate_u_csamul_cla32_and7_8(.a(a[7]), .b(b[8]), .out(u_csamul_cla32_and7_8));
  fa fa_u_csamul_cla32_fa7_8_out(.a(u_csamul_cla32_and7_8[0]), .b(u_csamul_cla32_fa8_7_xor1[0]), .cin(u_csamul_cla32_fa7_7_or0[0]), .fa_xor1(u_csamul_cla32_fa7_8_xor1), .fa_or0(u_csamul_cla32_fa7_8_or0));
  and_gate and_gate_u_csamul_cla32_and8_8(.a(a[8]), .b(b[8]), .out(u_csamul_cla32_and8_8));
  fa fa_u_csamul_cla32_fa8_8_out(.a(u_csamul_cla32_and8_8[0]), .b(u_csamul_cla32_fa9_7_xor1[0]), .cin(u_csamul_cla32_fa8_7_or0[0]), .fa_xor1(u_csamul_cla32_fa8_8_xor1), .fa_or0(u_csamul_cla32_fa8_8_or0));
  and_gate and_gate_u_csamul_cla32_and9_8(.a(a[9]), .b(b[8]), .out(u_csamul_cla32_and9_8));
  fa fa_u_csamul_cla32_fa9_8_out(.a(u_csamul_cla32_and9_8[0]), .b(u_csamul_cla32_fa10_7_xor1[0]), .cin(u_csamul_cla32_fa9_7_or0[0]), .fa_xor1(u_csamul_cla32_fa9_8_xor1), .fa_or0(u_csamul_cla32_fa9_8_or0));
  and_gate and_gate_u_csamul_cla32_and10_8(.a(a[10]), .b(b[8]), .out(u_csamul_cla32_and10_8));
  fa fa_u_csamul_cla32_fa10_8_out(.a(u_csamul_cla32_and10_8[0]), .b(u_csamul_cla32_fa11_7_xor1[0]), .cin(u_csamul_cla32_fa10_7_or0[0]), .fa_xor1(u_csamul_cla32_fa10_8_xor1), .fa_or0(u_csamul_cla32_fa10_8_or0));
  and_gate and_gate_u_csamul_cla32_and11_8(.a(a[11]), .b(b[8]), .out(u_csamul_cla32_and11_8));
  fa fa_u_csamul_cla32_fa11_8_out(.a(u_csamul_cla32_and11_8[0]), .b(u_csamul_cla32_fa12_7_xor1[0]), .cin(u_csamul_cla32_fa11_7_or0[0]), .fa_xor1(u_csamul_cla32_fa11_8_xor1), .fa_or0(u_csamul_cla32_fa11_8_or0));
  and_gate and_gate_u_csamul_cla32_and12_8(.a(a[12]), .b(b[8]), .out(u_csamul_cla32_and12_8));
  fa fa_u_csamul_cla32_fa12_8_out(.a(u_csamul_cla32_and12_8[0]), .b(u_csamul_cla32_fa13_7_xor1[0]), .cin(u_csamul_cla32_fa12_7_or0[0]), .fa_xor1(u_csamul_cla32_fa12_8_xor1), .fa_or0(u_csamul_cla32_fa12_8_or0));
  and_gate and_gate_u_csamul_cla32_and13_8(.a(a[13]), .b(b[8]), .out(u_csamul_cla32_and13_8));
  fa fa_u_csamul_cla32_fa13_8_out(.a(u_csamul_cla32_and13_8[0]), .b(u_csamul_cla32_fa14_7_xor1[0]), .cin(u_csamul_cla32_fa13_7_or0[0]), .fa_xor1(u_csamul_cla32_fa13_8_xor1), .fa_or0(u_csamul_cla32_fa13_8_or0));
  and_gate and_gate_u_csamul_cla32_and14_8(.a(a[14]), .b(b[8]), .out(u_csamul_cla32_and14_8));
  fa fa_u_csamul_cla32_fa14_8_out(.a(u_csamul_cla32_and14_8[0]), .b(u_csamul_cla32_fa15_7_xor1[0]), .cin(u_csamul_cla32_fa14_7_or0[0]), .fa_xor1(u_csamul_cla32_fa14_8_xor1), .fa_or0(u_csamul_cla32_fa14_8_or0));
  and_gate and_gate_u_csamul_cla32_and15_8(.a(a[15]), .b(b[8]), .out(u_csamul_cla32_and15_8));
  fa fa_u_csamul_cla32_fa15_8_out(.a(u_csamul_cla32_and15_8[0]), .b(u_csamul_cla32_fa16_7_xor1[0]), .cin(u_csamul_cla32_fa15_7_or0[0]), .fa_xor1(u_csamul_cla32_fa15_8_xor1), .fa_or0(u_csamul_cla32_fa15_8_or0));
  and_gate and_gate_u_csamul_cla32_and16_8(.a(a[16]), .b(b[8]), .out(u_csamul_cla32_and16_8));
  fa fa_u_csamul_cla32_fa16_8_out(.a(u_csamul_cla32_and16_8[0]), .b(u_csamul_cla32_fa17_7_xor1[0]), .cin(u_csamul_cla32_fa16_7_or0[0]), .fa_xor1(u_csamul_cla32_fa16_8_xor1), .fa_or0(u_csamul_cla32_fa16_8_or0));
  and_gate and_gate_u_csamul_cla32_and17_8(.a(a[17]), .b(b[8]), .out(u_csamul_cla32_and17_8));
  fa fa_u_csamul_cla32_fa17_8_out(.a(u_csamul_cla32_and17_8[0]), .b(u_csamul_cla32_fa18_7_xor1[0]), .cin(u_csamul_cla32_fa17_7_or0[0]), .fa_xor1(u_csamul_cla32_fa17_8_xor1), .fa_or0(u_csamul_cla32_fa17_8_or0));
  and_gate and_gate_u_csamul_cla32_and18_8(.a(a[18]), .b(b[8]), .out(u_csamul_cla32_and18_8));
  fa fa_u_csamul_cla32_fa18_8_out(.a(u_csamul_cla32_and18_8[0]), .b(u_csamul_cla32_fa19_7_xor1[0]), .cin(u_csamul_cla32_fa18_7_or0[0]), .fa_xor1(u_csamul_cla32_fa18_8_xor1), .fa_or0(u_csamul_cla32_fa18_8_or0));
  and_gate and_gate_u_csamul_cla32_and19_8(.a(a[19]), .b(b[8]), .out(u_csamul_cla32_and19_8));
  fa fa_u_csamul_cla32_fa19_8_out(.a(u_csamul_cla32_and19_8[0]), .b(u_csamul_cla32_fa20_7_xor1[0]), .cin(u_csamul_cla32_fa19_7_or0[0]), .fa_xor1(u_csamul_cla32_fa19_8_xor1), .fa_or0(u_csamul_cla32_fa19_8_or0));
  and_gate and_gate_u_csamul_cla32_and20_8(.a(a[20]), .b(b[8]), .out(u_csamul_cla32_and20_8));
  fa fa_u_csamul_cla32_fa20_8_out(.a(u_csamul_cla32_and20_8[0]), .b(u_csamul_cla32_fa21_7_xor1[0]), .cin(u_csamul_cla32_fa20_7_or0[0]), .fa_xor1(u_csamul_cla32_fa20_8_xor1), .fa_or0(u_csamul_cla32_fa20_8_or0));
  and_gate and_gate_u_csamul_cla32_and21_8(.a(a[21]), .b(b[8]), .out(u_csamul_cla32_and21_8));
  fa fa_u_csamul_cla32_fa21_8_out(.a(u_csamul_cla32_and21_8[0]), .b(u_csamul_cla32_fa22_7_xor1[0]), .cin(u_csamul_cla32_fa21_7_or0[0]), .fa_xor1(u_csamul_cla32_fa21_8_xor1), .fa_or0(u_csamul_cla32_fa21_8_or0));
  and_gate and_gate_u_csamul_cla32_and22_8(.a(a[22]), .b(b[8]), .out(u_csamul_cla32_and22_8));
  fa fa_u_csamul_cla32_fa22_8_out(.a(u_csamul_cla32_and22_8[0]), .b(u_csamul_cla32_fa23_7_xor1[0]), .cin(u_csamul_cla32_fa22_7_or0[0]), .fa_xor1(u_csamul_cla32_fa22_8_xor1), .fa_or0(u_csamul_cla32_fa22_8_or0));
  and_gate and_gate_u_csamul_cla32_and23_8(.a(a[23]), .b(b[8]), .out(u_csamul_cla32_and23_8));
  fa fa_u_csamul_cla32_fa23_8_out(.a(u_csamul_cla32_and23_8[0]), .b(u_csamul_cla32_fa24_7_xor1[0]), .cin(u_csamul_cla32_fa23_7_or0[0]), .fa_xor1(u_csamul_cla32_fa23_8_xor1), .fa_or0(u_csamul_cla32_fa23_8_or0));
  and_gate and_gate_u_csamul_cla32_and24_8(.a(a[24]), .b(b[8]), .out(u_csamul_cla32_and24_8));
  fa fa_u_csamul_cla32_fa24_8_out(.a(u_csamul_cla32_and24_8[0]), .b(u_csamul_cla32_fa25_7_xor1[0]), .cin(u_csamul_cla32_fa24_7_or0[0]), .fa_xor1(u_csamul_cla32_fa24_8_xor1), .fa_or0(u_csamul_cla32_fa24_8_or0));
  and_gate and_gate_u_csamul_cla32_and25_8(.a(a[25]), .b(b[8]), .out(u_csamul_cla32_and25_8));
  fa fa_u_csamul_cla32_fa25_8_out(.a(u_csamul_cla32_and25_8[0]), .b(u_csamul_cla32_fa26_7_xor1[0]), .cin(u_csamul_cla32_fa25_7_or0[0]), .fa_xor1(u_csamul_cla32_fa25_8_xor1), .fa_or0(u_csamul_cla32_fa25_8_or0));
  and_gate and_gate_u_csamul_cla32_and26_8(.a(a[26]), .b(b[8]), .out(u_csamul_cla32_and26_8));
  fa fa_u_csamul_cla32_fa26_8_out(.a(u_csamul_cla32_and26_8[0]), .b(u_csamul_cla32_fa27_7_xor1[0]), .cin(u_csamul_cla32_fa26_7_or0[0]), .fa_xor1(u_csamul_cla32_fa26_8_xor1), .fa_or0(u_csamul_cla32_fa26_8_or0));
  and_gate and_gate_u_csamul_cla32_and27_8(.a(a[27]), .b(b[8]), .out(u_csamul_cla32_and27_8));
  fa fa_u_csamul_cla32_fa27_8_out(.a(u_csamul_cla32_and27_8[0]), .b(u_csamul_cla32_fa28_7_xor1[0]), .cin(u_csamul_cla32_fa27_7_or0[0]), .fa_xor1(u_csamul_cla32_fa27_8_xor1), .fa_or0(u_csamul_cla32_fa27_8_or0));
  and_gate and_gate_u_csamul_cla32_and28_8(.a(a[28]), .b(b[8]), .out(u_csamul_cla32_and28_8));
  fa fa_u_csamul_cla32_fa28_8_out(.a(u_csamul_cla32_and28_8[0]), .b(u_csamul_cla32_fa29_7_xor1[0]), .cin(u_csamul_cla32_fa28_7_or0[0]), .fa_xor1(u_csamul_cla32_fa28_8_xor1), .fa_or0(u_csamul_cla32_fa28_8_or0));
  and_gate and_gate_u_csamul_cla32_and29_8(.a(a[29]), .b(b[8]), .out(u_csamul_cla32_and29_8));
  fa fa_u_csamul_cla32_fa29_8_out(.a(u_csamul_cla32_and29_8[0]), .b(u_csamul_cla32_fa30_7_xor1[0]), .cin(u_csamul_cla32_fa29_7_or0[0]), .fa_xor1(u_csamul_cla32_fa29_8_xor1), .fa_or0(u_csamul_cla32_fa29_8_or0));
  and_gate and_gate_u_csamul_cla32_and30_8(.a(a[30]), .b(b[8]), .out(u_csamul_cla32_and30_8));
  fa fa_u_csamul_cla32_fa30_8_out(.a(u_csamul_cla32_and30_8[0]), .b(u_csamul_cla32_and31_7[0]), .cin(u_csamul_cla32_fa30_7_or0[0]), .fa_xor1(u_csamul_cla32_fa30_8_xor1), .fa_or0(u_csamul_cla32_fa30_8_or0));
  and_gate and_gate_u_csamul_cla32_and31_8(.a(a[31]), .b(b[8]), .out(u_csamul_cla32_and31_8));
  and_gate and_gate_u_csamul_cla32_and0_9(.a(a[0]), .b(b[9]), .out(u_csamul_cla32_and0_9));
  fa fa_u_csamul_cla32_fa0_9_out(.a(u_csamul_cla32_and0_9[0]), .b(u_csamul_cla32_fa1_8_xor1[0]), .cin(u_csamul_cla32_fa0_8_or0[0]), .fa_xor1(u_csamul_cla32_fa0_9_xor1), .fa_or0(u_csamul_cla32_fa0_9_or0));
  and_gate and_gate_u_csamul_cla32_and1_9(.a(a[1]), .b(b[9]), .out(u_csamul_cla32_and1_9));
  fa fa_u_csamul_cla32_fa1_9_out(.a(u_csamul_cla32_and1_9[0]), .b(u_csamul_cla32_fa2_8_xor1[0]), .cin(u_csamul_cla32_fa1_8_or0[0]), .fa_xor1(u_csamul_cla32_fa1_9_xor1), .fa_or0(u_csamul_cla32_fa1_9_or0));
  and_gate and_gate_u_csamul_cla32_and2_9(.a(a[2]), .b(b[9]), .out(u_csamul_cla32_and2_9));
  fa fa_u_csamul_cla32_fa2_9_out(.a(u_csamul_cla32_and2_9[0]), .b(u_csamul_cla32_fa3_8_xor1[0]), .cin(u_csamul_cla32_fa2_8_or0[0]), .fa_xor1(u_csamul_cla32_fa2_9_xor1), .fa_or0(u_csamul_cla32_fa2_9_or0));
  and_gate and_gate_u_csamul_cla32_and3_9(.a(a[3]), .b(b[9]), .out(u_csamul_cla32_and3_9));
  fa fa_u_csamul_cla32_fa3_9_out(.a(u_csamul_cla32_and3_9[0]), .b(u_csamul_cla32_fa4_8_xor1[0]), .cin(u_csamul_cla32_fa3_8_or0[0]), .fa_xor1(u_csamul_cla32_fa3_9_xor1), .fa_or0(u_csamul_cla32_fa3_9_or0));
  and_gate and_gate_u_csamul_cla32_and4_9(.a(a[4]), .b(b[9]), .out(u_csamul_cla32_and4_9));
  fa fa_u_csamul_cla32_fa4_9_out(.a(u_csamul_cla32_and4_9[0]), .b(u_csamul_cla32_fa5_8_xor1[0]), .cin(u_csamul_cla32_fa4_8_or0[0]), .fa_xor1(u_csamul_cla32_fa4_9_xor1), .fa_or0(u_csamul_cla32_fa4_9_or0));
  and_gate and_gate_u_csamul_cla32_and5_9(.a(a[5]), .b(b[9]), .out(u_csamul_cla32_and5_9));
  fa fa_u_csamul_cla32_fa5_9_out(.a(u_csamul_cla32_and5_9[0]), .b(u_csamul_cla32_fa6_8_xor1[0]), .cin(u_csamul_cla32_fa5_8_or0[0]), .fa_xor1(u_csamul_cla32_fa5_9_xor1), .fa_or0(u_csamul_cla32_fa5_9_or0));
  and_gate and_gate_u_csamul_cla32_and6_9(.a(a[6]), .b(b[9]), .out(u_csamul_cla32_and6_9));
  fa fa_u_csamul_cla32_fa6_9_out(.a(u_csamul_cla32_and6_9[0]), .b(u_csamul_cla32_fa7_8_xor1[0]), .cin(u_csamul_cla32_fa6_8_or0[0]), .fa_xor1(u_csamul_cla32_fa6_9_xor1), .fa_or0(u_csamul_cla32_fa6_9_or0));
  and_gate and_gate_u_csamul_cla32_and7_9(.a(a[7]), .b(b[9]), .out(u_csamul_cla32_and7_9));
  fa fa_u_csamul_cla32_fa7_9_out(.a(u_csamul_cla32_and7_9[0]), .b(u_csamul_cla32_fa8_8_xor1[0]), .cin(u_csamul_cla32_fa7_8_or0[0]), .fa_xor1(u_csamul_cla32_fa7_9_xor1), .fa_or0(u_csamul_cla32_fa7_9_or0));
  and_gate and_gate_u_csamul_cla32_and8_9(.a(a[8]), .b(b[9]), .out(u_csamul_cla32_and8_9));
  fa fa_u_csamul_cla32_fa8_9_out(.a(u_csamul_cla32_and8_9[0]), .b(u_csamul_cla32_fa9_8_xor1[0]), .cin(u_csamul_cla32_fa8_8_or0[0]), .fa_xor1(u_csamul_cla32_fa8_9_xor1), .fa_or0(u_csamul_cla32_fa8_9_or0));
  and_gate and_gate_u_csamul_cla32_and9_9(.a(a[9]), .b(b[9]), .out(u_csamul_cla32_and9_9));
  fa fa_u_csamul_cla32_fa9_9_out(.a(u_csamul_cla32_and9_9[0]), .b(u_csamul_cla32_fa10_8_xor1[0]), .cin(u_csamul_cla32_fa9_8_or0[0]), .fa_xor1(u_csamul_cla32_fa9_9_xor1), .fa_or0(u_csamul_cla32_fa9_9_or0));
  and_gate and_gate_u_csamul_cla32_and10_9(.a(a[10]), .b(b[9]), .out(u_csamul_cla32_and10_9));
  fa fa_u_csamul_cla32_fa10_9_out(.a(u_csamul_cla32_and10_9[0]), .b(u_csamul_cla32_fa11_8_xor1[0]), .cin(u_csamul_cla32_fa10_8_or0[0]), .fa_xor1(u_csamul_cla32_fa10_9_xor1), .fa_or0(u_csamul_cla32_fa10_9_or0));
  and_gate and_gate_u_csamul_cla32_and11_9(.a(a[11]), .b(b[9]), .out(u_csamul_cla32_and11_9));
  fa fa_u_csamul_cla32_fa11_9_out(.a(u_csamul_cla32_and11_9[0]), .b(u_csamul_cla32_fa12_8_xor1[0]), .cin(u_csamul_cla32_fa11_8_or0[0]), .fa_xor1(u_csamul_cla32_fa11_9_xor1), .fa_or0(u_csamul_cla32_fa11_9_or0));
  and_gate and_gate_u_csamul_cla32_and12_9(.a(a[12]), .b(b[9]), .out(u_csamul_cla32_and12_9));
  fa fa_u_csamul_cla32_fa12_9_out(.a(u_csamul_cla32_and12_9[0]), .b(u_csamul_cla32_fa13_8_xor1[0]), .cin(u_csamul_cla32_fa12_8_or0[0]), .fa_xor1(u_csamul_cla32_fa12_9_xor1), .fa_or0(u_csamul_cla32_fa12_9_or0));
  and_gate and_gate_u_csamul_cla32_and13_9(.a(a[13]), .b(b[9]), .out(u_csamul_cla32_and13_9));
  fa fa_u_csamul_cla32_fa13_9_out(.a(u_csamul_cla32_and13_9[0]), .b(u_csamul_cla32_fa14_8_xor1[0]), .cin(u_csamul_cla32_fa13_8_or0[0]), .fa_xor1(u_csamul_cla32_fa13_9_xor1), .fa_or0(u_csamul_cla32_fa13_9_or0));
  and_gate and_gate_u_csamul_cla32_and14_9(.a(a[14]), .b(b[9]), .out(u_csamul_cla32_and14_9));
  fa fa_u_csamul_cla32_fa14_9_out(.a(u_csamul_cla32_and14_9[0]), .b(u_csamul_cla32_fa15_8_xor1[0]), .cin(u_csamul_cla32_fa14_8_or0[0]), .fa_xor1(u_csamul_cla32_fa14_9_xor1), .fa_or0(u_csamul_cla32_fa14_9_or0));
  and_gate and_gate_u_csamul_cla32_and15_9(.a(a[15]), .b(b[9]), .out(u_csamul_cla32_and15_9));
  fa fa_u_csamul_cla32_fa15_9_out(.a(u_csamul_cla32_and15_9[0]), .b(u_csamul_cla32_fa16_8_xor1[0]), .cin(u_csamul_cla32_fa15_8_or0[0]), .fa_xor1(u_csamul_cla32_fa15_9_xor1), .fa_or0(u_csamul_cla32_fa15_9_or0));
  and_gate and_gate_u_csamul_cla32_and16_9(.a(a[16]), .b(b[9]), .out(u_csamul_cla32_and16_9));
  fa fa_u_csamul_cla32_fa16_9_out(.a(u_csamul_cla32_and16_9[0]), .b(u_csamul_cla32_fa17_8_xor1[0]), .cin(u_csamul_cla32_fa16_8_or0[0]), .fa_xor1(u_csamul_cla32_fa16_9_xor1), .fa_or0(u_csamul_cla32_fa16_9_or0));
  and_gate and_gate_u_csamul_cla32_and17_9(.a(a[17]), .b(b[9]), .out(u_csamul_cla32_and17_9));
  fa fa_u_csamul_cla32_fa17_9_out(.a(u_csamul_cla32_and17_9[0]), .b(u_csamul_cla32_fa18_8_xor1[0]), .cin(u_csamul_cla32_fa17_8_or0[0]), .fa_xor1(u_csamul_cla32_fa17_9_xor1), .fa_or0(u_csamul_cla32_fa17_9_or0));
  and_gate and_gate_u_csamul_cla32_and18_9(.a(a[18]), .b(b[9]), .out(u_csamul_cla32_and18_9));
  fa fa_u_csamul_cla32_fa18_9_out(.a(u_csamul_cla32_and18_9[0]), .b(u_csamul_cla32_fa19_8_xor1[0]), .cin(u_csamul_cla32_fa18_8_or0[0]), .fa_xor1(u_csamul_cla32_fa18_9_xor1), .fa_or0(u_csamul_cla32_fa18_9_or0));
  and_gate and_gate_u_csamul_cla32_and19_9(.a(a[19]), .b(b[9]), .out(u_csamul_cla32_and19_9));
  fa fa_u_csamul_cla32_fa19_9_out(.a(u_csamul_cla32_and19_9[0]), .b(u_csamul_cla32_fa20_8_xor1[0]), .cin(u_csamul_cla32_fa19_8_or0[0]), .fa_xor1(u_csamul_cla32_fa19_9_xor1), .fa_or0(u_csamul_cla32_fa19_9_or0));
  and_gate and_gate_u_csamul_cla32_and20_9(.a(a[20]), .b(b[9]), .out(u_csamul_cla32_and20_9));
  fa fa_u_csamul_cla32_fa20_9_out(.a(u_csamul_cla32_and20_9[0]), .b(u_csamul_cla32_fa21_8_xor1[0]), .cin(u_csamul_cla32_fa20_8_or0[0]), .fa_xor1(u_csamul_cla32_fa20_9_xor1), .fa_or0(u_csamul_cla32_fa20_9_or0));
  and_gate and_gate_u_csamul_cla32_and21_9(.a(a[21]), .b(b[9]), .out(u_csamul_cla32_and21_9));
  fa fa_u_csamul_cla32_fa21_9_out(.a(u_csamul_cla32_and21_9[0]), .b(u_csamul_cla32_fa22_8_xor1[0]), .cin(u_csamul_cla32_fa21_8_or0[0]), .fa_xor1(u_csamul_cla32_fa21_9_xor1), .fa_or0(u_csamul_cla32_fa21_9_or0));
  and_gate and_gate_u_csamul_cla32_and22_9(.a(a[22]), .b(b[9]), .out(u_csamul_cla32_and22_9));
  fa fa_u_csamul_cla32_fa22_9_out(.a(u_csamul_cla32_and22_9[0]), .b(u_csamul_cla32_fa23_8_xor1[0]), .cin(u_csamul_cla32_fa22_8_or0[0]), .fa_xor1(u_csamul_cla32_fa22_9_xor1), .fa_or0(u_csamul_cla32_fa22_9_or0));
  and_gate and_gate_u_csamul_cla32_and23_9(.a(a[23]), .b(b[9]), .out(u_csamul_cla32_and23_9));
  fa fa_u_csamul_cla32_fa23_9_out(.a(u_csamul_cla32_and23_9[0]), .b(u_csamul_cla32_fa24_8_xor1[0]), .cin(u_csamul_cla32_fa23_8_or0[0]), .fa_xor1(u_csamul_cla32_fa23_9_xor1), .fa_or0(u_csamul_cla32_fa23_9_or0));
  and_gate and_gate_u_csamul_cla32_and24_9(.a(a[24]), .b(b[9]), .out(u_csamul_cla32_and24_9));
  fa fa_u_csamul_cla32_fa24_9_out(.a(u_csamul_cla32_and24_9[0]), .b(u_csamul_cla32_fa25_8_xor1[0]), .cin(u_csamul_cla32_fa24_8_or0[0]), .fa_xor1(u_csamul_cla32_fa24_9_xor1), .fa_or0(u_csamul_cla32_fa24_9_or0));
  and_gate and_gate_u_csamul_cla32_and25_9(.a(a[25]), .b(b[9]), .out(u_csamul_cla32_and25_9));
  fa fa_u_csamul_cla32_fa25_9_out(.a(u_csamul_cla32_and25_9[0]), .b(u_csamul_cla32_fa26_8_xor1[0]), .cin(u_csamul_cla32_fa25_8_or0[0]), .fa_xor1(u_csamul_cla32_fa25_9_xor1), .fa_or0(u_csamul_cla32_fa25_9_or0));
  and_gate and_gate_u_csamul_cla32_and26_9(.a(a[26]), .b(b[9]), .out(u_csamul_cla32_and26_9));
  fa fa_u_csamul_cla32_fa26_9_out(.a(u_csamul_cla32_and26_9[0]), .b(u_csamul_cla32_fa27_8_xor1[0]), .cin(u_csamul_cla32_fa26_8_or0[0]), .fa_xor1(u_csamul_cla32_fa26_9_xor1), .fa_or0(u_csamul_cla32_fa26_9_or0));
  and_gate and_gate_u_csamul_cla32_and27_9(.a(a[27]), .b(b[9]), .out(u_csamul_cla32_and27_9));
  fa fa_u_csamul_cla32_fa27_9_out(.a(u_csamul_cla32_and27_9[0]), .b(u_csamul_cla32_fa28_8_xor1[0]), .cin(u_csamul_cla32_fa27_8_or0[0]), .fa_xor1(u_csamul_cla32_fa27_9_xor1), .fa_or0(u_csamul_cla32_fa27_9_or0));
  and_gate and_gate_u_csamul_cla32_and28_9(.a(a[28]), .b(b[9]), .out(u_csamul_cla32_and28_9));
  fa fa_u_csamul_cla32_fa28_9_out(.a(u_csamul_cla32_and28_9[0]), .b(u_csamul_cla32_fa29_8_xor1[0]), .cin(u_csamul_cla32_fa28_8_or0[0]), .fa_xor1(u_csamul_cla32_fa28_9_xor1), .fa_or0(u_csamul_cla32_fa28_9_or0));
  and_gate and_gate_u_csamul_cla32_and29_9(.a(a[29]), .b(b[9]), .out(u_csamul_cla32_and29_9));
  fa fa_u_csamul_cla32_fa29_9_out(.a(u_csamul_cla32_and29_9[0]), .b(u_csamul_cla32_fa30_8_xor1[0]), .cin(u_csamul_cla32_fa29_8_or0[0]), .fa_xor1(u_csamul_cla32_fa29_9_xor1), .fa_or0(u_csamul_cla32_fa29_9_or0));
  and_gate and_gate_u_csamul_cla32_and30_9(.a(a[30]), .b(b[9]), .out(u_csamul_cla32_and30_9));
  fa fa_u_csamul_cla32_fa30_9_out(.a(u_csamul_cla32_and30_9[0]), .b(u_csamul_cla32_and31_8[0]), .cin(u_csamul_cla32_fa30_8_or0[0]), .fa_xor1(u_csamul_cla32_fa30_9_xor1), .fa_or0(u_csamul_cla32_fa30_9_or0));
  and_gate and_gate_u_csamul_cla32_and31_9(.a(a[31]), .b(b[9]), .out(u_csamul_cla32_and31_9));
  and_gate and_gate_u_csamul_cla32_and0_10(.a(a[0]), .b(b[10]), .out(u_csamul_cla32_and0_10));
  fa fa_u_csamul_cla32_fa0_10_out(.a(u_csamul_cla32_and0_10[0]), .b(u_csamul_cla32_fa1_9_xor1[0]), .cin(u_csamul_cla32_fa0_9_or0[0]), .fa_xor1(u_csamul_cla32_fa0_10_xor1), .fa_or0(u_csamul_cla32_fa0_10_or0));
  and_gate and_gate_u_csamul_cla32_and1_10(.a(a[1]), .b(b[10]), .out(u_csamul_cla32_and1_10));
  fa fa_u_csamul_cla32_fa1_10_out(.a(u_csamul_cla32_and1_10[0]), .b(u_csamul_cla32_fa2_9_xor1[0]), .cin(u_csamul_cla32_fa1_9_or0[0]), .fa_xor1(u_csamul_cla32_fa1_10_xor1), .fa_or0(u_csamul_cla32_fa1_10_or0));
  and_gate and_gate_u_csamul_cla32_and2_10(.a(a[2]), .b(b[10]), .out(u_csamul_cla32_and2_10));
  fa fa_u_csamul_cla32_fa2_10_out(.a(u_csamul_cla32_and2_10[0]), .b(u_csamul_cla32_fa3_9_xor1[0]), .cin(u_csamul_cla32_fa2_9_or0[0]), .fa_xor1(u_csamul_cla32_fa2_10_xor1), .fa_or0(u_csamul_cla32_fa2_10_or0));
  and_gate and_gate_u_csamul_cla32_and3_10(.a(a[3]), .b(b[10]), .out(u_csamul_cla32_and3_10));
  fa fa_u_csamul_cla32_fa3_10_out(.a(u_csamul_cla32_and3_10[0]), .b(u_csamul_cla32_fa4_9_xor1[0]), .cin(u_csamul_cla32_fa3_9_or0[0]), .fa_xor1(u_csamul_cla32_fa3_10_xor1), .fa_or0(u_csamul_cla32_fa3_10_or0));
  and_gate and_gate_u_csamul_cla32_and4_10(.a(a[4]), .b(b[10]), .out(u_csamul_cla32_and4_10));
  fa fa_u_csamul_cla32_fa4_10_out(.a(u_csamul_cla32_and4_10[0]), .b(u_csamul_cla32_fa5_9_xor1[0]), .cin(u_csamul_cla32_fa4_9_or0[0]), .fa_xor1(u_csamul_cla32_fa4_10_xor1), .fa_or0(u_csamul_cla32_fa4_10_or0));
  and_gate and_gate_u_csamul_cla32_and5_10(.a(a[5]), .b(b[10]), .out(u_csamul_cla32_and5_10));
  fa fa_u_csamul_cla32_fa5_10_out(.a(u_csamul_cla32_and5_10[0]), .b(u_csamul_cla32_fa6_9_xor1[0]), .cin(u_csamul_cla32_fa5_9_or0[0]), .fa_xor1(u_csamul_cla32_fa5_10_xor1), .fa_or0(u_csamul_cla32_fa5_10_or0));
  and_gate and_gate_u_csamul_cla32_and6_10(.a(a[6]), .b(b[10]), .out(u_csamul_cla32_and6_10));
  fa fa_u_csamul_cla32_fa6_10_out(.a(u_csamul_cla32_and6_10[0]), .b(u_csamul_cla32_fa7_9_xor1[0]), .cin(u_csamul_cla32_fa6_9_or0[0]), .fa_xor1(u_csamul_cla32_fa6_10_xor1), .fa_or0(u_csamul_cla32_fa6_10_or0));
  and_gate and_gate_u_csamul_cla32_and7_10(.a(a[7]), .b(b[10]), .out(u_csamul_cla32_and7_10));
  fa fa_u_csamul_cla32_fa7_10_out(.a(u_csamul_cla32_and7_10[0]), .b(u_csamul_cla32_fa8_9_xor1[0]), .cin(u_csamul_cla32_fa7_9_or0[0]), .fa_xor1(u_csamul_cla32_fa7_10_xor1), .fa_or0(u_csamul_cla32_fa7_10_or0));
  and_gate and_gate_u_csamul_cla32_and8_10(.a(a[8]), .b(b[10]), .out(u_csamul_cla32_and8_10));
  fa fa_u_csamul_cla32_fa8_10_out(.a(u_csamul_cla32_and8_10[0]), .b(u_csamul_cla32_fa9_9_xor1[0]), .cin(u_csamul_cla32_fa8_9_or0[0]), .fa_xor1(u_csamul_cla32_fa8_10_xor1), .fa_or0(u_csamul_cla32_fa8_10_or0));
  and_gate and_gate_u_csamul_cla32_and9_10(.a(a[9]), .b(b[10]), .out(u_csamul_cla32_and9_10));
  fa fa_u_csamul_cla32_fa9_10_out(.a(u_csamul_cla32_and9_10[0]), .b(u_csamul_cla32_fa10_9_xor1[0]), .cin(u_csamul_cla32_fa9_9_or0[0]), .fa_xor1(u_csamul_cla32_fa9_10_xor1), .fa_or0(u_csamul_cla32_fa9_10_or0));
  and_gate and_gate_u_csamul_cla32_and10_10(.a(a[10]), .b(b[10]), .out(u_csamul_cla32_and10_10));
  fa fa_u_csamul_cla32_fa10_10_out(.a(u_csamul_cla32_and10_10[0]), .b(u_csamul_cla32_fa11_9_xor1[0]), .cin(u_csamul_cla32_fa10_9_or0[0]), .fa_xor1(u_csamul_cla32_fa10_10_xor1), .fa_or0(u_csamul_cla32_fa10_10_or0));
  and_gate and_gate_u_csamul_cla32_and11_10(.a(a[11]), .b(b[10]), .out(u_csamul_cla32_and11_10));
  fa fa_u_csamul_cla32_fa11_10_out(.a(u_csamul_cla32_and11_10[0]), .b(u_csamul_cla32_fa12_9_xor1[0]), .cin(u_csamul_cla32_fa11_9_or0[0]), .fa_xor1(u_csamul_cla32_fa11_10_xor1), .fa_or0(u_csamul_cla32_fa11_10_or0));
  and_gate and_gate_u_csamul_cla32_and12_10(.a(a[12]), .b(b[10]), .out(u_csamul_cla32_and12_10));
  fa fa_u_csamul_cla32_fa12_10_out(.a(u_csamul_cla32_and12_10[0]), .b(u_csamul_cla32_fa13_9_xor1[0]), .cin(u_csamul_cla32_fa12_9_or0[0]), .fa_xor1(u_csamul_cla32_fa12_10_xor1), .fa_or0(u_csamul_cla32_fa12_10_or0));
  and_gate and_gate_u_csamul_cla32_and13_10(.a(a[13]), .b(b[10]), .out(u_csamul_cla32_and13_10));
  fa fa_u_csamul_cla32_fa13_10_out(.a(u_csamul_cla32_and13_10[0]), .b(u_csamul_cla32_fa14_9_xor1[0]), .cin(u_csamul_cla32_fa13_9_or0[0]), .fa_xor1(u_csamul_cla32_fa13_10_xor1), .fa_or0(u_csamul_cla32_fa13_10_or0));
  and_gate and_gate_u_csamul_cla32_and14_10(.a(a[14]), .b(b[10]), .out(u_csamul_cla32_and14_10));
  fa fa_u_csamul_cla32_fa14_10_out(.a(u_csamul_cla32_and14_10[0]), .b(u_csamul_cla32_fa15_9_xor1[0]), .cin(u_csamul_cla32_fa14_9_or0[0]), .fa_xor1(u_csamul_cla32_fa14_10_xor1), .fa_or0(u_csamul_cla32_fa14_10_or0));
  and_gate and_gate_u_csamul_cla32_and15_10(.a(a[15]), .b(b[10]), .out(u_csamul_cla32_and15_10));
  fa fa_u_csamul_cla32_fa15_10_out(.a(u_csamul_cla32_and15_10[0]), .b(u_csamul_cla32_fa16_9_xor1[0]), .cin(u_csamul_cla32_fa15_9_or0[0]), .fa_xor1(u_csamul_cla32_fa15_10_xor1), .fa_or0(u_csamul_cla32_fa15_10_or0));
  and_gate and_gate_u_csamul_cla32_and16_10(.a(a[16]), .b(b[10]), .out(u_csamul_cla32_and16_10));
  fa fa_u_csamul_cla32_fa16_10_out(.a(u_csamul_cla32_and16_10[0]), .b(u_csamul_cla32_fa17_9_xor1[0]), .cin(u_csamul_cla32_fa16_9_or0[0]), .fa_xor1(u_csamul_cla32_fa16_10_xor1), .fa_or0(u_csamul_cla32_fa16_10_or0));
  and_gate and_gate_u_csamul_cla32_and17_10(.a(a[17]), .b(b[10]), .out(u_csamul_cla32_and17_10));
  fa fa_u_csamul_cla32_fa17_10_out(.a(u_csamul_cla32_and17_10[0]), .b(u_csamul_cla32_fa18_9_xor1[0]), .cin(u_csamul_cla32_fa17_9_or0[0]), .fa_xor1(u_csamul_cla32_fa17_10_xor1), .fa_or0(u_csamul_cla32_fa17_10_or0));
  and_gate and_gate_u_csamul_cla32_and18_10(.a(a[18]), .b(b[10]), .out(u_csamul_cla32_and18_10));
  fa fa_u_csamul_cla32_fa18_10_out(.a(u_csamul_cla32_and18_10[0]), .b(u_csamul_cla32_fa19_9_xor1[0]), .cin(u_csamul_cla32_fa18_9_or0[0]), .fa_xor1(u_csamul_cla32_fa18_10_xor1), .fa_or0(u_csamul_cla32_fa18_10_or0));
  and_gate and_gate_u_csamul_cla32_and19_10(.a(a[19]), .b(b[10]), .out(u_csamul_cla32_and19_10));
  fa fa_u_csamul_cla32_fa19_10_out(.a(u_csamul_cla32_and19_10[0]), .b(u_csamul_cla32_fa20_9_xor1[0]), .cin(u_csamul_cla32_fa19_9_or0[0]), .fa_xor1(u_csamul_cla32_fa19_10_xor1), .fa_or0(u_csamul_cla32_fa19_10_or0));
  and_gate and_gate_u_csamul_cla32_and20_10(.a(a[20]), .b(b[10]), .out(u_csamul_cla32_and20_10));
  fa fa_u_csamul_cla32_fa20_10_out(.a(u_csamul_cla32_and20_10[0]), .b(u_csamul_cla32_fa21_9_xor1[0]), .cin(u_csamul_cla32_fa20_9_or0[0]), .fa_xor1(u_csamul_cla32_fa20_10_xor1), .fa_or0(u_csamul_cla32_fa20_10_or0));
  and_gate and_gate_u_csamul_cla32_and21_10(.a(a[21]), .b(b[10]), .out(u_csamul_cla32_and21_10));
  fa fa_u_csamul_cla32_fa21_10_out(.a(u_csamul_cla32_and21_10[0]), .b(u_csamul_cla32_fa22_9_xor1[0]), .cin(u_csamul_cla32_fa21_9_or0[0]), .fa_xor1(u_csamul_cla32_fa21_10_xor1), .fa_or0(u_csamul_cla32_fa21_10_or0));
  and_gate and_gate_u_csamul_cla32_and22_10(.a(a[22]), .b(b[10]), .out(u_csamul_cla32_and22_10));
  fa fa_u_csamul_cla32_fa22_10_out(.a(u_csamul_cla32_and22_10[0]), .b(u_csamul_cla32_fa23_9_xor1[0]), .cin(u_csamul_cla32_fa22_9_or0[0]), .fa_xor1(u_csamul_cla32_fa22_10_xor1), .fa_or0(u_csamul_cla32_fa22_10_or0));
  and_gate and_gate_u_csamul_cla32_and23_10(.a(a[23]), .b(b[10]), .out(u_csamul_cla32_and23_10));
  fa fa_u_csamul_cla32_fa23_10_out(.a(u_csamul_cla32_and23_10[0]), .b(u_csamul_cla32_fa24_9_xor1[0]), .cin(u_csamul_cla32_fa23_9_or0[0]), .fa_xor1(u_csamul_cla32_fa23_10_xor1), .fa_or0(u_csamul_cla32_fa23_10_or0));
  and_gate and_gate_u_csamul_cla32_and24_10(.a(a[24]), .b(b[10]), .out(u_csamul_cla32_and24_10));
  fa fa_u_csamul_cla32_fa24_10_out(.a(u_csamul_cla32_and24_10[0]), .b(u_csamul_cla32_fa25_9_xor1[0]), .cin(u_csamul_cla32_fa24_9_or0[0]), .fa_xor1(u_csamul_cla32_fa24_10_xor1), .fa_or0(u_csamul_cla32_fa24_10_or0));
  and_gate and_gate_u_csamul_cla32_and25_10(.a(a[25]), .b(b[10]), .out(u_csamul_cla32_and25_10));
  fa fa_u_csamul_cla32_fa25_10_out(.a(u_csamul_cla32_and25_10[0]), .b(u_csamul_cla32_fa26_9_xor1[0]), .cin(u_csamul_cla32_fa25_9_or0[0]), .fa_xor1(u_csamul_cla32_fa25_10_xor1), .fa_or0(u_csamul_cla32_fa25_10_or0));
  and_gate and_gate_u_csamul_cla32_and26_10(.a(a[26]), .b(b[10]), .out(u_csamul_cla32_and26_10));
  fa fa_u_csamul_cla32_fa26_10_out(.a(u_csamul_cla32_and26_10[0]), .b(u_csamul_cla32_fa27_9_xor1[0]), .cin(u_csamul_cla32_fa26_9_or0[0]), .fa_xor1(u_csamul_cla32_fa26_10_xor1), .fa_or0(u_csamul_cla32_fa26_10_or0));
  and_gate and_gate_u_csamul_cla32_and27_10(.a(a[27]), .b(b[10]), .out(u_csamul_cla32_and27_10));
  fa fa_u_csamul_cla32_fa27_10_out(.a(u_csamul_cla32_and27_10[0]), .b(u_csamul_cla32_fa28_9_xor1[0]), .cin(u_csamul_cla32_fa27_9_or0[0]), .fa_xor1(u_csamul_cla32_fa27_10_xor1), .fa_or0(u_csamul_cla32_fa27_10_or0));
  and_gate and_gate_u_csamul_cla32_and28_10(.a(a[28]), .b(b[10]), .out(u_csamul_cla32_and28_10));
  fa fa_u_csamul_cla32_fa28_10_out(.a(u_csamul_cla32_and28_10[0]), .b(u_csamul_cla32_fa29_9_xor1[0]), .cin(u_csamul_cla32_fa28_9_or0[0]), .fa_xor1(u_csamul_cla32_fa28_10_xor1), .fa_or0(u_csamul_cla32_fa28_10_or0));
  and_gate and_gate_u_csamul_cla32_and29_10(.a(a[29]), .b(b[10]), .out(u_csamul_cla32_and29_10));
  fa fa_u_csamul_cla32_fa29_10_out(.a(u_csamul_cla32_and29_10[0]), .b(u_csamul_cla32_fa30_9_xor1[0]), .cin(u_csamul_cla32_fa29_9_or0[0]), .fa_xor1(u_csamul_cla32_fa29_10_xor1), .fa_or0(u_csamul_cla32_fa29_10_or0));
  and_gate and_gate_u_csamul_cla32_and30_10(.a(a[30]), .b(b[10]), .out(u_csamul_cla32_and30_10));
  fa fa_u_csamul_cla32_fa30_10_out(.a(u_csamul_cla32_and30_10[0]), .b(u_csamul_cla32_and31_9[0]), .cin(u_csamul_cla32_fa30_9_or0[0]), .fa_xor1(u_csamul_cla32_fa30_10_xor1), .fa_or0(u_csamul_cla32_fa30_10_or0));
  and_gate and_gate_u_csamul_cla32_and31_10(.a(a[31]), .b(b[10]), .out(u_csamul_cla32_and31_10));
  and_gate and_gate_u_csamul_cla32_and0_11(.a(a[0]), .b(b[11]), .out(u_csamul_cla32_and0_11));
  fa fa_u_csamul_cla32_fa0_11_out(.a(u_csamul_cla32_and0_11[0]), .b(u_csamul_cla32_fa1_10_xor1[0]), .cin(u_csamul_cla32_fa0_10_or0[0]), .fa_xor1(u_csamul_cla32_fa0_11_xor1), .fa_or0(u_csamul_cla32_fa0_11_or0));
  and_gate and_gate_u_csamul_cla32_and1_11(.a(a[1]), .b(b[11]), .out(u_csamul_cla32_and1_11));
  fa fa_u_csamul_cla32_fa1_11_out(.a(u_csamul_cla32_and1_11[0]), .b(u_csamul_cla32_fa2_10_xor1[0]), .cin(u_csamul_cla32_fa1_10_or0[0]), .fa_xor1(u_csamul_cla32_fa1_11_xor1), .fa_or0(u_csamul_cla32_fa1_11_or0));
  and_gate and_gate_u_csamul_cla32_and2_11(.a(a[2]), .b(b[11]), .out(u_csamul_cla32_and2_11));
  fa fa_u_csamul_cla32_fa2_11_out(.a(u_csamul_cla32_and2_11[0]), .b(u_csamul_cla32_fa3_10_xor1[0]), .cin(u_csamul_cla32_fa2_10_or0[0]), .fa_xor1(u_csamul_cla32_fa2_11_xor1), .fa_or0(u_csamul_cla32_fa2_11_or0));
  and_gate and_gate_u_csamul_cla32_and3_11(.a(a[3]), .b(b[11]), .out(u_csamul_cla32_and3_11));
  fa fa_u_csamul_cla32_fa3_11_out(.a(u_csamul_cla32_and3_11[0]), .b(u_csamul_cla32_fa4_10_xor1[0]), .cin(u_csamul_cla32_fa3_10_or0[0]), .fa_xor1(u_csamul_cla32_fa3_11_xor1), .fa_or0(u_csamul_cla32_fa3_11_or0));
  and_gate and_gate_u_csamul_cla32_and4_11(.a(a[4]), .b(b[11]), .out(u_csamul_cla32_and4_11));
  fa fa_u_csamul_cla32_fa4_11_out(.a(u_csamul_cla32_and4_11[0]), .b(u_csamul_cla32_fa5_10_xor1[0]), .cin(u_csamul_cla32_fa4_10_or0[0]), .fa_xor1(u_csamul_cla32_fa4_11_xor1), .fa_or0(u_csamul_cla32_fa4_11_or0));
  and_gate and_gate_u_csamul_cla32_and5_11(.a(a[5]), .b(b[11]), .out(u_csamul_cla32_and5_11));
  fa fa_u_csamul_cla32_fa5_11_out(.a(u_csamul_cla32_and5_11[0]), .b(u_csamul_cla32_fa6_10_xor1[0]), .cin(u_csamul_cla32_fa5_10_or0[0]), .fa_xor1(u_csamul_cla32_fa5_11_xor1), .fa_or0(u_csamul_cla32_fa5_11_or0));
  and_gate and_gate_u_csamul_cla32_and6_11(.a(a[6]), .b(b[11]), .out(u_csamul_cla32_and6_11));
  fa fa_u_csamul_cla32_fa6_11_out(.a(u_csamul_cla32_and6_11[0]), .b(u_csamul_cla32_fa7_10_xor1[0]), .cin(u_csamul_cla32_fa6_10_or0[0]), .fa_xor1(u_csamul_cla32_fa6_11_xor1), .fa_or0(u_csamul_cla32_fa6_11_or0));
  and_gate and_gate_u_csamul_cla32_and7_11(.a(a[7]), .b(b[11]), .out(u_csamul_cla32_and7_11));
  fa fa_u_csamul_cla32_fa7_11_out(.a(u_csamul_cla32_and7_11[0]), .b(u_csamul_cla32_fa8_10_xor1[0]), .cin(u_csamul_cla32_fa7_10_or0[0]), .fa_xor1(u_csamul_cla32_fa7_11_xor1), .fa_or0(u_csamul_cla32_fa7_11_or0));
  and_gate and_gate_u_csamul_cla32_and8_11(.a(a[8]), .b(b[11]), .out(u_csamul_cla32_and8_11));
  fa fa_u_csamul_cla32_fa8_11_out(.a(u_csamul_cla32_and8_11[0]), .b(u_csamul_cla32_fa9_10_xor1[0]), .cin(u_csamul_cla32_fa8_10_or0[0]), .fa_xor1(u_csamul_cla32_fa8_11_xor1), .fa_or0(u_csamul_cla32_fa8_11_or0));
  and_gate and_gate_u_csamul_cla32_and9_11(.a(a[9]), .b(b[11]), .out(u_csamul_cla32_and9_11));
  fa fa_u_csamul_cla32_fa9_11_out(.a(u_csamul_cla32_and9_11[0]), .b(u_csamul_cla32_fa10_10_xor1[0]), .cin(u_csamul_cla32_fa9_10_or0[0]), .fa_xor1(u_csamul_cla32_fa9_11_xor1), .fa_or0(u_csamul_cla32_fa9_11_or0));
  and_gate and_gate_u_csamul_cla32_and10_11(.a(a[10]), .b(b[11]), .out(u_csamul_cla32_and10_11));
  fa fa_u_csamul_cla32_fa10_11_out(.a(u_csamul_cla32_and10_11[0]), .b(u_csamul_cla32_fa11_10_xor1[0]), .cin(u_csamul_cla32_fa10_10_or0[0]), .fa_xor1(u_csamul_cla32_fa10_11_xor1), .fa_or0(u_csamul_cla32_fa10_11_or0));
  and_gate and_gate_u_csamul_cla32_and11_11(.a(a[11]), .b(b[11]), .out(u_csamul_cla32_and11_11));
  fa fa_u_csamul_cla32_fa11_11_out(.a(u_csamul_cla32_and11_11[0]), .b(u_csamul_cla32_fa12_10_xor1[0]), .cin(u_csamul_cla32_fa11_10_or0[0]), .fa_xor1(u_csamul_cla32_fa11_11_xor1), .fa_or0(u_csamul_cla32_fa11_11_or0));
  and_gate and_gate_u_csamul_cla32_and12_11(.a(a[12]), .b(b[11]), .out(u_csamul_cla32_and12_11));
  fa fa_u_csamul_cla32_fa12_11_out(.a(u_csamul_cla32_and12_11[0]), .b(u_csamul_cla32_fa13_10_xor1[0]), .cin(u_csamul_cla32_fa12_10_or0[0]), .fa_xor1(u_csamul_cla32_fa12_11_xor1), .fa_or0(u_csamul_cla32_fa12_11_or0));
  and_gate and_gate_u_csamul_cla32_and13_11(.a(a[13]), .b(b[11]), .out(u_csamul_cla32_and13_11));
  fa fa_u_csamul_cla32_fa13_11_out(.a(u_csamul_cla32_and13_11[0]), .b(u_csamul_cla32_fa14_10_xor1[0]), .cin(u_csamul_cla32_fa13_10_or0[0]), .fa_xor1(u_csamul_cla32_fa13_11_xor1), .fa_or0(u_csamul_cla32_fa13_11_or0));
  and_gate and_gate_u_csamul_cla32_and14_11(.a(a[14]), .b(b[11]), .out(u_csamul_cla32_and14_11));
  fa fa_u_csamul_cla32_fa14_11_out(.a(u_csamul_cla32_and14_11[0]), .b(u_csamul_cla32_fa15_10_xor1[0]), .cin(u_csamul_cla32_fa14_10_or0[0]), .fa_xor1(u_csamul_cla32_fa14_11_xor1), .fa_or0(u_csamul_cla32_fa14_11_or0));
  and_gate and_gate_u_csamul_cla32_and15_11(.a(a[15]), .b(b[11]), .out(u_csamul_cla32_and15_11));
  fa fa_u_csamul_cla32_fa15_11_out(.a(u_csamul_cla32_and15_11[0]), .b(u_csamul_cla32_fa16_10_xor1[0]), .cin(u_csamul_cla32_fa15_10_or0[0]), .fa_xor1(u_csamul_cla32_fa15_11_xor1), .fa_or0(u_csamul_cla32_fa15_11_or0));
  and_gate and_gate_u_csamul_cla32_and16_11(.a(a[16]), .b(b[11]), .out(u_csamul_cla32_and16_11));
  fa fa_u_csamul_cla32_fa16_11_out(.a(u_csamul_cla32_and16_11[0]), .b(u_csamul_cla32_fa17_10_xor1[0]), .cin(u_csamul_cla32_fa16_10_or0[0]), .fa_xor1(u_csamul_cla32_fa16_11_xor1), .fa_or0(u_csamul_cla32_fa16_11_or0));
  and_gate and_gate_u_csamul_cla32_and17_11(.a(a[17]), .b(b[11]), .out(u_csamul_cla32_and17_11));
  fa fa_u_csamul_cla32_fa17_11_out(.a(u_csamul_cla32_and17_11[0]), .b(u_csamul_cla32_fa18_10_xor1[0]), .cin(u_csamul_cla32_fa17_10_or0[0]), .fa_xor1(u_csamul_cla32_fa17_11_xor1), .fa_or0(u_csamul_cla32_fa17_11_or0));
  and_gate and_gate_u_csamul_cla32_and18_11(.a(a[18]), .b(b[11]), .out(u_csamul_cla32_and18_11));
  fa fa_u_csamul_cla32_fa18_11_out(.a(u_csamul_cla32_and18_11[0]), .b(u_csamul_cla32_fa19_10_xor1[0]), .cin(u_csamul_cla32_fa18_10_or0[0]), .fa_xor1(u_csamul_cla32_fa18_11_xor1), .fa_or0(u_csamul_cla32_fa18_11_or0));
  and_gate and_gate_u_csamul_cla32_and19_11(.a(a[19]), .b(b[11]), .out(u_csamul_cla32_and19_11));
  fa fa_u_csamul_cla32_fa19_11_out(.a(u_csamul_cla32_and19_11[0]), .b(u_csamul_cla32_fa20_10_xor1[0]), .cin(u_csamul_cla32_fa19_10_or0[0]), .fa_xor1(u_csamul_cla32_fa19_11_xor1), .fa_or0(u_csamul_cla32_fa19_11_or0));
  and_gate and_gate_u_csamul_cla32_and20_11(.a(a[20]), .b(b[11]), .out(u_csamul_cla32_and20_11));
  fa fa_u_csamul_cla32_fa20_11_out(.a(u_csamul_cla32_and20_11[0]), .b(u_csamul_cla32_fa21_10_xor1[0]), .cin(u_csamul_cla32_fa20_10_or0[0]), .fa_xor1(u_csamul_cla32_fa20_11_xor1), .fa_or0(u_csamul_cla32_fa20_11_or0));
  and_gate and_gate_u_csamul_cla32_and21_11(.a(a[21]), .b(b[11]), .out(u_csamul_cla32_and21_11));
  fa fa_u_csamul_cla32_fa21_11_out(.a(u_csamul_cla32_and21_11[0]), .b(u_csamul_cla32_fa22_10_xor1[0]), .cin(u_csamul_cla32_fa21_10_or0[0]), .fa_xor1(u_csamul_cla32_fa21_11_xor1), .fa_or0(u_csamul_cla32_fa21_11_or0));
  and_gate and_gate_u_csamul_cla32_and22_11(.a(a[22]), .b(b[11]), .out(u_csamul_cla32_and22_11));
  fa fa_u_csamul_cla32_fa22_11_out(.a(u_csamul_cla32_and22_11[0]), .b(u_csamul_cla32_fa23_10_xor1[0]), .cin(u_csamul_cla32_fa22_10_or0[0]), .fa_xor1(u_csamul_cla32_fa22_11_xor1), .fa_or0(u_csamul_cla32_fa22_11_or0));
  and_gate and_gate_u_csamul_cla32_and23_11(.a(a[23]), .b(b[11]), .out(u_csamul_cla32_and23_11));
  fa fa_u_csamul_cla32_fa23_11_out(.a(u_csamul_cla32_and23_11[0]), .b(u_csamul_cla32_fa24_10_xor1[0]), .cin(u_csamul_cla32_fa23_10_or0[0]), .fa_xor1(u_csamul_cla32_fa23_11_xor1), .fa_or0(u_csamul_cla32_fa23_11_or0));
  and_gate and_gate_u_csamul_cla32_and24_11(.a(a[24]), .b(b[11]), .out(u_csamul_cla32_and24_11));
  fa fa_u_csamul_cla32_fa24_11_out(.a(u_csamul_cla32_and24_11[0]), .b(u_csamul_cla32_fa25_10_xor1[0]), .cin(u_csamul_cla32_fa24_10_or0[0]), .fa_xor1(u_csamul_cla32_fa24_11_xor1), .fa_or0(u_csamul_cla32_fa24_11_or0));
  and_gate and_gate_u_csamul_cla32_and25_11(.a(a[25]), .b(b[11]), .out(u_csamul_cla32_and25_11));
  fa fa_u_csamul_cla32_fa25_11_out(.a(u_csamul_cla32_and25_11[0]), .b(u_csamul_cla32_fa26_10_xor1[0]), .cin(u_csamul_cla32_fa25_10_or0[0]), .fa_xor1(u_csamul_cla32_fa25_11_xor1), .fa_or0(u_csamul_cla32_fa25_11_or0));
  and_gate and_gate_u_csamul_cla32_and26_11(.a(a[26]), .b(b[11]), .out(u_csamul_cla32_and26_11));
  fa fa_u_csamul_cla32_fa26_11_out(.a(u_csamul_cla32_and26_11[0]), .b(u_csamul_cla32_fa27_10_xor1[0]), .cin(u_csamul_cla32_fa26_10_or0[0]), .fa_xor1(u_csamul_cla32_fa26_11_xor1), .fa_or0(u_csamul_cla32_fa26_11_or0));
  and_gate and_gate_u_csamul_cla32_and27_11(.a(a[27]), .b(b[11]), .out(u_csamul_cla32_and27_11));
  fa fa_u_csamul_cla32_fa27_11_out(.a(u_csamul_cla32_and27_11[0]), .b(u_csamul_cla32_fa28_10_xor1[0]), .cin(u_csamul_cla32_fa27_10_or0[0]), .fa_xor1(u_csamul_cla32_fa27_11_xor1), .fa_or0(u_csamul_cla32_fa27_11_or0));
  and_gate and_gate_u_csamul_cla32_and28_11(.a(a[28]), .b(b[11]), .out(u_csamul_cla32_and28_11));
  fa fa_u_csamul_cla32_fa28_11_out(.a(u_csamul_cla32_and28_11[0]), .b(u_csamul_cla32_fa29_10_xor1[0]), .cin(u_csamul_cla32_fa28_10_or0[0]), .fa_xor1(u_csamul_cla32_fa28_11_xor1), .fa_or0(u_csamul_cla32_fa28_11_or0));
  and_gate and_gate_u_csamul_cla32_and29_11(.a(a[29]), .b(b[11]), .out(u_csamul_cla32_and29_11));
  fa fa_u_csamul_cla32_fa29_11_out(.a(u_csamul_cla32_and29_11[0]), .b(u_csamul_cla32_fa30_10_xor1[0]), .cin(u_csamul_cla32_fa29_10_or0[0]), .fa_xor1(u_csamul_cla32_fa29_11_xor1), .fa_or0(u_csamul_cla32_fa29_11_or0));
  and_gate and_gate_u_csamul_cla32_and30_11(.a(a[30]), .b(b[11]), .out(u_csamul_cla32_and30_11));
  fa fa_u_csamul_cla32_fa30_11_out(.a(u_csamul_cla32_and30_11[0]), .b(u_csamul_cla32_and31_10[0]), .cin(u_csamul_cla32_fa30_10_or0[0]), .fa_xor1(u_csamul_cla32_fa30_11_xor1), .fa_or0(u_csamul_cla32_fa30_11_or0));
  and_gate and_gate_u_csamul_cla32_and31_11(.a(a[31]), .b(b[11]), .out(u_csamul_cla32_and31_11));
  and_gate and_gate_u_csamul_cla32_and0_12(.a(a[0]), .b(b[12]), .out(u_csamul_cla32_and0_12));
  fa fa_u_csamul_cla32_fa0_12_out(.a(u_csamul_cla32_and0_12[0]), .b(u_csamul_cla32_fa1_11_xor1[0]), .cin(u_csamul_cla32_fa0_11_or0[0]), .fa_xor1(u_csamul_cla32_fa0_12_xor1), .fa_or0(u_csamul_cla32_fa0_12_or0));
  and_gate and_gate_u_csamul_cla32_and1_12(.a(a[1]), .b(b[12]), .out(u_csamul_cla32_and1_12));
  fa fa_u_csamul_cla32_fa1_12_out(.a(u_csamul_cla32_and1_12[0]), .b(u_csamul_cla32_fa2_11_xor1[0]), .cin(u_csamul_cla32_fa1_11_or0[0]), .fa_xor1(u_csamul_cla32_fa1_12_xor1), .fa_or0(u_csamul_cla32_fa1_12_or0));
  and_gate and_gate_u_csamul_cla32_and2_12(.a(a[2]), .b(b[12]), .out(u_csamul_cla32_and2_12));
  fa fa_u_csamul_cla32_fa2_12_out(.a(u_csamul_cla32_and2_12[0]), .b(u_csamul_cla32_fa3_11_xor1[0]), .cin(u_csamul_cla32_fa2_11_or0[0]), .fa_xor1(u_csamul_cla32_fa2_12_xor1), .fa_or0(u_csamul_cla32_fa2_12_or0));
  and_gate and_gate_u_csamul_cla32_and3_12(.a(a[3]), .b(b[12]), .out(u_csamul_cla32_and3_12));
  fa fa_u_csamul_cla32_fa3_12_out(.a(u_csamul_cla32_and3_12[0]), .b(u_csamul_cla32_fa4_11_xor1[0]), .cin(u_csamul_cla32_fa3_11_or0[0]), .fa_xor1(u_csamul_cla32_fa3_12_xor1), .fa_or0(u_csamul_cla32_fa3_12_or0));
  and_gate and_gate_u_csamul_cla32_and4_12(.a(a[4]), .b(b[12]), .out(u_csamul_cla32_and4_12));
  fa fa_u_csamul_cla32_fa4_12_out(.a(u_csamul_cla32_and4_12[0]), .b(u_csamul_cla32_fa5_11_xor1[0]), .cin(u_csamul_cla32_fa4_11_or0[0]), .fa_xor1(u_csamul_cla32_fa4_12_xor1), .fa_or0(u_csamul_cla32_fa4_12_or0));
  and_gate and_gate_u_csamul_cla32_and5_12(.a(a[5]), .b(b[12]), .out(u_csamul_cla32_and5_12));
  fa fa_u_csamul_cla32_fa5_12_out(.a(u_csamul_cla32_and5_12[0]), .b(u_csamul_cla32_fa6_11_xor1[0]), .cin(u_csamul_cla32_fa5_11_or0[0]), .fa_xor1(u_csamul_cla32_fa5_12_xor1), .fa_or0(u_csamul_cla32_fa5_12_or0));
  and_gate and_gate_u_csamul_cla32_and6_12(.a(a[6]), .b(b[12]), .out(u_csamul_cla32_and6_12));
  fa fa_u_csamul_cla32_fa6_12_out(.a(u_csamul_cla32_and6_12[0]), .b(u_csamul_cla32_fa7_11_xor1[0]), .cin(u_csamul_cla32_fa6_11_or0[0]), .fa_xor1(u_csamul_cla32_fa6_12_xor1), .fa_or0(u_csamul_cla32_fa6_12_or0));
  and_gate and_gate_u_csamul_cla32_and7_12(.a(a[7]), .b(b[12]), .out(u_csamul_cla32_and7_12));
  fa fa_u_csamul_cla32_fa7_12_out(.a(u_csamul_cla32_and7_12[0]), .b(u_csamul_cla32_fa8_11_xor1[0]), .cin(u_csamul_cla32_fa7_11_or0[0]), .fa_xor1(u_csamul_cla32_fa7_12_xor1), .fa_or0(u_csamul_cla32_fa7_12_or0));
  and_gate and_gate_u_csamul_cla32_and8_12(.a(a[8]), .b(b[12]), .out(u_csamul_cla32_and8_12));
  fa fa_u_csamul_cla32_fa8_12_out(.a(u_csamul_cla32_and8_12[0]), .b(u_csamul_cla32_fa9_11_xor1[0]), .cin(u_csamul_cla32_fa8_11_or0[0]), .fa_xor1(u_csamul_cla32_fa8_12_xor1), .fa_or0(u_csamul_cla32_fa8_12_or0));
  and_gate and_gate_u_csamul_cla32_and9_12(.a(a[9]), .b(b[12]), .out(u_csamul_cla32_and9_12));
  fa fa_u_csamul_cla32_fa9_12_out(.a(u_csamul_cla32_and9_12[0]), .b(u_csamul_cla32_fa10_11_xor1[0]), .cin(u_csamul_cla32_fa9_11_or0[0]), .fa_xor1(u_csamul_cla32_fa9_12_xor1), .fa_or0(u_csamul_cla32_fa9_12_or0));
  and_gate and_gate_u_csamul_cla32_and10_12(.a(a[10]), .b(b[12]), .out(u_csamul_cla32_and10_12));
  fa fa_u_csamul_cla32_fa10_12_out(.a(u_csamul_cla32_and10_12[0]), .b(u_csamul_cla32_fa11_11_xor1[0]), .cin(u_csamul_cla32_fa10_11_or0[0]), .fa_xor1(u_csamul_cla32_fa10_12_xor1), .fa_or0(u_csamul_cla32_fa10_12_or0));
  and_gate and_gate_u_csamul_cla32_and11_12(.a(a[11]), .b(b[12]), .out(u_csamul_cla32_and11_12));
  fa fa_u_csamul_cla32_fa11_12_out(.a(u_csamul_cla32_and11_12[0]), .b(u_csamul_cla32_fa12_11_xor1[0]), .cin(u_csamul_cla32_fa11_11_or0[0]), .fa_xor1(u_csamul_cla32_fa11_12_xor1), .fa_or0(u_csamul_cla32_fa11_12_or0));
  and_gate and_gate_u_csamul_cla32_and12_12(.a(a[12]), .b(b[12]), .out(u_csamul_cla32_and12_12));
  fa fa_u_csamul_cla32_fa12_12_out(.a(u_csamul_cla32_and12_12[0]), .b(u_csamul_cla32_fa13_11_xor1[0]), .cin(u_csamul_cla32_fa12_11_or0[0]), .fa_xor1(u_csamul_cla32_fa12_12_xor1), .fa_or0(u_csamul_cla32_fa12_12_or0));
  and_gate and_gate_u_csamul_cla32_and13_12(.a(a[13]), .b(b[12]), .out(u_csamul_cla32_and13_12));
  fa fa_u_csamul_cla32_fa13_12_out(.a(u_csamul_cla32_and13_12[0]), .b(u_csamul_cla32_fa14_11_xor1[0]), .cin(u_csamul_cla32_fa13_11_or0[0]), .fa_xor1(u_csamul_cla32_fa13_12_xor1), .fa_or0(u_csamul_cla32_fa13_12_or0));
  and_gate and_gate_u_csamul_cla32_and14_12(.a(a[14]), .b(b[12]), .out(u_csamul_cla32_and14_12));
  fa fa_u_csamul_cla32_fa14_12_out(.a(u_csamul_cla32_and14_12[0]), .b(u_csamul_cla32_fa15_11_xor1[0]), .cin(u_csamul_cla32_fa14_11_or0[0]), .fa_xor1(u_csamul_cla32_fa14_12_xor1), .fa_or0(u_csamul_cla32_fa14_12_or0));
  and_gate and_gate_u_csamul_cla32_and15_12(.a(a[15]), .b(b[12]), .out(u_csamul_cla32_and15_12));
  fa fa_u_csamul_cla32_fa15_12_out(.a(u_csamul_cla32_and15_12[0]), .b(u_csamul_cla32_fa16_11_xor1[0]), .cin(u_csamul_cla32_fa15_11_or0[0]), .fa_xor1(u_csamul_cla32_fa15_12_xor1), .fa_or0(u_csamul_cla32_fa15_12_or0));
  and_gate and_gate_u_csamul_cla32_and16_12(.a(a[16]), .b(b[12]), .out(u_csamul_cla32_and16_12));
  fa fa_u_csamul_cla32_fa16_12_out(.a(u_csamul_cla32_and16_12[0]), .b(u_csamul_cla32_fa17_11_xor1[0]), .cin(u_csamul_cla32_fa16_11_or0[0]), .fa_xor1(u_csamul_cla32_fa16_12_xor1), .fa_or0(u_csamul_cla32_fa16_12_or0));
  and_gate and_gate_u_csamul_cla32_and17_12(.a(a[17]), .b(b[12]), .out(u_csamul_cla32_and17_12));
  fa fa_u_csamul_cla32_fa17_12_out(.a(u_csamul_cla32_and17_12[0]), .b(u_csamul_cla32_fa18_11_xor1[0]), .cin(u_csamul_cla32_fa17_11_or0[0]), .fa_xor1(u_csamul_cla32_fa17_12_xor1), .fa_or0(u_csamul_cla32_fa17_12_or0));
  and_gate and_gate_u_csamul_cla32_and18_12(.a(a[18]), .b(b[12]), .out(u_csamul_cla32_and18_12));
  fa fa_u_csamul_cla32_fa18_12_out(.a(u_csamul_cla32_and18_12[0]), .b(u_csamul_cla32_fa19_11_xor1[0]), .cin(u_csamul_cla32_fa18_11_or0[0]), .fa_xor1(u_csamul_cla32_fa18_12_xor1), .fa_or0(u_csamul_cla32_fa18_12_or0));
  and_gate and_gate_u_csamul_cla32_and19_12(.a(a[19]), .b(b[12]), .out(u_csamul_cla32_and19_12));
  fa fa_u_csamul_cla32_fa19_12_out(.a(u_csamul_cla32_and19_12[0]), .b(u_csamul_cla32_fa20_11_xor1[0]), .cin(u_csamul_cla32_fa19_11_or0[0]), .fa_xor1(u_csamul_cla32_fa19_12_xor1), .fa_or0(u_csamul_cla32_fa19_12_or0));
  and_gate and_gate_u_csamul_cla32_and20_12(.a(a[20]), .b(b[12]), .out(u_csamul_cla32_and20_12));
  fa fa_u_csamul_cla32_fa20_12_out(.a(u_csamul_cla32_and20_12[0]), .b(u_csamul_cla32_fa21_11_xor1[0]), .cin(u_csamul_cla32_fa20_11_or0[0]), .fa_xor1(u_csamul_cla32_fa20_12_xor1), .fa_or0(u_csamul_cla32_fa20_12_or0));
  and_gate and_gate_u_csamul_cla32_and21_12(.a(a[21]), .b(b[12]), .out(u_csamul_cla32_and21_12));
  fa fa_u_csamul_cla32_fa21_12_out(.a(u_csamul_cla32_and21_12[0]), .b(u_csamul_cla32_fa22_11_xor1[0]), .cin(u_csamul_cla32_fa21_11_or0[0]), .fa_xor1(u_csamul_cla32_fa21_12_xor1), .fa_or0(u_csamul_cla32_fa21_12_or0));
  and_gate and_gate_u_csamul_cla32_and22_12(.a(a[22]), .b(b[12]), .out(u_csamul_cla32_and22_12));
  fa fa_u_csamul_cla32_fa22_12_out(.a(u_csamul_cla32_and22_12[0]), .b(u_csamul_cla32_fa23_11_xor1[0]), .cin(u_csamul_cla32_fa22_11_or0[0]), .fa_xor1(u_csamul_cla32_fa22_12_xor1), .fa_or0(u_csamul_cla32_fa22_12_or0));
  and_gate and_gate_u_csamul_cla32_and23_12(.a(a[23]), .b(b[12]), .out(u_csamul_cla32_and23_12));
  fa fa_u_csamul_cla32_fa23_12_out(.a(u_csamul_cla32_and23_12[0]), .b(u_csamul_cla32_fa24_11_xor1[0]), .cin(u_csamul_cla32_fa23_11_or0[0]), .fa_xor1(u_csamul_cla32_fa23_12_xor1), .fa_or0(u_csamul_cla32_fa23_12_or0));
  and_gate and_gate_u_csamul_cla32_and24_12(.a(a[24]), .b(b[12]), .out(u_csamul_cla32_and24_12));
  fa fa_u_csamul_cla32_fa24_12_out(.a(u_csamul_cla32_and24_12[0]), .b(u_csamul_cla32_fa25_11_xor1[0]), .cin(u_csamul_cla32_fa24_11_or0[0]), .fa_xor1(u_csamul_cla32_fa24_12_xor1), .fa_or0(u_csamul_cla32_fa24_12_or0));
  and_gate and_gate_u_csamul_cla32_and25_12(.a(a[25]), .b(b[12]), .out(u_csamul_cla32_and25_12));
  fa fa_u_csamul_cla32_fa25_12_out(.a(u_csamul_cla32_and25_12[0]), .b(u_csamul_cla32_fa26_11_xor1[0]), .cin(u_csamul_cla32_fa25_11_or0[0]), .fa_xor1(u_csamul_cla32_fa25_12_xor1), .fa_or0(u_csamul_cla32_fa25_12_or0));
  and_gate and_gate_u_csamul_cla32_and26_12(.a(a[26]), .b(b[12]), .out(u_csamul_cla32_and26_12));
  fa fa_u_csamul_cla32_fa26_12_out(.a(u_csamul_cla32_and26_12[0]), .b(u_csamul_cla32_fa27_11_xor1[0]), .cin(u_csamul_cla32_fa26_11_or0[0]), .fa_xor1(u_csamul_cla32_fa26_12_xor1), .fa_or0(u_csamul_cla32_fa26_12_or0));
  and_gate and_gate_u_csamul_cla32_and27_12(.a(a[27]), .b(b[12]), .out(u_csamul_cla32_and27_12));
  fa fa_u_csamul_cla32_fa27_12_out(.a(u_csamul_cla32_and27_12[0]), .b(u_csamul_cla32_fa28_11_xor1[0]), .cin(u_csamul_cla32_fa27_11_or0[0]), .fa_xor1(u_csamul_cla32_fa27_12_xor1), .fa_or0(u_csamul_cla32_fa27_12_or0));
  and_gate and_gate_u_csamul_cla32_and28_12(.a(a[28]), .b(b[12]), .out(u_csamul_cla32_and28_12));
  fa fa_u_csamul_cla32_fa28_12_out(.a(u_csamul_cla32_and28_12[0]), .b(u_csamul_cla32_fa29_11_xor1[0]), .cin(u_csamul_cla32_fa28_11_or0[0]), .fa_xor1(u_csamul_cla32_fa28_12_xor1), .fa_or0(u_csamul_cla32_fa28_12_or0));
  and_gate and_gate_u_csamul_cla32_and29_12(.a(a[29]), .b(b[12]), .out(u_csamul_cla32_and29_12));
  fa fa_u_csamul_cla32_fa29_12_out(.a(u_csamul_cla32_and29_12[0]), .b(u_csamul_cla32_fa30_11_xor1[0]), .cin(u_csamul_cla32_fa29_11_or0[0]), .fa_xor1(u_csamul_cla32_fa29_12_xor1), .fa_or0(u_csamul_cla32_fa29_12_or0));
  and_gate and_gate_u_csamul_cla32_and30_12(.a(a[30]), .b(b[12]), .out(u_csamul_cla32_and30_12));
  fa fa_u_csamul_cla32_fa30_12_out(.a(u_csamul_cla32_and30_12[0]), .b(u_csamul_cla32_and31_11[0]), .cin(u_csamul_cla32_fa30_11_or0[0]), .fa_xor1(u_csamul_cla32_fa30_12_xor1), .fa_or0(u_csamul_cla32_fa30_12_or0));
  and_gate and_gate_u_csamul_cla32_and31_12(.a(a[31]), .b(b[12]), .out(u_csamul_cla32_and31_12));
  and_gate and_gate_u_csamul_cla32_and0_13(.a(a[0]), .b(b[13]), .out(u_csamul_cla32_and0_13));
  fa fa_u_csamul_cla32_fa0_13_out(.a(u_csamul_cla32_and0_13[0]), .b(u_csamul_cla32_fa1_12_xor1[0]), .cin(u_csamul_cla32_fa0_12_or0[0]), .fa_xor1(u_csamul_cla32_fa0_13_xor1), .fa_or0(u_csamul_cla32_fa0_13_or0));
  and_gate and_gate_u_csamul_cla32_and1_13(.a(a[1]), .b(b[13]), .out(u_csamul_cla32_and1_13));
  fa fa_u_csamul_cla32_fa1_13_out(.a(u_csamul_cla32_and1_13[0]), .b(u_csamul_cla32_fa2_12_xor1[0]), .cin(u_csamul_cla32_fa1_12_or0[0]), .fa_xor1(u_csamul_cla32_fa1_13_xor1), .fa_or0(u_csamul_cla32_fa1_13_or0));
  and_gate and_gate_u_csamul_cla32_and2_13(.a(a[2]), .b(b[13]), .out(u_csamul_cla32_and2_13));
  fa fa_u_csamul_cla32_fa2_13_out(.a(u_csamul_cla32_and2_13[0]), .b(u_csamul_cla32_fa3_12_xor1[0]), .cin(u_csamul_cla32_fa2_12_or0[0]), .fa_xor1(u_csamul_cla32_fa2_13_xor1), .fa_or0(u_csamul_cla32_fa2_13_or0));
  and_gate and_gate_u_csamul_cla32_and3_13(.a(a[3]), .b(b[13]), .out(u_csamul_cla32_and3_13));
  fa fa_u_csamul_cla32_fa3_13_out(.a(u_csamul_cla32_and3_13[0]), .b(u_csamul_cla32_fa4_12_xor1[0]), .cin(u_csamul_cla32_fa3_12_or0[0]), .fa_xor1(u_csamul_cla32_fa3_13_xor1), .fa_or0(u_csamul_cla32_fa3_13_or0));
  and_gate and_gate_u_csamul_cla32_and4_13(.a(a[4]), .b(b[13]), .out(u_csamul_cla32_and4_13));
  fa fa_u_csamul_cla32_fa4_13_out(.a(u_csamul_cla32_and4_13[0]), .b(u_csamul_cla32_fa5_12_xor1[0]), .cin(u_csamul_cla32_fa4_12_or0[0]), .fa_xor1(u_csamul_cla32_fa4_13_xor1), .fa_or0(u_csamul_cla32_fa4_13_or0));
  and_gate and_gate_u_csamul_cla32_and5_13(.a(a[5]), .b(b[13]), .out(u_csamul_cla32_and5_13));
  fa fa_u_csamul_cla32_fa5_13_out(.a(u_csamul_cla32_and5_13[0]), .b(u_csamul_cla32_fa6_12_xor1[0]), .cin(u_csamul_cla32_fa5_12_or0[0]), .fa_xor1(u_csamul_cla32_fa5_13_xor1), .fa_or0(u_csamul_cla32_fa5_13_or0));
  and_gate and_gate_u_csamul_cla32_and6_13(.a(a[6]), .b(b[13]), .out(u_csamul_cla32_and6_13));
  fa fa_u_csamul_cla32_fa6_13_out(.a(u_csamul_cla32_and6_13[0]), .b(u_csamul_cla32_fa7_12_xor1[0]), .cin(u_csamul_cla32_fa6_12_or0[0]), .fa_xor1(u_csamul_cla32_fa6_13_xor1), .fa_or0(u_csamul_cla32_fa6_13_or0));
  and_gate and_gate_u_csamul_cla32_and7_13(.a(a[7]), .b(b[13]), .out(u_csamul_cla32_and7_13));
  fa fa_u_csamul_cla32_fa7_13_out(.a(u_csamul_cla32_and7_13[0]), .b(u_csamul_cla32_fa8_12_xor1[0]), .cin(u_csamul_cla32_fa7_12_or0[0]), .fa_xor1(u_csamul_cla32_fa7_13_xor1), .fa_or0(u_csamul_cla32_fa7_13_or0));
  and_gate and_gate_u_csamul_cla32_and8_13(.a(a[8]), .b(b[13]), .out(u_csamul_cla32_and8_13));
  fa fa_u_csamul_cla32_fa8_13_out(.a(u_csamul_cla32_and8_13[0]), .b(u_csamul_cla32_fa9_12_xor1[0]), .cin(u_csamul_cla32_fa8_12_or0[0]), .fa_xor1(u_csamul_cla32_fa8_13_xor1), .fa_or0(u_csamul_cla32_fa8_13_or0));
  and_gate and_gate_u_csamul_cla32_and9_13(.a(a[9]), .b(b[13]), .out(u_csamul_cla32_and9_13));
  fa fa_u_csamul_cla32_fa9_13_out(.a(u_csamul_cla32_and9_13[0]), .b(u_csamul_cla32_fa10_12_xor1[0]), .cin(u_csamul_cla32_fa9_12_or0[0]), .fa_xor1(u_csamul_cla32_fa9_13_xor1), .fa_or0(u_csamul_cla32_fa9_13_or0));
  and_gate and_gate_u_csamul_cla32_and10_13(.a(a[10]), .b(b[13]), .out(u_csamul_cla32_and10_13));
  fa fa_u_csamul_cla32_fa10_13_out(.a(u_csamul_cla32_and10_13[0]), .b(u_csamul_cla32_fa11_12_xor1[0]), .cin(u_csamul_cla32_fa10_12_or0[0]), .fa_xor1(u_csamul_cla32_fa10_13_xor1), .fa_or0(u_csamul_cla32_fa10_13_or0));
  and_gate and_gate_u_csamul_cla32_and11_13(.a(a[11]), .b(b[13]), .out(u_csamul_cla32_and11_13));
  fa fa_u_csamul_cla32_fa11_13_out(.a(u_csamul_cla32_and11_13[0]), .b(u_csamul_cla32_fa12_12_xor1[0]), .cin(u_csamul_cla32_fa11_12_or0[0]), .fa_xor1(u_csamul_cla32_fa11_13_xor1), .fa_or0(u_csamul_cla32_fa11_13_or0));
  and_gate and_gate_u_csamul_cla32_and12_13(.a(a[12]), .b(b[13]), .out(u_csamul_cla32_and12_13));
  fa fa_u_csamul_cla32_fa12_13_out(.a(u_csamul_cla32_and12_13[0]), .b(u_csamul_cla32_fa13_12_xor1[0]), .cin(u_csamul_cla32_fa12_12_or0[0]), .fa_xor1(u_csamul_cla32_fa12_13_xor1), .fa_or0(u_csamul_cla32_fa12_13_or0));
  and_gate and_gate_u_csamul_cla32_and13_13(.a(a[13]), .b(b[13]), .out(u_csamul_cla32_and13_13));
  fa fa_u_csamul_cla32_fa13_13_out(.a(u_csamul_cla32_and13_13[0]), .b(u_csamul_cla32_fa14_12_xor1[0]), .cin(u_csamul_cla32_fa13_12_or0[0]), .fa_xor1(u_csamul_cla32_fa13_13_xor1), .fa_or0(u_csamul_cla32_fa13_13_or0));
  and_gate and_gate_u_csamul_cla32_and14_13(.a(a[14]), .b(b[13]), .out(u_csamul_cla32_and14_13));
  fa fa_u_csamul_cla32_fa14_13_out(.a(u_csamul_cla32_and14_13[0]), .b(u_csamul_cla32_fa15_12_xor1[0]), .cin(u_csamul_cla32_fa14_12_or0[0]), .fa_xor1(u_csamul_cla32_fa14_13_xor1), .fa_or0(u_csamul_cla32_fa14_13_or0));
  and_gate and_gate_u_csamul_cla32_and15_13(.a(a[15]), .b(b[13]), .out(u_csamul_cla32_and15_13));
  fa fa_u_csamul_cla32_fa15_13_out(.a(u_csamul_cla32_and15_13[0]), .b(u_csamul_cla32_fa16_12_xor1[0]), .cin(u_csamul_cla32_fa15_12_or0[0]), .fa_xor1(u_csamul_cla32_fa15_13_xor1), .fa_or0(u_csamul_cla32_fa15_13_or0));
  and_gate and_gate_u_csamul_cla32_and16_13(.a(a[16]), .b(b[13]), .out(u_csamul_cla32_and16_13));
  fa fa_u_csamul_cla32_fa16_13_out(.a(u_csamul_cla32_and16_13[0]), .b(u_csamul_cla32_fa17_12_xor1[0]), .cin(u_csamul_cla32_fa16_12_or0[0]), .fa_xor1(u_csamul_cla32_fa16_13_xor1), .fa_or0(u_csamul_cla32_fa16_13_or0));
  and_gate and_gate_u_csamul_cla32_and17_13(.a(a[17]), .b(b[13]), .out(u_csamul_cla32_and17_13));
  fa fa_u_csamul_cla32_fa17_13_out(.a(u_csamul_cla32_and17_13[0]), .b(u_csamul_cla32_fa18_12_xor1[0]), .cin(u_csamul_cla32_fa17_12_or0[0]), .fa_xor1(u_csamul_cla32_fa17_13_xor1), .fa_or0(u_csamul_cla32_fa17_13_or0));
  and_gate and_gate_u_csamul_cla32_and18_13(.a(a[18]), .b(b[13]), .out(u_csamul_cla32_and18_13));
  fa fa_u_csamul_cla32_fa18_13_out(.a(u_csamul_cla32_and18_13[0]), .b(u_csamul_cla32_fa19_12_xor1[0]), .cin(u_csamul_cla32_fa18_12_or0[0]), .fa_xor1(u_csamul_cla32_fa18_13_xor1), .fa_or0(u_csamul_cla32_fa18_13_or0));
  and_gate and_gate_u_csamul_cla32_and19_13(.a(a[19]), .b(b[13]), .out(u_csamul_cla32_and19_13));
  fa fa_u_csamul_cla32_fa19_13_out(.a(u_csamul_cla32_and19_13[0]), .b(u_csamul_cla32_fa20_12_xor1[0]), .cin(u_csamul_cla32_fa19_12_or0[0]), .fa_xor1(u_csamul_cla32_fa19_13_xor1), .fa_or0(u_csamul_cla32_fa19_13_or0));
  and_gate and_gate_u_csamul_cla32_and20_13(.a(a[20]), .b(b[13]), .out(u_csamul_cla32_and20_13));
  fa fa_u_csamul_cla32_fa20_13_out(.a(u_csamul_cla32_and20_13[0]), .b(u_csamul_cla32_fa21_12_xor1[0]), .cin(u_csamul_cla32_fa20_12_or0[0]), .fa_xor1(u_csamul_cla32_fa20_13_xor1), .fa_or0(u_csamul_cla32_fa20_13_or0));
  and_gate and_gate_u_csamul_cla32_and21_13(.a(a[21]), .b(b[13]), .out(u_csamul_cla32_and21_13));
  fa fa_u_csamul_cla32_fa21_13_out(.a(u_csamul_cla32_and21_13[0]), .b(u_csamul_cla32_fa22_12_xor1[0]), .cin(u_csamul_cla32_fa21_12_or0[0]), .fa_xor1(u_csamul_cla32_fa21_13_xor1), .fa_or0(u_csamul_cla32_fa21_13_or0));
  and_gate and_gate_u_csamul_cla32_and22_13(.a(a[22]), .b(b[13]), .out(u_csamul_cla32_and22_13));
  fa fa_u_csamul_cla32_fa22_13_out(.a(u_csamul_cla32_and22_13[0]), .b(u_csamul_cla32_fa23_12_xor1[0]), .cin(u_csamul_cla32_fa22_12_or0[0]), .fa_xor1(u_csamul_cla32_fa22_13_xor1), .fa_or0(u_csamul_cla32_fa22_13_or0));
  and_gate and_gate_u_csamul_cla32_and23_13(.a(a[23]), .b(b[13]), .out(u_csamul_cla32_and23_13));
  fa fa_u_csamul_cla32_fa23_13_out(.a(u_csamul_cla32_and23_13[0]), .b(u_csamul_cla32_fa24_12_xor1[0]), .cin(u_csamul_cla32_fa23_12_or0[0]), .fa_xor1(u_csamul_cla32_fa23_13_xor1), .fa_or0(u_csamul_cla32_fa23_13_or0));
  and_gate and_gate_u_csamul_cla32_and24_13(.a(a[24]), .b(b[13]), .out(u_csamul_cla32_and24_13));
  fa fa_u_csamul_cla32_fa24_13_out(.a(u_csamul_cla32_and24_13[0]), .b(u_csamul_cla32_fa25_12_xor1[0]), .cin(u_csamul_cla32_fa24_12_or0[0]), .fa_xor1(u_csamul_cla32_fa24_13_xor1), .fa_or0(u_csamul_cla32_fa24_13_or0));
  and_gate and_gate_u_csamul_cla32_and25_13(.a(a[25]), .b(b[13]), .out(u_csamul_cla32_and25_13));
  fa fa_u_csamul_cla32_fa25_13_out(.a(u_csamul_cla32_and25_13[0]), .b(u_csamul_cla32_fa26_12_xor1[0]), .cin(u_csamul_cla32_fa25_12_or0[0]), .fa_xor1(u_csamul_cla32_fa25_13_xor1), .fa_or0(u_csamul_cla32_fa25_13_or0));
  and_gate and_gate_u_csamul_cla32_and26_13(.a(a[26]), .b(b[13]), .out(u_csamul_cla32_and26_13));
  fa fa_u_csamul_cla32_fa26_13_out(.a(u_csamul_cla32_and26_13[0]), .b(u_csamul_cla32_fa27_12_xor1[0]), .cin(u_csamul_cla32_fa26_12_or0[0]), .fa_xor1(u_csamul_cla32_fa26_13_xor1), .fa_or0(u_csamul_cla32_fa26_13_or0));
  and_gate and_gate_u_csamul_cla32_and27_13(.a(a[27]), .b(b[13]), .out(u_csamul_cla32_and27_13));
  fa fa_u_csamul_cla32_fa27_13_out(.a(u_csamul_cla32_and27_13[0]), .b(u_csamul_cla32_fa28_12_xor1[0]), .cin(u_csamul_cla32_fa27_12_or0[0]), .fa_xor1(u_csamul_cla32_fa27_13_xor1), .fa_or0(u_csamul_cla32_fa27_13_or0));
  and_gate and_gate_u_csamul_cla32_and28_13(.a(a[28]), .b(b[13]), .out(u_csamul_cla32_and28_13));
  fa fa_u_csamul_cla32_fa28_13_out(.a(u_csamul_cla32_and28_13[0]), .b(u_csamul_cla32_fa29_12_xor1[0]), .cin(u_csamul_cla32_fa28_12_or0[0]), .fa_xor1(u_csamul_cla32_fa28_13_xor1), .fa_or0(u_csamul_cla32_fa28_13_or0));
  and_gate and_gate_u_csamul_cla32_and29_13(.a(a[29]), .b(b[13]), .out(u_csamul_cla32_and29_13));
  fa fa_u_csamul_cla32_fa29_13_out(.a(u_csamul_cla32_and29_13[0]), .b(u_csamul_cla32_fa30_12_xor1[0]), .cin(u_csamul_cla32_fa29_12_or0[0]), .fa_xor1(u_csamul_cla32_fa29_13_xor1), .fa_or0(u_csamul_cla32_fa29_13_or0));
  and_gate and_gate_u_csamul_cla32_and30_13(.a(a[30]), .b(b[13]), .out(u_csamul_cla32_and30_13));
  fa fa_u_csamul_cla32_fa30_13_out(.a(u_csamul_cla32_and30_13[0]), .b(u_csamul_cla32_and31_12[0]), .cin(u_csamul_cla32_fa30_12_or0[0]), .fa_xor1(u_csamul_cla32_fa30_13_xor1), .fa_or0(u_csamul_cla32_fa30_13_or0));
  and_gate and_gate_u_csamul_cla32_and31_13(.a(a[31]), .b(b[13]), .out(u_csamul_cla32_and31_13));
  and_gate and_gate_u_csamul_cla32_and0_14(.a(a[0]), .b(b[14]), .out(u_csamul_cla32_and0_14));
  fa fa_u_csamul_cla32_fa0_14_out(.a(u_csamul_cla32_and0_14[0]), .b(u_csamul_cla32_fa1_13_xor1[0]), .cin(u_csamul_cla32_fa0_13_or0[0]), .fa_xor1(u_csamul_cla32_fa0_14_xor1), .fa_or0(u_csamul_cla32_fa0_14_or0));
  and_gate and_gate_u_csamul_cla32_and1_14(.a(a[1]), .b(b[14]), .out(u_csamul_cla32_and1_14));
  fa fa_u_csamul_cla32_fa1_14_out(.a(u_csamul_cla32_and1_14[0]), .b(u_csamul_cla32_fa2_13_xor1[0]), .cin(u_csamul_cla32_fa1_13_or0[0]), .fa_xor1(u_csamul_cla32_fa1_14_xor1), .fa_or0(u_csamul_cla32_fa1_14_or0));
  and_gate and_gate_u_csamul_cla32_and2_14(.a(a[2]), .b(b[14]), .out(u_csamul_cla32_and2_14));
  fa fa_u_csamul_cla32_fa2_14_out(.a(u_csamul_cla32_and2_14[0]), .b(u_csamul_cla32_fa3_13_xor1[0]), .cin(u_csamul_cla32_fa2_13_or0[0]), .fa_xor1(u_csamul_cla32_fa2_14_xor1), .fa_or0(u_csamul_cla32_fa2_14_or0));
  and_gate and_gate_u_csamul_cla32_and3_14(.a(a[3]), .b(b[14]), .out(u_csamul_cla32_and3_14));
  fa fa_u_csamul_cla32_fa3_14_out(.a(u_csamul_cla32_and3_14[0]), .b(u_csamul_cla32_fa4_13_xor1[0]), .cin(u_csamul_cla32_fa3_13_or0[0]), .fa_xor1(u_csamul_cla32_fa3_14_xor1), .fa_or0(u_csamul_cla32_fa3_14_or0));
  and_gate and_gate_u_csamul_cla32_and4_14(.a(a[4]), .b(b[14]), .out(u_csamul_cla32_and4_14));
  fa fa_u_csamul_cla32_fa4_14_out(.a(u_csamul_cla32_and4_14[0]), .b(u_csamul_cla32_fa5_13_xor1[0]), .cin(u_csamul_cla32_fa4_13_or0[0]), .fa_xor1(u_csamul_cla32_fa4_14_xor1), .fa_or0(u_csamul_cla32_fa4_14_or0));
  and_gate and_gate_u_csamul_cla32_and5_14(.a(a[5]), .b(b[14]), .out(u_csamul_cla32_and5_14));
  fa fa_u_csamul_cla32_fa5_14_out(.a(u_csamul_cla32_and5_14[0]), .b(u_csamul_cla32_fa6_13_xor1[0]), .cin(u_csamul_cla32_fa5_13_or0[0]), .fa_xor1(u_csamul_cla32_fa5_14_xor1), .fa_or0(u_csamul_cla32_fa5_14_or0));
  and_gate and_gate_u_csamul_cla32_and6_14(.a(a[6]), .b(b[14]), .out(u_csamul_cla32_and6_14));
  fa fa_u_csamul_cla32_fa6_14_out(.a(u_csamul_cla32_and6_14[0]), .b(u_csamul_cla32_fa7_13_xor1[0]), .cin(u_csamul_cla32_fa6_13_or0[0]), .fa_xor1(u_csamul_cla32_fa6_14_xor1), .fa_or0(u_csamul_cla32_fa6_14_or0));
  and_gate and_gate_u_csamul_cla32_and7_14(.a(a[7]), .b(b[14]), .out(u_csamul_cla32_and7_14));
  fa fa_u_csamul_cla32_fa7_14_out(.a(u_csamul_cla32_and7_14[0]), .b(u_csamul_cla32_fa8_13_xor1[0]), .cin(u_csamul_cla32_fa7_13_or0[0]), .fa_xor1(u_csamul_cla32_fa7_14_xor1), .fa_or0(u_csamul_cla32_fa7_14_or0));
  and_gate and_gate_u_csamul_cla32_and8_14(.a(a[8]), .b(b[14]), .out(u_csamul_cla32_and8_14));
  fa fa_u_csamul_cla32_fa8_14_out(.a(u_csamul_cla32_and8_14[0]), .b(u_csamul_cla32_fa9_13_xor1[0]), .cin(u_csamul_cla32_fa8_13_or0[0]), .fa_xor1(u_csamul_cla32_fa8_14_xor1), .fa_or0(u_csamul_cla32_fa8_14_or0));
  and_gate and_gate_u_csamul_cla32_and9_14(.a(a[9]), .b(b[14]), .out(u_csamul_cla32_and9_14));
  fa fa_u_csamul_cla32_fa9_14_out(.a(u_csamul_cla32_and9_14[0]), .b(u_csamul_cla32_fa10_13_xor1[0]), .cin(u_csamul_cla32_fa9_13_or0[0]), .fa_xor1(u_csamul_cla32_fa9_14_xor1), .fa_or0(u_csamul_cla32_fa9_14_or0));
  and_gate and_gate_u_csamul_cla32_and10_14(.a(a[10]), .b(b[14]), .out(u_csamul_cla32_and10_14));
  fa fa_u_csamul_cla32_fa10_14_out(.a(u_csamul_cla32_and10_14[0]), .b(u_csamul_cla32_fa11_13_xor1[0]), .cin(u_csamul_cla32_fa10_13_or0[0]), .fa_xor1(u_csamul_cla32_fa10_14_xor1), .fa_or0(u_csamul_cla32_fa10_14_or0));
  and_gate and_gate_u_csamul_cla32_and11_14(.a(a[11]), .b(b[14]), .out(u_csamul_cla32_and11_14));
  fa fa_u_csamul_cla32_fa11_14_out(.a(u_csamul_cla32_and11_14[0]), .b(u_csamul_cla32_fa12_13_xor1[0]), .cin(u_csamul_cla32_fa11_13_or0[0]), .fa_xor1(u_csamul_cla32_fa11_14_xor1), .fa_or0(u_csamul_cla32_fa11_14_or0));
  and_gate and_gate_u_csamul_cla32_and12_14(.a(a[12]), .b(b[14]), .out(u_csamul_cla32_and12_14));
  fa fa_u_csamul_cla32_fa12_14_out(.a(u_csamul_cla32_and12_14[0]), .b(u_csamul_cla32_fa13_13_xor1[0]), .cin(u_csamul_cla32_fa12_13_or0[0]), .fa_xor1(u_csamul_cla32_fa12_14_xor1), .fa_or0(u_csamul_cla32_fa12_14_or0));
  and_gate and_gate_u_csamul_cla32_and13_14(.a(a[13]), .b(b[14]), .out(u_csamul_cla32_and13_14));
  fa fa_u_csamul_cla32_fa13_14_out(.a(u_csamul_cla32_and13_14[0]), .b(u_csamul_cla32_fa14_13_xor1[0]), .cin(u_csamul_cla32_fa13_13_or0[0]), .fa_xor1(u_csamul_cla32_fa13_14_xor1), .fa_or0(u_csamul_cla32_fa13_14_or0));
  and_gate and_gate_u_csamul_cla32_and14_14(.a(a[14]), .b(b[14]), .out(u_csamul_cla32_and14_14));
  fa fa_u_csamul_cla32_fa14_14_out(.a(u_csamul_cla32_and14_14[0]), .b(u_csamul_cla32_fa15_13_xor1[0]), .cin(u_csamul_cla32_fa14_13_or0[0]), .fa_xor1(u_csamul_cla32_fa14_14_xor1), .fa_or0(u_csamul_cla32_fa14_14_or0));
  and_gate and_gate_u_csamul_cla32_and15_14(.a(a[15]), .b(b[14]), .out(u_csamul_cla32_and15_14));
  fa fa_u_csamul_cla32_fa15_14_out(.a(u_csamul_cla32_and15_14[0]), .b(u_csamul_cla32_fa16_13_xor1[0]), .cin(u_csamul_cla32_fa15_13_or0[0]), .fa_xor1(u_csamul_cla32_fa15_14_xor1), .fa_or0(u_csamul_cla32_fa15_14_or0));
  and_gate and_gate_u_csamul_cla32_and16_14(.a(a[16]), .b(b[14]), .out(u_csamul_cla32_and16_14));
  fa fa_u_csamul_cla32_fa16_14_out(.a(u_csamul_cla32_and16_14[0]), .b(u_csamul_cla32_fa17_13_xor1[0]), .cin(u_csamul_cla32_fa16_13_or0[0]), .fa_xor1(u_csamul_cla32_fa16_14_xor1), .fa_or0(u_csamul_cla32_fa16_14_or0));
  and_gate and_gate_u_csamul_cla32_and17_14(.a(a[17]), .b(b[14]), .out(u_csamul_cla32_and17_14));
  fa fa_u_csamul_cla32_fa17_14_out(.a(u_csamul_cla32_and17_14[0]), .b(u_csamul_cla32_fa18_13_xor1[0]), .cin(u_csamul_cla32_fa17_13_or0[0]), .fa_xor1(u_csamul_cla32_fa17_14_xor1), .fa_or0(u_csamul_cla32_fa17_14_or0));
  and_gate and_gate_u_csamul_cla32_and18_14(.a(a[18]), .b(b[14]), .out(u_csamul_cla32_and18_14));
  fa fa_u_csamul_cla32_fa18_14_out(.a(u_csamul_cla32_and18_14[0]), .b(u_csamul_cla32_fa19_13_xor1[0]), .cin(u_csamul_cla32_fa18_13_or0[0]), .fa_xor1(u_csamul_cla32_fa18_14_xor1), .fa_or0(u_csamul_cla32_fa18_14_or0));
  and_gate and_gate_u_csamul_cla32_and19_14(.a(a[19]), .b(b[14]), .out(u_csamul_cla32_and19_14));
  fa fa_u_csamul_cla32_fa19_14_out(.a(u_csamul_cla32_and19_14[0]), .b(u_csamul_cla32_fa20_13_xor1[0]), .cin(u_csamul_cla32_fa19_13_or0[0]), .fa_xor1(u_csamul_cla32_fa19_14_xor1), .fa_or0(u_csamul_cla32_fa19_14_or0));
  and_gate and_gate_u_csamul_cla32_and20_14(.a(a[20]), .b(b[14]), .out(u_csamul_cla32_and20_14));
  fa fa_u_csamul_cla32_fa20_14_out(.a(u_csamul_cla32_and20_14[0]), .b(u_csamul_cla32_fa21_13_xor1[0]), .cin(u_csamul_cla32_fa20_13_or0[0]), .fa_xor1(u_csamul_cla32_fa20_14_xor1), .fa_or0(u_csamul_cla32_fa20_14_or0));
  and_gate and_gate_u_csamul_cla32_and21_14(.a(a[21]), .b(b[14]), .out(u_csamul_cla32_and21_14));
  fa fa_u_csamul_cla32_fa21_14_out(.a(u_csamul_cla32_and21_14[0]), .b(u_csamul_cla32_fa22_13_xor1[0]), .cin(u_csamul_cla32_fa21_13_or0[0]), .fa_xor1(u_csamul_cla32_fa21_14_xor1), .fa_or0(u_csamul_cla32_fa21_14_or0));
  and_gate and_gate_u_csamul_cla32_and22_14(.a(a[22]), .b(b[14]), .out(u_csamul_cla32_and22_14));
  fa fa_u_csamul_cla32_fa22_14_out(.a(u_csamul_cla32_and22_14[0]), .b(u_csamul_cla32_fa23_13_xor1[0]), .cin(u_csamul_cla32_fa22_13_or0[0]), .fa_xor1(u_csamul_cla32_fa22_14_xor1), .fa_or0(u_csamul_cla32_fa22_14_or0));
  and_gate and_gate_u_csamul_cla32_and23_14(.a(a[23]), .b(b[14]), .out(u_csamul_cla32_and23_14));
  fa fa_u_csamul_cla32_fa23_14_out(.a(u_csamul_cla32_and23_14[0]), .b(u_csamul_cla32_fa24_13_xor1[0]), .cin(u_csamul_cla32_fa23_13_or0[0]), .fa_xor1(u_csamul_cla32_fa23_14_xor1), .fa_or0(u_csamul_cla32_fa23_14_or0));
  and_gate and_gate_u_csamul_cla32_and24_14(.a(a[24]), .b(b[14]), .out(u_csamul_cla32_and24_14));
  fa fa_u_csamul_cla32_fa24_14_out(.a(u_csamul_cla32_and24_14[0]), .b(u_csamul_cla32_fa25_13_xor1[0]), .cin(u_csamul_cla32_fa24_13_or0[0]), .fa_xor1(u_csamul_cla32_fa24_14_xor1), .fa_or0(u_csamul_cla32_fa24_14_or0));
  and_gate and_gate_u_csamul_cla32_and25_14(.a(a[25]), .b(b[14]), .out(u_csamul_cla32_and25_14));
  fa fa_u_csamul_cla32_fa25_14_out(.a(u_csamul_cla32_and25_14[0]), .b(u_csamul_cla32_fa26_13_xor1[0]), .cin(u_csamul_cla32_fa25_13_or0[0]), .fa_xor1(u_csamul_cla32_fa25_14_xor1), .fa_or0(u_csamul_cla32_fa25_14_or0));
  and_gate and_gate_u_csamul_cla32_and26_14(.a(a[26]), .b(b[14]), .out(u_csamul_cla32_and26_14));
  fa fa_u_csamul_cla32_fa26_14_out(.a(u_csamul_cla32_and26_14[0]), .b(u_csamul_cla32_fa27_13_xor1[0]), .cin(u_csamul_cla32_fa26_13_or0[0]), .fa_xor1(u_csamul_cla32_fa26_14_xor1), .fa_or0(u_csamul_cla32_fa26_14_or0));
  and_gate and_gate_u_csamul_cla32_and27_14(.a(a[27]), .b(b[14]), .out(u_csamul_cla32_and27_14));
  fa fa_u_csamul_cla32_fa27_14_out(.a(u_csamul_cla32_and27_14[0]), .b(u_csamul_cla32_fa28_13_xor1[0]), .cin(u_csamul_cla32_fa27_13_or0[0]), .fa_xor1(u_csamul_cla32_fa27_14_xor1), .fa_or0(u_csamul_cla32_fa27_14_or0));
  and_gate and_gate_u_csamul_cla32_and28_14(.a(a[28]), .b(b[14]), .out(u_csamul_cla32_and28_14));
  fa fa_u_csamul_cla32_fa28_14_out(.a(u_csamul_cla32_and28_14[0]), .b(u_csamul_cla32_fa29_13_xor1[0]), .cin(u_csamul_cla32_fa28_13_or0[0]), .fa_xor1(u_csamul_cla32_fa28_14_xor1), .fa_or0(u_csamul_cla32_fa28_14_or0));
  and_gate and_gate_u_csamul_cla32_and29_14(.a(a[29]), .b(b[14]), .out(u_csamul_cla32_and29_14));
  fa fa_u_csamul_cla32_fa29_14_out(.a(u_csamul_cla32_and29_14[0]), .b(u_csamul_cla32_fa30_13_xor1[0]), .cin(u_csamul_cla32_fa29_13_or0[0]), .fa_xor1(u_csamul_cla32_fa29_14_xor1), .fa_or0(u_csamul_cla32_fa29_14_or0));
  and_gate and_gate_u_csamul_cla32_and30_14(.a(a[30]), .b(b[14]), .out(u_csamul_cla32_and30_14));
  fa fa_u_csamul_cla32_fa30_14_out(.a(u_csamul_cla32_and30_14[0]), .b(u_csamul_cla32_and31_13[0]), .cin(u_csamul_cla32_fa30_13_or0[0]), .fa_xor1(u_csamul_cla32_fa30_14_xor1), .fa_or0(u_csamul_cla32_fa30_14_or0));
  and_gate and_gate_u_csamul_cla32_and31_14(.a(a[31]), .b(b[14]), .out(u_csamul_cla32_and31_14));
  and_gate and_gate_u_csamul_cla32_and0_15(.a(a[0]), .b(b[15]), .out(u_csamul_cla32_and0_15));
  fa fa_u_csamul_cla32_fa0_15_out(.a(u_csamul_cla32_and0_15[0]), .b(u_csamul_cla32_fa1_14_xor1[0]), .cin(u_csamul_cla32_fa0_14_or0[0]), .fa_xor1(u_csamul_cla32_fa0_15_xor1), .fa_or0(u_csamul_cla32_fa0_15_or0));
  and_gate and_gate_u_csamul_cla32_and1_15(.a(a[1]), .b(b[15]), .out(u_csamul_cla32_and1_15));
  fa fa_u_csamul_cla32_fa1_15_out(.a(u_csamul_cla32_and1_15[0]), .b(u_csamul_cla32_fa2_14_xor1[0]), .cin(u_csamul_cla32_fa1_14_or0[0]), .fa_xor1(u_csamul_cla32_fa1_15_xor1), .fa_or0(u_csamul_cla32_fa1_15_or0));
  and_gate and_gate_u_csamul_cla32_and2_15(.a(a[2]), .b(b[15]), .out(u_csamul_cla32_and2_15));
  fa fa_u_csamul_cla32_fa2_15_out(.a(u_csamul_cla32_and2_15[0]), .b(u_csamul_cla32_fa3_14_xor1[0]), .cin(u_csamul_cla32_fa2_14_or0[0]), .fa_xor1(u_csamul_cla32_fa2_15_xor1), .fa_or0(u_csamul_cla32_fa2_15_or0));
  and_gate and_gate_u_csamul_cla32_and3_15(.a(a[3]), .b(b[15]), .out(u_csamul_cla32_and3_15));
  fa fa_u_csamul_cla32_fa3_15_out(.a(u_csamul_cla32_and3_15[0]), .b(u_csamul_cla32_fa4_14_xor1[0]), .cin(u_csamul_cla32_fa3_14_or0[0]), .fa_xor1(u_csamul_cla32_fa3_15_xor1), .fa_or0(u_csamul_cla32_fa3_15_or0));
  and_gate and_gate_u_csamul_cla32_and4_15(.a(a[4]), .b(b[15]), .out(u_csamul_cla32_and4_15));
  fa fa_u_csamul_cla32_fa4_15_out(.a(u_csamul_cla32_and4_15[0]), .b(u_csamul_cla32_fa5_14_xor1[0]), .cin(u_csamul_cla32_fa4_14_or0[0]), .fa_xor1(u_csamul_cla32_fa4_15_xor1), .fa_or0(u_csamul_cla32_fa4_15_or0));
  and_gate and_gate_u_csamul_cla32_and5_15(.a(a[5]), .b(b[15]), .out(u_csamul_cla32_and5_15));
  fa fa_u_csamul_cla32_fa5_15_out(.a(u_csamul_cla32_and5_15[0]), .b(u_csamul_cla32_fa6_14_xor1[0]), .cin(u_csamul_cla32_fa5_14_or0[0]), .fa_xor1(u_csamul_cla32_fa5_15_xor1), .fa_or0(u_csamul_cla32_fa5_15_or0));
  and_gate and_gate_u_csamul_cla32_and6_15(.a(a[6]), .b(b[15]), .out(u_csamul_cla32_and6_15));
  fa fa_u_csamul_cla32_fa6_15_out(.a(u_csamul_cla32_and6_15[0]), .b(u_csamul_cla32_fa7_14_xor1[0]), .cin(u_csamul_cla32_fa6_14_or0[0]), .fa_xor1(u_csamul_cla32_fa6_15_xor1), .fa_or0(u_csamul_cla32_fa6_15_or0));
  and_gate and_gate_u_csamul_cla32_and7_15(.a(a[7]), .b(b[15]), .out(u_csamul_cla32_and7_15));
  fa fa_u_csamul_cla32_fa7_15_out(.a(u_csamul_cla32_and7_15[0]), .b(u_csamul_cla32_fa8_14_xor1[0]), .cin(u_csamul_cla32_fa7_14_or0[0]), .fa_xor1(u_csamul_cla32_fa7_15_xor1), .fa_or0(u_csamul_cla32_fa7_15_or0));
  and_gate and_gate_u_csamul_cla32_and8_15(.a(a[8]), .b(b[15]), .out(u_csamul_cla32_and8_15));
  fa fa_u_csamul_cla32_fa8_15_out(.a(u_csamul_cla32_and8_15[0]), .b(u_csamul_cla32_fa9_14_xor1[0]), .cin(u_csamul_cla32_fa8_14_or0[0]), .fa_xor1(u_csamul_cla32_fa8_15_xor1), .fa_or0(u_csamul_cla32_fa8_15_or0));
  and_gate and_gate_u_csamul_cla32_and9_15(.a(a[9]), .b(b[15]), .out(u_csamul_cla32_and9_15));
  fa fa_u_csamul_cla32_fa9_15_out(.a(u_csamul_cla32_and9_15[0]), .b(u_csamul_cla32_fa10_14_xor1[0]), .cin(u_csamul_cla32_fa9_14_or0[0]), .fa_xor1(u_csamul_cla32_fa9_15_xor1), .fa_or0(u_csamul_cla32_fa9_15_or0));
  and_gate and_gate_u_csamul_cla32_and10_15(.a(a[10]), .b(b[15]), .out(u_csamul_cla32_and10_15));
  fa fa_u_csamul_cla32_fa10_15_out(.a(u_csamul_cla32_and10_15[0]), .b(u_csamul_cla32_fa11_14_xor1[0]), .cin(u_csamul_cla32_fa10_14_or0[0]), .fa_xor1(u_csamul_cla32_fa10_15_xor1), .fa_or0(u_csamul_cla32_fa10_15_or0));
  and_gate and_gate_u_csamul_cla32_and11_15(.a(a[11]), .b(b[15]), .out(u_csamul_cla32_and11_15));
  fa fa_u_csamul_cla32_fa11_15_out(.a(u_csamul_cla32_and11_15[0]), .b(u_csamul_cla32_fa12_14_xor1[0]), .cin(u_csamul_cla32_fa11_14_or0[0]), .fa_xor1(u_csamul_cla32_fa11_15_xor1), .fa_or0(u_csamul_cla32_fa11_15_or0));
  and_gate and_gate_u_csamul_cla32_and12_15(.a(a[12]), .b(b[15]), .out(u_csamul_cla32_and12_15));
  fa fa_u_csamul_cla32_fa12_15_out(.a(u_csamul_cla32_and12_15[0]), .b(u_csamul_cla32_fa13_14_xor1[0]), .cin(u_csamul_cla32_fa12_14_or0[0]), .fa_xor1(u_csamul_cla32_fa12_15_xor1), .fa_or0(u_csamul_cla32_fa12_15_or0));
  and_gate and_gate_u_csamul_cla32_and13_15(.a(a[13]), .b(b[15]), .out(u_csamul_cla32_and13_15));
  fa fa_u_csamul_cla32_fa13_15_out(.a(u_csamul_cla32_and13_15[0]), .b(u_csamul_cla32_fa14_14_xor1[0]), .cin(u_csamul_cla32_fa13_14_or0[0]), .fa_xor1(u_csamul_cla32_fa13_15_xor1), .fa_or0(u_csamul_cla32_fa13_15_or0));
  and_gate and_gate_u_csamul_cla32_and14_15(.a(a[14]), .b(b[15]), .out(u_csamul_cla32_and14_15));
  fa fa_u_csamul_cla32_fa14_15_out(.a(u_csamul_cla32_and14_15[0]), .b(u_csamul_cla32_fa15_14_xor1[0]), .cin(u_csamul_cla32_fa14_14_or0[0]), .fa_xor1(u_csamul_cla32_fa14_15_xor1), .fa_or0(u_csamul_cla32_fa14_15_or0));
  and_gate and_gate_u_csamul_cla32_and15_15(.a(a[15]), .b(b[15]), .out(u_csamul_cla32_and15_15));
  fa fa_u_csamul_cla32_fa15_15_out(.a(u_csamul_cla32_and15_15[0]), .b(u_csamul_cla32_fa16_14_xor1[0]), .cin(u_csamul_cla32_fa15_14_or0[0]), .fa_xor1(u_csamul_cla32_fa15_15_xor1), .fa_or0(u_csamul_cla32_fa15_15_or0));
  and_gate and_gate_u_csamul_cla32_and16_15(.a(a[16]), .b(b[15]), .out(u_csamul_cla32_and16_15));
  fa fa_u_csamul_cla32_fa16_15_out(.a(u_csamul_cla32_and16_15[0]), .b(u_csamul_cla32_fa17_14_xor1[0]), .cin(u_csamul_cla32_fa16_14_or0[0]), .fa_xor1(u_csamul_cla32_fa16_15_xor1), .fa_or0(u_csamul_cla32_fa16_15_or0));
  and_gate and_gate_u_csamul_cla32_and17_15(.a(a[17]), .b(b[15]), .out(u_csamul_cla32_and17_15));
  fa fa_u_csamul_cla32_fa17_15_out(.a(u_csamul_cla32_and17_15[0]), .b(u_csamul_cla32_fa18_14_xor1[0]), .cin(u_csamul_cla32_fa17_14_or0[0]), .fa_xor1(u_csamul_cla32_fa17_15_xor1), .fa_or0(u_csamul_cla32_fa17_15_or0));
  and_gate and_gate_u_csamul_cla32_and18_15(.a(a[18]), .b(b[15]), .out(u_csamul_cla32_and18_15));
  fa fa_u_csamul_cla32_fa18_15_out(.a(u_csamul_cla32_and18_15[0]), .b(u_csamul_cla32_fa19_14_xor1[0]), .cin(u_csamul_cla32_fa18_14_or0[0]), .fa_xor1(u_csamul_cla32_fa18_15_xor1), .fa_or0(u_csamul_cla32_fa18_15_or0));
  and_gate and_gate_u_csamul_cla32_and19_15(.a(a[19]), .b(b[15]), .out(u_csamul_cla32_and19_15));
  fa fa_u_csamul_cla32_fa19_15_out(.a(u_csamul_cla32_and19_15[0]), .b(u_csamul_cla32_fa20_14_xor1[0]), .cin(u_csamul_cla32_fa19_14_or0[0]), .fa_xor1(u_csamul_cla32_fa19_15_xor1), .fa_or0(u_csamul_cla32_fa19_15_or0));
  and_gate and_gate_u_csamul_cla32_and20_15(.a(a[20]), .b(b[15]), .out(u_csamul_cla32_and20_15));
  fa fa_u_csamul_cla32_fa20_15_out(.a(u_csamul_cla32_and20_15[0]), .b(u_csamul_cla32_fa21_14_xor1[0]), .cin(u_csamul_cla32_fa20_14_or0[0]), .fa_xor1(u_csamul_cla32_fa20_15_xor1), .fa_or0(u_csamul_cla32_fa20_15_or0));
  and_gate and_gate_u_csamul_cla32_and21_15(.a(a[21]), .b(b[15]), .out(u_csamul_cla32_and21_15));
  fa fa_u_csamul_cla32_fa21_15_out(.a(u_csamul_cla32_and21_15[0]), .b(u_csamul_cla32_fa22_14_xor1[0]), .cin(u_csamul_cla32_fa21_14_or0[0]), .fa_xor1(u_csamul_cla32_fa21_15_xor1), .fa_or0(u_csamul_cla32_fa21_15_or0));
  and_gate and_gate_u_csamul_cla32_and22_15(.a(a[22]), .b(b[15]), .out(u_csamul_cla32_and22_15));
  fa fa_u_csamul_cla32_fa22_15_out(.a(u_csamul_cla32_and22_15[0]), .b(u_csamul_cla32_fa23_14_xor1[0]), .cin(u_csamul_cla32_fa22_14_or0[0]), .fa_xor1(u_csamul_cla32_fa22_15_xor1), .fa_or0(u_csamul_cla32_fa22_15_or0));
  and_gate and_gate_u_csamul_cla32_and23_15(.a(a[23]), .b(b[15]), .out(u_csamul_cla32_and23_15));
  fa fa_u_csamul_cla32_fa23_15_out(.a(u_csamul_cla32_and23_15[0]), .b(u_csamul_cla32_fa24_14_xor1[0]), .cin(u_csamul_cla32_fa23_14_or0[0]), .fa_xor1(u_csamul_cla32_fa23_15_xor1), .fa_or0(u_csamul_cla32_fa23_15_or0));
  and_gate and_gate_u_csamul_cla32_and24_15(.a(a[24]), .b(b[15]), .out(u_csamul_cla32_and24_15));
  fa fa_u_csamul_cla32_fa24_15_out(.a(u_csamul_cla32_and24_15[0]), .b(u_csamul_cla32_fa25_14_xor1[0]), .cin(u_csamul_cla32_fa24_14_or0[0]), .fa_xor1(u_csamul_cla32_fa24_15_xor1), .fa_or0(u_csamul_cla32_fa24_15_or0));
  and_gate and_gate_u_csamul_cla32_and25_15(.a(a[25]), .b(b[15]), .out(u_csamul_cla32_and25_15));
  fa fa_u_csamul_cla32_fa25_15_out(.a(u_csamul_cla32_and25_15[0]), .b(u_csamul_cla32_fa26_14_xor1[0]), .cin(u_csamul_cla32_fa25_14_or0[0]), .fa_xor1(u_csamul_cla32_fa25_15_xor1), .fa_or0(u_csamul_cla32_fa25_15_or0));
  and_gate and_gate_u_csamul_cla32_and26_15(.a(a[26]), .b(b[15]), .out(u_csamul_cla32_and26_15));
  fa fa_u_csamul_cla32_fa26_15_out(.a(u_csamul_cla32_and26_15[0]), .b(u_csamul_cla32_fa27_14_xor1[0]), .cin(u_csamul_cla32_fa26_14_or0[0]), .fa_xor1(u_csamul_cla32_fa26_15_xor1), .fa_or0(u_csamul_cla32_fa26_15_or0));
  and_gate and_gate_u_csamul_cla32_and27_15(.a(a[27]), .b(b[15]), .out(u_csamul_cla32_and27_15));
  fa fa_u_csamul_cla32_fa27_15_out(.a(u_csamul_cla32_and27_15[0]), .b(u_csamul_cla32_fa28_14_xor1[0]), .cin(u_csamul_cla32_fa27_14_or0[0]), .fa_xor1(u_csamul_cla32_fa27_15_xor1), .fa_or0(u_csamul_cla32_fa27_15_or0));
  and_gate and_gate_u_csamul_cla32_and28_15(.a(a[28]), .b(b[15]), .out(u_csamul_cla32_and28_15));
  fa fa_u_csamul_cla32_fa28_15_out(.a(u_csamul_cla32_and28_15[0]), .b(u_csamul_cla32_fa29_14_xor1[0]), .cin(u_csamul_cla32_fa28_14_or0[0]), .fa_xor1(u_csamul_cla32_fa28_15_xor1), .fa_or0(u_csamul_cla32_fa28_15_or0));
  and_gate and_gate_u_csamul_cla32_and29_15(.a(a[29]), .b(b[15]), .out(u_csamul_cla32_and29_15));
  fa fa_u_csamul_cla32_fa29_15_out(.a(u_csamul_cla32_and29_15[0]), .b(u_csamul_cla32_fa30_14_xor1[0]), .cin(u_csamul_cla32_fa29_14_or0[0]), .fa_xor1(u_csamul_cla32_fa29_15_xor1), .fa_or0(u_csamul_cla32_fa29_15_or0));
  and_gate and_gate_u_csamul_cla32_and30_15(.a(a[30]), .b(b[15]), .out(u_csamul_cla32_and30_15));
  fa fa_u_csamul_cla32_fa30_15_out(.a(u_csamul_cla32_and30_15[0]), .b(u_csamul_cla32_and31_14[0]), .cin(u_csamul_cla32_fa30_14_or0[0]), .fa_xor1(u_csamul_cla32_fa30_15_xor1), .fa_or0(u_csamul_cla32_fa30_15_or0));
  and_gate and_gate_u_csamul_cla32_and31_15(.a(a[31]), .b(b[15]), .out(u_csamul_cla32_and31_15));
  and_gate and_gate_u_csamul_cla32_and0_16(.a(a[0]), .b(b[16]), .out(u_csamul_cla32_and0_16));
  fa fa_u_csamul_cla32_fa0_16_out(.a(u_csamul_cla32_and0_16[0]), .b(u_csamul_cla32_fa1_15_xor1[0]), .cin(u_csamul_cla32_fa0_15_or0[0]), .fa_xor1(u_csamul_cla32_fa0_16_xor1), .fa_or0(u_csamul_cla32_fa0_16_or0));
  and_gate and_gate_u_csamul_cla32_and1_16(.a(a[1]), .b(b[16]), .out(u_csamul_cla32_and1_16));
  fa fa_u_csamul_cla32_fa1_16_out(.a(u_csamul_cla32_and1_16[0]), .b(u_csamul_cla32_fa2_15_xor1[0]), .cin(u_csamul_cla32_fa1_15_or0[0]), .fa_xor1(u_csamul_cla32_fa1_16_xor1), .fa_or0(u_csamul_cla32_fa1_16_or0));
  and_gate and_gate_u_csamul_cla32_and2_16(.a(a[2]), .b(b[16]), .out(u_csamul_cla32_and2_16));
  fa fa_u_csamul_cla32_fa2_16_out(.a(u_csamul_cla32_and2_16[0]), .b(u_csamul_cla32_fa3_15_xor1[0]), .cin(u_csamul_cla32_fa2_15_or0[0]), .fa_xor1(u_csamul_cla32_fa2_16_xor1), .fa_or0(u_csamul_cla32_fa2_16_or0));
  and_gate and_gate_u_csamul_cla32_and3_16(.a(a[3]), .b(b[16]), .out(u_csamul_cla32_and3_16));
  fa fa_u_csamul_cla32_fa3_16_out(.a(u_csamul_cla32_and3_16[0]), .b(u_csamul_cla32_fa4_15_xor1[0]), .cin(u_csamul_cla32_fa3_15_or0[0]), .fa_xor1(u_csamul_cla32_fa3_16_xor1), .fa_or0(u_csamul_cla32_fa3_16_or0));
  and_gate and_gate_u_csamul_cla32_and4_16(.a(a[4]), .b(b[16]), .out(u_csamul_cla32_and4_16));
  fa fa_u_csamul_cla32_fa4_16_out(.a(u_csamul_cla32_and4_16[0]), .b(u_csamul_cla32_fa5_15_xor1[0]), .cin(u_csamul_cla32_fa4_15_or0[0]), .fa_xor1(u_csamul_cla32_fa4_16_xor1), .fa_or0(u_csamul_cla32_fa4_16_or0));
  and_gate and_gate_u_csamul_cla32_and5_16(.a(a[5]), .b(b[16]), .out(u_csamul_cla32_and5_16));
  fa fa_u_csamul_cla32_fa5_16_out(.a(u_csamul_cla32_and5_16[0]), .b(u_csamul_cla32_fa6_15_xor1[0]), .cin(u_csamul_cla32_fa5_15_or0[0]), .fa_xor1(u_csamul_cla32_fa5_16_xor1), .fa_or0(u_csamul_cla32_fa5_16_or0));
  and_gate and_gate_u_csamul_cla32_and6_16(.a(a[6]), .b(b[16]), .out(u_csamul_cla32_and6_16));
  fa fa_u_csamul_cla32_fa6_16_out(.a(u_csamul_cla32_and6_16[0]), .b(u_csamul_cla32_fa7_15_xor1[0]), .cin(u_csamul_cla32_fa6_15_or0[0]), .fa_xor1(u_csamul_cla32_fa6_16_xor1), .fa_or0(u_csamul_cla32_fa6_16_or0));
  and_gate and_gate_u_csamul_cla32_and7_16(.a(a[7]), .b(b[16]), .out(u_csamul_cla32_and7_16));
  fa fa_u_csamul_cla32_fa7_16_out(.a(u_csamul_cla32_and7_16[0]), .b(u_csamul_cla32_fa8_15_xor1[0]), .cin(u_csamul_cla32_fa7_15_or0[0]), .fa_xor1(u_csamul_cla32_fa7_16_xor1), .fa_or0(u_csamul_cla32_fa7_16_or0));
  and_gate and_gate_u_csamul_cla32_and8_16(.a(a[8]), .b(b[16]), .out(u_csamul_cla32_and8_16));
  fa fa_u_csamul_cla32_fa8_16_out(.a(u_csamul_cla32_and8_16[0]), .b(u_csamul_cla32_fa9_15_xor1[0]), .cin(u_csamul_cla32_fa8_15_or0[0]), .fa_xor1(u_csamul_cla32_fa8_16_xor1), .fa_or0(u_csamul_cla32_fa8_16_or0));
  and_gate and_gate_u_csamul_cla32_and9_16(.a(a[9]), .b(b[16]), .out(u_csamul_cla32_and9_16));
  fa fa_u_csamul_cla32_fa9_16_out(.a(u_csamul_cla32_and9_16[0]), .b(u_csamul_cla32_fa10_15_xor1[0]), .cin(u_csamul_cla32_fa9_15_or0[0]), .fa_xor1(u_csamul_cla32_fa9_16_xor1), .fa_or0(u_csamul_cla32_fa9_16_or0));
  and_gate and_gate_u_csamul_cla32_and10_16(.a(a[10]), .b(b[16]), .out(u_csamul_cla32_and10_16));
  fa fa_u_csamul_cla32_fa10_16_out(.a(u_csamul_cla32_and10_16[0]), .b(u_csamul_cla32_fa11_15_xor1[0]), .cin(u_csamul_cla32_fa10_15_or0[0]), .fa_xor1(u_csamul_cla32_fa10_16_xor1), .fa_or0(u_csamul_cla32_fa10_16_or0));
  and_gate and_gate_u_csamul_cla32_and11_16(.a(a[11]), .b(b[16]), .out(u_csamul_cla32_and11_16));
  fa fa_u_csamul_cla32_fa11_16_out(.a(u_csamul_cla32_and11_16[0]), .b(u_csamul_cla32_fa12_15_xor1[0]), .cin(u_csamul_cla32_fa11_15_or0[0]), .fa_xor1(u_csamul_cla32_fa11_16_xor1), .fa_or0(u_csamul_cla32_fa11_16_or0));
  and_gate and_gate_u_csamul_cla32_and12_16(.a(a[12]), .b(b[16]), .out(u_csamul_cla32_and12_16));
  fa fa_u_csamul_cla32_fa12_16_out(.a(u_csamul_cla32_and12_16[0]), .b(u_csamul_cla32_fa13_15_xor1[0]), .cin(u_csamul_cla32_fa12_15_or0[0]), .fa_xor1(u_csamul_cla32_fa12_16_xor1), .fa_or0(u_csamul_cla32_fa12_16_or0));
  and_gate and_gate_u_csamul_cla32_and13_16(.a(a[13]), .b(b[16]), .out(u_csamul_cla32_and13_16));
  fa fa_u_csamul_cla32_fa13_16_out(.a(u_csamul_cla32_and13_16[0]), .b(u_csamul_cla32_fa14_15_xor1[0]), .cin(u_csamul_cla32_fa13_15_or0[0]), .fa_xor1(u_csamul_cla32_fa13_16_xor1), .fa_or0(u_csamul_cla32_fa13_16_or0));
  and_gate and_gate_u_csamul_cla32_and14_16(.a(a[14]), .b(b[16]), .out(u_csamul_cla32_and14_16));
  fa fa_u_csamul_cla32_fa14_16_out(.a(u_csamul_cla32_and14_16[0]), .b(u_csamul_cla32_fa15_15_xor1[0]), .cin(u_csamul_cla32_fa14_15_or0[0]), .fa_xor1(u_csamul_cla32_fa14_16_xor1), .fa_or0(u_csamul_cla32_fa14_16_or0));
  and_gate and_gate_u_csamul_cla32_and15_16(.a(a[15]), .b(b[16]), .out(u_csamul_cla32_and15_16));
  fa fa_u_csamul_cla32_fa15_16_out(.a(u_csamul_cla32_and15_16[0]), .b(u_csamul_cla32_fa16_15_xor1[0]), .cin(u_csamul_cla32_fa15_15_or0[0]), .fa_xor1(u_csamul_cla32_fa15_16_xor1), .fa_or0(u_csamul_cla32_fa15_16_or0));
  and_gate and_gate_u_csamul_cla32_and16_16(.a(a[16]), .b(b[16]), .out(u_csamul_cla32_and16_16));
  fa fa_u_csamul_cla32_fa16_16_out(.a(u_csamul_cla32_and16_16[0]), .b(u_csamul_cla32_fa17_15_xor1[0]), .cin(u_csamul_cla32_fa16_15_or0[0]), .fa_xor1(u_csamul_cla32_fa16_16_xor1), .fa_or0(u_csamul_cla32_fa16_16_or0));
  and_gate and_gate_u_csamul_cla32_and17_16(.a(a[17]), .b(b[16]), .out(u_csamul_cla32_and17_16));
  fa fa_u_csamul_cla32_fa17_16_out(.a(u_csamul_cla32_and17_16[0]), .b(u_csamul_cla32_fa18_15_xor1[0]), .cin(u_csamul_cla32_fa17_15_or0[0]), .fa_xor1(u_csamul_cla32_fa17_16_xor1), .fa_or0(u_csamul_cla32_fa17_16_or0));
  and_gate and_gate_u_csamul_cla32_and18_16(.a(a[18]), .b(b[16]), .out(u_csamul_cla32_and18_16));
  fa fa_u_csamul_cla32_fa18_16_out(.a(u_csamul_cla32_and18_16[0]), .b(u_csamul_cla32_fa19_15_xor1[0]), .cin(u_csamul_cla32_fa18_15_or0[0]), .fa_xor1(u_csamul_cla32_fa18_16_xor1), .fa_or0(u_csamul_cla32_fa18_16_or0));
  and_gate and_gate_u_csamul_cla32_and19_16(.a(a[19]), .b(b[16]), .out(u_csamul_cla32_and19_16));
  fa fa_u_csamul_cla32_fa19_16_out(.a(u_csamul_cla32_and19_16[0]), .b(u_csamul_cla32_fa20_15_xor1[0]), .cin(u_csamul_cla32_fa19_15_or0[0]), .fa_xor1(u_csamul_cla32_fa19_16_xor1), .fa_or0(u_csamul_cla32_fa19_16_or0));
  and_gate and_gate_u_csamul_cla32_and20_16(.a(a[20]), .b(b[16]), .out(u_csamul_cla32_and20_16));
  fa fa_u_csamul_cla32_fa20_16_out(.a(u_csamul_cla32_and20_16[0]), .b(u_csamul_cla32_fa21_15_xor1[0]), .cin(u_csamul_cla32_fa20_15_or0[0]), .fa_xor1(u_csamul_cla32_fa20_16_xor1), .fa_or0(u_csamul_cla32_fa20_16_or0));
  and_gate and_gate_u_csamul_cla32_and21_16(.a(a[21]), .b(b[16]), .out(u_csamul_cla32_and21_16));
  fa fa_u_csamul_cla32_fa21_16_out(.a(u_csamul_cla32_and21_16[0]), .b(u_csamul_cla32_fa22_15_xor1[0]), .cin(u_csamul_cla32_fa21_15_or0[0]), .fa_xor1(u_csamul_cla32_fa21_16_xor1), .fa_or0(u_csamul_cla32_fa21_16_or0));
  and_gate and_gate_u_csamul_cla32_and22_16(.a(a[22]), .b(b[16]), .out(u_csamul_cla32_and22_16));
  fa fa_u_csamul_cla32_fa22_16_out(.a(u_csamul_cla32_and22_16[0]), .b(u_csamul_cla32_fa23_15_xor1[0]), .cin(u_csamul_cla32_fa22_15_or0[0]), .fa_xor1(u_csamul_cla32_fa22_16_xor1), .fa_or0(u_csamul_cla32_fa22_16_or0));
  and_gate and_gate_u_csamul_cla32_and23_16(.a(a[23]), .b(b[16]), .out(u_csamul_cla32_and23_16));
  fa fa_u_csamul_cla32_fa23_16_out(.a(u_csamul_cla32_and23_16[0]), .b(u_csamul_cla32_fa24_15_xor1[0]), .cin(u_csamul_cla32_fa23_15_or0[0]), .fa_xor1(u_csamul_cla32_fa23_16_xor1), .fa_or0(u_csamul_cla32_fa23_16_or0));
  and_gate and_gate_u_csamul_cla32_and24_16(.a(a[24]), .b(b[16]), .out(u_csamul_cla32_and24_16));
  fa fa_u_csamul_cla32_fa24_16_out(.a(u_csamul_cla32_and24_16[0]), .b(u_csamul_cla32_fa25_15_xor1[0]), .cin(u_csamul_cla32_fa24_15_or0[0]), .fa_xor1(u_csamul_cla32_fa24_16_xor1), .fa_or0(u_csamul_cla32_fa24_16_or0));
  and_gate and_gate_u_csamul_cla32_and25_16(.a(a[25]), .b(b[16]), .out(u_csamul_cla32_and25_16));
  fa fa_u_csamul_cla32_fa25_16_out(.a(u_csamul_cla32_and25_16[0]), .b(u_csamul_cla32_fa26_15_xor1[0]), .cin(u_csamul_cla32_fa25_15_or0[0]), .fa_xor1(u_csamul_cla32_fa25_16_xor1), .fa_or0(u_csamul_cla32_fa25_16_or0));
  and_gate and_gate_u_csamul_cla32_and26_16(.a(a[26]), .b(b[16]), .out(u_csamul_cla32_and26_16));
  fa fa_u_csamul_cla32_fa26_16_out(.a(u_csamul_cla32_and26_16[0]), .b(u_csamul_cla32_fa27_15_xor1[0]), .cin(u_csamul_cla32_fa26_15_or0[0]), .fa_xor1(u_csamul_cla32_fa26_16_xor1), .fa_or0(u_csamul_cla32_fa26_16_or0));
  and_gate and_gate_u_csamul_cla32_and27_16(.a(a[27]), .b(b[16]), .out(u_csamul_cla32_and27_16));
  fa fa_u_csamul_cla32_fa27_16_out(.a(u_csamul_cla32_and27_16[0]), .b(u_csamul_cla32_fa28_15_xor1[0]), .cin(u_csamul_cla32_fa27_15_or0[0]), .fa_xor1(u_csamul_cla32_fa27_16_xor1), .fa_or0(u_csamul_cla32_fa27_16_or0));
  and_gate and_gate_u_csamul_cla32_and28_16(.a(a[28]), .b(b[16]), .out(u_csamul_cla32_and28_16));
  fa fa_u_csamul_cla32_fa28_16_out(.a(u_csamul_cla32_and28_16[0]), .b(u_csamul_cla32_fa29_15_xor1[0]), .cin(u_csamul_cla32_fa28_15_or0[0]), .fa_xor1(u_csamul_cla32_fa28_16_xor1), .fa_or0(u_csamul_cla32_fa28_16_or0));
  and_gate and_gate_u_csamul_cla32_and29_16(.a(a[29]), .b(b[16]), .out(u_csamul_cla32_and29_16));
  fa fa_u_csamul_cla32_fa29_16_out(.a(u_csamul_cla32_and29_16[0]), .b(u_csamul_cla32_fa30_15_xor1[0]), .cin(u_csamul_cla32_fa29_15_or0[0]), .fa_xor1(u_csamul_cla32_fa29_16_xor1), .fa_or0(u_csamul_cla32_fa29_16_or0));
  and_gate and_gate_u_csamul_cla32_and30_16(.a(a[30]), .b(b[16]), .out(u_csamul_cla32_and30_16));
  fa fa_u_csamul_cla32_fa30_16_out(.a(u_csamul_cla32_and30_16[0]), .b(u_csamul_cla32_and31_15[0]), .cin(u_csamul_cla32_fa30_15_or0[0]), .fa_xor1(u_csamul_cla32_fa30_16_xor1), .fa_or0(u_csamul_cla32_fa30_16_or0));
  and_gate and_gate_u_csamul_cla32_and31_16(.a(a[31]), .b(b[16]), .out(u_csamul_cla32_and31_16));
  and_gate and_gate_u_csamul_cla32_and0_17(.a(a[0]), .b(b[17]), .out(u_csamul_cla32_and0_17));
  fa fa_u_csamul_cla32_fa0_17_out(.a(u_csamul_cla32_and0_17[0]), .b(u_csamul_cla32_fa1_16_xor1[0]), .cin(u_csamul_cla32_fa0_16_or0[0]), .fa_xor1(u_csamul_cla32_fa0_17_xor1), .fa_or0(u_csamul_cla32_fa0_17_or0));
  and_gate and_gate_u_csamul_cla32_and1_17(.a(a[1]), .b(b[17]), .out(u_csamul_cla32_and1_17));
  fa fa_u_csamul_cla32_fa1_17_out(.a(u_csamul_cla32_and1_17[0]), .b(u_csamul_cla32_fa2_16_xor1[0]), .cin(u_csamul_cla32_fa1_16_or0[0]), .fa_xor1(u_csamul_cla32_fa1_17_xor1), .fa_or0(u_csamul_cla32_fa1_17_or0));
  and_gate and_gate_u_csamul_cla32_and2_17(.a(a[2]), .b(b[17]), .out(u_csamul_cla32_and2_17));
  fa fa_u_csamul_cla32_fa2_17_out(.a(u_csamul_cla32_and2_17[0]), .b(u_csamul_cla32_fa3_16_xor1[0]), .cin(u_csamul_cla32_fa2_16_or0[0]), .fa_xor1(u_csamul_cla32_fa2_17_xor1), .fa_or0(u_csamul_cla32_fa2_17_or0));
  and_gate and_gate_u_csamul_cla32_and3_17(.a(a[3]), .b(b[17]), .out(u_csamul_cla32_and3_17));
  fa fa_u_csamul_cla32_fa3_17_out(.a(u_csamul_cla32_and3_17[0]), .b(u_csamul_cla32_fa4_16_xor1[0]), .cin(u_csamul_cla32_fa3_16_or0[0]), .fa_xor1(u_csamul_cla32_fa3_17_xor1), .fa_or0(u_csamul_cla32_fa3_17_or0));
  and_gate and_gate_u_csamul_cla32_and4_17(.a(a[4]), .b(b[17]), .out(u_csamul_cla32_and4_17));
  fa fa_u_csamul_cla32_fa4_17_out(.a(u_csamul_cla32_and4_17[0]), .b(u_csamul_cla32_fa5_16_xor1[0]), .cin(u_csamul_cla32_fa4_16_or0[0]), .fa_xor1(u_csamul_cla32_fa4_17_xor1), .fa_or0(u_csamul_cla32_fa4_17_or0));
  and_gate and_gate_u_csamul_cla32_and5_17(.a(a[5]), .b(b[17]), .out(u_csamul_cla32_and5_17));
  fa fa_u_csamul_cla32_fa5_17_out(.a(u_csamul_cla32_and5_17[0]), .b(u_csamul_cla32_fa6_16_xor1[0]), .cin(u_csamul_cla32_fa5_16_or0[0]), .fa_xor1(u_csamul_cla32_fa5_17_xor1), .fa_or0(u_csamul_cla32_fa5_17_or0));
  and_gate and_gate_u_csamul_cla32_and6_17(.a(a[6]), .b(b[17]), .out(u_csamul_cla32_and6_17));
  fa fa_u_csamul_cla32_fa6_17_out(.a(u_csamul_cla32_and6_17[0]), .b(u_csamul_cla32_fa7_16_xor1[0]), .cin(u_csamul_cla32_fa6_16_or0[0]), .fa_xor1(u_csamul_cla32_fa6_17_xor1), .fa_or0(u_csamul_cla32_fa6_17_or0));
  and_gate and_gate_u_csamul_cla32_and7_17(.a(a[7]), .b(b[17]), .out(u_csamul_cla32_and7_17));
  fa fa_u_csamul_cla32_fa7_17_out(.a(u_csamul_cla32_and7_17[0]), .b(u_csamul_cla32_fa8_16_xor1[0]), .cin(u_csamul_cla32_fa7_16_or0[0]), .fa_xor1(u_csamul_cla32_fa7_17_xor1), .fa_or0(u_csamul_cla32_fa7_17_or0));
  and_gate and_gate_u_csamul_cla32_and8_17(.a(a[8]), .b(b[17]), .out(u_csamul_cla32_and8_17));
  fa fa_u_csamul_cla32_fa8_17_out(.a(u_csamul_cla32_and8_17[0]), .b(u_csamul_cla32_fa9_16_xor1[0]), .cin(u_csamul_cla32_fa8_16_or0[0]), .fa_xor1(u_csamul_cla32_fa8_17_xor1), .fa_or0(u_csamul_cla32_fa8_17_or0));
  and_gate and_gate_u_csamul_cla32_and9_17(.a(a[9]), .b(b[17]), .out(u_csamul_cla32_and9_17));
  fa fa_u_csamul_cla32_fa9_17_out(.a(u_csamul_cla32_and9_17[0]), .b(u_csamul_cla32_fa10_16_xor1[0]), .cin(u_csamul_cla32_fa9_16_or0[0]), .fa_xor1(u_csamul_cla32_fa9_17_xor1), .fa_or0(u_csamul_cla32_fa9_17_or0));
  and_gate and_gate_u_csamul_cla32_and10_17(.a(a[10]), .b(b[17]), .out(u_csamul_cla32_and10_17));
  fa fa_u_csamul_cla32_fa10_17_out(.a(u_csamul_cla32_and10_17[0]), .b(u_csamul_cla32_fa11_16_xor1[0]), .cin(u_csamul_cla32_fa10_16_or0[0]), .fa_xor1(u_csamul_cla32_fa10_17_xor1), .fa_or0(u_csamul_cla32_fa10_17_or0));
  and_gate and_gate_u_csamul_cla32_and11_17(.a(a[11]), .b(b[17]), .out(u_csamul_cla32_and11_17));
  fa fa_u_csamul_cla32_fa11_17_out(.a(u_csamul_cla32_and11_17[0]), .b(u_csamul_cla32_fa12_16_xor1[0]), .cin(u_csamul_cla32_fa11_16_or0[0]), .fa_xor1(u_csamul_cla32_fa11_17_xor1), .fa_or0(u_csamul_cla32_fa11_17_or0));
  and_gate and_gate_u_csamul_cla32_and12_17(.a(a[12]), .b(b[17]), .out(u_csamul_cla32_and12_17));
  fa fa_u_csamul_cla32_fa12_17_out(.a(u_csamul_cla32_and12_17[0]), .b(u_csamul_cla32_fa13_16_xor1[0]), .cin(u_csamul_cla32_fa12_16_or0[0]), .fa_xor1(u_csamul_cla32_fa12_17_xor1), .fa_or0(u_csamul_cla32_fa12_17_or0));
  and_gate and_gate_u_csamul_cla32_and13_17(.a(a[13]), .b(b[17]), .out(u_csamul_cla32_and13_17));
  fa fa_u_csamul_cla32_fa13_17_out(.a(u_csamul_cla32_and13_17[0]), .b(u_csamul_cla32_fa14_16_xor1[0]), .cin(u_csamul_cla32_fa13_16_or0[0]), .fa_xor1(u_csamul_cla32_fa13_17_xor1), .fa_or0(u_csamul_cla32_fa13_17_or0));
  and_gate and_gate_u_csamul_cla32_and14_17(.a(a[14]), .b(b[17]), .out(u_csamul_cla32_and14_17));
  fa fa_u_csamul_cla32_fa14_17_out(.a(u_csamul_cla32_and14_17[0]), .b(u_csamul_cla32_fa15_16_xor1[0]), .cin(u_csamul_cla32_fa14_16_or0[0]), .fa_xor1(u_csamul_cla32_fa14_17_xor1), .fa_or0(u_csamul_cla32_fa14_17_or0));
  and_gate and_gate_u_csamul_cla32_and15_17(.a(a[15]), .b(b[17]), .out(u_csamul_cla32_and15_17));
  fa fa_u_csamul_cla32_fa15_17_out(.a(u_csamul_cla32_and15_17[0]), .b(u_csamul_cla32_fa16_16_xor1[0]), .cin(u_csamul_cla32_fa15_16_or0[0]), .fa_xor1(u_csamul_cla32_fa15_17_xor1), .fa_or0(u_csamul_cla32_fa15_17_or0));
  and_gate and_gate_u_csamul_cla32_and16_17(.a(a[16]), .b(b[17]), .out(u_csamul_cla32_and16_17));
  fa fa_u_csamul_cla32_fa16_17_out(.a(u_csamul_cla32_and16_17[0]), .b(u_csamul_cla32_fa17_16_xor1[0]), .cin(u_csamul_cla32_fa16_16_or0[0]), .fa_xor1(u_csamul_cla32_fa16_17_xor1), .fa_or0(u_csamul_cla32_fa16_17_or0));
  and_gate and_gate_u_csamul_cla32_and17_17(.a(a[17]), .b(b[17]), .out(u_csamul_cla32_and17_17));
  fa fa_u_csamul_cla32_fa17_17_out(.a(u_csamul_cla32_and17_17[0]), .b(u_csamul_cla32_fa18_16_xor1[0]), .cin(u_csamul_cla32_fa17_16_or0[0]), .fa_xor1(u_csamul_cla32_fa17_17_xor1), .fa_or0(u_csamul_cla32_fa17_17_or0));
  and_gate and_gate_u_csamul_cla32_and18_17(.a(a[18]), .b(b[17]), .out(u_csamul_cla32_and18_17));
  fa fa_u_csamul_cla32_fa18_17_out(.a(u_csamul_cla32_and18_17[0]), .b(u_csamul_cla32_fa19_16_xor1[0]), .cin(u_csamul_cla32_fa18_16_or0[0]), .fa_xor1(u_csamul_cla32_fa18_17_xor1), .fa_or0(u_csamul_cla32_fa18_17_or0));
  and_gate and_gate_u_csamul_cla32_and19_17(.a(a[19]), .b(b[17]), .out(u_csamul_cla32_and19_17));
  fa fa_u_csamul_cla32_fa19_17_out(.a(u_csamul_cla32_and19_17[0]), .b(u_csamul_cla32_fa20_16_xor1[0]), .cin(u_csamul_cla32_fa19_16_or0[0]), .fa_xor1(u_csamul_cla32_fa19_17_xor1), .fa_or0(u_csamul_cla32_fa19_17_or0));
  and_gate and_gate_u_csamul_cla32_and20_17(.a(a[20]), .b(b[17]), .out(u_csamul_cla32_and20_17));
  fa fa_u_csamul_cla32_fa20_17_out(.a(u_csamul_cla32_and20_17[0]), .b(u_csamul_cla32_fa21_16_xor1[0]), .cin(u_csamul_cla32_fa20_16_or0[0]), .fa_xor1(u_csamul_cla32_fa20_17_xor1), .fa_or0(u_csamul_cla32_fa20_17_or0));
  and_gate and_gate_u_csamul_cla32_and21_17(.a(a[21]), .b(b[17]), .out(u_csamul_cla32_and21_17));
  fa fa_u_csamul_cla32_fa21_17_out(.a(u_csamul_cla32_and21_17[0]), .b(u_csamul_cla32_fa22_16_xor1[0]), .cin(u_csamul_cla32_fa21_16_or0[0]), .fa_xor1(u_csamul_cla32_fa21_17_xor1), .fa_or0(u_csamul_cla32_fa21_17_or0));
  and_gate and_gate_u_csamul_cla32_and22_17(.a(a[22]), .b(b[17]), .out(u_csamul_cla32_and22_17));
  fa fa_u_csamul_cla32_fa22_17_out(.a(u_csamul_cla32_and22_17[0]), .b(u_csamul_cla32_fa23_16_xor1[0]), .cin(u_csamul_cla32_fa22_16_or0[0]), .fa_xor1(u_csamul_cla32_fa22_17_xor1), .fa_or0(u_csamul_cla32_fa22_17_or0));
  and_gate and_gate_u_csamul_cla32_and23_17(.a(a[23]), .b(b[17]), .out(u_csamul_cla32_and23_17));
  fa fa_u_csamul_cla32_fa23_17_out(.a(u_csamul_cla32_and23_17[0]), .b(u_csamul_cla32_fa24_16_xor1[0]), .cin(u_csamul_cla32_fa23_16_or0[0]), .fa_xor1(u_csamul_cla32_fa23_17_xor1), .fa_or0(u_csamul_cla32_fa23_17_or0));
  and_gate and_gate_u_csamul_cla32_and24_17(.a(a[24]), .b(b[17]), .out(u_csamul_cla32_and24_17));
  fa fa_u_csamul_cla32_fa24_17_out(.a(u_csamul_cla32_and24_17[0]), .b(u_csamul_cla32_fa25_16_xor1[0]), .cin(u_csamul_cla32_fa24_16_or0[0]), .fa_xor1(u_csamul_cla32_fa24_17_xor1), .fa_or0(u_csamul_cla32_fa24_17_or0));
  and_gate and_gate_u_csamul_cla32_and25_17(.a(a[25]), .b(b[17]), .out(u_csamul_cla32_and25_17));
  fa fa_u_csamul_cla32_fa25_17_out(.a(u_csamul_cla32_and25_17[0]), .b(u_csamul_cla32_fa26_16_xor1[0]), .cin(u_csamul_cla32_fa25_16_or0[0]), .fa_xor1(u_csamul_cla32_fa25_17_xor1), .fa_or0(u_csamul_cla32_fa25_17_or0));
  and_gate and_gate_u_csamul_cla32_and26_17(.a(a[26]), .b(b[17]), .out(u_csamul_cla32_and26_17));
  fa fa_u_csamul_cla32_fa26_17_out(.a(u_csamul_cla32_and26_17[0]), .b(u_csamul_cla32_fa27_16_xor1[0]), .cin(u_csamul_cla32_fa26_16_or0[0]), .fa_xor1(u_csamul_cla32_fa26_17_xor1), .fa_or0(u_csamul_cla32_fa26_17_or0));
  and_gate and_gate_u_csamul_cla32_and27_17(.a(a[27]), .b(b[17]), .out(u_csamul_cla32_and27_17));
  fa fa_u_csamul_cla32_fa27_17_out(.a(u_csamul_cla32_and27_17[0]), .b(u_csamul_cla32_fa28_16_xor1[0]), .cin(u_csamul_cla32_fa27_16_or0[0]), .fa_xor1(u_csamul_cla32_fa27_17_xor1), .fa_or0(u_csamul_cla32_fa27_17_or0));
  and_gate and_gate_u_csamul_cla32_and28_17(.a(a[28]), .b(b[17]), .out(u_csamul_cla32_and28_17));
  fa fa_u_csamul_cla32_fa28_17_out(.a(u_csamul_cla32_and28_17[0]), .b(u_csamul_cla32_fa29_16_xor1[0]), .cin(u_csamul_cla32_fa28_16_or0[0]), .fa_xor1(u_csamul_cla32_fa28_17_xor1), .fa_or0(u_csamul_cla32_fa28_17_or0));
  and_gate and_gate_u_csamul_cla32_and29_17(.a(a[29]), .b(b[17]), .out(u_csamul_cla32_and29_17));
  fa fa_u_csamul_cla32_fa29_17_out(.a(u_csamul_cla32_and29_17[0]), .b(u_csamul_cla32_fa30_16_xor1[0]), .cin(u_csamul_cla32_fa29_16_or0[0]), .fa_xor1(u_csamul_cla32_fa29_17_xor1), .fa_or0(u_csamul_cla32_fa29_17_or0));
  and_gate and_gate_u_csamul_cla32_and30_17(.a(a[30]), .b(b[17]), .out(u_csamul_cla32_and30_17));
  fa fa_u_csamul_cla32_fa30_17_out(.a(u_csamul_cla32_and30_17[0]), .b(u_csamul_cla32_and31_16[0]), .cin(u_csamul_cla32_fa30_16_or0[0]), .fa_xor1(u_csamul_cla32_fa30_17_xor1), .fa_or0(u_csamul_cla32_fa30_17_or0));
  and_gate and_gate_u_csamul_cla32_and31_17(.a(a[31]), .b(b[17]), .out(u_csamul_cla32_and31_17));
  and_gate and_gate_u_csamul_cla32_and0_18(.a(a[0]), .b(b[18]), .out(u_csamul_cla32_and0_18));
  fa fa_u_csamul_cla32_fa0_18_out(.a(u_csamul_cla32_and0_18[0]), .b(u_csamul_cla32_fa1_17_xor1[0]), .cin(u_csamul_cla32_fa0_17_or0[0]), .fa_xor1(u_csamul_cla32_fa0_18_xor1), .fa_or0(u_csamul_cla32_fa0_18_or0));
  and_gate and_gate_u_csamul_cla32_and1_18(.a(a[1]), .b(b[18]), .out(u_csamul_cla32_and1_18));
  fa fa_u_csamul_cla32_fa1_18_out(.a(u_csamul_cla32_and1_18[0]), .b(u_csamul_cla32_fa2_17_xor1[0]), .cin(u_csamul_cla32_fa1_17_or0[0]), .fa_xor1(u_csamul_cla32_fa1_18_xor1), .fa_or0(u_csamul_cla32_fa1_18_or0));
  and_gate and_gate_u_csamul_cla32_and2_18(.a(a[2]), .b(b[18]), .out(u_csamul_cla32_and2_18));
  fa fa_u_csamul_cla32_fa2_18_out(.a(u_csamul_cla32_and2_18[0]), .b(u_csamul_cla32_fa3_17_xor1[0]), .cin(u_csamul_cla32_fa2_17_or0[0]), .fa_xor1(u_csamul_cla32_fa2_18_xor1), .fa_or0(u_csamul_cla32_fa2_18_or0));
  and_gate and_gate_u_csamul_cla32_and3_18(.a(a[3]), .b(b[18]), .out(u_csamul_cla32_and3_18));
  fa fa_u_csamul_cla32_fa3_18_out(.a(u_csamul_cla32_and3_18[0]), .b(u_csamul_cla32_fa4_17_xor1[0]), .cin(u_csamul_cla32_fa3_17_or0[0]), .fa_xor1(u_csamul_cla32_fa3_18_xor1), .fa_or0(u_csamul_cla32_fa3_18_or0));
  and_gate and_gate_u_csamul_cla32_and4_18(.a(a[4]), .b(b[18]), .out(u_csamul_cla32_and4_18));
  fa fa_u_csamul_cla32_fa4_18_out(.a(u_csamul_cla32_and4_18[0]), .b(u_csamul_cla32_fa5_17_xor1[0]), .cin(u_csamul_cla32_fa4_17_or0[0]), .fa_xor1(u_csamul_cla32_fa4_18_xor1), .fa_or0(u_csamul_cla32_fa4_18_or0));
  and_gate and_gate_u_csamul_cla32_and5_18(.a(a[5]), .b(b[18]), .out(u_csamul_cla32_and5_18));
  fa fa_u_csamul_cla32_fa5_18_out(.a(u_csamul_cla32_and5_18[0]), .b(u_csamul_cla32_fa6_17_xor1[0]), .cin(u_csamul_cla32_fa5_17_or0[0]), .fa_xor1(u_csamul_cla32_fa5_18_xor1), .fa_or0(u_csamul_cla32_fa5_18_or0));
  and_gate and_gate_u_csamul_cla32_and6_18(.a(a[6]), .b(b[18]), .out(u_csamul_cla32_and6_18));
  fa fa_u_csamul_cla32_fa6_18_out(.a(u_csamul_cla32_and6_18[0]), .b(u_csamul_cla32_fa7_17_xor1[0]), .cin(u_csamul_cla32_fa6_17_or0[0]), .fa_xor1(u_csamul_cla32_fa6_18_xor1), .fa_or0(u_csamul_cla32_fa6_18_or0));
  and_gate and_gate_u_csamul_cla32_and7_18(.a(a[7]), .b(b[18]), .out(u_csamul_cla32_and7_18));
  fa fa_u_csamul_cla32_fa7_18_out(.a(u_csamul_cla32_and7_18[0]), .b(u_csamul_cla32_fa8_17_xor1[0]), .cin(u_csamul_cla32_fa7_17_or0[0]), .fa_xor1(u_csamul_cla32_fa7_18_xor1), .fa_or0(u_csamul_cla32_fa7_18_or0));
  and_gate and_gate_u_csamul_cla32_and8_18(.a(a[8]), .b(b[18]), .out(u_csamul_cla32_and8_18));
  fa fa_u_csamul_cla32_fa8_18_out(.a(u_csamul_cla32_and8_18[0]), .b(u_csamul_cla32_fa9_17_xor1[0]), .cin(u_csamul_cla32_fa8_17_or0[0]), .fa_xor1(u_csamul_cla32_fa8_18_xor1), .fa_or0(u_csamul_cla32_fa8_18_or0));
  and_gate and_gate_u_csamul_cla32_and9_18(.a(a[9]), .b(b[18]), .out(u_csamul_cla32_and9_18));
  fa fa_u_csamul_cla32_fa9_18_out(.a(u_csamul_cla32_and9_18[0]), .b(u_csamul_cla32_fa10_17_xor1[0]), .cin(u_csamul_cla32_fa9_17_or0[0]), .fa_xor1(u_csamul_cla32_fa9_18_xor1), .fa_or0(u_csamul_cla32_fa9_18_or0));
  and_gate and_gate_u_csamul_cla32_and10_18(.a(a[10]), .b(b[18]), .out(u_csamul_cla32_and10_18));
  fa fa_u_csamul_cla32_fa10_18_out(.a(u_csamul_cla32_and10_18[0]), .b(u_csamul_cla32_fa11_17_xor1[0]), .cin(u_csamul_cla32_fa10_17_or0[0]), .fa_xor1(u_csamul_cla32_fa10_18_xor1), .fa_or0(u_csamul_cla32_fa10_18_or0));
  and_gate and_gate_u_csamul_cla32_and11_18(.a(a[11]), .b(b[18]), .out(u_csamul_cla32_and11_18));
  fa fa_u_csamul_cla32_fa11_18_out(.a(u_csamul_cla32_and11_18[0]), .b(u_csamul_cla32_fa12_17_xor1[0]), .cin(u_csamul_cla32_fa11_17_or0[0]), .fa_xor1(u_csamul_cla32_fa11_18_xor1), .fa_or0(u_csamul_cla32_fa11_18_or0));
  and_gate and_gate_u_csamul_cla32_and12_18(.a(a[12]), .b(b[18]), .out(u_csamul_cla32_and12_18));
  fa fa_u_csamul_cla32_fa12_18_out(.a(u_csamul_cla32_and12_18[0]), .b(u_csamul_cla32_fa13_17_xor1[0]), .cin(u_csamul_cla32_fa12_17_or0[0]), .fa_xor1(u_csamul_cla32_fa12_18_xor1), .fa_or0(u_csamul_cla32_fa12_18_or0));
  and_gate and_gate_u_csamul_cla32_and13_18(.a(a[13]), .b(b[18]), .out(u_csamul_cla32_and13_18));
  fa fa_u_csamul_cla32_fa13_18_out(.a(u_csamul_cla32_and13_18[0]), .b(u_csamul_cla32_fa14_17_xor1[0]), .cin(u_csamul_cla32_fa13_17_or0[0]), .fa_xor1(u_csamul_cla32_fa13_18_xor1), .fa_or0(u_csamul_cla32_fa13_18_or0));
  and_gate and_gate_u_csamul_cla32_and14_18(.a(a[14]), .b(b[18]), .out(u_csamul_cla32_and14_18));
  fa fa_u_csamul_cla32_fa14_18_out(.a(u_csamul_cla32_and14_18[0]), .b(u_csamul_cla32_fa15_17_xor1[0]), .cin(u_csamul_cla32_fa14_17_or0[0]), .fa_xor1(u_csamul_cla32_fa14_18_xor1), .fa_or0(u_csamul_cla32_fa14_18_or0));
  and_gate and_gate_u_csamul_cla32_and15_18(.a(a[15]), .b(b[18]), .out(u_csamul_cla32_and15_18));
  fa fa_u_csamul_cla32_fa15_18_out(.a(u_csamul_cla32_and15_18[0]), .b(u_csamul_cla32_fa16_17_xor1[0]), .cin(u_csamul_cla32_fa15_17_or0[0]), .fa_xor1(u_csamul_cla32_fa15_18_xor1), .fa_or0(u_csamul_cla32_fa15_18_or0));
  and_gate and_gate_u_csamul_cla32_and16_18(.a(a[16]), .b(b[18]), .out(u_csamul_cla32_and16_18));
  fa fa_u_csamul_cla32_fa16_18_out(.a(u_csamul_cla32_and16_18[0]), .b(u_csamul_cla32_fa17_17_xor1[0]), .cin(u_csamul_cla32_fa16_17_or0[0]), .fa_xor1(u_csamul_cla32_fa16_18_xor1), .fa_or0(u_csamul_cla32_fa16_18_or0));
  and_gate and_gate_u_csamul_cla32_and17_18(.a(a[17]), .b(b[18]), .out(u_csamul_cla32_and17_18));
  fa fa_u_csamul_cla32_fa17_18_out(.a(u_csamul_cla32_and17_18[0]), .b(u_csamul_cla32_fa18_17_xor1[0]), .cin(u_csamul_cla32_fa17_17_or0[0]), .fa_xor1(u_csamul_cla32_fa17_18_xor1), .fa_or0(u_csamul_cla32_fa17_18_or0));
  and_gate and_gate_u_csamul_cla32_and18_18(.a(a[18]), .b(b[18]), .out(u_csamul_cla32_and18_18));
  fa fa_u_csamul_cla32_fa18_18_out(.a(u_csamul_cla32_and18_18[0]), .b(u_csamul_cla32_fa19_17_xor1[0]), .cin(u_csamul_cla32_fa18_17_or0[0]), .fa_xor1(u_csamul_cla32_fa18_18_xor1), .fa_or0(u_csamul_cla32_fa18_18_or0));
  and_gate and_gate_u_csamul_cla32_and19_18(.a(a[19]), .b(b[18]), .out(u_csamul_cla32_and19_18));
  fa fa_u_csamul_cla32_fa19_18_out(.a(u_csamul_cla32_and19_18[0]), .b(u_csamul_cla32_fa20_17_xor1[0]), .cin(u_csamul_cla32_fa19_17_or0[0]), .fa_xor1(u_csamul_cla32_fa19_18_xor1), .fa_or0(u_csamul_cla32_fa19_18_or0));
  and_gate and_gate_u_csamul_cla32_and20_18(.a(a[20]), .b(b[18]), .out(u_csamul_cla32_and20_18));
  fa fa_u_csamul_cla32_fa20_18_out(.a(u_csamul_cla32_and20_18[0]), .b(u_csamul_cla32_fa21_17_xor1[0]), .cin(u_csamul_cla32_fa20_17_or0[0]), .fa_xor1(u_csamul_cla32_fa20_18_xor1), .fa_or0(u_csamul_cla32_fa20_18_or0));
  and_gate and_gate_u_csamul_cla32_and21_18(.a(a[21]), .b(b[18]), .out(u_csamul_cla32_and21_18));
  fa fa_u_csamul_cla32_fa21_18_out(.a(u_csamul_cla32_and21_18[0]), .b(u_csamul_cla32_fa22_17_xor1[0]), .cin(u_csamul_cla32_fa21_17_or0[0]), .fa_xor1(u_csamul_cla32_fa21_18_xor1), .fa_or0(u_csamul_cla32_fa21_18_or0));
  and_gate and_gate_u_csamul_cla32_and22_18(.a(a[22]), .b(b[18]), .out(u_csamul_cla32_and22_18));
  fa fa_u_csamul_cla32_fa22_18_out(.a(u_csamul_cla32_and22_18[0]), .b(u_csamul_cla32_fa23_17_xor1[0]), .cin(u_csamul_cla32_fa22_17_or0[0]), .fa_xor1(u_csamul_cla32_fa22_18_xor1), .fa_or0(u_csamul_cla32_fa22_18_or0));
  and_gate and_gate_u_csamul_cla32_and23_18(.a(a[23]), .b(b[18]), .out(u_csamul_cla32_and23_18));
  fa fa_u_csamul_cla32_fa23_18_out(.a(u_csamul_cla32_and23_18[0]), .b(u_csamul_cla32_fa24_17_xor1[0]), .cin(u_csamul_cla32_fa23_17_or0[0]), .fa_xor1(u_csamul_cla32_fa23_18_xor1), .fa_or0(u_csamul_cla32_fa23_18_or0));
  and_gate and_gate_u_csamul_cla32_and24_18(.a(a[24]), .b(b[18]), .out(u_csamul_cla32_and24_18));
  fa fa_u_csamul_cla32_fa24_18_out(.a(u_csamul_cla32_and24_18[0]), .b(u_csamul_cla32_fa25_17_xor1[0]), .cin(u_csamul_cla32_fa24_17_or0[0]), .fa_xor1(u_csamul_cla32_fa24_18_xor1), .fa_or0(u_csamul_cla32_fa24_18_or0));
  and_gate and_gate_u_csamul_cla32_and25_18(.a(a[25]), .b(b[18]), .out(u_csamul_cla32_and25_18));
  fa fa_u_csamul_cla32_fa25_18_out(.a(u_csamul_cla32_and25_18[0]), .b(u_csamul_cla32_fa26_17_xor1[0]), .cin(u_csamul_cla32_fa25_17_or0[0]), .fa_xor1(u_csamul_cla32_fa25_18_xor1), .fa_or0(u_csamul_cla32_fa25_18_or0));
  and_gate and_gate_u_csamul_cla32_and26_18(.a(a[26]), .b(b[18]), .out(u_csamul_cla32_and26_18));
  fa fa_u_csamul_cla32_fa26_18_out(.a(u_csamul_cla32_and26_18[0]), .b(u_csamul_cla32_fa27_17_xor1[0]), .cin(u_csamul_cla32_fa26_17_or0[0]), .fa_xor1(u_csamul_cla32_fa26_18_xor1), .fa_or0(u_csamul_cla32_fa26_18_or0));
  and_gate and_gate_u_csamul_cla32_and27_18(.a(a[27]), .b(b[18]), .out(u_csamul_cla32_and27_18));
  fa fa_u_csamul_cla32_fa27_18_out(.a(u_csamul_cla32_and27_18[0]), .b(u_csamul_cla32_fa28_17_xor1[0]), .cin(u_csamul_cla32_fa27_17_or0[0]), .fa_xor1(u_csamul_cla32_fa27_18_xor1), .fa_or0(u_csamul_cla32_fa27_18_or0));
  and_gate and_gate_u_csamul_cla32_and28_18(.a(a[28]), .b(b[18]), .out(u_csamul_cla32_and28_18));
  fa fa_u_csamul_cla32_fa28_18_out(.a(u_csamul_cla32_and28_18[0]), .b(u_csamul_cla32_fa29_17_xor1[0]), .cin(u_csamul_cla32_fa28_17_or0[0]), .fa_xor1(u_csamul_cla32_fa28_18_xor1), .fa_or0(u_csamul_cla32_fa28_18_or0));
  and_gate and_gate_u_csamul_cla32_and29_18(.a(a[29]), .b(b[18]), .out(u_csamul_cla32_and29_18));
  fa fa_u_csamul_cla32_fa29_18_out(.a(u_csamul_cla32_and29_18[0]), .b(u_csamul_cla32_fa30_17_xor1[0]), .cin(u_csamul_cla32_fa29_17_or0[0]), .fa_xor1(u_csamul_cla32_fa29_18_xor1), .fa_or0(u_csamul_cla32_fa29_18_or0));
  and_gate and_gate_u_csamul_cla32_and30_18(.a(a[30]), .b(b[18]), .out(u_csamul_cla32_and30_18));
  fa fa_u_csamul_cla32_fa30_18_out(.a(u_csamul_cla32_and30_18[0]), .b(u_csamul_cla32_and31_17[0]), .cin(u_csamul_cla32_fa30_17_or0[0]), .fa_xor1(u_csamul_cla32_fa30_18_xor1), .fa_or0(u_csamul_cla32_fa30_18_or0));
  and_gate and_gate_u_csamul_cla32_and31_18(.a(a[31]), .b(b[18]), .out(u_csamul_cla32_and31_18));
  and_gate and_gate_u_csamul_cla32_and0_19(.a(a[0]), .b(b[19]), .out(u_csamul_cla32_and0_19));
  fa fa_u_csamul_cla32_fa0_19_out(.a(u_csamul_cla32_and0_19[0]), .b(u_csamul_cla32_fa1_18_xor1[0]), .cin(u_csamul_cla32_fa0_18_or0[0]), .fa_xor1(u_csamul_cla32_fa0_19_xor1), .fa_or0(u_csamul_cla32_fa0_19_or0));
  and_gate and_gate_u_csamul_cla32_and1_19(.a(a[1]), .b(b[19]), .out(u_csamul_cla32_and1_19));
  fa fa_u_csamul_cla32_fa1_19_out(.a(u_csamul_cla32_and1_19[0]), .b(u_csamul_cla32_fa2_18_xor1[0]), .cin(u_csamul_cla32_fa1_18_or0[0]), .fa_xor1(u_csamul_cla32_fa1_19_xor1), .fa_or0(u_csamul_cla32_fa1_19_or0));
  and_gate and_gate_u_csamul_cla32_and2_19(.a(a[2]), .b(b[19]), .out(u_csamul_cla32_and2_19));
  fa fa_u_csamul_cla32_fa2_19_out(.a(u_csamul_cla32_and2_19[0]), .b(u_csamul_cla32_fa3_18_xor1[0]), .cin(u_csamul_cla32_fa2_18_or0[0]), .fa_xor1(u_csamul_cla32_fa2_19_xor1), .fa_or0(u_csamul_cla32_fa2_19_or0));
  and_gate and_gate_u_csamul_cla32_and3_19(.a(a[3]), .b(b[19]), .out(u_csamul_cla32_and3_19));
  fa fa_u_csamul_cla32_fa3_19_out(.a(u_csamul_cla32_and3_19[0]), .b(u_csamul_cla32_fa4_18_xor1[0]), .cin(u_csamul_cla32_fa3_18_or0[0]), .fa_xor1(u_csamul_cla32_fa3_19_xor1), .fa_or0(u_csamul_cla32_fa3_19_or0));
  and_gate and_gate_u_csamul_cla32_and4_19(.a(a[4]), .b(b[19]), .out(u_csamul_cla32_and4_19));
  fa fa_u_csamul_cla32_fa4_19_out(.a(u_csamul_cla32_and4_19[0]), .b(u_csamul_cla32_fa5_18_xor1[0]), .cin(u_csamul_cla32_fa4_18_or0[0]), .fa_xor1(u_csamul_cla32_fa4_19_xor1), .fa_or0(u_csamul_cla32_fa4_19_or0));
  and_gate and_gate_u_csamul_cla32_and5_19(.a(a[5]), .b(b[19]), .out(u_csamul_cla32_and5_19));
  fa fa_u_csamul_cla32_fa5_19_out(.a(u_csamul_cla32_and5_19[0]), .b(u_csamul_cla32_fa6_18_xor1[0]), .cin(u_csamul_cla32_fa5_18_or0[0]), .fa_xor1(u_csamul_cla32_fa5_19_xor1), .fa_or0(u_csamul_cla32_fa5_19_or0));
  and_gate and_gate_u_csamul_cla32_and6_19(.a(a[6]), .b(b[19]), .out(u_csamul_cla32_and6_19));
  fa fa_u_csamul_cla32_fa6_19_out(.a(u_csamul_cla32_and6_19[0]), .b(u_csamul_cla32_fa7_18_xor1[0]), .cin(u_csamul_cla32_fa6_18_or0[0]), .fa_xor1(u_csamul_cla32_fa6_19_xor1), .fa_or0(u_csamul_cla32_fa6_19_or0));
  and_gate and_gate_u_csamul_cla32_and7_19(.a(a[7]), .b(b[19]), .out(u_csamul_cla32_and7_19));
  fa fa_u_csamul_cla32_fa7_19_out(.a(u_csamul_cla32_and7_19[0]), .b(u_csamul_cla32_fa8_18_xor1[0]), .cin(u_csamul_cla32_fa7_18_or0[0]), .fa_xor1(u_csamul_cla32_fa7_19_xor1), .fa_or0(u_csamul_cla32_fa7_19_or0));
  and_gate and_gate_u_csamul_cla32_and8_19(.a(a[8]), .b(b[19]), .out(u_csamul_cla32_and8_19));
  fa fa_u_csamul_cla32_fa8_19_out(.a(u_csamul_cla32_and8_19[0]), .b(u_csamul_cla32_fa9_18_xor1[0]), .cin(u_csamul_cla32_fa8_18_or0[0]), .fa_xor1(u_csamul_cla32_fa8_19_xor1), .fa_or0(u_csamul_cla32_fa8_19_or0));
  and_gate and_gate_u_csamul_cla32_and9_19(.a(a[9]), .b(b[19]), .out(u_csamul_cla32_and9_19));
  fa fa_u_csamul_cla32_fa9_19_out(.a(u_csamul_cla32_and9_19[0]), .b(u_csamul_cla32_fa10_18_xor1[0]), .cin(u_csamul_cla32_fa9_18_or0[0]), .fa_xor1(u_csamul_cla32_fa9_19_xor1), .fa_or0(u_csamul_cla32_fa9_19_or0));
  and_gate and_gate_u_csamul_cla32_and10_19(.a(a[10]), .b(b[19]), .out(u_csamul_cla32_and10_19));
  fa fa_u_csamul_cla32_fa10_19_out(.a(u_csamul_cla32_and10_19[0]), .b(u_csamul_cla32_fa11_18_xor1[0]), .cin(u_csamul_cla32_fa10_18_or0[0]), .fa_xor1(u_csamul_cla32_fa10_19_xor1), .fa_or0(u_csamul_cla32_fa10_19_or0));
  and_gate and_gate_u_csamul_cla32_and11_19(.a(a[11]), .b(b[19]), .out(u_csamul_cla32_and11_19));
  fa fa_u_csamul_cla32_fa11_19_out(.a(u_csamul_cla32_and11_19[0]), .b(u_csamul_cla32_fa12_18_xor1[0]), .cin(u_csamul_cla32_fa11_18_or0[0]), .fa_xor1(u_csamul_cla32_fa11_19_xor1), .fa_or0(u_csamul_cla32_fa11_19_or0));
  and_gate and_gate_u_csamul_cla32_and12_19(.a(a[12]), .b(b[19]), .out(u_csamul_cla32_and12_19));
  fa fa_u_csamul_cla32_fa12_19_out(.a(u_csamul_cla32_and12_19[0]), .b(u_csamul_cla32_fa13_18_xor1[0]), .cin(u_csamul_cla32_fa12_18_or0[0]), .fa_xor1(u_csamul_cla32_fa12_19_xor1), .fa_or0(u_csamul_cla32_fa12_19_or0));
  and_gate and_gate_u_csamul_cla32_and13_19(.a(a[13]), .b(b[19]), .out(u_csamul_cla32_and13_19));
  fa fa_u_csamul_cla32_fa13_19_out(.a(u_csamul_cla32_and13_19[0]), .b(u_csamul_cla32_fa14_18_xor1[0]), .cin(u_csamul_cla32_fa13_18_or0[0]), .fa_xor1(u_csamul_cla32_fa13_19_xor1), .fa_or0(u_csamul_cla32_fa13_19_or0));
  and_gate and_gate_u_csamul_cla32_and14_19(.a(a[14]), .b(b[19]), .out(u_csamul_cla32_and14_19));
  fa fa_u_csamul_cla32_fa14_19_out(.a(u_csamul_cla32_and14_19[0]), .b(u_csamul_cla32_fa15_18_xor1[0]), .cin(u_csamul_cla32_fa14_18_or0[0]), .fa_xor1(u_csamul_cla32_fa14_19_xor1), .fa_or0(u_csamul_cla32_fa14_19_or0));
  and_gate and_gate_u_csamul_cla32_and15_19(.a(a[15]), .b(b[19]), .out(u_csamul_cla32_and15_19));
  fa fa_u_csamul_cla32_fa15_19_out(.a(u_csamul_cla32_and15_19[0]), .b(u_csamul_cla32_fa16_18_xor1[0]), .cin(u_csamul_cla32_fa15_18_or0[0]), .fa_xor1(u_csamul_cla32_fa15_19_xor1), .fa_or0(u_csamul_cla32_fa15_19_or0));
  and_gate and_gate_u_csamul_cla32_and16_19(.a(a[16]), .b(b[19]), .out(u_csamul_cla32_and16_19));
  fa fa_u_csamul_cla32_fa16_19_out(.a(u_csamul_cla32_and16_19[0]), .b(u_csamul_cla32_fa17_18_xor1[0]), .cin(u_csamul_cla32_fa16_18_or0[0]), .fa_xor1(u_csamul_cla32_fa16_19_xor1), .fa_or0(u_csamul_cla32_fa16_19_or0));
  and_gate and_gate_u_csamul_cla32_and17_19(.a(a[17]), .b(b[19]), .out(u_csamul_cla32_and17_19));
  fa fa_u_csamul_cla32_fa17_19_out(.a(u_csamul_cla32_and17_19[0]), .b(u_csamul_cla32_fa18_18_xor1[0]), .cin(u_csamul_cla32_fa17_18_or0[0]), .fa_xor1(u_csamul_cla32_fa17_19_xor1), .fa_or0(u_csamul_cla32_fa17_19_or0));
  and_gate and_gate_u_csamul_cla32_and18_19(.a(a[18]), .b(b[19]), .out(u_csamul_cla32_and18_19));
  fa fa_u_csamul_cla32_fa18_19_out(.a(u_csamul_cla32_and18_19[0]), .b(u_csamul_cla32_fa19_18_xor1[0]), .cin(u_csamul_cla32_fa18_18_or0[0]), .fa_xor1(u_csamul_cla32_fa18_19_xor1), .fa_or0(u_csamul_cla32_fa18_19_or0));
  and_gate and_gate_u_csamul_cla32_and19_19(.a(a[19]), .b(b[19]), .out(u_csamul_cla32_and19_19));
  fa fa_u_csamul_cla32_fa19_19_out(.a(u_csamul_cla32_and19_19[0]), .b(u_csamul_cla32_fa20_18_xor1[0]), .cin(u_csamul_cla32_fa19_18_or0[0]), .fa_xor1(u_csamul_cla32_fa19_19_xor1), .fa_or0(u_csamul_cla32_fa19_19_or0));
  and_gate and_gate_u_csamul_cla32_and20_19(.a(a[20]), .b(b[19]), .out(u_csamul_cla32_and20_19));
  fa fa_u_csamul_cla32_fa20_19_out(.a(u_csamul_cla32_and20_19[0]), .b(u_csamul_cla32_fa21_18_xor1[0]), .cin(u_csamul_cla32_fa20_18_or0[0]), .fa_xor1(u_csamul_cla32_fa20_19_xor1), .fa_or0(u_csamul_cla32_fa20_19_or0));
  and_gate and_gate_u_csamul_cla32_and21_19(.a(a[21]), .b(b[19]), .out(u_csamul_cla32_and21_19));
  fa fa_u_csamul_cla32_fa21_19_out(.a(u_csamul_cla32_and21_19[0]), .b(u_csamul_cla32_fa22_18_xor1[0]), .cin(u_csamul_cla32_fa21_18_or0[0]), .fa_xor1(u_csamul_cla32_fa21_19_xor1), .fa_or0(u_csamul_cla32_fa21_19_or0));
  and_gate and_gate_u_csamul_cla32_and22_19(.a(a[22]), .b(b[19]), .out(u_csamul_cla32_and22_19));
  fa fa_u_csamul_cla32_fa22_19_out(.a(u_csamul_cla32_and22_19[0]), .b(u_csamul_cla32_fa23_18_xor1[0]), .cin(u_csamul_cla32_fa22_18_or0[0]), .fa_xor1(u_csamul_cla32_fa22_19_xor1), .fa_or0(u_csamul_cla32_fa22_19_or0));
  and_gate and_gate_u_csamul_cla32_and23_19(.a(a[23]), .b(b[19]), .out(u_csamul_cla32_and23_19));
  fa fa_u_csamul_cla32_fa23_19_out(.a(u_csamul_cla32_and23_19[0]), .b(u_csamul_cla32_fa24_18_xor1[0]), .cin(u_csamul_cla32_fa23_18_or0[0]), .fa_xor1(u_csamul_cla32_fa23_19_xor1), .fa_or0(u_csamul_cla32_fa23_19_or0));
  and_gate and_gate_u_csamul_cla32_and24_19(.a(a[24]), .b(b[19]), .out(u_csamul_cla32_and24_19));
  fa fa_u_csamul_cla32_fa24_19_out(.a(u_csamul_cla32_and24_19[0]), .b(u_csamul_cla32_fa25_18_xor1[0]), .cin(u_csamul_cla32_fa24_18_or0[0]), .fa_xor1(u_csamul_cla32_fa24_19_xor1), .fa_or0(u_csamul_cla32_fa24_19_or0));
  and_gate and_gate_u_csamul_cla32_and25_19(.a(a[25]), .b(b[19]), .out(u_csamul_cla32_and25_19));
  fa fa_u_csamul_cla32_fa25_19_out(.a(u_csamul_cla32_and25_19[0]), .b(u_csamul_cla32_fa26_18_xor1[0]), .cin(u_csamul_cla32_fa25_18_or0[0]), .fa_xor1(u_csamul_cla32_fa25_19_xor1), .fa_or0(u_csamul_cla32_fa25_19_or0));
  and_gate and_gate_u_csamul_cla32_and26_19(.a(a[26]), .b(b[19]), .out(u_csamul_cla32_and26_19));
  fa fa_u_csamul_cla32_fa26_19_out(.a(u_csamul_cla32_and26_19[0]), .b(u_csamul_cla32_fa27_18_xor1[0]), .cin(u_csamul_cla32_fa26_18_or0[0]), .fa_xor1(u_csamul_cla32_fa26_19_xor1), .fa_or0(u_csamul_cla32_fa26_19_or0));
  and_gate and_gate_u_csamul_cla32_and27_19(.a(a[27]), .b(b[19]), .out(u_csamul_cla32_and27_19));
  fa fa_u_csamul_cla32_fa27_19_out(.a(u_csamul_cla32_and27_19[0]), .b(u_csamul_cla32_fa28_18_xor1[0]), .cin(u_csamul_cla32_fa27_18_or0[0]), .fa_xor1(u_csamul_cla32_fa27_19_xor1), .fa_or0(u_csamul_cla32_fa27_19_or0));
  and_gate and_gate_u_csamul_cla32_and28_19(.a(a[28]), .b(b[19]), .out(u_csamul_cla32_and28_19));
  fa fa_u_csamul_cla32_fa28_19_out(.a(u_csamul_cla32_and28_19[0]), .b(u_csamul_cla32_fa29_18_xor1[0]), .cin(u_csamul_cla32_fa28_18_or0[0]), .fa_xor1(u_csamul_cla32_fa28_19_xor1), .fa_or0(u_csamul_cla32_fa28_19_or0));
  and_gate and_gate_u_csamul_cla32_and29_19(.a(a[29]), .b(b[19]), .out(u_csamul_cla32_and29_19));
  fa fa_u_csamul_cla32_fa29_19_out(.a(u_csamul_cla32_and29_19[0]), .b(u_csamul_cla32_fa30_18_xor1[0]), .cin(u_csamul_cla32_fa29_18_or0[0]), .fa_xor1(u_csamul_cla32_fa29_19_xor1), .fa_or0(u_csamul_cla32_fa29_19_or0));
  and_gate and_gate_u_csamul_cla32_and30_19(.a(a[30]), .b(b[19]), .out(u_csamul_cla32_and30_19));
  fa fa_u_csamul_cla32_fa30_19_out(.a(u_csamul_cla32_and30_19[0]), .b(u_csamul_cla32_and31_18[0]), .cin(u_csamul_cla32_fa30_18_or0[0]), .fa_xor1(u_csamul_cla32_fa30_19_xor1), .fa_or0(u_csamul_cla32_fa30_19_or0));
  and_gate and_gate_u_csamul_cla32_and31_19(.a(a[31]), .b(b[19]), .out(u_csamul_cla32_and31_19));
  and_gate and_gate_u_csamul_cla32_and0_20(.a(a[0]), .b(b[20]), .out(u_csamul_cla32_and0_20));
  fa fa_u_csamul_cla32_fa0_20_out(.a(u_csamul_cla32_and0_20[0]), .b(u_csamul_cla32_fa1_19_xor1[0]), .cin(u_csamul_cla32_fa0_19_or0[0]), .fa_xor1(u_csamul_cla32_fa0_20_xor1), .fa_or0(u_csamul_cla32_fa0_20_or0));
  and_gate and_gate_u_csamul_cla32_and1_20(.a(a[1]), .b(b[20]), .out(u_csamul_cla32_and1_20));
  fa fa_u_csamul_cla32_fa1_20_out(.a(u_csamul_cla32_and1_20[0]), .b(u_csamul_cla32_fa2_19_xor1[0]), .cin(u_csamul_cla32_fa1_19_or0[0]), .fa_xor1(u_csamul_cla32_fa1_20_xor1), .fa_or0(u_csamul_cla32_fa1_20_or0));
  and_gate and_gate_u_csamul_cla32_and2_20(.a(a[2]), .b(b[20]), .out(u_csamul_cla32_and2_20));
  fa fa_u_csamul_cla32_fa2_20_out(.a(u_csamul_cla32_and2_20[0]), .b(u_csamul_cla32_fa3_19_xor1[0]), .cin(u_csamul_cla32_fa2_19_or0[0]), .fa_xor1(u_csamul_cla32_fa2_20_xor1), .fa_or0(u_csamul_cla32_fa2_20_or0));
  and_gate and_gate_u_csamul_cla32_and3_20(.a(a[3]), .b(b[20]), .out(u_csamul_cla32_and3_20));
  fa fa_u_csamul_cla32_fa3_20_out(.a(u_csamul_cla32_and3_20[0]), .b(u_csamul_cla32_fa4_19_xor1[0]), .cin(u_csamul_cla32_fa3_19_or0[0]), .fa_xor1(u_csamul_cla32_fa3_20_xor1), .fa_or0(u_csamul_cla32_fa3_20_or0));
  and_gate and_gate_u_csamul_cla32_and4_20(.a(a[4]), .b(b[20]), .out(u_csamul_cla32_and4_20));
  fa fa_u_csamul_cla32_fa4_20_out(.a(u_csamul_cla32_and4_20[0]), .b(u_csamul_cla32_fa5_19_xor1[0]), .cin(u_csamul_cla32_fa4_19_or0[0]), .fa_xor1(u_csamul_cla32_fa4_20_xor1), .fa_or0(u_csamul_cla32_fa4_20_or0));
  and_gate and_gate_u_csamul_cla32_and5_20(.a(a[5]), .b(b[20]), .out(u_csamul_cla32_and5_20));
  fa fa_u_csamul_cla32_fa5_20_out(.a(u_csamul_cla32_and5_20[0]), .b(u_csamul_cla32_fa6_19_xor1[0]), .cin(u_csamul_cla32_fa5_19_or0[0]), .fa_xor1(u_csamul_cla32_fa5_20_xor1), .fa_or0(u_csamul_cla32_fa5_20_or0));
  and_gate and_gate_u_csamul_cla32_and6_20(.a(a[6]), .b(b[20]), .out(u_csamul_cla32_and6_20));
  fa fa_u_csamul_cla32_fa6_20_out(.a(u_csamul_cla32_and6_20[0]), .b(u_csamul_cla32_fa7_19_xor1[0]), .cin(u_csamul_cla32_fa6_19_or0[0]), .fa_xor1(u_csamul_cla32_fa6_20_xor1), .fa_or0(u_csamul_cla32_fa6_20_or0));
  and_gate and_gate_u_csamul_cla32_and7_20(.a(a[7]), .b(b[20]), .out(u_csamul_cla32_and7_20));
  fa fa_u_csamul_cla32_fa7_20_out(.a(u_csamul_cla32_and7_20[0]), .b(u_csamul_cla32_fa8_19_xor1[0]), .cin(u_csamul_cla32_fa7_19_or0[0]), .fa_xor1(u_csamul_cla32_fa7_20_xor1), .fa_or0(u_csamul_cla32_fa7_20_or0));
  and_gate and_gate_u_csamul_cla32_and8_20(.a(a[8]), .b(b[20]), .out(u_csamul_cla32_and8_20));
  fa fa_u_csamul_cla32_fa8_20_out(.a(u_csamul_cla32_and8_20[0]), .b(u_csamul_cla32_fa9_19_xor1[0]), .cin(u_csamul_cla32_fa8_19_or0[0]), .fa_xor1(u_csamul_cla32_fa8_20_xor1), .fa_or0(u_csamul_cla32_fa8_20_or0));
  and_gate and_gate_u_csamul_cla32_and9_20(.a(a[9]), .b(b[20]), .out(u_csamul_cla32_and9_20));
  fa fa_u_csamul_cla32_fa9_20_out(.a(u_csamul_cla32_and9_20[0]), .b(u_csamul_cla32_fa10_19_xor1[0]), .cin(u_csamul_cla32_fa9_19_or0[0]), .fa_xor1(u_csamul_cla32_fa9_20_xor1), .fa_or0(u_csamul_cla32_fa9_20_or0));
  and_gate and_gate_u_csamul_cla32_and10_20(.a(a[10]), .b(b[20]), .out(u_csamul_cla32_and10_20));
  fa fa_u_csamul_cla32_fa10_20_out(.a(u_csamul_cla32_and10_20[0]), .b(u_csamul_cla32_fa11_19_xor1[0]), .cin(u_csamul_cla32_fa10_19_or0[0]), .fa_xor1(u_csamul_cla32_fa10_20_xor1), .fa_or0(u_csamul_cla32_fa10_20_or0));
  and_gate and_gate_u_csamul_cla32_and11_20(.a(a[11]), .b(b[20]), .out(u_csamul_cla32_and11_20));
  fa fa_u_csamul_cla32_fa11_20_out(.a(u_csamul_cla32_and11_20[0]), .b(u_csamul_cla32_fa12_19_xor1[0]), .cin(u_csamul_cla32_fa11_19_or0[0]), .fa_xor1(u_csamul_cla32_fa11_20_xor1), .fa_or0(u_csamul_cla32_fa11_20_or0));
  and_gate and_gate_u_csamul_cla32_and12_20(.a(a[12]), .b(b[20]), .out(u_csamul_cla32_and12_20));
  fa fa_u_csamul_cla32_fa12_20_out(.a(u_csamul_cla32_and12_20[0]), .b(u_csamul_cla32_fa13_19_xor1[0]), .cin(u_csamul_cla32_fa12_19_or0[0]), .fa_xor1(u_csamul_cla32_fa12_20_xor1), .fa_or0(u_csamul_cla32_fa12_20_or0));
  and_gate and_gate_u_csamul_cla32_and13_20(.a(a[13]), .b(b[20]), .out(u_csamul_cla32_and13_20));
  fa fa_u_csamul_cla32_fa13_20_out(.a(u_csamul_cla32_and13_20[0]), .b(u_csamul_cla32_fa14_19_xor1[0]), .cin(u_csamul_cla32_fa13_19_or0[0]), .fa_xor1(u_csamul_cla32_fa13_20_xor1), .fa_or0(u_csamul_cla32_fa13_20_or0));
  and_gate and_gate_u_csamul_cla32_and14_20(.a(a[14]), .b(b[20]), .out(u_csamul_cla32_and14_20));
  fa fa_u_csamul_cla32_fa14_20_out(.a(u_csamul_cla32_and14_20[0]), .b(u_csamul_cla32_fa15_19_xor1[0]), .cin(u_csamul_cla32_fa14_19_or0[0]), .fa_xor1(u_csamul_cla32_fa14_20_xor1), .fa_or0(u_csamul_cla32_fa14_20_or0));
  and_gate and_gate_u_csamul_cla32_and15_20(.a(a[15]), .b(b[20]), .out(u_csamul_cla32_and15_20));
  fa fa_u_csamul_cla32_fa15_20_out(.a(u_csamul_cla32_and15_20[0]), .b(u_csamul_cla32_fa16_19_xor1[0]), .cin(u_csamul_cla32_fa15_19_or0[0]), .fa_xor1(u_csamul_cla32_fa15_20_xor1), .fa_or0(u_csamul_cla32_fa15_20_or0));
  and_gate and_gate_u_csamul_cla32_and16_20(.a(a[16]), .b(b[20]), .out(u_csamul_cla32_and16_20));
  fa fa_u_csamul_cla32_fa16_20_out(.a(u_csamul_cla32_and16_20[0]), .b(u_csamul_cla32_fa17_19_xor1[0]), .cin(u_csamul_cla32_fa16_19_or0[0]), .fa_xor1(u_csamul_cla32_fa16_20_xor1), .fa_or0(u_csamul_cla32_fa16_20_or0));
  and_gate and_gate_u_csamul_cla32_and17_20(.a(a[17]), .b(b[20]), .out(u_csamul_cla32_and17_20));
  fa fa_u_csamul_cla32_fa17_20_out(.a(u_csamul_cla32_and17_20[0]), .b(u_csamul_cla32_fa18_19_xor1[0]), .cin(u_csamul_cla32_fa17_19_or0[0]), .fa_xor1(u_csamul_cla32_fa17_20_xor1), .fa_or0(u_csamul_cla32_fa17_20_or0));
  and_gate and_gate_u_csamul_cla32_and18_20(.a(a[18]), .b(b[20]), .out(u_csamul_cla32_and18_20));
  fa fa_u_csamul_cla32_fa18_20_out(.a(u_csamul_cla32_and18_20[0]), .b(u_csamul_cla32_fa19_19_xor1[0]), .cin(u_csamul_cla32_fa18_19_or0[0]), .fa_xor1(u_csamul_cla32_fa18_20_xor1), .fa_or0(u_csamul_cla32_fa18_20_or0));
  and_gate and_gate_u_csamul_cla32_and19_20(.a(a[19]), .b(b[20]), .out(u_csamul_cla32_and19_20));
  fa fa_u_csamul_cla32_fa19_20_out(.a(u_csamul_cla32_and19_20[0]), .b(u_csamul_cla32_fa20_19_xor1[0]), .cin(u_csamul_cla32_fa19_19_or0[0]), .fa_xor1(u_csamul_cla32_fa19_20_xor1), .fa_or0(u_csamul_cla32_fa19_20_or0));
  and_gate and_gate_u_csamul_cla32_and20_20(.a(a[20]), .b(b[20]), .out(u_csamul_cla32_and20_20));
  fa fa_u_csamul_cla32_fa20_20_out(.a(u_csamul_cla32_and20_20[0]), .b(u_csamul_cla32_fa21_19_xor1[0]), .cin(u_csamul_cla32_fa20_19_or0[0]), .fa_xor1(u_csamul_cla32_fa20_20_xor1), .fa_or0(u_csamul_cla32_fa20_20_or0));
  and_gate and_gate_u_csamul_cla32_and21_20(.a(a[21]), .b(b[20]), .out(u_csamul_cla32_and21_20));
  fa fa_u_csamul_cla32_fa21_20_out(.a(u_csamul_cla32_and21_20[0]), .b(u_csamul_cla32_fa22_19_xor1[0]), .cin(u_csamul_cla32_fa21_19_or0[0]), .fa_xor1(u_csamul_cla32_fa21_20_xor1), .fa_or0(u_csamul_cla32_fa21_20_or0));
  and_gate and_gate_u_csamul_cla32_and22_20(.a(a[22]), .b(b[20]), .out(u_csamul_cla32_and22_20));
  fa fa_u_csamul_cla32_fa22_20_out(.a(u_csamul_cla32_and22_20[0]), .b(u_csamul_cla32_fa23_19_xor1[0]), .cin(u_csamul_cla32_fa22_19_or0[0]), .fa_xor1(u_csamul_cla32_fa22_20_xor1), .fa_or0(u_csamul_cla32_fa22_20_or0));
  and_gate and_gate_u_csamul_cla32_and23_20(.a(a[23]), .b(b[20]), .out(u_csamul_cla32_and23_20));
  fa fa_u_csamul_cla32_fa23_20_out(.a(u_csamul_cla32_and23_20[0]), .b(u_csamul_cla32_fa24_19_xor1[0]), .cin(u_csamul_cla32_fa23_19_or0[0]), .fa_xor1(u_csamul_cla32_fa23_20_xor1), .fa_or0(u_csamul_cla32_fa23_20_or0));
  and_gate and_gate_u_csamul_cla32_and24_20(.a(a[24]), .b(b[20]), .out(u_csamul_cla32_and24_20));
  fa fa_u_csamul_cla32_fa24_20_out(.a(u_csamul_cla32_and24_20[0]), .b(u_csamul_cla32_fa25_19_xor1[0]), .cin(u_csamul_cla32_fa24_19_or0[0]), .fa_xor1(u_csamul_cla32_fa24_20_xor1), .fa_or0(u_csamul_cla32_fa24_20_or0));
  and_gate and_gate_u_csamul_cla32_and25_20(.a(a[25]), .b(b[20]), .out(u_csamul_cla32_and25_20));
  fa fa_u_csamul_cla32_fa25_20_out(.a(u_csamul_cla32_and25_20[0]), .b(u_csamul_cla32_fa26_19_xor1[0]), .cin(u_csamul_cla32_fa25_19_or0[0]), .fa_xor1(u_csamul_cla32_fa25_20_xor1), .fa_or0(u_csamul_cla32_fa25_20_or0));
  and_gate and_gate_u_csamul_cla32_and26_20(.a(a[26]), .b(b[20]), .out(u_csamul_cla32_and26_20));
  fa fa_u_csamul_cla32_fa26_20_out(.a(u_csamul_cla32_and26_20[0]), .b(u_csamul_cla32_fa27_19_xor1[0]), .cin(u_csamul_cla32_fa26_19_or0[0]), .fa_xor1(u_csamul_cla32_fa26_20_xor1), .fa_or0(u_csamul_cla32_fa26_20_or0));
  and_gate and_gate_u_csamul_cla32_and27_20(.a(a[27]), .b(b[20]), .out(u_csamul_cla32_and27_20));
  fa fa_u_csamul_cla32_fa27_20_out(.a(u_csamul_cla32_and27_20[0]), .b(u_csamul_cla32_fa28_19_xor1[0]), .cin(u_csamul_cla32_fa27_19_or0[0]), .fa_xor1(u_csamul_cla32_fa27_20_xor1), .fa_or0(u_csamul_cla32_fa27_20_or0));
  and_gate and_gate_u_csamul_cla32_and28_20(.a(a[28]), .b(b[20]), .out(u_csamul_cla32_and28_20));
  fa fa_u_csamul_cla32_fa28_20_out(.a(u_csamul_cla32_and28_20[0]), .b(u_csamul_cla32_fa29_19_xor1[0]), .cin(u_csamul_cla32_fa28_19_or0[0]), .fa_xor1(u_csamul_cla32_fa28_20_xor1), .fa_or0(u_csamul_cla32_fa28_20_or0));
  and_gate and_gate_u_csamul_cla32_and29_20(.a(a[29]), .b(b[20]), .out(u_csamul_cla32_and29_20));
  fa fa_u_csamul_cla32_fa29_20_out(.a(u_csamul_cla32_and29_20[0]), .b(u_csamul_cla32_fa30_19_xor1[0]), .cin(u_csamul_cla32_fa29_19_or0[0]), .fa_xor1(u_csamul_cla32_fa29_20_xor1), .fa_or0(u_csamul_cla32_fa29_20_or0));
  and_gate and_gate_u_csamul_cla32_and30_20(.a(a[30]), .b(b[20]), .out(u_csamul_cla32_and30_20));
  fa fa_u_csamul_cla32_fa30_20_out(.a(u_csamul_cla32_and30_20[0]), .b(u_csamul_cla32_and31_19[0]), .cin(u_csamul_cla32_fa30_19_or0[0]), .fa_xor1(u_csamul_cla32_fa30_20_xor1), .fa_or0(u_csamul_cla32_fa30_20_or0));
  and_gate and_gate_u_csamul_cla32_and31_20(.a(a[31]), .b(b[20]), .out(u_csamul_cla32_and31_20));
  and_gate and_gate_u_csamul_cla32_and0_21(.a(a[0]), .b(b[21]), .out(u_csamul_cla32_and0_21));
  fa fa_u_csamul_cla32_fa0_21_out(.a(u_csamul_cla32_and0_21[0]), .b(u_csamul_cla32_fa1_20_xor1[0]), .cin(u_csamul_cla32_fa0_20_or0[0]), .fa_xor1(u_csamul_cla32_fa0_21_xor1), .fa_or0(u_csamul_cla32_fa0_21_or0));
  and_gate and_gate_u_csamul_cla32_and1_21(.a(a[1]), .b(b[21]), .out(u_csamul_cla32_and1_21));
  fa fa_u_csamul_cla32_fa1_21_out(.a(u_csamul_cla32_and1_21[0]), .b(u_csamul_cla32_fa2_20_xor1[0]), .cin(u_csamul_cla32_fa1_20_or0[0]), .fa_xor1(u_csamul_cla32_fa1_21_xor1), .fa_or0(u_csamul_cla32_fa1_21_or0));
  and_gate and_gate_u_csamul_cla32_and2_21(.a(a[2]), .b(b[21]), .out(u_csamul_cla32_and2_21));
  fa fa_u_csamul_cla32_fa2_21_out(.a(u_csamul_cla32_and2_21[0]), .b(u_csamul_cla32_fa3_20_xor1[0]), .cin(u_csamul_cla32_fa2_20_or0[0]), .fa_xor1(u_csamul_cla32_fa2_21_xor1), .fa_or0(u_csamul_cla32_fa2_21_or0));
  and_gate and_gate_u_csamul_cla32_and3_21(.a(a[3]), .b(b[21]), .out(u_csamul_cla32_and3_21));
  fa fa_u_csamul_cla32_fa3_21_out(.a(u_csamul_cla32_and3_21[0]), .b(u_csamul_cla32_fa4_20_xor1[0]), .cin(u_csamul_cla32_fa3_20_or0[0]), .fa_xor1(u_csamul_cla32_fa3_21_xor1), .fa_or0(u_csamul_cla32_fa3_21_or0));
  and_gate and_gate_u_csamul_cla32_and4_21(.a(a[4]), .b(b[21]), .out(u_csamul_cla32_and4_21));
  fa fa_u_csamul_cla32_fa4_21_out(.a(u_csamul_cla32_and4_21[0]), .b(u_csamul_cla32_fa5_20_xor1[0]), .cin(u_csamul_cla32_fa4_20_or0[0]), .fa_xor1(u_csamul_cla32_fa4_21_xor1), .fa_or0(u_csamul_cla32_fa4_21_or0));
  and_gate and_gate_u_csamul_cla32_and5_21(.a(a[5]), .b(b[21]), .out(u_csamul_cla32_and5_21));
  fa fa_u_csamul_cla32_fa5_21_out(.a(u_csamul_cla32_and5_21[0]), .b(u_csamul_cla32_fa6_20_xor1[0]), .cin(u_csamul_cla32_fa5_20_or0[0]), .fa_xor1(u_csamul_cla32_fa5_21_xor1), .fa_or0(u_csamul_cla32_fa5_21_or0));
  and_gate and_gate_u_csamul_cla32_and6_21(.a(a[6]), .b(b[21]), .out(u_csamul_cla32_and6_21));
  fa fa_u_csamul_cla32_fa6_21_out(.a(u_csamul_cla32_and6_21[0]), .b(u_csamul_cla32_fa7_20_xor1[0]), .cin(u_csamul_cla32_fa6_20_or0[0]), .fa_xor1(u_csamul_cla32_fa6_21_xor1), .fa_or0(u_csamul_cla32_fa6_21_or0));
  and_gate and_gate_u_csamul_cla32_and7_21(.a(a[7]), .b(b[21]), .out(u_csamul_cla32_and7_21));
  fa fa_u_csamul_cla32_fa7_21_out(.a(u_csamul_cla32_and7_21[0]), .b(u_csamul_cla32_fa8_20_xor1[0]), .cin(u_csamul_cla32_fa7_20_or0[0]), .fa_xor1(u_csamul_cla32_fa7_21_xor1), .fa_or0(u_csamul_cla32_fa7_21_or0));
  and_gate and_gate_u_csamul_cla32_and8_21(.a(a[8]), .b(b[21]), .out(u_csamul_cla32_and8_21));
  fa fa_u_csamul_cla32_fa8_21_out(.a(u_csamul_cla32_and8_21[0]), .b(u_csamul_cla32_fa9_20_xor1[0]), .cin(u_csamul_cla32_fa8_20_or0[0]), .fa_xor1(u_csamul_cla32_fa8_21_xor1), .fa_or0(u_csamul_cla32_fa8_21_or0));
  and_gate and_gate_u_csamul_cla32_and9_21(.a(a[9]), .b(b[21]), .out(u_csamul_cla32_and9_21));
  fa fa_u_csamul_cla32_fa9_21_out(.a(u_csamul_cla32_and9_21[0]), .b(u_csamul_cla32_fa10_20_xor1[0]), .cin(u_csamul_cla32_fa9_20_or0[0]), .fa_xor1(u_csamul_cla32_fa9_21_xor1), .fa_or0(u_csamul_cla32_fa9_21_or0));
  and_gate and_gate_u_csamul_cla32_and10_21(.a(a[10]), .b(b[21]), .out(u_csamul_cla32_and10_21));
  fa fa_u_csamul_cla32_fa10_21_out(.a(u_csamul_cla32_and10_21[0]), .b(u_csamul_cla32_fa11_20_xor1[0]), .cin(u_csamul_cla32_fa10_20_or0[0]), .fa_xor1(u_csamul_cla32_fa10_21_xor1), .fa_or0(u_csamul_cla32_fa10_21_or0));
  and_gate and_gate_u_csamul_cla32_and11_21(.a(a[11]), .b(b[21]), .out(u_csamul_cla32_and11_21));
  fa fa_u_csamul_cla32_fa11_21_out(.a(u_csamul_cla32_and11_21[0]), .b(u_csamul_cla32_fa12_20_xor1[0]), .cin(u_csamul_cla32_fa11_20_or0[0]), .fa_xor1(u_csamul_cla32_fa11_21_xor1), .fa_or0(u_csamul_cla32_fa11_21_or0));
  and_gate and_gate_u_csamul_cla32_and12_21(.a(a[12]), .b(b[21]), .out(u_csamul_cla32_and12_21));
  fa fa_u_csamul_cla32_fa12_21_out(.a(u_csamul_cla32_and12_21[0]), .b(u_csamul_cla32_fa13_20_xor1[0]), .cin(u_csamul_cla32_fa12_20_or0[0]), .fa_xor1(u_csamul_cla32_fa12_21_xor1), .fa_or0(u_csamul_cla32_fa12_21_or0));
  and_gate and_gate_u_csamul_cla32_and13_21(.a(a[13]), .b(b[21]), .out(u_csamul_cla32_and13_21));
  fa fa_u_csamul_cla32_fa13_21_out(.a(u_csamul_cla32_and13_21[0]), .b(u_csamul_cla32_fa14_20_xor1[0]), .cin(u_csamul_cla32_fa13_20_or0[0]), .fa_xor1(u_csamul_cla32_fa13_21_xor1), .fa_or0(u_csamul_cla32_fa13_21_or0));
  and_gate and_gate_u_csamul_cla32_and14_21(.a(a[14]), .b(b[21]), .out(u_csamul_cla32_and14_21));
  fa fa_u_csamul_cla32_fa14_21_out(.a(u_csamul_cla32_and14_21[0]), .b(u_csamul_cla32_fa15_20_xor1[0]), .cin(u_csamul_cla32_fa14_20_or0[0]), .fa_xor1(u_csamul_cla32_fa14_21_xor1), .fa_or0(u_csamul_cla32_fa14_21_or0));
  and_gate and_gate_u_csamul_cla32_and15_21(.a(a[15]), .b(b[21]), .out(u_csamul_cla32_and15_21));
  fa fa_u_csamul_cla32_fa15_21_out(.a(u_csamul_cla32_and15_21[0]), .b(u_csamul_cla32_fa16_20_xor1[0]), .cin(u_csamul_cla32_fa15_20_or0[0]), .fa_xor1(u_csamul_cla32_fa15_21_xor1), .fa_or0(u_csamul_cla32_fa15_21_or0));
  and_gate and_gate_u_csamul_cla32_and16_21(.a(a[16]), .b(b[21]), .out(u_csamul_cla32_and16_21));
  fa fa_u_csamul_cla32_fa16_21_out(.a(u_csamul_cla32_and16_21[0]), .b(u_csamul_cla32_fa17_20_xor1[0]), .cin(u_csamul_cla32_fa16_20_or0[0]), .fa_xor1(u_csamul_cla32_fa16_21_xor1), .fa_or0(u_csamul_cla32_fa16_21_or0));
  and_gate and_gate_u_csamul_cla32_and17_21(.a(a[17]), .b(b[21]), .out(u_csamul_cla32_and17_21));
  fa fa_u_csamul_cla32_fa17_21_out(.a(u_csamul_cla32_and17_21[0]), .b(u_csamul_cla32_fa18_20_xor1[0]), .cin(u_csamul_cla32_fa17_20_or0[0]), .fa_xor1(u_csamul_cla32_fa17_21_xor1), .fa_or0(u_csamul_cla32_fa17_21_or0));
  and_gate and_gate_u_csamul_cla32_and18_21(.a(a[18]), .b(b[21]), .out(u_csamul_cla32_and18_21));
  fa fa_u_csamul_cla32_fa18_21_out(.a(u_csamul_cla32_and18_21[0]), .b(u_csamul_cla32_fa19_20_xor1[0]), .cin(u_csamul_cla32_fa18_20_or0[0]), .fa_xor1(u_csamul_cla32_fa18_21_xor1), .fa_or0(u_csamul_cla32_fa18_21_or0));
  and_gate and_gate_u_csamul_cla32_and19_21(.a(a[19]), .b(b[21]), .out(u_csamul_cla32_and19_21));
  fa fa_u_csamul_cla32_fa19_21_out(.a(u_csamul_cla32_and19_21[0]), .b(u_csamul_cla32_fa20_20_xor1[0]), .cin(u_csamul_cla32_fa19_20_or0[0]), .fa_xor1(u_csamul_cla32_fa19_21_xor1), .fa_or0(u_csamul_cla32_fa19_21_or0));
  and_gate and_gate_u_csamul_cla32_and20_21(.a(a[20]), .b(b[21]), .out(u_csamul_cla32_and20_21));
  fa fa_u_csamul_cla32_fa20_21_out(.a(u_csamul_cla32_and20_21[0]), .b(u_csamul_cla32_fa21_20_xor1[0]), .cin(u_csamul_cla32_fa20_20_or0[0]), .fa_xor1(u_csamul_cla32_fa20_21_xor1), .fa_or0(u_csamul_cla32_fa20_21_or0));
  and_gate and_gate_u_csamul_cla32_and21_21(.a(a[21]), .b(b[21]), .out(u_csamul_cla32_and21_21));
  fa fa_u_csamul_cla32_fa21_21_out(.a(u_csamul_cla32_and21_21[0]), .b(u_csamul_cla32_fa22_20_xor1[0]), .cin(u_csamul_cla32_fa21_20_or0[0]), .fa_xor1(u_csamul_cla32_fa21_21_xor1), .fa_or0(u_csamul_cla32_fa21_21_or0));
  and_gate and_gate_u_csamul_cla32_and22_21(.a(a[22]), .b(b[21]), .out(u_csamul_cla32_and22_21));
  fa fa_u_csamul_cla32_fa22_21_out(.a(u_csamul_cla32_and22_21[0]), .b(u_csamul_cla32_fa23_20_xor1[0]), .cin(u_csamul_cla32_fa22_20_or0[0]), .fa_xor1(u_csamul_cla32_fa22_21_xor1), .fa_or0(u_csamul_cla32_fa22_21_or0));
  and_gate and_gate_u_csamul_cla32_and23_21(.a(a[23]), .b(b[21]), .out(u_csamul_cla32_and23_21));
  fa fa_u_csamul_cla32_fa23_21_out(.a(u_csamul_cla32_and23_21[0]), .b(u_csamul_cla32_fa24_20_xor1[0]), .cin(u_csamul_cla32_fa23_20_or0[0]), .fa_xor1(u_csamul_cla32_fa23_21_xor1), .fa_or0(u_csamul_cla32_fa23_21_or0));
  and_gate and_gate_u_csamul_cla32_and24_21(.a(a[24]), .b(b[21]), .out(u_csamul_cla32_and24_21));
  fa fa_u_csamul_cla32_fa24_21_out(.a(u_csamul_cla32_and24_21[0]), .b(u_csamul_cla32_fa25_20_xor1[0]), .cin(u_csamul_cla32_fa24_20_or0[0]), .fa_xor1(u_csamul_cla32_fa24_21_xor1), .fa_or0(u_csamul_cla32_fa24_21_or0));
  and_gate and_gate_u_csamul_cla32_and25_21(.a(a[25]), .b(b[21]), .out(u_csamul_cla32_and25_21));
  fa fa_u_csamul_cla32_fa25_21_out(.a(u_csamul_cla32_and25_21[0]), .b(u_csamul_cla32_fa26_20_xor1[0]), .cin(u_csamul_cla32_fa25_20_or0[0]), .fa_xor1(u_csamul_cla32_fa25_21_xor1), .fa_or0(u_csamul_cla32_fa25_21_or0));
  and_gate and_gate_u_csamul_cla32_and26_21(.a(a[26]), .b(b[21]), .out(u_csamul_cla32_and26_21));
  fa fa_u_csamul_cla32_fa26_21_out(.a(u_csamul_cla32_and26_21[0]), .b(u_csamul_cla32_fa27_20_xor1[0]), .cin(u_csamul_cla32_fa26_20_or0[0]), .fa_xor1(u_csamul_cla32_fa26_21_xor1), .fa_or0(u_csamul_cla32_fa26_21_or0));
  and_gate and_gate_u_csamul_cla32_and27_21(.a(a[27]), .b(b[21]), .out(u_csamul_cla32_and27_21));
  fa fa_u_csamul_cla32_fa27_21_out(.a(u_csamul_cla32_and27_21[0]), .b(u_csamul_cla32_fa28_20_xor1[0]), .cin(u_csamul_cla32_fa27_20_or0[0]), .fa_xor1(u_csamul_cla32_fa27_21_xor1), .fa_or0(u_csamul_cla32_fa27_21_or0));
  and_gate and_gate_u_csamul_cla32_and28_21(.a(a[28]), .b(b[21]), .out(u_csamul_cla32_and28_21));
  fa fa_u_csamul_cla32_fa28_21_out(.a(u_csamul_cla32_and28_21[0]), .b(u_csamul_cla32_fa29_20_xor1[0]), .cin(u_csamul_cla32_fa28_20_or0[0]), .fa_xor1(u_csamul_cla32_fa28_21_xor1), .fa_or0(u_csamul_cla32_fa28_21_or0));
  and_gate and_gate_u_csamul_cla32_and29_21(.a(a[29]), .b(b[21]), .out(u_csamul_cla32_and29_21));
  fa fa_u_csamul_cla32_fa29_21_out(.a(u_csamul_cla32_and29_21[0]), .b(u_csamul_cla32_fa30_20_xor1[0]), .cin(u_csamul_cla32_fa29_20_or0[0]), .fa_xor1(u_csamul_cla32_fa29_21_xor1), .fa_or0(u_csamul_cla32_fa29_21_or0));
  and_gate and_gate_u_csamul_cla32_and30_21(.a(a[30]), .b(b[21]), .out(u_csamul_cla32_and30_21));
  fa fa_u_csamul_cla32_fa30_21_out(.a(u_csamul_cla32_and30_21[0]), .b(u_csamul_cla32_and31_20[0]), .cin(u_csamul_cla32_fa30_20_or0[0]), .fa_xor1(u_csamul_cla32_fa30_21_xor1), .fa_or0(u_csamul_cla32_fa30_21_or0));
  and_gate and_gate_u_csamul_cla32_and31_21(.a(a[31]), .b(b[21]), .out(u_csamul_cla32_and31_21));
  and_gate and_gate_u_csamul_cla32_and0_22(.a(a[0]), .b(b[22]), .out(u_csamul_cla32_and0_22));
  fa fa_u_csamul_cla32_fa0_22_out(.a(u_csamul_cla32_and0_22[0]), .b(u_csamul_cla32_fa1_21_xor1[0]), .cin(u_csamul_cla32_fa0_21_or0[0]), .fa_xor1(u_csamul_cla32_fa0_22_xor1), .fa_or0(u_csamul_cla32_fa0_22_or0));
  and_gate and_gate_u_csamul_cla32_and1_22(.a(a[1]), .b(b[22]), .out(u_csamul_cla32_and1_22));
  fa fa_u_csamul_cla32_fa1_22_out(.a(u_csamul_cla32_and1_22[0]), .b(u_csamul_cla32_fa2_21_xor1[0]), .cin(u_csamul_cla32_fa1_21_or0[0]), .fa_xor1(u_csamul_cla32_fa1_22_xor1), .fa_or0(u_csamul_cla32_fa1_22_or0));
  and_gate and_gate_u_csamul_cla32_and2_22(.a(a[2]), .b(b[22]), .out(u_csamul_cla32_and2_22));
  fa fa_u_csamul_cla32_fa2_22_out(.a(u_csamul_cla32_and2_22[0]), .b(u_csamul_cla32_fa3_21_xor1[0]), .cin(u_csamul_cla32_fa2_21_or0[0]), .fa_xor1(u_csamul_cla32_fa2_22_xor1), .fa_or0(u_csamul_cla32_fa2_22_or0));
  and_gate and_gate_u_csamul_cla32_and3_22(.a(a[3]), .b(b[22]), .out(u_csamul_cla32_and3_22));
  fa fa_u_csamul_cla32_fa3_22_out(.a(u_csamul_cla32_and3_22[0]), .b(u_csamul_cla32_fa4_21_xor1[0]), .cin(u_csamul_cla32_fa3_21_or0[0]), .fa_xor1(u_csamul_cla32_fa3_22_xor1), .fa_or0(u_csamul_cla32_fa3_22_or0));
  and_gate and_gate_u_csamul_cla32_and4_22(.a(a[4]), .b(b[22]), .out(u_csamul_cla32_and4_22));
  fa fa_u_csamul_cla32_fa4_22_out(.a(u_csamul_cla32_and4_22[0]), .b(u_csamul_cla32_fa5_21_xor1[0]), .cin(u_csamul_cla32_fa4_21_or0[0]), .fa_xor1(u_csamul_cla32_fa4_22_xor1), .fa_or0(u_csamul_cla32_fa4_22_or0));
  and_gate and_gate_u_csamul_cla32_and5_22(.a(a[5]), .b(b[22]), .out(u_csamul_cla32_and5_22));
  fa fa_u_csamul_cla32_fa5_22_out(.a(u_csamul_cla32_and5_22[0]), .b(u_csamul_cla32_fa6_21_xor1[0]), .cin(u_csamul_cla32_fa5_21_or0[0]), .fa_xor1(u_csamul_cla32_fa5_22_xor1), .fa_or0(u_csamul_cla32_fa5_22_or0));
  and_gate and_gate_u_csamul_cla32_and6_22(.a(a[6]), .b(b[22]), .out(u_csamul_cla32_and6_22));
  fa fa_u_csamul_cla32_fa6_22_out(.a(u_csamul_cla32_and6_22[0]), .b(u_csamul_cla32_fa7_21_xor1[0]), .cin(u_csamul_cla32_fa6_21_or0[0]), .fa_xor1(u_csamul_cla32_fa6_22_xor1), .fa_or0(u_csamul_cla32_fa6_22_or0));
  and_gate and_gate_u_csamul_cla32_and7_22(.a(a[7]), .b(b[22]), .out(u_csamul_cla32_and7_22));
  fa fa_u_csamul_cla32_fa7_22_out(.a(u_csamul_cla32_and7_22[0]), .b(u_csamul_cla32_fa8_21_xor1[0]), .cin(u_csamul_cla32_fa7_21_or0[0]), .fa_xor1(u_csamul_cla32_fa7_22_xor1), .fa_or0(u_csamul_cla32_fa7_22_or0));
  and_gate and_gate_u_csamul_cla32_and8_22(.a(a[8]), .b(b[22]), .out(u_csamul_cla32_and8_22));
  fa fa_u_csamul_cla32_fa8_22_out(.a(u_csamul_cla32_and8_22[0]), .b(u_csamul_cla32_fa9_21_xor1[0]), .cin(u_csamul_cla32_fa8_21_or0[0]), .fa_xor1(u_csamul_cla32_fa8_22_xor1), .fa_or0(u_csamul_cla32_fa8_22_or0));
  and_gate and_gate_u_csamul_cla32_and9_22(.a(a[9]), .b(b[22]), .out(u_csamul_cla32_and9_22));
  fa fa_u_csamul_cla32_fa9_22_out(.a(u_csamul_cla32_and9_22[0]), .b(u_csamul_cla32_fa10_21_xor1[0]), .cin(u_csamul_cla32_fa9_21_or0[0]), .fa_xor1(u_csamul_cla32_fa9_22_xor1), .fa_or0(u_csamul_cla32_fa9_22_or0));
  and_gate and_gate_u_csamul_cla32_and10_22(.a(a[10]), .b(b[22]), .out(u_csamul_cla32_and10_22));
  fa fa_u_csamul_cla32_fa10_22_out(.a(u_csamul_cla32_and10_22[0]), .b(u_csamul_cla32_fa11_21_xor1[0]), .cin(u_csamul_cla32_fa10_21_or0[0]), .fa_xor1(u_csamul_cla32_fa10_22_xor1), .fa_or0(u_csamul_cla32_fa10_22_or0));
  and_gate and_gate_u_csamul_cla32_and11_22(.a(a[11]), .b(b[22]), .out(u_csamul_cla32_and11_22));
  fa fa_u_csamul_cla32_fa11_22_out(.a(u_csamul_cla32_and11_22[0]), .b(u_csamul_cla32_fa12_21_xor1[0]), .cin(u_csamul_cla32_fa11_21_or0[0]), .fa_xor1(u_csamul_cla32_fa11_22_xor1), .fa_or0(u_csamul_cla32_fa11_22_or0));
  and_gate and_gate_u_csamul_cla32_and12_22(.a(a[12]), .b(b[22]), .out(u_csamul_cla32_and12_22));
  fa fa_u_csamul_cla32_fa12_22_out(.a(u_csamul_cla32_and12_22[0]), .b(u_csamul_cla32_fa13_21_xor1[0]), .cin(u_csamul_cla32_fa12_21_or0[0]), .fa_xor1(u_csamul_cla32_fa12_22_xor1), .fa_or0(u_csamul_cla32_fa12_22_or0));
  and_gate and_gate_u_csamul_cla32_and13_22(.a(a[13]), .b(b[22]), .out(u_csamul_cla32_and13_22));
  fa fa_u_csamul_cla32_fa13_22_out(.a(u_csamul_cla32_and13_22[0]), .b(u_csamul_cla32_fa14_21_xor1[0]), .cin(u_csamul_cla32_fa13_21_or0[0]), .fa_xor1(u_csamul_cla32_fa13_22_xor1), .fa_or0(u_csamul_cla32_fa13_22_or0));
  and_gate and_gate_u_csamul_cla32_and14_22(.a(a[14]), .b(b[22]), .out(u_csamul_cla32_and14_22));
  fa fa_u_csamul_cla32_fa14_22_out(.a(u_csamul_cla32_and14_22[0]), .b(u_csamul_cla32_fa15_21_xor1[0]), .cin(u_csamul_cla32_fa14_21_or0[0]), .fa_xor1(u_csamul_cla32_fa14_22_xor1), .fa_or0(u_csamul_cla32_fa14_22_or0));
  and_gate and_gate_u_csamul_cla32_and15_22(.a(a[15]), .b(b[22]), .out(u_csamul_cla32_and15_22));
  fa fa_u_csamul_cla32_fa15_22_out(.a(u_csamul_cla32_and15_22[0]), .b(u_csamul_cla32_fa16_21_xor1[0]), .cin(u_csamul_cla32_fa15_21_or0[0]), .fa_xor1(u_csamul_cla32_fa15_22_xor1), .fa_or0(u_csamul_cla32_fa15_22_or0));
  and_gate and_gate_u_csamul_cla32_and16_22(.a(a[16]), .b(b[22]), .out(u_csamul_cla32_and16_22));
  fa fa_u_csamul_cla32_fa16_22_out(.a(u_csamul_cla32_and16_22[0]), .b(u_csamul_cla32_fa17_21_xor1[0]), .cin(u_csamul_cla32_fa16_21_or0[0]), .fa_xor1(u_csamul_cla32_fa16_22_xor1), .fa_or0(u_csamul_cla32_fa16_22_or0));
  and_gate and_gate_u_csamul_cla32_and17_22(.a(a[17]), .b(b[22]), .out(u_csamul_cla32_and17_22));
  fa fa_u_csamul_cla32_fa17_22_out(.a(u_csamul_cla32_and17_22[0]), .b(u_csamul_cla32_fa18_21_xor1[0]), .cin(u_csamul_cla32_fa17_21_or0[0]), .fa_xor1(u_csamul_cla32_fa17_22_xor1), .fa_or0(u_csamul_cla32_fa17_22_or0));
  and_gate and_gate_u_csamul_cla32_and18_22(.a(a[18]), .b(b[22]), .out(u_csamul_cla32_and18_22));
  fa fa_u_csamul_cla32_fa18_22_out(.a(u_csamul_cla32_and18_22[0]), .b(u_csamul_cla32_fa19_21_xor1[0]), .cin(u_csamul_cla32_fa18_21_or0[0]), .fa_xor1(u_csamul_cla32_fa18_22_xor1), .fa_or0(u_csamul_cla32_fa18_22_or0));
  and_gate and_gate_u_csamul_cla32_and19_22(.a(a[19]), .b(b[22]), .out(u_csamul_cla32_and19_22));
  fa fa_u_csamul_cla32_fa19_22_out(.a(u_csamul_cla32_and19_22[0]), .b(u_csamul_cla32_fa20_21_xor1[0]), .cin(u_csamul_cla32_fa19_21_or0[0]), .fa_xor1(u_csamul_cla32_fa19_22_xor1), .fa_or0(u_csamul_cla32_fa19_22_or0));
  and_gate and_gate_u_csamul_cla32_and20_22(.a(a[20]), .b(b[22]), .out(u_csamul_cla32_and20_22));
  fa fa_u_csamul_cla32_fa20_22_out(.a(u_csamul_cla32_and20_22[0]), .b(u_csamul_cla32_fa21_21_xor1[0]), .cin(u_csamul_cla32_fa20_21_or0[0]), .fa_xor1(u_csamul_cla32_fa20_22_xor1), .fa_or0(u_csamul_cla32_fa20_22_or0));
  and_gate and_gate_u_csamul_cla32_and21_22(.a(a[21]), .b(b[22]), .out(u_csamul_cla32_and21_22));
  fa fa_u_csamul_cla32_fa21_22_out(.a(u_csamul_cla32_and21_22[0]), .b(u_csamul_cla32_fa22_21_xor1[0]), .cin(u_csamul_cla32_fa21_21_or0[0]), .fa_xor1(u_csamul_cla32_fa21_22_xor1), .fa_or0(u_csamul_cla32_fa21_22_or0));
  and_gate and_gate_u_csamul_cla32_and22_22(.a(a[22]), .b(b[22]), .out(u_csamul_cla32_and22_22));
  fa fa_u_csamul_cla32_fa22_22_out(.a(u_csamul_cla32_and22_22[0]), .b(u_csamul_cla32_fa23_21_xor1[0]), .cin(u_csamul_cla32_fa22_21_or0[0]), .fa_xor1(u_csamul_cla32_fa22_22_xor1), .fa_or0(u_csamul_cla32_fa22_22_or0));
  and_gate and_gate_u_csamul_cla32_and23_22(.a(a[23]), .b(b[22]), .out(u_csamul_cla32_and23_22));
  fa fa_u_csamul_cla32_fa23_22_out(.a(u_csamul_cla32_and23_22[0]), .b(u_csamul_cla32_fa24_21_xor1[0]), .cin(u_csamul_cla32_fa23_21_or0[0]), .fa_xor1(u_csamul_cla32_fa23_22_xor1), .fa_or0(u_csamul_cla32_fa23_22_or0));
  and_gate and_gate_u_csamul_cla32_and24_22(.a(a[24]), .b(b[22]), .out(u_csamul_cla32_and24_22));
  fa fa_u_csamul_cla32_fa24_22_out(.a(u_csamul_cla32_and24_22[0]), .b(u_csamul_cla32_fa25_21_xor1[0]), .cin(u_csamul_cla32_fa24_21_or0[0]), .fa_xor1(u_csamul_cla32_fa24_22_xor1), .fa_or0(u_csamul_cla32_fa24_22_or0));
  and_gate and_gate_u_csamul_cla32_and25_22(.a(a[25]), .b(b[22]), .out(u_csamul_cla32_and25_22));
  fa fa_u_csamul_cla32_fa25_22_out(.a(u_csamul_cla32_and25_22[0]), .b(u_csamul_cla32_fa26_21_xor1[0]), .cin(u_csamul_cla32_fa25_21_or0[0]), .fa_xor1(u_csamul_cla32_fa25_22_xor1), .fa_or0(u_csamul_cla32_fa25_22_or0));
  and_gate and_gate_u_csamul_cla32_and26_22(.a(a[26]), .b(b[22]), .out(u_csamul_cla32_and26_22));
  fa fa_u_csamul_cla32_fa26_22_out(.a(u_csamul_cla32_and26_22[0]), .b(u_csamul_cla32_fa27_21_xor1[0]), .cin(u_csamul_cla32_fa26_21_or0[0]), .fa_xor1(u_csamul_cla32_fa26_22_xor1), .fa_or0(u_csamul_cla32_fa26_22_or0));
  and_gate and_gate_u_csamul_cla32_and27_22(.a(a[27]), .b(b[22]), .out(u_csamul_cla32_and27_22));
  fa fa_u_csamul_cla32_fa27_22_out(.a(u_csamul_cla32_and27_22[0]), .b(u_csamul_cla32_fa28_21_xor1[0]), .cin(u_csamul_cla32_fa27_21_or0[0]), .fa_xor1(u_csamul_cla32_fa27_22_xor1), .fa_or0(u_csamul_cla32_fa27_22_or0));
  and_gate and_gate_u_csamul_cla32_and28_22(.a(a[28]), .b(b[22]), .out(u_csamul_cla32_and28_22));
  fa fa_u_csamul_cla32_fa28_22_out(.a(u_csamul_cla32_and28_22[0]), .b(u_csamul_cla32_fa29_21_xor1[0]), .cin(u_csamul_cla32_fa28_21_or0[0]), .fa_xor1(u_csamul_cla32_fa28_22_xor1), .fa_or0(u_csamul_cla32_fa28_22_or0));
  and_gate and_gate_u_csamul_cla32_and29_22(.a(a[29]), .b(b[22]), .out(u_csamul_cla32_and29_22));
  fa fa_u_csamul_cla32_fa29_22_out(.a(u_csamul_cla32_and29_22[0]), .b(u_csamul_cla32_fa30_21_xor1[0]), .cin(u_csamul_cla32_fa29_21_or0[0]), .fa_xor1(u_csamul_cla32_fa29_22_xor1), .fa_or0(u_csamul_cla32_fa29_22_or0));
  and_gate and_gate_u_csamul_cla32_and30_22(.a(a[30]), .b(b[22]), .out(u_csamul_cla32_and30_22));
  fa fa_u_csamul_cla32_fa30_22_out(.a(u_csamul_cla32_and30_22[0]), .b(u_csamul_cla32_and31_21[0]), .cin(u_csamul_cla32_fa30_21_or0[0]), .fa_xor1(u_csamul_cla32_fa30_22_xor1), .fa_or0(u_csamul_cla32_fa30_22_or0));
  and_gate and_gate_u_csamul_cla32_and31_22(.a(a[31]), .b(b[22]), .out(u_csamul_cla32_and31_22));
  and_gate and_gate_u_csamul_cla32_and0_23(.a(a[0]), .b(b[23]), .out(u_csamul_cla32_and0_23));
  fa fa_u_csamul_cla32_fa0_23_out(.a(u_csamul_cla32_and0_23[0]), .b(u_csamul_cla32_fa1_22_xor1[0]), .cin(u_csamul_cla32_fa0_22_or0[0]), .fa_xor1(u_csamul_cla32_fa0_23_xor1), .fa_or0(u_csamul_cla32_fa0_23_or0));
  and_gate and_gate_u_csamul_cla32_and1_23(.a(a[1]), .b(b[23]), .out(u_csamul_cla32_and1_23));
  fa fa_u_csamul_cla32_fa1_23_out(.a(u_csamul_cla32_and1_23[0]), .b(u_csamul_cla32_fa2_22_xor1[0]), .cin(u_csamul_cla32_fa1_22_or0[0]), .fa_xor1(u_csamul_cla32_fa1_23_xor1), .fa_or0(u_csamul_cla32_fa1_23_or0));
  and_gate and_gate_u_csamul_cla32_and2_23(.a(a[2]), .b(b[23]), .out(u_csamul_cla32_and2_23));
  fa fa_u_csamul_cla32_fa2_23_out(.a(u_csamul_cla32_and2_23[0]), .b(u_csamul_cla32_fa3_22_xor1[0]), .cin(u_csamul_cla32_fa2_22_or0[0]), .fa_xor1(u_csamul_cla32_fa2_23_xor1), .fa_or0(u_csamul_cla32_fa2_23_or0));
  and_gate and_gate_u_csamul_cla32_and3_23(.a(a[3]), .b(b[23]), .out(u_csamul_cla32_and3_23));
  fa fa_u_csamul_cla32_fa3_23_out(.a(u_csamul_cla32_and3_23[0]), .b(u_csamul_cla32_fa4_22_xor1[0]), .cin(u_csamul_cla32_fa3_22_or0[0]), .fa_xor1(u_csamul_cla32_fa3_23_xor1), .fa_or0(u_csamul_cla32_fa3_23_or0));
  and_gate and_gate_u_csamul_cla32_and4_23(.a(a[4]), .b(b[23]), .out(u_csamul_cla32_and4_23));
  fa fa_u_csamul_cla32_fa4_23_out(.a(u_csamul_cla32_and4_23[0]), .b(u_csamul_cla32_fa5_22_xor1[0]), .cin(u_csamul_cla32_fa4_22_or0[0]), .fa_xor1(u_csamul_cla32_fa4_23_xor1), .fa_or0(u_csamul_cla32_fa4_23_or0));
  and_gate and_gate_u_csamul_cla32_and5_23(.a(a[5]), .b(b[23]), .out(u_csamul_cla32_and5_23));
  fa fa_u_csamul_cla32_fa5_23_out(.a(u_csamul_cla32_and5_23[0]), .b(u_csamul_cla32_fa6_22_xor1[0]), .cin(u_csamul_cla32_fa5_22_or0[0]), .fa_xor1(u_csamul_cla32_fa5_23_xor1), .fa_or0(u_csamul_cla32_fa5_23_or0));
  and_gate and_gate_u_csamul_cla32_and6_23(.a(a[6]), .b(b[23]), .out(u_csamul_cla32_and6_23));
  fa fa_u_csamul_cla32_fa6_23_out(.a(u_csamul_cla32_and6_23[0]), .b(u_csamul_cla32_fa7_22_xor1[0]), .cin(u_csamul_cla32_fa6_22_or0[0]), .fa_xor1(u_csamul_cla32_fa6_23_xor1), .fa_or0(u_csamul_cla32_fa6_23_or0));
  and_gate and_gate_u_csamul_cla32_and7_23(.a(a[7]), .b(b[23]), .out(u_csamul_cla32_and7_23));
  fa fa_u_csamul_cla32_fa7_23_out(.a(u_csamul_cla32_and7_23[0]), .b(u_csamul_cla32_fa8_22_xor1[0]), .cin(u_csamul_cla32_fa7_22_or0[0]), .fa_xor1(u_csamul_cla32_fa7_23_xor1), .fa_or0(u_csamul_cla32_fa7_23_or0));
  and_gate and_gate_u_csamul_cla32_and8_23(.a(a[8]), .b(b[23]), .out(u_csamul_cla32_and8_23));
  fa fa_u_csamul_cla32_fa8_23_out(.a(u_csamul_cla32_and8_23[0]), .b(u_csamul_cla32_fa9_22_xor1[0]), .cin(u_csamul_cla32_fa8_22_or0[0]), .fa_xor1(u_csamul_cla32_fa8_23_xor1), .fa_or0(u_csamul_cla32_fa8_23_or0));
  and_gate and_gate_u_csamul_cla32_and9_23(.a(a[9]), .b(b[23]), .out(u_csamul_cla32_and9_23));
  fa fa_u_csamul_cla32_fa9_23_out(.a(u_csamul_cla32_and9_23[0]), .b(u_csamul_cla32_fa10_22_xor1[0]), .cin(u_csamul_cla32_fa9_22_or0[0]), .fa_xor1(u_csamul_cla32_fa9_23_xor1), .fa_or0(u_csamul_cla32_fa9_23_or0));
  and_gate and_gate_u_csamul_cla32_and10_23(.a(a[10]), .b(b[23]), .out(u_csamul_cla32_and10_23));
  fa fa_u_csamul_cla32_fa10_23_out(.a(u_csamul_cla32_and10_23[0]), .b(u_csamul_cla32_fa11_22_xor1[0]), .cin(u_csamul_cla32_fa10_22_or0[0]), .fa_xor1(u_csamul_cla32_fa10_23_xor1), .fa_or0(u_csamul_cla32_fa10_23_or0));
  and_gate and_gate_u_csamul_cla32_and11_23(.a(a[11]), .b(b[23]), .out(u_csamul_cla32_and11_23));
  fa fa_u_csamul_cla32_fa11_23_out(.a(u_csamul_cla32_and11_23[0]), .b(u_csamul_cla32_fa12_22_xor1[0]), .cin(u_csamul_cla32_fa11_22_or0[0]), .fa_xor1(u_csamul_cla32_fa11_23_xor1), .fa_or0(u_csamul_cla32_fa11_23_or0));
  and_gate and_gate_u_csamul_cla32_and12_23(.a(a[12]), .b(b[23]), .out(u_csamul_cla32_and12_23));
  fa fa_u_csamul_cla32_fa12_23_out(.a(u_csamul_cla32_and12_23[0]), .b(u_csamul_cla32_fa13_22_xor1[0]), .cin(u_csamul_cla32_fa12_22_or0[0]), .fa_xor1(u_csamul_cla32_fa12_23_xor1), .fa_or0(u_csamul_cla32_fa12_23_or0));
  and_gate and_gate_u_csamul_cla32_and13_23(.a(a[13]), .b(b[23]), .out(u_csamul_cla32_and13_23));
  fa fa_u_csamul_cla32_fa13_23_out(.a(u_csamul_cla32_and13_23[0]), .b(u_csamul_cla32_fa14_22_xor1[0]), .cin(u_csamul_cla32_fa13_22_or0[0]), .fa_xor1(u_csamul_cla32_fa13_23_xor1), .fa_or0(u_csamul_cla32_fa13_23_or0));
  and_gate and_gate_u_csamul_cla32_and14_23(.a(a[14]), .b(b[23]), .out(u_csamul_cla32_and14_23));
  fa fa_u_csamul_cla32_fa14_23_out(.a(u_csamul_cla32_and14_23[0]), .b(u_csamul_cla32_fa15_22_xor1[0]), .cin(u_csamul_cla32_fa14_22_or0[0]), .fa_xor1(u_csamul_cla32_fa14_23_xor1), .fa_or0(u_csamul_cla32_fa14_23_or0));
  and_gate and_gate_u_csamul_cla32_and15_23(.a(a[15]), .b(b[23]), .out(u_csamul_cla32_and15_23));
  fa fa_u_csamul_cla32_fa15_23_out(.a(u_csamul_cla32_and15_23[0]), .b(u_csamul_cla32_fa16_22_xor1[0]), .cin(u_csamul_cla32_fa15_22_or0[0]), .fa_xor1(u_csamul_cla32_fa15_23_xor1), .fa_or0(u_csamul_cla32_fa15_23_or0));
  and_gate and_gate_u_csamul_cla32_and16_23(.a(a[16]), .b(b[23]), .out(u_csamul_cla32_and16_23));
  fa fa_u_csamul_cla32_fa16_23_out(.a(u_csamul_cla32_and16_23[0]), .b(u_csamul_cla32_fa17_22_xor1[0]), .cin(u_csamul_cla32_fa16_22_or0[0]), .fa_xor1(u_csamul_cla32_fa16_23_xor1), .fa_or0(u_csamul_cla32_fa16_23_or0));
  and_gate and_gate_u_csamul_cla32_and17_23(.a(a[17]), .b(b[23]), .out(u_csamul_cla32_and17_23));
  fa fa_u_csamul_cla32_fa17_23_out(.a(u_csamul_cla32_and17_23[0]), .b(u_csamul_cla32_fa18_22_xor1[0]), .cin(u_csamul_cla32_fa17_22_or0[0]), .fa_xor1(u_csamul_cla32_fa17_23_xor1), .fa_or0(u_csamul_cla32_fa17_23_or0));
  and_gate and_gate_u_csamul_cla32_and18_23(.a(a[18]), .b(b[23]), .out(u_csamul_cla32_and18_23));
  fa fa_u_csamul_cla32_fa18_23_out(.a(u_csamul_cla32_and18_23[0]), .b(u_csamul_cla32_fa19_22_xor1[0]), .cin(u_csamul_cla32_fa18_22_or0[0]), .fa_xor1(u_csamul_cla32_fa18_23_xor1), .fa_or0(u_csamul_cla32_fa18_23_or0));
  and_gate and_gate_u_csamul_cla32_and19_23(.a(a[19]), .b(b[23]), .out(u_csamul_cla32_and19_23));
  fa fa_u_csamul_cla32_fa19_23_out(.a(u_csamul_cla32_and19_23[0]), .b(u_csamul_cla32_fa20_22_xor1[0]), .cin(u_csamul_cla32_fa19_22_or0[0]), .fa_xor1(u_csamul_cla32_fa19_23_xor1), .fa_or0(u_csamul_cla32_fa19_23_or0));
  and_gate and_gate_u_csamul_cla32_and20_23(.a(a[20]), .b(b[23]), .out(u_csamul_cla32_and20_23));
  fa fa_u_csamul_cla32_fa20_23_out(.a(u_csamul_cla32_and20_23[0]), .b(u_csamul_cla32_fa21_22_xor1[0]), .cin(u_csamul_cla32_fa20_22_or0[0]), .fa_xor1(u_csamul_cla32_fa20_23_xor1), .fa_or0(u_csamul_cla32_fa20_23_or0));
  and_gate and_gate_u_csamul_cla32_and21_23(.a(a[21]), .b(b[23]), .out(u_csamul_cla32_and21_23));
  fa fa_u_csamul_cla32_fa21_23_out(.a(u_csamul_cla32_and21_23[0]), .b(u_csamul_cla32_fa22_22_xor1[0]), .cin(u_csamul_cla32_fa21_22_or0[0]), .fa_xor1(u_csamul_cla32_fa21_23_xor1), .fa_or0(u_csamul_cla32_fa21_23_or0));
  and_gate and_gate_u_csamul_cla32_and22_23(.a(a[22]), .b(b[23]), .out(u_csamul_cla32_and22_23));
  fa fa_u_csamul_cla32_fa22_23_out(.a(u_csamul_cla32_and22_23[0]), .b(u_csamul_cla32_fa23_22_xor1[0]), .cin(u_csamul_cla32_fa22_22_or0[0]), .fa_xor1(u_csamul_cla32_fa22_23_xor1), .fa_or0(u_csamul_cla32_fa22_23_or0));
  and_gate and_gate_u_csamul_cla32_and23_23(.a(a[23]), .b(b[23]), .out(u_csamul_cla32_and23_23));
  fa fa_u_csamul_cla32_fa23_23_out(.a(u_csamul_cla32_and23_23[0]), .b(u_csamul_cla32_fa24_22_xor1[0]), .cin(u_csamul_cla32_fa23_22_or0[0]), .fa_xor1(u_csamul_cla32_fa23_23_xor1), .fa_or0(u_csamul_cla32_fa23_23_or0));
  and_gate and_gate_u_csamul_cla32_and24_23(.a(a[24]), .b(b[23]), .out(u_csamul_cla32_and24_23));
  fa fa_u_csamul_cla32_fa24_23_out(.a(u_csamul_cla32_and24_23[0]), .b(u_csamul_cla32_fa25_22_xor1[0]), .cin(u_csamul_cla32_fa24_22_or0[0]), .fa_xor1(u_csamul_cla32_fa24_23_xor1), .fa_or0(u_csamul_cla32_fa24_23_or0));
  and_gate and_gate_u_csamul_cla32_and25_23(.a(a[25]), .b(b[23]), .out(u_csamul_cla32_and25_23));
  fa fa_u_csamul_cla32_fa25_23_out(.a(u_csamul_cla32_and25_23[0]), .b(u_csamul_cla32_fa26_22_xor1[0]), .cin(u_csamul_cla32_fa25_22_or0[0]), .fa_xor1(u_csamul_cla32_fa25_23_xor1), .fa_or0(u_csamul_cla32_fa25_23_or0));
  and_gate and_gate_u_csamul_cla32_and26_23(.a(a[26]), .b(b[23]), .out(u_csamul_cla32_and26_23));
  fa fa_u_csamul_cla32_fa26_23_out(.a(u_csamul_cla32_and26_23[0]), .b(u_csamul_cla32_fa27_22_xor1[0]), .cin(u_csamul_cla32_fa26_22_or0[0]), .fa_xor1(u_csamul_cla32_fa26_23_xor1), .fa_or0(u_csamul_cla32_fa26_23_or0));
  and_gate and_gate_u_csamul_cla32_and27_23(.a(a[27]), .b(b[23]), .out(u_csamul_cla32_and27_23));
  fa fa_u_csamul_cla32_fa27_23_out(.a(u_csamul_cla32_and27_23[0]), .b(u_csamul_cla32_fa28_22_xor1[0]), .cin(u_csamul_cla32_fa27_22_or0[0]), .fa_xor1(u_csamul_cla32_fa27_23_xor1), .fa_or0(u_csamul_cla32_fa27_23_or0));
  and_gate and_gate_u_csamul_cla32_and28_23(.a(a[28]), .b(b[23]), .out(u_csamul_cla32_and28_23));
  fa fa_u_csamul_cla32_fa28_23_out(.a(u_csamul_cla32_and28_23[0]), .b(u_csamul_cla32_fa29_22_xor1[0]), .cin(u_csamul_cla32_fa28_22_or0[0]), .fa_xor1(u_csamul_cla32_fa28_23_xor1), .fa_or0(u_csamul_cla32_fa28_23_or0));
  and_gate and_gate_u_csamul_cla32_and29_23(.a(a[29]), .b(b[23]), .out(u_csamul_cla32_and29_23));
  fa fa_u_csamul_cla32_fa29_23_out(.a(u_csamul_cla32_and29_23[0]), .b(u_csamul_cla32_fa30_22_xor1[0]), .cin(u_csamul_cla32_fa29_22_or0[0]), .fa_xor1(u_csamul_cla32_fa29_23_xor1), .fa_or0(u_csamul_cla32_fa29_23_or0));
  and_gate and_gate_u_csamul_cla32_and30_23(.a(a[30]), .b(b[23]), .out(u_csamul_cla32_and30_23));
  fa fa_u_csamul_cla32_fa30_23_out(.a(u_csamul_cla32_and30_23[0]), .b(u_csamul_cla32_and31_22[0]), .cin(u_csamul_cla32_fa30_22_or0[0]), .fa_xor1(u_csamul_cla32_fa30_23_xor1), .fa_or0(u_csamul_cla32_fa30_23_or0));
  and_gate and_gate_u_csamul_cla32_and31_23(.a(a[31]), .b(b[23]), .out(u_csamul_cla32_and31_23));
  and_gate and_gate_u_csamul_cla32_and0_24(.a(a[0]), .b(b[24]), .out(u_csamul_cla32_and0_24));
  fa fa_u_csamul_cla32_fa0_24_out(.a(u_csamul_cla32_and0_24[0]), .b(u_csamul_cla32_fa1_23_xor1[0]), .cin(u_csamul_cla32_fa0_23_or0[0]), .fa_xor1(u_csamul_cla32_fa0_24_xor1), .fa_or0(u_csamul_cla32_fa0_24_or0));
  and_gate and_gate_u_csamul_cla32_and1_24(.a(a[1]), .b(b[24]), .out(u_csamul_cla32_and1_24));
  fa fa_u_csamul_cla32_fa1_24_out(.a(u_csamul_cla32_and1_24[0]), .b(u_csamul_cla32_fa2_23_xor1[0]), .cin(u_csamul_cla32_fa1_23_or0[0]), .fa_xor1(u_csamul_cla32_fa1_24_xor1), .fa_or0(u_csamul_cla32_fa1_24_or0));
  and_gate and_gate_u_csamul_cla32_and2_24(.a(a[2]), .b(b[24]), .out(u_csamul_cla32_and2_24));
  fa fa_u_csamul_cla32_fa2_24_out(.a(u_csamul_cla32_and2_24[0]), .b(u_csamul_cla32_fa3_23_xor1[0]), .cin(u_csamul_cla32_fa2_23_or0[0]), .fa_xor1(u_csamul_cla32_fa2_24_xor1), .fa_or0(u_csamul_cla32_fa2_24_or0));
  and_gate and_gate_u_csamul_cla32_and3_24(.a(a[3]), .b(b[24]), .out(u_csamul_cla32_and3_24));
  fa fa_u_csamul_cla32_fa3_24_out(.a(u_csamul_cla32_and3_24[0]), .b(u_csamul_cla32_fa4_23_xor1[0]), .cin(u_csamul_cla32_fa3_23_or0[0]), .fa_xor1(u_csamul_cla32_fa3_24_xor1), .fa_or0(u_csamul_cla32_fa3_24_or0));
  and_gate and_gate_u_csamul_cla32_and4_24(.a(a[4]), .b(b[24]), .out(u_csamul_cla32_and4_24));
  fa fa_u_csamul_cla32_fa4_24_out(.a(u_csamul_cla32_and4_24[0]), .b(u_csamul_cla32_fa5_23_xor1[0]), .cin(u_csamul_cla32_fa4_23_or0[0]), .fa_xor1(u_csamul_cla32_fa4_24_xor1), .fa_or0(u_csamul_cla32_fa4_24_or0));
  and_gate and_gate_u_csamul_cla32_and5_24(.a(a[5]), .b(b[24]), .out(u_csamul_cla32_and5_24));
  fa fa_u_csamul_cla32_fa5_24_out(.a(u_csamul_cla32_and5_24[0]), .b(u_csamul_cla32_fa6_23_xor1[0]), .cin(u_csamul_cla32_fa5_23_or0[0]), .fa_xor1(u_csamul_cla32_fa5_24_xor1), .fa_or0(u_csamul_cla32_fa5_24_or0));
  and_gate and_gate_u_csamul_cla32_and6_24(.a(a[6]), .b(b[24]), .out(u_csamul_cla32_and6_24));
  fa fa_u_csamul_cla32_fa6_24_out(.a(u_csamul_cla32_and6_24[0]), .b(u_csamul_cla32_fa7_23_xor1[0]), .cin(u_csamul_cla32_fa6_23_or0[0]), .fa_xor1(u_csamul_cla32_fa6_24_xor1), .fa_or0(u_csamul_cla32_fa6_24_or0));
  and_gate and_gate_u_csamul_cla32_and7_24(.a(a[7]), .b(b[24]), .out(u_csamul_cla32_and7_24));
  fa fa_u_csamul_cla32_fa7_24_out(.a(u_csamul_cla32_and7_24[0]), .b(u_csamul_cla32_fa8_23_xor1[0]), .cin(u_csamul_cla32_fa7_23_or0[0]), .fa_xor1(u_csamul_cla32_fa7_24_xor1), .fa_or0(u_csamul_cla32_fa7_24_or0));
  and_gate and_gate_u_csamul_cla32_and8_24(.a(a[8]), .b(b[24]), .out(u_csamul_cla32_and8_24));
  fa fa_u_csamul_cla32_fa8_24_out(.a(u_csamul_cla32_and8_24[0]), .b(u_csamul_cla32_fa9_23_xor1[0]), .cin(u_csamul_cla32_fa8_23_or0[0]), .fa_xor1(u_csamul_cla32_fa8_24_xor1), .fa_or0(u_csamul_cla32_fa8_24_or0));
  and_gate and_gate_u_csamul_cla32_and9_24(.a(a[9]), .b(b[24]), .out(u_csamul_cla32_and9_24));
  fa fa_u_csamul_cla32_fa9_24_out(.a(u_csamul_cla32_and9_24[0]), .b(u_csamul_cla32_fa10_23_xor1[0]), .cin(u_csamul_cla32_fa9_23_or0[0]), .fa_xor1(u_csamul_cla32_fa9_24_xor1), .fa_or0(u_csamul_cla32_fa9_24_or0));
  and_gate and_gate_u_csamul_cla32_and10_24(.a(a[10]), .b(b[24]), .out(u_csamul_cla32_and10_24));
  fa fa_u_csamul_cla32_fa10_24_out(.a(u_csamul_cla32_and10_24[0]), .b(u_csamul_cla32_fa11_23_xor1[0]), .cin(u_csamul_cla32_fa10_23_or0[0]), .fa_xor1(u_csamul_cla32_fa10_24_xor1), .fa_or0(u_csamul_cla32_fa10_24_or0));
  and_gate and_gate_u_csamul_cla32_and11_24(.a(a[11]), .b(b[24]), .out(u_csamul_cla32_and11_24));
  fa fa_u_csamul_cla32_fa11_24_out(.a(u_csamul_cla32_and11_24[0]), .b(u_csamul_cla32_fa12_23_xor1[0]), .cin(u_csamul_cla32_fa11_23_or0[0]), .fa_xor1(u_csamul_cla32_fa11_24_xor1), .fa_or0(u_csamul_cla32_fa11_24_or0));
  and_gate and_gate_u_csamul_cla32_and12_24(.a(a[12]), .b(b[24]), .out(u_csamul_cla32_and12_24));
  fa fa_u_csamul_cla32_fa12_24_out(.a(u_csamul_cla32_and12_24[0]), .b(u_csamul_cla32_fa13_23_xor1[0]), .cin(u_csamul_cla32_fa12_23_or0[0]), .fa_xor1(u_csamul_cla32_fa12_24_xor1), .fa_or0(u_csamul_cla32_fa12_24_or0));
  and_gate and_gate_u_csamul_cla32_and13_24(.a(a[13]), .b(b[24]), .out(u_csamul_cla32_and13_24));
  fa fa_u_csamul_cla32_fa13_24_out(.a(u_csamul_cla32_and13_24[0]), .b(u_csamul_cla32_fa14_23_xor1[0]), .cin(u_csamul_cla32_fa13_23_or0[0]), .fa_xor1(u_csamul_cla32_fa13_24_xor1), .fa_or0(u_csamul_cla32_fa13_24_or0));
  and_gate and_gate_u_csamul_cla32_and14_24(.a(a[14]), .b(b[24]), .out(u_csamul_cla32_and14_24));
  fa fa_u_csamul_cla32_fa14_24_out(.a(u_csamul_cla32_and14_24[0]), .b(u_csamul_cla32_fa15_23_xor1[0]), .cin(u_csamul_cla32_fa14_23_or0[0]), .fa_xor1(u_csamul_cla32_fa14_24_xor1), .fa_or0(u_csamul_cla32_fa14_24_or0));
  and_gate and_gate_u_csamul_cla32_and15_24(.a(a[15]), .b(b[24]), .out(u_csamul_cla32_and15_24));
  fa fa_u_csamul_cla32_fa15_24_out(.a(u_csamul_cla32_and15_24[0]), .b(u_csamul_cla32_fa16_23_xor1[0]), .cin(u_csamul_cla32_fa15_23_or0[0]), .fa_xor1(u_csamul_cla32_fa15_24_xor1), .fa_or0(u_csamul_cla32_fa15_24_or0));
  and_gate and_gate_u_csamul_cla32_and16_24(.a(a[16]), .b(b[24]), .out(u_csamul_cla32_and16_24));
  fa fa_u_csamul_cla32_fa16_24_out(.a(u_csamul_cla32_and16_24[0]), .b(u_csamul_cla32_fa17_23_xor1[0]), .cin(u_csamul_cla32_fa16_23_or0[0]), .fa_xor1(u_csamul_cla32_fa16_24_xor1), .fa_or0(u_csamul_cla32_fa16_24_or0));
  and_gate and_gate_u_csamul_cla32_and17_24(.a(a[17]), .b(b[24]), .out(u_csamul_cla32_and17_24));
  fa fa_u_csamul_cla32_fa17_24_out(.a(u_csamul_cla32_and17_24[0]), .b(u_csamul_cla32_fa18_23_xor1[0]), .cin(u_csamul_cla32_fa17_23_or0[0]), .fa_xor1(u_csamul_cla32_fa17_24_xor1), .fa_or0(u_csamul_cla32_fa17_24_or0));
  and_gate and_gate_u_csamul_cla32_and18_24(.a(a[18]), .b(b[24]), .out(u_csamul_cla32_and18_24));
  fa fa_u_csamul_cla32_fa18_24_out(.a(u_csamul_cla32_and18_24[0]), .b(u_csamul_cla32_fa19_23_xor1[0]), .cin(u_csamul_cla32_fa18_23_or0[0]), .fa_xor1(u_csamul_cla32_fa18_24_xor1), .fa_or0(u_csamul_cla32_fa18_24_or0));
  and_gate and_gate_u_csamul_cla32_and19_24(.a(a[19]), .b(b[24]), .out(u_csamul_cla32_and19_24));
  fa fa_u_csamul_cla32_fa19_24_out(.a(u_csamul_cla32_and19_24[0]), .b(u_csamul_cla32_fa20_23_xor1[0]), .cin(u_csamul_cla32_fa19_23_or0[0]), .fa_xor1(u_csamul_cla32_fa19_24_xor1), .fa_or0(u_csamul_cla32_fa19_24_or0));
  and_gate and_gate_u_csamul_cla32_and20_24(.a(a[20]), .b(b[24]), .out(u_csamul_cla32_and20_24));
  fa fa_u_csamul_cla32_fa20_24_out(.a(u_csamul_cla32_and20_24[0]), .b(u_csamul_cla32_fa21_23_xor1[0]), .cin(u_csamul_cla32_fa20_23_or0[0]), .fa_xor1(u_csamul_cla32_fa20_24_xor1), .fa_or0(u_csamul_cla32_fa20_24_or0));
  and_gate and_gate_u_csamul_cla32_and21_24(.a(a[21]), .b(b[24]), .out(u_csamul_cla32_and21_24));
  fa fa_u_csamul_cla32_fa21_24_out(.a(u_csamul_cla32_and21_24[0]), .b(u_csamul_cla32_fa22_23_xor1[0]), .cin(u_csamul_cla32_fa21_23_or0[0]), .fa_xor1(u_csamul_cla32_fa21_24_xor1), .fa_or0(u_csamul_cla32_fa21_24_or0));
  and_gate and_gate_u_csamul_cla32_and22_24(.a(a[22]), .b(b[24]), .out(u_csamul_cla32_and22_24));
  fa fa_u_csamul_cla32_fa22_24_out(.a(u_csamul_cla32_and22_24[0]), .b(u_csamul_cla32_fa23_23_xor1[0]), .cin(u_csamul_cla32_fa22_23_or0[0]), .fa_xor1(u_csamul_cla32_fa22_24_xor1), .fa_or0(u_csamul_cla32_fa22_24_or0));
  and_gate and_gate_u_csamul_cla32_and23_24(.a(a[23]), .b(b[24]), .out(u_csamul_cla32_and23_24));
  fa fa_u_csamul_cla32_fa23_24_out(.a(u_csamul_cla32_and23_24[0]), .b(u_csamul_cla32_fa24_23_xor1[0]), .cin(u_csamul_cla32_fa23_23_or0[0]), .fa_xor1(u_csamul_cla32_fa23_24_xor1), .fa_or0(u_csamul_cla32_fa23_24_or0));
  and_gate and_gate_u_csamul_cla32_and24_24(.a(a[24]), .b(b[24]), .out(u_csamul_cla32_and24_24));
  fa fa_u_csamul_cla32_fa24_24_out(.a(u_csamul_cla32_and24_24[0]), .b(u_csamul_cla32_fa25_23_xor1[0]), .cin(u_csamul_cla32_fa24_23_or0[0]), .fa_xor1(u_csamul_cla32_fa24_24_xor1), .fa_or0(u_csamul_cla32_fa24_24_or0));
  and_gate and_gate_u_csamul_cla32_and25_24(.a(a[25]), .b(b[24]), .out(u_csamul_cla32_and25_24));
  fa fa_u_csamul_cla32_fa25_24_out(.a(u_csamul_cla32_and25_24[0]), .b(u_csamul_cla32_fa26_23_xor1[0]), .cin(u_csamul_cla32_fa25_23_or0[0]), .fa_xor1(u_csamul_cla32_fa25_24_xor1), .fa_or0(u_csamul_cla32_fa25_24_or0));
  and_gate and_gate_u_csamul_cla32_and26_24(.a(a[26]), .b(b[24]), .out(u_csamul_cla32_and26_24));
  fa fa_u_csamul_cla32_fa26_24_out(.a(u_csamul_cla32_and26_24[0]), .b(u_csamul_cla32_fa27_23_xor1[0]), .cin(u_csamul_cla32_fa26_23_or0[0]), .fa_xor1(u_csamul_cla32_fa26_24_xor1), .fa_or0(u_csamul_cla32_fa26_24_or0));
  and_gate and_gate_u_csamul_cla32_and27_24(.a(a[27]), .b(b[24]), .out(u_csamul_cla32_and27_24));
  fa fa_u_csamul_cla32_fa27_24_out(.a(u_csamul_cla32_and27_24[0]), .b(u_csamul_cla32_fa28_23_xor1[0]), .cin(u_csamul_cla32_fa27_23_or0[0]), .fa_xor1(u_csamul_cla32_fa27_24_xor1), .fa_or0(u_csamul_cla32_fa27_24_or0));
  and_gate and_gate_u_csamul_cla32_and28_24(.a(a[28]), .b(b[24]), .out(u_csamul_cla32_and28_24));
  fa fa_u_csamul_cla32_fa28_24_out(.a(u_csamul_cla32_and28_24[0]), .b(u_csamul_cla32_fa29_23_xor1[0]), .cin(u_csamul_cla32_fa28_23_or0[0]), .fa_xor1(u_csamul_cla32_fa28_24_xor1), .fa_or0(u_csamul_cla32_fa28_24_or0));
  and_gate and_gate_u_csamul_cla32_and29_24(.a(a[29]), .b(b[24]), .out(u_csamul_cla32_and29_24));
  fa fa_u_csamul_cla32_fa29_24_out(.a(u_csamul_cla32_and29_24[0]), .b(u_csamul_cla32_fa30_23_xor1[0]), .cin(u_csamul_cla32_fa29_23_or0[0]), .fa_xor1(u_csamul_cla32_fa29_24_xor1), .fa_or0(u_csamul_cla32_fa29_24_or0));
  and_gate and_gate_u_csamul_cla32_and30_24(.a(a[30]), .b(b[24]), .out(u_csamul_cla32_and30_24));
  fa fa_u_csamul_cla32_fa30_24_out(.a(u_csamul_cla32_and30_24[0]), .b(u_csamul_cla32_and31_23[0]), .cin(u_csamul_cla32_fa30_23_or0[0]), .fa_xor1(u_csamul_cla32_fa30_24_xor1), .fa_or0(u_csamul_cla32_fa30_24_or0));
  and_gate and_gate_u_csamul_cla32_and31_24(.a(a[31]), .b(b[24]), .out(u_csamul_cla32_and31_24));
  and_gate and_gate_u_csamul_cla32_and0_25(.a(a[0]), .b(b[25]), .out(u_csamul_cla32_and0_25));
  fa fa_u_csamul_cla32_fa0_25_out(.a(u_csamul_cla32_and0_25[0]), .b(u_csamul_cla32_fa1_24_xor1[0]), .cin(u_csamul_cla32_fa0_24_or0[0]), .fa_xor1(u_csamul_cla32_fa0_25_xor1), .fa_or0(u_csamul_cla32_fa0_25_or0));
  and_gate and_gate_u_csamul_cla32_and1_25(.a(a[1]), .b(b[25]), .out(u_csamul_cla32_and1_25));
  fa fa_u_csamul_cla32_fa1_25_out(.a(u_csamul_cla32_and1_25[0]), .b(u_csamul_cla32_fa2_24_xor1[0]), .cin(u_csamul_cla32_fa1_24_or0[0]), .fa_xor1(u_csamul_cla32_fa1_25_xor1), .fa_or0(u_csamul_cla32_fa1_25_or0));
  and_gate and_gate_u_csamul_cla32_and2_25(.a(a[2]), .b(b[25]), .out(u_csamul_cla32_and2_25));
  fa fa_u_csamul_cla32_fa2_25_out(.a(u_csamul_cla32_and2_25[0]), .b(u_csamul_cla32_fa3_24_xor1[0]), .cin(u_csamul_cla32_fa2_24_or0[0]), .fa_xor1(u_csamul_cla32_fa2_25_xor1), .fa_or0(u_csamul_cla32_fa2_25_or0));
  and_gate and_gate_u_csamul_cla32_and3_25(.a(a[3]), .b(b[25]), .out(u_csamul_cla32_and3_25));
  fa fa_u_csamul_cla32_fa3_25_out(.a(u_csamul_cla32_and3_25[0]), .b(u_csamul_cla32_fa4_24_xor1[0]), .cin(u_csamul_cla32_fa3_24_or0[0]), .fa_xor1(u_csamul_cla32_fa3_25_xor1), .fa_or0(u_csamul_cla32_fa3_25_or0));
  and_gate and_gate_u_csamul_cla32_and4_25(.a(a[4]), .b(b[25]), .out(u_csamul_cla32_and4_25));
  fa fa_u_csamul_cla32_fa4_25_out(.a(u_csamul_cla32_and4_25[0]), .b(u_csamul_cla32_fa5_24_xor1[0]), .cin(u_csamul_cla32_fa4_24_or0[0]), .fa_xor1(u_csamul_cla32_fa4_25_xor1), .fa_or0(u_csamul_cla32_fa4_25_or0));
  and_gate and_gate_u_csamul_cla32_and5_25(.a(a[5]), .b(b[25]), .out(u_csamul_cla32_and5_25));
  fa fa_u_csamul_cla32_fa5_25_out(.a(u_csamul_cla32_and5_25[0]), .b(u_csamul_cla32_fa6_24_xor1[0]), .cin(u_csamul_cla32_fa5_24_or0[0]), .fa_xor1(u_csamul_cla32_fa5_25_xor1), .fa_or0(u_csamul_cla32_fa5_25_or0));
  and_gate and_gate_u_csamul_cla32_and6_25(.a(a[6]), .b(b[25]), .out(u_csamul_cla32_and6_25));
  fa fa_u_csamul_cla32_fa6_25_out(.a(u_csamul_cla32_and6_25[0]), .b(u_csamul_cla32_fa7_24_xor1[0]), .cin(u_csamul_cla32_fa6_24_or0[0]), .fa_xor1(u_csamul_cla32_fa6_25_xor1), .fa_or0(u_csamul_cla32_fa6_25_or0));
  and_gate and_gate_u_csamul_cla32_and7_25(.a(a[7]), .b(b[25]), .out(u_csamul_cla32_and7_25));
  fa fa_u_csamul_cla32_fa7_25_out(.a(u_csamul_cla32_and7_25[0]), .b(u_csamul_cla32_fa8_24_xor1[0]), .cin(u_csamul_cla32_fa7_24_or0[0]), .fa_xor1(u_csamul_cla32_fa7_25_xor1), .fa_or0(u_csamul_cla32_fa7_25_or0));
  and_gate and_gate_u_csamul_cla32_and8_25(.a(a[8]), .b(b[25]), .out(u_csamul_cla32_and8_25));
  fa fa_u_csamul_cla32_fa8_25_out(.a(u_csamul_cla32_and8_25[0]), .b(u_csamul_cla32_fa9_24_xor1[0]), .cin(u_csamul_cla32_fa8_24_or0[0]), .fa_xor1(u_csamul_cla32_fa8_25_xor1), .fa_or0(u_csamul_cla32_fa8_25_or0));
  and_gate and_gate_u_csamul_cla32_and9_25(.a(a[9]), .b(b[25]), .out(u_csamul_cla32_and9_25));
  fa fa_u_csamul_cla32_fa9_25_out(.a(u_csamul_cla32_and9_25[0]), .b(u_csamul_cla32_fa10_24_xor1[0]), .cin(u_csamul_cla32_fa9_24_or0[0]), .fa_xor1(u_csamul_cla32_fa9_25_xor1), .fa_or0(u_csamul_cla32_fa9_25_or0));
  and_gate and_gate_u_csamul_cla32_and10_25(.a(a[10]), .b(b[25]), .out(u_csamul_cla32_and10_25));
  fa fa_u_csamul_cla32_fa10_25_out(.a(u_csamul_cla32_and10_25[0]), .b(u_csamul_cla32_fa11_24_xor1[0]), .cin(u_csamul_cla32_fa10_24_or0[0]), .fa_xor1(u_csamul_cla32_fa10_25_xor1), .fa_or0(u_csamul_cla32_fa10_25_or0));
  and_gate and_gate_u_csamul_cla32_and11_25(.a(a[11]), .b(b[25]), .out(u_csamul_cla32_and11_25));
  fa fa_u_csamul_cla32_fa11_25_out(.a(u_csamul_cla32_and11_25[0]), .b(u_csamul_cla32_fa12_24_xor1[0]), .cin(u_csamul_cla32_fa11_24_or0[0]), .fa_xor1(u_csamul_cla32_fa11_25_xor1), .fa_or0(u_csamul_cla32_fa11_25_or0));
  and_gate and_gate_u_csamul_cla32_and12_25(.a(a[12]), .b(b[25]), .out(u_csamul_cla32_and12_25));
  fa fa_u_csamul_cla32_fa12_25_out(.a(u_csamul_cla32_and12_25[0]), .b(u_csamul_cla32_fa13_24_xor1[0]), .cin(u_csamul_cla32_fa12_24_or0[0]), .fa_xor1(u_csamul_cla32_fa12_25_xor1), .fa_or0(u_csamul_cla32_fa12_25_or0));
  and_gate and_gate_u_csamul_cla32_and13_25(.a(a[13]), .b(b[25]), .out(u_csamul_cla32_and13_25));
  fa fa_u_csamul_cla32_fa13_25_out(.a(u_csamul_cla32_and13_25[0]), .b(u_csamul_cla32_fa14_24_xor1[0]), .cin(u_csamul_cla32_fa13_24_or0[0]), .fa_xor1(u_csamul_cla32_fa13_25_xor1), .fa_or0(u_csamul_cla32_fa13_25_or0));
  and_gate and_gate_u_csamul_cla32_and14_25(.a(a[14]), .b(b[25]), .out(u_csamul_cla32_and14_25));
  fa fa_u_csamul_cla32_fa14_25_out(.a(u_csamul_cla32_and14_25[0]), .b(u_csamul_cla32_fa15_24_xor1[0]), .cin(u_csamul_cla32_fa14_24_or0[0]), .fa_xor1(u_csamul_cla32_fa14_25_xor1), .fa_or0(u_csamul_cla32_fa14_25_or0));
  and_gate and_gate_u_csamul_cla32_and15_25(.a(a[15]), .b(b[25]), .out(u_csamul_cla32_and15_25));
  fa fa_u_csamul_cla32_fa15_25_out(.a(u_csamul_cla32_and15_25[0]), .b(u_csamul_cla32_fa16_24_xor1[0]), .cin(u_csamul_cla32_fa15_24_or0[0]), .fa_xor1(u_csamul_cla32_fa15_25_xor1), .fa_or0(u_csamul_cla32_fa15_25_or0));
  and_gate and_gate_u_csamul_cla32_and16_25(.a(a[16]), .b(b[25]), .out(u_csamul_cla32_and16_25));
  fa fa_u_csamul_cla32_fa16_25_out(.a(u_csamul_cla32_and16_25[0]), .b(u_csamul_cla32_fa17_24_xor1[0]), .cin(u_csamul_cla32_fa16_24_or0[0]), .fa_xor1(u_csamul_cla32_fa16_25_xor1), .fa_or0(u_csamul_cla32_fa16_25_or0));
  and_gate and_gate_u_csamul_cla32_and17_25(.a(a[17]), .b(b[25]), .out(u_csamul_cla32_and17_25));
  fa fa_u_csamul_cla32_fa17_25_out(.a(u_csamul_cla32_and17_25[0]), .b(u_csamul_cla32_fa18_24_xor1[0]), .cin(u_csamul_cla32_fa17_24_or0[0]), .fa_xor1(u_csamul_cla32_fa17_25_xor1), .fa_or0(u_csamul_cla32_fa17_25_or0));
  and_gate and_gate_u_csamul_cla32_and18_25(.a(a[18]), .b(b[25]), .out(u_csamul_cla32_and18_25));
  fa fa_u_csamul_cla32_fa18_25_out(.a(u_csamul_cla32_and18_25[0]), .b(u_csamul_cla32_fa19_24_xor1[0]), .cin(u_csamul_cla32_fa18_24_or0[0]), .fa_xor1(u_csamul_cla32_fa18_25_xor1), .fa_or0(u_csamul_cla32_fa18_25_or0));
  and_gate and_gate_u_csamul_cla32_and19_25(.a(a[19]), .b(b[25]), .out(u_csamul_cla32_and19_25));
  fa fa_u_csamul_cla32_fa19_25_out(.a(u_csamul_cla32_and19_25[0]), .b(u_csamul_cla32_fa20_24_xor1[0]), .cin(u_csamul_cla32_fa19_24_or0[0]), .fa_xor1(u_csamul_cla32_fa19_25_xor1), .fa_or0(u_csamul_cla32_fa19_25_or0));
  and_gate and_gate_u_csamul_cla32_and20_25(.a(a[20]), .b(b[25]), .out(u_csamul_cla32_and20_25));
  fa fa_u_csamul_cla32_fa20_25_out(.a(u_csamul_cla32_and20_25[0]), .b(u_csamul_cla32_fa21_24_xor1[0]), .cin(u_csamul_cla32_fa20_24_or0[0]), .fa_xor1(u_csamul_cla32_fa20_25_xor1), .fa_or0(u_csamul_cla32_fa20_25_or0));
  and_gate and_gate_u_csamul_cla32_and21_25(.a(a[21]), .b(b[25]), .out(u_csamul_cla32_and21_25));
  fa fa_u_csamul_cla32_fa21_25_out(.a(u_csamul_cla32_and21_25[0]), .b(u_csamul_cla32_fa22_24_xor1[0]), .cin(u_csamul_cla32_fa21_24_or0[0]), .fa_xor1(u_csamul_cla32_fa21_25_xor1), .fa_or0(u_csamul_cla32_fa21_25_or0));
  and_gate and_gate_u_csamul_cla32_and22_25(.a(a[22]), .b(b[25]), .out(u_csamul_cla32_and22_25));
  fa fa_u_csamul_cla32_fa22_25_out(.a(u_csamul_cla32_and22_25[0]), .b(u_csamul_cla32_fa23_24_xor1[0]), .cin(u_csamul_cla32_fa22_24_or0[0]), .fa_xor1(u_csamul_cla32_fa22_25_xor1), .fa_or0(u_csamul_cla32_fa22_25_or0));
  and_gate and_gate_u_csamul_cla32_and23_25(.a(a[23]), .b(b[25]), .out(u_csamul_cla32_and23_25));
  fa fa_u_csamul_cla32_fa23_25_out(.a(u_csamul_cla32_and23_25[0]), .b(u_csamul_cla32_fa24_24_xor1[0]), .cin(u_csamul_cla32_fa23_24_or0[0]), .fa_xor1(u_csamul_cla32_fa23_25_xor1), .fa_or0(u_csamul_cla32_fa23_25_or0));
  and_gate and_gate_u_csamul_cla32_and24_25(.a(a[24]), .b(b[25]), .out(u_csamul_cla32_and24_25));
  fa fa_u_csamul_cla32_fa24_25_out(.a(u_csamul_cla32_and24_25[0]), .b(u_csamul_cla32_fa25_24_xor1[0]), .cin(u_csamul_cla32_fa24_24_or0[0]), .fa_xor1(u_csamul_cla32_fa24_25_xor1), .fa_or0(u_csamul_cla32_fa24_25_or0));
  and_gate and_gate_u_csamul_cla32_and25_25(.a(a[25]), .b(b[25]), .out(u_csamul_cla32_and25_25));
  fa fa_u_csamul_cla32_fa25_25_out(.a(u_csamul_cla32_and25_25[0]), .b(u_csamul_cla32_fa26_24_xor1[0]), .cin(u_csamul_cla32_fa25_24_or0[0]), .fa_xor1(u_csamul_cla32_fa25_25_xor1), .fa_or0(u_csamul_cla32_fa25_25_or0));
  and_gate and_gate_u_csamul_cla32_and26_25(.a(a[26]), .b(b[25]), .out(u_csamul_cla32_and26_25));
  fa fa_u_csamul_cla32_fa26_25_out(.a(u_csamul_cla32_and26_25[0]), .b(u_csamul_cla32_fa27_24_xor1[0]), .cin(u_csamul_cla32_fa26_24_or0[0]), .fa_xor1(u_csamul_cla32_fa26_25_xor1), .fa_or0(u_csamul_cla32_fa26_25_or0));
  and_gate and_gate_u_csamul_cla32_and27_25(.a(a[27]), .b(b[25]), .out(u_csamul_cla32_and27_25));
  fa fa_u_csamul_cla32_fa27_25_out(.a(u_csamul_cla32_and27_25[0]), .b(u_csamul_cla32_fa28_24_xor1[0]), .cin(u_csamul_cla32_fa27_24_or0[0]), .fa_xor1(u_csamul_cla32_fa27_25_xor1), .fa_or0(u_csamul_cla32_fa27_25_or0));
  and_gate and_gate_u_csamul_cla32_and28_25(.a(a[28]), .b(b[25]), .out(u_csamul_cla32_and28_25));
  fa fa_u_csamul_cla32_fa28_25_out(.a(u_csamul_cla32_and28_25[0]), .b(u_csamul_cla32_fa29_24_xor1[0]), .cin(u_csamul_cla32_fa28_24_or0[0]), .fa_xor1(u_csamul_cla32_fa28_25_xor1), .fa_or0(u_csamul_cla32_fa28_25_or0));
  and_gate and_gate_u_csamul_cla32_and29_25(.a(a[29]), .b(b[25]), .out(u_csamul_cla32_and29_25));
  fa fa_u_csamul_cla32_fa29_25_out(.a(u_csamul_cla32_and29_25[0]), .b(u_csamul_cla32_fa30_24_xor1[0]), .cin(u_csamul_cla32_fa29_24_or0[0]), .fa_xor1(u_csamul_cla32_fa29_25_xor1), .fa_or0(u_csamul_cla32_fa29_25_or0));
  and_gate and_gate_u_csamul_cla32_and30_25(.a(a[30]), .b(b[25]), .out(u_csamul_cla32_and30_25));
  fa fa_u_csamul_cla32_fa30_25_out(.a(u_csamul_cla32_and30_25[0]), .b(u_csamul_cla32_and31_24[0]), .cin(u_csamul_cla32_fa30_24_or0[0]), .fa_xor1(u_csamul_cla32_fa30_25_xor1), .fa_or0(u_csamul_cla32_fa30_25_or0));
  and_gate and_gate_u_csamul_cla32_and31_25(.a(a[31]), .b(b[25]), .out(u_csamul_cla32_and31_25));
  and_gate and_gate_u_csamul_cla32_and0_26(.a(a[0]), .b(b[26]), .out(u_csamul_cla32_and0_26));
  fa fa_u_csamul_cla32_fa0_26_out(.a(u_csamul_cla32_and0_26[0]), .b(u_csamul_cla32_fa1_25_xor1[0]), .cin(u_csamul_cla32_fa0_25_or0[0]), .fa_xor1(u_csamul_cla32_fa0_26_xor1), .fa_or0(u_csamul_cla32_fa0_26_or0));
  and_gate and_gate_u_csamul_cla32_and1_26(.a(a[1]), .b(b[26]), .out(u_csamul_cla32_and1_26));
  fa fa_u_csamul_cla32_fa1_26_out(.a(u_csamul_cla32_and1_26[0]), .b(u_csamul_cla32_fa2_25_xor1[0]), .cin(u_csamul_cla32_fa1_25_or0[0]), .fa_xor1(u_csamul_cla32_fa1_26_xor1), .fa_or0(u_csamul_cla32_fa1_26_or0));
  and_gate and_gate_u_csamul_cla32_and2_26(.a(a[2]), .b(b[26]), .out(u_csamul_cla32_and2_26));
  fa fa_u_csamul_cla32_fa2_26_out(.a(u_csamul_cla32_and2_26[0]), .b(u_csamul_cla32_fa3_25_xor1[0]), .cin(u_csamul_cla32_fa2_25_or0[0]), .fa_xor1(u_csamul_cla32_fa2_26_xor1), .fa_or0(u_csamul_cla32_fa2_26_or0));
  and_gate and_gate_u_csamul_cla32_and3_26(.a(a[3]), .b(b[26]), .out(u_csamul_cla32_and3_26));
  fa fa_u_csamul_cla32_fa3_26_out(.a(u_csamul_cla32_and3_26[0]), .b(u_csamul_cla32_fa4_25_xor1[0]), .cin(u_csamul_cla32_fa3_25_or0[0]), .fa_xor1(u_csamul_cla32_fa3_26_xor1), .fa_or0(u_csamul_cla32_fa3_26_or0));
  and_gate and_gate_u_csamul_cla32_and4_26(.a(a[4]), .b(b[26]), .out(u_csamul_cla32_and4_26));
  fa fa_u_csamul_cla32_fa4_26_out(.a(u_csamul_cla32_and4_26[0]), .b(u_csamul_cla32_fa5_25_xor1[0]), .cin(u_csamul_cla32_fa4_25_or0[0]), .fa_xor1(u_csamul_cla32_fa4_26_xor1), .fa_or0(u_csamul_cla32_fa4_26_or0));
  and_gate and_gate_u_csamul_cla32_and5_26(.a(a[5]), .b(b[26]), .out(u_csamul_cla32_and5_26));
  fa fa_u_csamul_cla32_fa5_26_out(.a(u_csamul_cla32_and5_26[0]), .b(u_csamul_cla32_fa6_25_xor1[0]), .cin(u_csamul_cla32_fa5_25_or0[0]), .fa_xor1(u_csamul_cla32_fa5_26_xor1), .fa_or0(u_csamul_cla32_fa5_26_or0));
  and_gate and_gate_u_csamul_cla32_and6_26(.a(a[6]), .b(b[26]), .out(u_csamul_cla32_and6_26));
  fa fa_u_csamul_cla32_fa6_26_out(.a(u_csamul_cla32_and6_26[0]), .b(u_csamul_cla32_fa7_25_xor1[0]), .cin(u_csamul_cla32_fa6_25_or0[0]), .fa_xor1(u_csamul_cla32_fa6_26_xor1), .fa_or0(u_csamul_cla32_fa6_26_or0));
  and_gate and_gate_u_csamul_cla32_and7_26(.a(a[7]), .b(b[26]), .out(u_csamul_cla32_and7_26));
  fa fa_u_csamul_cla32_fa7_26_out(.a(u_csamul_cla32_and7_26[0]), .b(u_csamul_cla32_fa8_25_xor1[0]), .cin(u_csamul_cla32_fa7_25_or0[0]), .fa_xor1(u_csamul_cla32_fa7_26_xor1), .fa_or0(u_csamul_cla32_fa7_26_or0));
  and_gate and_gate_u_csamul_cla32_and8_26(.a(a[8]), .b(b[26]), .out(u_csamul_cla32_and8_26));
  fa fa_u_csamul_cla32_fa8_26_out(.a(u_csamul_cla32_and8_26[0]), .b(u_csamul_cla32_fa9_25_xor1[0]), .cin(u_csamul_cla32_fa8_25_or0[0]), .fa_xor1(u_csamul_cla32_fa8_26_xor1), .fa_or0(u_csamul_cla32_fa8_26_or0));
  and_gate and_gate_u_csamul_cla32_and9_26(.a(a[9]), .b(b[26]), .out(u_csamul_cla32_and9_26));
  fa fa_u_csamul_cla32_fa9_26_out(.a(u_csamul_cla32_and9_26[0]), .b(u_csamul_cla32_fa10_25_xor1[0]), .cin(u_csamul_cla32_fa9_25_or0[0]), .fa_xor1(u_csamul_cla32_fa9_26_xor1), .fa_or0(u_csamul_cla32_fa9_26_or0));
  and_gate and_gate_u_csamul_cla32_and10_26(.a(a[10]), .b(b[26]), .out(u_csamul_cla32_and10_26));
  fa fa_u_csamul_cla32_fa10_26_out(.a(u_csamul_cla32_and10_26[0]), .b(u_csamul_cla32_fa11_25_xor1[0]), .cin(u_csamul_cla32_fa10_25_or0[0]), .fa_xor1(u_csamul_cla32_fa10_26_xor1), .fa_or0(u_csamul_cla32_fa10_26_or0));
  and_gate and_gate_u_csamul_cla32_and11_26(.a(a[11]), .b(b[26]), .out(u_csamul_cla32_and11_26));
  fa fa_u_csamul_cla32_fa11_26_out(.a(u_csamul_cla32_and11_26[0]), .b(u_csamul_cla32_fa12_25_xor1[0]), .cin(u_csamul_cla32_fa11_25_or0[0]), .fa_xor1(u_csamul_cla32_fa11_26_xor1), .fa_or0(u_csamul_cla32_fa11_26_or0));
  and_gate and_gate_u_csamul_cla32_and12_26(.a(a[12]), .b(b[26]), .out(u_csamul_cla32_and12_26));
  fa fa_u_csamul_cla32_fa12_26_out(.a(u_csamul_cla32_and12_26[0]), .b(u_csamul_cla32_fa13_25_xor1[0]), .cin(u_csamul_cla32_fa12_25_or0[0]), .fa_xor1(u_csamul_cla32_fa12_26_xor1), .fa_or0(u_csamul_cla32_fa12_26_or0));
  and_gate and_gate_u_csamul_cla32_and13_26(.a(a[13]), .b(b[26]), .out(u_csamul_cla32_and13_26));
  fa fa_u_csamul_cla32_fa13_26_out(.a(u_csamul_cla32_and13_26[0]), .b(u_csamul_cla32_fa14_25_xor1[0]), .cin(u_csamul_cla32_fa13_25_or0[0]), .fa_xor1(u_csamul_cla32_fa13_26_xor1), .fa_or0(u_csamul_cla32_fa13_26_or0));
  and_gate and_gate_u_csamul_cla32_and14_26(.a(a[14]), .b(b[26]), .out(u_csamul_cla32_and14_26));
  fa fa_u_csamul_cla32_fa14_26_out(.a(u_csamul_cla32_and14_26[0]), .b(u_csamul_cla32_fa15_25_xor1[0]), .cin(u_csamul_cla32_fa14_25_or0[0]), .fa_xor1(u_csamul_cla32_fa14_26_xor1), .fa_or0(u_csamul_cla32_fa14_26_or0));
  and_gate and_gate_u_csamul_cla32_and15_26(.a(a[15]), .b(b[26]), .out(u_csamul_cla32_and15_26));
  fa fa_u_csamul_cla32_fa15_26_out(.a(u_csamul_cla32_and15_26[0]), .b(u_csamul_cla32_fa16_25_xor1[0]), .cin(u_csamul_cla32_fa15_25_or0[0]), .fa_xor1(u_csamul_cla32_fa15_26_xor1), .fa_or0(u_csamul_cla32_fa15_26_or0));
  and_gate and_gate_u_csamul_cla32_and16_26(.a(a[16]), .b(b[26]), .out(u_csamul_cla32_and16_26));
  fa fa_u_csamul_cla32_fa16_26_out(.a(u_csamul_cla32_and16_26[0]), .b(u_csamul_cla32_fa17_25_xor1[0]), .cin(u_csamul_cla32_fa16_25_or0[0]), .fa_xor1(u_csamul_cla32_fa16_26_xor1), .fa_or0(u_csamul_cla32_fa16_26_or0));
  and_gate and_gate_u_csamul_cla32_and17_26(.a(a[17]), .b(b[26]), .out(u_csamul_cla32_and17_26));
  fa fa_u_csamul_cla32_fa17_26_out(.a(u_csamul_cla32_and17_26[0]), .b(u_csamul_cla32_fa18_25_xor1[0]), .cin(u_csamul_cla32_fa17_25_or0[0]), .fa_xor1(u_csamul_cla32_fa17_26_xor1), .fa_or0(u_csamul_cla32_fa17_26_or0));
  and_gate and_gate_u_csamul_cla32_and18_26(.a(a[18]), .b(b[26]), .out(u_csamul_cla32_and18_26));
  fa fa_u_csamul_cla32_fa18_26_out(.a(u_csamul_cla32_and18_26[0]), .b(u_csamul_cla32_fa19_25_xor1[0]), .cin(u_csamul_cla32_fa18_25_or0[0]), .fa_xor1(u_csamul_cla32_fa18_26_xor1), .fa_or0(u_csamul_cla32_fa18_26_or0));
  and_gate and_gate_u_csamul_cla32_and19_26(.a(a[19]), .b(b[26]), .out(u_csamul_cla32_and19_26));
  fa fa_u_csamul_cla32_fa19_26_out(.a(u_csamul_cla32_and19_26[0]), .b(u_csamul_cla32_fa20_25_xor1[0]), .cin(u_csamul_cla32_fa19_25_or0[0]), .fa_xor1(u_csamul_cla32_fa19_26_xor1), .fa_or0(u_csamul_cla32_fa19_26_or0));
  and_gate and_gate_u_csamul_cla32_and20_26(.a(a[20]), .b(b[26]), .out(u_csamul_cla32_and20_26));
  fa fa_u_csamul_cla32_fa20_26_out(.a(u_csamul_cla32_and20_26[0]), .b(u_csamul_cla32_fa21_25_xor1[0]), .cin(u_csamul_cla32_fa20_25_or0[0]), .fa_xor1(u_csamul_cla32_fa20_26_xor1), .fa_or0(u_csamul_cla32_fa20_26_or0));
  and_gate and_gate_u_csamul_cla32_and21_26(.a(a[21]), .b(b[26]), .out(u_csamul_cla32_and21_26));
  fa fa_u_csamul_cla32_fa21_26_out(.a(u_csamul_cla32_and21_26[0]), .b(u_csamul_cla32_fa22_25_xor1[0]), .cin(u_csamul_cla32_fa21_25_or0[0]), .fa_xor1(u_csamul_cla32_fa21_26_xor1), .fa_or0(u_csamul_cla32_fa21_26_or0));
  and_gate and_gate_u_csamul_cla32_and22_26(.a(a[22]), .b(b[26]), .out(u_csamul_cla32_and22_26));
  fa fa_u_csamul_cla32_fa22_26_out(.a(u_csamul_cla32_and22_26[0]), .b(u_csamul_cla32_fa23_25_xor1[0]), .cin(u_csamul_cla32_fa22_25_or0[0]), .fa_xor1(u_csamul_cla32_fa22_26_xor1), .fa_or0(u_csamul_cla32_fa22_26_or0));
  and_gate and_gate_u_csamul_cla32_and23_26(.a(a[23]), .b(b[26]), .out(u_csamul_cla32_and23_26));
  fa fa_u_csamul_cla32_fa23_26_out(.a(u_csamul_cla32_and23_26[0]), .b(u_csamul_cla32_fa24_25_xor1[0]), .cin(u_csamul_cla32_fa23_25_or0[0]), .fa_xor1(u_csamul_cla32_fa23_26_xor1), .fa_or0(u_csamul_cla32_fa23_26_or0));
  and_gate and_gate_u_csamul_cla32_and24_26(.a(a[24]), .b(b[26]), .out(u_csamul_cla32_and24_26));
  fa fa_u_csamul_cla32_fa24_26_out(.a(u_csamul_cla32_and24_26[0]), .b(u_csamul_cla32_fa25_25_xor1[0]), .cin(u_csamul_cla32_fa24_25_or0[0]), .fa_xor1(u_csamul_cla32_fa24_26_xor1), .fa_or0(u_csamul_cla32_fa24_26_or0));
  and_gate and_gate_u_csamul_cla32_and25_26(.a(a[25]), .b(b[26]), .out(u_csamul_cla32_and25_26));
  fa fa_u_csamul_cla32_fa25_26_out(.a(u_csamul_cla32_and25_26[0]), .b(u_csamul_cla32_fa26_25_xor1[0]), .cin(u_csamul_cla32_fa25_25_or0[0]), .fa_xor1(u_csamul_cla32_fa25_26_xor1), .fa_or0(u_csamul_cla32_fa25_26_or0));
  and_gate and_gate_u_csamul_cla32_and26_26(.a(a[26]), .b(b[26]), .out(u_csamul_cla32_and26_26));
  fa fa_u_csamul_cla32_fa26_26_out(.a(u_csamul_cla32_and26_26[0]), .b(u_csamul_cla32_fa27_25_xor1[0]), .cin(u_csamul_cla32_fa26_25_or0[0]), .fa_xor1(u_csamul_cla32_fa26_26_xor1), .fa_or0(u_csamul_cla32_fa26_26_or0));
  and_gate and_gate_u_csamul_cla32_and27_26(.a(a[27]), .b(b[26]), .out(u_csamul_cla32_and27_26));
  fa fa_u_csamul_cla32_fa27_26_out(.a(u_csamul_cla32_and27_26[0]), .b(u_csamul_cla32_fa28_25_xor1[0]), .cin(u_csamul_cla32_fa27_25_or0[0]), .fa_xor1(u_csamul_cla32_fa27_26_xor1), .fa_or0(u_csamul_cla32_fa27_26_or0));
  and_gate and_gate_u_csamul_cla32_and28_26(.a(a[28]), .b(b[26]), .out(u_csamul_cla32_and28_26));
  fa fa_u_csamul_cla32_fa28_26_out(.a(u_csamul_cla32_and28_26[0]), .b(u_csamul_cla32_fa29_25_xor1[0]), .cin(u_csamul_cla32_fa28_25_or0[0]), .fa_xor1(u_csamul_cla32_fa28_26_xor1), .fa_or0(u_csamul_cla32_fa28_26_or0));
  and_gate and_gate_u_csamul_cla32_and29_26(.a(a[29]), .b(b[26]), .out(u_csamul_cla32_and29_26));
  fa fa_u_csamul_cla32_fa29_26_out(.a(u_csamul_cla32_and29_26[0]), .b(u_csamul_cla32_fa30_25_xor1[0]), .cin(u_csamul_cla32_fa29_25_or0[0]), .fa_xor1(u_csamul_cla32_fa29_26_xor1), .fa_or0(u_csamul_cla32_fa29_26_or0));
  and_gate and_gate_u_csamul_cla32_and30_26(.a(a[30]), .b(b[26]), .out(u_csamul_cla32_and30_26));
  fa fa_u_csamul_cla32_fa30_26_out(.a(u_csamul_cla32_and30_26[0]), .b(u_csamul_cla32_and31_25[0]), .cin(u_csamul_cla32_fa30_25_or0[0]), .fa_xor1(u_csamul_cla32_fa30_26_xor1), .fa_or0(u_csamul_cla32_fa30_26_or0));
  and_gate and_gate_u_csamul_cla32_and31_26(.a(a[31]), .b(b[26]), .out(u_csamul_cla32_and31_26));
  and_gate and_gate_u_csamul_cla32_and0_27(.a(a[0]), .b(b[27]), .out(u_csamul_cla32_and0_27));
  fa fa_u_csamul_cla32_fa0_27_out(.a(u_csamul_cla32_and0_27[0]), .b(u_csamul_cla32_fa1_26_xor1[0]), .cin(u_csamul_cla32_fa0_26_or0[0]), .fa_xor1(u_csamul_cla32_fa0_27_xor1), .fa_or0(u_csamul_cla32_fa0_27_or0));
  and_gate and_gate_u_csamul_cla32_and1_27(.a(a[1]), .b(b[27]), .out(u_csamul_cla32_and1_27));
  fa fa_u_csamul_cla32_fa1_27_out(.a(u_csamul_cla32_and1_27[0]), .b(u_csamul_cla32_fa2_26_xor1[0]), .cin(u_csamul_cla32_fa1_26_or0[0]), .fa_xor1(u_csamul_cla32_fa1_27_xor1), .fa_or0(u_csamul_cla32_fa1_27_or0));
  and_gate and_gate_u_csamul_cla32_and2_27(.a(a[2]), .b(b[27]), .out(u_csamul_cla32_and2_27));
  fa fa_u_csamul_cla32_fa2_27_out(.a(u_csamul_cla32_and2_27[0]), .b(u_csamul_cla32_fa3_26_xor1[0]), .cin(u_csamul_cla32_fa2_26_or0[0]), .fa_xor1(u_csamul_cla32_fa2_27_xor1), .fa_or0(u_csamul_cla32_fa2_27_or0));
  and_gate and_gate_u_csamul_cla32_and3_27(.a(a[3]), .b(b[27]), .out(u_csamul_cla32_and3_27));
  fa fa_u_csamul_cla32_fa3_27_out(.a(u_csamul_cla32_and3_27[0]), .b(u_csamul_cla32_fa4_26_xor1[0]), .cin(u_csamul_cla32_fa3_26_or0[0]), .fa_xor1(u_csamul_cla32_fa3_27_xor1), .fa_or0(u_csamul_cla32_fa3_27_or0));
  and_gate and_gate_u_csamul_cla32_and4_27(.a(a[4]), .b(b[27]), .out(u_csamul_cla32_and4_27));
  fa fa_u_csamul_cla32_fa4_27_out(.a(u_csamul_cla32_and4_27[0]), .b(u_csamul_cla32_fa5_26_xor1[0]), .cin(u_csamul_cla32_fa4_26_or0[0]), .fa_xor1(u_csamul_cla32_fa4_27_xor1), .fa_or0(u_csamul_cla32_fa4_27_or0));
  and_gate and_gate_u_csamul_cla32_and5_27(.a(a[5]), .b(b[27]), .out(u_csamul_cla32_and5_27));
  fa fa_u_csamul_cla32_fa5_27_out(.a(u_csamul_cla32_and5_27[0]), .b(u_csamul_cla32_fa6_26_xor1[0]), .cin(u_csamul_cla32_fa5_26_or0[0]), .fa_xor1(u_csamul_cla32_fa5_27_xor1), .fa_or0(u_csamul_cla32_fa5_27_or0));
  and_gate and_gate_u_csamul_cla32_and6_27(.a(a[6]), .b(b[27]), .out(u_csamul_cla32_and6_27));
  fa fa_u_csamul_cla32_fa6_27_out(.a(u_csamul_cla32_and6_27[0]), .b(u_csamul_cla32_fa7_26_xor1[0]), .cin(u_csamul_cla32_fa6_26_or0[0]), .fa_xor1(u_csamul_cla32_fa6_27_xor1), .fa_or0(u_csamul_cla32_fa6_27_or0));
  and_gate and_gate_u_csamul_cla32_and7_27(.a(a[7]), .b(b[27]), .out(u_csamul_cla32_and7_27));
  fa fa_u_csamul_cla32_fa7_27_out(.a(u_csamul_cla32_and7_27[0]), .b(u_csamul_cla32_fa8_26_xor1[0]), .cin(u_csamul_cla32_fa7_26_or0[0]), .fa_xor1(u_csamul_cla32_fa7_27_xor1), .fa_or0(u_csamul_cla32_fa7_27_or0));
  and_gate and_gate_u_csamul_cla32_and8_27(.a(a[8]), .b(b[27]), .out(u_csamul_cla32_and8_27));
  fa fa_u_csamul_cla32_fa8_27_out(.a(u_csamul_cla32_and8_27[0]), .b(u_csamul_cla32_fa9_26_xor1[0]), .cin(u_csamul_cla32_fa8_26_or0[0]), .fa_xor1(u_csamul_cla32_fa8_27_xor1), .fa_or0(u_csamul_cla32_fa8_27_or0));
  and_gate and_gate_u_csamul_cla32_and9_27(.a(a[9]), .b(b[27]), .out(u_csamul_cla32_and9_27));
  fa fa_u_csamul_cla32_fa9_27_out(.a(u_csamul_cla32_and9_27[0]), .b(u_csamul_cla32_fa10_26_xor1[0]), .cin(u_csamul_cla32_fa9_26_or0[0]), .fa_xor1(u_csamul_cla32_fa9_27_xor1), .fa_or0(u_csamul_cla32_fa9_27_or0));
  and_gate and_gate_u_csamul_cla32_and10_27(.a(a[10]), .b(b[27]), .out(u_csamul_cla32_and10_27));
  fa fa_u_csamul_cla32_fa10_27_out(.a(u_csamul_cla32_and10_27[0]), .b(u_csamul_cla32_fa11_26_xor1[0]), .cin(u_csamul_cla32_fa10_26_or0[0]), .fa_xor1(u_csamul_cla32_fa10_27_xor1), .fa_or0(u_csamul_cla32_fa10_27_or0));
  and_gate and_gate_u_csamul_cla32_and11_27(.a(a[11]), .b(b[27]), .out(u_csamul_cla32_and11_27));
  fa fa_u_csamul_cla32_fa11_27_out(.a(u_csamul_cla32_and11_27[0]), .b(u_csamul_cla32_fa12_26_xor1[0]), .cin(u_csamul_cla32_fa11_26_or0[0]), .fa_xor1(u_csamul_cla32_fa11_27_xor1), .fa_or0(u_csamul_cla32_fa11_27_or0));
  and_gate and_gate_u_csamul_cla32_and12_27(.a(a[12]), .b(b[27]), .out(u_csamul_cla32_and12_27));
  fa fa_u_csamul_cla32_fa12_27_out(.a(u_csamul_cla32_and12_27[0]), .b(u_csamul_cla32_fa13_26_xor1[0]), .cin(u_csamul_cla32_fa12_26_or0[0]), .fa_xor1(u_csamul_cla32_fa12_27_xor1), .fa_or0(u_csamul_cla32_fa12_27_or0));
  and_gate and_gate_u_csamul_cla32_and13_27(.a(a[13]), .b(b[27]), .out(u_csamul_cla32_and13_27));
  fa fa_u_csamul_cla32_fa13_27_out(.a(u_csamul_cla32_and13_27[0]), .b(u_csamul_cla32_fa14_26_xor1[0]), .cin(u_csamul_cla32_fa13_26_or0[0]), .fa_xor1(u_csamul_cla32_fa13_27_xor1), .fa_or0(u_csamul_cla32_fa13_27_or0));
  and_gate and_gate_u_csamul_cla32_and14_27(.a(a[14]), .b(b[27]), .out(u_csamul_cla32_and14_27));
  fa fa_u_csamul_cla32_fa14_27_out(.a(u_csamul_cla32_and14_27[0]), .b(u_csamul_cla32_fa15_26_xor1[0]), .cin(u_csamul_cla32_fa14_26_or0[0]), .fa_xor1(u_csamul_cla32_fa14_27_xor1), .fa_or0(u_csamul_cla32_fa14_27_or0));
  and_gate and_gate_u_csamul_cla32_and15_27(.a(a[15]), .b(b[27]), .out(u_csamul_cla32_and15_27));
  fa fa_u_csamul_cla32_fa15_27_out(.a(u_csamul_cla32_and15_27[0]), .b(u_csamul_cla32_fa16_26_xor1[0]), .cin(u_csamul_cla32_fa15_26_or0[0]), .fa_xor1(u_csamul_cla32_fa15_27_xor1), .fa_or0(u_csamul_cla32_fa15_27_or0));
  and_gate and_gate_u_csamul_cla32_and16_27(.a(a[16]), .b(b[27]), .out(u_csamul_cla32_and16_27));
  fa fa_u_csamul_cla32_fa16_27_out(.a(u_csamul_cla32_and16_27[0]), .b(u_csamul_cla32_fa17_26_xor1[0]), .cin(u_csamul_cla32_fa16_26_or0[0]), .fa_xor1(u_csamul_cla32_fa16_27_xor1), .fa_or0(u_csamul_cla32_fa16_27_or0));
  and_gate and_gate_u_csamul_cla32_and17_27(.a(a[17]), .b(b[27]), .out(u_csamul_cla32_and17_27));
  fa fa_u_csamul_cla32_fa17_27_out(.a(u_csamul_cla32_and17_27[0]), .b(u_csamul_cla32_fa18_26_xor1[0]), .cin(u_csamul_cla32_fa17_26_or0[0]), .fa_xor1(u_csamul_cla32_fa17_27_xor1), .fa_or0(u_csamul_cla32_fa17_27_or0));
  and_gate and_gate_u_csamul_cla32_and18_27(.a(a[18]), .b(b[27]), .out(u_csamul_cla32_and18_27));
  fa fa_u_csamul_cla32_fa18_27_out(.a(u_csamul_cla32_and18_27[0]), .b(u_csamul_cla32_fa19_26_xor1[0]), .cin(u_csamul_cla32_fa18_26_or0[0]), .fa_xor1(u_csamul_cla32_fa18_27_xor1), .fa_or0(u_csamul_cla32_fa18_27_or0));
  and_gate and_gate_u_csamul_cla32_and19_27(.a(a[19]), .b(b[27]), .out(u_csamul_cla32_and19_27));
  fa fa_u_csamul_cla32_fa19_27_out(.a(u_csamul_cla32_and19_27[0]), .b(u_csamul_cla32_fa20_26_xor1[0]), .cin(u_csamul_cla32_fa19_26_or0[0]), .fa_xor1(u_csamul_cla32_fa19_27_xor1), .fa_or0(u_csamul_cla32_fa19_27_or0));
  and_gate and_gate_u_csamul_cla32_and20_27(.a(a[20]), .b(b[27]), .out(u_csamul_cla32_and20_27));
  fa fa_u_csamul_cla32_fa20_27_out(.a(u_csamul_cla32_and20_27[0]), .b(u_csamul_cla32_fa21_26_xor1[0]), .cin(u_csamul_cla32_fa20_26_or0[0]), .fa_xor1(u_csamul_cla32_fa20_27_xor1), .fa_or0(u_csamul_cla32_fa20_27_or0));
  and_gate and_gate_u_csamul_cla32_and21_27(.a(a[21]), .b(b[27]), .out(u_csamul_cla32_and21_27));
  fa fa_u_csamul_cla32_fa21_27_out(.a(u_csamul_cla32_and21_27[0]), .b(u_csamul_cla32_fa22_26_xor1[0]), .cin(u_csamul_cla32_fa21_26_or0[0]), .fa_xor1(u_csamul_cla32_fa21_27_xor1), .fa_or0(u_csamul_cla32_fa21_27_or0));
  and_gate and_gate_u_csamul_cla32_and22_27(.a(a[22]), .b(b[27]), .out(u_csamul_cla32_and22_27));
  fa fa_u_csamul_cla32_fa22_27_out(.a(u_csamul_cla32_and22_27[0]), .b(u_csamul_cla32_fa23_26_xor1[0]), .cin(u_csamul_cla32_fa22_26_or0[0]), .fa_xor1(u_csamul_cla32_fa22_27_xor1), .fa_or0(u_csamul_cla32_fa22_27_or0));
  and_gate and_gate_u_csamul_cla32_and23_27(.a(a[23]), .b(b[27]), .out(u_csamul_cla32_and23_27));
  fa fa_u_csamul_cla32_fa23_27_out(.a(u_csamul_cla32_and23_27[0]), .b(u_csamul_cla32_fa24_26_xor1[0]), .cin(u_csamul_cla32_fa23_26_or0[0]), .fa_xor1(u_csamul_cla32_fa23_27_xor1), .fa_or0(u_csamul_cla32_fa23_27_or0));
  and_gate and_gate_u_csamul_cla32_and24_27(.a(a[24]), .b(b[27]), .out(u_csamul_cla32_and24_27));
  fa fa_u_csamul_cla32_fa24_27_out(.a(u_csamul_cla32_and24_27[0]), .b(u_csamul_cla32_fa25_26_xor1[0]), .cin(u_csamul_cla32_fa24_26_or0[0]), .fa_xor1(u_csamul_cla32_fa24_27_xor1), .fa_or0(u_csamul_cla32_fa24_27_or0));
  and_gate and_gate_u_csamul_cla32_and25_27(.a(a[25]), .b(b[27]), .out(u_csamul_cla32_and25_27));
  fa fa_u_csamul_cla32_fa25_27_out(.a(u_csamul_cla32_and25_27[0]), .b(u_csamul_cla32_fa26_26_xor1[0]), .cin(u_csamul_cla32_fa25_26_or0[0]), .fa_xor1(u_csamul_cla32_fa25_27_xor1), .fa_or0(u_csamul_cla32_fa25_27_or0));
  and_gate and_gate_u_csamul_cla32_and26_27(.a(a[26]), .b(b[27]), .out(u_csamul_cla32_and26_27));
  fa fa_u_csamul_cla32_fa26_27_out(.a(u_csamul_cla32_and26_27[0]), .b(u_csamul_cla32_fa27_26_xor1[0]), .cin(u_csamul_cla32_fa26_26_or0[0]), .fa_xor1(u_csamul_cla32_fa26_27_xor1), .fa_or0(u_csamul_cla32_fa26_27_or0));
  and_gate and_gate_u_csamul_cla32_and27_27(.a(a[27]), .b(b[27]), .out(u_csamul_cla32_and27_27));
  fa fa_u_csamul_cla32_fa27_27_out(.a(u_csamul_cla32_and27_27[0]), .b(u_csamul_cla32_fa28_26_xor1[0]), .cin(u_csamul_cla32_fa27_26_or0[0]), .fa_xor1(u_csamul_cla32_fa27_27_xor1), .fa_or0(u_csamul_cla32_fa27_27_or0));
  and_gate and_gate_u_csamul_cla32_and28_27(.a(a[28]), .b(b[27]), .out(u_csamul_cla32_and28_27));
  fa fa_u_csamul_cla32_fa28_27_out(.a(u_csamul_cla32_and28_27[0]), .b(u_csamul_cla32_fa29_26_xor1[0]), .cin(u_csamul_cla32_fa28_26_or0[0]), .fa_xor1(u_csamul_cla32_fa28_27_xor1), .fa_or0(u_csamul_cla32_fa28_27_or0));
  and_gate and_gate_u_csamul_cla32_and29_27(.a(a[29]), .b(b[27]), .out(u_csamul_cla32_and29_27));
  fa fa_u_csamul_cla32_fa29_27_out(.a(u_csamul_cla32_and29_27[0]), .b(u_csamul_cla32_fa30_26_xor1[0]), .cin(u_csamul_cla32_fa29_26_or0[0]), .fa_xor1(u_csamul_cla32_fa29_27_xor1), .fa_or0(u_csamul_cla32_fa29_27_or0));
  and_gate and_gate_u_csamul_cla32_and30_27(.a(a[30]), .b(b[27]), .out(u_csamul_cla32_and30_27));
  fa fa_u_csamul_cla32_fa30_27_out(.a(u_csamul_cla32_and30_27[0]), .b(u_csamul_cla32_and31_26[0]), .cin(u_csamul_cla32_fa30_26_or0[0]), .fa_xor1(u_csamul_cla32_fa30_27_xor1), .fa_or0(u_csamul_cla32_fa30_27_or0));
  and_gate and_gate_u_csamul_cla32_and31_27(.a(a[31]), .b(b[27]), .out(u_csamul_cla32_and31_27));
  and_gate and_gate_u_csamul_cla32_and0_28(.a(a[0]), .b(b[28]), .out(u_csamul_cla32_and0_28));
  fa fa_u_csamul_cla32_fa0_28_out(.a(u_csamul_cla32_and0_28[0]), .b(u_csamul_cla32_fa1_27_xor1[0]), .cin(u_csamul_cla32_fa0_27_or0[0]), .fa_xor1(u_csamul_cla32_fa0_28_xor1), .fa_or0(u_csamul_cla32_fa0_28_or0));
  and_gate and_gate_u_csamul_cla32_and1_28(.a(a[1]), .b(b[28]), .out(u_csamul_cla32_and1_28));
  fa fa_u_csamul_cla32_fa1_28_out(.a(u_csamul_cla32_and1_28[0]), .b(u_csamul_cla32_fa2_27_xor1[0]), .cin(u_csamul_cla32_fa1_27_or0[0]), .fa_xor1(u_csamul_cla32_fa1_28_xor1), .fa_or0(u_csamul_cla32_fa1_28_or0));
  and_gate and_gate_u_csamul_cla32_and2_28(.a(a[2]), .b(b[28]), .out(u_csamul_cla32_and2_28));
  fa fa_u_csamul_cla32_fa2_28_out(.a(u_csamul_cla32_and2_28[0]), .b(u_csamul_cla32_fa3_27_xor1[0]), .cin(u_csamul_cla32_fa2_27_or0[0]), .fa_xor1(u_csamul_cla32_fa2_28_xor1), .fa_or0(u_csamul_cla32_fa2_28_or0));
  and_gate and_gate_u_csamul_cla32_and3_28(.a(a[3]), .b(b[28]), .out(u_csamul_cla32_and3_28));
  fa fa_u_csamul_cla32_fa3_28_out(.a(u_csamul_cla32_and3_28[0]), .b(u_csamul_cla32_fa4_27_xor1[0]), .cin(u_csamul_cla32_fa3_27_or0[0]), .fa_xor1(u_csamul_cla32_fa3_28_xor1), .fa_or0(u_csamul_cla32_fa3_28_or0));
  and_gate and_gate_u_csamul_cla32_and4_28(.a(a[4]), .b(b[28]), .out(u_csamul_cla32_and4_28));
  fa fa_u_csamul_cla32_fa4_28_out(.a(u_csamul_cla32_and4_28[0]), .b(u_csamul_cla32_fa5_27_xor1[0]), .cin(u_csamul_cla32_fa4_27_or0[0]), .fa_xor1(u_csamul_cla32_fa4_28_xor1), .fa_or0(u_csamul_cla32_fa4_28_or0));
  and_gate and_gate_u_csamul_cla32_and5_28(.a(a[5]), .b(b[28]), .out(u_csamul_cla32_and5_28));
  fa fa_u_csamul_cla32_fa5_28_out(.a(u_csamul_cla32_and5_28[0]), .b(u_csamul_cla32_fa6_27_xor1[0]), .cin(u_csamul_cla32_fa5_27_or0[0]), .fa_xor1(u_csamul_cla32_fa5_28_xor1), .fa_or0(u_csamul_cla32_fa5_28_or0));
  and_gate and_gate_u_csamul_cla32_and6_28(.a(a[6]), .b(b[28]), .out(u_csamul_cla32_and6_28));
  fa fa_u_csamul_cla32_fa6_28_out(.a(u_csamul_cla32_and6_28[0]), .b(u_csamul_cla32_fa7_27_xor1[0]), .cin(u_csamul_cla32_fa6_27_or0[0]), .fa_xor1(u_csamul_cla32_fa6_28_xor1), .fa_or0(u_csamul_cla32_fa6_28_or0));
  and_gate and_gate_u_csamul_cla32_and7_28(.a(a[7]), .b(b[28]), .out(u_csamul_cla32_and7_28));
  fa fa_u_csamul_cla32_fa7_28_out(.a(u_csamul_cla32_and7_28[0]), .b(u_csamul_cla32_fa8_27_xor1[0]), .cin(u_csamul_cla32_fa7_27_or0[0]), .fa_xor1(u_csamul_cla32_fa7_28_xor1), .fa_or0(u_csamul_cla32_fa7_28_or0));
  and_gate and_gate_u_csamul_cla32_and8_28(.a(a[8]), .b(b[28]), .out(u_csamul_cla32_and8_28));
  fa fa_u_csamul_cla32_fa8_28_out(.a(u_csamul_cla32_and8_28[0]), .b(u_csamul_cla32_fa9_27_xor1[0]), .cin(u_csamul_cla32_fa8_27_or0[0]), .fa_xor1(u_csamul_cla32_fa8_28_xor1), .fa_or0(u_csamul_cla32_fa8_28_or0));
  and_gate and_gate_u_csamul_cla32_and9_28(.a(a[9]), .b(b[28]), .out(u_csamul_cla32_and9_28));
  fa fa_u_csamul_cla32_fa9_28_out(.a(u_csamul_cla32_and9_28[0]), .b(u_csamul_cla32_fa10_27_xor1[0]), .cin(u_csamul_cla32_fa9_27_or0[0]), .fa_xor1(u_csamul_cla32_fa9_28_xor1), .fa_or0(u_csamul_cla32_fa9_28_or0));
  and_gate and_gate_u_csamul_cla32_and10_28(.a(a[10]), .b(b[28]), .out(u_csamul_cla32_and10_28));
  fa fa_u_csamul_cla32_fa10_28_out(.a(u_csamul_cla32_and10_28[0]), .b(u_csamul_cla32_fa11_27_xor1[0]), .cin(u_csamul_cla32_fa10_27_or0[0]), .fa_xor1(u_csamul_cla32_fa10_28_xor1), .fa_or0(u_csamul_cla32_fa10_28_or0));
  and_gate and_gate_u_csamul_cla32_and11_28(.a(a[11]), .b(b[28]), .out(u_csamul_cla32_and11_28));
  fa fa_u_csamul_cla32_fa11_28_out(.a(u_csamul_cla32_and11_28[0]), .b(u_csamul_cla32_fa12_27_xor1[0]), .cin(u_csamul_cla32_fa11_27_or0[0]), .fa_xor1(u_csamul_cla32_fa11_28_xor1), .fa_or0(u_csamul_cla32_fa11_28_or0));
  and_gate and_gate_u_csamul_cla32_and12_28(.a(a[12]), .b(b[28]), .out(u_csamul_cla32_and12_28));
  fa fa_u_csamul_cla32_fa12_28_out(.a(u_csamul_cla32_and12_28[0]), .b(u_csamul_cla32_fa13_27_xor1[0]), .cin(u_csamul_cla32_fa12_27_or0[0]), .fa_xor1(u_csamul_cla32_fa12_28_xor1), .fa_or0(u_csamul_cla32_fa12_28_or0));
  and_gate and_gate_u_csamul_cla32_and13_28(.a(a[13]), .b(b[28]), .out(u_csamul_cla32_and13_28));
  fa fa_u_csamul_cla32_fa13_28_out(.a(u_csamul_cla32_and13_28[0]), .b(u_csamul_cla32_fa14_27_xor1[0]), .cin(u_csamul_cla32_fa13_27_or0[0]), .fa_xor1(u_csamul_cla32_fa13_28_xor1), .fa_or0(u_csamul_cla32_fa13_28_or0));
  and_gate and_gate_u_csamul_cla32_and14_28(.a(a[14]), .b(b[28]), .out(u_csamul_cla32_and14_28));
  fa fa_u_csamul_cla32_fa14_28_out(.a(u_csamul_cla32_and14_28[0]), .b(u_csamul_cla32_fa15_27_xor1[0]), .cin(u_csamul_cla32_fa14_27_or0[0]), .fa_xor1(u_csamul_cla32_fa14_28_xor1), .fa_or0(u_csamul_cla32_fa14_28_or0));
  and_gate and_gate_u_csamul_cla32_and15_28(.a(a[15]), .b(b[28]), .out(u_csamul_cla32_and15_28));
  fa fa_u_csamul_cla32_fa15_28_out(.a(u_csamul_cla32_and15_28[0]), .b(u_csamul_cla32_fa16_27_xor1[0]), .cin(u_csamul_cla32_fa15_27_or0[0]), .fa_xor1(u_csamul_cla32_fa15_28_xor1), .fa_or0(u_csamul_cla32_fa15_28_or0));
  and_gate and_gate_u_csamul_cla32_and16_28(.a(a[16]), .b(b[28]), .out(u_csamul_cla32_and16_28));
  fa fa_u_csamul_cla32_fa16_28_out(.a(u_csamul_cla32_and16_28[0]), .b(u_csamul_cla32_fa17_27_xor1[0]), .cin(u_csamul_cla32_fa16_27_or0[0]), .fa_xor1(u_csamul_cla32_fa16_28_xor1), .fa_or0(u_csamul_cla32_fa16_28_or0));
  and_gate and_gate_u_csamul_cla32_and17_28(.a(a[17]), .b(b[28]), .out(u_csamul_cla32_and17_28));
  fa fa_u_csamul_cla32_fa17_28_out(.a(u_csamul_cla32_and17_28[0]), .b(u_csamul_cla32_fa18_27_xor1[0]), .cin(u_csamul_cla32_fa17_27_or0[0]), .fa_xor1(u_csamul_cla32_fa17_28_xor1), .fa_or0(u_csamul_cla32_fa17_28_or0));
  and_gate and_gate_u_csamul_cla32_and18_28(.a(a[18]), .b(b[28]), .out(u_csamul_cla32_and18_28));
  fa fa_u_csamul_cla32_fa18_28_out(.a(u_csamul_cla32_and18_28[0]), .b(u_csamul_cla32_fa19_27_xor1[0]), .cin(u_csamul_cla32_fa18_27_or0[0]), .fa_xor1(u_csamul_cla32_fa18_28_xor1), .fa_or0(u_csamul_cla32_fa18_28_or0));
  and_gate and_gate_u_csamul_cla32_and19_28(.a(a[19]), .b(b[28]), .out(u_csamul_cla32_and19_28));
  fa fa_u_csamul_cla32_fa19_28_out(.a(u_csamul_cla32_and19_28[0]), .b(u_csamul_cla32_fa20_27_xor1[0]), .cin(u_csamul_cla32_fa19_27_or0[0]), .fa_xor1(u_csamul_cla32_fa19_28_xor1), .fa_or0(u_csamul_cla32_fa19_28_or0));
  and_gate and_gate_u_csamul_cla32_and20_28(.a(a[20]), .b(b[28]), .out(u_csamul_cla32_and20_28));
  fa fa_u_csamul_cla32_fa20_28_out(.a(u_csamul_cla32_and20_28[0]), .b(u_csamul_cla32_fa21_27_xor1[0]), .cin(u_csamul_cla32_fa20_27_or0[0]), .fa_xor1(u_csamul_cla32_fa20_28_xor1), .fa_or0(u_csamul_cla32_fa20_28_or0));
  and_gate and_gate_u_csamul_cla32_and21_28(.a(a[21]), .b(b[28]), .out(u_csamul_cla32_and21_28));
  fa fa_u_csamul_cla32_fa21_28_out(.a(u_csamul_cla32_and21_28[0]), .b(u_csamul_cla32_fa22_27_xor1[0]), .cin(u_csamul_cla32_fa21_27_or0[0]), .fa_xor1(u_csamul_cla32_fa21_28_xor1), .fa_or0(u_csamul_cla32_fa21_28_or0));
  and_gate and_gate_u_csamul_cla32_and22_28(.a(a[22]), .b(b[28]), .out(u_csamul_cla32_and22_28));
  fa fa_u_csamul_cla32_fa22_28_out(.a(u_csamul_cla32_and22_28[0]), .b(u_csamul_cla32_fa23_27_xor1[0]), .cin(u_csamul_cla32_fa22_27_or0[0]), .fa_xor1(u_csamul_cla32_fa22_28_xor1), .fa_or0(u_csamul_cla32_fa22_28_or0));
  and_gate and_gate_u_csamul_cla32_and23_28(.a(a[23]), .b(b[28]), .out(u_csamul_cla32_and23_28));
  fa fa_u_csamul_cla32_fa23_28_out(.a(u_csamul_cla32_and23_28[0]), .b(u_csamul_cla32_fa24_27_xor1[0]), .cin(u_csamul_cla32_fa23_27_or0[0]), .fa_xor1(u_csamul_cla32_fa23_28_xor1), .fa_or0(u_csamul_cla32_fa23_28_or0));
  and_gate and_gate_u_csamul_cla32_and24_28(.a(a[24]), .b(b[28]), .out(u_csamul_cla32_and24_28));
  fa fa_u_csamul_cla32_fa24_28_out(.a(u_csamul_cla32_and24_28[0]), .b(u_csamul_cla32_fa25_27_xor1[0]), .cin(u_csamul_cla32_fa24_27_or0[0]), .fa_xor1(u_csamul_cla32_fa24_28_xor1), .fa_or0(u_csamul_cla32_fa24_28_or0));
  and_gate and_gate_u_csamul_cla32_and25_28(.a(a[25]), .b(b[28]), .out(u_csamul_cla32_and25_28));
  fa fa_u_csamul_cla32_fa25_28_out(.a(u_csamul_cla32_and25_28[0]), .b(u_csamul_cla32_fa26_27_xor1[0]), .cin(u_csamul_cla32_fa25_27_or0[0]), .fa_xor1(u_csamul_cla32_fa25_28_xor1), .fa_or0(u_csamul_cla32_fa25_28_or0));
  and_gate and_gate_u_csamul_cla32_and26_28(.a(a[26]), .b(b[28]), .out(u_csamul_cla32_and26_28));
  fa fa_u_csamul_cla32_fa26_28_out(.a(u_csamul_cla32_and26_28[0]), .b(u_csamul_cla32_fa27_27_xor1[0]), .cin(u_csamul_cla32_fa26_27_or0[0]), .fa_xor1(u_csamul_cla32_fa26_28_xor1), .fa_or0(u_csamul_cla32_fa26_28_or0));
  and_gate and_gate_u_csamul_cla32_and27_28(.a(a[27]), .b(b[28]), .out(u_csamul_cla32_and27_28));
  fa fa_u_csamul_cla32_fa27_28_out(.a(u_csamul_cla32_and27_28[0]), .b(u_csamul_cla32_fa28_27_xor1[0]), .cin(u_csamul_cla32_fa27_27_or0[0]), .fa_xor1(u_csamul_cla32_fa27_28_xor1), .fa_or0(u_csamul_cla32_fa27_28_or0));
  and_gate and_gate_u_csamul_cla32_and28_28(.a(a[28]), .b(b[28]), .out(u_csamul_cla32_and28_28));
  fa fa_u_csamul_cla32_fa28_28_out(.a(u_csamul_cla32_and28_28[0]), .b(u_csamul_cla32_fa29_27_xor1[0]), .cin(u_csamul_cla32_fa28_27_or0[0]), .fa_xor1(u_csamul_cla32_fa28_28_xor1), .fa_or0(u_csamul_cla32_fa28_28_or0));
  and_gate and_gate_u_csamul_cla32_and29_28(.a(a[29]), .b(b[28]), .out(u_csamul_cla32_and29_28));
  fa fa_u_csamul_cla32_fa29_28_out(.a(u_csamul_cla32_and29_28[0]), .b(u_csamul_cla32_fa30_27_xor1[0]), .cin(u_csamul_cla32_fa29_27_or0[0]), .fa_xor1(u_csamul_cla32_fa29_28_xor1), .fa_or0(u_csamul_cla32_fa29_28_or0));
  and_gate and_gate_u_csamul_cla32_and30_28(.a(a[30]), .b(b[28]), .out(u_csamul_cla32_and30_28));
  fa fa_u_csamul_cla32_fa30_28_out(.a(u_csamul_cla32_and30_28[0]), .b(u_csamul_cla32_and31_27[0]), .cin(u_csamul_cla32_fa30_27_or0[0]), .fa_xor1(u_csamul_cla32_fa30_28_xor1), .fa_or0(u_csamul_cla32_fa30_28_or0));
  and_gate and_gate_u_csamul_cla32_and31_28(.a(a[31]), .b(b[28]), .out(u_csamul_cla32_and31_28));
  and_gate and_gate_u_csamul_cla32_and0_29(.a(a[0]), .b(b[29]), .out(u_csamul_cla32_and0_29));
  fa fa_u_csamul_cla32_fa0_29_out(.a(u_csamul_cla32_and0_29[0]), .b(u_csamul_cla32_fa1_28_xor1[0]), .cin(u_csamul_cla32_fa0_28_or0[0]), .fa_xor1(u_csamul_cla32_fa0_29_xor1), .fa_or0(u_csamul_cla32_fa0_29_or0));
  and_gate and_gate_u_csamul_cla32_and1_29(.a(a[1]), .b(b[29]), .out(u_csamul_cla32_and1_29));
  fa fa_u_csamul_cla32_fa1_29_out(.a(u_csamul_cla32_and1_29[0]), .b(u_csamul_cla32_fa2_28_xor1[0]), .cin(u_csamul_cla32_fa1_28_or0[0]), .fa_xor1(u_csamul_cla32_fa1_29_xor1), .fa_or0(u_csamul_cla32_fa1_29_or0));
  and_gate and_gate_u_csamul_cla32_and2_29(.a(a[2]), .b(b[29]), .out(u_csamul_cla32_and2_29));
  fa fa_u_csamul_cla32_fa2_29_out(.a(u_csamul_cla32_and2_29[0]), .b(u_csamul_cla32_fa3_28_xor1[0]), .cin(u_csamul_cla32_fa2_28_or0[0]), .fa_xor1(u_csamul_cla32_fa2_29_xor1), .fa_or0(u_csamul_cla32_fa2_29_or0));
  and_gate and_gate_u_csamul_cla32_and3_29(.a(a[3]), .b(b[29]), .out(u_csamul_cla32_and3_29));
  fa fa_u_csamul_cla32_fa3_29_out(.a(u_csamul_cla32_and3_29[0]), .b(u_csamul_cla32_fa4_28_xor1[0]), .cin(u_csamul_cla32_fa3_28_or0[0]), .fa_xor1(u_csamul_cla32_fa3_29_xor1), .fa_or0(u_csamul_cla32_fa3_29_or0));
  and_gate and_gate_u_csamul_cla32_and4_29(.a(a[4]), .b(b[29]), .out(u_csamul_cla32_and4_29));
  fa fa_u_csamul_cla32_fa4_29_out(.a(u_csamul_cla32_and4_29[0]), .b(u_csamul_cla32_fa5_28_xor1[0]), .cin(u_csamul_cla32_fa4_28_or0[0]), .fa_xor1(u_csamul_cla32_fa4_29_xor1), .fa_or0(u_csamul_cla32_fa4_29_or0));
  and_gate and_gate_u_csamul_cla32_and5_29(.a(a[5]), .b(b[29]), .out(u_csamul_cla32_and5_29));
  fa fa_u_csamul_cla32_fa5_29_out(.a(u_csamul_cla32_and5_29[0]), .b(u_csamul_cla32_fa6_28_xor1[0]), .cin(u_csamul_cla32_fa5_28_or0[0]), .fa_xor1(u_csamul_cla32_fa5_29_xor1), .fa_or0(u_csamul_cla32_fa5_29_or0));
  and_gate and_gate_u_csamul_cla32_and6_29(.a(a[6]), .b(b[29]), .out(u_csamul_cla32_and6_29));
  fa fa_u_csamul_cla32_fa6_29_out(.a(u_csamul_cla32_and6_29[0]), .b(u_csamul_cla32_fa7_28_xor1[0]), .cin(u_csamul_cla32_fa6_28_or0[0]), .fa_xor1(u_csamul_cla32_fa6_29_xor1), .fa_or0(u_csamul_cla32_fa6_29_or0));
  and_gate and_gate_u_csamul_cla32_and7_29(.a(a[7]), .b(b[29]), .out(u_csamul_cla32_and7_29));
  fa fa_u_csamul_cla32_fa7_29_out(.a(u_csamul_cla32_and7_29[0]), .b(u_csamul_cla32_fa8_28_xor1[0]), .cin(u_csamul_cla32_fa7_28_or0[0]), .fa_xor1(u_csamul_cla32_fa7_29_xor1), .fa_or0(u_csamul_cla32_fa7_29_or0));
  and_gate and_gate_u_csamul_cla32_and8_29(.a(a[8]), .b(b[29]), .out(u_csamul_cla32_and8_29));
  fa fa_u_csamul_cla32_fa8_29_out(.a(u_csamul_cla32_and8_29[0]), .b(u_csamul_cla32_fa9_28_xor1[0]), .cin(u_csamul_cla32_fa8_28_or0[0]), .fa_xor1(u_csamul_cla32_fa8_29_xor1), .fa_or0(u_csamul_cla32_fa8_29_or0));
  and_gate and_gate_u_csamul_cla32_and9_29(.a(a[9]), .b(b[29]), .out(u_csamul_cla32_and9_29));
  fa fa_u_csamul_cla32_fa9_29_out(.a(u_csamul_cla32_and9_29[0]), .b(u_csamul_cla32_fa10_28_xor1[0]), .cin(u_csamul_cla32_fa9_28_or0[0]), .fa_xor1(u_csamul_cla32_fa9_29_xor1), .fa_or0(u_csamul_cla32_fa9_29_or0));
  and_gate and_gate_u_csamul_cla32_and10_29(.a(a[10]), .b(b[29]), .out(u_csamul_cla32_and10_29));
  fa fa_u_csamul_cla32_fa10_29_out(.a(u_csamul_cla32_and10_29[0]), .b(u_csamul_cla32_fa11_28_xor1[0]), .cin(u_csamul_cla32_fa10_28_or0[0]), .fa_xor1(u_csamul_cla32_fa10_29_xor1), .fa_or0(u_csamul_cla32_fa10_29_or0));
  and_gate and_gate_u_csamul_cla32_and11_29(.a(a[11]), .b(b[29]), .out(u_csamul_cla32_and11_29));
  fa fa_u_csamul_cla32_fa11_29_out(.a(u_csamul_cla32_and11_29[0]), .b(u_csamul_cla32_fa12_28_xor1[0]), .cin(u_csamul_cla32_fa11_28_or0[0]), .fa_xor1(u_csamul_cla32_fa11_29_xor1), .fa_or0(u_csamul_cla32_fa11_29_or0));
  and_gate and_gate_u_csamul_cla32_and12_29(.a(a[12]), .b(b[29]), .out(u_csamul_cla32_and12_29));
  fa fa_u_csamul_cla32_fa12_29_out(.a(u_csamul_cla32_and12_29[0]), .b(u_csamul_cla32_fa13_28_xor1[0]), .cin(u_csamul_cla32_fa12_28_or0[0]), .fa_xor1(u_csamul_cla32_fa12_29_xor1), .fa_or0(u_csamul_cla32_fa12_29_or0));
  and_gate and_gate_u_csamul_cla32_and13_29(.a(a[13]), .b(b[29]), .out(u_csamul_cla32_and13_29));
  fa fa_u_csamul_cla32_fa13_29_out(.a(u_csamul_cla32_and13_29[0]), .b(u_csamul_cla32_fa14_28_xor1[0]), .cin(u_csamul_cla32_fa13_28_or0[0]), .fa_xor1(u_csamul_cla32_fa13_29_xor1), .fa_or0(u_csamul_cla32_fa13_29_or0));
  and_gate and_gate_u_csamul_cla32_and14_29(.a(a[14]), .b(b[29]), .out(u_csamul_cla32_and14_29));
  fa fa_u_csamul_cla32_fa14_29_out(.a(u_csamul_cla32_and14_29[0]), .b(u_csamul_cla32_fa15_28_xor1[0]), .cin(u_csamul_cla32_fa14_28_or0[0]), .fa_xor1(u_csamul_cla32_fa14_29_xor1), .fa_or0(u_csamul_cla32_fa14_29_or0));
  and_gate and_gate_u_csamul_cla32_and15_29(.a(a[15]), .b(b[29]), .out(u_csamul_cla32_and15_29));
  fa fa_u_csamul_cla32_fa15_29_out(.a(u_csamul_cla32_and15_29[0]), .b(u_csamul_cla32_fa16_28_xor1[0]), .cin(u_csamul_cla32_fa15_28_or0[0]), .fa_xor1(u_csamul_cla32_fa15_29_xor1), .fa_or0(u_csamul_cla32_fa15_29_or0));
  and_gate and_gate_u_csamul_cla32_and16_29(.a(a[16]), .b(b[29]), .out(u_csamul_cla32_and16_29));
  fa fa_u_csamul_cla32_fa16_29_out(.a(u_csamul_cla32_and16_29[0]), .b(u_csamul_cla32_fa17_28_xor1[0]), .cin(u_csamul_cla32_fa16_28_or0[0]), .fa_xor1(u_csamul_cla32_fa16_29_xor1), .fa_or0(u_csamul_cla32_fa16_29_or0));
  and_gate and_gate_u_csamul_cla32_and17_29(.a(a[17]), .b(b[29]), .out(u_csamul_cla32_and17_29));
  fa fa_u_csamul_cla32_fa17_29_out(.a(u_csamul_cla32_and17_29[0]), .b(u_csamul_cla32_fa18_28_xor1[0]), .cin(u_csamul_cla32_fa17_28_or0[0]), .fa_xor1(u_csamul_cla32_fa17_29_xor1), .fa_or0(u_csamul_cla32_fa17_29_or0));
  and_gate and_gate_u_csamul_cla32_and18_29(.a(a[18]), .b(b[29]), .out(u_csamul_cla32_and18_29));
  fa fa_u_csamul_cla32_fa18_29_out(.a(u_csamul_cla32_and18_29[0]), .b(u_csamul_cla32_fa19_28_xor1[0]), .cin(u_csamul_cla32_fa18_28_or0[0]), .fa_xor1(u_csamul_cla32_fa18_29_xor1), .fa_or0(u_csamul_cla32_fa18_29_or0));
  and_gate and_gate_u_csamul_cla32_and19_29(.a(a[19]), .b(b[29]), .out(u_csamul_cla32_and19_29));
  fa fa_u_csamul_cla32_fa19_29_out(.a(u_csamul_cla32_and19_29[0]), .b(u_csamul_cla32_fa20_28_xor1[0]), .cin(u_csamul_cla32_fa19_28_or0[0]), .fa_xor1(u_csamul_cla32_fa19_29_xor1), .fa_or0(u_csamul_cla32_fa19_29_or0));
  and_gate and_gate_u_csamul_cla32_and20_29(.a(a[20]), .b(b[29]), .out(u_csamul_cla32_and20_29));
  fa fa_u_csamul_cla32_fa20_29_out(.a(u_csamul_cla32_and20_29[0]), .b(u_csamul_cla32_fa21_28_xor1[0]), .cin(u_csamul_cla32_fa20_28_or0[0]), .fa_xor1(u_csamul_cla32_fa20_29_xor1), .fa_or0(u_csamul_cla32_fa20_29_or0));
  and_gate and_gate_u_csamul_cla32_and21_29(.a(a[21]), .b(b[29]), .out(u_csamul_cla32_and21_29));
  fa fa_u_csamul_cla32_fa21_29_out(.a(u_csamul_cla32_and21_29[0]), .b(u_csamul_cla32_fa22_28_xor1[0]), .cin(u_csamul_cla32_fa21_28_or0[0]), .fa_xor1(u_csamul_cla32_fa21_29_xor1), .fa_or0(u_csamul_cla32_fa21_29_or0));
  and_gate and_gate_u_csamul_cla32_and22_29(.a(a[22]), .b(b[29]), .out(u_csamul_cla32_and22_29));
  fa fa_u_csamul_cla32_fa22_29_out(.a(u_csamul_cla32_and22_29[0]), .b(u_csamul_cla32_fa23_28_xor1[0]), .cin(u_csamul_cla32_fa22_28_or0[0]), .fa_xor1(u_csamul_cla32_fa22_29_xor1), .fa_or0(u_csamul_cla32_fa22_29_or0));
  and_gate and_gate_u_csamul_cla32_and23_29(.a(a[23]), .b(b[29]), .out(u_csamul_cla32_and23_29));
  fa fa_u_csamul_cla32_fa23_29_out(.a(u_csamul_cla32_and23_29[0]), .b(u_csamul_cla32_fa24_28_xor1[0]), .cin(u_csamul_cla32_fa23_28_or0[0]), .fa_xor1(u_csamul_cla32_fa23_29_xor1), .fa_or0(u_csamul_cla32_fa23_29_or0));
  and_gate and_gate_u_csamul_cla32_and24_29(.a(a[24]), .b(b[29]), .out(u_csamul_cla32_and24_29));
  fa fa_u_csamul_cla32_fa24_29_out(.a(u_csamul_cla32_and24_29[0]), .b(u_csamul_cla32_fa25_28_xor1[0]), .cin(u_csamul_cla32_fa24_28_or0[0]), .fa_xor1(u_csamul_cla32_fa24_29_xor1), .fa_or0(u_csamul_cla32_fa24_29_or0));
  and_gate and_gate_u_csamul_cla32_and25_29(.a(a[25]), .b(b[29]), .out(u_csamul_cla32_and25_29));
  fa fa_u_csamul_cla32_fa25_29_out(.a(u_csamul_cla32_and25_29[0]), .b(u_csamul_cla32_fa26_28_xor1[0]), .cin(u_csamul_cla32_fa25_28_or0[0]), .fa_xor1(u_csamul_cla32_fa25_29_xor1), .fa_or0(u_csamul_cla32_fa25_29_or0));
  and_gate and_gate_u_csamul_cla32_and26_29(.a(a[26]), .b(b[29]), .out(u_csamul_cla32_and26_29));
  fa fa_u_csamul_cla32_fa26_29_out(.a(u_csamul_cla32_and26_29[0]), .b(u_csamul_cla32_fa27_28_xor1[0]), .cin(u_csamul_cla32_fa26_28_or0[0]), .fa_xor1(u_csamul_cla32_fa26_29_xor1), .fa_or0(u_csamul_cla32_fa26_29_or0));
  and_gate and_gate_u_csamul_cla32_and27_29(.a(a[27]), .b(b[29]), .out(u_csamul_cla32_and27_29));
  fa fa_u_csamul_cla32_fa27_29_out(.a(u_csamul_cla32_and27_29[0]), .b(u_csamul_cla32_fa28_28_xor1[0]), .cin(u_csamul_cla32_fa27_28_or0[0]), .fa_xor1(u_csamul_cla32_fa27_29_xor1), .fa_or0(u_csamul_cla32_fa27_29_or0));
  and_gate and_gate_u_csamul_cla32_and28_29(.a(a[28]), .b(b[29]), .out(u_csamul_cla32_and28_29));
  fa fa_u_csamul_cla32_fa28_29_out(.a(u_csamul_cla32_and28_29[0]), .b(u_csamul_cla32_fa29_28_xor1[0]), .cin(u_csamul_cla32_fa28_28_or0[0]), .fa_xor1(u_csamul_cla32_fa28_29_xor1), .fa_or0(u_csamul_cla32_fa28_29_or0));
  and_gate and_gate_u_csamul_cla32_and29_29(.a(a[29]), .b(b[29]), .out(u_csamul_cla32_and29_29));
  fa fa_u_csamul_cla32_fa29_29_out(.a(u_csamul_cla32_and29_29[0]), .b(u_csamul_cla32_fa30_28_xor1[0]), .cin(u_csamul_cla32_fa29_28_or0[0]), .fa_xor1(u_csamul_cla32_fa29_29_xor1), .fa_or0(u_csamul_cla32_fa29_29_or0));
  and_gate and_gate_u_csamul_cla32_and30_29(.a(a[30]), .b(b[29]), .out(u_csamul_cla32_and30_29));
  fa fa_u_csamul_cla32_fa30_29_out(.a(u_csamul_cla32_and30_29[0]), .b(u_csamul_cla32_and31_28[0]), .cin(u_csamul_cla32_fa30_28_or0[0]), .fa_xor1(u_csamul_cla32_fa30_29_xor1), .fa_or0(u_csamul_cla32_fa30_29_or0));
  and_gate and_gate_u_csamul_cla32_and31_29(.a(a[31]), .b(b[29]), .out(u_csamul_cla32_and31_29));
  and_gate and_gate_u_csamul_cla32_and0_30(.a(a[0]), .b(b[30]), .out(u_csamul_cla32_and0_30));
  fa fa_u_csamul_cla32_fa0_30_out(.a(u_csamul_cla32_and0_30[0]), .b(u_csamul_cla32_fa1_29_xor1[0]), .cin(u_csamul_cla32_fa0_29_or0[0]), .fa_xor1(u_csamul_cla32_fa0_30_xor1), .fa_or0(u_csamul_cla32_fa0_30_or0));
  and_gate and_gate_u_csamul_cla32_and1_30(.a(a[1]), .b(b[30]), .out(u_csamul_cla32_and1_30));
  fa fa_u_csamul_cla32_fa1_30_out(.a(u_csamul_cla32_and1_30[0]), .b(u_csamul_cla32_fa2_29_xor1[0]), .cin(u_csamul_cla32_fa1_29_or0[0]), .fa_xor1(u_csamul_cla32_fa1_30_xor1), .fa_or0(u_csamul_cla32_fa1_30_or0));
  and_gate and_gate_u_csamul_cla32_and2_30(.a(a[2]), .b(b[30]), .out(u_csamul_cla32_and2_30));
  fa fa_u_csamul_cla32_fa2_30_out(.a(u_csamul_cla32_and2_30[0]), .b(u_csamul_cla32_fa3_29_xor1[0]), .cin(u_csamul_cla32_fa2_29_or0[0]), .fa_xor1(u_csamul_cla32_fa2_30_xor1), .fa_or0(u_csamul_cla32_fa2_30_or0));
  and_gate and_gate_u_csamul_cla32_and3_30(.a(a[3]), .b(b[30]), .out(u_csamul_cla32_and3_30));
  fa fa_u_csamul_cla32_fa3_30_out(.a(u_csamul_cla32_and3_30[0]), .b(u_csamul_cla32_fa4_29_xor1[0]), .cin(u_csamul_cla32_fa3_29_or0[0]), .fa_xor1(u_csamul_cla32_fa3_30_xor1), .fa_or0(u_csamul_cla32_fa3_30_or0));
  and_gate and_gate_u_csamul_cla32_and4_30(.a(a[4]), .b(b[30]), .out(u_csamul_cla32_and4_30));
  fa fa_u_csamul_cla32_fa4_30_out(.a(u_csamul_cla32_and4_30[0]), .b(u_csamul_cla32_fa5_29_xor1[0]), .cin(u_csamul_cla32_fa4_29_or0[0]), .fa_xor1(u_csamul_cla32_fa4_30_xor1), .fa_or0(u_csamul_cla32_fa4_30_or0));
  and_gate and_gate_u_csamul_cla32_and5_30(.a(a[5]), .b(b[30]), .out(u_csamul_cla32_and5_30));
  fa fa_u_csamul_cla32_fa5_30_out(.a(u_csamul_cla32_and5_30[0]), .b(u_csamul_cla32_fa6_29_xor1[0]), .cin(u_csamul_cla32_fa5_29_or0[0]), .fa_xor1(u_csamul_cla32_fa5_30_xor1), .fa_or0(u_csamul_cla32_fa5_30_or0));
  and_gate and_gate_u_csamul_cla32_and6_30(.a(a[6]), .b(b[30]), .out(u_csamul_cla32_and6_30));
  fa fa_u_csamul_cla32_fa6_30_out(.a(u_csamul_cla32_and6_30[0]), .b(u_csamul_cla32_fa7_29_xor1[0]), .cin(u_csamul_cla32_fa6_29_or0[0]), .fa_xor1(u_csamul_cla32_fa6_30_xor1), .fa_or0(u_csamul_cla32_fa6_30_or0));
  and_gate and_gate_u_csamul_cla32_and7_30(.a(a[7]), .b(b[30]), .out(u_csamul_cla32_and7_30));
  fa fa_u_csamul_cla32_fa7_30_out(.a(u_csamul_cla32_and7_30[0]), .b(u_csamul_cla32_fa8_29_xor1[0]), .cin(u_csamul_cla32_fa7_29_or0[0]), .fa_xor1(u_csamul_cla32_fa7_30_xor1), .fa_or0(u_csamul_cla32_fa7_30_or0));
  and_gate and_gate_u_csamul_cla32_and8_30(.a(a[8]), .b(b[30]), .out(u_csamul_cla32_and8_30));
  fa fa_u_csamul_cla32_fa8_30_out(.a(u_csamul_cla32_and8_30[0]), .b(u_csamul_cla32_fa9_29_xor1[0]), .cin(u_csamul_cla32_fa8_29_or0[0]), .fa_xor1(u_csamul_cla32_fa8_30_xor1), .fa_or0(u_csamul_cla32_fa8_30_or0));
  and_gate and_gate_u_csamul_cla32_and9_30(.a(a[9]), .b(b[30]), .out(u_csamul_cla32_and9_30));
  fa fa_u_csamul_cla32_fa9_30_out(.a(u_csamul_cla32_and9_30[0]), .b(u_csamul_cla32_fa10_29_xor1[0]), .cin(u_csamul_cla32_fa9_29_or0[0]), .fa_xor1(u_csamul_cla32_fa9_30_xor1), .fa_or0(u_csamul_cla32_fa9_30_or0));
  and_gate and_gate_u_csamul_cla32_and10_30(.a(a[10]), .b(b[30]), .out(u_csamul_cla32_and10_30));
  fa fa_u_csamul_cla32_fa10_30_out(.a(u_csamul_cla32_and10_30[0]), .b(u_csamul_cla32_fa11_29_xor1[0]), .cin(u_csamul_cla32_fa10_29_or0[0]), .fa_xor1(u_csamul_cla32_fa10_30_xor1), .fa_or0(u_csamul_cla32_fa10_30_or0));
  and_gate and_gate_u_csamul_cla32_and11_30(.a(a[11]), .b(b[30]), .out(u_csamul_cla32_and11_30));
  fa fa_u_csamul_cla32_fa11_30_out(.a(u_csamul_cla32_and11_30[0]), .b(u_csamul_cla32_fa12_29_xor1[0]), .cin(u_csamul_cla32_fa11_29_or0[0]), .fa_xor1(u_csamul_cla32_fa11_30_xor1), .fa_or0(u_csamul_cla32_fa11_30_or0));
  and_gate and_gate_u_csamul_cla32_and12_30(.a(a[12]), .b(b[30]), .out(u_csamul_cla32_and12_30));
  fa fa_u_csamul_cla32_fa12_30_out(.a(u_csamul_cla32_and12_30[0]), .b(u_csamul_cla32_fa13_29_xor1[0]), .cin(u_csamul_cla32_fa12_29_or0[0]), .fa_xor1(u_csamul_cla32_fa12_30_xor1), .fa_or0(u_csamul_cla32_fa12_30_or0));
  and_gate and_gate_u_csamul_cla32_and13_30(.a(a[13]), .b(b[30]), .out(u_csamul_cla32_and13_30));
  fa fa_u_csamul_cla32_fa13_30_out(.a(u_csamul_cla32_and13_30[0]), .b(u_csamul_cla32_fa14_29_xor1[0]), .cin(u_csamul_cla32_fa13_29_or0[0]), .fa_xor1(u_csamul_cla32_fa13_30_xor1), .fa_or0(u_csamul_cla32_fa13_30_or0));
  and_gate and_gate_u_csamul_cla32_and14_30(.a(a[14]), .b(b[30]), .out(u_csamul_cla32_and14_30));
  fa fa_u_csamul_cla32_fa14_30_out(.a(u_csamul_cla32_and14_30[0]), .b(u_csamul_cla32_fa15_29_xor1[0]), .cin(u_csamul_cla32_fa14_29_or0[0]), .fa_xor1(u_csamul_cla32_fa14_30_xor1), .fa_or0(u_csamul_cla32_fa14_30_or0));
  and_gate and_gate_u_csamul_cla32_and15_30(.a(a[15]), .b(b[30]), .out(u_csamul_cla32_and15_30));
  fa fa_u_csamul_cla32_fa15_30_out(.a(u_csamul_cla32_and15_30[0]), .b(u_csamul_cla32_fa16_29_xor1[0]), .cin(u_csamul_cla32_fa15_29_or0[0]), .fa_xor1(u_csamul_cla32_fa15_30_xor1), .fa_or0(u_csamul_cla32_fa15_30_or0));
  and_gate and_gate_u_csamul_cla32_and16_30(.a(a[16]), .b(b[30]), .out(u_csamul_cla32_and16_30));
  fa fa_u_csamul_cla32_fa16_30_out(.a(u_csamul_cla32_and16_30[0]), .b(u_csamul_cla32_fa17_29_xor1[0]), .cin(u_csamul_cla32_fa16_29_or0[0]), .fa_xor1(u_csamul_cla32_fa16_30_xor1), .fa_or0(u_csamul_cla32_fa16_30_or0));
  and_gate and_gate_u_csamul_cla32_and17_30(.a(a[17]), .b(b[30]), .out(u_csamul_cla32_and17_30));
  fa fa_u_csamul_cla32_fa17_30_out(.a(u_csamul_cla32_and17_30[0]), .b(u_csamul_cla32_fa18_29_xor1[0]), .cin(u_csamul_cla32_fa17_29_or0[0]), .fa_xor1(u_csamul_cla32_fa17_30_xor1), .fa_or0(u_csamul_cla32_fa17_30_or0));
  and_gate and_gate_u_csamul_cla32_and18_30(.a(a[18]), .b(b[30]), .out(u_csamul_cla32_and18_30));
  fa fa_u_csamul_cla32_fa18_30_out(.a(u_csamul_cla32_and18_30[0]), .b(u_csamul_cla32_fa19_29_xor1[0]), .cin(u_csamul_cla32_fa18_29_or0[0]), .fa_xor1(u_csamul_cla32_fa18_30_xor1), .fa_or0(u_csamul_cla32_fa18_30_or0));
  and_gate and_gate_u_csamul_cla32_and19_30(.a(a[19]), .b(b[30]), .out(u_csamul_cla32_and19_30));
  fa fa_u_csamul_cla32_fa19_30_out(.a(u_csamul_cla32_and19_30[0]), .b(u_csamul_cla32_fa20_29_xor1[0]), .cin(u_csamul_cla32_fa19_29_or0[0]), .fa_xor1(u_csamul_cla32_fa19_30_xor1), .fa_or0(u_csamul_cla32_fa19_30_or0));
  and_gate and_gate_u_csamul_cla32_and20_30(.a(a[20]), .b(b[30]), .out(u_csamul_cla32_and20_30));
  fa fa_u_csamul_cla32_fa20_30_out(.a(u_csamul_cla32_and20_30[0]), .b(u_csamul_cla32_fa21_29_xor1[0]), .cin(u_csamul_cla32_fa20_29_or0[0]), .fa_xor1(u_csamul_cla32_fa20_30_xor1), .fa_or0(u_csamul_cla32_fa20_30_or0));
  and_gate and_gate_u_csamul_cla32_and21_30(.a(a[21]), .b(b[30]), .out(u_csamul_cla32_and21_30));
  fa fa_u_csamul_cla32_fa21_30_out(.a(u_csamul_cla32_and21_30[0]), .b(u_csamul_cla32_fa22_29_xor1[0]), .cin(u_csamul_cla32_fa21_29_or0[0]), .fa_xor1(u_csamul_cla32_fa21_30_xor1), .fa_or0(u_csamul_cla32_fa21_30_or0));
  and_gate and_gate_u_csamul_cla32_and22_30(.a(a[22]), .b(b[30]), .out(u_csamul_cla32_and22_30));
  fa fa_u_csamul_cla32_fa22_30_out(.a(u_csamul_cla32_and22_30[0]), .b(u_csamul_cla32_fa23_29_xor1[0]), .cin(u_csamul_cla32_fa22_29_or0[0]), .fa_xor1(u_csamul_cla32_fa22_30_xor1), .fa_or0(u_csamul_cla32_fa22_30_or0));
  and_gate and_gate_u_csamul_cla32_and23_30(.a(a[23]), .b(b[30]), .out(u_csamul_cla32_and23_30));
  fa fa_u_csamul_cla32_fa23_30_out(.a(u_csamul_cla32_and23_30[0]), .b(u_csamul_cla32_fa24_29_xor1[0]), .cin(u_csamul_cla32_fa23_29_or0[0]), .fa_xor1(u_csamul_cla32_fa23_30_xor1), .fa_or0(u_csamul_cla32_fa23_30_or0));
  and_gate and_gate_u_csamul_cla32_and24_30(.a(a[24]), .b(b[30]), .out(u_csamul_cla32_and24_30));
  fa fa_u_csamul_cla32_fa24_30_out(.a(u_csamul_cla32_and24_30[0]), .b(u_csamul_cla32_fa25_29_xor1[0]), .cin(u_csamul_cla32_fa24_29_or0[0]), .fa_xor1(u_csamul_cla32_fa24_30_xor1), .fa_or0(u_csamul_cla32_fa24_30_or0));
  and_gate and_gate_u_csamul_cla32_and25_30(.a(a[25]), .b(b[30]), .out(u_csamul_cla32_and25_30));
  fa fa_u_csamul_cla32_fa25_30_out(.a(u_csamul_cla32_and25_30[0]), .b(u_csamul_cla32_fa26_29_xor1[0]), .cin(u_csamul_cla32_fa25_29_or0[0]), .fa_xor1(u_csamul_cla32_fa25_30_xor1), .fa_or0(u_csamul_cla32_fa25_30_or0));
  and_gate and_gate_u_csamul_cla32_and26_30(.a(a[26]), .b(b[30]), .out(u_csamul_cla32_and26_30));
  fa fa_u_csamul_cla32_fa26_30_out(.a(u_csamul_cla32_and26_30[0]), .b(u_csamul_cla32_fa27_29_xor1[0]), .cin(u_csamul_cla32_fa26_29_or0[0]), .fa_xor1(u_csamul_cla32_fa26_30_xor1), .fa_or0(u_csamul_cla32_fa26_30_or0));
  and_gate and_gate_u_csamul_cla32_and27_30(.a(a[27]), .b(b[30]), .out(u_csamul_cla32_and27_30));
  fa fa_u_csamul_cla32_fa27_30_out(.a(u_csamul_cla32_and27_30[0]), .b(u_csamul_cla32_fa28_29_xor1[0]), .cin(u_csamul_cla32_fa27_29_or0[0]), .fa_xor1(u_csamul_cla32_fa27_30_xor1), .fa_or0(u_csamul_cla32_fa27_30_or0));
  and_gate and_gate_u_csamul_cla32_and28_30(.a(a[28]), .b(b[30]), .out(u_csamul_cla32_and28_30));
  fa fa_u_csamul_cla32_fa28_30_out(.a(u_csamul_cla32_and28_30[0]), .b(u_csamul_cla32_fa29_29_xor1[0]), .cin(u_csamul_cla32_fa28_29_or0[0]), .fa_xor1(u_csamul_cla32_fa28_30_xor1), .fa_or0(u_csamul_cla32_fa28_30_or0));
  and_gate and_gate_u_csamul_cla32_and29_30(.a(a[29]), .b(b[30]), .out(u_csamul_cla32_and29_30));
  fa fa_u_csamul_cla32_fa29_30_out(.a(u_csamul_cla32_and29_30[0]), .b(u_csamul_cla32_fa30_29_xor1[0]), .cin(u_csamul_cla32_fa29_29_or0[0]), .fa_xor1(u_csamul_cla32_fa29_30_xor1), .fa_or0(u_csamul_cla32_fa29_30_or0));
  and_gate and_gate_u_csamul_cla32_and30_30(.a(a[30]), .b(b[30]), .out(u_csamul_cla32_and30_30));
  fa fa_u_csamul_cla32_fa30_30_out(.a(u_csamul_cla32_and30_30[0]), .b(u_csamul_cla32_and31_29[0]), .cin(u_csamul_cla32_fa30_29_or0[0]), .fa_xor1(u_csamul_cla32_fa30_30_xor1), .fa_or0(u_csamul_cla32_fa30_30_or0));
  and_gate and_gate_u_csamul_cla32_and31_30(.a(a[31]), .b(b[30]), .out(u_csamul_cla32_and31_30));
  and_gate and_gate_u_csamul_cla32_and0_31(.a(a[0]), .b(b[31]), .out(u_csamul_cla32_and0_31));
  fa fa_u_csamul_cla32_fa0_31_out(.a(u_csamul_cla32_and0_31[0]), .b(u_csamul_cla32_fa1_30_xor1[0]), .cin(u_csamul_cla32_fa0_30_or0[0]), .fa_xor1(u_csamul_cla32_fa0_31_xor1), .fa_or0(u_csamul_cla32_fa0_31_or0));
  and_gate and_gate_u_csamul_cla32_and1_31(.a(a[1]), .b(b[31]), .out(u_csamul_cla32_and1_31));
  fa fa_u_csamul_cla32_fa1_31_out(.a(u_csamul_cla32_and1_31[0]), .b(u_csamul_cla32_fa2_30_xor1[0]), .cin(u_csamul_cla32_fa1_30_or0[0]), .fa_xor1(u_csamul_cla32_fa1_31_xor1), .fa_or0(u_csamul_cla32_fa1_31_or0));
  and_gate and_gate_u_csamul_cla32_and2_31(.a(a[2]), .b(b[31]), .out(u_csamul_cla32_and2_31));
  fa fa_u_csamul_cla32_fa2_31_out(.a(u_csamul_cla32_and2_31[0]), .b(u_csamul_cla32_fa3_30_xor1[0]), .cin(u_csamul_cla32_fa2_30_or0[0]), .fa_xor1(u_csamul_cla32_fa2_31_xor1), .fa_or0(u_csamul_cla32_fa2_31_or0));
  and_gate and_gate_u_csamul_cla32_and3_31(.a(a[3]), .b(b[31]), .out(u_csamul_cla32_and3_31));
  fa fa_u_csamul_cla32_fa3_31_out(.a(u_csamul_cla32_and3_31[0]), .b(u_csamul_cla32_fa4_30_xor1[0]), .cin(u_csamul_cla32_fa3_30_or0[0]), .fa_xor1(u_csamul_cla32_fa3_31_xor1), .fa_or0(u_csamul_cla32_fa3_31_or0));
  and_gate and_gate_u_csamul_cla32_and4_31(.a(a[4]), .b(b[31]), .out(u_csamul_cla32_and4_31));
  fa fa_u_csamul_cla32_fa4_31_out(.a(u_csamul_cla32_and4_31[0]), .b(u_csamul_cla32_fa5_30_xor1[0]), .cin(u_csamul_cla32_fa4_30_or0[0]), .fa_xor1(u_csamul_cla32_fa4_31_xor1), .fa_or0(u_csamul_cla32_fa4_31_or0));
  and_gate and_gate_u_csamul_cla32_and5_31(.a(a[5]), .b(b[31]), .out(u_csamul_cla32_and5_31));
  fa fa_u_csamul_cla32_fa5_31_out(.a(u_csamul_cla32_and5_31[0]), .b(u_csamul_cla32_fa6_30_xor1[0]), .cin(u_csamul_cla32_fa5_30_or0[0]), .fa_xor1(u_csamul_cla32_fa5_31_xor1), .fa_or0(u_csamul_cla32_fa5_31_or0));
  and_gate and_gate_u_csamul_cla32_and6_31(.a(a[6]), .b(b[31]), .out(u_csamul_cla32_and6_31));
  fa fa_u_csamul_cla32_fa6_31_out(.a(u_csamul_cla32_and6_31[0]), .b(u_csamul_cla32_fa7_30_xor1[0]), .cin(u_csamul_cla32_fa6_30_or0[0]), .fa_xor1(u_csamul_cla32_fa6_31_xor1), .fa_or0(u_csamul_cla32_fa6_31_or0));
  and_gate and_gate_u_csamul_cla32_and7_31(.a(a[7]), .b(b[31]), .out(u_csamul_cla32_and7_31));
  fa fa_u_csamul_cla32_fa7_31_out(.a(u_csamul_cla32_and7_31[0]), .b(u_csamul_cla32_fa8_30_xor1[0]), .cin(u_csamul_cla32_fa7_30_or0[0]), .fa_xor1(u_csamul_cla32_fa7_31_xor1), .fa_or0(u_csamul_cla32_fa7_31_or0));
  and_gate and_gate_u_csamul_cla32_and8_31(.a(a[8]), .b(b[31]), .out(u_csamul_cla32_and8_31));
  fa fa_u_csamul_cla32_fa8_31_out(.a(u_csamul_cla32_and8_31[0]), .b(u_csamul_cla32_fa9_30_xor1[0]), .cin(u_csamul_cla32_fa8_30_or0[0]), .fa_xor1(u_csamul_cla32_fa8_31_xor1), .fa_or0(u_csamul_cla32_fa8_31_or0));
  and_gate and_gate_u_csamul_cla32_and9_31(.a(a[9]), .b(b[31]), .out(u_csamul_cla32_and9_31));
  fa fa_u_csamul_cla32_fa9_31_out(.a(u_csamul_cla32_and9_31[0]), .b(u_csamul_cla32_fa10_30_xor1[0]), .cin(u_csamul_cla32_fa9_30_or0[0]), .fa_xor1(u_csamul_cla32_fa9_31_xor1), .fa_or0(u_csamul_cla32_fa9_31_or0));
  and_gate and_gate_u_csamul_cla32_and10_31(.a(a[10]), .b(b[31]), .out(u_csamul_cla32_and10_31));
  fa fa_u_csamul_cla32_fa10_31_out(.a(u_csamul_cla32_and10_31[0]), .b(u_csamul_cla32_fa11_30_xor1[0]), .cin(u_csamul_cla32_fa10_30_or0[0]), .fa_xor1(u_csamul_cla32_fa10_31_xor1), .fa_or0(u_csamul_cla32_fa10_31_or0));
  and_gate and_gate_u_csamul_cla32_and11_31(.a(a[11]), .b(b[31]), .out(u_csamul_cla32_and11_31));
  fa fa_u_csamul_cla32_fa11_31_out(.a(u_csamul_cla32_and11_31[0]), .b(u_csamul_cla32_fa12_30_xor1[0]), .cin(u_csamul_cla32_fa11_30_or0[0]), .fa_xor1(u_csamul_cla32_fa11_31_xor1), .fa_or0(u_csamul_cla32_fa11_31_or0));
  and_gate and_gate_u_csamul_cla32_and12_31(.a(a[12]), .b(b[31]), .out(u_csamul_cla32_and12_31));
  fa fa_u_csamul_cla32_fa12_31_out(.a(u_csamul_cla32_and12_31[0]), .b(u_csamul_cla32_fa13_30_xor1[0]), .cin(u_csamul_cla32_fa12_30_or0[0]), .fa_xor1(u_csamul_cla32_fa12_31_xor1), .fa_or0(u_csamul_cla32_fa12_31_or0));
  and_gate and_gate_u_csamul_cla32_and13_31(.a(a[13]), .b(b[31]), .out(u_csamul_cla32_and13_31));
  fa fa_u_csamul_cla32_fa13_31_out(.a(u_csamul_cla32_and13_31[0]), .b(u_csamul_cla32_fa14_30_xor1[0]), .cin(u_csamul_cla32_fa13_30_or0[0]), .fa_xor1(u_csamul_cla32_fa13_31_xor1), .fa_or0(u_csamul_cla32_fa13_31_or0));
  and_gate and_gate_u_csamul_cla32_and14_31(.a(a[14]), .b(b[31]), .out(u_csamul_cla32_and14_31));
  fa fa_u_csamul_cla32_fa14_31_out(.a(u_csamul_cla32_and14_31[0]), .b(u_csamul_cla32_fa15_30_xor1[0]), .cin(u_csamul_cla32_fa14_30_or0[0]), .fa_xor1(u_csamul_cla32_fa14_31_xor1), .fa_or0(u_csamul_cla32_fa14_31_or0));
  and_gate and_gate_u_csamul_cla32_and15_31(.a(a[15]), .b(b[31]), .out(u_csamul_cla32_and15_31));
  fa fa_u_csamul_cla32_fa15_31_out(.a(u_csamul_cla32_and15_31[0]), .b(u_csamul_cla32_fa16_30_xor1[0]), .cin(u_csamul_cla32_fa15_30_or0[0]), .fa_xor1(u_csamul_cla32_fa15_31_xor1), .fa_or0(u_csamul_cla32_fa15_31_or0));
  and_gate and_gate_u_csamul_cla32_and16_31(.a(a[16]), .b(b[31]), .out(u_csamul_cla32_and16_31));
  fa fa_u_csamul_cla32_fa16_31_out(.a(u_csamul_cla32_and16_31[0]), .b(u_csamul_cla32_fa17_30_xor1[0]), .cin(u_csamul_cla32_fa16_30_or0[0]), .fa_xor1(u_csamul_cla32_fa16_31_xor1), .fa_or0(u_csamul_cla32_fa16_31_or0));
  and_gate and_gate_u_csamul_cla32_and17_31(.a(a[17]), .b(b[31]), .out(u_csamul_cla32_and17_31));
  fa fa_u_csamul_cla32_fa17_31_out(.a(u_csamul_cla32_and17_31[0]), .b(u_csamul_cla32_fa18_30_xor1[0]), .cin(u_csamul_cla32_fa17_30_or0[0]), .fa_xor1(u_csamul_cla32_fa17_31_xor1), .fa_or0(u_csamul_cla32_fa17_31_or0));
  and_gate and_gate_u_csamul_cla32_and18_31(.a(a[18]), .b(b[31]), .out(u_csamul_cla32_and18_31));
  fa fa_u_csamul_cla32_fa18_31_out(.a(u_csamul_cla32_and18_31[0]), .b(u_csamul_cla32_fa19_30_xor1[0]), .cin(u_csamul_cla32_fa18_30_or0[0]), .fa_xor1(u_csamul_cla32_fa18_31_xor1), .fa_or0(u_csamul_cla32_fa18_31_or0));
  and_gate and_gate_u_csamul_cla32_and19_31(.a(a[19]), .b(b[31]), .out(u_csamul_cla32_and19_31));
  fa fa_u_csamul_cla32_fa19_31_out(.a(u_csamul_cla32_and19_31[0]), .b(u_csamul_cla32_fa20_30_xor1[0]), .cin(u_csamul_cla32_fa19_30_or0[0]), .fa_xor1(u_csamul_cla32_fa19_31_xor1), .fa_or0(u_csamul_cla32_fa19_31_or0));
  and_gate and_gate_u_csamul_cla32_and20_31(.a(a[20]), .b(b[31]), .out(u_csamul_cla32_and20_31));
  fa fa_u_csamul_cla32_fa20_31_out(.a(u_csamul_cla32_and20_31[0]), .b(u_csamul_cla32_fa21_30_xor1[0]), .cin(u_csamul_cla32_fa20_30_or0[0]), .fa_xor1(u_csamul_cla32_fa20_31_xor1), .fa_or0(u_csamul_cla32_fa20_31_or0));
  and_gate and_gate_u_csamul_cla32_and21_31(.a(a[21]), .b(b[31]), .out(u_csamul_cla32_and21_31));
  fa fa_u_csamul_cla32_fa21_31_out(.a(u_csamul_cla32_and21_31[0]), .b(u_csamul_cla32_fa22_30_xor1[0]), .cin(u_csamul_cla32_fa21_30_or0[0]), .fa_xor1(u_csamul_cla32_fa21_31_xor1), .fa_or0(u_csamul_cla32_fa21_31_or0));
  and_gate and_gate_u_csamul_cla32_and22_31(.a(a[22]), .b(b[31]), .out(u_csamul_cla32_and22_31));
  fa fa_u_csamul_cla32_fa22_31_out(.a(u_csamul_cla32_and22_31[0]), .b(u_csamul_cla32_fa23_30_xor1[0]), .cin(u_csamul_cla32_fa22_30_or0[0]), .fa_xor1(u_csamul_cla32_fa22_31_xor1), .fa_or0(u_csamul_cla32_fa22_31_or0));
  and_gate and_gate_u_csamul_cla32_and23_31(.a(a[23]), .b(b[31]), .out(u_csamul_cla32_and23_31));
  fa fa_u_csamul_cla32_fa23_31_out(.a(u_csamul_cla32_and23_31[0]), .b(u_csamul_cla32_fa24_30_xor1[0]), .cin(u_csamul_cla32_fa23_30_or0[0]), .fa_xor1(u_csamul_cla32_fa23_31_xor1), .fa_or0(u_csamul_cla32_fa23_31_or0));
  and_gate and_gate_u_csamul_cla32_and24_31(.a(a[24]), .b(b[31]), .out(u_csamul_cla32_and24_31));
  fa fa_u_csamul_cla32_fa24_31_out(.a(u_csamul_cla32_and24_31[0]), .b(u_csamul_cla32_fa25_30_xor1[0]), .cin(u_csamul_cla32_fa24_30_or0[0]), .fa_xor1(u_csamul_cla32_fa24_31_xor1), .fa_or0(u_csamul_cla32_fa24_31_or0));
  and_gate and_gate_u_csamul_cla32_and25_31(.a(a[25]), .b(b[31]), .out(u_csamul_cla32_and25_31));
  fa fa_u_csamul_cla32_fa25_31_out(.a(u_csamul_cla32_and25_31[0]), .b(u_csamul_cla32_fa26_30_xor1[0]), .cin(u_csamul_cla32_fa25_30_or0[0]), .fa_xor1(u_csamul_cla32_fa25_31_xor1), .fa_or0(u_csamul_cla32_fa25_31_or0));
  and_gate and_gate_u_csamul_cla32_and26_31(.a(a[26]), .b(b[31]), .out(u_csamul_cla32_and26_31));
  fa fa_u_csamul_cla32_fa26_31_out(.a(u_csamul_cla32_and26_31[0]), .b(u_csamul_cla32_fa27_30_xor1[0]), .cin(u_csamul_cla32_fa26_30_or0[0]), .fa_xor1(u_csamul_cla32_fa26_31_xor1), .fa_or0(u_csamul_cla32_fa26_31_or0));
  and_gate and_gate_u_csamul_cla32_and27_31(.a(a[27]), .b(b[31]), .out(u_csamul_cla32_and27_31));
  fa fa_u_csamul_cla32_fa27_31_out(.a(u_csamul_cla32_and27_31[0]), .b(u_csamul_cla32_fa28_30_xor1[0]), .cin(u_csamul_cla32_fa27_30_or0[0]), .fa_xor1(u_csamul_cla32_fa27_31_xor1), .fa_or0(u_csamul_cla32_fa27_31_or0));
  and_gate and_gate_u_csamul_cla32_and28_31(.a(a[28]), .b(b[31]), .out(u_csamul_cla32_and28_31));
  fa fa_u_csamul_cla32_fa28_31_out(.a(u_csamul_cla32_and28_31[0]), .b(u_csamul_cla32_fa29_30_xor1[0]), .cin(u_csamul_cla32_fa28_30_or0[0]), .fa_xor1(u_csamul_cla32_fa28_31_xor1), .fa_or0(u_csamul_cla32_fa28_31_or0));
  and_gate and_gate_u_csamul_cla32_and29_31(.a(a[29]), .b(b[31]), .out(u_csamul_cla32_and29_31));
  fa fa_u_csamul_cla32_fa29_31_out(.a(u_csamul_cla32_and29_31[0]), .b(u_csamul_cla32_fa30_30_xor1[0]), .cin(u_csamul_cla32_fa29_30_or0[0]), .fa_xor1(u_csamul_cla32_fa29_31_xor1), .fa_or0(u_csamul_cla32_fa29_31_or0));
  and_gate and_gate_u_csamul_cla32_and30_31(.a(a[30]), .b(b[31]), .out(u_csamul_cla32_and30_31));
  fa fa_u_csamul_cla32_fa30_31_out(.a(u_csamul_cla32_and30_31[0]), .b(u_csamul_cla32_and31_30[0]), .cin(u_csamul_cla32_fa30_30_or0[0]), .fa_xor1(u_csamul_cla32_fa30_31_xor1), .fa_or0(u_csamul_cla32_fa30_31_or0));
  and_gate and_gate_u_csamul_cla32_and31_31(.a(a[31]), .b(b[31]), .out(u_csamul_cla32_and31_31));
  assign u_csamul_cla32_u_cla32_a[0] = u_csamul_cla32_fa1_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[1] = u_csamul_cla32_fa2_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[2] = u_csamul_cla32_fa3_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[3] = u_csamul_cla32_fa4_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[4] = u_csamul_cla32_fa5_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[5] = u_csamul_cla32_fa6_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[6] = u_csamul_cla32_fa7_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[7] = u_csamul_cla32_fa8_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[8] = u_csamul_cla32_fa9_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[9] = u_csamul_cla32_fa10_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[10] = u_csamul_cla32_fa11_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[11] = u_csamul_cla32_fa12_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[12] = u_csamul_cla32_fa13_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[13] = u_csamul_cla32_fa14_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[14] = u_csamul_cla32_fa15_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[15] = u_csamul_cla32_fa16_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[16] = u_csamul_cla32_fa17_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[17] = u_csamul_cla32_fa18_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[18] = u_csamul_cla32_fa19_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[19] = u_csamul_cla32_fa20_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[20] = u_csamul_cla32_fa21_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[21] = u_csamul_cla32_fa22_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[22] = u_csamul_cla32_fa23_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[23] = u_csamul_cla32_fa24_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[24] = u_csamul_cla32_fa25_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[25] = u_csamul_cla32_fa26_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[26] = u_csamul_cla32_fa27_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[27] = u_csamul_cla32_fa28_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[28] = u_csamul_cla32_fa29_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[29] = u_csamul_cla32_fa30_31_xor1[0];
  assign u_csamul_cla32_u_cla32_a[30] = u_csamul_cla32_and31_31[0];
  assign u_csamul_cla32_u_cla32_a[31] = 1'b0;
  assign u_csamul_cla32_u_cla32_b[0] = u_csamul_cla32_fa0_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[1] = u_csamul_cla32_fa1_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[2] = u_csamul_cla32_fa2_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[3] = u_csamul_cla32_fa3_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[4] = u_csamul_cla32_fa4_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[5] = u_csamul_cla32_fa5_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[6] = u_csamul_cla32_fa6_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[7] = u_csamul_cla32_fa7_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[8] = u_csamul_cla32_fa8_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[9] = u_csamul_cla32_fa9_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[10] = u_csamul_cla32_fa10_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[11] = u_csamul_cla32_fa11_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[12] = u_csamul_cla32_fa12_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[13] = u_csamul_cla32_fa13_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[14] = u_csamul_cla32_fa14_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[15] = u_csamul_cla32_fa15_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[16] = u_csamul_cla32_fa16_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[17] = u_csamul_cla32_fa17_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[18] = u_csamul_cla32_fa18_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[19] = u_csamul_cla32_fa19_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[20] = u_csamul_cla32_fa20_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[21] = u_csamul_cla32_fa21_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[22] = u_csamul_cla32_fa22_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[23] = u_csamul_cla32_fa23_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[24] = u_csamul_cla32_fa24_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[25] = u_csamul_cla32_fa25_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[26] = u_csamul_cla32_fa26_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[27] = u_csamul_cla32_fa27_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[28] = u_csamul_cla32_fa28_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[29] = u_csamul_cla32_fa29_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[30] = u_csamul_cla32_fa30_31_or0[0];
  assign u_csamul_cla32_u_cla32_b[31] = 1'b0;
  u_cla32 u_cla32_u_csamul_cla32_u_cla32_out(.a(u_csamul_cla32_u_cla32_a), .b(u_csamul_cla32_u_cla32_b), .u_cla32_out(u_csamul_cla32_u_cla32_out));

  assign u_csamul_cla32_out[0] = u_csamul_cla32_and0_0[0];
  assign u_csamul_cla32_out[1] = u_csamul_cla32_ha0_1_xor0[0];
  assign u_csamul_cla32_out[2] = u_csamul_cla32_fa0_2_xor1[0];
  assign u_csamul_cla32_out[3] = u_csamul_cla32_fa0_3_xor1[0];
  assign u_csamul_cla32_out[4] = u_csamul_cla32_fa0_4_xor1[0];
  assign u_csamul_cla32_out[5] = u_csamul_cla32_fa0_5_xor1[0];
  assign u_csamul_cla32_out[6] = u_csamul_cla32_fa0_6_xor1[0];
  assign u_csamul_cla32_out[7] = u_csamul_cla32_fa0_7_xor1[0];
  assign u_csamul_cla32_out[8] = u_csamul_cla32_fa0_8_xor1[0];
  assign u_csamul_cla32_out[9] = u_csamul_cla32_fa0_9_xor1[0];
  assign u_csamul_cla32_out[10] = u_csamul_cla32_fa0_10_xor1[0];
  assign u_csamul_cla32_out[11] = u_csamul_cla32_fa0_11_xor1[0];
  assign u_csamul_cla32_out[12] = u_csamul_cla32_fa0_12_xor1[0];
  assign u_csamul_cla32_out[13] = u_csamul_cla32_fa0_13_xor1[0];
  assign u_csamul_cla32_out[14] = u_csamul_cla32_fa0_14_xor1[0];
  assign u_csamul_cla32_out[15] = u_csamul_cla32_fa0_15_xor1[0];
  assign u_csamul_cla32_out[16] = u_csamul_cla32_fa0_16_xor1[0];
  assign u_csamul_cla32_out[17] = u_csamul_cla32_fa0_17_xor1[0];
  assign u_csamul_cla32_out[18] = u_csamul_cla32_fa0_18_xor1[0];
  assign u_csamul_cla32_out[19] = u_csamul_cla32_fa0_19_xor1[0];
  assign u_csamul_cla32_out[20] = u_csamul_cla32_fa0_20_xor1[0];
  assign u_csamul_cla32_out[21] = u_csamul_cla32_fa0_21_xor1[0];
  assign u_csamul_cla32_out[22] = u_csamul_cla32_fa0_22_xor1[0];
  assign u_csamul_cla32_out[23] = u_csamul_cla32_fa0_23_xor1[0];
  assign u_csamul_cla32_out[24] = u_csamul_cla32_fa0_24_xor1[0];
  assign u_csamul_cla32_out[25] = u_csamul_cla32_fa0_25_xor1[0];
  assign u_csamul_cla32_out[26] = u_csamul_cla32_fa0_26_xor1[0];
  assign u_csamul_cla32_out[27] = u_csamul_cla32_fa0_27_xor1[0];
  assign u_csamul_cla32_out[28] = u_csamul_cla32_fa0_28_xor1[0];
  assign u_csamul_cla32_out[29] = u_csamul_cla32_fa0_29_xor1[0];
  assign u_csamul_cla32_out[30] = u_csamul_cla32_fa0_30_xor1[0];
  assign u_csamul_cla32_out[31] = u_csamul_cla32_fa0_31_xor1[0];
  assign u_csamul_cla32_out[32] = u_csamul_cla32_u_cla32_out[0];
  assign u_csamul_cla32_out[33] = u_csamul_cla32_u_cla32_out[1];
  assign u_csamul_cla32_out[34] = u_csamul_cla32_u_cla32_out[2];
  assign u_csamul_cla32_out[35] = u_csamul_cla32_u_cla32_out[3];
  assign u_csamul_cla32_out[36] = u_csamul_cla32_u_cla32_out[4];
  assign u_csamul_cla32_out[37] = u_csamul_cla32_u_cla32_out[5];
  assign u_csamul_cla32_out[38] = u_csamul_cla32_u_cla32_out[6];
  assign u_csamul_cla32_out[39] = u_csamul_cla32_u_cla32_out[7];
  assign u_csamul_cla32_out[40] = u_csamul_cla32_u_cla32_out[8];
  assign u_csamul_cla32_out[41] = u_csamul_cla32_u_cla32_out[9];
  assign u_csamul_cla32_out[42] = u_csamul_cla32_u_cla32_out[10];
  assign u_csamul_cla32_out[43] = u_csamul_cla32_u_cla32_out[11];
  assign u_csamul_cla32_out[44] = u_csamul_cla32_u_cla32_out[12];
  assign u_csamul_cla32_out[45] = u_csamul_cla32_u_cla32_out[13];
  assign u_csamul_cla32_out[46] = u_csamul_cla32_u_cla32_out[14];
  assign u_csamul_cla32_out[47] = u_csamul_cla32_u_cla32_out[15];
  assign u_csamul_cla32_out[48] = u_csamul_cla32_u_cla32_out[16];
  assign u_csamul_cla32_out[49] = u_csamul_cla32_u_cla32_out[17];
  assign u_csamul_cla32_out[50] = u_csamul_cla32_u_cla32_out[18];
  assign u_csamul_cla32_out[51] = u_csamul_cla32_u_cla32_out[19];
  assign u_csamul_cla32_out[52] = u_csamul_cla32_u_cla32_out[20];
  assign u_csamul_cla32_out[53] = u_csamul_cla32_u_cla32_out[21];
  assign u_csamul_cla32_out[54] = u_csamul_cla32_u_cla32_out[22];
  assign u_csamul_cla32_out[55] = u_csamul_cla32_u_cla32_out[23];
  assign u_csamul_cla32_out[56] = u_csamul_cla32_u_cla32_out[24];
  assign u_csamul_cla32_out[57] = u_csamul_cla32_u_cla32_out[25];
  assign u_csamul_cla32_out[58] = u_csamul_cla32_u_cla32_out[26];
  assign u_csamul_cla32_out[59] = u_csamul_cla32_u_cla32_out[27];
  assign u_csamul_cla32_out[60] = u_csamul_cla32_u_cla32_out[28];
  assign u_csamul_cla32_out[61] = u_csamul_cla32_u_cla32_out[29];
  assign u_csamul_cla32_out[62] = u_csamul_cla32_u_cla32_out[30];
  assign u_csamul_cla32_out[63] = u_csamul_cla32_u_cla32_out[31];
endmodule