module f_u_cska12(input [11:0] a, input [11:0] b, output [12:0] f_u_cska12_out);
  wire f_u_cska12_xor0;
  wire f_u_cska12_ha0_xor0;
  wire f_u_cska12_ha0_and0;
  wire f_u_cska12_xor1;
  wire f_u_cska12_fa0_xor0;
  wire f_u_cska12_fa0_and0;
  wire f_u_cska12_fa0_xor1;
  wire f_u_cska12_fa0_and1;
  wire f_u_cska12_fa0_or0;
  wire f_u_cska12_xor2;
  wire f_u_cska12_fa1_xor0;
  wire f_u_cska12_fa1_and0;
  wire f_u_cska12_fa1_xor1;
  wire f_u_cska12_fa1_and1;
  wire f_u_cska12_fa1_or0;
  wire f_u_cska12_xor3;
  wire f_u_cska12_fa2_xor0;
  wire f_u_cska12_fa2_and0;
  wire f_u_cska12_fa2_xor1;
  wire f_u_cska12_fa2_and1;
  wire f_u_cska12_fa2_or0;
  wire f_u_cska12_and_propagate00;
  wire f_u_cska12_and_propagate01;
  wire f_u_cska12_and_propagate02;
  wire f_u_cska12_mux2to10_not0;
  wire f_u_cska12_mux2to10_and1;
  wire f_u_cska12_xor4;
  wire f_u_cska12_fa3_xor0;
  wire f_u_cska12_fa3_and0;
  wire f_u_cska12_fa3_xor1;
  wire f_u_cska12_fa3_and1;
  wire f_u_cska12_fa3_or0;
  wire f_u_cska12_xor5;
  wire f_u_cska12_fa4_xor0;
  wire f_u_cska12_fa4_and0;
  wire f_u_cska12_fa4_xor1;
  wire f_u_cska12_fa4_and1;
  wire f_u_cska12_fa4_or0;
  wire f_u_cska12_xor6;
  wire f_u_cska12_fa5_xor0;
  wire f_u_cska12_fa5_and0;
  wire f_u_cska12_fa5_xor1;
  wire f_u_cska12_fa5_and1;
  wire f_u_cska12_fa5_or0;
  wire f_u_cska12_xor7;
  wire f_u_cska12_fa6_xor0;
  wire f_u_cska12_fa6_and0;
  wire f_u_cska12_fa6_xor1;
  wire f_u_cska12_fa6_and1;
  wire f_u_cska12_fa6_or0;
  wire f_u_cska12_and_propagate13;
  wire f_u_cska12_and_propagate14;
  wire f_u_cska12_and_propagate15;
  wire f_u_cska12_mux2to11_and0;
  wire f_u_cska12_mux2to11_not0;
  wire f_u_cska12_mux2to11_and1;
  wire f_u_cska12_mux2to11_xor0;
  wire f_u_cska12_xor8;
  wire f_u_cska12_fa7_xor0;
  wire f_u_cska12_fa7_and0;
  wire f_u_cska12_fa7_xor1;
  wire f_u_cska12_fa7_and1;
  wire f_u_cska12_fa7_or0;
  wire f_u_cska12_xor9;
  wire f_u_cska12_fa8_xor0;
  wire f_u_cska12_fa8_and0;
  wire f_u_cska12_fa8_xor1;
  wire f_u_cska12_fa8_and1;
  wire f_u_cska12_fa8_or0;
  wire f_u_cska12_xor10;
  wire f_u_cska12_fa9_xor0;
  wire f_u_cska12_fa9_and0;
  wire f_u_cska12_fa9_xor1;
  wire f_u_cska12_fa9_and1;
  wire f_u_cska12_fa9_or0;
  wire f_u_cska12_xor11;
  wire f_u_cska12_fa10_xor0;
  wire f_u_cska12_fa10_and0;
  wire f_u_cska12_fa10_xor1;
  wire f_u_cska12_fa10_and1;
  wire f_u_cska12_fa10_or0;
  wire f_u_cska12_and_propagate26;
  wire f_u_cska12_and_propagate27;
  wire f_u_cska12_and_propagate28;
  wire f_u_cska12_mux2to12_and0;
  wire f_u_cska12_mux2to12_not0;
  wire f_u_cska12_mux2to12_and1;
  wire f_u_cska12_mux2to12_xor0;

  assign f_u_cska12_xor0 = a[0] ^ b[0];
  assign f_u_cska12_ha0_xor0 = a[0] ^ b[0];
  assign f_u_cska12_ha0_and0 = a[0] & b[0];
  assign f_u_cska12_xor1 = a[1] ^ b[1];
  assign f_u_cska12_fa0_xor0 = a[1] ^ b[1];
  assign f_u_cska12_fa0_and0 = a[1] & b[1];
  assign f_u_cska12_fa0_xor1 = f_u_cska12_fa0_xor0 ^ f_u_cska12_ha0_and0;
  assign f_u_cska12_fa0_and1 = f_u_cska12_fa0_xor0 & f_u_cska12_ha0_and0;
  assign f_u_cska12_fa0_or0 = f_u_cska12_fa0_and0 | f_u_cska12_fa0_and1;
  assign f_u_cska12_xor2 = a[2] ^ b[2];
  assign f_u_cska12_fa1_xor0 = a[2] ^ b[2];
  assign f_u_cska12_fa1_and0 = a[2] & b[2];
  assign f_u_cska12_fa1_xor1 = f_u_cska12_fa1_xor0 ^ f_u_cska12_fa0_or0;
  assign f_u_cska12_fa1_and1 = f_u_cska12_fa1_xor0 & f_u_cska12_fa0_or0;
  assign f_u_cska12_fa1_or0 = f_u_cska12_fa1_and0 | f_u_cska12_fa1_and1;
  assign f_u_cska12_xor3 = a[3] ^ b[3];
  assign f_u_cska12_fa2_xor0 = a[3] ^ b[3];
  assign f_u_cska12_fa2_and0 = a[3] & b[3];
  assign f_u_cska12_fa2_xor1 = f_u_cska12_fa2_xor0 ^ f_u_cska12_fa1_or0;
  assign f_u_cska12_fa2_and1 = f_u_cska12_fa2_xor0 & f_u_cska12_fa1_or0;
  assign f_u_cska12_fa2_or0 = f_u_cska12_fa2_and0 | f_u_cska12_fa2_and1;
  assign f_u_cska12_and_propagate00 = f_u_cska12_xor0 & f_u_cska12_xor2;
  assign f_u_cska12_and_propagate01 = f_u_cska12_xor1 & f_u_cska12_xor3;
  assign f_u_cska12_and_propagate02 = f_u_cska12_and_propagate00 & f_u_cska12_and_propagate01;
  assign f_u_cska12_mux2to10_not0 = ~f_u_cska12_and_propagate02;
  assign f_u_cska12_mux2to10_and1 = f_u_cska12_fa2_or0 & f_u_cska12_mux2to10_not0;
  assign f_u_cska12_xor4 = a[4] ^ b[4];
  assign f_u_cska12_fa3_xor0 = a[4] ^ b[4];
  assign f_u_cska12_fa3_and0 = a[4] & b[4];
  assign f_u_cska12_fa3_xor1 = f_u_cska12_fa3_xor0 ^ f_u_cska12_mux2to10_and1;
  assign f_u_cska12_fa3_and1 = f_u_cska12_fa3_xor0 & f_u_cska12_mux2to10_and1;
  assign f_u_cska12_fa3_or0 = f_u_cska12_fa3_and0 | f_u_cska12_fa3_and1;
  assign f_u_cska12_xor5 = a[5] ^ b[5];
  assign f_u_cska12_fa4_xor0 = a[5] ^ b[5];
  assign f_u_cska12_fa4_and0 = a[5] & b[5];
  assign f_u_cska12_fa4_xor1 = f_u_cska12_fa4_xor0 ^ f_u_cska12_fa3_or0;
  assign f_u_cska12_fa4_and1 = f_u_cska12_fa4_xor0 & f_u_cska12_fa3_or0;
  assign f_u_cska12_fa4_or0 = f_u_cska12_fa4_and0 | f_u_cska12_fa4_and1;
  assign f_u_cska12_xor6 = a[6] ^ b[6];
  assign f_u_cska12_fa5_xor0 = a[6] ^ b[6];
  assign f_u_cska12_fa5_and0 = a[6] & b[6];
  assign f_u_cska12_fa5_xor1 = f_u_cska12_fa5_xor0 ^ f_u_cska12_fa4_or0;
  assign f_u_cska12_fa5_and1 = f_u_cska12_fa5_xor0 & f_u_cska12_fa4_or0;
  assign f_u_cska12_fa5_or0 = f_u_cska12_fa5_and0 | f_u_cska12_fa5_and1;
  assign f_u_cska12_xor7 = a[7] ^ b[7];
  assign f_u_cska12_fa6_xor0 = a[7] ^ b[7];
  assign f_u_cska12_fa6_and0 = a[7] & b[7];
  assign f_u_cska12_fa6_xor1 = f_u_cska12_fa6_xor0 ^ f_u_cska12_fa5_or0;
  assign f_u_cska12_fa6_and1 = f_u_cska12_fa6_xor0 & f_u_cska12_fa5_or0;
  assign f_u_cska12_fa6_or0 = f_u_cska12_fa6_and0 | f_u_cska12_fa6_and1;
  assign f_u_cska12_and_propagate13 = f_u_cska12_xor4 & f_u_cska12_xor6;
  assign f_u_cska12_and_propagate14 = f_u_cska12_xor5 & f_u_cska12_xor7;
  assign f_u_cska12_and_propagate15 = f_u_cska12_and_propagate13 & f_u_cska12_and_propagate14;
  assign f_u_cska12_mux2to11_and0 = f_u_cska12_mux2to10_and1 & f_u_cska12_and_propagate15;
  assign f_u_cska12_mux2to11_not0 = ~f_u_cska12_and_propagate15;
  assign f_u_cska12_mux2to11_and1 = f_u_cska12_fa6_or0 & f_u_cska12_mux2to11_not0;
  assign f_u_cska12_mux2to11_xor0 = f_u_cska12_mux2to11_and0 ^ f_u_cska12_mux2to11_and1;
  assign f_u_cska12_xor8 = a[8] ^ b[8];
  assign f_u_cska12_fa7_xor0 = a[8] ^ b[8];
  assign f_u_cska12_fa7_and0 = a[8] & b[8];
  assign f_u_cska12_fa7_xor1 = f_u_cska12_fa7_xor0 ^ f_u_cska12_mux2to11_xor0;
  assign f_u_cska12_fa7_and1 = f_u_cska12_fa7_xor0 & f_u_cska12_mux2to11_xor0;
  assign f_u_cska12_fa7_or0 = f_u_cska12_fa7_and0 | f_u_cska12_fa7_and1;
  assign f_u_cska12_xor9 = a[9] ^ b[9];
  assign f_u_cska12_fa8_xor0 = a[9] ^ b[9];
  assign f_u_cska12_fa8_and0 = a[9] & b[9];
  assign f_u_cska12_fa8_xor1 = f_u_cska12_fa8_xor0 ^ f_u_cska12_fa7_or0;
  assign f_u_cska12_fa8_and1 = f_u_cska12_fa8_xor0 & f_u_cska12_fa7_or0;
  assign f_u_cska12_fa8_or0 = f_u_cska12_fa8_and0 | f_u_cska12_fa8_and1;
  assign f_u_cska12_xor10 = a[10] ^ b[10];
  assign f_u_cska12_fa9_xor0 = a[10] ^ b[10];
  assign f_u_cska12_fa9_and0 = a[10] & b[10];
  assign f_u_cska12_fa9_xor1 = f_u_cska12_fa9_xor0 ^ f_u_cska12_fa8_or0;
  assign f_u_cska12_fa9_and1 = f_u_cska12_fa9_xor0 & f_u_cska12_fa8_or0;
  assign f_u_cska12_fa9_or0 = f_u_cska12_fa9_and0 | f_u_cska12_fa9_and1;
  assign f_u_cska12_xor11 = a[11] ^ b[11];
  assign f_u_cska12_fa10_xor0 = a[11] ^ b[11];
  assign f_u_cska12_fa10_and0 = a[11] & b[11];
  assign f_u_cska12_fa10_xor1 = f_u_cska12_fa10_xor0 ^ f_u_cska12_fa9_or0;
  assign f_u_cska12_fa10_and1 = f_u_cska12_fa10_xor0 & f_u_cska12_fa9_or0;
  assign f_u_cska12_fa10_or0 = f_u_cska12_fa10_and0 | f_u_cska12_fa10_and1;
  assign f_u_cska12_and_propagate26 = f_u_cska12_xor8 & f_u_cska12_xor10;
  assign f_u_cska12_and_propagate27 = f_u_cska12_xor9 & f_u_cska12_xor11;
  assign f_u_cska12_and_propagate28 = f_u_cska12_and_propagate26 & f_u_cska12_and_propagate27;
  assign f_u_cska12_mux2to12_and0 = f_u_cska12_mux2to11_xor0 & f_u_cska12_and_propagate28;
  assign f_u_cska12_mux2to12_not0 = ~f_u_cska12_and_propagate28;
  assign f_u_cska12_mux2to12_and1 = f_u_cska12_fa10_or0 & f_u_cska12_mux2to12_not0;
  assign f_u_cska12_mux2to12_xor0 = f_u_cska12_mux2to12_and0 ^ f_u_cska12_mux2to12_and1;

  assign f_u_cska12_out[0] = f_u_cska12_ha0_xor0;
  assign f_u_cska12_out[1] = f_u_cska12_fa0_xor1;
  assign f_u_cska12_out[2] = f_u_cska12_fa1_xor1;
  assign f_u_cska12_out[3] = f_u_cska12_fa2_xor1;
  assign f_u_cska12_out[4] = f_u_cska12_fa3_xor1;
  assign f_u_cska12_out[5] = f_u_cska12_fa4_xor1;
  assign f_u_cska12_out[6] = f_u_cska12_fa5_xor1;
  assign f_u_cska12_out[7] = f_u_cska12_fa6_xor1;
  assign f_u_cska12_out[8] = f_u_cska12_fa7_xor1;
  assign f_u_cska12_out[9] = f_u_cska12_fa8_xor1;
  assign f_u_cska12_out[10] = f_u_cska12_fa9_xor1;
  assign f_u_cska12_out[11] = f_u_cska12_fa10_xor1;
  assign f_u_cska12_out[12] = f_u_cska12_mux2to12_xor0;
endmodule