module f_u_cla32(input [31:0] a, input [31:0] b, output [32:0] f_u_cla32_out);
  wire f_u_cla32_pg_logic0_or0;
  wire f_u_cla32_pg_logic0_and0;
  wire f_u_cla32_pg_logic0_xor0;
  wire f_u_cla32_pg_logic1_or0;
  wire f_u_cla32_pg_logic1_and0;
  wire f_u_cla32_pg_logic1_xor0;
  wire f_u_cla32_xor1;
  wire f_u_cla32_and0;
  wire f_u_cla32_or0;
  wire f_u_cla32_pg_logic2_or0;
  wire f_u_cla32_pg_logic2_and0;
  wire f_u_cla32_pg_logic2_xor0;
  wire f_u_cla32_xor2;
  wire f_u_cla32_and1;
  wire f_u_cla32_and2;
  wire f_u_cla32_and3;
  wire f_u_cla32_and4;
  wire f_u_cla32_or1;
  wire f_u_cla32_or2;
  wire f_u_cla32_pg_logic3_or0;
  wire f_u_cla32_pg_logic3_and0;
  wire f_u_cla32_pg_logic3_xor0;
  wire f_u_cla32_xor3;
  wire f_u_cla32_and5;
  wire f_u_cla32_and6;
  wire f_u_cla32_and7;
  wire f_u_cla32_and8;
  wire f_u_cla32_and9;
  wire f_u_cla32_and10;
  wire f_u_cla32_and11;
  wire f_u_cla32_or3;
  wire f_u_cla32_or4;
  wire f_u_cla32_or5;
  wire f_u_cla32_pg_logic4_or0;
  wire f_u_cla32_pg_logic4_and0;
  wire f_u_cla32_pg_logic4_xor0;
  wire f_u_cla32_xor4;
  wire f_u_cla32_and12;
  wire f_u_cla32_or6;
  wire f_u_cla32_pg_logic5_or0;
  wire f_u_cla32_pg_logic5_and0;
  wire f_u_cla32_pg_logic5_xor0;
  wire f_u_cla32_xor5;
  wire f_u_cla32_and13;
  wire f_u_cla32_and14;
  wire f_u_cla32_and15;
  wire f_u_cla32_or7;
  wire f_u_cla32_or8;
  wire f_u_cla32_pg_logic6_or0;
  wire f_u_cla32_pg_logic6_and0;
  wire f_u_cla32_pg_logic6_xor0;
  wire f_u_cla32_xor6;
  wire f_u_cla32_and16;
  wire f_u_cla32_and17;
  wire f_u_cla32_and18;
  wire f_u_cla32_and19;
  wire f_u_cla32_and20;
  wire f_u_cla32_and21;
  wire f_u_cla32_or9;
  wire f_u_cla32_or10;
  wire f_u_cla32_or11;
  wire f_u_cla32_pg_logic7_or0;
  wire f_u_cla32_pg_logic7_and0;
  wire f_u_cla32_pg_logic7_xor0;
  wire f_u_cla32_xor7;
  wire f_u_cla32_and22;
  wire f_u_cla32_and23;
  wire f_u_cla32_and24;
  wire f_u_cla32_and25;
  wire f_u_cla32_and26;
  wire f_u_cla32_and27;
  wire f_u_cla32_and28;
  wire f_u_cla32_and29;
  wire f_u_cla32_and30;
  wire f_u_cla32_and31;
  wire f_u_cla32_or12;
  wire f_u_cla32_or13;
  wire f_u_cla32_or14;
  wire f_u_cla32_or15;
  wire f_u_cla32_pg_logic8_or0;
  wire f_u_cla32_pg_logic8_and0;
  wire f_u_cla32_pg_logic8_xor0;
  wire f_u_cla32_xor8;
  wire f_u_cla32_and32;
  wire f_u_cla32_or16;
  wire f_u_cla32_pg_logic9_or0;
  wire f_u_cla32_pg_logic9_and0;
  wire f_u_cla32_pg_logic9_xor0;
  wire f_u_cla32_xor9;
  wire f_u_cla32_and33;
  wire f_u_cla32_and34;
  wire f_u_cla32_and35;
  wire f_u_cla32_or17;
  wire f_u_cla32_or18;
  wire f_u_cla32_pg_logic10_or0;
  wire f_u_cla32_pg_logic10_and0;
  wire f_u_cla32_pg_logic10_xor0;
  wire f_u_cla32_xor10;
  wire f_u_cla32_and36;
  wire f_u_cla32_and37;
  wire f_u_cla32_and38;
  wire f_u_cla32_and39;
  wire f_u_cla32_and40;
  wire f_u_cla32_and41;
  wire f_u_cla32_or19;
  wire f_u_cla32_or20;
  wire f_u_cla32_or21;
  wire f_u_cla32_pg_logic11_or0;
  wire f_u_cla32_pg_logic11_and0;
  wire f_u_cla32_pg_logic11_xor0;
  wire f_u_cla32_xor11;
  wire f_u_cla32_and42;
  wire f_u_cla32_and43;
  wire f_u_cla32_and44;
  wire f_u_cla32_and45;
  wire f_u_cla32_and46;
  wire f_u_cla32_and47;
  wire f_u_cla32_and48;
  wire f_u_cla32_and49;
  wire f_u_cla32_and50;
  wire f_u_cla32_and51;
  wire f_u_cla32_or22;
  wire f_u_cla32_or23;
  wire f_u_cla32_or24;
  wire f_u_cla32_or25;
  wire f_u_cla32_pg_logic12_or0;
  wire f_u_cla32_pg_logic12_and0;
  wire f_u_cla32_pg_logic12_xor0;
  wire f_u_cla32_xor12;
  wire f_u_cla32_and52;
  wire f_u_cla32_or26;
  wire f_u_cla32_pg_logic13_or0;
  wire f_u_cla32_pg_logic13_and0;
  wire f_u_cla32_pg_logic13_xor0;
  wire f_u_cla32_xor13;
  wire f_u_cla32_and53;
  wire f_u_cla32_and54;
  wire f_u_cla32_and55;
  wire f_u_cla32_or27;
  wire f_u_cla32_or28;
  wire f_u_cla32_pg_logic14_or0;
  wire f_u_cla32_pg_logic14_and0;
  wire f_u_cla32_pg_logic14_xor0;
  wire f_u_cla32_xor14;
  wire f_u_cla32_and56;
  wire f_u_cla32_and57;
  wire f_u_cla32_and58;
  wire f_u_cla32_and59;
  wire f_u_cla32_and60;
  wire f_u_cla32_and61;
  wire f_u_cla32_or29;
  wire f_u_cla32_or30;
  wire f_u_cla32_or31;
  wire f_u_cla32_pg_logic15_or0;
  wire f_u_cla32_pg_logic15_and0;
  wire f_u_cla32_pg_logic15_xor0;
  wire f_u_cla32_xor15;
  wire f_u_cla32_and62;
  wire f_u_cla32_and63;
  wire f_u_cla32_and64;
  wire f_u_cla32_and65;
  wire f_u_cla32_and66;
  wire f_u_cla32_and67;
  wire f_u_cla32_and68;
  wire f_u_cla32_and69;
  wire f_u_cla32_and70;
  wire f_u_cla32_and71;
  wire f_u_cla32_or32;
  wire f_u_cla32_or33;
  wire f_u_cla32_or34;
  wire f_u_cla32_or35;
  wire f_u_cla32_pg_logic16_or0;
  wire f_u_cla32_pg_logic16_and0;
  wire f_u_cla32_pg_logic16_xor0;
  wire f_u_cla32_xor16;
  wire f_u_cla32_and72;
  wire f_u_cla32_or36;
  wire f_u_cla32_pg_logic17_or0;
  wire f_u_cla32_pg_logic17_and0;
  wire f_u_cla32_pg_logic17_xor0;
  wire f_u_cla32_xor17;
  wire f_u_cla32_and73;
  wire f_u_cla32_and74;
  wire f_u_cla32_and75;
  wire f_u_cla32_or37;
  wire f_u_cla32_or38;
  wire f_u_cla32_pg_logic18_or0;
  wire f_u_cla32_pg_logic18_and0;
  wire f_u_cla32_pg_logic18_xor0;
  wire f_u_cla32_xor18;
  wire f_u_cla32_and76;
  wire f_u_cla32_and77;
  wire f_u_cla32_and78;
  wire f_u_cla32_and79;
  wire f_u_cla32_and80;
  wire f_u_cla32_and81;
  wire f_u_cla32_or39;
  wire f_u_cla32_or40;
  wire f_u_cla32_or41;
  wire f_u_cla32_pg_logic19_or0;
  wire f_u_cla32_pg_logic19_and0;
  wire f_u_cla32_pg_logic19_xor0;
  wire f_u_cla32_xor19;
  wire f_u_cla32_and82;
  wire f_u_cla32_and83;
  wire f_u_cla32_and84;
  wire f_u_cla32_and85;
  wire f_u_cla32_and86;
  wire f_u_cla32_and87;
  wire f_u_cla32_and88;
  wire f_u_cla32_and89;
  wire f_u_cla32_and90;
  wire f_u_cla32_and91;
  wire f_u_cla32_or42;
  wire f_u_cla32_or43;
  wire f_u_cla32_or44;
  wire f_u_cla32_or45;
  wire f_u_cla32_pg_logic20_or0;
  wire f_u_cla32_pg_logic20_and0;
  wire f_u_cla32_pg_logic20_xor0;
  wire f_u_cla32_xor20;
  wire f_u_cla32_and92;
  wire f_u_cla32_or46;
  wire f_u_cla32_pg_logic21_or0;
  wire f_u_cla32_pg_logic21_and0;
  wire f_u_cla32_pg_logic21_xor0;
  wire f_u_cla32_xor21;
  wire f_u_cla32_and93;
  wire f_u_cla32_and94;
  wire f_u_cla32_and95;
  wire f_u_cla32_or47;
  wire f_u_cla32_or48;
  wire f_u_cla32_pg_logic22_or0;
  wire f_u_cla32_pg_logic22_and0;
  wire f_u_cla32_pg_logic22_xor0;
  wire f_u_cla32_xor22;
  wire f_u_cla32_and96;
  wire f_u_cla32_and97;
  wire f_u_cla32_and98;
  wire f_u_cla32_and99;
  wire f_u_cla32_and100;
  wire f_u_cla32_and101;
  wire f_u_cla32_or49;
  wire f_u_cla32_or50;
  wire f_u_cla32_or51;
  wire f_u_cla32_pg_logic23_or0;
  wire f_u_cla32_pg_logic23_and0;
  wire f_u_cla32_pg_logic23_xor0;
  wire f_u_cla32_xor23;
  wire f_u_cla32_and102;
  wire f_u_cla32_and103;
  wire f_u_cla32_and104;
  wire f_u_cla32_and105;
  wire f_u_cla32_and106;
  wire f_u_cla32_and107;
  wire f_u_cla32_and108;
  wire f_u_cla32_and109;
  wire f_u_cla32_and110;
  wire f_u_cla32_and111;
  wire f_u_cla32_or52;
  wire f_u_cla32_or53;
  wire f_u_cla32_or54;
  wire f_u_cla32_or55;
  wire f_u_cla32_pg_logic24_or0;
  wire f_u_cla32_pg_logic24_and0;
  wire f_u_cla32_pg_logic24_xor0;
  wire f_u_cla32_xor24;
  wire f_u_cla32_and112;
  wire f_u_cla32_or56;
  wire f_u_cla32_pg_logic25_or0;
  wire f_u_cla32_pg_logic25_and0;
  wire f_u_cla32_pg_logic25_xor0;
  wire f_u_cla32_xor25;
  wire f_u_cla32_and113;
  wire f_u_cla32_and114;
  wire f_u_cla32_and115;
  wire f_u_cla32_or57;
  wire f_u_cla32_or58;
  wire f_u_cla32_pg_logic26_or0;
  wire f_u_cla32_pg_logic26_and0;
  wire f_u_cla32_pg_logic26_xor0;
  wire f_u_cla32_xor26;
  wire f_u_cla32_and116;
  wire f_u_cla32_and117;
  wire f_u_cla32_and118;
  wire f_u_cla32_and119;
  wire f_u_cla32_and120;
  wire f_u_cla32_and121;
  wire f_u_cla32_or59;
  wire f_u_cla32_or60;
  wire f_u_cla32_or61;
  wire f_u_cla32_pg_logic27_or0;
  wire f_u_cla32_pg_logic27_and0;
  wire f_u_cla32_pg_logic27_xor0;
  wire f_u_cla32_xor27;
  wire f_u_cla32_and122;
  wire f_u_cla32_and123;
  wire f_u_cla32_and124;
  wire f_u_cla32_and125;
  wire f_u_cla32_and126;
  wire f_u_cla32_and127;
  wire f_u_cla32_and128;
  wire f_u_cla32_and129;
  wire f_u_cla32_and130;
  wire f_u_cla32_and131;
  wire f_u_cla32_or62;
  wire f_u_cla32_or63;
  wire f_u_cla32_or64;
  wire f_u_cla32_or65;
  wire f_u_cla32_pg_logic28_or0;
  wire f_u_cla32_pg_logic28_and0;
  wire f_u_cla32_pg_logic28_xor0;
  wire f_u_cla32_xor28;
  wire f_u_cla32_and132;
  wire f_u_cla32_or66;
  wire f_u_cla32_pg_logic29_or0;
  wire f_u_cla32_pg_logic29_and0;
  wire f_u_cla32_pg_logic29_xor0;
  wire f_u_cla32_xor29;
  wire f_u_cla32_and133;
  wire f_u_cla32_and134;
  wire f_u_cla32_and135;
  wire f_u_cla32_or67;
  wire f_u_cla32_or68;
  wire f_u_cla32_pg_logic30_or0;
  wire f_u_cla32_pg_logic30_and0;
  wire f_u_cla32_pg_logic30_xor0;
  wire f_u_cla32_xor30;
  wire f_u_cla32_and136;
  wire f_u_cla32_and137;
  wire f_u_cla32_and138;
  wire f_u_cla32_and139;
  wire f_u_cla32_and140;
  wire f_u_cla32_and141;
  wire f_u_cla32_or69;
  wire f_u_cla32_or70;
  wire f_u_cla32_or71;
  wire f_u_cla32_pg_logic31_or0;
  wire f_u_cla32_pg_logic31_and0;
  wire f_u_cla32_pg_logic31_xor0;
  wire f_u_cla32_xor31;
  wire f_u_cla32_and142;
  wire f_u_cla32_and143;
  wire f_u_cla32_and144;
  wire f_u_cla32_and145;
  wire f_u_cla32_and146;
  wire f_u_cla32_and147;
  wire f_u_cla32_and148;
  wire f_u_cla32_and149;
  wire f_u_cla32_and150;
  wire f_u_cla32_and151;
  wire f_u_cla32_or72;
  wire f_u_cla32_or73;
  wire f_u_cla32_or74;
  wire f_u_cla32_or75;

  assign f_u_cla32_pg_logic0_or0 = a[0] | b[0];
  assign f_u_cla32_pg_logic0_and0 = a[0] & b[0];
  assign f_u_cla32_pg_logic0_xor0 = a[0] ^ b[0];
  assign f_u_cla32_pg_logic1_or0 = a[1] | b[1];
  assign f_u_cla32_pg_logic1_and0 = a[1] & b[1];
  assign f_u_cla32_pg_logic1_xor0 = a[1] ^ b[1];
  assign f_u_cla32_xor1 = f_u_cla32_pg_logic1_xor0 ^ f_u_cla32_pg_logic0_and0;
  assign f_u_cla32_and0 = f_u_cla32_pg_logic0_and0 & f_u_cla32_pg_logic1_or0;
  assign f_u_cla32_or0 = f_u_cla32_pg_logic1_and0 | f_u_cla32_and0;
  assign f_u_cla32_pg_logic2_or0 = a[2] | b[2];
  assign f_u_cla32_pg_logic2_and0 = a[2] & b[2];
  assign f_u_cla32_pg_logic2_xor0 = a[2] ^ b[2];
  assign f_u_cla32_xor2 = f_u_cla32_pg_logic2_xor0 ^ f_u_cla32_or0;
  assign f_u_cla32_and1 = f_u_cla32_pg_logic2_or0 & f_u_cla32_pg_logic0_or0;
  assign f_u_cla32_and2 = f_u_cla32_pg_logic0_and0 & f_u_cla32_pg_logic2_or0;
  assign f_u_cla32_and3 = f_u_cla32_and2 & f_u_cla32_pg_logic1_or0;
  assign f_u_cla32_and4 = f_u_cla32_pg_logic1_and0 & f_u_cla32_pg_logic2_or0;
  assign f_u_cla32_or1 = f_u_cla32_and3 | f_u_cla32_and4;
  assign f_u_cla32_or2 = f_u_cla32_pg_logic2_and0 | f_u_cla32_or1;
  assign f_u_cla32_pg_logic3_or0 = a[3] | b[3];
  assign f_u_cla32_pg_logic3_and0 = a[3] & b[3];
  assign f_u_cla32_pg_logic3_xor0 = a[3] ^ b[3];
  assign f_u_cla32_xor3 = f_u_cla32_pg_logic3_xor0 ^ f_u_cla32_or2;
  assign f_u_cla32_and5 = f_u_cla32_pg_logic3_or0 & f_u_cla32_pg_logic1_or0;
  assign f_u_cla32_and6 = f_u_cla32_pg_logic0_and0 & f_u_cla32_pg_logic2_or0;
  assign f_u_cla32_and7 = f_u_cla32_pg_logic3_or0 & f_u_cla32_pg_logic1_or0;
  assign f_u_cla32_and8 = f_u_cla32_and6 & f_u_cla32_and7;
  assign f_u_cla32_and9 = f_u_cla32_pg_logic1_and0 & f_u_cla32_pg_logic3_or0;
  assign f_u_cla32_and10 = f_u_cla32_and9 & f_u_cla32_pg_logic2_or0;
  assign f_u_cla32_and11 = f_u_cla32_pg_logic2_and0 & f_u_cla32_pg_logic3_or0;
  assign f_u_cla32_or3 = f_u_cla32_and8 | f_u_cla32_and11;
  assign f_u_cla32_or4 = f_u_cla32_and10 | f_u_cla32_or3;
  assign f_u_cla32_or5 = f_u_cla32_pg_logic3_and0 | f_u_cla32_or4;
  assign f_u_cla32_pg_logic4_or0 = a[4] | b[4];
  assign f_u_cla32_pg_logic4_and0 = a[4] & b[4];
  assign f_u_cla32_pg_logic4_xor0 = a[4] ^ b[4];
  assign f_u_cla32_xor4 = f_u_cla32_pg_logic4_xor0 ^ f_u_cla32_or5;
  assign f_u_cla32_and12 = f_u_cla32_or5 & f_u_cla32_pg_logic4_or0;
  assign f_u_cla32_or6 = f_u_cla32_pg_logic4_and0 | f_u_cla32_and12;
  assign f_u_cla32_pg_logic5_or0 = a[5] | b[5];
  assign f_u_cla32_pg_logic5_and0 = a[5] & b[5];
  assign f_u_cla32_pg_logic5_xor0 = a[5] ^ b[5];
  assign f_u_cla32_xor5 = f_u_cla32_pg_logic5_xor0 ^ f_u_cla32_or6;
  assign f_u_cla32_and13 = f_u_cla32_or5 & f_u_cla32_pg_logic5_or0;
  assign f_u_cla32_and14 = f_u_cla32_and13 & f_u_cla32_pg_logic4_or0;
  assign f_u_cla32_and15 = f_u_cla32_pg_logic4_and0 & f_u_cla32_pg_logic5_or0;
  assign f_u_cla32_or7 = f_u_cla32_and14 | f_u_cla32_and15;
  assign f_u_cla32_or8 = f_u_cla32_pg_logic5_and0 | f_u_cla32_or7;
  assign f_u_cla32_pg_logic6_or0 = a[6] | b[6];
  assign f_u_cla32_pg_logic6_and0 = a[6] & b[6];
  assign f_u_cla32_pg_logic6_xor0 = a[6] ^ b[6];
  assign f_u_cla32_xor6 = f_u_cla32_pg_logic6_xor0 ^ f_u_cla32_or8;
  assign f_u_cla32_and16 = f_u_cla32_or5 & f_u_cla32_pg_logic5_or0;
  assign f_u_cla32_and17 = f_u_cla32_pg_logic6_or0 & f_u_cla32_pg_logic4_or0;
  assign f_u_cla32_and18 = f_u_cla32_and16 & f_u_cla32_and17;
  assign f_u_cla32_and19 = f_u_cla32_pg_logic4_and0 & f_u_cla32_pg_logic6_or0;
  assign f_u_cla32_and20 = f_u_cla32_and19 & f_u_cla32_pg_logic5_or0;
  assign f_u_cla32_and21 = f_u_cla32_pg_logic5_and0 & f_u_cla32_pg_logic6_or0;
  assign f_u_cla32_or9 = f_u_cla32_and18 | f_u_cla32_and20;
  assign f_u_cla32_or10 = f_u_cla32_or9 | f_u_cla32_and21;
  assign f_u_cla32_or11 = f_u_cla32_pg_logic6_and0 | f_u_cla32_or10;
  assign f_u_cla32_pg_logic7_or0 = a[7] | b[7];
  assign f_u_cla32_pg_logic7_and0 = a[7] & b[7];
  assign f_u_cla32_pg_logic7_xor0 = a[7] ^ b[7];
  assign f_u_cla32_xor7 = f_u_cla32_pg_logic7_xor0 ^ f_u_cla32_or11;
  assign f_u_cla32_and22 = f_u_cla32_or5 & f_u_cla32_pg_logic6_or0;
  assign f_u_cla32_and23 = f_u_cla32_pg_logic7_or0 & f_u_cla32_pg_logic5_or0;
  assign f_u_cla32_and24 = f_u_cla32_and22 & f_u_cla32_and23;
  assign f_u_cla32_and25 = f_u_cla32_and24 & f_u_cla32_pg_logic4_or0;
  assign f_u_cla32_and26 = f_u_cla32_pg_logic4_and0 & f_u_cla32_pg_logic6_or0;
  assign f_u_cla32_and27 = f_u_cla32_pg_logic7_or0 & f_u_cla32_pg_logic5_or0;
  assign f_u_cla32_and28 = f_u_cla32_and26 & f_u_cla32_and27;
  assign f_u_cla32_and29 = f_u_cla32_pg_logic5_and0 & f_u_cla32_pg_logic7_or0;
  assign f_u_cla32_and30 = f_u_cla32_and29 & f_u_cla32_pg_logic6_or0;
  assign f_u_cla32_and31 = f_u_cla32_pg_logic6_and0 & f_u_cla32_pg_logic7_or0;
  assign f_u_cla32_or12 = f_u_cla32_and25 | f_u_cla32_and30;
  assign f_u_cla32_or13 = f_u_cla32_and28 | f_u_cla32_and31;
  assign f_u_cla32_or14 = f_u_cla32_or12 | f_u_cla32_or13;
  assign f_u_cla32_or15 = f_u_cla32_pg_logic7_and0 | f_u_cla32_or14;
  assign f_u_cla32_pg_logic8_or0 = a[8] | b[8];
  assign f_u_cla32_pg_logic8_and0 = a[8] & b[8];
  assign f_u_cla32_pg_logic8_xor0 = a[8] ^ b[8];
  assign f_u_cla32_xor8 = f_u_cla32_pg_logic8_xor0 ^ f_u_cla32_or15;
  assign f_u_cla32_and32 = f_u_cla32_or15 & f_u_cla32_pg_logic8_or0;
  assign f_u_cla32_or16 = f_u_cla32_pg_logic8_and0 | f_u_cla32_and32;
  assign f_u_cla32_pg_logic9_or0 = a[9] | b[9];
  assign f_u_cla32_pg_logic9_and0 = a[9] & b[9];
  assign f_u_cla32_pg_logic9_xor0 = a[9] ^ b[9];
  assign f_u_cla32_xor9 = f_u_cla32_pg_logic9_xor0 ^ f_u_cla32_or16;
  assign f_u_cla32_and33 = f_u_cla32_or15 & f_u_cla32_pg_logic9_or0;
  assign f_u_cla32_and34 = f_u_cla32_and33 & f_u_cla32_pg_logic8_or0;
  assign f_u_cla32_and35 = f_u_cla32_pg_logic8_and0 & f_u_cla32_pg_logic9_or0;
  assign f_u_cla32_or17 = f_u_cla32_and34 | f_u_cla32_and35;
  assign f_u_cla32_or18 = f_u_cla32_pg_logic9_and0 | f_u_cla32_or17;
  assign f_u_cla32_pg_logic10_or0 = a[10] | b[10];
  assign f_u_cla32_pg_logic10_and0 = a[10] & b[10];
  assign f_u_cla32_pg_logic10_xor0 = a[10] ^ b[10];
  assign f_u_cla32_xor10 = f_u_cla32_pg_logic10_xor0 ^ f_u_cla32_or18;
  assign f_u_cla32_and36 = f_u_cla32_or15 & f_u_cla32_pg_logic9_or0;
  assign f_u_cla32_and37 = f_u_cla32_pg_logic10_or0 & f_u_cla32_pg_logic8_or0;
  assign f_u_cla32_and38 = f_u_cla32_and36 & f_u_cla32_and37;
  assign f_u_cla32_and39 = f_u_cla32_pg_logic8_and0 & f_u_cla32_pg_logic10_or0;
  assign f_u_cla32_and40 = f_u_cla32_and39 & f_u_cla32_pg_logic9_or0;
  assign f_u_cla32_and41 = f_u_cla32_pg_logic9_and0 & f_u_cla32_pg_logic10_or0;
  assign f_u_cla32_or19 = f_u_cla32_and38 | f_u_cla32_and40;
  assign f_u_cla32_or20 = f_u_cla32_or19 | f_u_cla32_and41;
  assign f_u_cla32_or21 = f_u_cla32_pg_logic10_and0 | f_u_cla32_or20;
  assign f_u_cla32_pg_logic11_or0 = a[11] | b[11];
  assign f_u_cla32_pg_logic11_and0 = a[11] & b[11];
  assign f_u_cla32_pg_logic11_xor0 = a[11] ^ b[11];
  assign f_u_cla32_xor11 = f_u_cla32_pg_logic11_xor0 ^ f_u_cla32_or21;
  assign f_u_cla32_and42 = f_u_cla32_or15 & f_u_cla32_pg_logic10_or0;
  assign f_u_cla32_and43 = f_u_cla32_pg_logic11_or0 & f_u_cla32_pg_logic9_or0;
  assign f_u_cla32_and44 = f_u_cla32_and42 & f_u_cla32_and43;
  assign f_u_cla32_and45 = f_u_cla32_and44 & f_u_cla32_pg_logic8_or0;
  assign f_u_cla32_and46 = f_u_cla32_pg_logic8_and0 & f_u_cla32_pg_logic10_or0;
  assign f_u_cla32_and47 = f_u_cla32_pg_logic11_or0 & f_u_cla32_pg_logic9_or0;
  assign f_u_cla32_and48 = f_u_cla32_and46 & f_u_cla32_and47;
  assign f_u_cla32_and49 = f_u_cla32_pg_logic9_and0 & f_u_cla32_pg_logic11_or0;
  assign f_u_cla32_and50 = f_u_cla32_and49 & f_u_cla32_pg_logic10_or0;
  assign f_u_cla32_and51 = f_u_cla32_pg_logic10_and0 & f_u_cla32_pg_logic11_or0;
  assign f_u_cla32_or22 = f_u_cla32_and45 | f_u_cla32_and50;
  assign f_u_cla32_or23 = f_u_cla32_and48 | f_u_cla32_and51;
  assign f_u_cla32_or24 = f_u_cla32_or22 | f_u_cla32_or23;
  assign f_u_cla32_or25 = f_u_cla32_pg_logic11_and0 | f_u_cla32_or24;
  assign f_u_cla32_pg_logic12_or0 = a[12] | b[12];
  assign f_u_cla32_pg_logic12_and0 = a[12] & b[12];
  assign f_u_cla32_pg_logic12_xor0 = a[12] ^ b[12];
  assign f_u_cla32_xor12 = f_u_cla32_pg_logic12_xor0 ^ f_u_cla32_or25;
  assign f_u_cla32_and52 = f_u_cla32_or25 & f_u_cla32_pg_logic12_or0;
  assign f_u_cla32_or26 = f_u_cla32_pg_logic12_and0 | f_u_cla32_and52;
  assign f_u_cla32_pg_logic13_or0 = a[13] | b[13];
  assign f_u_cla32_pg_logic13_and0 = a[13] & b[13];
  assign f_u_cla32_pg_logic13_xor0 = a[13] ^ b[13];
  assign f_u_cla32_xor13 = f_u_cla32_pg_logic13_xor0 ^ f_u_cla32_or26;
  assign f_u_cla32_and53 = f_u_cla32_or25 & f_u_cla32_pg_logic13_or0;
  assign f_u_cla32_and54 = f_u_cla32_and53 & f_u_cla32_pg_logic12_or0;
  assign f_u_cla32_and55 = f_u_cla32_pg_logic12_and0 & f_u_cla32_pg_logic13_or0;
  assign f_u_cla32_or27 = f_u_cla32_and54 | f_u_cla32_and55;
  assign f_u_cla32_or28 = f_u_cla32_pg_logic13_and0 | f_u_cla32_or27;
  assign f_u_cla32_pg_logic14_or0 = a[14] | b[14];
  assign f_u_cla32_pg_logic14_and0 = a[14] & b[14];
  assign f_u_cla32_pg_logic14_xor0 = a[14] ^ b[14];
  assign f_u_cla32_xor14 = f_u_cla32_pg_logic14_xor0 ^ f_u_cla32_or28;
  assign f_u_cla32_and56 = f_u_cla32_or25 & f_u_cla32_pg_logic13_or0;
  assign f_u_cla32_and57 = f_u_cla32_pg_logic14_or0 & f_u_cla32_pg_logic12_or0;
  assign f_u_cla32_and58 = f_u_cla32_and56 & f_u_cla32_and57;
  assign f_u_cla32_and59 = f_u_cla32_pg_logic12_and0 & f_u_cla32_pg_logic14_or0;
  assign f_u_cla32_and60 = f_u_cla32_and59 & f_u_cla32_pg_logic13_or0;
  assign f_u_cla32_and61 = f_u_cla32_pg_logic13_and0 & f_u_cla32_pg_logic14_or0;
  assign f_u_cla32_or29 = f_u_cla32_and58 | f_u_cla32_and60;
  assign f_u_cla32_or30 = f_u_cla32_or29 | f_u_cla32_and61;
  assign f_u_cla32_or31 = f_u_cla32_pg_logic14_and0 | f_u_cla32_or30;
  assign f_u_cla32_pg_logic15_or0 = a[15] | b[15];
  assign f_u_cla32_pg_logic15_and0 = a[15] & b[15];
  assign f_u_cla32_pg_logic15_xor0 = a[15] ^ b[15];
  assign f_u_cla32_xor15 = f_u_cla32_pg_logic15_xor0 ^ f_u_cla32_or31;
  assign f_u_cla32_and62 = f_u_cla32_or25 & f_u_cla32_pg_logic14_or0;
  assign f_u_cla32_and63 = f_u_cla32_pg_logic15_or0 & f_u_cla32_pg_logic13_or0;
  assign f_u_cla32_and64 = f_u_cla32_and62 & f_u_cla32_and63;
  assign f_u_cla32_and65 = f_u_cla32_and64 & f_u_cla32_pg_logic12_or0;
  assign f_u_cla32_and66 = f_u_cla32_pg_logic12_and0 & f_u_cla32_pg_logic14_or0;
  assign f_u_cla32_and67 = f_u_cla32_pg_logic15_or0 & f_u_cla32_pg_logic13_or0;
  assign f_u_cla32_and68 = f_u_cla32_and66 & f_u_cla32_and67;
  assign f_u_cla32_and69 = f_u_cla32_pg_logic13_and0 & f_u_cla32_pg_logic15_or0;
  assign f_u_cla32_and70 = f_u_cla32_and69 & f_u_cla32_pg_logic14_or0;
  assign f_u_cla32_and71 = f_u_cla32_pg_logic14_and0 & f_u_cla32_pg_logic15_or0;
  assign f_u_cla32_or32 = f_u_cla32_and65 | f_u_cla32_and70;
  assign f_u_cla32_or33 = f_u_cla32_and68 | f_u_cla32_and71;
  assign f_u_cla32_or34 = f_u_cla32_or32 | f_u_cla32_or33;
  assign f_u_cla32_or35 = f_u_cla32_pg_logic15_and0 | f_u_cla32_or34;
  assign f_u_cla32_pg_logic16_or0 = a[16] | b[16];
  assign f_u_cla32_pg_logic16_and0 = a[16] & b[16];
  assign f_u_cla32_pg_logic16_xor0 = a[16] ^ b[16];
  assign f_u_cla32_xor16 = f_u_cla32_pg_logic16_xor0 ^ f_u_cla32_or35;
  assign f_u_cla32_and72 = f_u_cla32_or35 & f_u_cla32_pg_logic16_or0;
  assign f_u_cla32_or36 = f_u_cla32_pg_logic16_and0 | f_u_cla32_and72;
  assign f_u_cla32_pg_logic17_or0 = a[17] | b[17];
  assign f_u_cla32_pg_logic17_and0 = a[17] & b[17];
  assign f_u_cla32_pg_logic17_xor0 = a[17] ^ b[17];
  assign f_u_cla32_xor17 = f_u_cla32_pg_logic17_xor0 ^ f_u_cla32_or36;
  assign f_u_cla32_and73 = f_u_cla32_or35 & f_u_cla32_pg_logic17_or0;
  assign f_u_cla32_and74 = f_u_cla32_and73 & f_u_cla32_pg_logic16_or0;
  assign f_u_cla32_and75 = f_u_cla32_pg_logic16_and0 & f_u_cla32_pg_logic17_or0;
  assign f_u_cla32_or37 = f_u_cla32_and74 | f_u_cla32_and75;
  assign f_u_cla32_or38 = f_u_cla32_pg_logic17_and0 | f_u_cla32_or37;
  assign f_u_cla32_pg_logic18_or0 = a[18] | b[18];
  assign f_u_cla32_pg_logic18_and0 = a[18] & b[18];
  assign f_u_cla32_pg_logic18_xor0 = a[18] ^ b[18];
  assign f_u_cla32_xor18 = f_u_cla32_pg_logic18_xor0 ^ f_u_cla32_or38;
  assign f_u_cla32_and76 = f_u_cla32_or35 & f_u_cla32_pg_logic17_or0;
  assign f_u_cla32_and77 = f_u_cla32_pg_logic18_or0 & f_u_cla32_pg_logic16_or0;
  assign f_u_cla32_and78 = f_u_cla32_and76 & f_u_cla32_and77;
  assign f_u_cla32_and79 = f_u_cla32_pg_logic16_and0 & f_u_cla32_pg_logic18_or0;
  assign f_u_cla32_and80 = f_u_cla32_and79 & f_u_cla32_pg_logic17_or0;
  assign f_u_cla32_and81 = f_u_cla32_pg_logic17_and0 & f_u_cla32_pg_logic18_or0;
  assign f_u_cla32_or39 = f_u_cla32_and78 | f_u_cla32_and80;
  assign f_u_cla32_or40 = f_u_cla32_or39 | f_u_cla32_and81;
  assign f_u_cla32_or41 = f_u_cla32_pg_logic18_and0 | f_u_cla32_or40;
  assign f_u_cla32_pg_logic19_or0 = a[19] | b[19];
  assign f_u_cla32_pg_logic19_and0 = a[19] & b[19];
  assign f_u_cla32_pg_logic19_xor0 = a[19] ^ b[19];
  assign f_u_cla32_xor19 = f_u_cla32_pg_logic19_xor0 ^ f_u_cla32_or41;
  assign f_u_cla32_and82 = f_u_cla32_or35 & f_u_cla32_pg_logic18_or0;
  assign f_u_cla32_and83 = f_u_cla32_pg_logic19_or0 & f_u_cla32_pg_logic17_or0;
  assign f_u_cla32_and84 = f_u_cla32_and82 & f_u_cla32_and83;
  assign f_u_cla32_and85 = f_u_cla32_and84 & f_u_cla32_pg_logic16_or0;
  assign f_u_cla32_and86 = f_u_cla32_pg_logic16_and0 & f_u_cla32_pg_logic18_or0;
  assign f_u_cla32_and87 = f_u_cla32_pg_logic19_or0 & f_u_cla32_pg_logic17_or0;
  assign f_u_cla32_and88 = f_u_cla32_and86 & f_u_cla32_and87;
  assign f_u_cla32_and89 = f_u_cla32_pg_logic17_and0 & f_u_cla32_pg_logic19_or0;
  assign f_u_cla32_and90 = f_u_cla32_and89 & f_u_cla32_pg_logic18_or0;
  assign f_u_cla32_and91 = f_u_cla32_pg_logic18_and0 & f_u_cla32_pg_logic19_or0;
  assign f_u_cla32_or42 = f_u_cla32_and85 | f_u_cla32_and90;
  assign f_u_cla32_or43 = f_u_cla32_and88 | f_u_cla32_and91;
  assign f_u_cla32_or44 = f_u_cla32_or42 | f_u_cla32_or43;
  assign f_u_cla32_or45 = f_u_cla32_pg_logic19_and0 | f_u_cla32_or44;
  assign f_u_cla32_pg_logic20_or0 = a[20] | b[20];
  assign f_u_cla32_pg_logic20_and0 = a[20] & b[20];
  assign f_u_cla32_pg_logic20_xor0 = a[20] ^ b[20];
  assign f_u_cla32_xor20 = f_u_cla32_pg_logic20_xor0 ^ f_u_cla32_or45;
  assign f_u_cla32_and92 = f_u_cla32_or45 & f_u_cla32_pg_logic20_or0;
  assign f_u_cla32_or46 = f_u_cla32_pg_logic20_and0 | f_u_cla32_and92;
  assign f_u_cla32_pg_logic21_or0 = a[21] | b[21];
  assign f_u_cla32_pg_logic21_and0 = a[21] & b[21];
  assign f_u_cla32_pg_logic21_xor0 = a[21] ^ b[21];
  assign f_u_cla32_xor21 = f_u_cla32_pg_logic21_xor0 ^ f_u_cla32_or46;
  assign f_u_cla32_and93 = f_u_cla32_or45 & f_u_cla32_pg_logic21_or0;
  assign f_u_cla32_and94 = f_u_cla32_and93 & f_u_cla32_pg_logic20_or0;
  assign f_u_cla32_and95 = f_u_cla32_pg_logic20_and0 & f_u_cla32_pg_logic21_or0;
  assign f_u_cla32_or47 = f_u_cla32_and94 | f_u_cla32_and95;
  assign f_u_cla32_or48 = f_u_cla32_pg_logic21_and0 | f_u_cla32_or47;
  assign f_u_cla32_pg_logic22_or0 = a[22] | b[22];
  assign f_u_cla32_pg_logic22_and0 = a[22] & b[22];
  assign f_u_cla32_pg_logic22_xor0 = a[22] ^ b[22];
  assign f_u_cla32_xor22 = f_u_cla32_pg_logic22_xor0 ^ f_u_cla32_or48;
  assign f_u_cla32_and96 = f_u_cla32_or45 & f_u_cla32_pg_logic21_or0;
  assign f_u_cla32_and97 = f_u_cla32_pg_logic22_or0 & f_u_cla32_pg_logic20_or0;
  assign f_u_cla32_and98 = f_u_cla32_and96 & f_u_cla32_and97;
  assign f_u_cla32_and99 = f_u_cla32_pg_logic20_and0 & f_u_cla32_pg_logic22_or0;
  assign f_u_cla32_and100 = f_u_cla32_and99 & f_u_cla32_pg_logic21_or0;
  assign f_u_cla32_and101 = f_u_cla32_pg_logic21_and0 & f_u_cla32_pg_logic22_or0;
  assign f_u_cla32_or49 = f_u_cla32_and98 | f_u_cla32_and100;
  assign f_u_cla32_or50 = f_u_cla32_or49 | f_u_cla32_and101;
  assign f_u_cla32_or51 = f_u_cla32_pg_logic22_and0 | f_u_cla32_or50;
  assign f_u_cla32_pg_logic23_or0 = a[23] | b[23];
  assign f_u_cla32_pg_logic23_and0 = a[23] & b[23];
  assign f_u_cla32_pg_logic23_xor0 = a[23] ^ b[23];
  assign f_u_cla32_xor23 = f_u_cla32_pg_logic23_xor0 ^ f_u_cla32_or51;
  assign f_u_cla32_and102 = f_u_cla32_or45 & f_u_cla32_pg_logic22_or0;
  assign f_u_cla32_and103 = f_u_cla32_pg_logic23_or0 & f_u_cla32_pg_logic21_or0;
  assign f_u_cla32_and104 = f_u_cla32_and102 & f_u_cla32_and103;
  assign f_u_cla32_and105 = f_u_cla32_and104 & f_u_cla32_pg_logic20_or0;
  assign f_u_cla32_and106 = f_u_cla32_pg_logic20_and0 & f_u_cla32_pg_logic22_or0;
  assign f_u_cla32_and107 = f_u_cla32_pg_logic23_or0 & f_u_cla32_pg_logic21_or0;
  assign f_u_cla32_and108 = f_u_cla32_and106 & f_u_cla32_and107;
  assign f_u_cla32_and109 = f_u_cla32_pg_logic21_and0 & f_u_cla32_pg_logic23_or0;
  assign f_u_cla32_and110 = f_u_cla32_and109 & f_u_cla32_pg_logic22_or0;
  assign f_u_cla32_and111 = f_u_cla32_pg_logic22_and0 & f_u_cla32_pg_logic23_or0;
  assign f_u_cla32_or52 = f_u_cla32_and105 | f_u_cla32_and110;
  assign f_u_cla32_or53 = f_u_cla32_and108 | f_u_cla32_and111;
  assign f_u_cla32_or54 = f_u_cla32_or52 | f_u_cla32_or53;
  assign f_u_cla32_or55 = f_u_cla32_pg_logic23_and0 | f_u_cla32_or54;
  assign f_u_cla32_pg_logic24_or0 = a[24] | b[24];
  assign f_u_cla32_pg_logic24_and0 = a[24] & b[24];
  assign f_u_cla32_pg_logic24_xor0 = a[24] ^ b[24];
  assign f_u_cla32_xor24 = f_u_cla32_pg_logic24_xor0 ^ f_u_cla32_or55;
  assign f_u_cla32_and112 = f_u_cla32_or55 & f_u_cla32_pg_logic24_or0;
  assign f_u_cla32_or56 = f_u_cla32_pg_logic24_and0 | f_u_cla32_and112;
  assign f_u_cla32_pg_logic25_or0 = a[25] | b[25];
  assign f_u_cla32_pg_logic25_and0 = a[25] & b[25];
  assign f_u_cla32_pg_logic25_xor0 = a[25] ^ b[25];
  assign f_u_cla32_xor25 = f_u_cla32_pg_logic25_xor0 ^ f_u_cla32_or56;
  assign f_u_cla32_and113 = f_u_cla32_or55 & f_u_cla32_pg_logic25_or0;
  assign f_u_cla32_and114 = f_u_cla32_and113 & f_u_cla32_pg_logic24_or0;
  assign f_u_cla32_and115 = f_u_cla32_pg_logic24_and0 & f_u_cla32_pg_logic25_or0;
  assign f_u_cla32_or57 = f_u_cla32_and114 | f_u_cla32_and115;
  assign f_u_cla32_or58 = f_u_cla32_pg_logic25_and0 | f_u_cla32_or57;
  assign f_u_cla32_pg_logic26_or0 = a[26] | b[26];
  assign f_u_cla32_pg_logic26_and0 = a[26] & b[26];
  assign f_u_cla32_pg_logic26_xor0 = a[26] ^ b[26];
  assign f_u_cla32_xor26 = f_u_cla32_pg_logic26_xor0 ^ f_u_cla32_or58;
  assign f_u_cla32_and116 = f_u_cla32_or55 & f_u_cla32_pg_logic25_or0;
  assign f_u_cla32_and117 = f_u_cla32_pg_logic26_or0 & f_u_cla32_pg_logic24_or0;
  assign f_u_cla32_and118 = f_u_cla32_and116 & f_u_cla32_and117;
  assign f_u_cla32_and119 = f_u_cla32_pg_logic24_and0 & f_u_cla32_pg_logic26_or0;
  assign f_u_cla32_and120 = f_u_cla32_and119 & f_u_cla32_pg_logic25_or0;
  assign f_u_cla32_and121 = f_u_cla32_pg_logic25_and0 & f_u_cla32_pg_logic26_or0;
  assign f_u_cla32_or59 = f_u_cla32_and118 | f_u_cla32_and120;
  assign f_u_cla32_or60 = f_u_cla32_or59 | f_u_cla32_and121;
  assign f_u_cla32_or61 = f_u_cla32_pg_logic26_and0 | f_u_cla32_or60;
  assign f_u_cla32_pg_logic27_or0 = a[27] | b[27];
  assign f_u_cla32_pg_logic27_and0 = a[27] & b[27];
  assign f_u_cla32_pg_logic27_xor0 = a[27] ^ b[27];
  assign f_u_cla32_xor27 = f_u_cla32_pg_logic27_xor0 ^ f_u_cla32_or61;
  assign f_u_cla32_and122 = f_u_cla32_or55 & f_u_cla32_pg_logic26_or0;
  assign f_u_cla32_and123 = f_u_cla32_pg_logic27_or0 & f_u_cla32_pg_logic25_or0;
  assign f_u_cla32_and124 = f_u_cla32_and122 & f_u_cla32_and123;
  assign f_u_cla32_and125 = f_u_cla32_and124 & f_u_cla32_pg_logic24_or0;
  assign f_u_cla32_and126 = f_u_cla32_pg_logic24_and0 & f_u_cla32_pg_logic26_or0;
  assign f_u_cla32_and127 = f_u_cla32_pg_logic27_or0 & f_u_cla32_pg_logic25_or0;
  assign f_u_cla32_and128 = f_u_cla32_and126 & f_u_cla32_and127;
  assign f_u_cla32_and129 = f_u_cla32_pg_logic25_and0 & f_u_cla32_pg_logic27_or0;
  assign f_u_cla32_and130 = f_u_cla32_and129 & f_u_cla32_pg_logic26_or0;
  assign f_u_cla32_and131 = f_u_cla32_pg_logic26_and0 & f_u_cla32_pg_logic27_or0;
  assign f_u_cla32_or62 = f_u_cla32_and125 | f_u_cla32_and130;
  assign f_u_cla32_or63 = f_u_cla32_and128 | f_u_cla32_and131;
  assign f_u_cla32_or64 = f_u_cla32_or62 | f_u_cla32_or63;
  assign f_u_cla32_or65 = f_u_cla32_pg_logic27_and0 | f_u_cla32_or64;
  assign f_u_cla32_pg_logic28_or0 = a[28] | b[28];
  assign f_u_cla32_pg_logic28_and0 = a[28] & b[28];
  assign f_u_cla32_pg_logic28_xor0 = a[28] ^ b[28];
  assign f_u_cla32_xor28 = f_u_cla32_pg_logic28_xor0 ^ f_u_cla32_or65;
  assign f_u_cla32_and132 = f_u_cla32_or65 & f_u_cla32_pg_logic28_or0;
  assign f_u_cla32_or66 = f_u_cla32_pg_logic28_and0 | f_u_cla32_and132;
  assign f_u_cla32_pg_logic29_or0 = a[29] | b[29];
  assign f_u_cla32_pg_logic29_and0 = a[29] & b[29];
  assign f_u_cla32_pg_logic29_xor0 = a[29] ^ b[29];
  assign f_u_cla32_xor29 = f_u_cla32_pg_logic29_xor0 ^ f_u_cla32_or66;
  assign f_u_cla32_and133 = f_u_cla32_or65 & f_u_cla32_pg_logic29_or0;
  assign f_u_cla32_and134 = f_u_cla32_and133 & f_u_cla32_pg_logic28_or0;
  assign f_u_cla32_and135 = f_u_cla32_pg_logic28_and0 & f_u_cla32_pg_logic29_or0;
  assign f_u_cla32_or67 = f_u_cla32_and134 | f_u_cla32_and135;
  assign f_u_cla32_or68 = f_u_cla32_pg_logic29_and0 | f_u_cla32_or67;
  assign f_u_cla32_pg_logic30_or0 = a[30] | b[30];
  assign f_u_cla32_pg_logic30_and0 = a[30] & b[30];
  assign f_u_cla32_pg_logic30_xor0 = a[30] ^ b[30];
  assign f_u_cla32_xor30 = f_u_cla32_pg_logic30_xor0 ^ f_u_cla32_or68;
  assign f_u_cla32_and136 = f_u_cla32_or65 & f_u_cla32_pg_logic29_or0;
  assign f_u_cla32_and137 = f_u_cla32_pg_logic30_or0 & f_u_cla32_pg_logic28_or0;
  assign f_u_cla32_and138 = f_u_cla32_and136 & f_u_cla32_and137;
  assign f_u_cla32_and139 = f_u_cla32_pg_logic28_and0 & f_u_cla32_pg_logic30_or0;
  assign f_u_cla32_and140 = f_u_cla32_and139 & f_u_cla32_pg_logic29_or0;
  assign f_u_cla32_and141 = f_u_cla32_pg_logic29_and0 & f_u_cla32_pg_logic30_or0;
  assign f_u_cla32_or69 = f_u_cla32_and138 | f_u_cla32_and140;
  assign f_u_cla32_or70 = f_u_cla32_or69 | f_u_cla32_and141;
  assign f_u_cla32_or71 = f_u_cla32_pg_logic30_and0 | f_u_cla32_or70;
  assign f_u_cla32_pg_logic31_or0 = a[31] | b[31];
  assign f_u_cla32_pg_logic31_and0 = a[31] & b[31];
  assign f_u_cla32_pg_logic31_xor0 = a[31] ^ b[31];
  assign f_u_cla32_xor31 = f_u_cla32_pg_logic31_xor0 ^ f_u_cla32_or71;
  assign f_u_cla32_and142 = f_u_cla32_or65 & f_u_cla32_pg_logic30_or0;
  assign f_u_cla32_and143 = f_u_cla32_pg_logic31_or0 & f_u_cla32_pg_logic29_or0;
  assign f_u_cla32_and144 = f_u_cla32_and142 & f_u_cla32_and143;
  assign f_u_cla32_and145 = f_u_cla32_and144 & f_u_cla32_pg_logic28_or0;
  assign f_u_cla32_and146 = f_u_cla32_pg_logic28_and0 & f_u_cla32_pg_logic30_or0;
  assign f_u_cla32_and147 = f_u_cla32_pg_logic31_or0 & f_u_cla32_pg_logic29_or0;
  assign f_u_cla32_and148 = f_u_cla32_and146 & f_u_cla32_and147;
  assign f_u_cla32_and149 = f_u_cla32_pg_logic29_and0 & f_u_cla32_pg_logic31_or0;
  assign f_u_cla32_and150 = f_u_cla32_and149 & f_u_cla32_pg_logic30_or0;
  assign f_u_cla32_and151 = f_u_cla32_pg_logic30_and0 & f_u_cla32_pg_logic31_or0;
  assign f_u_cla32_or72 = f_u_cla32_and145 | f_u_cla32_and150;
  assign f_u_cla32_or73 = f_u_cla32_and148 | f_u_cla32_and151;
  assign f_u_cla32_or74 = f_u_cla32_or72 | f_u_cla32_or73;
  assign f_u_cla32_or75 = f_u_cla32_pg_logic31_and0 | f_u_cla32_or74;

  assign f_u_cla32_out[0] = f_u_cla32_pg_logic0_xor0;
  assign f_u_cla32_out[1] = f_u_cla32_xor1;
  assign f_u_cla32_out[2] = f_u_cla32_xor2;
  assign f_u_cla32_out[3] = f_u_cla32_xor3;
  assign f_u_cla32_out[4] = f_u_cla32_xor4;
  assign f_u_cla32_out[5] = f_u_cla32_xor5;
  assign f_u_cla32_out[6] = f_u_cla32_xor6;
  assign f_u_cla32_out[7] = f_u_cla32_xor7;
  assign f_u_cla32_out[8] = f_u_cla32_xor8;
  assign f_u_cla32_out[9] = f_u_cla32_xor9;
  assign f_u_cla32_out[10] = f_u_cla32_xor10;
  assign f_u_cla32_out[11] = f_u_cla32_xor11;
  assign f_u_cla32_out[12] = f_u_cla32_xor12;
  assign f_u_cla32_out[13] = f_u_cla32_xor13;
  assign f_u_cla32_out[14] = f_u_cla32_xor14;
  assign f_u_cla32_out[15] = f_u_cla32_xor15;
  assign f_u_cla32_out[16] = f_u_cla32_xor16;
  assign f_u_cla32_out[17] = f_u_cla32_xor17;
  assign f_u_cla32_out[18] = f_u_cla32_xor18;
  assign f_u_cla32_out[19] = f_u_cla32_xor19;
  assign f_u_cla32_out[20] = f_u_cla32_xor20;
  assign f_u_cla32_out[21] = f_u_cla32_xor21;
  assign f_u_cla32_out[22] = f_u_cla32_xor22;
  assign f_u_cla32_out[23] = f_u_cla32_xor23;
  assign f_u_cla32_out[24] = f_u_cla32_xor24;
  assign f_u_cla32_out[25] = f_u_cla32_xor25;
  assign f_u_cla32_out[26] = f_u_cla32_xor26;
  assign f_u_cla32_out[27] = f_u_cla32_xor27;
  assign f_u_cla32_out[28] = f_u_cla32_xor28;
  assign f_u_cla32_out[29] = f_u_cla32_xor29;
  assign f_u_cla32_out[30] = f_u_cla32_xor30;
  assign f_u_cla32_out[31] = f_u_cla32_xor31;
  assign f_u_cla32_out[32] = f_u_cla32_or75;
endmodule