module s_wallace_cla8(input [7:0] a, input [7:0] b, output [15:0] s_wallace_cla8_out);
  wire s_wallace_cla8_and_2_0;
  wire s_wallace_cla8_and_1_1;
  wire s_wallace_cla8_ha0_xor0;
  wire s_wallace_cla8_ha0_and0;
  wire s_wallace_cla8_and_3_0;
  wire s_wallace_cla8_and_2_1;
  wire s_wallace_cla8_fa0_xor0;
  wire s_wallace_cla8_fa0_and0;
  wire s_wallace_cla8_fa0_xor1;
  wire s_wallace_cla8_fa0_and1;
  wire s_wallace_cla8_fa0_or0;
  wire s_wallace_cla8_and_4_0;
  wire s_wallace_cla8_and_3_1;
  wire s_wallace_cla8_fa1_xor0;
  wire s_wallace_cla8_fa1_and0;
  wire s_wallace_cla8_fa1_xor1;
  wire s_wallace_cla8_fa1_and1;
  wire s_wallace_cla8_fa1_or0;
  wire s_wallace_cla8_and_5_0;
  wire s_wallace_cla8_and_4_1;
  wire s_wallace_cla8_fa2_xor0;
  wire s_wallace_cla8_fa2_and0;
  wire s_wallace_cla8_fa2_xor1;
  wire s_wallace_cla8_fa2_and1;
  wire s_wallace_cla8_fa2_or0;
  wire s_wallace_cla8_and_6_0;
  wire s_wallace_cla8_and_5_1;
  wire s_wallace_cla8_fa3_xor0;
  wire s_wallace_cla8_fa3_and0;
  wire s_wallace_cla8_fa3_xor1;
  wire s_wallace_cla8_fa3_and1;
  wire s_wallace_cla8_fa3_or0;
  wire s_wallace_cla8_nand_7_0;
  wire s_wallace_cla8_and_6_1;
  wire s_wallace_cla8_fa4_xor0;
  wire s_wallace_cla8_fa4_and0;
  wire s_wallace_cla8_fa4_xor1;
  wire s_wallace_cla8_fa4_and1;
  wire s_wallace_cla8_fa4_or0;
  wire s_wallace_cla8_nand_7_1;
  wire s_wallace_cla8_fa5_xor0;
  wire s_wallace_cla8_fa5_xor1;
  wire s_wallace_cla8_fa5_and1;
  wire s_wallace_cla8_fa5_or0;
  wire s_wallace_cla8_nand_7_2;
  wire s_wallace_cla8_and_6_3;
  wire s_wallace_cla8_fa6_xor0;
  wire s_wallace_cla8_fa6_and0;
  wire s_wallace_cla8_fa6_xor1;
  wire s_wallace_cla8_fa6_and1;
  wire s_wallace_cla8_fa6_or0;
  wire s_wallace_cla8_nand_7_3;
  wire s_wallace_cla8_and_6_4;
  wire s_wallace_cla8_fa7_xor0;
  wire s_wallace_cla8_fa7_and0;
  wire s_wallace_cla8_fa7_xor1;
  wire s_wallace_cla8_fa7_and1;
  wire s_wallace_cla8_fa7_or0;
  wire s_wallace_cla8_nand_7_4;
  wire s_wallace_cla8_and_6_5;
  wire s_wallace_cla8_fa8_xor0;
  wire s_wallace_cla8_fa8_and0;
  wire s_wallace_cla8_fa8_xor1;
  wire s_wallace_cla8_fa8_and1;
  wire s_wallace_cla8_fa8_or0;
  wire s_wallace_cla8_nand_7_5;
  wire s_wallace_cla8_and_6_6;
  wire s_wallace_cla8_fa9_xor0;
  wire s_wallace_cla8_fa9_and0;
  wire s_wallace_cla8_fa9_xor1;
  wire s_wallace_cla8_fa9_and1;
  wire s_wallace_cla8_fa9_or0;
  wire s_wallace_cla8_and_1_2;
  wire s_wallace_cla8_and_0_3;
  wire s_wallace_cla8_ha1_xor0;
  wire s_wallace_cla8_ha1_and0;
  wire s_wallace_cla8_and_2_2;
  wire s_wallace_cla8_and_1_3;
  wire s_wallace_cla8_fa10_xor0;
  wire s_wallace_cla8_fa10_and0;
  wire s_wallace_cla8_fa10_xor1;
  wire s_wallace_cla8_fa10_and1;
  wire s_wallace_cla8_fa10_or0;
  wire s_wallace_cla8_and_3_2;
  wire s_wallace_cla8_and_2_3;
  wire s_wallace_cla8_fa11_xor0;
  wire s_wallace_cla8_fa11_and0;
  wire s_wallace_cla8_fa11_xor1;
  wire s_wallace_cla8_fa11_and1;
  wire s_wallace_cla8_fa11_or0;
  wire s_wallace_cla8_and_4_2;
  wire s_wallace_cla8_and_3_3;
  wire s_wallace_cla8_fa12_xor0;
  wire s_wallace_cla8_fa12_and0;
  wire s_wallace_cla8_fa12_xor1;
  wire s_wallace_cla8_fa12_and1;
  wire s_wallace_cla8_fa12_or0;
  wire s_wallace_cla8_and_5_2;
  wire s_wallace_cla8_and_4_3;
  wire s_wallace_cla8_fa13_xor0;
  wire s_wallace_cla8_fa13_and0;
  wire s_wallace_cla8_fa13_xor1;
  wire s_wallace_cla8_fa13_and1;
  wire s_wallace_cla8_fa13_or0;
  wire s_wallace_cla8_and_6_2;
  wire s_wallace_cla8_and_5_3;
  wire s_wallace_cla8_fa14_xor0;
  wire s_wallace_cla8_fa14_and0;
  wire s_wallace_cla8_fa14_xor1;
  wire s_wallace_cla8_fa14_and1;
  wire s_wallace_cla8_fa14_or0;
  wire s_wallace_cla8_and_5_4;
  wire s_wallace_cla8_and_4_5;
  wire s_wallace_cla8_fa15_xor0;
  wire s_wallace_cla8_fa15_and0;
  wire s_wallace_cla8_fa15_xor1;
  wire s_wallace_cla8_fa15_and1;
  wire s_wallace_cla8_fa15_or0;
  wire s_wallace_cla8_and_5_5;
  wire s_wallace_cla8_and_4_6;
  wire s_wallace_cla8_fa16_xor0;
  wire s_wallace_cla8_fa16_and0;
  wire s_wallace_cla8_fa16_xor1;
  wire s_wallace_cla8_fa16_and1;
  wire s_wallace_cla8_fa16_or0;
  wire s_wallace_cla8_and_5_6;
  wire s_wallace_cla8_nand_4_7;
  wire s_wallace_cla8_fa17_xor0;
  wire s_wallace_cla8_fa17_and0;
  wire s_wallace_cla8_fa17_xor1;
  wire s_wallace_cla8_fa17_and1;
  wire s_wallace_cla8_fa17_or0;
  wire s_wallace_cla8_and_0_4;
  wire s_wallace_cla8_ha2_xor0;
  wire s_wallace_cla8_ha2_and0;
  wire s_wallace_cla8_and_1_4;
  wire s_wallace_cla8_and_0_5;
  wire s_wallace_cla8_fa18_xor0;
  wire s_wallace_cla8_fa18_and0;
  wire s_wallace_cla8_fa18_xor1;
  wire s_wallace_cla8_fa18_and1;
  wire s_wallace_cla8_fa18_or0;
  wire s_wallace_cla8_and_2_4;
  wire s_wallace_cla8_and_1_5;
  wire s_wallace_cla8_fa19_xor0;
  wire s_wallace_cla8_fa19_and0;
  wire s_wallace_cla8_fa19_xor1;
  wire s_wallace_cla8_fa19_and1;
  wire s_wallace_cla8_fa19_or0;
  wire s_wallace_cla8_and_3_4;
  wire s_wallace_cla8_and_2_5;
  wire s_wallace_cla8_fa20_xor0;
  wire s_wallace_cla8_fa20_and0;
  wire s_wallace_cla8_fa20_xor1;
  wire s_wallace_cla8_fa20_and1;
  wire s_wallace_cla8_fa20_or0;
  wire s_wallace_cla8_and_4_4;
  wire s_wallace_cla8_and_3_5;
  wire s_wallace_cla8_fa21_xor0;
  wire s_wallace_cla8_fa21_and0;
  wire s_wallace_cla8_fa21_xor1;
  wire s_wallace_cla8_fa21_and1;
  wire s_wallace_cla8_fa21_or0;
  wire s_wallace_cla8_and_3_6;
  wire s_wallace_cla8_nand_2_7;
  wire s_wallace_cla8_fa22_xor0;
  wire s_wallace_cla8_fa22_and0;
  wire s_wallace_cla8_fa22_xor1;
  wire s_wallace_cla8_fa22_and1;
  wire s_wallace_cla8_fa22_or0;
  wire s_wallace_cla8_nand_3_7;
  wire s_wallace_cla8_fa23_xor0;
  wire s_wallace_cla8_fa23_and0;
  wire s_wallace_cla8_fa23_xor1;
  wire s_wallace_cla8_fa23_and1;
  wire s_wallace_cla8_fa23_or0;
  wire s_wallace_cla8_ha3_xor0;
  wire s_wallace_cla8_ha3_and0;
  wire s_wallace_cla8_and_0_6;
  wire s_wallace_cla8_fa24_xor0;
  wire s_wallace_cla8_fa24_and0;
  wire s_wallace_cla8_fa24_xor1;
  wire s_wallace_cla8_fa24_and1;
  wire s_wallace_cla8_fa24_or0;
  wire s_wallace_cla8_and_1_6;
  wire s_wallace_cla8_nand_0_7;
  wire s_wallace_cla8_fa25_xor0;
  wire s_wallace_cla8_fa25_and0;
  wire s_wallace_cla8_fa25_xor1;
  wire s_wallace_cla8_fa25_and1;
  wire s_wallace_cla8_fa25_or0;
  wire s_wallace_cla8_and_2_6;
  wire s_wallace_cla8_nand_1_7;
  wire s_wallace_cla8_fa26_xor0;
  wire s_wallace_cla8_fa26_and0;
  wire s_wallace_cla8_fa26_xor1;
  wire s_wallace_cla8_fa26_and1;
  wire s_wallace_cla8_fa26_or0;
  wire s_wallace_cla8_fa27_xor0;
  wire s_wallace_cla8_fa27_and0;
  wire s_wallace_cla8_fa27_xor1;
  wire s_wallace_cla8_fa27_and1;
  wire s_wallace_cla8_fa27_or0;
  wire s_wallace_cla8_ha4_xor0;
  wire s_wallace_cla8_ha4_and0;
  wire s_wallace_cla8_fa28_xor0;
  wire s_wallace_cla8_fa28_and0;
  wire s_wallace_cla8_fa28_xor1;
  wire s_wallace_cla8_fa28_and1;
  wire s_wallace_cla8_fa28_or0;
  wire s_wallace_cla8_fa29_xor0;
  wire s_wallace_cla8_fa29_and0;
  wire s_wallace_cla8_fa29_xor1;
  wire s_wallace_cla8_fa29_and1;
  wire s_wallace_cla8_fa29_or0;
  wire s_wallace_cla8_ha5_xor0;
  wire s_wallace_cla8_ha5_and0;
  wire s_wallace_cla8_fa30_xor0;
  wire s_wallace_cla8_fa30_and0;
  wire s_wallace_cla8_fa30_xor1;
  wire s_wallace_cla8_fa30_and1;
  wire s_wallace_cla8_fa30_or0;
  wire s_wallace_cla8_fa31_xor0;
  wire s_wallace_cla8_fa31_and0;
  wire s_wallace_cla8_fa31_xor1;
  wire s_wallace_cla8_fa31_and1;
  wire s_wallace_cla8_fa31_or0;
  wire s_wallace_cla8_fa32_xor0;
  wire s_wallace_cla8_fa32_and0;
  wire s_wallace_cla8_fa32_xor1;
  wire s_wallace_cla8_fa32_and1;
  wire s_wallace_cla8_fa32_or0;
  wire s_wallace_cla8_fa33_xor0;
  wire s_wallace_cla8_fa33_and0;
  wire s_wallace_cla8_fa33_xor1;
  wire s_wallace_cla8_fa33_and1;
  wire s_wallace_cla8_fa33_or0;
  wire s_wallace_cla8_nand_5_7;
  wire s_wallace_cla8_fa34_xor0;
  wire s_wallace_cla8_fa34_and0;
  wire s_wallace_cla8_fa34_xor1;
  wire s_wallace_cla8_fa34_and1;
  wire s_wallace_cla8_fa34_or0;
  wire s_wallace_cla8_nand_7_6;
  wire s_wallace_cla8_fa35_xor0;
  wire s_wallace_cla8_fa35_and0;
  wire s_wallace_cla8_fa35_xor1;
  wire s_wallace_cla8_fa35_and1;
  wire s_wallace_cla8_fa35_or0;
  wire s_wallace_cla8_and_0_0;
  wire s_wallace_cla8_and_1_0;
  wire s_wallace_cla8_and_0_2;
  wire s_wallace_cla8_nand_6_7;
  wire s_wallace_cla8_and_0_1;
  wire s_wallace_cla8_and_7_7;
  wire s_wallace_cla8_u_cla14_pg_logic0_or0;
  wire s_wallace_cla8_u_cla14_pg_logic0_and0;
  wire s_wallace_cla8_u_cla14_pg_logic0_xor0;
  wire s_wallace_cla8_u_cla14_pg_logic1_or0;
  wire s_wallace_cla8_u_cla14_pg_logic1_and0;
  wire s_wallace_cla8_u_cla14_pg_logic1_xor0;
  wire s_wallace_cla8_u_cla14_xor1;
  wire s_wallace_cla8_u_cla14_and0;
  wire s_wallace_cla8_u_cla14_or0;
  wire s_wallace_cla8_u_cla14_pg_logic2_or0;
  wire s_wallace_cla8_u_cla14_pg_logic2_and0;
  wire s_wallace_cla8_u_cla14_pg_logic2_xor0;
  wire s_wallace_cla8_u_cla14_xor2;
  wire s_wallace_cla8_u_cla14_and1;
  wire s_wallace_cla8_u_cla14_and2;
  wire s_wallace_cla8_u_cla14_and3;
  wire s_wallace_cla8_u_cla14_and4;
  wire s_wallace_cla8_u_cla14_or1;
  wire s_wallace_cla8_u_cla14_or2;
  wire s_wallace_cla8_u_cla14_pg_logic3_or0;
  wire s_wallace_cla8_u_cla14_pg_logic3_and0;
  wire s_wallace_cla8_u_cla14_pg_logic3_xor0;
  wire s_wallace_cla8_u_cla14_xor3;
  wire s_wallace_cla8_u_cla14_and5;
  wire s_wallace_cla8_u_cla14_and6;
  wire s_wallace_cla8_u_cla14_and7;
  wire s_wallace_cla8_u_cla14_and8;
  wire s_wallace_cla8_u_cla14_and9;
  wire s_wallace_cla8_u_cla14_and10;
  wire s_wallace_cla8_u_cla14_and11;
  wire s_wallace_cla8_u_cla14_or3;
  wire s_wallace_cla8_u_cla14_or4;
  wire s_wallace_cla8_u_cla14_or5;
  wire s_wallace_cla8_u_cla14_pg_logic4_or0;
  wire s_wallace_cla8_u_cla14_pg_logic4_and0;
  wire s_wallace_cla8_u_cla14_pg_logic4_xor0;
  wire s_wallace_cla8_u_cla14_xor4;
  wire s_wallace_cla8_u_cla14_and12;
  wire s_wallace_cla8_u_cla14_or6;
  wire s_wallace_cla8_u_cla14_pg_logic5_or0;
  wire s_wallace_cla8_u_cla14_pg_logic5_and0;
  wire s_wallace_cla8_u_cla14_pg_logic5_xor0;
  wire s_wallace_cla8_u_cla14_xor5;
  wire s_wallace_cla8_u_cla14_and13;
  wire s_wallace_cla8_u_cla14_and14;
  wire s_wallace_cla8_u_cla14_and15;
  wire s_wallace_cla8_u_cla14_or7;
  wire s_wallace_cla8_u_cla14_or8;
  wire s_wallace_cla8_u_cla14_pg_logic6_or0;
  wire s_wallace_cla8_u_cla14_pg_logic6_and0;
  wire s_wallace_cla8_u_cla14_pg_logic6_xor0;
  wire s_wallace_cla8_u_cla14_xor6;
  wire s_wallace_cla8_u_cla14_and16;
  wire s_wallace_cla8_u_cla14_and17;
  wire s_wallace_cla8_u_cla14_and18;
  wire s_wallace_cla8_u_cla14_and19;
  wire s_wallace_cla8_u_cla14_and20;
  wire s_wallace_cla8_u_cla14_and21;
  wire s_wallace_cla8_u_cla14_or9;
  wire s_wallace_cla8_u_cla14_or10;
  wire s_wallace_cla8_u_cla14_or11;
  wire s_wallace_cla8_u_cla14_pg_logic7_or0;
  wire s_wallace_cla8_u_cla14_pg_logic7_and0;
  wire s_wallace_cla8_u_cla14_pg_logic7_xor0;
  wire s_wallace_cla8_u_cla14_xor7;
  wire s_wallace_cla8_u_cla14_and22;
  wire s_wallace_cla8_u_cla14_and23;
  wire s_wallace_cla8_u_cla14_and24;
  wire s_wallace_cla8_u_cla14_and25;
  wire s_wallace_cla8_u_cla14_and26;
  wire s_wallace_cla8_u_cla14_and27;
  wire s_wallace_cla8_u_cla14_and28;
  wire s_wallace_cla8_u_cla14_and29;
  wire s_wallace_cla8_u_cla14_and30;
  wire s_wallace_cla8_u_cla14_and31;
  wire s_wallace_cla8_u_cla14_or12;
  wire s_wallace_cla8_u_cla14_or13;
  wire s_wallace_cla8_u_cla14_or14;
  wire s_wallace_cla8_u_cla14_or15;
  wire s_wallace_cla8_u_cla14_pg_logic8_or0;
  wire s_wallace_cla8_u_cla14_pg_logic8_and0;
  wire s_wallace_cla8_u_cla14_pg_logic8_xor0;
  wire s_wallace_cla8_u_cla14_xor8;
  wire s_wallace_cla8_u_cla14_and32;
  wire s_wallace_cla8_u_cla14_or16;
  wire s_wallace_cla8_u_cla14_pg_logic9_or0;
  wire s_wallace_cla8_u_cla14_pg_logic9_and0;
  wire s_wallace_cla8_u_cla14_pg_logic9_xor0;
  wire s_wallace_cla8_u_cla14_xor9;
  wire s_wallace_cla8_u_cla14_and33;
  wire s_wallace_cla8_u_cla14_and34;
  wire s_wallace_cla8_u_cla14_and35;
  wire s_wallace_cla8_u_cla14_or17;
  wire s_wallace_cla8_u_cla14_or18;
  wire s_wallace_cla8_u_cla14_pg_logic10_or0;
  wire s_wallace_cla8_u_cla14_pg_logic10_and0;
  wire s_wallace_cla8_u_cla14_pg_logic10_xor0;
  wire s_wallace_cla8_u_cla14_xor10;
  wire s_wallace_cla8_u_cla14_and36;
  wire s_wallace_cla8_u_cla14_and37;
  wire s_wallace_cla8_u_cla14_and38;
  wire s_wallace_cla8_u_cla14_and39;
  wire s_wallace_cla8_u_cla14_and40;
  wire s_wallace_cla8_u_cla14_and41;
  wire s_wallace_cla8_u_cla14_or19;
  wire s_wallace_cla8_u_cla14_or20;
  wire s_wallace_cla8_u_cla14_or21;
  wire s_wallace_cla8_u_cla14_pg_logic11_or0;
  wire s_wallace_cla8_u_cla14_pg_logic11_and0;
  wire s_wallace_cla8_u_cla14_pg_logic11_xor0;
  wire s_wallace_cla8_u_cla14_xor11;
  wire s_wallace_cla8_u_cla14_and42;
  wire s_wallace_cla8_u_cla14_and43;
  wire s_wallace_cla8_u_cla14_and44;
  wire s_wallace_cla8_u_cla14_and45;
  wire s_wallace_cla8_u_cla14_and46;
  wire s_wallace_cla8_u_cla14_and47;
  wire s_wallace_cla8_u_cla14_and48;
  wire s_wallace_cla8_u_cla14_and49;
  wire s_wallace_cla8_u_cla14_and50;
  wire s_wallace_cla8_u_cla14_and51;
  wire s_wallace_cla8_u_cla14_or22;
  wire s_wallace_cla8_u_cla14_or23;
  wire s_wallace_cla8_u_cla14_or24;
  wire s_wallace_cla8_u_cla14_or25;
  wire s_wallace_cla8_u_cla14_pg_logic12_or0;
  wire s_wallace_cla8_u_cla14_pg_logic12_and0;
  wire s_wallace_cla8_u_cla14_pg_logic12_xor0;
  wire s_wallace_cla8_u_cla14_xor12;
  wire s_wallace_cla8_u_cla14_and52;
  wire s_wallace_cla8_u_cla14_or26;
  wire s_wallace_cla8_u_cla14_pg_logic13_or0;
  wire s_wallace_cla8_u_cla14_pg_logic13_and0;
  wire s_wallace_cla8_u_cla14_pg_logic13_xor0;
  wire s_wallace_cla8_u_cla14_xor13;
  wire s_wallace_cla8_u_cla14_and53;
  wire s_wallace_cla8_u_cla14_and54;
  wire s_wallace_cla8_u_cla14_and55;
  wire s_wallace_cla8_u_cla14_or27;
  wire s_wallace_cla8_u_cla14_or28;
  wire s_wallace_cla8_xor0;

  assign s_wallace_cla8_and_2_0 = a[2] & b[0];
  assign s_wallace_cla8_and_1_1 = a[1] & b[1];
  assign s_wallace_cla8_ha0_xor0 = s_wallace_cla8_and_2_0 ^ s_wallace_cla8_and_1_1;
  assign s_wallace_cla8_ha0_and0 = s_wallace_cla8_and_2_0 & s_wallace_cla8_and_1_1;
  assign s_wallace_cla8_and_3_0 = a[3] & b[0];
  assign s_wallace_cla8_and_2_1 = a[2] & b[1];
  assign s_wallace_cla8_fa0_xor0 = s_wallace_cla8_ha0_and0 ^ s_wallace_cla8_and_3_0;
  assign s_wallace_cla8_fa0_and0 = s_wallace_cla8_ha0_and0 & s_wallace_cla8_and_3_0;
  assign s_wallace_cla8_fa0_xor1 = s_wallace_cla8_fa0_xor0 ^ s_wallace_cla8_and_2_1;
  assign s_wallace_cla8_fa0_and1 = s_wallace_cla8_fa0_xor0 & s_wallace_cla8_and_2_1;
  assign s_wallace_cla8_fa0_or0 = s_wallace_cla8_fa0_and0 | s_wallace_cla8_fa0_and1;
  assign s_wallace_cla8_and_4_0 = a[4] & b[0];
  assign s_wallace_cla8_and_3_1 = a[3] & b[1];
  assign s_wallace_cla8_fa1_xor0 = s_wallace_cla8_fa0_or0 ^ s_wallace_cla8_and_4_0;
  assign s_wallace_cla8_fa1_and0 = s_wallace_cla8_fa0_or0 & s_wallace_cla8_and_4_0;
  assign s_wallace_cla8_fa1_xor1 = s_wallace_cla8_fa1_xor0 ^ s_wallace_cla8_and_3_1;
  assign s_wallace_cla8_fa1_and1 = s_wallace_cla8_fa1_xor0 & s_wallace_cla8_and_3_1;
  assign s_wallace_cla8_fa1_or0 = s_wallace_cla8_fa1_and0 | s_wallace_cla8_fa1_and1;
  assign s_wallace_cla8_and_5_0 = a[5] & b[0];
  assign s_wallace_cla8_and_4_1 = a[4] & b[1];
  assign s_wallace_cla8_fa2_xor0 = s_wallace_cla8_fa1_or0 ^ s_wallace_cla8_and_5_0;
  assign s_wallace_cla8_fa2_and0 = s_wallace_cla8_fa1_or0 & s_wallace_cla8_and_5_0;
  assign s_wallace_cla8_fa2_xor1 = s_wallace_cla8_fa2_xor0 ^ s_wallace_cla8_and_4_1;
  assign s_wallace_cla8_fa2_and1 = s_wallace_cla8_fa2_xor0 & s_wallace_cla8_and_4_1;
  assign s_wallace_cla8_fa2_or0 = s_wallace_cla8_fa2_and0 | s_wallace_cla8_fa2_and1;
  assign s_wallace_cla8_and_6_0 = a[6] & b[0];
  assign s_wallace_cla8_and_5_1 = a[5] & b[1];
  assign s_wallace_cla8_fa3_xor0 = s_wallace_cla8_fa2_or0 ^ s_wallace_cla8_and_6_0;
  assign s_wallace_cla8_fa3_and0 = s_wallace_cla8_fa2_or0 & s_wallace_cla8_and_6_0;
  assign s_wallace_cla8_fa3_xor1 = s_wallace_cla8_fa3_xor0 ^ s_wallace_cla8_and_5_1;
  assign s_wallace_cla8_fa3_and1 = s_wallace_cla8_fa3_xor0 & s_wallace_cla8_and_5_1;
  assign s_wallace_cla8_fa3_or0 = s_wallace_cla8_fa3_and0 | s_wallace_cla8_fa3_and1;
  assign s_wallace_cla8_nand_7_0 = ~(a[7] & b[0]);
  assign s_wallace_cla8_and_6_1 = a[6] & b[1];
  assign s_wallace_cla8_fa4_xor0 = s_wallace_cla8_fa3_or0 ^ s_wallace_cla8_nand_7_0;
  assign s_wallace_cla8_fa4_and0 = s_wallace_cla8_fa3_or0 & s_wallace_cla8_nand_7_0;
  assign s_wallace_cla8_fa4_xor1 = s_wallace_cla8_fa4_xor0 ^ s_wallace_cla8_and_6_1;
  assign s_wallace_cla8_fa4_and1 = s_wallace_cla8_fa4_xor0 & s_wallace_cla8_and_6_1;
  assign s_wallace_cla8_fa4_or0 = s_wallace_cla8_fa4_and0 | s_wallace_cla8_fa4_and1;
  assign s_wallace_cla8_nand_7_1 = ~(a[7] & b[1]);
  assign s_wallace_cla8_fa5_xor0 = ~s_wallace_cla8_fa4_or0;
  assign s_wallace_cla8_fa5_xor1 = s_wallace_cla8_fa5_xor0 ^ s_wallace_cla8_nand_7_1;
  assign s_wallace_cla8_fa5_and1 = s_wallace_cla8_fa5_xor0 & s_wallace_cla8_nand_7_1;
  assign s_wallace_cla8_fa5_or0 = s_wallace_cla8_fa4_or0 | s_wallace_cla8_fa5_and1;
  assign s_wallace_cla8_nand_7_2 = ~(a[7] & b[2]);
  assign s_wallace_cla8_and_6_3 = a[6] & b[3];
  assign s_wallace_cla8_fa6_xor0 = s_wallace_cla8_fa5_or0 ^ s_wallace_cla8_nand_7_2;
  assign s_wallace_cla8_fa6_and0 = s_wallace_cla8_fa5_or0 & s_wallace_cla8_nand_7_2;
  assign s_wallace_cla8_fa6_xor1 = s_wallace_cla8_fa6_xor0 ^ s_wallace_cla8_and_6_3;
  assign s_wallace_cla8_fa6_and1 = s_wallace_cla8_fa6_xor0 & s_wallace_cla8_and_6_3;
  assign s_wallace_cla8_fa6_or0 = s_wallace_cla8_fa6_and0 | s_wallace_cla8_fa6_and1;
  assign s_wallace_cla8_nand_7_3 = ~(a[7] & b[3]);
  assign s_wallace_cla8_and_6_4 = a[6] & b[4];
  assign s_wallace_cla8_fa7_xor0 = s_wallace_cla8_fa6_or0 ^ s_wallace_cla8_nand_7_3;
  assign s_wallace_cla8_fa7_and0 = s_wallace_cla8_fa6_or0 & s_wallace_cla8_nand_7_3;
  assign s_wallace_cla8_fa7_xor1 = s_wallace_cla8_fa7_xor0 ^ s_wallace_cla8_and_6_4;
  assign s_wallace_cla8_fa7_and1 = s_wallace_cla8_fa7_xor0 & s_wallace_cla8_and_6_4;
  assign s_wallace_cla8_fa7_or0 = s_wallace_cla8_fa7_and0 | s_wallace_cla8_fa7_and1;
  assign s_wallace_cla8_nand_7_4 = ~(a[7] & b[4]);
  assign s_wallace_cla8_and_6_5 = a[6] & b[5];
  assign s_wallace_cla8_fa8_xor0 = s_wallace_cla8_fa7_or0 ^ s_wallace_cla8_nand_7_4;
  assign s_wallace_cla8_fa8_and0 = s_wallace_cla8_fa7_or0 & s_wallace_cla8_nand_7_4;
  assign s_wallace_cla8_fa8_xor1 = s_wallace_cla8_fa8_xor0 ^ s_wallace_cla8_and_6_5;
  assign s_wallace_cla8_fa8_and1 = s_wallace_cla8_fa8_xor0 & s_wallace_cla8_and_6_5;
  assign s_wallace_cla8_fa8_or0 = s_wallace_cla8_fa8_and0 | s_wallace_cla8_fa8_and1;
  assign s_wallace_cla8_nand_7_5 = ~(a[7] & b[5]);
  assign s_wallace_cla8_and_6_6 = a[6] & b[6];
  assign s_wallace_cla8_fa9_xor0 = s_wallace_cla8_fa8_or0 ^ s_wallace_cla8_nand_7_5;
  assign s_wallace_cla8_fa9_and0 = s_wallace_cla8_fa8_or0 & s_wallace_cla8_nand_7_5;
  assign s_wallace_cla8_fa9_xor1 = s_wallace_cla8_fa9_xor0 ^ s_wallace_cla8_and_6_6;
  assign s_wallace_cla8_fa9_and1 = s_wallace_cla8_fa9_xor0 & s_wallace_cla8_and_6_6;
  assign s_wallace_cla8_fa9_or0 = s_wallace_cla8_fa9_and0 | s_wallace_cla8_fa9_and1;
  assign s_wallace_cla8_and_1_2 = a[1] & b[2];
  assign s_wallace_cla8_and_0_3 = a[0] & b[3];
  assign s_wallace_cla8_ha1_xor0 = s_wallace_cla8_and_1_2 ^ s_wallace_cla8_and_0_3;
  assign s_wallace_cla8_ha1_and0 = s_wallace_cla8_and_1_2 & s_wallace_cla8_and_0_3;
  assign s_wallace_cla8_and_2_2 = a[2] & b[2];
  assign s_wallace_cla8_and_1_3 = a[1] & b[3];
  assign s_wallace_cla8_fa10_xor0 = s_wallace_cla8_ha1_and0 ^ s_wallace_cla8_and_2_2;
  assign s_wallace_cla8_fa10_and0 = s_wallace_cla8_ha1_and0 & s_wallace_cla8_and_2_2;
  assign s_wallace_cla8_fa10_xor1 = s_wallace_cla8_fa10_xor0 ^ s_wallace_cla8_and_1_3;
  assign s_wallace_cla8_fa10_and1 = s_wallace_cla8_fa10_xor0 & s_wallace_cla8_and_1_3;
  assign s_wallace_cla8_fa10_or0 = s_wallace_cla8_fa10_and0 | s_wallace_cla8_fa10_and1;
  assign s_wallace_cla8_and_3_2 = a[3] & b[2];
  assign s_wallace_cla8_and_2_3 = a[2] & b[3];
  assign s_wallace_cla8_fa11_xor0 = s_wallace_cla8_fa10_or0 ^ s_wallace_cla8_and_3_2;
  assign s_wallace_cla8_fa11_and0 = s_wallace_cla8_fa10_or0 & s_wallace_cla8_and_3_2;
  assign s_wallace_cla8_fa11_xor1 = s_wallace_cla8_fa11_xor0 ^ s_wallace_cla8_and_2_3;
  assign s_wallace_cla8_fa11_and1 = s_wallace_cla8_fa11_xor0 & s_wallace_cla8_and_2_3;
  assign s_wallace_cla8_fa11_or0 = s_wallace_cla8_fa11_and0 | s_wallace_cla8_fa11_and1;
  assign s_wallace_cla8_and_4_2 = a[4] & b[2];
  assign s_wallace_cla8_and_3_3 = a[3] & b[3];
  assign s_wallace_cla8_fa12_xor0 = s_wallace_cla8_fa11_or0 ^ s_wallace_cla8_and_4_2;
  assign s_wallace_cla8_fa12_and0 = s_wallace_cla8_fa11_or0 & s_wallace_cla8_and_4_2;
  assign s_wallace_cla8_fa12_xor1 = s_wallace_cla8_fa12_xor0 ^ s_wallace_cla8_and_3_3;
  assign s_wallace_cla8_fa12_and1 = s_wallace_cla8_fa12_xor0 & s_wallace_cla8_and_3_3;
  assign s_wallace_cla8_fa12_or0 = s_wallace_cla8_fa12_and0 | s_wallace_cla8_fa12_and1;
  assign s_wallace_cla8_and_5_2 = a[5] & b[2];
  assign s_wallace_cla8_and_4_3 = a[4] & b[3];
  assign s_wallace_cla8_fa13_xor0 = s_wallace_cla8_fa12_or0 ^ s_wallace_cla8_and_5_2;
  assign s_wallace_cla8_fa13_and0 = s_wallace_cla8_fa12_or0 & s_wallace_cla8_and_5_2;
  assign s_wallace_cla8_fa13_xor1 = s_wallace_cla8_fa13_xor0 ^ s_wallace_cla8_and_4_3;
  assign s_wallace_cla8_fa13_and1 = s_wallace_cla8_fa13_xor0 & s_wallace_cla8_and_4_3;
  assign s_wallace_cla8_fa13_or0 = s_wallace_cla8_fa13_and0 | s_wallace_cla8_fa13_and1;
  assign s_wallace_cla8_and_6_2 = a[6] & b[2];
  assign s_wallace_cla8_and_5_3 = a[5] & b[3];
  assign s_wallace_cla8_fa14_xor0 = s_wallace_cla8_fa13_or0 ^ s_wallace_cla8_and_6_2;
  assign s_wallace_cla8_fa14_and0 = s_wallace_cla8_fa13_or0 & s_wallace_cla8_and_6_2;
  assign s_wallace_cla8_fa14_xor1 = s_wallace_cla8_fa14_xor0 ^ s_wallace_cla8_and_5_3;
  assign s_wallace_cla8_fa14_and1 = s_wallace_cla8_fa14_xor0 & s_wallace_cla8_and_5_3;
  assign s_wallace_cla8_fa14_or0 = s_wallace_cla8_fa14_and0 | s_wallace_cla8_fa14_and1;
  assign s_wallace_cla8_and_5_4 = a[5] & b[4];
  assign s_wallace_cla8_and_4_5 = a[4] & b[5];
  assign s_wallace_cla8_fa15_xor0 = s_wallace_cla8_fa14_or0 ^ s_wallace_cla8_and_5_4;
  assign s_wallace_cla8_fa15_and0 = s_wallace_cla8_fa14_or0 & s_wallace_cla8_and_5_4;
  assign s_wallace_cla8_fa15_xor1 = s_wallace_cla8_fa15_xor0 ^ s_wallace_cla8_and_4_5;
  assign s_wallace_cla8_fa15_and1 = s_wallace_cla8_fa15_xor0 & s_wallace_cla8_and_4_5;
  assign s_wallace_cla8_fa15_or0 = s_wallace_cla8_fa15_and0 | s_wallace_cla8_fa15_and1;
  assign s_wallace_cla8_and_5_5 = a[5] & b[5];
  assign s_wallace_cla8_and_4_6 = a[4] & b[6];
  assign s_wallace_cla8_fa16_xor0 = s_wallace_cla8_fa15_or0 ^ s_wallace_cla8_and_5_5;
  assign s_wallace_cla8_fa16_and0 = s_wallace_cla8_fa15_or0 & s_wallace_cla8_and_5_5;
  assign s_wallace_cla8_fa16_xor1 = s_wallace_cla8_fa16_xor0 ^ s_wallace_cla8_and_4_6;
  assign s_wallace_cla8_fa16_and1 = s_wallace_cla8_fa16_xor0 & s_wallace_cla8_and_4_6;
  assign s_wallace_cla8_fa16_or0 = s_wallace_cla8_fa16_and0 | s_wallace_cla8_fa16_and1;
  assign s_wallace_cla8_and_5_6 = a[5] & b[6];
  assign s_wallace_cla8_nand_4_7 = ~(a[4] & b[7]);
  assign s_wallace_cla8_fa17_xor0 = s_wallace_cla8_fa16_or0 ^ s_wallace_cla8_and_5_6;
  assign s_wallace_cla8_fa17_and0 = s_wallace_cla8_fa16_or0 & s_wallace_cla8_and_5_6;
  assign s_wallace_cla8_fa17_xor1 = s_wallace_cla8_fa17_xor0 ^ s_wallace_cla8_nand_4_7;
  assign s_wallace_cla8_fa17_and1 = s_wallace_cla8_fa17_xor0 & s_wallace_cla8_nand_4_7;
  assign s_wallace_cla8_fa17_or0 = s_wallace_cla8_fa17_and0 | s_wallace_cla8_fa17_and1;
  assign s_wallace_cla8_and_0_4 = a[0] & b[4];
  assign s_wallace_cla8_ha2_xor0 = s_wallace_cla8_and_0_4 ^ s_wallace_cla8_fa1_xor1;
  assign s_wallace_cla8_ha2_and0 = s_wallace_cla8_and_0_4 & s_wallace_cla8_fa1_xor1;
  assign s_wallace_cla8_and_1_4 = a[1] & b[4];
  assign s_wallace_cla8_and_0_5 = a[0] & b[5];
  assign s_wallace_cla8_fa18_xor0 = s_wallace_cla8_ha2_and0 ^ s_wallace_cla8_and_1_4;
  assign s_wallace_cla8_fa18_and0 = s_wallace_cla8_ha2_and0 & s_wallace_cla8_and_1_4;
  assign s_wallace_cla8_fa18_xor1 = s_wallace_cla8_fa18_xor0 ^ s_wallace_cla8_and_0_5;
  assign s_wallace_cla8_fa18_and1 = s_wallace_cla8_fa18_xor0 & s_wallace_cla8_and_0_5;
  assign s_wallace_cla8_fa18_or0 = s_wallace_cla8_fa18_and0 | s_wallace_cla8_fa18_and1;
  assign s_wallace_cla8_and_2_4 = a[2] & b[4];
  assign s_wallace_cla8_and_1_5 = a[1] & b[5];
  assign s_wallace_cla8_fa19_xor0 = s_wallace_cla8_fa18_or0 ^ s_wallace_cla8_and_2_4;
  assign s_wallace_cla8_fa19_and0 = s_wallace_cla8_fa18_or0 & s_wallace_cla8_and_2_4;
  assign s_wallace_cla8_fa19_xor1 = s_wallace_cla8_fa19_xor0 ^ s_wallace_cla8_and_1_5;
  assign s_wallace_cla8_fa19_and1 = s_wallace_cla8_fa19_xor0 & s_wallace_cla8_and_1_5;
  assign s_wallace_cla8_fa19_or0 = s_wallace_cla8_fa19_and0 | s_wallace_cla8_fa19_and1;
  assign s_wallace_cla8_and_3_4 = a[3] & b[4];
  assign s_wallace_cla8_and_2_5 = a[2] & b[5];
  assign s_wallace_cla8_fa20_xor0 = s_wallace_cla8_fa19_or0 ^ s_wallace_cla8_and_3_4;
  assign s_wallace_cla8_fa20_and0 = s_wallace_cla8_fa19_or0 & s_wallace_cla8_and_3_4;
  assign s_wallace_cla8_fa20_xor1 = s_wallace_cla8_fa20_xor0 ^ s_wallace_cla8_and_2_5;
  assign s_wallace_cla8_fa20_and1 = s_wallace_cla8_fa20_xor0 & s_wallace_cla8_and_2_5;
  assign s_wallace_cla8_fa20_or0 = s_wallace_cla8_fa20_and0 | s_wallace_cla8_fa20_and1;
  assign s_wallace_cla8_and_4_4 = a[4] & b[4];
  assign s_wallace_cla8_and_3_5 = a[3] & b[5];
  assign s_wallace_cla8_fa21_xor0 = s_wallace_cla8_fa20_or0 ^ s_wallace_cla8_and_4_4;
  assign s_wallace_cla8_fa21_and0 = s_wallace_cla8_fa20_or0 & s_wallace_cla8_and_4_4;
  assign s_wallace_cla8_fa21_xor1 = s_wallace_cla8_fa21_xor0 ^ s_wallace_cla8_and_3_5;
  assign s_wallace_cla8_fa21_and1 = s_wallace_cla8_fa21_xor0 & s_wallace_cla8_and_3_5;
  assign s_wallace_cla8_fa21_or0 = s_wallace_cla8_fa21_and0 | s_wallace_cla8_fa21_and1;
  assign s_wallace_cla8_and_3_6 = a[3] & b[6];
  assign s_wallace_cla8_nand_2_7 = ~(a[2] & b[7]);
  assign s_wallace_cla8_fa22_xor0 = s_wallace_cla8_fa21_or0 ^ s_wallace_cla8_and_3_6;
  assign s_wallace_cla8_fa22_and0 = s_wallace_cla8_fa21_or0 & s_wallace_cla8_and_3_6;
  assign s_wallace_cla8_fa22_xor1 = s_wallace_cla8_fa22_xor0 ^ s_wallace_cla8_nand_2_7;
  assign s_wallace_cla8_fa22_and1 = s_wallace_cla8_fa22_xor0 & s_wallace_cla8_nand_2_7;
  assign s_wallace_cla8_fa22_or0 = s_wallace_cla8_fa22_and0 | s_wallace_cla8_fa22_and1;
  assign s_wallace_cla8_nand_3_7 = ~(a[3] & b[7]);
  assign s_wallace_cla8_fa23_xor0 = s_wallace_cla8_fa22_or0 ^ s_wallace_cla8_nand_3_7;
  assign s_wallace_cla8_fa23_and0 = s_wallace_cla8_fa22_or0 & s_wallace_cla8_nand_3_7;
  assign s_wallace_cla8_fa23_xor1 = s_wallace_cla8_fa23_xor0 ^ s_wallace_cla8_fa7_xor1;
  assign s_wallace_cla8_fa23_and1 = s_wallace_cla8_fa23_xor0 & s_wallace_cla8_fa7_xor1;
  assign s_wallace_cla8_fa23_or0 = s_wallace_cla8_fa23_and0 | s_wallace_cla8_fa23_and1;
  assign s_wallace_cla8_ha3_xor0 = s_wallace_cla8_fa2_xor1 ^ s_wallace_cla8_fa11_xor1;
  assign s_wallace_cla8_ha3_and0 = s_wallace_cla8_fa2_xor1 & s_wallace_cla8_fa11_xor1;
  assign s_wallace_cla8_and_0_6 = a[0] & b[6];
  assign s_wallace_cla8_fa24_xor0 = s_wallace_cla8_ha3_and0 ^ s_wallace_cla8_and_0_6;
  assign s_wallace_cla8_fa24_and0 = s_wallace_cla8_ha3_and0 & s_wallace_cla8_and_0_6;
  assign s_wallace_cla8_fa24_xor1 = s_wallace_cla8_fa24_xor0 ^ s_wallace_cla8_fa3_xor1;
  assign s_wallace_cla8_fa24_and1 = s_wallace_cla8_fa24_xor0 & s_wallace_cla8_fa3_xor1;
  assign s_wallace_cla8_fa24_or0 = s_wallace_cla8_fa24_and0 | s_wallace_cla8_fa24_and1;
  assign s_wallace_cla8_and_1_6 = a[1] & b[6];
  assign s_wallace_cla8_nand_0_7 = ~(a[0] & b[7]);
  assign s_wallace_cla8_fa25_xor0 = s_wallace_cla8_fa24_or0 ^ s_wallace_cla8_and_1_6;
  assign s_wallace_cla8_fa25_and0 = s_wallace_cla8_fa24_or0 & s_wallace_cla8_and_1_6;
  assign s_wallace_cla8_fa25_xor1 = s_wallace_cla8_fa25_xor0 ^ s_wallace_cla8_nand_0_7;
  assign s_wallace_cla8_fa25_and1 = s_wallace_cla8_fa25_xor0 & s_wallace_cla8_nand_0_7;
  assign s_wallace_cla8_fa25_or0 = s_wallace_cla8_fa25_and0 | s_wallace_cla8_fa25_and1;
  assign s_wallace_cla8_and_2_6 = a[2] & b[6];
  assign s_wallace_cla8_nand_1_7 = ~(a[1] & b[7]);
  assign s_wallace_cla8_fa26_xor0 = s_wallace_cla8_fa25_or0 ^ s_wallace_cla8_and_2_6;
  assign s_wallace_cla8_fa26_and0 = s_wallace_cla8_fa25_or0 & s_wallace_cla8_and_2_6;
  assign s_wallace_cla8_fa26_xor1 = s_wallace_cla8_fa26_xor0 ^ s_wallace_cla8_nand_1_7;
  assign s_wallace_cla8_fa26_and1 = s_wallace_cla8_fa26_xor0 & s_wallace_cla8_nand_1_7;
  assign s_wallace_cla8_fa26_or0 = s_wallace_cla8_fa26_and0 | s_wallace_cla8_fa26_and1;
  assign s_wallace_cla8_fa27_xor0 = s_wallace_cla8_fa26_or0 ^ s_wallace_cla8_fa6_xor1;
  assign s_wallace_cla8_fa27_and0 = s_wallace_cla8_fa26_or0 & s_wallace_cla8_fa6_xor1;
  assign s_wallace_cla8_fa27_xor1 = s_wallace_cla8_fa27_xor0 ^ s_wallace_cla8_fa15_xor1;
  assign s_wallace_cla8_fa27_and1 = s_wallace_cla8_fa27_xor0 & s_wallace_cla8_fa15_xor1;
  assign s_wallace_cla8_fa27_or0 = s_wallace_cla8_fa27_and0 | s_wallace_cla8_fa27_and1;
  assign s_wallace_cla8_ha4_xor0 = s_wallace_cla8_fa12_xor1 ^ s_wallace_cla8_fa19_xor1;
  assign s_wallace_cla8_ha4_and0 = s_wallace_cla8_fa12_xor1 & s_wallace_cla8_fa19_xor1;
  assign s_wallace_cla8_fa28_xor0 = s_wallace_cla8_ha4_and0 ^ s_wallace_cla8_fa4_xor1;
  assign s_wallace_cla8_fa28_and0 = s_wallace_cla8_ha4_and0 & s_wallace_cla8_fa4_xor1;
  assign s_wallace_cla8_fa28_xor1 = s_wallace_cla8_fa28_xor0 ^ s_wallace_cla8_fa13_xor1;
  assign s_wallace_cla8_fa28_and1 = s_wallace_cla8_fa28_xor0 & s_wallace_cla8_fa13_xor1;
  assign s_wallace_cla8_fa28_or0 = s_wallace_cla8_fa28_and0 | s_wallace_cla8_fa28_and1;
  assign s_wallace_cla8_fa29_xor0 = s_wallace_cla8_fa28_or0 ^ s_wallace_cla8_fa5_xor1;
  assign s_wallace_cla8_fa29_and0 = s_wallace_cla8_fa28_or0 & s_wallace_cla8_fa5_xor1;
  assign s_wallace_cla8_fa29_xor1 = s_wallace_cla8_fa29_xor0 ^ s_wallace_cla8_fa14_xor1;
  assign s_wallace_cla8_fa29_and1 = s_wallace_cla8_fa29_xor0 & s_wallace_cla8_fa14_xor1;
  assign s_wallace_cla8_fa29_or0 = s_wallace_cla8_fa29_and0 | s_wallace_cla8_fa29_and1;
  assign s_wallace_cla8_ha5_xor0 = s_wallace_cla8_fa20_xor1 ^ s_wallace_cla8_fa25_xor1;
  assign s_wallace_cla8_ha5_and0 = s_wallace_cla8_fa20_xor1 & s_wallace_cla8_fa25_xor1;
  assign s_wallace_cla8_fa30_xor0 = s_wallace_cla8_ha5_and0 ^ s_wallace_cla8_fa21_xor1;
  assign s_wallace_cla8_fa30_and0 = s_wallace_cla8_ha5_and0 & s_wallace_cla8_fa21_xor1;
  assign s_wallace_cla8_fa30_xor1 = s_wallace_cla8_fa30_xor0 ^ s_wallace_cla8_fa26_xor1;
  assign s_wallace_cla8_fa30_and1 = s_wallace_cla8_fa30_xor0 & s_wallace_cla8_fa26_xor1;
  assign s_wallace_cla8_fa30_or0 = s_wallace_cla8_fa30_and0 | s_wallace_cla8_fa30_and1;
  assign s_wallace_cla8_fa31_xor0 = s_wallace_cla8_fa30_or0 ^ s_wallace_cla8_fa29_or0;
  assign s_wallace_cla8_fa31_and0 = s_wallace_cla8_fa30_or0 & s_wallace_cla8_fa29_or0;
  assign s_wallace_cla8_fa31_xor1 = s_wallace_cla8_fa31_xor0 ^ s_wallace_cla8_fa22_xor1;
  assign s_wallace_cla8_fa31_and1 = s_wallace_cla8_fa31_xor0 & s_wallace_cla8_fa22_xor1;
  assign s_wallace_cla8_fa31_or0 = s_wallace_cla8_fa31_and0 | s_wallace_cla8_fa31_and1;
  assign s_wallace_cla8_fa32_xor0 = s_wallace_cla8_fa31_or0 ^ s_wallace_cla8_fa27_or0;
  assign s_wallace_cla8_fa32_and0 = s_wallace_cla8_fa31_or0 & s_wallace_cla8_fa27_or0;
  assign s_wallace_cla8_fa32_xor1 = s_wallace_cla8_fa32_xor0 ^ s_wallace_cla8_fa16_xor1;
  assign s_wallace_cla8_fa32_and1 = s_wallace_cla8_fa32_xor0 & s_wallace_cla8_fa16_xor1;
  assign s_wallace_cla8_fa32_or0 = s_wallace_cla8_fa32_and0 | s_wallace_cla8_fa32_and1;
  assign s_wallace_cla8_fa33_xor0 = s_wallace_cla8_fa32_or0 ^ s_wallace_cla8_fa23_or0;
  assign s_wallace_cla8_fa33_and0 = s_wallace_cla8_fa32_or0 & s_wallace_cla8_fa23_or0;
  assign s_wallace_cla8_fa33_xor1 = s_wallace_cla8_fa33_xor0 ^ s_wallace_cla8_fa8_xor1;
  assign s_wallace_cla8_fa33_and1 = s_wallace_cla8_fa33_xor0 & s_wallace_cla8_fa8_xor1;
  assign s_wallace_cla8_fa33_or0 = s_wallace_cla8_fa33_and0 | s_wallace_cla8_fa33_and1;
  assign s_wallace_cla8_nand_5_7 = ~(a[5] & b[7]);
  assign s_wallace_cla8_fa34_xor0 = s_wallace_cla8_fa33_or0 ^ s_wallace_cla8_fa17_or0;
  assign s_wallace_cla8_fa34_and0 = s_wallace_cla8_fa33_or0 & s_wallace_cla8_fa17_or0;
  assign s_wallace_cla8_fa34_xor1 = s_wallace_cla8_fa34_xor0 ^ s_wallace_cla8_nand_5_7;
  assign s_wallace_cla8_fa34_and1 = s_wallace_cla8_fa34_xor0 & s_wallace_cla8_nand_5_7;
  assign s_wallace_cla8_fa34_or0 = s_wallace_cla8_fa34_and0 | s_wallace_cla8_fa34_and1;
  assign s_wallace_cla8_nand_7_6 = ~(a[7] & b[6]);
  assign s_wallace_cla8_fa35_xor0 = s_wallace_cla8_fa34_or0 ^ s_wallace_cla8_fa9_or0;
  assign s_wallace_cla8_fa35_and0 = s_wallace_cla8_fa34_or0 & s_wallace_cla8_fa9_or0;
  assign s_wallace_cla8_fa35_xor1 = s_wallace_cla8_fa35_xor0 ^ s_wallace_cla8_nand_7_6;
  assign s_wallace_cla8_fa35_and1 = s_wallace_cla8_fa35_xor0 & s_wallace_cla8_nand_7_6;
  assign s_wallace_cla8_fa35_or0 = s_wallace_cla8_fa35_and0 | s_wallace_cla8_fa35_and1;
  assign s_wallace_cla8_and_0_0 = a[0] & b[0];
  assign s_wallace_cla8_and_1_0 = a[1] & b[0];
  assign s_wallace_cla8_and_0_2 = a[0] & b[2];
  assign s_wallace_cla8_nand_6_7 = ~(a[6] & b[7]);
  assign s_wallace_cla8_and_0_1 = a[0] & b[1];
  assign s_wallace_cla8_and_7_7 = a[7] & b[7];
  assign s_wallace_cla8_u_cla14_pg_logic0_or0 = s_wallace_cla8_and_1_0 | s_wallace_cla8_and_0_1;
  assign s_wallace_cla8_u_cla14_pg_logic0_and0 = s_wallace_cla8_and_1_0 & s_wallace_cla8_and_0_1;
  assign s_wallace_cla8_u_cla14_pg_logic0_xor0 = s_wallace_cla8_and_1_0 ^ s_wallace_cla8_and_0_1;
  assign s_wallace_cla8_u_cla14_pg_logic1_or0 = s_wallace_cla8_and_0_2 | s_wallace_cla8_ha0_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic1_and0 = s_wallace_cla8_and_0_2 & s_wallace_cla8_ha0_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic1_xor0 = s_wallace_cla8_and_0_2 ^ s_wallace_cla8_ha0_xor0;
  assign s_wallace_cla8_u_cla14_xor1 = s_wallace_cla8_u_cla14_pg_logic1_xor0 ^ s_wallace_cla8_u_cla14_pg_logic0_and0;
  assign s_wallace_cla8_u_cla14_and0 = s_wallace_cla8_u_cla14_pg_logic0_and0 & s_wallace_cla8_u_cla14_pg_logic1_or0;
  assign s_wallace_cla8_u_cla14_or0 = s_wallace_cla8_u_cla14_pg_logic1_and0 | s_wallace_cla8_u_cla14_and0;
  assign s_wallace_cla8_u_cla14_pg_logic2_or0 = s_wallace_cla8_fa0_xor1 | s_wallace_cla8_ha1_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic2_and0 = s_wallace_cla8_fa0_xor1 & s_wallace_cla8_ha1_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic2_xor0 = s_wallace_cla8_fa0_xor1 ^ s_wallace_cla8_ha1_xor0;
  assign s_wallace_cla8_u_cla14_xor2 = s_wallace_cla8_u_cla14_pg_logic2_xor0 ^ s_wallace_cla8_u_cla14_or0;
  assign s_wallace_cla8_u_cla14_and1 = s_wallace_cla8_u_cla14_pg_logic2_or0 & s_wallace_cla8_u_cla14_pg_logic0_or0;
  assign s_wallace_cla8_u_cla14_and2 = s_wallace_cla8_u_cla14_pg_logic0_and0 & s_wallace_cla8_u_cla14_pg_logic2_or0;
  assign s_wallace_cla8_u_cla14_and3 = s_wallace_cla8_u_cla14_and2 & s_wallace_cla8_u_cla14_pg_logic1_or0;
  assign s_wallace_cla8_u_cla14_and4 = s_wallace_cla8_u_cla14_pg_logic1_and0 & s_wallace_cla8_u_cla14_pg_logic2_or0;
  assign s_wallace_cla8_u_cla14_or1 = s_wallace_cla8_u_cla14_and3 | s_wallace_cla8_u_cla14_and4;
  assign s_wallace_cla8_u_cla14_or2 = s_wallace_cla8_u_cla14_pg_logic2_and0 | s_wallace_cla8_u_cla14_or1;
  assign s_wallace_cla8_u_cla14_pg_logic3_or0 = s_wallace_cla8_fa10_xor1 | s_wallace_cla8_ha2_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic3_and0 = s_wallace_cla8_fa10_xor1 & s_wallace_cla8_ha2_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic3_xor0 = s_wallace_cla8_fa10_xor1 ^ s_wallace_cla8_ha2_xor0;
  assign s_wallace_cla8_u_cla14_xor3 = s_wallace_cla8_u_cla14_pg_logic3_xor0 ^ s_wallace_cla8_u_cla14_or2;
  assign s_wallace_cla8_u_cla14_and5 = s_wallace_cla8_u_cla14_pg_logic3_or0 & s_wallace_cla8_u_cla14_pg_logic1_or0;
  assign s_wallace_cla8_u_cla14_and6 = s_wallace_cla8_u_cla14_pg_logic0_and0 & s_wallace_cla8_u_cla14_pg_logic2_or0;
  assign s_wallace_cla8_u_cla14_and7 = s_wallace_cla8_u_cla14_pg_logic3_or0 & s_wallace_cla8_u_cla14_pg_logic1_or0;
  assign s_wallace_cla8_u_cla14_and8 = s_wallace_cla8_u_cla14_and6 & s_wallace_cla8_u_cla14_and7;
  assign s_wallace_cla8_u_cla14_and9 = s_wallace_cla8_u_cla14_pg_logic1_and0 & s_wallace_cla8_u_cla14_pg_logic3_or0;
  assign s_wallace_cla8_u_cla14_and10 = s_wallace_cla8_u_cla14_and9 & s_wallace_cla8_u_cla14_pg_logic2_or0;
  assign s_wallace_cla8_u_cla14_and11 = s_wallace_cla8_u_cla14_pg_logic2_and0 & s_wallace_cla8_u_cla14_pg_logic3_or0;
  assign s_wallace_cla8_u_cla14_or3 = s_wallace_cla8_u_cla14_and8 | s_wallace_cla8_u_cla14_and11;
  assign s_wallace_cla8_u_cla14_or4 = s_wallace_cla8_u_cla14_and10 | s_wallace_cla8_u_cla14_or3;
  assign s_wallace_cla8_u_cla14_or5 = s_wallace_cla8_u_cla14_pg_logic3_and0 | s_wallace_cla8_u_cla14_or4;
  assign s_wallace_cla8_u_cla14_pg_logic4_or0 = s_wallace_cla8_fa18_xor1 | s_wallace_cla8_ha3_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic4_and0 = s_wallace_cla8_fa18_xor1 & s_wallace_cla8_ha3_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic4_xor0 = s_wallace_cla8_fa18_xor1 ^ s_wallace_cla8_ha3_xor0;
  assign s_wallace_cla8_u_cla14_xor4 = s_wallace_cla8_u_cla14_pg_logic4_xor0 ^ s_wallace_cla8_u_cla14_or5;
  assign s_wallace_cla8_u_cla14_and12 = s_wallace_cla8_u_cla14_or5 & s_wallace_cla8_u_cla14_pg_logic4_or0;
  assign s_wallace_cla8_u_cla14_or6 = s_wallace_cla8_u_cla14_pg_logic4_and0 | s_wallace_cla8_u_cla14_and12;
  assign s_wallace_cla8_u_cla14_pg_logic5_or0 = s_wallace_cla8_fa24_xor1 | s_wallace_cla8_ha4_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic5_and0 = s_wallace_cla8_fa24_xor1 & s_wallace_cla8_ha4_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic5_xor0 = s_wallace_cla8_fa24_xor1 ^ s_wallace_cla8_ha4_xor0;
  assign s_wallace_cla8_u_cla14_xor5 = s_wallace_cla8_u_cla14_pg_logic5_xor0 ^ s_wallace_cla8_u_cla14_or6;
  assign s_wallace_cla8_u_cla14_and13 = s_wallace_cla8_u_cla14_or5 & s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign s_wallace_cla8_u_cla14_and14 = s_wallace_cla8_u_cla14_and13 & s_wallace_cla8_u_cla14_pg_logic4_or0;
  assign s_wallace_cla8_u_cla14_and15 = s_wallace_cla8_u_cla14_pg_logic4_and0 & s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign s_wallace_cla8_u_cla14_or7 = s_wallace_cla8_u_cla14_and14 | s_wallace_cla8_u_cla14_and15;
  assign s_wallace_cla8_u_cla14_or8 = s_wallace_cla8_u_cla14_pg_logic5_and0 | s_wallace_cla8_u_cla14_or7;
  assign s_wallace_cla8_u_cla14_pg_logic6_or0 = s_wallace_cla8_fa28_xor1 | s_wallace_cla8_ha5_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic6_and0 = s_wallace_cla8_fa28_xor1 & s_wallace_cla8_ha5_xor0;
  assign s_wallace_cla8_u_cla14_pg_logic6_xor0 = s_wallace_cla8_fa28_xor1 ^ s_wallace_cla8_ha5_xor0;
  assign s_wallace_cla8_u_cla14_xor6 = s_wallace_cla8_u_cla14_pg_logic6_xor0 ^ s_wallace_cla8_u_cla14_or8;
  assign s_wallace_cla8_u_cla14_and16 = s_wallace_cla8_u_cla14_or5 & s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign s_wallace_cla8_u_cla14_and17 = s_wallace_cla8_u_cla14_pg_logic6_or0 & s_wallace_cla8_u_cla14_pg_logic4_or0;
  assign s_wallace_cla8_u_cla14_and18 = s_wallace_cla8_u_cla14_and16 & s_wallace_cla8_u_cla14_and17;
  assign s_wallace_cla8_u_cla14_and19 = s_wallace_cla8_u_cla14_pg_logic4_and0 & s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign s_wallace_cla8_u_cla14_and20 = s_wallace_cla8_u_cla14_and19 & s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign s_wallace_cla8_u_cla14_and21 = s_wallace_cla8_u_cla14_pg_logic5_and0 & s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign s_wallace_cla8_u_cla14_or9 = s_wallace_cla8_u_cla14_and18 | s_wallace_cla8_u_cla14_and20;
  assign s_wallace_cla8_u_cla14_or10 = s_wallace_cla8_u_cla14_or9 | s_wallace_cla8_u_cla14_and21;
  assign s_wallace_cla8_u_cla14_or11 = s_wallace_cla8_u_cla14_pg_logic6_and0 | s_wallace_cla8_u_cla14_or10;
  assign s_wallace_cla8_u_cla14_pg_logic7_or0 = s_wallace_cla8_fa29_xor1 | s_wallace_cla8_fa30_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic7_and0 = s_wallace_cla8_fa29_xor1 & s_wallace_cla8_fa30_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic7_xor0 = s_wallace_cla8_fa29_xor1 ^ s_wallace_cla8_fa30_xor1;
  assign s_wallace_cla8_u_cla14_xor7 = s_wallace_cla8_u_cla14_pg_logic7_xor0 ^ s_wallace_cla8_u_cla14_or11;
  assign s_wallace_cla8_u_cla14_and22 = s_wallace_cla8_u_cla14_or5 & s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign s_wallace_cla8_u_cla14_and23 = s_wallace_cla8_u_cla14_pg_logic7_or0 & s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign s_wallace_cla8_u_cla14_and24 = s_wallace_cla8_u_cla14_and22 & s_wallace_cla8_u_cla14_and23;
  assign s_wallace_cla8_u_cla14_and25 = s_wallace_cla8_u_cla14_and24 & s_wallace_cla8_u_cla14_pg_logic4_or0;
  assign s_wallace_cla8_u_cla14_and26 = s_wallace_cla8_u_cla14_pg_logic4_and0 & s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign s_wallace_cla8_u_cla14_and27 = s_wallace_cla8_u_cla14_pg_logic7_or0 & s_wallace_cla8_u_cla14_pg_logic5_or0;
  assign s_wallace_cla8_u_cla14_and28 = s_wallace_cla8_u_cla14_and26 & s_wallace_cla8_u_cla14_and27;
  assign s_wallace_cla8_u_cla14_and29 = s_wallace_cla8_u_cla14_pg_logic5_and0 & s_wallace_cla8_u_cla14_pg_logic7_or0;
  assign s_wallace_cla8_u_cla14_and30 = s_wallace_cla8_u_cla14_and29 & s_wallace_cla8_u_cla14_pg_logic6_or0;
  assign s_wallace_cla8_u_cla14_and31 = s_wallace_cla8_u_cla14_pg_logic6_and0 & s_wallace_cla8_u_cla14_pg_logic7_or0;
  assign s_wallace_cla8_u_cla14_or12 = s_wallace_cla8_u_cla14_and25 | s_wallace_cla8_u_cla14_and30;
  assign s_wallace_cla8_u_cla14_or13 = s_wallace_cla8_u_cla14_and28 | s_wallace_cla8_u_cla14_and31;
  assign s_wallace_cla8_u_cla14_or14 = s_wallace_cla8_u_cla14_or12 | s_wallace_cla8_u_cla14_or13;
  assign s_wallace_cla8_u_cla14_or15 = s_wallace_cla8_u_cla14_pg_logic7_and0 | s_wallace_cla8_u_cla14_or14;
  assign s_wallace_cla8_u_cla14_pg_logic8_or0 = s_wallace_cla8_fa27_xor1 | s_wallace_cla8_fa31_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic8_and0 = s_wallace_cla8_fa27_xor1 & s_wallace_cla8_fa31_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic8_xor0 = s_wallace_cla8_fa27_xor1 ^ s_wallace_cla8_fa31_xor1;
  assign s_wallace_cla8_u_cla14_xor8 = s_wallace_cla8_u_cla14_pg_logic8_xor0 ^ s_wallace_cla8_u_cla14_or15;
  assign s_wallace_cla8_u_cla14_and32 = s_wallace_cla8_u_cla14_or15 & s_wallace_cla8_u_cla14_pg_logic8_or0;
  assign s_wallace_cla8_u_cla14_or16 = s_wallace_cla8_u_cla14_pg_logic8_and0 | s_wallace_cla8_u_cla14_and32;
  assign s_wallace_cla8_u_cla14_pg_logic9_or0 = s_wallace_cla8_fa23_xor1 | s_wallace_cla8_fa32_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic9_and0 = s_wallace_cla8_fa23_xor1 & s_wallace_cla8_fa32_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic9_xor0 = s_wallace_cla8_fa23_xor1 ^ s_wallace_cla8_fa32_xor1;
  assign s_wallace_cla8_u_cla14_xor9 = s_wallace_cla8_u_cla14_pg_logic9_xor0 ^ s_wallace_cla8_u_cla14_or16;
  assign s_wallace_cla8_u_cla14_and33 = s_wallace_cla8_u_cla14_or15 & s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign s_wallace_cla8_u_cla14_and34 = s_wallace_cla8_u_cla14_and33 & s_wallace_cla8_u_cla14_pg_logic8_or0;
  assign s_wallace_cla8_u_cla14_and35 = s_wallace_cla8_u_cla14_pg_logic8_and0 & s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign s_wallace_cla8_u_cla14_or17 = s_wallace_cla8_u_cla14_and34 | s_wallace_cla8_u_cla14_and35;
  assign s_wallace_cla8_u_cla14_or18 = s_wallace_cla8_u_cla14_pg_logic9_and0 | s_wallace_cla8_u_cla14_or17;
  assign s_wallace_cla8_u_cla14_pg_logic10_or0 = s_wallace_cla8_fa17_xor1 | s_wallace_cla8_fa33_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic10_and0 = s_wallace_cla8_fa17_xor1 & s_wallace_cla8_fa33_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic10_xor0 = s_wallace_cla8_fa17_xor1 ^ s_wallace_cla8_fa33_xor1;
  assign s_wallace_cla8_u_cla14_xor10 = s_wallace_cla8_u_cla14_pg_logic10_xor0 ^ s_wallace_cla8_u_cla14_or18;
  assign s_wallace_cla8_u_cla14_and36 = s_wallace_cla8_u_cla14_or15 & s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign s_wallace_cla8_u_cla14_and37 = s_wallace_cla8_u_cla14_pg_logic10_or0 & s_wallace_cla8_u_cla14_pg_logic8_or0;
  assign s_wallace_cla8_u_cla14_and38 = s_wallace_cla8_u_cla14_and36 & s_wallace_cla8_u_cla14_and37;
  assign s_wallace_cla8_u_cla14_and39 = s_wallace_cla8_u_cla14_pg_logic8_and0 & s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign s_wallace_cla8_u_cla14_and40 = s_wallace_cla8_u_cla14_and39 & s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign s_wallace_cla8_u_cla14_and41 = s_wallace_cla8_u_cla14_pg_logic9_and0 & s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign s_wallace_cla8_u_cla14_or19 = s_wallace_cla8_u_cla14_and38 | s_wallace_cla8_u_cla14_and40;
  assign s_wallace_cla8_u_cla14_or20 = s_wallace_cla8_u_cla14_or19 | s_wallace_cla8_u_cla14_and41;
  assign s_wallace_cla8_u_cla14_or21 = s_wallace_cla8_u_cla14_pg_logic10_and0 | s_wallace_cla8_u_cla14_or20;
  assign s_wallace_cla8_u_cla14_pg_logic11_or0 = s_wallace_cla8_fa9_xor1 | s_wallace_cla8_fa34_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic11_and0 = s_wallace_cla8_fa9_xor1 & s_wallace_cla8_fa34_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic11_xor0 = s_wallace_cla8_fa9_xor1 ^ s_wallace_cla8_fa34_xor1;
  assign s_wallace_cla8_u_cla14_xor11 = s_wallace_cla8_u_cla14_pg_logic11_xor0 ^ s_wallace_cla8_u_cla14_or21;
  assign s_wallace_cla8_u_cla14_and42 = s_wallace_cla8_u_cla14_or15 & s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign s_wallace_cla8_u_cla14_and43 = s_wallace_cla8_u_cla14_pg_logic11_or0 & s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign s_wallace_cla8_u_cla14_and44 = s_wallace_cla8_u_cla14_and42 & s_wallace_cla8_u_cla14_and43;
  assign s_wallace_cla8_u_cla14_and45 = s_wallace_cla8_u_cla14_and44 & s_wallace_cla8_u_cla14_pg_logic8_or0;
  assign s_wallace_cla8_u_cla14_and46 = s_wallace_cla8_u_cla14_pg_logic8_and0 & s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign s_wallace_cla8_u_cla14_and47 = s_wallace_cla8_u_cla14_pg_logic11_or0 & s_wallace_cla8_u_cla14_pg_logic9_or0;
  assign s_wallace_cla8_u_cla14_and48 = s_wallace_cla8_u_cla14_and46 & s_wallace_cla8_u_cla14_and47;
  assign s_wallace_cla8_u_cla14_and49 = s_wallace_cla8_u_cla14_pg_logic9_and0 & s_wallace_cla8_u_cla14_pg_logic11_or0;
  assign s_wallace_cla8_u_cla14_and50 = s_wallace_cla8_u_cla14_and49 & s_wallace_cla8_u_cla14_pg_logic10_or0;
  assign s_wallace_cla8_u_cla14_and51 = s_wallace_cla8_u_cla14_pg_logic10_and0 & s_wallace_cla8_u_cla14_pg_logic11_or0;
  assign s_wallace_cla8_u_cla14_or22 = s_wallace_cla8_u_cla14_and45 | s_wallace_cla8_u_cla14_and50;
  assign s_wallace_cla8_u_cla14_or23 = s_wallace_cla8_u_cla14_and48 | s_wallace_cla8_u_cla14_and51;
  assign s_wallace_cla8_u_cla14_or24 = s_wallace_cla8_u_cla14_or22 | s_wallace_cla8_u_cla14_or23;
  assign s_wallace_cla8_u_cla14_or25 = s_wallace_cla8_u_cla14_pg_logic11_and0 | s_wallace_cla8_u_cla14_or24;
  assign s_wallace_cla8_u_cla14_pg_logic12_or0 = s_wallace_cla8_nand_6_7 | s_wallace_cla8_fa35_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic12_and0 = s_wallace_cla8_nand_6_7 & s_wallace_cla8_fa35_xor1;
  assign s_wallace_cla8_u_cla14_pg_logic12_xor0 = s_wallace_cla8_nand_6_7 ^ s_wallace_cla8_fa35_xor1;
  assign s_wallace_cla8_u_cla14_xor12 = s_wallace_cla8_u_cla14_pg_logic12_xor0 ^ s_wallace_cla8_u_cla14_or25;
  assign s_wallace_cla8_u_cla14_and52 = s_wallace_cla8_u_cla14_or25 & s_wallace_cla8_u_cla14_pg_logic12_or0;
  assign s_wallace_cla8_u_cla14_or26 = s_wallace_cla8_u_cla14_pg_logic12_and0 | s_wallace_cla8_u_cla14_and52;
  assign s_wallace_cla8_u_cla14_pg_logic13_or0 = s_wallace_cla8_fa35_or0 | s_wallace_cla8_and_7_7;
  assign s_wallace_cla8_u_cla14_pg_logic13_and0 = s_wallace_cla8_fa35_or0 & s_wallace_cla8_and_7_7;
  assign s_wallace_cla8_u_cla14_pg_logic13_xor0 = s_wallace_cla8_fa35_or0 ^ s_wallace_cla8_and_7_7;
  assign s_wallace_cla8_u_cla14_xor13 = s_wallace_cla8_u_cla14_pg_logic13_xor0 ^ s_wallace_cla8_u_cla14_or26;
  assign s_wallace_cla8_u_cla14_and53 = s_wallace_cla8_u_cla14_or25 & s_wallace_cla8_u_cla14_pg_logic13_or0;
  assign s_wallace_cla8_u_cla14_and54 = s_wallace_cla8_u_cla14_and53 & s_wallace_cla8_u_cla14_pg_logic12_or0;
  assign s_wallace_cla8_u_cla14_and55 = s_wallace_cla8_u_cla14_pg_logic12_and0 & s_wallace_cla8_u_cla14_pg_logic13_or0;
  assign s_wallace_cla8_u_cla14_or27 = s_wallace_cla8_u_cla14_and54 | s_wallace_cla8_u_cla14_and55;
  assign s_wallace_cla8_u_cla14_or28 = s_wallace_cla8_u_cla14_pg_logic13_and0 | s_wallace_cla8_u_cla14_or27;
  assign s_wallace_cla8_xor0 = ~s_wallace_cla8_u_cla14_or28;

  assign s_wallace_cla8_out[0] = s_wallace_cla8_and_0_0;
  assign s_wallace_cla8_out[1] = s_wallace_cla8_u_cla14_pg_logic0_xor0;
  assign s_wallace_cla8_out[2] = s_wallace_cla8_u_cla14_xor1;
  assign s_wallace_cla8_out[3] = s_wallace_cla8_u_cla14_xor2;
  assign s_wallace_cla8_out[4] = s_wallace_cla8_u_cla14_xor3;
  assign s_wallace_cla8_out[5] = s_wallace_cla8_u_cla14_xor4;
  assign s_wallace_cla8_out[6] = s_wallace_cla8_u_cla14_xor5;
  assign s_wallace_cla8_out[7] = s_wallace_cla8_u_cla14_xor6;
  assign s_wallace_cla8_out[8] = s_wallace_cla8_u_cla14_xor7;
  assign s_wallace_cla8_out[9] = s_wallace_cla8_u_cla14_xor8;
  assign s_wallace_cla8_out[10] = s_wallace_cla8_u_cla14_xor9;
  assign s_wallace_cla8_out[11] = s_wallace_cla8_u_cla14_xor10;
  assign s_wallace_cla8_out[12] = s_wallace_cla8_u_cla14_xor11;
  assign s_wallace_cla8_out[13] = s_wallace_cla8_u_cla14_xor12;
  assign s_wallace_cla8_out[14] = s_wallace_cla8_u_cla14_xor13;
  assign s_wallace_cla8_out[15] = s_wallace_cla8_xor0;
endmodule