module s_csamul_rca16(input [15:0] a, input [15:0] b, output [31:0] s_csamul_rca16_out);
  wire s_csamul_rca16_and0_0;
  wire s_csamul_rca16_and1_0;
  wire s_csamul_rca16_and2_0;
  wire s_csamul_rca16_and3_0;
  wire s_csamul_rca16_and4_0;
  wire s_csamul_rca16_and5_0;
  wire s_csamul_rca16_and6_0;
  wire s_csamul_rca16_and7_0;
  wire s_csamul_rca16_and8_0;
  wire s_csamul_rca16_and9_0;
  wire s_csamul_rca16_and10_0;
  wire s_csamul_rca16_and11_0;
  wire s_csamul_rca16_and12_0;
  wire s_csamul_rca16_and13_0;
  wire s_csamul_rca16_and14_0;
  wire s_csamul_rca16_nand15_0;
  wire s_csamul_rca16_and0_1;
  wire s_csamul_rca16_ha0_1_xor0;
  wire s_csamul_rca16_ha0_1_and0;
  wire s_csamul_rca16_and1_1;
  wire s_csamul_rca16_ha1_1_xor0;
  wire s_csamul_rca16_ha1_1_and0;
  wire s_csamul_rca16_and2_1;
  wire s_csamul_rca16_ha2_1_xor0;
  wire s_csamul_rca16_ha2_1_and0;
  wire s_csamul_rca16_and3_1;
  wire s_csamul_rca16_ha3_1_xor0;
  wire s_csamul_rca16_ha3_1_and0;
  wire s_csamul_rca16_and4_1;
  wire s_csamul_rca16_ha4_1_xor0;
  wire s_csamul_rca16_ha4_1_and0;
  wire s_csamul_rca16_and5_1;
  wire s_csamul_rca16_ha5_1_xor0;
  wire s_csamul_rca16_ha5_1_and0;
  wire s_csamul_rca16_and6_1;
  wire s_csamul_rca16_ha6_1_xor0;
  wire s_csamul_rca16_ha6_1_and0;
  wire s_csamul_rca16_and7_1;
  wire s_csamul_rca16_ha7_1_xor0;
  wire s_csamul_rca16_ha7_1_and0;
  wire s_csamul_rca16_and8_1;
  wire s_csamul_rca16_ha8_1_xor0;
  wire s_csamul_rca16_ha8_1_and0;
  wire s_csamul_rca16_and9_1;
  wire s_csamul_rca16_ha9_1_xor0;
  wire s_csamul_rca16_ha9_1_and0;
  wire s_csamul_rca16_and10_1;
  wire s_csamul_rca16_ha10_1_xor0;
  wire s_csamul_rca16_ha10_1_and0;
  wire s_csamul_rca16_and11_1;
  wire s_csamul_rca16_ha11_1_xor0;
  wire s_csamul_rca16_ha11_1_and0;
  wire s_csamul_rca16_and12_1;
  wire s_csamul_rca16_ha12_1_xor0;
  wire s_csamul_rca16_ha12_1_and0;
  wire s_csamul_rca16_and13_1;
  wire s_csamul_rca16_ha13_1_xor0;
  wire s_csamul_rca16_ha13_1_and0;
  wire s_csamul_rca16_and14_1;
  wire s_csamul_rca16_ha14_1_xor0;
  wire s_csamul_rca16_ha14_1_and0;
  wire s_csamul_rca16_nand15_1;
  wire s_csamul_rca16_ha15_1_xor0;
  wire s_csamul_rca16_and0_2;
  wire s_csamul_rca16_fa0_2_xor0;
  wire s_csamul_rca16_fa0_2_and0;
  wire s_csamul_rca16_fa0_2_xor1;
  wire s_csamul_rca16_fa0_2_and1;
  wire s_csamul_rca16_fa0_2_or0;
  wire s_csamul_rca16_and1_2;
  wire s_csamul_rca16_fa1_2_xor0;
  wire s_csamul_rca16_fa1_2_and0;
  wire s_csamul_rca16_fa1_2_xor1;
  wire s_csamul_rca16_fa1_2_and1;
  wire s_csamul_rca16_fa1_2_or0;
  wire s_csamul_rca16_and2_2;
  wire s_csamul_rca16_fa2_2_xor0;
  wire s_csamul_rca16_fa2_2_and0;
  wire s_csamul_rca16_fa2_2_xor1;
  wire s_csamul_rca16_fa2_2_and1;
  wire s_csamul_rca16_fa2_2_or0;
  wire s_csamul_rca16_and3_2;
  wire s_csamul_rca16_fa3_2_xor0;
  wire s_csamul_rca16_fa3_2_and0;
  wire s_csamul_rca16_fa3_2_xor1;
  wire s_csamul_rca16_fa3_2_and1;
  wire s_csamul_rca16_fa3_2_or0;
  wire s_csamul_rca16_and4_2;
  wire s_csamul_rca16_fa4_2_xor0;
  wire s_csamul_rca16_fa4_2_and0;
  wire s_csamul_rca16_fa4_2_xor1;
  wire s_csamul_rca16_fa4_2_and1;
  wire s_csamul_rca16_fa4_2_or0;
  wire s_csamul_rca16_and5_2;
  wire s_csamul_rca16_fa5_2_xor0;
  wire s_csamul_rca16_fa5_2_and0;
  wire s_csamul_rca16_fa5_2_xor1;
  wire s_csamul_rca16_fa5_2_and1;
  wire s_csamul_rca16_fa5_2_or0;
  wire s_csamul_rca16_and6_2;
  wire s_csamul_rca16_fa6_2_xor0;
  wire s_csamul_rca16_fa6_2_and0;
  wire s_csamul_rca16_fa6_2_xor1;
  wire s_csamul_rca16_fa6_2_and1;
  wire s_csamul_rca16_fa6_2_or0;
  wire s_csamul_rca16_and7_2;
  wire s_csamul_rca16_fa7_2_xor0;
  wire s_csamul_rca16_fa7_2_and0;
  wire s_csamul_rca16_fa7_2_xor1;
  wire s_csamul_rca16_fa7_2_and1;
  wire s_csamul_rca16_fa7_2_or0;
  wire s_csamul_rca16_and8_2;
  wire s_csamul_rca16_fa8_2_xor0;
  wire s_csamul_rca16_fa8_2_and0;
  wire s_csamul_rca16_fa8_2_xor1;
  wire s_csamul_rca16_fa8_2_and1;
  wire s_csamul_rca16_fa8_2_or0;
  wire s_csamul_rca16_and9_2;
  wire s_csamul_rca16_fa9_2_xor0;
  wire s_csamul_rca16_fa9_2_and0;
  wire s_csamul_rca16_fa9_2_xor1;
  wire s_csamul_rca16_fa9_2_and1;
  wire s_csamul_rca16_fa9_2_or0;
  wire s_csamul_rca16_and10_2;
  wire s_csamul_rca16_fa10_2_xor0;
  wire s_csamul_rca16_fa10_2_and0;
  wire s_csamul_rca16_fa10_2_xor1;
  wire s_csamul_rca16_fa10_2_and1;
  wire s_csamul_rca16_fa10_2_or0;
  wire s_csamul_rca16_and11_2;
  wire s_csamul_rca16_fa11_2_xor0;
  wire s_csamul_rca16_fa11_2_and0;
  wire s_csamul_rca16_fa11_2_xor1;
  wire s_csamul_rca16_fa11_2_and1;
  wire s_csamul_rca16_fa11_2_or0;
  wire s_csamul_rca16_and12_2;
  wire s_csamul_rca16_fa12_2_xor0;
  wire s_csamul_rca16_fa12_2_and0;
  wire s_csamul_rca16_fa12_2_xor1;
  wire s_csamul_rca16_fa12_2_and1;
  wire s_csamul_rca16_fa12_2_or0;
  wire s_csamul_rca16_and13_2;
  wire s_csamul_rca16_fa13_2_xor0;
  wire s_csamul_rca16_fa13_2_and0;
  wire s_csamul_rca16_fa13_2_xor1;
  wire s_csamul_rca16_fa13_2_and1;
  wire s_csamul_rca16_fa13_2_or0;
  wire s_csamul_rca16_and14_2;
  wire s_csamul_rca16_fa14_2_xor0;
  wire s_csamul_rca16_fa14_2_and0;
  wire s_csamul_rca16_fa14_2_xor1;
  wire s_csamul_rca16_fa14_2_and1;
  wire s_csamul_rca16_fa14_2_or0;
  wire s_csamul_rca16_nand15_2;
  wire s_csamul_rca16_ha15_2_xor0;
  wire s_csamul_rca16_ha15_2_and0;
  wire s_csamul_rca16_and0_3;
  wire s_csamul_rca16_fa0_3_xor0;
  wire s_csamul_rca16_fa0_3_and0;
  wire s_csamul_rca16_fa0_3_xor1;
  wire s_csamul_rca16_fa0_3_and1;
  wire s_csamul_rca16_fa0_3_or0;
  wire s_csamul_rca16_and1_3;
  wire s_csamul_rca16_fa1_3_xor0;
  wire s_csamul_rca16_fa1_3_and0;
  wire s_csamul_rca16_fa1_3_xor1;
  wire s_csamul_rca16_fa1_3_and1;
  wire s_csamul_rca16_fa1_3_or0;
  wire s_csamul_rca16_and2_3;
  wire s_csamul_rca16_fa2_3_xor0;
  wire s_csamul_rca16_fa2_3_and0;
  wire s_csamul_rca16_fa2_3_xor1;
  wire s_csamul_rca16_fa2_3_and1;
  wire s_csamul_rca16_fa2_3_or0;
  wire s_csamul_rca16_and3_3;
  wire s_csamul_rca16_fa3_3_xor0;
  wire s_csamul_rca16_fa3_3_and0;
  wire s_csamul_rca16_fa3_3_xor1;
  wire s_csamul_rca16_fa3_3_and1;
  wire s_csamul_rca16_fa3_3_or0;
  wire s_csamul_rca16_and4_3;
  wire s_csamul_rca16_fa4_3_xor0;
  wire s_csamul_rca16_fa4_3_and0;
  wire s_csamul_rca16_fa4_3_xor1;
  wire s_csamul_rca16_fa4_3_and1;
  wire s_csamul_rca16_fa4_3_or0;
  wire s_csamul_rca16_and5_3;
  wire s_csamul_rca16_fa5_3_xor0;
  wire s_csamul_rca16_fa5_3_and0;
  wire s_csamul_rca16_fa5_3_xor1;
  wire s_csamul_rca16_fa5_3_and1;
  wire s_csamul_rca16_fa5_3_or0;
  wire s_csamul_rca16_and6_3;
  wire s_csamul_rca16_fa6_3_xor0;
  wire s_csamul_rca16_fa6_3_and0;
  wire s_csamul_rca16_fa6_3_xor1;
  wire s_csamul_rca16_fa6_3_and1;
  wire s_csamul_rca16_fa6_3_or0;
  wire s_csamul_rca16_and7_3;
  wire s_csamul_rca16_fa7_3_xor0;
  wire s_csamul_rca16_fa7_3_and0;
  wire s_csamul_rca16_fa7_3_xor1;
  wire s_csamul_rca16_fa7_3_and1;
  wire s_csamul_rca16_fa7_3_or0;
  wire s_csamul_rca16_and8_3;
  wire s_csamul_rca16_fa8_3_xor0;
  wire s_csamul_rca16_fa8_3_and0;
  wire s_csamul_rca16_fa8_3_xor1;
  wire s_csamul_rca16_fa8_3_and1;
  wire s_csamul_rca16_fa8_3_or0;
  wire s_csamul_rca16_and9_3;
  wire s_csamul_rca16_fa9_3_xor0;
  wire s_csamul_rca16_fa9_3_and0;
  wire s_csamul_rca16_fa9_3_xor1;
  wire s_csamul_rca16_fa9_3_and1;
  wire s_csamul_rca16_fa9_3_or0;
  wire s_csamul_rca16_and10_3;
  wire s_csamul_rca16_fa10_3_xor0;
  wire s_csamul_rca16_fa10_3_and0;
  wire s_csamul_rca16_fa10_3_xor1;
  wire s_csamul_rca16_fa10_3_and1;
  wire s_csamul_rca16_fa10_3_or0;
  wire s_csamul_rca16_and11_3;
  wire s_csamul_rca16_fa11_3_xor0;
  wire s_csamul_rca16_fa11_3_and0;
  wire s_csamul_rca16_fa11_3_xor1;
  wire s_csamul_rca16_fa11_3_and1;
  wire s_csamul_rca16_fa11_3_or0;
  wire s_csamul_rca16_and12_3;
  wire s_csamul_rca16_fa12_3_xor0;
  wire s_csamul_rca16_fa12_3_and0;
  wire s_csamul_rca16_fa12_3_xor1;
  wire s_csamul_rca16_fa12_3_and1;
  wire s_csamul_rca16_fa12_3_or0;
  wire s_csamul_rca16_and13_3;
  wire s_csamul_rca16_fa13_3_xor0;
  wire s_csamul_rca16_fa13_3_and0;
  wire s_csamul_rca16_fa13_3_xor1;
  wire s_csamul_rca16_fa13_3_and1;
  wire s_csamul_rca16_fa13_3_or0;
  wire s_csamul_rca16_and14_3;
  wire s_csamul_rca16_fa14_3_xor0;
  wire s_csamul_rca16_fa14_3_and0;
  wire s_csamul_rca16_fa14_3_xor1;
  wire s_csamul_rca16_fa14_3_and1;
  wire s_csamul_rca16_fa14_3_or0;
  wire s_csamul_rca16_nand15_3;
  wire s_csamul_rca16_ha15_3_xor0;
  wire s_csamul_rca16_ha15_3_and0;
  wire s_csamul_rca16_and0_4;
  wire s_csamul_rca16_fa0_4_xor0;
  wire s_csamul_rca16_fa0_4_and0;
  wire s_csamul_rca16_fa0_4_xor1;
  wire s_csamul_rca16_fa0_4_and1;
  wire s_csamul_rca16_fa0_4_or0;
  wire s_csamul_rca16_and1_4;
  wire s_csamul_rca16_fa1_4_xor0;
  wire s_csamul_rca16_fa1_4_and0;
  wire s_csamul_rca16_fa1_4_xor1;
  wire s_csamul_rca16_fa1_4_and1;
  wire s_csamul_rca16_fa1_4_or0;
  wire s_csamul_rca16_and2_4;
  wire s_csamul_rca16_fa2_4_xor0;
  wire s_csamul_rca16_fa2_4_and0;
  wire s_csamul_rca16_fa2_4_xor1;
  wire s_csamul_rca16_fa2_4_and1;
  wire s_csamul_rca16_fa2_4_or0;
  wire s_csamul_rca16_and3_4;
  wire s_csamul_rca16_fa3_4_xor0;
  wire s_csamul_rca16_fa3_4_and0;
  wire s_csamul_rca16_fa3_4_xor1;
  wire s_csamul_rca16_fa3_4_and1;
  wire s_csamul_rca16_fa3_4_or0;
  wire s_csamul_rca16_and4_4;
  wire s_csamul_rca16_fa4_4_xor0;
  wire s_csamul_rca16_fa4_4_and0;
  wire s_csamul_rca16_fa4_4_xor1;
  wire s_csamul_rca16_fa4_4_and1;
  wire s_csamul_rca16_fa4_4_or0;
  wire s_csamul_rca16_and5_4;
  wire s_csamul_rca16_fa5_4_xor0;
  wire s_csamul_rca16_fa5_4_and0;
  wire s_csamul_rca16_fa5_4_xor1;
  wire s_csamul_rca16_fa5_4_and1;
  wire s_csamul_rca16_fa5_4_or0;
  wire s_csamul_rca16_and6_4;
  wire s_csamul_rca16_fa6_4_xor0;
  wire s_csamul_rca16_fa6_4_and0;
  wire s_csamul_rca16_fa6_4_xor1;
  wire s_csamul_rca16_fa6_4_and1;
  wire s_csamul_rca16_fa6_4_or0;
  wire s_csamul_rca16_and7_4;
  wire s_csamul_rca16_fa7_4_xor0;
  wire s_csamul_rca16_fa7_4_and0;
  wire s_csamul_rca16_fa7_4_xor1;
  wire s_csamul_rca16_fa7_4_and1;
  wire s_csamul_rca16_fa7_4_or0;
  wire s_csamul_rca16_and8_4;
  wire s_csamul_rca16_fa8_4_xor0;
  wire s_csamul_rca16_fa8_4_and0;
  wire s_csamul_rca16_fa8_4_xor1;
  wire s_csamul_rca16_fa8_4_and1;
  wire s_csamul_rca16_fa8_4_or0;
  wire s_csamul_rca16_and9_4;
  wire s_csamul_rca16_fa9_4_xor0;
  wire s_csamul_rca16_fa9_4_and0;
  wire s_csamul_rca16_fa9_4_xor1;
  wire s_csamul_rca16_fa9_4_and1;
  wire s_csamul_rca16_fa9_4_or0;
  wire s_csamul_rca16_and10_4;
  wire s_csamul_rca16_fa10_4_xor0;
  wire s_csamul_rca16_fa10_4_and0;
  wire s_csamul_rca16_fa10_4_xor1;
  wire s_csamul_rca16_fa10_4_and1;
  wire s_csamul_rca16_fa10_4_or0;
  wire s_csamul_rca16_and11_4;
  wire s_csamul_rca16_fa11_4_xor0;
  wire s_csamul_rca16_fa11_4_and0;
  wire s_csamul_rca16_fa11_4_xor1;
  wire s_csamul_rca16_fa11_4_and1;
  wire s_csamul_rca16_fa11_4_or0;
  wire s_csamul_rca16_and12_4;
  wire s_csamul_rca16_fa12_4_xor0;
  wire s_csamul_rca16_fa12_4_and0;
  wire s_csamul_rca16_fa12_4_xor1;
  wire s_csamul_rca16_fa12_4_and1;
  wire s_csamul_rca16_fa12_4_or0;
  wire s_csamul_rca16_and13_4;
  wire s_csamul_rca16_fa13_4_xor0;
  wire s_csamul_rca16_fa13_4_and0;
  wire s_csamul_rca16_fa13_4_xor1;
  wire s_csamul_rca16_fa13_4_and1;
  wire s_csamul_rca16_fa13_4_or0;
  wire s_csamul_rca16_and14_4;
  wire s_csamul_rca16_fa14_4_xor0;
  wire s_csamul_rca16_fa14_4_and0;
  wire s_csamul_rca16_fa14_4_xor1;
  wire s_csamul_rca16_fa14_4_and1;
  wire s_csamul_rca16_fa14_4_or0;
  wire s_csamul_rca16_nand15_4;
  wire s_csamul_rca16_ha15_4_xor0;
  wire s_csamul_rca16_ha15_4_and0;
  wire s_csamul_rca16_and0_5;
  wire s_csamul_rca16_fa0_5_xor0;
  wire s_csamul_rca16_fa0_5_and0;
  wire s_csamul_rca16_fa0_5_xor1;
  wire s_csamul_rca16_fa0_5_and1;
  wire s_csamul_rca16_fa0_5_or0;
  wire s_csamul_rca16_and1_5;
  wire s_csamul_rca16_fa1_5_xor0;
  wire s_csamul_rca16_fa1_5_and0;
  wire s_csamul_rca16_fa1_5_xor1;
  wire s_csamul_rca16_fa1_5_and1;
  wire s_csamul_rca16_fa1_5_or0;
  wire s_csamul_rca16_and2_5;
  wire s_csamul_rca16_fa2_5_xor0;
  wire s_csamul_rca16_fa2_5_and0;
  wire s_csamul_rca16_fa2_5_xor1;
  wire s_csamul_rca16_fa2_5_and1;
  wire s_csamul_rca16_fa2_5_or0;
  wire s_csamul_rca16_and3_5;
  wire s_csamul_rca16_fa3_5_xor0;
  wire s_csamul_rca16_fa3_5_and0;
  wire s_csamul_rca16_fa3_5_xor1;
  wire s_csamul_rca16_fa3_5_and1;
  wire s_csamul_rca16_fa3_5_or0;
  wire s_csamul_rca16_and4_5;
  wire s_csamul_rca16_fa4_5_xor0;
  wire s_csamul_rca16_fa4_5_and0;
  wire s_csamul_rca16_fa4_5_xor1;
  wire s_csamul_rca16_fa4_5_and1;
  wire s_csamul_rca16_fa4_5_or0;
  wire s_csamul_rca16_and5_5;
  wire s_csamul_rca16_fa5_5_xor0;
  wire s_csamul_rca16_fa5_5_and0;
  wire s_csamul_rca16_fa5_5_xor1;
  wire s_csamul_rca16_fa5_5_and1;
  wire s_csamul_rca16_fa5_5_or0;
  wire s_csamul_rca16_and6_5;
  wire s_csamul_rca16_fa6_5_xor0;
  wire s_csamul_rca16_fa6_5_and0;
  wire s_csamul_rca16_fa6_5_xor1;
  wire s_csamul_rca16_fa6_5_and1;
  wire s_csamul_rca16_fa6_5_or0;
  wire s_csamul_rca16_and7_5;
  wire s_csamul_rca16_fa7_5_xor0;
  wire s_csamul_rca16_fa7_5_and0;
  wire s_csamul_rca16_fa7_5_xor1;
  wire s_csamul_rca16_fa7_5_and1;
  wire s_csamul_rca16_fa7_5_or0;
  wire s_csamul_rca16_and8_5;
  wire s_csamul_rca16_fa8_5_xor0;
  wire s_csamul_rca16_fa8_5_and0;
  wire s_csamul_rca16_fa8_5_xor1;
  wire s_csamul_rca16_fa8_5_and1;
  wire s_csamul_rca16_fa8_5_or0;
  wire s_csamul_rca16_and9_5;
  wire s_csamul_rca16_fa9_5_xor0;
  wire s_csamul_rca16_fa9_5_and0;
  wire s_csamul_rca16_fa9_5_xor1;
  wire s_csamul_rca16_fa9_5_and1;
  wire s_csamul_rca16_fa9_5_or0;
  wire s_csamul_rca16_and10_5;
  wire s_csamul_rca16_fa10_5_xor0;
  wire s_csamul_rca16_fa10_5_and0;
  wire s_csamul_rca16_fa10_5_xor1;
  wire s_csamul_rca16_fa10_5_and1;
  wire s_csamul_rca16_fa10_5_or0;
  wire s_csamul_rca16_and11_5;
  wire s_csamul_rca16_fa11_5_xor0;
  wire s_csamul_rca16_fa11_5_and0;
  wire s_csamul_rca16_fa11_5_xor1;
  wire s_csamul_rca16_fa11_5_and1;
  wire s_csamul_rca16_fa11_5_or0;
  wire s_csamul_rca16_and12_5;
  wire s_csamul_rca16_fa12_5_xor0;
  wire s_csamul_rca16_fa12_5_and0;
  wire s_csamul_rca16_fa12_5_xor1;
  wire s_csamul_rca16_fa12_5_and1;
  wire s_csamul_rca16_fa12_5_or0;
  wire s_csamul_rca16_and13_5;
  wire s_csamul_rca16_fa13_5_xor0;
  wire s_csamul_rca16_fa13_5_and0;
  wire s_csamul_rca16_fa13_5_xor1;
  wire s_csamul_rca16_fa13_5_and1;
  wire s_csamul_rca16_fa13_5_or0;
  wire s_csamul_rca16_and14_5;
  wire s_csamul_rca16_fa14_5_xor0;
  wire s_csamul_rca16_fa14_5_and0;
  wire s_csamul_rca16_fa14_5_xor1;
  wire s_csamul_rca16_fa14_5_and1;
  wire s_csamul_rca16_fa14_5_or0;
  wire s_csamul_rca16_nand15_5;
  wire s_csamul_rca16_ha15_5_xor0;
  wire s_csamul_rca16_ha15_5_and0;
  wire s_csamul_rca16_and0_6;
  wire s_csamul_rca16_fa0_6_xor0;
  wire s_csamul_rca16_fa0_6_and0;
  wire s_csamul_rca16_fa0_6_xor1;
  wire s_csamul_rca16_fa0_6_and1;
  wire s_csamul_rca16_fa0_6_or0;
  wire s_csamul_rca16_and1_6;
  wire s_csamul_rca16_fa1_6_xor0;
  wire s_csamul_rca16_fa1_6_and0;
  wire s_csamul_rca16_fa1_6_xor1;
  wire s_csamul_rca16_fa1_6_and1;
  wire s_csamul_rca16_fa1_6_or0;
  wire s_csamul_rca16_and2_6;
  wire s_csamul_rca16_fa2_6_xor0;
  wire s_csamul_rca16_fa2_6_and0;
  wire s_csamul_rca16_fa2_6_xor1;
  wire s_csamul_rca16_fa2_6_and1;
  wire s_csamul_rca16_fa2_6_or0;
  wire s_csamul_rca16_and3_6;
  wire s_csamul_rca16_fa3_6_xor0;
  wire s_csamul_rca16_fa3_6_and0;
  wire s_csamul_rca16_fa3_6_xor1;
  wire s_csamul_rca16_fa3_6_and1;
  wire s_csamul_rca16_fa3_6_or0;
  wire s_csamul_rca16_and4_6;
  wire s_csamul_rca16_fa4_6_xor0;
  wire s_csamul_rca16_fa4_6_and0;
  wire s_csamul_rca16_fa4_6_xor1;
  wire s_csamul_rca16_fa4_6_and1;
  wire s_csamul_rca16_fa4_6_or0;
  wire s_csamul_rca16_and5_6;
  wire s_csamul_rca16_fa5_6_xor0;
  wire s_csamul_rca16_fa5_6_and0;
  wire s_csamul_rca16_fa5_6_xor1;
  wire s_csamul_rca16_fa5_6_and1;
  wire s_csamul_rca16_fa5_6_or0;
  wire s_csamul_rca16_and6_6;
  wire s_csamul_rca16_fa6_6_xor0;
  wire s_csamul_rca16_fa6_6_and0;
  wire s_csamul_rca16_fa6_6_xor1;
  wire s_csamul_rca16_fa6_6_and1;
  wire s_csamul_rca16_fa6_6_or0;
  wire s_csamul_rca16_and7_6;
  wire s_csamul_rca16_fa7_6_xor0;
  wire s_csamul_rca16_fa7_6_and0;
  wire s_csamul_rca16_fa7_6_xor1;
  wire s_csamul_rca16_fa7_6_and1;
  wire s_csamul_rca16_fa7_6_or0;
  wire s_csamul_rca16_and8_6;
  wire s_csamul_rca16_fa8_6_xor0;
  wire s_csamul_rca16_fa8_6_and0;
  wire s_csamul_rca16_fa8_6_xor1;
  wire s_csamul_rca16_fa8_6_and1;
  wire s_csamul_rca16_fa8_6_or0;
  wire s_csamul_rca16_and9_6;
  wire s_csamul_rca16_fa9_6_xor0;
  wire s_csamul_rca16_fa9_6_and0;
  wire s_csamul_rca16_fa9_6_xor1;
  wire s_csamul_rca16_fa9_6_and1;
  wire s_csamul_rca16_fa9_6_or0;
  wire s_csamul_rca16_and10_6;
  wire s_csamul_rca16_fa10_6_xor0;
  wire s_csamul_rca16_fa10_6_and0;
  wire s_csamul_rca16_fa10_6_xor1;
  wire s_csamul_rca16_fa10_6_and1;
  wire s_csamul_rca16_fa10_6_or0;
  wire s_csamul_rca16_and11_6;
  wire s_csamul_rca16_fa11_6_xor0;
  wire s_csamul_rca16_fa11_6_and0;
  wire s_csamul_rca16_fa11_6_xor1;
  wire s_csamul_rca16_fa11_6_and1;
  wire s_csamul_rca16_fa11_6_or0;
  wire s_csamul_rca16_and12_6;
  wire s_csamul_rca16_fa12_6_xor0;
  wire s_csamul_rca16_fa12_6_and0;
  wire s_csamul_rca16_fa12_6_xor1;
  wire s_csamul_rca16_fa12_6_and1;
  wire s_csamul_rca16_fa12_6_or0;
  wire s_csamul_rca16_and13_6;
  wire s_csamul_rca16_fa13_6_xor0;
  wire s_csamul_rca16_fa13_6_and0;
  wire s_csamul_rca16_fa13_6_xor1;
  wire s_csamul_rca16_fa13_6_and1;
  wire s_csamul_rca16_fa13_6_or0;
  wire s_csamul_rca16_and14_6;
  wire s_csamul_rca16_fa14_6_xor0;
  wire s_csamul_rca16_fa14_6_and0;
  wire s_csamul_rca16_fa14_6_xor1;
  wire s_csamul_rca16_fa14_6_and1;
  wire s_csamul_rca16_fa14_6_or0;
  wire s_csamul_rca16_nand15_6;
  wire s_csamul_rca16_ha15_6_xor0;
  wire s_csamul_rca16_ha15_6_and0;
  wire s_csamul_rca16_and0_7;
  wire s_csamul_rca16_fa0_7_xor0;
  wire s_csamul_rca16_fa0_7_and0;
  wire s_csamul_rca16_fa0_7_xor1;
  wire s_csamul_rca16_fa0_7_and1;
  wire s_csamul_rca16_fa0_7_or0;
  wire s_csamul_rca16_and1_7;
  wire s_csamul_rca16_fa1_7_xor0;
  wire s_csamul_rca16_fa1_7_and0;
  wire s_csamul_rca16_fa1_7_xor1;
  wire s_csamul_rca16_fa1_7_and1;
  wire s_csamul_rca16_fa1_7_or0;
  wire s_csamul_rca16_and2_7;
  wire s_csamul_rca16_fa2_7_xor0;
  wire s_csamul_rca16_fa2_7_and0;
  wire s_csamul_rca16_fa2_7_xor1;
  wire s_csamul_rca16_fa2_7_and1;
  wire s_csamul_rca16_fa2_7_or0;
  wire s_csamul_rca16_and3_7;
  wire s_csamul_rca16_fa3_7_xor0;
  wire s_csamul_rca16_fa3_7_and0;
  wire s_csamul_rca16_fa3_7_xor1;
  wire s_csamul_rca16_fa3_7_and1;
  wire s_csamul_rca16_fa3_7_or0;
  wire s_csamul_rca16_and4_7;
  wire s_csamul_rca16_fa4_7_xor0;
  wire s_csamul_rca16_fa4_7_and0;
  wire s_csamul_rca16_fa4_7_xor1;
  wire s_csamul_rca16_fa4_7_and1;
  wire s_csamul_rca16_fa4_7_or0;
  wire s_csamul_rca16_and5_7;
  wire s_csamul_rca16_fa5_7_xor0;
  wire s_csamul_rca16_fa5_7_and0;
  wire s_csamul_rca16_fa5_7_xor1;
  wire s_csamul_rca16_fa5_7_and1;
  wire s_csamul_rca16_fa5_7_or0;
  wire s_csamul_rca16_and6_7;
  wire s_csamul_rca16_fa6_7_xor0;
  wire s_csamul_rca16_fa6_7_and0;
  wire s_csamul_rca16_fa6_7_xor1;
  wire s_csamul_rca16_fa6_7_and1;
  wire s_csamul_rca16_fa6_7_or0;
  wire s_csamul_rca16_and7_7;
  wire s_csamul_rca16_fa7_7_xor0;
  wire s_csamul_rca16_fa7_7_and0;
  wire s_csamul_rca16_fa7_7_xor1;
  wire s_csamul_rca16_fa7_7_and1;
  wire s_csamul_rca16_fa7_7_or0;
  wire s_csamul_rca16_and8_7;
  wire s_csamul_rca16_fa8_7_xor0;
  wire s_csamul_rca16_fa8_7_and0;
  wire s_csamul_rca16_fa8_7_xor1;
  wire s_csamul_rca16_fa8_7_and1;
  wire s_csamul_rca16_fa8_7_or0;
  wire s_csamul_rca16_and9_7;
  wire s_csamul_rca16_fa9_7_xor0;
  wire s_csamul_rca16_fa9_7_and0;
  wire s_csamul_rca16_fa9_7_xor1;
  wire s_csamul_rca16_fa9_7_and1;
  wire s_csamul_rca16_fa9_7_or0;
  wire s_csamul_rca16_and10_7;
  wire s_csamul_rca16_fa10_7_xor0;
  wire s_csamul_rca16_fa10_7_and0;
  wire s_csamul_rca16_fa10_7_xor1;
  wire s_csamul_rca16_fa10_7_and1;
  wire s_csamul_rca16_fa10_7_or0;
  wire s_csamul_rca16_and11_7;
  wire s_csamul_rca16_fa11_7_xor0;
  wire s_csamul_rca16_fa11_7_and0;
  wire s_csamul_rca16_fa11_7_xor1;
  wire s_csamul_rca16_fa11_7_and1;
  wire s_csamul_rca16_fa11_7_or0;
  wire s_csamul_rca16_and12_7;
  wire s_csamul_rca16_fa12_7_xor0;
  wire s_csamul_rca16_fa12_7_and0;
  wire s_csamul_rca16_fa12_7_xor1;
  wire s_csamul_rca16_fa12_7_and1;
  wire s_csamul_rca16_fa12_7_or0;
  wire s_csamul_rca16_and13_7;
  wire s_csamul_rca16_fa13_7_xor0;
  wire s_csamul_rca16_fa13_7_and0;
  wire s_csamul_rca16_fa13_7_xor1;
  wire s_csamul_rca16_fa13_7_and1;
  wire s_csamul_rca16_fa13_7_or0;
  wire s_csamul_rca16_and14_7;
  wire s_csamul_rca16_fa14_7_xor0;
  wire s_csamul_rca16_fa14_7_and0;
  wire s_csamul_rca16_fa14_7_xor1;
  wire s_csamul_rca16_fa14_7_and1;
  wire s_csamul_rca16_fa14_7_or0;
  wire s_csamul_rca16_nand15_7;
  wire s_csamul_rca16_ha15_7_xor0;
  wire s_csamul_rca16_ha15_7_and0;
  wire s_csamul_rca16_and0_8;
  wire s_csamul_rca16_fa0_8_xor0;
  wire s_csamul_rca16_fa0_8_and0;
  wire s_csamul_rca16_fa0_8_xor1;
  wire s_csamul_rca16_fa0_8_and1;
  wire s_csamul_rca16_fa0_8_or0;
  wire s_csamul_rca16_and1_8;
  wire s_csamul_rca16_fa1_8_xor0;
  wire s_csamul_rca16_fa1_8_and0;
  wire s_csamul_rca16_fa1_8_xor1;
  wire s_csamul_rca16_fa1_8_and1;
  wire s_csamul_rca16_fa1_8_or0;
  wire s_csamul_rca16_and2_8;
  wire s_csamul_rca16_fa2_8_xor0;
  wire s_csamul_rca16_fa2_8_and0;
  wire s_csamul_rca16_fa2_8_xor1;
  wire s_csamul_rca16_fa2_8_and1;
  wire s_csamul_rca16_fa2_8_or0;
  wire s_csamul_rca16_and3_8;
  wire s_csamul_rca16_fa3_8_xor0;
  wire s_csamul_rca16_fa3_8_and0;
  wire s_csamul_rca16_fa3_8_xor1;
  wire s_csamul_rca16_fa3_8_and1;
  wire s_csamul_rca16_fa3_8_or0;
  wire s_csamul_rca16_and4_8;
  wire s_csamul_rca16_fa4_8_xor0;
  wire s_csamul_rca16_fa4_8_and0;
  wire s_csamul_rca16_fa4_8_xor1;
  wire s_csamul_rca16_fa4_8_and1;
  wire s_csamul_rca16_fa4_8_or0;
  wire s_csamul_rca16_and5_8;
  wire s_csamul_rca16_fa5_8_xor0;
  wire s_csamul_rca16_fa5_8_and0;
  wire s_csamul_rca16_fa5_8_xor1;
  wire s_csamul_rca16_fa5_8_and1;
  wire s_csamul_rca16_fa5_8_or0;
  wire s_csamul_rca16_and6_8;
  wire s_csamul_rca16_fa6_8_xor0;
  wire s_csamul_rca16_fa6_8_and0;
  wire s_csamul_rca16_fa6_8_xor1;
  wire s_csamul_rca16_fa6_8_and1;
  wire s_csamul_rca16_fa6_8_or0;
  wire s_csamul_rca16_and7_8;
  wire s_csamul_rca16_fa7_8_xor0;
  wire s_csamul_rca16_fa7_8_and0;
  wire s_csamul_rca16_fa7_8_xor1;
  wire s_csamul_rca16_fa7_8_and1;
  wire s_csamul_rca16_fa7_8_or0;
  wire s_csamul_rca16_and8_8;
  wire s_csamul_rca16_fa8_8_xor0;
  wire s_csamul_rca16_fa8_8_and0;
  wire s_csamul_rca16_fa8_8_xor1;
  wire s_csamul_rca16_fa8_8_and1;
  wire s_csamul_rca16_fa8_8_or0;
  wire s_csamul_rca16_and9_8;
  wire s_csamul_rca16_fa9_8_xor0;
  wire s_csamul_rca16_fa9_8_and0;
  wire s_csamul_rca16_fa9_8_xor1;
  wire s_csamul_rca16_fa9_8_and1;
  wire s_csamul_rca16_fa9_8_or0;
  wire s_csamul_rca16_and10_8;
  wire s_csamul_rca16_fa10_8_xor0;
  wire s_csamul_rca16_fa10_8_and0;
  wire s_csamul_rca16_fa10_8_xor1;
  wire s_csamul_rca16_fa10_8_and1;
  wire s_csamul_rca16_fa10_8_or0;
  wire s_csamul_rca16_and11_8;
  wire s_csamul_rca16_fa11_8_xor0;
  wire s_csamul_rca16_fa11_8_and0;
  wire s_csamul_rca16_fa11_8_xor1;
  wire s_csamul_rca16_fa11_8_and1;
  wire s_csamul_rca16_fa11_8_or0;
  wire s_csamul_rca16_and12_8;
  wire s_csamul_rca16_fa12_8_xor0;
  wire s_csamul_rca16_fa12_8_and0;
  wire s_csamul_rca16_fa12_8_xor1;
  wire s_csamul_rca16_fa12_8_and1;
  wire s_csamul_rca16_fa12_8_or0;
  wire s_csamul_rca16_and13_8;
  wire s_csamul_rca16_fa13_8_xor0;
  wire s_csamul_rca16_fa13_8_and0;
  wire s_csamul_rca16_fa13_8_xor1;
  wire s_csamul_rca16_fa13_8_and1;
  wire s_csamul_rca16_fa13_8_or0;
  wire s_csamul_rca16_and14_8;
  wire s_csamul_rca16_fa14_8_xor0;
  wire s_csamul_rca16_fa14_8_and0;
  wire s_csamul_rca16_fa14_8_xor1;
  wire s_csamul_rca16_fa14_8_and1;
  wire s_csamul_rca16_fa14_8_or0;
  wire s_csamul_rca16_nand15_8;
  wire s_csamul_rca16_ha15_8_xor0;
  wire s_csamul_rca16_ha15_8_and0;
  wire s_csamul_rca16_and0_9;
  wire s_csamul_rca16_fa0_9_xor0;
  wire s_csamul_rca16_fa0_9_and0;
  wire s_csamul_rca16_fa0_9_xor1;
  wire s_csamul_rca16_fa0_9_and1;
  wire s_csamul_rca16_fa0_9_or0;
  wire s_csamul_rca16_and1_9;
  wire s_csamul_rca16_fa1_9_xor0;
  wire s_csamul_rca16_fa1_9_and0;
  wire s_csamul_rca16_fa1_9_xor1;
  wire s_csamul_rca16_fa1_9_and1;
  wire s_csamul_rca16_fa1_9_or0;
  wire s_csamul_rca16_and2_9;
  wire s_csamul_rca16_fa2_9_xor0;
  wire s_csamul_rca16_fa2_9_and0;
  wire s_csamul_rca16_fa2_9_xor1;
  wire s_csamul_rca16_fa2_9_and1;
  wire s_csamul_rca16_fa2_9_or0;
  wire s_csamul_rca16_and3_9;
  wire s_csamul_rca16_fa3_9_xor0;
  wire s_csamul_rca16_fa3_9_and0;
  wire s_csamul_rca16_fa3_9_xor1;
  wire s_csamul_rca16_fa3_9_and1;
  wire s_csamul_rca16_fa3_9_or0;
  wire s_csamul_rca16_and4_9;
  wire s_csamul_rca16_fa4_9_xor0;
  wire s_csamul_rca16_fa4_9_and0;
  wire s_csamul_rca16_fa4_9_xor1;
  wire s_csamul_rca16_fa4_9_and1;
  wire s_csamul_rca16_fa4_9_or0;
  wire s_csamul_rca16_and5_9;
  wire s_csamul_rca16_fa5_9_xor0;
  wire s_csamul_rca16_fa5_9_and0;
  wire s_csamul_rca16_fa5_9_xor1;
  wire s_csamul_rca16_fa5_9_and1;
  wire s_csamul_rca16_fa5_9_or0;
  wire s_csamul_rca16_and6_9;
  wire s_csamul_rca16_fa6_9_xor0;
  wire s_csamul_rca16_fa6_9_and0;
  wire s_csamul_rca16_fa6_9_xor1;
  wire s_csamul_rca16_fa6_9_and1;
  wire s_csamul_rca16_fa6_9_or0;
  wire s_csamul_rca16_and7_9;
  wire s_csamul_rca16_fa7_9_xor0;
  wire s_csamul_rca16_fa7_9_and0;
  wire s_csamul_rca16_fa7_9_xor1;
  wire s_csamul_rca16_fa7_9_and1;
  wire s_csamul_rca16_fa7_9_or0;
  wire s_csamul_rca16_and8_9;
  wire s_csamul_rca16_fa8_9_xor0;
  wire s_csamul_rca16_fa8_9_and0;
  wire s_csamul_rca16_fa8_9_xor1;
  wire s_csamul_rca16_fa8_9_and1;
  wire s_csamul_rca16_fa8_9_or0;
  wire s_csamul_rca16_and9_9;
  wire s_csamul_rca16_fa9_9_xor0;
  wire s_csamul_rca16_fa9_9_and0;
  wire s_csamul_rca16_fa9_9_xor1;
  wire s_csamul_rca16_fa9_9_and1;
  wire s_csamul_rca16_fa9_9_or0;
  wire s_csamul_rca16_and10_9;
  wire s_csamul_rca16_fa10_9_xor0;
  wire s_csamul_rca16_fa10_9_and0;
  wire s_csamul_rca16_fa10_9_xor1;
  wire s_csamul_rca16_fa10_9_and1;
  wire s_csamul_rca16_fa10_9_or0;
  wire s_csamul_rca16_and11_9;
  wire s_csamul_rca16_fa11_9_xor0;
  wire s_csamul_rca16_fa11_9_and0;
  wire s_csamul_rca16_fa11_9_xor1;
  wire s_csamul_rca16_fa11_9_and1;
  wire s_csamul_rca16_fa11_9_or0;
  wire s_csamul_rca16_and12_9;
  wire s_csamul_rca16_fa12_9_xor0;
  wire s_csamul_rca16_fa12_9_and0;
  wire s_csamul_rca16_fa12_9_xor1;
  wire s_csamul_rca16_fa12_9_and1;
  wire s_csamul_rca16_fa12_9_or0;
  wire s_csamul_rca16_and13_9;
  wire s_csamul_rca16_fa13_9_xor0;
  wire s_csamul_rca16_fa13_9_and0;
  wire s_csamul_rca16_fa13_9_xor1;
  wire s_csamul_rca16_fa13_9_and1;
  wire s_csamul_rca16_fa13_9_or0;
  wire s_csamul_rca16_and14_9;
  wire s_csamul_rca16_fa14_9_xor0;
  wire s_csamul_rca16_fa14_9_and0;
  wire s_csamul_rca16_fa14_9_xor1;
  wire s_csamul_rca16_fa14_9_and1;
  wire s_csamul_rca16_fa14_9_or0;
  wire s_csamul_rca16_nand15_9;
  wire s_csamul_rca16_ha15_9_xor0;
  wire s_csamul_rca16_ha15_9_and0;
  wire s_csamul_rca16_and0_10;
  wire s_csamul_rca16_fa0_10_xor0;
  wire s_csamul_rca16_fa0_10_and0;
  wire s_csamul_rca16_fa0_10_xor1;
  wire s_csamul_rca16_fa0_10_and1;
  wire s_csamul_rca16_fa0_10_or0;
  wire s_csamul_rca16_and1_10;
  wire s_csamul_rca16_fa1_10_xor0;
  wire s_csamul_rca16_fa1_10_and0;
  wire s_csamul_rca16_fa1_10_xor1;
  wire s_csamul_rca16_fa1_10_and1;
  wire s_csamul_rca16_fa1_10_or0;
  wire s_csamul_rca16_and2_10;
  wire s_csamul_rca16_fa2_10_xor0;
  wire s_csamul_rca16_fa2_10_and0;
  wire s_csamul_rca16_fa2_10_xor1;
  wire s_csamul_rca16_fa2_10_and1;
  wire s_csamul_rca16_fa2_10_or0;
  wire s_csamul_rca16_and3_10;
  wire s_csamul_rca16_fa3_10_xor0;
  wire s_csamul_rca16_fa3_10_and0;
  wire s_csamul_rca16_fa3_10_xor1;
  wire s_csamul_rca16_fa3_10_and1;
  wire s_csamul_rca16_fa3_10_or0;
  wire s_csamul_rca16_and4_10;
  wire s_csamul_rca16_fa4_10_xor0;
  wire s_csamul_rca16_fa4_10_and0;
  wire s_csamul_rca16_fa4_10_xor1;
  wire s_csamul_rca16_fa4_10_and1;
  wire s_csamul_rca16_fa4_10_or0;
  wire s_csamul_rca16_and5_10;
  wire s_csamul_rca16_fa5_10_xor0;
  wire s_csamul_rca16_fa5_10_and0;
  wire s_csamul_rca16_fa5_10_xor1;
  wire s_csamul_rca16_fa5_10_and1;
  wire s_csamul_rca16_fa5_10_or0;
  wire s_csamul_rca16_and6_10;
  wire s_csamul_rca16_fa6_10_xor0;
  wire s_csamul_rca16_fa6_10_and0;
  wire s_csamul_rca16_fa6_10_xor1;
  wire s_csamul_rca16_fa6_10_and1;
  wire s_csamul_rca16_fa6_10_or0;
  wire s_csamul_rca16_and7_10;
  wire s_csamul_rca16_fa7_10_xor0;
  wire s_csamul_rca16_fa7_10_and0;
  wire s_csamul_rca16_fa7_10_xor1;
  wire s_csamul_rca16_fa7_10_and1;
  wire s_csamul_rca16_fa7_10_or0;
  wire s_csamul_rca16_and8_10;
  wire s_csamul_rca16_fa8_10_xor0;
  wire s_csamul_rca16_fa8_10_and0;
  wire s_csamul_rca16_fa8_10_xor1;
  wire s_csamul_rca16_fa8_10_and1;
  wire s_csamul_rca16_fa8_10_or0;
  wire s_csamul_rca16_and9_10;
  wire s_csamul_rca16_fa9_10_xor0;
  wire s_csamul_rca16_fa9_10_and0;
  wire s_csamul_rca16_fa9_10_xor1;
  wire s_csamul_rca16_fa9_10_and1;
  wire s_csamul_rca16_fa9_10_or0;
  wire s_csamul_rca16_and10_10;
  wire s_csamul_rca16_fa10_10_xor0;
  wire s_csamul_rca16_fa10_10_and0;
  wire s_csamul_rca16_fa10_10_xor1;
  wire s_csamul_rca16_fa10_10_and1;
  wire s_csamul_rca16_fa10_10_or0;
  wire s_csamul_rca16_and11_10;
  wire s_csamul_rca16_fa11_10_xor0;
  wire s_csamul_rca16_fa11_10_and0;
  wire s_csamul_rca16_fa11_10_xor1;
  wire s_csamul_rca16_fa11_10_and1;
  wire s_csamul_rca16_fa11_10_or0;
  wire s_csamul_rca16_and12_10;
  wire s_csamul_rca16_fa12_10_xor0;
  wire s_csamul_rca16_fa12_10_and0;
  wire s_csamul_rca16_fa12_10_xor1;
  wire s_csamul_rca16_fa12_10_and1;
  wire s_csamul_rca16_fa12_10_or0;
  wire s_csamul_rca16_and13_10;
  wire s_csamul_rca16_fa13_10_xor0;
  wire s_csamul_rca16_fa13_10_and0;
  wire s_csamul_rca16_fa13_10_xor1;
  wire s_csamul_rca16_fa13_10_and1;
  wire s_csamul_rca16_fa13_10_or0;
  wire s_csamul_rca16_and14_10;
  wire s_csamul_rca16_fa14_10_xor0;
  wire s_csamul_rca16_fa14_10_and0;
  wire s_csamul_rca16_fa14_10_xor1;
  wire s_csamul_rca16_fa14_10_and1;
  wire s_csamul_rca16_fa14_10_or0;
  wire s_csamul_rca16_nand15_10;
  wire s_csamul_rca16_ha15_10_xor0;
  wire s_csamul_rca16_ha15_10_and0;
  wire s_csamul_rca16_and0_11;
  wire s_csamul_rca16_fa0_11_xor0;
  wire s_csamul_rca16_fa0_11_and0;
  wire s_csamul_rca16_fa0_11_xor1;
  wire s_csamul_rca16_fa0_11_and1;
  wire s_csamul_rca16_fa0_11_or0;
  wire s_csamul_rca16_and1_11;
  wire s_csamul_rca16_fa1_11_xor0;
  wire s_csamul_rca16_fa1_11_and0;
  wire s_csamul_rca16_fa1_11_xor1;
  wire s_csamul_rca16_fa1_11_and1;
  wire s_csamul_rca16_fa1_11_or0;
  wire s_csamul_rca16_and2_11;
  wire s_csamul_rca16_fa2_11_xor0;
  wire s_csamul_rca16_fa2_11_and0;
  wire s_csamul_rca16_fa2_11_xor1;
  wire s_csamul_rca16_fa2_11_and1;
  wire s_csamul_rca16_fa2_11_or0;
  wire s_csamul_rca16_and3_11;
  wire s_csamul_rca16_fa3_11_xor0;
  wire s_csamul_rca16_fa3_11_and0;
  wire s_csamul_rca16_fa3_11_xor1;
  wire s_csamul_rca16_fa3_11_and1;
  wire s_csamul_rca16_fa3_11_or0;
  wire s_csamul_rca16_and4_11;
  wire s_csamul_rca16_fa4_11_xor0;
  wire s_csamul_rca16_fa4_11_and0;
  wire s_csamul_rca16_fa4_11_xor1;
  wire s_csamul_rca16_fa4_11_and1;
  wire s_csamul_rca16_fa4_11_or0;
  wire s_csamul_rca16_and5_11;
  wire s_csamul_rca16_fa5_11_xor0;
  wire s_csamul_rca16_fa5_11_and0;
  wire s_csamul_rca16_fa5_11_xor1;
  wire s_csamul_rca16_fa5_11_and1;
  wire s_csamul_rca16_fa5_11_or0;
  wire s_csamul_rca16_and6_11;
  wire s_csamul_rca16_fa6_11_xor0;
  wire s_csamul_rca16_fa6_11_and0;
  wire s_csamul_rca16_fa6_11_xor1;
  wire s_csamul_rca16_fa6_11_and1;
  wire s_csamul_rca16_fa6_11_or0;
  wire s_csamul_rca16_and7_11;
  wire s_csamul_rca16_fa7_11_xor0;
  wire s_csamul_rca16_fa7_11_and0;
  wire s_csamul_rca16_fa7_11_xor1;
  wire s_csamul_rca16_fa7_11_and1;
  wire s_csamul_rca16_fa7_11_or0;
  wire s_csamul_rca16_and8_11;
  wire s_csamul_rca16_fa8_11_xor0;
  wire s_csamul_rca16_fa8_11_and0;
  wire s_csamul_rca16_fa8_11_xor1;
  wire s_csamul_rca16_fa8_11_and1;
  wire s_csamul_rca16_fa8_11_or0;
  wire s_csamul_rca16_and9_11;
  wire s_csamul_rca16_fa9_11_xor0;
  wire s_csamul_rca16_fa9_11_and0;
  wire s_csamul_rca16_fa9_11_xor1;
  wire s_csamul_rca16_fa9_11_and1;
  wire s_csamul_rca16_fa9_11_or0;
  wire s_csamul_rca16_and10_11;
  wire s_csamul_rca16_fa10_11_xor0;
  wire s_csamul_rca16_fa10_11_and0;
  wire s_csamul_rca16_fa10_11_xor1;
  wire s_csamul_rca16_fa10_11_and1;
  wire s_csamul_rca16_fa10_11_or0;
  wire s_csamul_rca16_and11_11;
  wire s_csamul_rca16_fa11_11_xor0;
  wire s_csamul_rca16_fa11_11_and0;
  wire s_csamul_rca16_fa11_11_xor1;
  wire s_csamul_rca16_fa11_11_and1;
  wire s_csamul_rca16_fa11_11_or0;
  wire s_csamul_rca16_and12_11;
  wire s_csamul_rca16_fa12_11_xor0;
  wire s_csamul_rca16_fa12_11_and0;
  wire s_csamul_rca16_fa12_11_xor1;
  wire s_csamul_rca16_fa12_11_and1;
  wire s_csamul_rca16_fa12_11_or0;
  wire s_csamul_rca16_and13_11;
  wire s_csamul_rca16_fa13_11_xor0;
  wire s_csamul_rca16_fa13_11_and0;
  wire s_csamul_rca16_fa13_11_xor1;
  wire s_csamul_rca16_fa13_11_and1;
  wire s_csamul_rca16_fa13_11_or0;
  wire s_csamul_rca16_and14_11;
  wire s_csamul_rca16_fa14_11_xor0;
  wire s_csamul_rca16_fa14_11_and0;
  wire s_csamul_rca16_fa14_11_xor1;
  wire s_csamul_rca16_fa14_11_and1;
  wire s_csamul_rca16_fa14_11_or0;
  wire s_csamul_rca16_nand15_11;
  wire s_csamul_rca16_ha15_11_xor0;
  wire s_csamul_rca16_ha15_11_and0;
  wire s_csamul_rca16_and0_12;
  wire s_csamul_rca16_fa0_12_xor0;
  wire s_csamul_rca16_fa0_12_and0;
  wire s_csamul_rca16_fa0_12_xor1;
  wire s_csamul_rca16_fa0_12_and1;
  wire s_csamul_rca16_fa0_12_or0;
  wire s_csamul_rca16_and1_12;
  wire s_csamul_rca16_fa1_12_xor0;
  wire s_csamul_rca16_fa1_12_and0;
  wire s_csamul_rca16_fa1_12_xor1;
  wire s_csamul_rca16_fa1_12_and1;
  wire s_csamul_rca16_fa1_12_or0;
  wire s_csamul_rca16_and2_12;
  wire s_csamul_rca16_fa2_12_xor0;
  wire s_csamul_rca16_fa2_12_and0;
  wire s_csamul_rca16_fa2_12_xor1;
  wire s_csamul_rca16_fa2_12_and1;
  wire s_csamul_rca16_fa2_12_or0;
  wire s_csamul_rca16_and3_12;
  wire s_csamul_rca16_fa3_12_xor0;
  wire s_csamul_rca16_fa3_12_and0;
  wire s_csamul_rca16_fa3_12_xor1;
  wire s_csamul_rca16_fa3_12_and1;
  wire s_csamul_rca16_fa3_12_or0;
  wire s_csamul_rca16_and4_12;
  wire s_csamul_rca16_fa4_12_xor0;
  wire s_csamul_rca16_fa4_12_and0;
  wire s_csamul_rca16_fa4_12_xor1;
  wire s_csamul_rca16_fa4_12_and1;
  wire s_csamul_rca16_fa4_12_or0;
  wire s_csamul_rca16_and5_12;
  wire s_csamul_rca16_fa5_12_xor0;
  wire s_csamul_rca16_fa5_12_and0;
  wire s_csamul_rca16_fa5_12_xor1;
  wire s_csamul_rca16_fa5_12_and1;
  wire s_csamul_rca16_fa5_12_or0;
  wire s_csamul_rca16_and6_12;
  wire s_csamul_rca16_fa6_12_xor0;
  wire s_csamul_rca16_fa6_12_and0;
  wire s_csamul_rca16_fa6_12_xor1;
  wire s_csamul_rca16_fa6_12_and1;
  wire s_csamul_rca16_fa6_12_or0;
  wire s_csamul_rca16_and7_12;
  wire s_csamul_rca16_fa7_12_xor0;
  wire s_csamul_rca16_fa7_12_and0;
  wire s_csamul_rca16_fa7_12_xor1;
  wire s_csamul_rca16_fa7_12_and1;
  wire s_csamul_rca16_fa7_12_or0;
  wire s_csamul_rca16_and8_12;
  wire s_csamul_rca16_fa8_12_xor0;
  wire s_csamul_rca16_fa8_12_and0;
  wire s_csamul_rca16_fa8_12_xor1;
  wire s_csamul_rca16_fa8_12_and1;
  wire s_csamul_rca16_fa8_12_or0;
  wire s_csamul_rca16_and9_12;
  wire s_csamul_rca16_fa9_12_xor0;
  wire s_csamul_rca16_fa9_12_and0;
  wire s_csamul_rca16_fa9_12_xor1;
  wire s_csamul_rca16_fa9_12_and1;
  wire s_csamul_rca16_fa9_12_or0;
  wire s_csamul_rca16_and10_12;
  wire s_csamul_rca16_fa10_12_xor0;
  wire s_csamul_rca16_fa10_12_and0;
  wire s_csamul_rca16_fa10_12_xor1;
  wire s_csamul_rca16_fa10_12_and1;
  wire s_csamul_rca16_fa10_12_or0;
  wire s_csamul_rca16_and11_12;
  wire s_csamul_rca16_fa11_12_xor0;
  wire s_csamul_rca16_fa11_12_and0;
  wire s_csamul_rca16_fa11_12_xor1;
  wire s_csamul_rca16_fa11_12_and1;
  wire s_csamul_rca16_fa11_12_or0;
  wire s_csamul_rca16_and12_12;
  wire s_csamul_rca16_fa12_12_xor0;
  wire s_csamul_rca16_fa12_12_and0;
  wire s_csamul_rca16_fa12_12_xor1;
  wire s_csamul_rca16_fa12_12_and1;
  wire s_csamul_rca16_fa12_12_or0;
  wire s_csamul_rca16_and13_12;
  wire s_csamul_rca16_fa13_12_xor0;
  wire s_csamul_rca16_fa13_12_and0;
  wire s_csamul_rca16_fa13_12_xor1;
  wire s_csamul_rca16_fa13_12_and1;
  wire s_csamul_rca16_fa13_12_or0;
  wire s_csamul_rca16_and14_12;
  wire s_csamul_rca16_fa14_12_xor0;
  wire s_csamul_rca16_fa14_12_and0;
  wire s_csamul_rca16_fa14_12_xor1;
  wire s_csamul_rca16_fa14_12_and1;
  wire s_csamul_rca16_fa14_12_or0;
  wire s_csamul_rca16_nand15_12;
  wire s_csamul_rca16_ha15_12_xor0;
  wire s_csamul_rca16_ha15_12_and0;
  wire s_csamul_rca16_and0_13;
  wire s_csamul_rca16_fa0_13_xor0;
  wire s_csamul_rca16_fa0_13_and0;
  wire s_csamul_rca16_fa0_13_xor1;
  wire s_csamul_rca16_fa0_13_and1;
  wire s_csamul_rca16_fa0_13_or0;
  wire s_csamul_rca16_and1_13;
  wire s_csamul_rca16_fa1_13_xor0;
  wire s_csamul_rca16_fa1_13_and0;
  wire s_csamul_rca16_fa1_13_xor1;
  wire s_csamul_rca16_fa1_13_and1;
  wire s_csamul_rca16_fa1_13_or0;
  wire s_csamul_rca16_and2_13;
  wire s_csamul_rca16_fa2_13_xor0;
  wire s_csamul_rca16_fa2_13_and0;
  wire s_csamul_rca16_fa2_13_xor1;
  wire s_csamul_rca16_fa2_13_and1;
  wire s_csamul_rca16_fa2_13_or0;
  wire s_csamul_rca16_and3_13;
  wire s_csamul_rca16_fa3_13_xor0;
  wire s_csamul_rca16_fa3_13_and0;
  wire s_csamul_rca16_fa3_13_xor1;
  wire s_csamul_rca16_fa3_13_and1;
  wire s_csamul_rca16_fa3_13_or0;
  wire s_csamul_rca16_and4_13;
  wire s_csamul_rca16_fa4_13_xor0;
  wire s_csamul_rca16_fa4_13_and0;
  wire s_csamul_rca16_fa4_13_xor1;
  wire s_csamul_rca16_fa4_13_and1;
  wire s_csamul_rca16_fa4_13_or0;
  wire s_csamul_rca16_and5_13;
  wire s_csamul_rca16_fa5_13_xor0;
  wire s_csamul_rca16_fa5_13_and0;
  wire s_csamul_rca16_fa5_13_xor1;
  wire s_csamul_rca16_fa5_13_and1;
  wire s_csamul_rca16_fa5_13_or0;
  wire s_csamul_rca16_and6_13;
  wire s_csamul_rca16_fa6_13_xor0;
  wire s_csamul_rca16_fa6_13_and0;
  wire s_csamul_rca16_fa6_13_xor1;
  wire s_csamul_rca16_fa6_13_and1;
  wire s_csamul_rca16_fa6_13_or0;
  wire s_csamul_rca16_and7_13;
  wire s_csamul_rca16_fa7_13_xor0;
  wire s_csamul_rca16_fa7_13_and0;
  wire s_csamul_rca16_fa7_13_xor1;
  wire s_csamul_rca16_fa7_13_and1;
  wire s_csamul_rca16_fa7_13_or0;
  wire s_csamul_rca16_and8_13;
  wire s_csamul_rca16_fa8_13_xor0;
  wire s_csamul_rca16_fa8_13_and0;
  wire s_csamul_rca16_fa8_13_xor1;
  wire s_csamul_rca16_fa8_13_and1;
  wire s_csamul_rca16_fa8_13_or0;
  wire s_csamul_rca16_and9_13;
  wire s_csamul_rca16_fa9_13_xor0;
  wire s_csamul_rca16_fa9_13_and0;
  wire s_csamul_rca16_fa9_13_xor1;
  wire s_csamul_rca16_fa9_13_and1;
  wire s_csamul_rca16_fa9_13_or0;
  wire s_csamul_rca16_and10_13;
  wire s_csamul_rca16_fa10_13_xor0;
  wire s_csamul_rca16_fa10_13_and0;
  wire s_csamul_rca16_fa10_13_xor1;
  wire s_csamul_rca16_fa10_13_and1;
  wire s_csamul_rca16_fa10_13_or0;
  wire s_csamul_rca16_and11_13;
  wire s_csamul_rca16_fa11_13_xor0;
  wire s_csamul_rca16_fa11_13_and0;
  wire s_csamul_rca16_fa11_13_xor1;
  wire s_csamul_rca16_fa11_13_and1;
  wire s_csamul_rca16_fa11_13_or0;
  wire s_csamul_rca16_and12_13;
  wire s_csamul_rca16_fa12_13_xor0;
  wire s_csamul_rca16_fa12_13_and0;
  wire s_csamul_rca16_fa12_13_xor1;
  wire s_csamul_rca16_fa12_13_and1;
  wire s_csamul_rca16_fa12_13_or0;
  wire s_csamul_rca16_and13_13;
  wire s_csamul_rca16_fa13_13_xor0;
  wire s_csamul_rca16_fa13_13_and0;
  wire s_csamul_rca16_fa13_13_xor1;
  wire s_csamul_rca16_fa13_13_and1;
  wire s_csamul_rca16_fa13_13_or0;
  wire s_csamul_rca16_and14_13;
  wire s_csamul_rca16_fa14_13_xor0;
  wire s_csamul_rca16_fa14_13_and0;
  wire s_csamul_rca16_fa14_13_xor1;
  wire s_csamul_rca16_fa14_13_and1;
  wire s_csamul_rca16_fa14_13_or0;
  wire s_csamul_rca16_nand15_13;
  wire s_csamul_rca16_ha15_13_xor0;
  wire s_csamul_rca16_ha15_13_and0;
  wire s_csamul_rca16_and0_14;
  wire s_csamul_rca16_fa0_14_xor0;
  wire s_csamul_rca16_fa0_14_and0;
  wire s_csamul_rca16_fa0_14_xor1;
  wire s_csamul_rca16_fa0_14_and1;
  wire s_csamul_rca16_fa0_14_or0;
  wire s_csamul_rca16_and1_14;
  wire s_csamul_rca16_fa1_14_xor0;
  wire s_csamul_rca16_fa1_14_and0;
  wire s_csamul_rca16_fa1_14_xor1;
  wire s_csamul_rca16_fa1_14_and1;
  wire s_csamul_rca16_fa1_14_or0;
  wire s_csamul_rca16_and2_14;
  wire s_csamul_rca16_fa2_14_xor0;
  wire s_csamul_rca16_fa2_14_and0;
  wire s_csamul_rca16_fa2_14_xor1;
  wire s_csamul_rca16_fa2_14_and1;
  wire s_csamul_rca16_fa2_14_or0;
  wire s_csamul_rca16_and3_14;
  wire s_csamul_rca16_fa3_14_xor0;
  wire s_csamul_rca16_fa3_14_and0;
  wire s_csamul_rca16_fa3_14_xor1;
  wire s_csamul_rca16_fa3_14_and1;
  wire s_csamul_rca16_fa3_14_or0;
  wire s_csamul_rca16_and4_14;
  wire s_csamul_rca16_fa4_14_xor0;
  wire s_csamul_rca16_fa4_14_and0;
  wire s_csamul_rca16_fa4_14_xor1;
  wire s_csamul_rca16_fa4_14_and1;
  wire s_csamul_rca16_fa4_14_or0;
  wire s_csamul_rca16_and5_14;
  wire s_csamul_rca16_fa5_14_xor0;
  wire s_csamul_rca16_fa5_14_and0;
  wire s_csamul_rca16_fa5_14_xor1;
  wire s_csamul_rca16_fa5_14_and1;
  wire s_csamul_rca16_fa5_14_or0;
  wire s_csamul_rca16_and6_14;
  wire s_csamul_rca16_fa6_14_xor0;
  wire s_csamul_rca16_fa6_14_and0;
  wire s_csamul_rca16_fa6_14_xor1;
  wire s_csamul_rca16_fa6_14_and1;
  wire s_csamul_rca16_fa6_14_or0;
  wire s_csamul_rca16_and7_14;
  wire s_csamul_rca16_fa7_14_xor0;
  wire s_csamul_rca16_fa7_14_and0;
  wire s_csamul_rca16_fa7_14_xor1;
  wire s_csamul_rca16_fa7_14_and1;
  wire s_csamul_rca16_fa7_14_or0;
  wire s_csamul_rca16_and8_14;
  wire s_csamul_rca16_fa8_14_xor0;
  wire s_csamul_rca16_fa8_14_and0;
  wire s_csamul_rca16_fa8_14_xor1;
  wire s_csamul_rca16_fa8_14_and1;
  wire s_csamul_rca16_fa8_14_or0;
  wire s_csamul_rca16_and9_14;
  wire s_csamul_rca16_fa9_14_xor0;
  wire s_csamul_rca16_fa9_14_and0;
  wire s_csamul_rca16_fa9_14_xor1;
  wire s_csamul_rca16_fa9_14_and1;
  wire s_csamul_rca16_fa9_14_or0;
  wire s_csamul_rca16_and10_14;
  wire s_csamul_rca16_fa10_14_xor0;
  wire s_csamul_rca16_fa10_14_and0;
  wire s_csamul_rca16_fa10_14_xor1;
  wire s_csamul_rca16_fa10_14_and1;
  wire s_csamul_rca16_fa10_14_or0;
  wire s_csamul_rca16_and11_14;
  wire s_csamul_rca16_fa11_14_xor0;
  wire s_csamul_rca16_fa11_14_and0;
  wire s_csamul_rca16_fa11_14_xor1;
  wire s_csamul_rca16_fa11_14_and1;
  wire s_csamul_rca16_fa11_14_or0;
  wire s_csamul_rca16_and12_14;
  wire s_csamul_rca16_fa12_14_xor0;
  wire s_csamul_rca16_fa12_14_and0;
  wire s_csamul_rca16_fa12_14_xor1;
  wire s_csamul_rca16_fa12_14_and1;
  wire s_csamul_rca16_fa12_14_or0;
  wire s_csamul_rca16_and13_14;
  wire s_csamul_rca16_fa13_14_xor0;
  wire s_csamul_rca16_fa13_14_and0;
  wire s_csamul_rca16_fa13_14_xor1;
  wire s_csamul_rca16_fa13_14_and1;
  wire s_csamul_rca16_fa13_14_or0;
  wire s_csamul_rca16_and14_14;
  wire s_csamul_rca16_fa14_14_xor0;
  wire s_csamul_rca16_fa14_14_and0;
  wire s_csamul_rca16_fa14_14_xor1;
  wire s_csamul_rca16_fa14_14_and1;
  wire s_csamul_rca16_fa14_14_or0;
  wire s_csamul_rca16_nand15_14;
  wire s_csamul_rca16_ha15_14_xor0;
  wire s_csamul_rca16_ha15_14_and0;
  wire s_csamul_rca16_nand0_15;
  wire s_csamul_rca16_fa0_15_xor0;
  wire s_csamul_rca16_fa0_15_and0;
  wire s_csamul_rca16_fa0_15_xor1;
  wire s_csamul_rca16_fa0_15_and1;
  wire s_csamul_rca16_fa0_15_or0;
  wire s_csamul_rca16_nand1_15;
  wire s_csamul_rca16_fa1_15_xor0;
  wire s_csamul_rca16_fa1_15_and0;
  wire s_csamul_rca16_fa1_15_xor1;
  wire s_csamul_rca16_fa1_15_and1;
  wire s_csamul_rca16_fa1_15_or0;
  wire s_csamul_rca16_nand2_15;
  wire s_csamul_rca16_fa2_15_xor0;
  wire s_csamul_rca16_fa2_15_and0;
  wire s_csamul_rca16_fa2_15_xor1;
  wire s_csamul_rca16_fa2_15_and1;
  wire s_csamul_rca16_fa2_15_or0;
  wire s_csamul_rca16_nand3_15;
  wire s_csamul_rca16_fa3_15_xor0;
  wire s_csamul_rca16_fa3_15_and0;
  wire s_csamul_rca16_fa3_15_xor1;
  wire s_csamul_rca16_fa3_15_and1;
  wire s_csamul_rca16_fa3_15_or0;
  wire s_csamul_rca16_nand4_15;
  wire s_csamul_rca16_fa4_15_xor0;
  wire s_csamul_rca16_fa4_15_and0;
  wire s_csamul_rca16_fa4_15_xor1;
  wire s_csamul_rca16_fa4_15_and1;
  wire s_csamul_rca16_fa4_15_or0;
  wire s_csamul_rca16_nand5_15;
  wire s_csamul_rca16_fa5_15_xor0;
  wire s_csamul_rca16_fa5_15_and0;
  wire s_csamul_rca16_fa5_15_xor1;
  wire s_csamul_rca16_fa5_15_and1;
  wire s_csamul_rca16_fa5_15_or0;
  wire s_csamul_rca16_nand6_15;
  wire s_csamul_rca16_fa6_15_xor0;
  wire s_csamul_rca16_fa6_15_and0;
  wire s_csamul_rca16_fa6_15_xor1;
  wire s_csamul_rca16_fa6_15_and1;
  wire s_csamul_rca16_fa6_15_or0;
  wire s_csamul_rca16_nand7_15;
  wire s_csamul_rca16_fa7_15_xor0;
  wire s_csamul_rca16_fa7_15_and0;
  wire s_csamul_rca16_fa7_15_xor1;
  wire s_csamul_rca16_fa7_15_and1;
  wire s_csamul_rca16_fa7_15_or0;
  wire s_csamul_rca16_nand8_15;
  wire s_csamul_rca16_fa8_15_xor0;
  wire s_csamul_rca16_fa8_15_and0;
  wire s_csamul_rca16_fa8_15_xor1;
  wire s_csamul_rca16_fa8_15_and1;
  wire s_csamul_rca16_fa8_15_or0;
  wire s_csamul_rca16_nand9_15;
  wire s_csamul_rca16_fa9_15_xor0;
  wire s_csamul_rca16_fa9_15_and0;
  wire s_csamul_rca16_fa9_15_xor1;
  wire s_csamul_rca16_fa9_15_and1;
  wire s_csamul_rca16_fa9_15_or0;
  wire s_csamul_rca16_nand10_15;
  wire s_csamul_rca16_fa10_15_xor0;
  wire s_csamul_rca16_fa10_15_and0;
  wire s_csamul_rca16_fa10_15_xor1;
  wire s_csamul_rca16_fa10_15_and1;
  wire s_csamul_rca16_fa10_15_or0;
  wire s_csamul_rca16_nand11_15;
  wire s_csamul_rca16_fa11_15_xor0;
  wire s_csamul_rca16_fa11_15_and0;
  wire s_csamul_rca16_fa11_15_xor1;
  wire s_csamul_rca16_fa11_15_and1;
  wire s_csamul_rca16_fa11_15_or0;
  wire s_csamul_rca16_nand12_15;
  wire s_csamul_rca16_fa12_15_xor0;
  wire s_csamul_rca16_fa12_15_and0;
  wire s_csamul_rca16_fa12_15_xor1;
  wire s_csamul_rca16_fa12_15_and1;
  wire s_csamul_rca16_fa12_15_or0;
  wire s_csamul_rca16_nand13_15;
  wire s_csamul_rca16_fa13_15_xor0;
  wire s_csamul_rca16_fa13_15_and0;
  wire s_csamul_rca16_fa13_15_xor1;
  wire s_csamul_rca16_fa13_15_and1;
  wire s_csamul_rca16_fa13_15_or0;
  wire s_csamul_rca16_nand14_15;
  wire s_csamul_rca16_fa14_15_xor0;
  wire s_csamul_rca16_fa14_15_and0;
  wire s_csamul_rca16_fa14_15_xor1;
  wire s_csamul_rca16_fa14_15_and1;
  wire s_csamul_rca16_fa14_15_or0;
  wire s_csamul_rca16_and15_15;
  wire s_csamul_rca16_ha15_15_xor0;
  wire s_csamul_rca16_ha15_15_and0;
  wire s_csamul_rca16_u_rca16_ha_xor0;
  wire s_csamul_rca16_u_rca16_ha_and0;
  wire s_csamul_rca16_u_rca16_fa1_xor0;
  wire s_csamul_rca16_u_rca16_fa1_and0;
  wire s_csamul_rca16_u_rca16_fa1_xor1;
  wire s_csamul_rca16_u_rca16_fa1_and1;
  wire s_csamul_rca16_u_rca16_fa1_or0;
  wire s_csamul_rca16_u_rca16_fa2_xor0;
  wire s_csamul_rca16_u_rca16_fa2_and0;
  wire s_csamul_rca16_u_rca16_fa2_xor1;
  wire s_csamul_rca16_u_rca16_fa2_and1;
  wire s_csamul_rca16_u_rca16_fa2_or0;
  wire s_csamul_rca16_u_rca16_fa3_xor0;
  wire s_csamul_rca16_u_rca16_fa3_and0;
  wire s_csamul_rca16_u_rca16_fa3_xor1;
  wire s_csamul_rca16_u_rca16_fa3_and1;
  wire s_csamul_rca16_u_rca16_fa3_or0;
  wire s_csamul_rca16_u_rca16_fa4_xor0;
  wire s_csamul_rca16_u_rca16_fa4_and0;
  wire s_csamul_rca16_u_rca16_fa4_xor1;
  wire s_csamul_rca16_u_rca16_fa4_and1;
  wire s_csamul_rca16_u_rca16_fa4_or0;
  wire s_csamul_rca16_u_rca16_fa5_xor0;
  wire s_csamul_rca16_u_rca16_fa5_and0;
  wire s_csamul_rca16_u_rca16_fa5_xor1;
  wire s_csamul_rca16_u_rca16_fa5_and1;
  wire s_csamul_rca16_u_rca16_fa5_or0;
  wire s_csamul_rca16_u_rca16_fa6_xor0;
  wire s_csamul_rca16_u_rca16_fa6_and0;
  wire s_csamul_rca16_u_rca16_fa6_xor1;
  wire s_csamul_rca16_u_rca16_fa6_and1;
  wire s_csamul_rca16_u_rca16_fa6_or0;
  wire s_csamul_rca16_u_rca16_fa7_xor0;
  wire s_csamul_rca16_u_rca16_fa7_and0;
  wire s_csamul_rca16_u_rca16_fa7_xor1;
  wire s_csamul_rca16_u_rca16_fa7_and1;
  wire s_csamul_rca16_u_rca16_fa7_or0;
  wire s_csamul_rca16_u_rca16_fa8_xor0;
  wire s_csamul_rca16_u_rca16_fa8_and0;
  wire s_csamul_rca16_u_rca16_fa8_xor1;
  wire s_csamul_rca16_u_rca16_fa8_and1;
  wire s_csamul_rca16_u_rca16_fa8_or0;
  wire s_csamul_rca16_u_rca16_fa9_xor0;
  wire s_csamul_rca16_u_rca16_fa9_and0;
  wire s_csamul_rca16_u_rca16_fa9_xor1;
  wire s_csamul_rca16_u_rca16_fa9_and1;
  wire s_csamul_rca16_u_rca16_fa9_or0;
  wire s_csamul_rca16_u_rca16_fa10_xor0;
  wire s_csamul_rca16_u_rca16_fa10_and0;
  wire s_csamul_rca16_u_rca16_fa10_xor1;
  wire s_csamul_rca16_u_rca16_fa10_and1;
  wire s_csamul_rca16_u_rca16_fa10_or0;
  wire s_csamul_rca16_u_rca16_fa11_xor0;
  wire s_csamul_rca16_u_rca16_fa11_and0;
  wire s_csamul_rca16_u_rca16_fa11_xor1;
  wire s_csamul_rca16_u_rca16_fa11_and1;
  wire s_csamul_rca16_u_rca16_fa11_or0;
  wire s_csamul_rca16_u_rca16_fa12_xor0;
  wire s_csamul_rca16_u_rca16_fa12_and0;
  wire s_csamul_rca16_u_rca16_fa12_xor1;
  wire s_csamul_rca16_u_rca16_fa12_and1;
  wire s_csamul_rca16_u_rca16_fa12_or0;
  wire s_csamul_rca16_u_rca16_fa13_xor0;
  wire s_csamul_rca16_u_rca16_fa13_and0;
  wire s_csamul_rca16_u_rca16_fa13_xor1;
  wire s_csamul_rca16_u_rca16_fa13_and1;
  wire s_csamul_rca16_u_rca16_fa13_or0;
  wire s_csamul_rca16_u_rca16_fa14_xor0;
  wire s_csamul_rca16_u_rca16_fa14_and0;
  wire s_csamul_rca16_u_rca16_fa14_xor1;
  wire s_csamul_rca16_u_rca16_fa14_and1;
  wire s_csamul_rca16_u_rca16_fa14_or0;
  wire s_csamul_rca16_u_rca16_fa15_xor0;
  wire s_csamul_rca16_u_rca16_fa15_xor1;
  wire s_csamul_rca16_u_rca16_fa15_and1;
  wire s_csamul_rca16_u_rca16_fa15_or0;

  assign s_csamul_rca16_and0_0 = a[0] & b[0];
  assign s_csamul_rca16_and1_0 = a[1] & b[0];
  assign s_csamul_rca16_and2_0 = a[2] & b[0];
  assign s_csamul_rca16_and3_0 = a[3] & b[0];
  assign s_csamul_rca16_and4_0 = a[4] & b[0];
  assign s_csamul_rca16_and5_0 = a[5] & b[0];
  assign s_csamul_rca16_and6_0 = a[6] & b[0];
  assign s_csamul_rca16_and7_0 = a[7] & b[0];
  assign s_csamul_rca16_and8_0 = a[8] & b[0];
  assign s_csamul_rca16_and9_0 = a[9] & b[0];
  assign s_csamul_rca16_and10_0 = a[10] & b[0];
  assign s_csamul_rca16_and11_0 = a[11] & b[0];
  assign s_csamul_rca16_and12_0 = a[12] & b[0];
  assign s_csamul_rca16_and13_0 = a[13] & b[0];
  assign s_csamul_rca16_and14_0 = a[14] & b[0];
  assign s_csamul_rca16_nand15_0 = ~(a[15] & b[0]);
  assign s_csamul_rca16_and0_1 = a[0] & b[1];
  assign s_csamul_rca16_ha0_1_xor0 = s_csamul_rca16_and0_1 ^ s_csamul_rca16_and1_0;
  assign s_csamul_rca16_ha0_1_and0 = s_csamul_rca16_and0_1 & s_csamul_rca16_and1_0;
  assign s_csamul_rca16_and1_1 = a[1] & b[1];
  assign s_csamul_rca16_ha1_1_xor0 = s_csamul_rca16_and1_1 ^ s_csamul_rca16_and2_0;
  assign s_csamul_rca16_ha1_1_and0 = s_csamul_rca16_and1_1 & s_csamul_rca16_and2_0;
  assign s_csamul_rca16_and2_1 = a[2] & b[1];
  assign s_csamul_rca16_ha2_1_xor0 = s_csamul_rca16_and2_1 ^ s_csamul_rca16_and3_0;
  assign s_csamul_rca16_ha2_1_and0 = s_csamul_rca16_and2_1 & s_csamul_rca16_and3_0;
  assign s_csamul_rca16_and3_1 = a[3] & b[1];
  assign s_csamul_rca16_ha3_1_xor0 = s_csamul_rca16_and3_1 ^ s_csamul_rca16_and4_0;
  assign s_csamul_rca16_ha3_1_and0 = s_csamul_rca16_and3_1 & s_csamul_rca16_and4_0;
  assign s_csamul_rca16_and4_1 = a[4] & b[1];
  assign s_csamul_rca16_ha4_1_xor0 = s_csamul_rca16_and4_1 ^ s_csamul_rca16_and5_0;
  assign s_csamul_rca16_ha4_1_and0 = s_csamul_rca16_and4_1 & s_csamul_rca16_and5_0;
  assign s_csamul_rca16_and5_1 = a[5] & b[1];
  assign s_csamul_rca16_ha5_1_xor0 = s_csamul_rca16_and5_1 ^ s_csamul_rca16_and6_0;
  assign s_csamul_rca16_ha5_1_and0 = s_csamul_rca16_and5_1 & s_csamul_rca16_and6_0;
  assign s_csamul_rca16_and6_1 = a[6] & b[1];
  assign s_csamul_rca16_ha6_1_xor0 = s_csamul_rca16_and6_1 ^ s_csamul_rca16_and7_0;
  assign s_csamul_rca16_ha6_1_and0 = s_csamul_rca16_and6_1 & s_csamul_rca16_and7_0;
  assign s_csamul_rca16_and7_1 = a[7] & b[1];
  assign s_csamul_rca16_ha7_1_xor0 = s_csamul_rca16_and7_1 ^ s_csamul_rca16_and8_0;
  assign s_csamul_rca16_ha7_1_and0 = s_csamul_rca16_and7_1 & s_csamul_rca16_and8_0;
  assign s_csamul_rca16_and8_1 = a[8] & b[1];
  assign s_csamul_rca16_ha8_1_xor0 = s_csamul_rca16_and8_1 ^ s_csamul_rca16_and9_0;
  assign s_csamul_rca16_ha8_1_and0 = s_csamul_rca16_and8_1 & s_csamul_rca16_and9_0;
  assign s_csamul_rca16_and9_1 = a[9] & b[1];
  assign s_csamul_rca16_ha9_1_xor0 = s_csamul_rca16_and9_1 ^ s_csamul_rca16_and10_0;
  assign s_csamul_rca16_ha9_1_and0 = s_csamul_rca16_and9_1 & s_csamul_rca16_and10_0;
  assign s_csamul_rca16_and10_1 = a[10] & b[1];
  assign s_csamul_rca16_ha10_1_xor0 = s_csamul_rca16_and10_1 ^ s_csamul_rca16_and11_0;
  assign s_csamul_rca16_ha10_1_and0 = s_csamul_rca16_and10_1 & s_csamul_rca16_and11_0;
  assign s_csamul_rca16_and11_1 = a[11] & b[1];
  assign s_csamul_rca16_ha11_1_xor0 = s_csamul_rca16_and11_1 ^ s_csamul_rca16_and12_0;
  assign s_csamul_rca16_ha11_1_and0 = s_csamul_rca16_and11_1 & s_csamul_rca16_and12_0;
  assign s_csamul_rca16_and12_1 = a[12] & b[1];
  assign s_csamul_rca16_ha12_1_xor0 = s_csamul_rca16_and12_1 ^ s_csamul_rca16_and13_0;
  assign s_csamul_rca16_ha12_1_and0 = s_csamul_rca16_and12_1 & s_csamul_rca16_and13_0;
  assign s_csamul_rca16_and13_1 = a[13] & b[1];
  assign s_csamul_rca16_ha13_1_xor0 = s_csamul_rca16_and13_1 ^ s_csamul_rca16_and14_0;
  assign s_csamul_rca16_ha13_1_and0 = s_csamul_rca16_and13_1 & s_csamul_rca16_and14_0;
  assign s_csamul_rca16_and14_1 = a[14] & b[1];
  assign s_csamul_rca16_ha14_1_xor0 = s_csamul_rca16_and14_1 ^ s_csamul_rca16_nand15_0;
  assign s_csamul_rca16_ha14_1_and0 = s_csamul_rca16_and14_1 & s_csamul_rca16_nand15_0;
  assign s_csamul_rca16_nand15_1 = ~(a[15] & b[1]);
  assign s_csamul_rca16_ha15_1_xor0 = ~s_csamul_rca16_nand15_1;
  assign s_csamul_rca16_and0_2 = a[0] & b[2];
  assign s_csamul_rca16_fa0_2_xor0 = s_csamul_rca16_and0_2 ^ s_csamul_rca16_ha1_1_xor0;
  assign s_csamul_rca16_fa0_2_and0 = s_csamul_rca16_and0_2 & s_csamul_rca16_ha1_1_xor0;
  assign s_csamul_rca16_fa0_2_xor1 = s_csamul_rca16_fa0_2_xor0 ^ s_csamul_rca16_ha0_1_and0;
  assign s_csamul_rca16_fa0_2_and1 = s_csamul_rca16_fa0_2_xor0 & s_csamul_rca16_ha0_1_and0;
  assign s_csamul_rca16_fa0_2_or0 = s_csamul_rca16_fa0_2_and0 | s_csamul_rca16_fa0_2_and1;
  assign s_csamul_rca16_and1_2 = a[1] & b[2];
  assign s_csamul_rca16_fa1_2_xor0 = s_csamul_rca16_and1_2 ^ s_csamul_rca16_ha2_1_xor0;
  assign s_csamul_rca16_fa1_2_and0 = s_csamul_rca16_and1_2 & s_csamul_rca16_ha2_1_xor0;
  assign s_csamul_rca16_fa1_2_xor1 = s_csamul_rca16_fa1_2_xor0 ^ s_csamul_rca16_ha1_1_and0;
  assign s_csamul_rca16_fa1_2_and1 = s_csamul_rca16_fa1_2_xor0 & s_csamul_rca16_ha1_1_and0;
  assign s_csamul_rca16_fa1_2_or0 = s_csamul_rca16_fa1_2_and0 | s_csamul_rca16_fa1_2_and1;
  assign s_csamul_rca16_and2_2 = a[2] & b[2];
  assign s_csamul_rca16_fa2_2_xor0 = s_csamul_rca16_and2_2 ^ s_csamul_rca16_ha3_1_xor0;
  assign s_csamul_rca16_fa2_2_and0 = s_csamul_rca16_and2_2 & s_csamul_rca16_ha3_1_xor0;
  assign s_csamul_rca16_fa2_2_xor1 = s_csamul_rca16_fa2_2_xor0 ^ s_csamul_rca16_ha2_1_and0;
  assign s_csamul_rca16_fa2_2_and1 = s_csamul_rca16_fa2_2_xor0 & s_csamul_rca16_ha2_1_and0;
  assign s_csamul_rca16_fa2_2_or0 = s_csamul_rca16_fa2_2_and0 | s_csamul_rca16_fa2_2_and1;
  assign s_csamul_rca16_and3_2 = a[3] & b[2];
  assign s_csamul_rca16_fa3_2_xor0 = s_csamul_rca16_and3_2 ^ s_csamul_rca16_ha4_1_xor0;
  assign s_csamul_rca16_fa3_2_and0 = s_csamul_rca16_and3_2 & s_csamul_rca16_ha4_1_xor0;
  assign s_csamul_rca16_fa3_2_xor1 = s_csamul_rca16_fa3_2_xor0 ^ s_csamul_rca16_ha3_1_and0;
  assign s_csamul_rca16_fa3_2_and1 = s_csamul_rca16_fa3_2_xor0 & s_csamul_rca16_ha3_1_and0;
  assign s_csamul_rca16_fa3_2_or0 = s_csamul_rca16_fa3_2_and0 | s_csamul_rca16_fa3_2_and1;
  assign s_csamul_rca16_and4_2 = a[4] & b[2];
  assign s_csamul_rca16_fa4_2_xor0 = s_csamul_rca16_and4_2 ^ s_csamul_rca16_ha5_1_xor0;
  assign s_csamul_rca16_fa4_2_and0 = s_csamul_rca16_and4_2 & s_csamul_rca16_ha5_1_xor0;
  assign s_csamul_rca16_fa4_2_xor1 = s_csamul_rca16_fa4_2_xor0 ^ s_csamul_rca16_ha4_1_and0;
  assign s_csamul_rca16_fa4_2_and1 = s_csamul_rca16_fa4_2_xor0 & s_csamul_rca16_ha4_1_and0;
  assign s_csamul_rca16_fa4_2_or0 = s_csamul_rca16_fa4_2_and0 | s_csamul_rca16_fa4_2_and1;
  assign s_csamul_rca16_and5_2 = a[5] & b[2];
  assign s_csamul_rca16_fa5_2_xor0 = s_csamul_rca16_and5_2 ^ s_csamul_rca16_ha6_1_xor0;
  assign s_csamul_rca16_fa5_2_and0 = s_csamul_rca16_and5_2 & s_csamul_rca16_ha6_1_xor0;
  assign s_csamul_rca16_fa5_2_xor1 = s_csamul_rca16_fa5_2_xor0 ^ s_csamul_rca16_ha5_1_and0;
  assign s_csamul_rca16_fa5_2_and1 = s_csamul_rca16_fa5_2_xor0 & s_csamul_rca16_ha5_1_and0;
  assign s_csamul_rca16_fa5_2_or0 = s_csamul_rca16_fa5_2_and0 | s_csamul_rca16_fa5_2_and1;
  assign s_csamul_rca16_and6_2 = a[6] & b[2];
  assign s_csamul_rca16_fa6_2_xor0 = s_csamul_rca16_and6_2 ^ s_csamul_rca16_ha7_1_xor0;
  assign s_csamul_rca16_fa6_2_and0 = s_csamul_rca16_and6_2 & s_csamul_rca16_ha7_1_xor0;
  assign s_csamul_rca16_fa6_2_xor1 = s_csamul_rca16_fa6_2_xor0 ^ s_csamul_rca16_ha6_1_and0;
  assign s_csamul_rca16_fa6_2_and1 = s_csamul_rca16_fa6_2_xor0 & s_csamul_rca16_ha6_1_and0;
  assign s_csamul_rca16_fa6_2_or0 = s_csamul_rca16_fa6_2_and0 | s_csamul_rca16_fa6_2_and1;
  assign s_csamul_rca16_and7_2 = a[7] & b[2];
  assign s_csamul_rca16_fa7_2_xor0 = s_csamul_rca16_and7_2 ^ s_csamul_rca16_ha8_1_xor0;
  assign s_csamul_rca16_fa7_2_and0 = s_csamul_rca16_and7_2 & s_csamul_rca16_ha8_1_xor0;
  assign s_csamul_rca16_fa7_2_xor1 = s_csamul_rca16_fa7_2_xor0 ^ s_csamul_rca16_ha7_1_and0;
  assign s_csamul_rca16_fa7_2_and1 = s_csamul_rca16_fa7_2_xor0 & s_csamul_rca16_ha7_1_and0;
  assign s_csamul_rca16_fa7_2_or0 = s_csamul_rca16_fa7_2_and0 | s_csamul_rca16_fa7_2_and1;
  assign s_csamul_rca16_and8_2 = a[8] & b[2];
  assign s_csamul_rca16_fa8_2_xor0 = s_csamul_rca16_and8_2 ^ s_csamul_rca16_ha9_1_xor0;
  assign s_csamul_rca16_fa8_2_and0 = s_csamul_rca16_and8_2 & s_csamul_rca16_ha9_1_xor0;
  assign s_csamul_rca16_fa8_2_xor1 = s_csamul_rca16_fa8_2_xor0 ^ s_csamul_rca16_ha8_1_and0;
  assign s_csamul_rca16_fa8_2_and1 = s_csamul_rca16_fa8_2_xor0 & s_csamul_rca16_ha8_1_and0;
  assign s_csamul_rca16_fa8_2_or0 = s_csamul_rca16_fa8_2_and0 | s_csamul_rca16_fa8_2_and1;
  assign s_csamul_rca16_and9_2 = a[9] & b[2];
  assign s_csamul_rca16_fa9_2_xor0 = s_csamul_rca16_and9_2 ^ s_csamul_rca16_ha10_1_xor0;
  assign s_csamul_rca16_fa9_2_and0 = s_csamul_rca16_and9_2 & s_csamul_rca16_ha10_1_xor0;
  assign s_csamul_rca16_fa9_2_xor1 = s_csamul_rca16_fa9_2_xor0 ^ s_csamul_rca16_ha9_1_and0;
  assign s_csamul_rca16_fa9_2_and1 = s_csamul_rca16_fa9_2_xor0 & s_csamul_rca16_ha9_1_and0;
  assign s_csamul_rca16_fa9_2_or0 = s_csamul_rca16_fa9_2_and0 | s_csamul_rca16_fa9_2_and1;
  assign s_csamul_rca16_and10_2 = a[10] & b[2];
  assign s_csamul_rca16_fa10_2_xor0 = s_csamul_rca16_and10_2 ^ s_csamul_rca16_ha11_1_xor0;
  assign s_csamul_rca16_fa10_2_and0 = s_csamul_rca16_and10_2 & s_csamul_rca16_ha11_1_xor0;
  assign s_csamul_rca16_fa10_2_xor1 = s_csamul_rca16_fa10_2_xor0 ^ s_csamul_rca16_ha10_1_and0;
  assign s_csamul_rca16_fa10_2_and1 = s_csamul_rca16_fa10_2_xor0 & s_csamul_rca16_ha10_1_and0;
  assign s_csamul_rca16_fa10_2_or0 = s_csamul_rca16_fa10_2_and0 | s_csamul_rca16_fa10_2_and1;
  assign s_csamul_rca16_and11_2 = a[11] & b[2];
  assign s_csamul_rca16_fa11_2_xor0 = s_csamul_rca16_and11_2 ^ s_csamul_rca16_ha12_1_xor0;
  assign s_csamul_rca16_fa11_2_and0 = s_csamul_rca16_and11_2 & s_csamul_rca16_ha12_1_xor0;
  assign s_csamul_rca16_fa11_2_xor1 = s_csamul_rca16_fa11_2_xor0 ^ s_csamul_rca16_ha11_1_and0;
  assign s_csamul_rca16_fa11_2_and1 = s_csamul_rca16_fa11_2_xor0 & s_csamul_rca16_ha11_1_and0;
  assign s_csamul_rca16_fa11_2_or0 = s_csamul_rca16_fa11_2_and0 | s_csamul_rca16_fa11_2_and1;
  assign s_csamul_rca16_and12_2 = a[12] & b[2];
  assign s_csamul_rca16_fa12_2_xor0 = s_csamul_rca16_and12_2 ^ s_csamul_rca16_ha13_1_xor0;
  assign s_csamul_rca16_fa12_2_and0 = s_csamul_rca16_and12_2 & s_csamul_rca16_ha13_1_xor0;
  assign s_csamul_rca16_fa12_2_xor1 = s_csamul_rca16_fa12_2_xor0 ^ s_csamul_rca16_ha12_1_and0;
  assign s_csamul_rca16_fa12_2_and1 = s_csamul_rca16_fa12_2_xor0 & s_csamul_rca16_ha12_1_and0;
  assign s_csamul_rca16_fa12_2_or0 = s_csamul_rca16_fa12_2_and0 | s_csamul_rca16_fa12_2_and1;
  assign s_csamul_rca16_and13_2 = a[13] & b[2];
  assign s_csamul_rca16_fa13_2_xor0 = s_csamul_rca16_and13_2 ^ s_csamul_rca16_ha14_1_xor0;
  assign s_csamul_rca16_fa13_2_and0 = s_csamul_rca16_and13_2 & s_csamul_rca16_ha14_1_xor0;
  assign s_csamul_rca16_fa13_2_xor1 = s_csamul_rca16_fa13_2_xor0 ^ s_csamul_rca16_ha13_1_and0;
  assign s_csamul_rca16_fa13_2_and1 = s_csamul_rca16_fa13_2_xor0 & s_csamul_rca16_ha13_1_and0;
  assign s_csamul_rca16_fa13_2_or0 = s_csamul_rca16_fa13_2_and0 | s_csamul_rca16_fa13_2_and1;
  assign s_csamul_rca16_and14_2 = a[14] & b[2];
  assign s_csamul_rca16_fa14_2_xor0 = s_csamul_rca16_and14_2 ^ s_csamul_rca16_ha15_1_xor0;
  assign s_csamul_rca16_fa14_2_and0 = s_csamul_rca16_and14_2 & s_csamul_rca16_ha15_1_xor0;
  assign s_csamul_rca16_fa14_2_xor1 = s_csamul_rca16_fa14_2_xor0 ^ s_csamul_rca16_ha14_1_and0;
  assign s_csamul_rca16_fa14_2_and1 = s_csamul_rca16_fa14_2_xor0 & s_csamul_rca16_ha14_1_and0;
  assign s_csamul_rca16_fa14_2_or0 = s_csamul_rca16_fa14_2_and0 | s_csamul_rca16_fa14_2_and1;
  assign s_csamul_rca16_nand15_2 = ~(a[15] & b[2]);
  assign s_csamul_rca16_ha15_2_xor0 = s_csamul_rca16_nand15_2 ^ s_csamul_rca16_nand15_1;
  assign s_csamul_rca16_ha15_2_and0 = s_csamul_rca16_nand15_2 & s_csamul_rca16_nand15_1;
  assign s_csamul_rca16_and0_3 = a[0] & b[3];
  assign s_csamul_rca16_fa0_3_xor0 = s_csamul_rca16_and0_3 ^ s_csamul_rca16_fa1_2_xor1;
  assign s_csamul_rca16_fa0_3_and0 = s_csamul_rca16_and0_3 & s_csamul_rca16_fa1_2_xor1;
  assign s_csamul_rca16_fa0_3_xor1 = s_csamul_rca16_fa0_3_xor0 ^ s_csamul_rca16_fa0_2_or0;
  assign s_csamul_rca16_fa0_3_and1 = s_csamul_rca16_fa0_3_xor0 & s_csamul_rca16_fa0_2_or0;
  assign s_csamul_rca16_fa0_3_or0 = s_csamul_rca16_fa0_3_and0 | s_csamul_rca16_fa0_3_and1;
  assign s_csamul_rca16_and1_3 = a[1] & b[3];
  assign s_csamul_rca16_fa1_3_xor0 = s_csamul_rca16_and1_3 ^ s_csamul_rca16_fa2_2_xor1;
  assign s_csamul_rca16_fa1_3_and0 = s_csamul_rca16_and1_3 & s_csamul_rca16_fa2_2_xor1;
  assign s_csamul_rca16_fa1_3_xor1 = s_csamul_rca16_fa1_3_xor0 ^ s_csamul_rca16_fa1_2_or0;
  assign s_csamul_rca16_fa1_3_and1 = s_csamul_rca16_fa1_3_xor0 & s_csamul_rca16_fa1_2_or0;
  assign s_csamul_rca16_fa1_3_or0 = s_csamul_rca16_fa1_3_and0 | s_csamul_rca16_fa1_3_and1;
  assign s_csamul_rca16_and2_3 = a[2] & b[3];
  assign s_csamul_rca16_fa2_3_xor0 = s_csamul_rca16_and2_3 ^ s_csamul_rca16_fa3_2_xor1;
  assign s_csamul_rca16_fa2_3_and0 = s_csamul_rca16_and2_3 & s_csamul_rca16_fa3_2_xor1;
  assign s_csamul_rca16_fa2_3_xor1 = s_csamul_rca16_fa2_3_xor0 ^ s_csamul_rca16_fa2_2_or0;
  assign s_csamul_rca16_fa2_3_and1 = s_csamul_rca16_fa2_3_xor0 & s_csamul_rca16_fa2_2_or0;
  assign s_csamul_rca16_fa2_3_or0 = s_csamul_rca16_fa2_3_and0 | s_csamul_rca16_fa2_3_and1;
  assign s_csamul_rca16_and3_3 = a[3] & b[3];
  assign s_csamul_rca16_fa3_3_xor0 = s_csamul_rca16_and3_3 ^ s_csamul_rca16_fa4_2_xor1;
  assign s_csamul_rca16_fa3_3_and0 = s_csamul_rca16_and3_3 & s_csamul_rca16_fa4_2_xor1;
  assign s_csamul_rca16_fa3_3_xor1 = s_csamul_rca16_fa3_3_xor0 ^ s_csamul_rca16_fa3_2_or0;
  assign s_csamul_rca16_fa3_3_and1 = s_csamul_rca16_fa3_3_xor0 & s_csamul_rca16_fa3_2_or0;
  assign s_csamul_rca16_fa3_3_or0 = s_csamul_rca16_fa3_3_and0 | s_csamul_rca16_fa3_3_and1;
  assign s_csamul_rca16_and4_3 = a[4] & b[3];
  assign s_csamul_rca16_fa4_3_xor0 = s_csamul_rca16_and4_3 ^ s_csamul_rca16_fa5_2_xor1;
  assign s_csamul_rca16_fa4_3_and0 = s_csamul_rca16_and4_3 & s_csamul_rca16_fa5_2_xor1;
  assign s_csamul_rca16_fa4_3_xor1 = s_csamul_rca16_fa4_3_xor0 ^ s_csamul_rca16_fa4_2_or0;
  assign s_csamul_rca16_fa4_3_and1 = s_csamul_rca16_fa4_3_xor0 & s_csamul_rca16_fa4_2_or0;
  assign s_csamul_rca16_fa4_3_or0 = s_csamul_rca16_fa4_3_and0 | s_csamul_rca16_fa4_3_and1;
  assign s_csamul_rca16_and5_3 = a[5] & b[3];
  assign s_csamul_rca16_fa5_3_xor0 = s_csamul_rca16_and5_3 ^ s_csamul_rca16_fa6_2_xor1;
  assign s_csamul_rca16_fa5_3_and0 = s_csamul_rca16_and5_3 & s_csamul_rca16_fa6_2_xor1;
  assign s_csamul_rca16_fa5_3_xor1 = s_csamul_rca16_fa5_3_xor0 ^ s_csamul_rca16_fa5_2_or0;
  assign s_csamul_rca16_fa5_3_and1 = s_csamul_rca16_fa5_3_xor0 & s_csamul_rca16_fa5_2_or0;
  assign s_csamul_rca16_fa5_3_or0 = s_csamul_rca16_fa5_3_and0 | s_csamul_rca16_fa5_3_and1;
  assign s_csamul_rca16_and6_3 = a[6] & b[3];
  assign s_csamul_rca16_fa6_3_xor0 = s_csamul_rca16_and6_3 ^ s_csamul_rca16_fa7_2_xor1;
  assign s_csamul_rca16_fa6_3_and0 = s_csamul_rca16_and6_3 & s_csamul_rca16_fa7_2_xor1;
  assign s_csamul_rca16_fa6_3_xor1 = s_csamul_rca16_fa6_3_xor0 ^ s_csamul_rca16_fa6_2_or0;
  assign s_csamul_rca16_fa6_3_and1 = s_csamul_rca16_fa6_3_xor0 & s_csamul_rca16_fa6_2_or0;
  assign s_csamul_rca16_fa6_3_or0 = s_csamul_rca16_fa6_3_and0 | s_csamul_rca16_fa6_3_and1;
  assign s_csamul_rca16_and7_3 = a[7] & b[3];
  assign s_csamul_rca16_fa7_3_xor0 = s_csamul_rca16_and7_3 ^ s_csamul_rca16_fa8_2_xor1;
  assign s_csamul_rca16_fa7_3_and0 = s_csamul_rca16_and7_3 & s_csamul_rca16_fa8_2_xor1;
  assign s_csamul_rca16_fa7_3_xor1 = s_csamul_rca16_fa7_3_xor0 ^ s_csamul_rca16_fa7_2_or0;
  assign s_csamul_rca16_fa7_3_and1 = s_csamul_rca16_fa7_3_xor0 & s_csamul_rca16_fa7_2_or0;
  assign s_csamul_rca16_fa7_3_or0 = s_csamul_rca16_fa7_3_and0 | s_csamul_rca16_fa7_3_and1;
  assign s_csamul_rca16_and8_3 = a[8] & b[3];
  assign s_csamul_rca16_fa8_3_xor0 = s_csamul_rca16_and8_3 ^ s_csamul_rca16_fa9_2_xor1;
  assign s_csamul_rca16_fa8_3_and0 = s_csamul_rca16_and8_3 & s_csamul_rca16_fa9_2_xor1;
  assign s_csamul_rca16_fa8_3_xor1 = s_csamul_rca16_fa8_3_xor0 ^ s_csamul_rca16_fa8_2_or0;
  assign s_csamul_rca16_fa8_3_and1 = s_csamul_rca16_fa8_3_xor0 & s_csamul_rca16_fa8_2_or0;
  assign s_csamul_rca16_fa8_3_or0 = s_csamul_rca16_fa8_3_and0 | s_csamul_rca16_fa8_3_and1;
  assign s_csamul_rca16_and9_3 = a[9] & b[3];
  assign s_csamul_rca16_fa9_3_xor0 = s_csamul_rca16_and9_3 ^ s_csamul_rca16_fa10_2_xor1;
  assign s_csamul_rca16_fa9_3_and0 = s_csamul_rca16_and9_3 & s_csamul_rca16_fa10_2_xor1;
  assign s_csamul_rca16_fa9_3_xor1 = s_csamul_rca16_fa9_3_xor0 ^ s_csamul_rca16_fa9_2_or0;
  assign s_csamul_rca16_fa9_3_and1 = s_csamul_rca16_fa9_3_xor0 & s_csamul_rca16_fa9_2_or0;
  assign s_csamul_rca16_fa9_3_or0 = s_csamul_rca16_fa9_3_and0 | s_csamul_rca16_fa9_3_and1;
  assign s_csamul_rca16_and10_3 = a[10] & b[3];
  assign s_csamul_rca16_fa10_3_xor0 = s_csamul_rca16_and10_3 ^ s_csamul_rca16_fa11_2_xor1;
  assign s_csamul_rca16_fa10_3_and0 = s_csamul_rca16_and10_3 & s_csamul_rca16_fa11_2_xor1;
  assign s_csamul_rca16_fa10_3_xor1 = s_csamul_rca16_fa10_3_xor0 ^ s_csamul_rca16_fa10_2_or0;
  assign s_csamul_rca16_fa10_3_and1 = s_csamul_rca16_fa10_3_xor0 & s_csamul_rca16_fa10_2_or0;
  assign s_csamul_rca16_fa10_3_or0 = s_csamul_rca16_fa10_3_and0 | s_csamul_rca16_fa10_3_and1;
  assign s_csamul_rca16_and11_3 = a[11] & b[3];
  assign s_csamul_rca16_fa11_3_xor0 = s_csamul_rca16_and11_3 ^ s_csamul_rca16_fa12_2_xor1;
  assign s_csamul_rca16_fa11_3_and0 = s_csamul_rca16_and11_3 & s_csamul_rca16_fa12_2_xor1;
  assign s_csamul_rca16_fa11_3_xor1 = s_csamul_rca16_fa11_3_xor0 ^ s_csamul_rca16_fa11_2_or0;
  assign s_csamul_rca16_fa11_3_and1 = s_csamul_rca16_fa11_3_xor0 & s_csamul_rca16_fa11_2_or0;
  assign s_csamul_rca16_fa11_3_or0 = s_csamul_rca16_fa11_3_and0 | s_csamul_rca16_fa11_3_and1;
  assign s_csamul_rca16_and12_3 = a[12] & b[3];
  assign s_csamul_rca16_fa12_3_xor0 = s_csamul_rca16_and12_3 ^ s_csamul_rca16_fa13_2_xor1;
  assign s_csamul_rca16_fa12_3_and0 = s_csamul_rca16_and12_3 & s_csamul_rca16_fa13_2_xor1;
  assign s_csamul_rca16_fa12_3_xor1 = s_csamul_rca16_fa12_3_xor0 ^ s_csamul_rca16_fa12_2_or0;
  assign s_csamul_rca16_fa12_3_and1 = s_csamul_rca16_fa12_3_xor0 & s_csamul_rca16_fa12_2_or0;
  assign s_csamul_rca16_fa12_3_or0 = s_csamul_rca16_fa12_3_and0 | s_csamul_rca16_fa12_3_and1;
  assign s_csamul_rca16_and13_3 = a[13] & b[3];
  assign s_csamul_rca16_fa13_3_xor0 = s_csamul_rca16_and13_3 ^ s_csamul_rca16_fa14_2_xor1;
  assign s_csamul_rca16_fa13_3_and0 = s_csamul_rca16_and13_3 & s_csamul_rca16_fa14_2_xor1;
  assign s_csamul_rca16_fa13_3_xor1 = s_csamul_rca16_fa13_3_xor0 ^ s_csamul_rca16_fa13_2_or0;
  assign s_csamul_rca16_fa13_3_and1 = s_csamul_rca16_fa13_3_xor0 & s_csamul_rca16_fa13_2_or0;
  assign s_csamul_rca16_fa13_3_or0 = s_csamul_rca16_fa13_3_and0 | s_csamul_rca16_fa13_3_and1;
  assign s_csamul_rca16_and14_3 = a[14] & b[3];
  assign s_csamul_rca16_fa14_3_xor0 = s_csamul_rca16_and14_3 ^ s_csamul_rca16_ha15_2_xor0;
  assign s_csamul_rca16_fa14_3_and0 = s_csamul_rca16_and14_3 & s_csamul_rca16_ha15_2_xor0;
  assign s_csamul_rca16_fa14_3_xor1 = s_csamul_rca16_fa14_3_xor0 ^ s_csamul_rca16_fa14_2_or0;
  assign s_csamul_rca16_fa14_3_and1 = s_csamul_rca16_fa14_3_xor0 & s_csamul_rca16_fa14_2_or0;
  assign s_csamul_rca16_fa14_3_or0 = s_csamul_rca16_fa14_3_and0 | s_csamul_rca16_fa14_3_and1;
  assign s_csamul_rca16_nand15_3 = ~(a[15] & b[3]);
  assign s_csamul_rca16_ha15_3_xor0 = s_csamul_rca16_nand15_3 ^ s_csamul_rca16_ha15_2_and0;
  assign s_csamul_rca16_ha15_3_and0 = s_csamul_rca16_nand15_3 & s_csamul_rca16_ha15_2_and0;
  assign s_csamul_rca16_and0_4 = a[0] & b[4];
  assign s_csamul_rca16_fa0_4_xor0 = s_csamul_rca16_and0_4 ^ s_csamul_rca16_fa1_3_xor1;
  assign s_csamul_rca16_fa0_4_and0 = s_csamul_rca16_and0_4 & s_csamul_rca16_fa1_3_xor1;
  assign s_csamul_rca16_fa0_4_xor1 = s_csamul_rca16_fa0_4_xor0 ^ s_csamul_rca16_fa0_3_or0;
  assign s_csamul_rca16_fa0_4_and1 = s_csamul_rca16_fa0_4_xor0 & s_csamul_rca16_fa0_3_or0;
  assign s_csamul_rca16_fa0_4_or0 = s_csamul_rca16_fa0_4_and0 | s_csamul_rca16_fa0_4_and1;
  assign s_csamul_rca16_and1_4 = a[1] & b[4];
  assign s_csamul_rca16_fa1_4_xor0 = s_csamul_rca16_and1_4 ^ s_csamul_rca16_fa2_3_xor1;
  assign s_csamul_rca16_fa1_4_and0 = s_csamul_rca16_and1_4 & s_csamul_rca16_fa2_3_xor1;
  assign s_csamul_rca16_fa1_4_xor1 = s_csamul_rca16_fa1_4_xor0 ^ s_csamul_rca16_fa1_3_or0;
  assign s_csamul_rca16_fa1_4_and1 = s_csamul_rca16_fa1_4_xor0 & s_csamul_rca16_fa1_3_or0;
  assign s_csamul_rca16_fa1_4_or0 = s_csamul_rca16_fa1_4_and0 | s_csamul_rca16_fa1_4_and1;
  assign s_csamul_rca16_and2_4 = a[2] & b[4];
  assign s_csamul_rca16_fa2_4_xor0 = s_csamul_rca16_and2_4 ^ s_csamul_rca16_fa3_3_xor1;
  assign s_csamul_rca16_fa2_4_and0 = s_csamul_rca16_and2_4 & s_csamul_rca16_fa3_3_xor1;
  assign s_csamul_rca16_fa2_4_xor1 = s_csamul_rca16_fa2_4_xor0 ^ s_csamul_rca16_fa2_3_or0;
  assign s_csamul_rca16_fa2_4_and1 = s_csamul_rca16_fa2_4_xor0 & s_csamul_rca16_fa2_3_or0;
  assign s_csamul_rca16_fa2_4_or0 = s_csamul_rca16_fa2_4_and0 | s_csamul_rca16_fa2_4_and1;
  assign s_csamul_rca16_and3_4 = a[3] & b[4];
  assign s_csamul_rca16_fa3_4_xor0 = s_csamul_rca16_and3_4 ^ s_csamul_rca16_fa4_3_xor1;
  assign s_csamul_rca16_fa3_4_and0 = s_csamul_rca16_and3_4 & s_csamul_rca16_fa4_3_xor1;
  assign s_csamul_rca16_fa3_4_xor1 = s_csamul_rca16_fa3_4_xor0 ^ s_csamul_rca16_fa3_3_or0;
  assign s_csamul_rca16_fa3_4_and1 = s_csamul_rca16_fa3_4_xor0 & s_csamul_rca16_fa3_3_or0;
  assign s_csamul_rca16_fa3_4_or0 = s_csamul_rca16_fa3_4_and0 | s_csamul_rca16_fa3_4_and1;
  assign s_csamul_rca16_and4_4 = a[4] & b[4];
  assign s_csamul_rca16_fa4_4_xor0 = s_csamul_rca16_and4_4 ^ s_csamul_rca16_fa5_3_xor1;
  assign s_csamul_rca16_fa4_4_and0 = s_csamul_rca16_and4_4 & s_csamul_rca16_fa5_3_xor1;
  assign s_csamul_rca16_fa4_4_xor1 = s_csamul_rca16_fa4_4_xor0 ^ s_csamul_rca16_fa4_3_or0;
  assign s_csamul_rca16_fa4_4_and1 = s_csamul_rca16_fa4_4_xor0 & s_csamul_rca16_fa4_3_or0;
  assign s_csamul_rca16_fa4_4_or0 = s_csamul_rca16_fa4_4_and0 | s_csamul_rca16_fa4_4_and1;
  assign s_csamul_rca16_and5_4 = a[5] & b[4];
  assign s_csamul_rca16_fa5_4_xor0 = s_csamul_rca16_and5_4 ^ s_csamul_rca16_fa6_3_xor1;
  assign s_csamul_rca16_fa5_4_and0 = s_csamul_rca16_and5_4 & s_csamul_rca16_fa6_3_xor1;
  assign s_csamul_rca16_fa5_4_xor1 = s_csamul_rca16_fa5_4_xor0 ^ s_csamul_rca16_fa5_3_or0;
  assign s_csamul_rca16_fa5_4_and1 = s_csamul_rca16_fa5_4_xor0 & s_csamul_rca16_fa5_3_or0;
  assign s_csamul_rca16_fa5_4_or0 = s_csamul_rca16_fa5_4_and0 | s_csamul_rca16_fa5_4_and1;
  assign s_csamul_rca16_and6_4 = a[6] & b[4];
  assign s_csamul_rca16_fa6_4_xor0 = s_csamul_rca16_and6_4 ^ s_csamul_rca16_fa7_3_xor1;
  assign s_csamul_rca16_fa6_4_and0 = s_csamul_rca16_and6_4 & s_csamul_rca16_fa7_3_xor1;
  assign s_csamul_rca16_fa6_4_xor1 = s_csamul_rca16_fa6_4_xor0 ^ s_csamul_rca16_fa6_3_or0;
  assign s_csamul_rca16_fa6_4_and1 = s_csamul_rca16_fa6_4_xor0 & s_csamul_rca16_fa6_3_or0;
  assign s_csamul_rca16_fa6_4_or0 = s_csamul_rca16_fa6_4_and0 | s_csamul_rca16_fa6_4_and1;
  assign s_csamul_rca16_and7_4 = a[7] & b[4];
  assign s_csamul_rca16_fa7_4_xor0 = s_csamul_rca16_and7_4 ^ s_csamul_rca16_fa8_3_xor1;
  assign s_csamul_rca16_fa7_4_and0 = s_csamul_rca16_and7_4 & s_csamul_rca16_fa8_3_xor1;
  assign s_csamul_rca16_fa7_4_xor1 = s_csamul_rca16_fa7_4_xor0 ^ s_csamul_rca16_fa7_3_or0;
  assign s_csamul_rca16_fa7_4_and1 = s_csamul_rca16_fa7_4_xor0 & s_csamul_rca16_fa7_3_or0;
  assign s_csamul_rca16_fa7_4_or0 = s_csamul_rca16_fa7_4_and0 | s_csamul_rca16_fa7_4_and1;
  assign s_csamul_rca16_and8_4 = a[8] & b[4];
  assign s_csamul_rca16_fa8_4_xor0 = s_csamul_rca16_and8_4 ^ s_csamul_rca16_fa9_3_xor1;
  assign s_csamul_rca16_fa8_4_and0 = s_csamul_rca16_and8_4 & s_csamul_rca16_fa9_3_xor1;
  assign s_csamul_rca16_fa8_4_xor1 = s_csamul_rca16_fa8_4_xor0 ^ s_csamul_rca16_fa8_3_or0;
  assign s_csamul_rca16_fa8_4_and1 = s_csamul_rca16_fa8_4_xor0 & s_csamul_rca16_fa8_3_or0;
  assign s_csamul_rca16_fa8_4_or0 = s_csamul_rca16_fa8_4_and0 | s_csamul_rca16_fa8_4_and1;
  assign s_csamul_rca16_and9_4 = a[9] & b[4];
  assign s_csamul_rca16_fa9_4_xor0 = s_csamul_rca16_and9_4 ^ s_csamul_rca16_fa10_3_xor1;
  assign s_csamul_rca16_fa9_4_and0 = s_csamul_rca16_and9_4 & s_csamul_rca16_fa10_3_xor1;
  assign s_csamul_rca16_fa9_4_xor1 = s_csamul_rca16_fa9_4_xor0 ^ s_csamul_rca16_fa9_3_or0;
  assign s_csamul_rca16_fa9_4_and1 = s_csamul_rca16_fa9_4_xor0 & s_csamul_rca16_fa9_3_or0;
  assign s_csamul_rca16_fa9_4_or0 = s_csamul_rca16_fa9_4_and0 | s_csamul_rca16_fa9_4_and1;
  assign s_csamul_rca16_and10_4 = a[10] & b[4];
  assign s_csamul_rca16_fa10_4_xor0 = s_csamul_rca16_and10_4 ^ s_csamul_rca16_fa11_3_xor1;
  assign s_csamul_rca16_fa10_4_and0 = s_csamul_rca16_and10_4 & s_csamul_rca16_fa11_3_xor1;
  assign s_csamul_rca16_fa10_4_xor1 = s_csamul_rca16_fa10_4_xor0 ^ s_csamul_rca16_fa10_3_or0;
  assign s_csamul_rca16_fa10_4_and1 = s_csamul_rca16_fa10_4_xor0 & s_csamul_rca16_fa10_3_or0;
  assign s_csamul_rca16_fa10_4_or0 = s_csamul_rca16_fa10_4_and0 | s_csamul_rca16_fa10_4_and1;
  assign s_csamul_rca16_and11_4 = a[11] & b[4];
  assign s_csamul_rca16_fa11_4_xor0 = s_csamul_rca16_and11_4 ^ s_csamul_rca16_fa12_3_xor1;
  assign s_csamul_rca16_fa11_4_and0 = s_csamul_rca16_and11_4 & s_csamul_rca16_fa12_3_xor1;
  assign s_csamul_rca16_fa11_4_xor1 = s_csamul_rca16_fa11_4_xor0 ^ s_csamul_rca16_fa11_3_or0;
  assign s_csamul_rca16_fa11_4_and1 = s_csamul_rca16_fa11_4_xor0 & s_csamul_rca16_fa11_3_or0;
  assign s_csamul_rca16_fa11_4_or0 = s_csamul_rca16_fa11_4_and0 | s_csamul_rca16_fa11_4_and1;
  assign s_csamul_rca16_and12_4 = a[12] & b[4];
  assign s_csamul_rca16_fa12_4_xor0 = s_csamul_rca16_and12_4 ^ s_csamul_rca16_fa13_3_xor1;
  assign s_csamul_rca16_fa12_4_and0 = s_csamul_rca16_and12_4 & s_csamul_rca16_fa13_3_xor1;
  assign s_csamul_rca16_fa12_4_xor1 = s_csamul_rca16_fa12_4_xor0 ^ s_csamul_rca16_fa12_3_or0;
  assign s_csamul_rca16_fa12_4_and1 = s_csamul_rca16_fa12_4_xor0 & s_csamul_rca16_fa12_3_or0;
  assign s_csamul_rca16_fa12_4_or0 = s_csamul_rca16_fa12_4_and0 | s_csamul_rca16_fa12_4_and1;
  assign s_csamul_rca16_and13_4 = a[13] & b[4];
  assign s_csamul_rca16_fa13_4_xor0 = s_csamul_rca16_and13_4 ^ s_csamul_rca16_fa14_3_xor1;
  assign s_csamul_rca16_fa13_4_and0 = s_csamul_rca16_and13_4 & s_csamul_rca16_fa14_3_xor1;
  assign s_csamul_rca16_fa13_4_xor1 = s_csamul_rca16_fa13_4_xor0 ^ s_csamul_rca16_fa13_3_or0;
  assign s_csamul_rca16_fa13_4_and1 = s_csamul_rca16_fa13_4_xor0 & s_csamul_rca16_fa13_3_or0;
  assign s_csamul_rca16_fa13_4_or0 = s_csamul_rca16_fa13_4_and0 | s_csamul_rca16_fa13_4_and1;
  assign s_csamul_rca16_and14_4 = a[14] & b[4];
  assign s_csamul_rca16_fa14_4_xor0 = s_csamul_rca16_and14_4 ^ s_csamul_rca16_ha15_3_xor0;
  assign s_csamul_rca16_fa14_4_and0 = s_csamul_rca16_and14_4 & s_csamul_rca16_ha15_3_xor0;
  assign s_csamul_rca16_fa14_4_xor1 = s_csamul_rca16_fa14_4_xor0 ^ s_csamul_rca16_fa14_3_or0;
  assign s_csamul_rca16_fa14_4_and1 = s_csamul_rca16_fa14_4_xor0 & s_csamul_rca16_fa14_3_or0;
  assign s_csamul_rca16_fa14_4_or0 = s_csamul_rca16_fa14_4_and0 | s_csamul_rca16_fa14_4_and1;
  assign s_csamul_rca16_nand15_4 = ~(a[15] & b[4]);
  assign s_csamul_rca16_ha15_4_xor0 = s_csamul_rca16_nand15_4 ^ s_csamul_rca16_ha15_3_and0;
  assign s_csamul_rca16_ha15_4_and0 = s_csamul_rca16_nand15_4 & s_csamul_rca16_ha15_3_and0;
  assign s_csamul_rca16_and0_5 = a[0] & b[5];
  assign s_csamul_rca16_fa0_5_xor0 = s_csamul_rca16_and0_5 ^ s_csamul_rca16_fa1_4_xor1;
  assign s_csamul_rca16_fa0_5_and0 = s_csamul_rca16_and0_5 & s_csamul_rca16_fa1_4_xor1;
  assign s_csamul_rca16_fa0_5_xor1 = s_csamul_rca16_fa0_5_xor0 ^ s_csamul_rca16_fa0_4_or0;
  assign s_csamul_rca16_fa0_5_and1 = s_csamul_rca16_fa0_5_xor0 & s_csamul_rca16_fa0_4_or0;
  assign s_csamul_rca16_fa0_5_or0 = s_csamul_rca16_fa0_5_and0 | s_csamul_rca16_fa0_5_and1;
  assign s_csamul_rca16_and1_5 = a[1] & b[5];
  assign s_csamul_rca16_fa1_5_xor0 = s_csamul_rca16_and1_5 ^ s_csamul_rca16_fa2_4_xor1;
  assign s_csamul_rca16_fa1_5_and0 = s_csamul_rca16_and1_5 & s_csamul_rca16_fa2_4_xor1;
  assign s_csamul_rca16_fa1_5_xor1 = s_csamul_rca16_fa1_5_xor0 ^ s_csamul_rca16_fa1_4_or0;
  assign s_csamul_rca16_fa1_5_and1 = s_csamul_rca16_fa1_5_xor0 & s_csamul_rca16_fa1_4_or0;
  assign s_csamul_rca16_fa1_5_or0 = s_csamul_rca16_fa1_5_and0 | s_csamul_rca16_fa1_5_and1;
  assign s_csamul_rca16_and2_5 = a[2] & b[5];
  assign s_csamul_rca16_fa2_5_xor0 = s_csamul_rca16_and2_5 ^ s_csamul_rca16_fa3_4_xor1;
  assign s_csamul_rca16_fa2_5_and0 = s_csamul_rca16_and2_5 & s_csamul_rca16_fa3_4_xor1;
  assign s_csamul_rca16_fa2_5_xor1 = s_csamul_rca16_fa2_5_xor0 ^ s_csamul_rca16_fa2_4_or0;
  assign s_csamul_rca16_fa2_5_and1 = s_csamul_rca16_fa2_5_xor0 & s_csamul_rca16_fa2_4_or0;
  assign s_csamul_rca16_fa2_5_or0 = s_csamul_rca16_fa2_5_and0 | s_csamul_rca16_fa2_5_and1;
  assign s_csamul_rca16_and3_5 = a[3] & b[5];
  assign s_csamul_rca16_fa3_5_xor0 = s_csamul_rca16_and3_5 ^ s_csamul_rca16_fa4_4_xor1;
  assign s_csamul_rca16_fa3_5_and0 = s_csamul_rca16_and3_5 & s_csamul_rca16_fa4_4_xor1;
  assign s_csamul_rca16_fa3_5_xor1 = s_csamul_rca16_fa3_5_xor0 ^ s_csamul_rca16_fa3_4_or0;
  assign s_csamul_rca16_fa3_5_and1 = s_csamul_rca16_fa3_5_xor0 & s_csamul_rca16_fa3_4_or0;
  assign s_csamul_rca16_fa3_5_or0 = s_csamul_rca16_fa3_5_and0 | s_csamul_rca16_fa3_5_and1;
  assign s_csamul_rca16_and4_5 = a[4] & b[5];
  assign s_csamul_rca16_fa4_5_xor0 = s_csamul_rca16_and4_5 ^ s_csamul_rca16_fa5_4_xor1;
  assign s_csamul_rca16_fa4_5_and0 = s_csamul_rca16_and4_5 & s_csamul_rca16_fa5_4_xor1;
  assign s_csamul_rca16_fa4_5_xor1 = s_csamul_rca16_fa4_5_xor0 ^ s_csamul_rca16_fa4_4_or0;
  assign s_csamul_rca16_fa4_5_and1 = s_csamul_rca16_fa4_5_xor0 & s_csamul_rca16_fa4_4_or0;
  assign s_csamul_rca16_fa4_5_or0 = s_csamul_rca16_fa4_5_and0 | s_csamul_rca16_fa4_5_and1;
  assign s_csamul_rca16_and5_5 = a[5] & b[5];
  assign s_csamul_rca16_fa5_5_xor0 = s_csamul_rca16_and5_5 ^ s_csamul_rca16_fa6_4_xor1;
  assign s_csamul_rca16_fa5_5_and0 = s_csamul_rca16_and5_5 & s_csamul_rca16_fa6_4_xor1;
  assign s_csamul_rca16_fa5_5_xor1 = s_csamul_rca16_fa5_5_xor0 ^ s_csamul_rca16_fa5_4_or0;
  assign s_csamul_rca16_fa5_5_and1 = s_csamul_rca16_fa5_5_xor0 & s_csamul_rca16_fa5_4_or0;
  assign s_csamul_rca16_fa5_5_or0 = s_csamul_rca16_fa5_5_and0 | s_csamul_rca16_fa5_5_and1;
  assign s_csamul_rca16_and6_5 = a[6] & b[5];
  assign s_csamul_rca16_fa6_5_xor0 = s_csamul_rca16_and6_5 ^ s_csamul_rca16_fa7_4_xor1;
  assign s_csamul_rca16_fa6_5_and0 = s_csamul_rca16_and6_5 & s_csamul_rca16_fa7_4_xor1;
  assign s_csamul_rca16_fa6_5_xor1 = s_csamul_rca16_fa6_5_xor0 ^ s_csamul_rca16_fa6_4_or0;
  assign s_csamul_rca16_fa6_5_and1 = s_csamul_rca16_fa6_5_xor0 & s_csamul_rca16_fa6_4_or0;
  assign s_csamul_rca16_fa6_5_or0 = s_csamul_rca16_fa6_5_and0 | s_csamul_rca16_fa6_5_and1;
  assign s_csamul_rca16_and7_5 = a[7] & b[5];
  assign s_csamul_rca16_fa7_5_xor0 = s_csamul_rca16_and7_5 ^ s_csamul_rca16_fa8_4_xor1;
  assign s_csamul_rca16_fa7_5_and0 = s_csamul_rca16_and7_5 & s_csamul_rca16_fa8_4_xor1;
  assign s_csamul_rca16_fa7_5_xor1 = s_csamul_rca16_fa7_5_xor0 ^ s_csamul_rca16_fa7_4_or0;
  assign s_csamul_rca16_fa7_5_and1 = s_csamul_rca16_fa7_5_xor0 & s_csamul_rca16_fa7_4_or0;
  assign s_csamul_rca16_fa7_5_or0 = s_csamul_rca16_fa7_5_and0 | s_csamul_rca16_fa7_5_and1;
  assign s_csamul_rca16_and8_5 = a[8] & b[5];
  assign s_csamul_rca16_fa8_5_xor0 = s_csamul_rca16_and8_5 ^ s_csamul_rca16_fa9_4_xor1;
  assign s_csamul_rca16_fa8_5_and0 = s_csamul_rca16_and8_5 & s_csamul_rca16_fa9_4_xor1;
  assign s_csamul_rca16_fa8_5_xor1 = s_csamul_rca16_fa8_5_xor0 ^ s_csamul_rca16_fa8_4_or0;
  assign s_csamul_rca16_fa8_5_and1 = s_csamul_rca16_fa8_5_xor0 & s_csamul_rca16_fa8_4_or0;
  assign s_csamul_rca16_fa8_5_or0 = s_csamul_rca16_fa8_5_and0 | s_csamul_rca16_fa8_5_and1;
  assign s_csamul_rca16_and9_5 = a[9] & b[5];
  assign s_csamul_rca16_fa9_5_xor0 = s_csamul_rca16_and9_5 ^ s_csamul_rca16_fa10_4_xor1;
  assign s_csamul_rca16_fa9_5_and0 = s_csamul_rca16_and9_5 & s_csamul_rca16_fa10_4_xor1;
  assign s_csamul_rca16_fa9_5_xor1 = s_csamul_rca16_fa9_5_xor0 ^ s_csamul_rca16_fa9_4_or0;
  assign s_csamul_rca16_fa9_5_and1 = s_csamul_rca16_fa9_5_xor0 & s_csamul_rca16_fa9_4_or0;
  assign s_csamul_rca16_fa9_5_or0 = s_csamul_rca16_fa9_5_and0 | s_csamul_rca16_fa9_5_and1;
  assign s_csamul_rca16_and10_5 = a[10] & b[5];
  assign s_csamul_rca16_fa10_5_xor0 = s_csamul_rca16_and10_5 ^ s_csamul_rca16_fa11_4_xor1;
  assign s_csamul_rca16_fa10_5_and0 = s_csamul_rca16_and10_5 & s_csamul_rca16_fa11_4_xor1;
  assign s_csamul_rca16_fa10_5_xor1 = s_csamul_rca16_fa10_5_xor0 ^ s_csamul_rca16_fa10_4_or0;
  assign s_csamul_rca16_fa10_5_and1 = s_csamul_rca16_fa10_5_xor0 & s_csamul_rca16_fa10_4_or0;
  assign s_csamul_rca16_fa10_5_or0 = s_csamul_rca16_fa10_5_and0 | s_csamul_rca16_fa10_5_and1;
  assign s_csamul_rca16_and11_5 = a[11] & b[5];
  assign s_csamul_rca16_fa11_5_xor0 = s_csamul_rca16_and11_5 ^ s_csamul_rca16_fa12_4_xor1;
  assign s_csamul_rca16_fa11_5_and0 = s_csamul_rca16_and11_5 & s_csamul_rca16_fa12_4_xor1;
  assign s_csamul_rca16_fa11_5_xor1 = s_csamul_rca16_fa11_5_xor0 ^ s_csamul_rca16_fa11_4_or0;
  assign s_csamul_rca16_fa11_5_and1 = s_csamul_rca16_fa11_5_xor0 & s_csamul_rca16_fa11_4_or0;
  assign s_csamul_rca16_fa11_5_or0 = s_csamul_rca16_fa11_5_and0 | s_csamul_rca16_fa11_5_and1;
  assign s_csamul_rca16_and12_5 = a[12] & b[5];
  assign s_csamul_rca16_fa12_5_xor0 = s_csamul_rca16_and12_5 ^ s_csamul_rca16_fa13_4_xor1;
  assign s_csamul_rca16_fa12_5_and0 = s_csamul_rca16_and12_5 & s_csamul_rca16_fa13_4_xor1;
  assign s_csamul_rca16_fa12_5_xor1 = s_csamul_rca16_fa12_5_xor0 ^ s_csamul_rca16_fa12_4_or0;
  assign s_csamul_rca16_fa12_5_and1 = s_csamul_rca16_fa12_5_xor0 & s_csamul_rca16_fa12_4_or0;
  assign s_csamul_rca16_fa12_5_or0 = s_csamul_rca16_fa12_5_and0 | s_csamul_rca16_fa12_5_and1;
  assign s_csamul_rca16_and13_5 = a[13] & b[5];
  assign s_csamul_rca16_fa13_5_xor0 = s_csamul_rca16_and13_5 ^ s_csamul_rca16_fa14_4_xor1;
  assign s_csamul_rca16_fa13_5_and0 = s_csamul_rca16_and13_5 & s_csamul_rca16_fa14_4_xor1;
  assign s_csamul_rca16_fa13_5_xor1 = s_csamul_rca16_fa13_5_xor0 ^ s_csamul_rca16_fa13_4_or0;
  assign s_csamul_rca16_fa13_5_and1 = s_csamul_rca16_fa13_5_xor0 & s_csamul_rca16_fa13_4_or0;
  assign s_csamul_rca16_fa13_5_or0 = s_csamul_rca16_fa13_5_and0 | s_csamul_rca16_fa13_5_and1;
  assign s_csamul_rca16_and14_5 = a[14] & b[5];
  assign s_csamul_rca16_fa14_5_xor0 = s_csamul_rca16_and14_5 ^ s_csamul_rca16_ha15_4_xor0;
  assign s_csamul_rca16_fa14_5_and0 = s_csamul_rca16_and14_5 & s_csamul_rca16_ha15_4_xor0;
  assign s_csamul_rca16_fa14_5_xor1 = s_csamul_rca16_fa14_5_xor0 ^ s_csamul_rca16_fa14_4_or0;
  assign s_csamul_rca16_fa14_5_and1 = s_csamul_rca16_fa14_5_xor0 & s_csamul_rca16_fa14_4_or0;
  assign s_csamul_rca16_fa14_5_or0 = s_csamul_rca16_fa14_5_and0 | s_csamul_rca16_fa14_5_and1;
  assign s_csamul_rca16_nand15_5 = ~(a[15] & b[5]);
  assign s_csamul_rca16_ha15_5_xor0 = s_csamul_rca16_nand15_5 ^ s_csamul_rca16_ha15_4_and0;
  assign s_csamul_rca16_ha15_5_and0 = s_csamul_rca16_nand15_5 & s_csamul_rca16_ha15_4_and0;
  assign s_csamul_rca16_and0_6 = a[0] & b[6];
  assign s_csamul_rca16_fa0_6_xor0 = s_csamul_rca16_and0_6 ^ s_csamul_rca16_fa1_5_xor1;
  assign s_csamul_rca16_fa0_6_and0 = s_csamul_rca16_and0_6 & s_csamul_rca16_fa1_5_xor1;
  assign s_csamul_rca16_fa0_6_xor1 = s_csamul_rca16_fa0_6_xor0 ^ s_csamul_rca16_fa0_5_or0;
  assign s_csamul_rca16_fa0_6_and1 = s_csamul_rca16_fa0_6_xor0 & s_csamul_rca16_fa0_5_or0;
  assign s_csamul_rca16_fa0_6_or0 = s_csamul_rca16_fa0_6_and0 | s_csamul_rca16_fa0_6_and1;
  assign s_csamul_rca16_and1_6 = a[1] & b[6];
  assign s_csamul_rca16_fa1_6_xor0 = s_csamul_rca16_and1_6 ^ s_csamul_rca16_fa2_5_xor1;
  assign s_csamul_rca16_fa1_6_and0 = s_csamul_rca16_and1_6 & s_csamul_rca16_fa2_5_xor1;
  assign s_csamul_rca16_fa1_6_xor1 = s_csamul_rca16_fa1_6_xor0 ^ s_csamul_rca16_fa1_5_or0;
  assign s_csamul_rca16_fa1_6_and1 = s_csamul_rca16_fa1_6_xor0 & s_csamul_rca16_fa1_5_or0;
  assign s_csamul_rca16_fa1_6_or0 = s_csamul_rca16_fa1_6_and0 | s_csamul_rca16_fa1_6_and1;
  assign s_csamul_rca16_and2_6 = a[2] & b[6];
  assign s_csamul_rca16_fa2_6_xor0 = s_csamul_rca16_and2_6 ^ s_csamul_rca16_fa3_5_xor1;
  assign s_csamul_rca16_fa2_6_and0 = s_csamul_rca16_and2_6 & s_csamul_rca16_fa3_5_xor1;
  assign s_csamul_rca16_fa2_6_xor1 = s_csamul_rca16_fa2_6_xor0 ^ s_csamul_rca16_fa2_5_or0;
  assign s_csamul_rca16_fa2_6_and1 = s_csamul_rca16_fa2_6_xor0 & s_csamul_rca16_fa2_5_or0;
  assign s_csamul_rca16_fa2_6_or0 = s_csamul_rca16_fa2_6_and0 | s_csamul_rca16_fa2_6_and1;
  assign s_csamul_rca16_and3_6 = a[3] & b[6];
  assign s_csamul_rca16_fa3_6_xor0 = s_csamul_rca16_and3_6 ^ s_csamul_rca16_fa4_5_xor1;
  assign s_csamul_rca16_fa3_6_and0 = s_csamul_rca16_and3_6 & s_csamul_rca16_fa4_5_xor1;
  assign s_csamul_rca16_fa3_6_xor1 = s_csamul_rca16_fa3_6_xor0 ^ s_csamul_rca16_fa3_5_or0;
  assign s_csamul_rca16_fa3_6_and1 = s_csamul_rca16_fa3_6_xor0 & s_csamul_rca16_fa3_5_or0;
  assign s_csamul_rca16_fa3_6_or0 = s_csamul_rca16_fa3_6_and0 | s_csamul_rca16_fa3_6_and1;
  assign s_csamul_rca16_and4_6 = a[4] & b[6];
  assign s_csamul_rca16_fa4_6_xor0 = s_csamul_rca16_and4_6 ^ s_csamul_rca16_fa5_5_xor1;
  assign s_csamul_rca16_fa4_6_and0 = s_csamul_rca16_and4_6 & s_csamul_rca16_fa5_5_xor1;
  assign s_csamul_rca16_fa4_6_xor1 = s_csamul_rca16_fa4_6_xor0 ^ s_csamul_rca16_fa4_5_or0;
  assign s_csamul_rca16_fa4_6_and1 = s_csamul_rca16_fa4_6_xor0 & s_csamul_rca16_fa4_5_or0;
  assign s_csamul_rca16_fa4_6_or0 = s_csamul_rca16_fa4_6_and0 | s_csamul_rca16_fa4_6_and1;
  assign s_csamul_rca16_and5_6 = a[5] & b[6];
  assign s_csamul_rca16_fa5_6_xor0 = s_csamul_rca16_and5_6 ^ s_csamul_rca16_fa6_5_xor1;
  assign s_csamul_rca16_fa5_6_and0 = s_csamul_rca16_and5_6 & s_csamul_rca16_fa6_5_xor1;
  assign s_csamul_rca16_fa5_6_xor1 = s_csamul_rca16_fa5_6_xor0 ^ s_csamul_rca16_fa5_5_or0;
  assign s_csamul_rca16_fa5_6_and1 = s_csamul_rca16_fa5_6_xor0 & s_csamul_rca16_fa5_5_or0;
  assign s_csamul_rca16_fa5_6_or0 = s_csamul_rca16_fa5_6_and0 | s_csamul_rca16_fa5_6_and1;
  assign s_csamul_rca16_and6_6 = a[6] & b[6];
  assign s_csamul_rca16_fa6_6_xor0 = s_csamul_rca16_and6_6 ^ s_csamul_rca16_fa7_5_xor1;
  assign s_csamul_rca16_fa6_6_and0 = s_csamul_rca16_and6_6 & s_csamul_rca16_fa7_5_xor1;
  assign s_csamul_rca16_fa6_6_xor1 = s_csamul_rca16_fa6_6_xor0 ^ s_csamul_rca16_fa6_5_or0;
  assign s_csamul_rca16_fa6_6_and1 = s_csamul_rca16_fa6_6_xor0 & s_csamul_rca16_fa6_5_or0;
  assign s_csamul_rca16_fa6_6_or0 = s_csamul_rca16_fa6_6_and0 | s_csamul_rca16_fa6_6_and1;
  assign s_csamul_rca16_and7_6 = a[7] & b[6];
  assign s_csamul_rca16_fa7_6_xor0 = s_csamul_rca16_and7_6 ^ s_csamul_rca16_fa8_5_xor1;
  assign s_csamul_rca16_fa7_6_and0 = s_csamul_rca16_and7_6 & s_csamul_rca16_fa8_5_xor1;
  assign s_csamul_rca16_fa7_6_xor1 = s_csamul_rca16_fa7_6_xor0 ^ s_csamul_rca16_fa7_5_or0;
  assign s_csamul_rca16_fa7_6_and1 = s_csamul_rca16_fa7_6_xor0 & s_csamul_rca16_fa7_5_or0;
  assign s_csamul_rca16_fa7_6_or0 = s_csamul_rca16_fa7_6_and0 | s_csamul_rca16_fa7_6_and1;
  assign s_csamul_rca16_and8_6 = a[8] & b[6];
  assign s_csamul_rca16_fa8_6_xor0 = s_csamul_rca16_and8_6 ^ s_csamul_rca16_fa9_5_xor1;
  assign s_csamul_rca16_fa8_6_and0 = s_csamul_rca16_and8_6 & s_csamul_rca16_fa9_5_xor1;
  assign s_csamul_rca16_fa8_6_xor1 = s_csamul_rca16_fa8_6_xor0 ^ s_csamul_rca16_fa8_5_or0;
  assign s_csamul_rca16_fa8_6_and1 = s_csamul_rca16_fa8_6_xor0 & s_csamul_rca16_fa8_5_or0;
  assign s_csamul_rca16_fa8_6_or0 = s_csamul_rca16_fa8_6_and0 | s_csamul_rca16_fa8_6_and1;
  assign s_csamul_rca16_and9_6 = a[9] & b[6];
  assign s_csamul_rca16_fa9_6_xor0 = s_csamul_rca16_and9_6 ^ s_csamul_rca16_fa10_5_xor1;
  assign s_csamul_rca16_fa9_6_and0 = s_csamul_rca16_and9_6 & s_csamul_rca16_fa10_5_xor1;
  assign s_csamul_rca16_fa9_6_xor1 = s_csamul_rca16_fa9_6_xor0 ^ s_csamul_rca16_fa9_5_or0;
  assign s_csamul_rca16_fa9_6_and1 = s_csamul_rca16_fa9_6_xor0 & s_csamul_rca16_fa9_5_or0;
  assign s_csamul_rca16_fa9_6_or0 = s_csamul_rca16_fa9_6_and0 | s_csamul_rca16_fa9_6_and1;
  assign s_csamul_rca16_and10_6 = a[10] & b[6];
  assign s_csamul_rca16_fa10_6_xor0 = s_csamul_rca16_and10_6 ^ s_csamul_rca16_fa11_5_xor1;
  assign s_csamul_rca16_fa10_6_and0 = s_csamul_rca16_and10_6 & s_csamul_rca16_fa11_5_xor1;
  assign s_csamul_rca16_fa10_6_xor1 = s_csamul_rca16_fa10_6_xor0 ^ s_csamul_rca16_fa10_5_or0;
  assign s_csamul_rca16_fa10_6_and1 = s_csamul_rca16_fa10_6_xor0 & s_csamul_rca16_fa10_5_or0;
  assign s_csamul_rca16_fa10_6_or0 = s_csamul_rca16_fa10_6_and0 | s_csamul_rca16_fa10_6_and1;
  assign s_csamul_rca16_and11_6 = a[11] & b[6];
  assign s_csamul_rca16_fa11_6_xor0 = s_csamul_rca16_and11_6 ^ s_csamul_rca16_fa12_5_xor1;
  assign s_csamul_rca16_fa11_6_and0 = s_csamul_rca16_and11_6 & s_csamul_rca16_fa12_5_xor1;
  assign s_csamul_rca16_fa11_6_xor1 = s_csamul_rca16_fa11_6_xor0 ^ s_csamul_rca16_fa11_5_or0;
  assign s_csamul_rca16_fa11_6_and1 = s_csamul_rca16_fa11_6_xor0 & s_csamul_rca16_fa11_5_or0;
  assign s_csamul_rca16_fa11_6_or0 = s_csamul_rca16_fa11_6_and0 | s_csamul_rca16_fa11_6_and1;
  assign s_csamul_rca16_and12_6 = a[12] & b[6];
  assign s_csamul_rca16_fa12_6_xor0 = s_csamul_rca16_and12_6 ^ s_csamul_rca16_fa13_5_xor1;
  assign s_csamul_rca16_fa12_6_and0 = s_csamul_rca16_and12_6 & s_csamul_rca16_fa13_5_xor1;
  assign s_csamul_rca16_fa12_6_xor1 = s_csamul_rca16_fa12_6_xor0 ^ s_csamul_rca16_fa12_5_or0;
  assign s_csamul_rca16_fa12_6_and1 = s_csamul_rca16_fa12_6_xor0 & s_csamul_rca16_fa12_5_or0;
  assign s_csamul_rca16_fa12_6_or0 = s_csamul_rca16_fa12_6_and0 | s_csamul_rca16_fa12_6_and1;
  assign s_csamul_rca16_and13_6 = a[13] & b[6];
  assign s_csamul_rca16_fa13_6_xor0 = s_csamul_rca16_and13_6 ^ s_csamul_rca16_fa14_5_xor1;
  assign s_csamul_rca16_fa13_6_and0 = s_csamul_rca16_and13_6 & s_csamul_rca16_fa14_5_xor1;
  assign s_csamul_rca16_fa13_6_xor1 = s_csamul_rca16_fa13_6_xor0 ^ s_csamul_rca16_fa13_5_or0;
  assign s_csamul_rca16_fa13_6_and1 = s_csamul_rca16_fa13_6_xor0 & s_csamul_rca16_fa13_5_or0;
  assign s_csamul_rca16_fa13_6_or0 = s_csamul_rca16_fa13_6_and0 | s_csamul_rca16_fa13_6_and1;
  assign s_csamul_rca16_and14_6 = a[14] & b[6];
  assign s_csamul_rca16_fa14_6_xor0 = s_csamul_rca16_and14_6 ^ s_csamul_rca16_ha15_5_xor0;
  assign s_csamul_rca16_fa14_6_and0 = s_csamul_rca16_and14_6 & s_csamul_rca16_ha15_5_xor0;
  assign s_csamul_rca16_fa14_6_xor1 = s_csamul_rca16_fa14_6_xor0 ^ s_csamul_rca16_fa14_5_or0;
  assign s_csamul_rca16_fa14_6_and1 = s_csamul_rca16_fa14_6_xor0 & s_csamul_rca16_fa14_5_or0;
  assign s_csamul_rca16_fa14_6_or0 = s_csamul_rca16_fa14_6_and0 | s_csamul_rca16_fa14_6_and1;
  assign s_csamul_rca16_nand15_6 = ~(a[15] & b[6]);
  assign s_csamul_rca16_ha15_6_xor0 = s_csamul_rca16_nand15_6 ^ s_csamul_rca16_ha15_5_and0;
  assign s_csamul_rca16_ha15_6_and0 = s_csamul_rca16_nand15_6 & s_csamul_rca16_ha15_5_and0;
  assign s_csamul_rca16_and0_7 = a[0] & b[7];
  assign s_csamul_rca16_fa0_7_xor0 = s_csamul_rca16_and0_7 ^ s_csamul_rca16_fa1_6_xor1;
  assign s_csamul_rca16_fa0_7_and0 = s_csamul_rca16_and0_7 & s_csamul_rca16_fa1_6_xor1;
  assign s_csamul_rca16_fa0_7_xor1 = s_csamul_rca16_fa0_7_xor0 ^ s_csamul_rca16_fa0_6_or0;
  assign s_csamul_rca16_fa0_7_and1 = s_csamul_rca16_fa0_7_xor0 & s_csamul_rca16_fa0_6_or0;
  assign s_csamul_rca16_fa0_7_or0 = s_csamul_rca16_fa0_7_and0 | s_csamul_rca16_fa0_7_and1;
  assign s_csamul_rca16_and1_7 = a[1] & b[7];
  assign s_csamul_rca16_fa1_7_xor0 = s_csamul_rca16_and1_7 ^ s_csamul_rca16_fa2_6_xor1;
  assign s_csamul_rca16_fa1_7_and0 = s_csamul_rca16_and1_7 & s_csamul_rca16_fa2_6_xor1;
  assign s_csamul_rca16_fa1_7_xor1 = s_csamul_rca16_fa1_7_xor0 ^ s_csamul_rca16_fa1_6_or0;
  assign s_csamul_rca16_fa1_7_and1 = s_csamul_rca16_fa1_7_xor0 & s_csamul_rca16_fa1_6_or0;
  assign s_csamul_rca16_fa1_7_or0 = s_csamul_rca16_fa1_7_and0 | s_csamul_rca16_fa1_7_and1;
  assign s_csamul_rca16_and2_7 = a[2] & b[7];
  assign s_csamul_rca16_fa2_7_xor0 = s_csamul_rca16_and2_7 ^ s_csamul_rca16_fa3_6_xor1;
  assign s_csamul_rca16_fa2_7_and0 = s_csamul_rca16_and2_7 & s_csamul_rca16_fa3_6_xor1;
  assign s_csamul_rca16_fa2_7_xor1 = s_csamul_rca16_fa2_7_xor0 ^ s_csamul_rca16_fa2_6_or0;
  assign s_csamul_rca16_fa2_7_and1 = s_csamul_rca16_fa2_7_xor0 & s_csamul_rca16_fa2_6_or0;
  assign s_csamul_rca16_fa2_7_or0 = s_csamul_rca16_fa2_7_and0 | s_csamul_rca16_fa2_7_and1;
  assign s_csamul_rca16_and3_7 = a[3] & b[7];
  assign s_csamul_rca16_fa3_7_xor0 = s_csamul_rca16_and3_7 ^ s_csamul_rca16_fa4_6_xor1;
  assign s_csamul_rca16_fa3_7_and0 = s_csamul_rca16_and3_7 & s_csamul_rca16_fa4_6_xor1;
  assign s_csamul_rca16_fa3_7_xor1 = s_csamul_rca16_fa3_7_xor0 ^ s_csamul_rca16_fa3_6_or0;
  assign s_csamul_rca16_fa3_7_and1 = s_csamul_rca16_fa3_7_xor0 & s_csamul_rca16_fa3_6_or0;
  assign s_csamul_rca16_fa3_7_or0 = s_csamul_rca16_fa3_7_and0 | s_csamul_rca16_fa3_7_and1;
  assign s_csamul_rca16_and4_7 = a[4] & b[7];
  assign s_csamul_rca16_fa4_7_xor0 = s_csamul_rca16_and4_7 ^ s_csamul_rca16_fa5_6_xor1;
  assign s_csamul_rca16_fa4_7_and0 = s_csamul_rca16_and4_7 & s_csamul_rca16_fa5_6_xor1;
  assign s_csamul_rca16_fa4_7_xor1 = s_csamul_rca16_fa4_7_xor0 ^ s_csamul_rca16_fa4_6_or0;
  assign s_csamul_rca16_fa4_7_and1 = s_csamul_rca16_fa4_7_xor0 & s_csamul_rca16_fa4_6_or0;
  assign s_csamul_rca16_fa4_7_or0 = s_csamul_rca16_fa4_7_and0 | s_csamul_rca16_fa4_7_and1;
  assign s_csamul_rca16_and5_7 = a[5] & b[7];
  assign s_csamul_rca16_fa5_7_xor0 = s_csamul_rca16_and5_7 ^ s_csamul_rca16_fa6_6_xor1;
  assign s_csamul_rca16_fa5_7_and0 = s_csamul_rca16_and5_7 & s_csamul_rca16_fa6_6_xor1;
  assign s_csamul_rca16_fa5_7_xor1 = s_csamul_rca16_fa5_7_xor0 ^ s_csamul_rca16_fa5_6_or0;
  assign s_csamul_rca16_fa5_7_and1 = s_csamul_rca16_fa5_7_xor0 & s_csamul_rca16_fa5_6_or0;
  assign s_csamul_rca16_fa5_7_or0 = s_csamul_rca16_fa5_7_and0 | s_csamul_rca16_fa5_7_and1;
  assign s_csamul_rca16_and6_7 = a[6] & b[7];
  assign s_csamul_rca16_fa6_7_xor0 = s_csamul_rca16_and6_7 ^ s_csamul_rca16_fa7_6_xor1;
  assign s_csamul_rca16_fa6_7_and0 = s_csamul_rca16_and6_7 & s_csamul_rca16_fa7_6_xor1;
  assign s_csamul_rca16_fa6_7_xor1 = s_csamul_rca16_fa6_7_xor0 ^ s_csamul_rca16_fa6_6_or0;
  assign s_csamul_rca16_fa6_7_and1 = s_csamul_rca16_fa6_7_xor0 & s_csamul_rca16_fa6_6_or0;
  assign s_csamul_rca16_fa6_7_or0 = s_csamul_rca16_fa6_7_and0 | s_csamul_rca16_fa6_7_and1;
  assign s_csamul_rca16_and7_7 = a[7] & b[7];
  assign s_csamul_rca16_fa7_7_xor0 = s_csamul_rca16_and7_7 ^ s_csamul_rca16_fa8_6_xor1;
  assign s_csamul_rca16_fa7_7_and0 = s_csamul_rca16_and7_7 & s_csamul_rca16_fa8_6_xor1;
  assign s_csamul_rca16_fa7_7_xor1 = s_csamul_rca16_fa7_7_xor0 ^ s_csamul_rca16_fa7_6_or0;
  assign s_csamul_rca16_fa7_7_and1 = s_csamul_rca16_fa7_7_xor0 & s_csamul_rca16_fa7_6_or0;
  assign s_csamul_rca16_fa7_7_or0 = s_csamul_rca16_fa7_7_and0 | s_csamul_rca16_fa7_7_and1;
  assign s_csamul_rca16_and8_7 = a[8] & b[7];
  assign s_csamul_rca16_fa8_7_xor0 = s_csamul_rca16_and8_7 ^ s_csamul_rca16_fa9_6_xor1;
  assign s_csamul_rca16_fa8_7_and0 = s_csamul_rca16_and8_7 & s_csamul_rca16_fa9_6_xor1;
  assign s_csamul_rca16_fa8_7_xor1 = s_csamul_rca16_fa8_7_xor0 ^ s_csamul_rca16_fa8_6_or0;
  assign s_csamul_rca16_fa8_7_and1 = s_csamul_rca16_fa8_7_xor0 & s_csamul_rca16_fa8_6_or0;
  assign s_csamul_rca16_fa8_7_or0 = s_csamul_rca16_fa8_7_and0 | s_csamul_rca16_fa8_7_and1;
  assign s_csamul_rca16_and9_7 = a[9] & b[7];
  assign s_csamul_rca16_fa9_7_xor0 = s_csamul_rca16_and9_7 ^ s_csamul_rca16_fa10_6_xor1;
  assign s_csamul_rca16_fa9_7_and0 = s_csamul_rca16_and9_7 & s_csamul_rca16_fa10_6_xor1;
  assign s_csamul_rca16_fa9_7_xor1 = s_csamul_rca16_fa9_7_xor0 ^ s_csamul_rca16_fa9_6_or0;
  assign s_csamul_rca16_fa9_7_and1 = s_csamul_rca16_fa9_7_xor0 & s_csamul_rca16_fa9_6_or0;
  assign s_csamul_rca16_fa9_7_or0 = s_csamul_rca16_fa9_7_and0 | s_csamul_rca16_fa9_7_and1;
  assign s_csamul_rca16_and10_7 = a[10] & b[7];
  assign s_csamul_rca16_fa10_7_xor0 = s_csamul_rca16_and10_7 ^ s_csamul_rca16_fa11_6_xor1;
  assign s_csamul_rca16_fa10_7_and0 = s_csamul_rca16_and10_7 & s_csamul_rca16_fa11_6_xor1;
  assign s_csamul_rca16_fa10_7_xor1 = s_csamul_rca16_fa10_7_xor0 ^ s_csamul_rca16_fa10_6_or0;
  assign s_csamul_rca16_fa10_7_and1 = s_csamul_rca16_fa10_7_xor0 & s_csamul_rca16_fa10_6_or0;
  assign s_csamul_rca16_fa10_7_or0 = s_csamul_rca16_fa10_7_and0 | s_csamul_rca16_fa10_7_and1;
  assign s_csamul_rca16_and11_7 = a[11] & b[7];
  assign s_csamul_rca16_fa11_7_xor0 = s_csamul_rca16_and11_7 ^ s_csamul_rca16_fa12_6_xor1;
  assign s_csamul_rca16_fa11_7_and0 = s_csamul_rca16_and11_7 & s_csamul_rca16_fa12_6_xor1;
  assign s_csamul_rca16_fa11_7_xor1 = s_csamul_rca16_fa11_7_xor0 ^ s_csamul_rca16_fa11_6_or0;
  assign s_csamul_rca16_fa11_7_and1 = s_csamul_rca16_fa11_7_xor0 & s_csamul_rca16_fa11_6_or0;
  assign s_csamul_rca16_fa11_7_or0 = s_csamul_rca16_fa11_7_and0 | s_csamul_rca16_fa11_7_and1;
  assign s_csamul_rca16_and12_7 = a[12] & b[7];
  assign s_csamul_rca16_fa12_7_xor0 = s_csamul_rca16_and12_7 ^ s_csamul_rca16_fa13_6_xor1;
  assign s_csamul_rca16_fa12_7_and0 = s_csamul_rca16_and12_7 & s_csamul_rca16_fa13_6_xor1;
  assign s_csamul_rca16_fa12_7_xor1 = s_csamul_rca16_fa12_7_xor0 ^ s_csamul_rca16_fa12_6_or0;
  assign s_csamul_rca16_fa12_7_and1 = s_csamul_rca16_fa12_7_xor0 & s_csamul_rca16_fa12_6_or0;
  assign s_csamul_rca16_fa12_7_or0 = s_csamul_rca16_fa12_7_and0 | s_csamul_rca16_fa12_7_and1;
  assign s_csamul_rca16_and13_7 = a[13] & b[7];
  assign s_csamul_rca16_fa13_7_xor0 = s_csamul_rca16_and13_7 ^ s_csamul_rca16_fa14_6_xor1;
  assign s_csamul_rca16_fa13_7_and0 = s_csamul_rca16_and13_7 & s_csamul_rca16_fa14_6_xor1;
  assign s_csamul_rca16_fa13_7_xor1 = s_csamul_rca16_fa13_7_xor0 ^ s_csamul_rca16_fa13_6_or0;
  assign s_csamul_rca16_fa13_7_and1 = s_csamul_rca16_fa13_7_xor0 & s_csamul_rca16_fa13_6_or0;
  assign s_csamul_rca16_fa13_7_or0 = s_csamul_rca16_fa13_7_and0 | s_csamul_rca16_fa13_7_and1;
  assign s_csamul_rca16_and14_7 = a[14] & b[7];
  assign s_csamul_rca16_fa14_7_xor0 = s_csamul_rca16_and14_7 ^ s_csamul_rca16_ha15_6_xor0;
  assign s_csamul_rca16_fa14_7_and0 = s_csamul_rca16_and14_7 & s_csamul_rca16_ha15_6_xor0;
  assign s_csamul_rca16_fa14_7_xor1 = s_csamul_rca16_fa14_7_xor0 ^ s_csamul_rca16_fa14_6_or0;
  assign s_csamul_rca16_fa14_7_and1 = s_csamul_rca16_fa14_7_xor0 & s_csamul_rca16_fa14_6_or0;
  assign s_csamul_rca16_fa14_7_or0 = s_csamul_rca16_fa14_7_and0 | s_csamul_rca16_fa14_7_and1;
  assign s_csamul_rca16_nand15_7 = ~(a[15] & b[7]);
  assign s_csamul_rca16_ha15_7_xor0 = s_csamul_rca16_nand15_7 ^ s_csamul_rca16_ha15_6_and0;
  assign s_csamul_rca16_ha15_7_and0 = s_csamul_rca16_nand15_7 & s_csamul_rca16_ha15_6_and0;
  assign s_csamul_rca16_and0_8 = a[0] & b[8];
  assign s_csamul_rca16_fa0_8_xor0 = s_csamul_rca16_and0_8 ^ s_csamul_rca16_fa1_7_xor1;
  assign s_csamul_rca16_fa0_8_and0 = s_csamul_rca16_and0_8 & s_csamul_rca16_fa1_7_xor1;
  assign s_csamul_rca16_fa0_8_xor1 = s_csamul_rca16_fa0_8_xor0 ^ s_csamul_rca16_fa0_7_or0;
  assign s_csamul_rca16_fa0_8_and1 = s_csamul_rca16_fa0_8_xor0 & s_csamul_rca16_fa0_7_or0;
  assign s_csamul_rca16_fa0_8_or0 = s_csamul_rca16_fa0_8_and0 | s_csamul_rca16_fa0_8_and1;
  assign s_csamul_rca16_and1_8 = a[1] & b[8];
  assign s_csamul_rca16_fa1_8_xor0 = s_csamul_rca16_and1_8 ^ s_csamul_rca16_fa2_7_xor1;
  assign s_csamul_rca16_fa1_8_and0 = s_csamul_rca16_and1_8 & s_csamul_rca16_fa2_7_xor1;
  assign s_csamul_rca16_fa1_8_xor1 = s_csamul_rca16_fa1_8_xor0 ^ s_csamul_rca16_fa1_7_or0;
  assign s_csamul_rca16_fa1_8_and1 = s_csamul_rca16_fa1_8_xor0 & s_csamul_rca16_fa1_7_or0;
  assign s_csamul_rca16_fa1_8_or0 = s_csamul_rca16_fa1_8_and0 | s_csamul_rca16_fa1_8_and1;
  assign s_csamul_rca16_and2_8 = a[2] & b[8];
  assign s_csamul_rca16_fa2_8_xor0 = s_csamul_rca16_and2_8 ^ s_csamul_rca16_fa3_7_xor1;
  assign s_csamul_rca16_fa2_8_and0 = s_csamul_rca16_and2_8 & s_csamul_rca16_fa3_7_xor1;
  assign s_csamul_rca16_fa2_8_xor1 = s_csamul_rca16_fa2_8_xor0 ^ s_csamul_rca16_fa2_7_or0;
  assign s_csamul_rca16_fa2_8_and1 = s_csamul_rca16_fa2_8_xor0 & s_csamul_rca16_fa2_7_or0;
  assign s_csamul_rca16_fa2_8_or0 = s_csamul_rca16_fa2_8_and0 | s_csamul_rca16_fa2_8_and1;
  assign s_csamul_rca16_and3_8 = a[3] & b[8];
  assign s_csamul_rca16_fa3_8_xor0 = s_csamul_rca16_and3_8 ^ s_csamul_rca16_fa4_7_xor1;
  assign s_csamul_rca16_fa3_8_and0 = s_csamul_rca16_and3_8 & s_csamul_rca16_fa4_7_xor1;
  assign s_csamul_rca16_fa3_8_xor1 = s_csamul_rca16_fa3_8_xor0 ^ s_csamul_rca16_fa3_7_or0;
  assign s_csamul_rca16_fa3_8_and1 = s_csamul_rca16_fa3_8_xor0 & s_csamul_rca16_fa3_7_or0;
  assign s_csamul_rca16_fa3_8_or0 = s_csamul_rca16_fa3_8_and0 | s_csamul_rca16_fa3_8_and1;
  assign s_csamul_rca16_and4_8 = a[4] & b[8];
  assign s_csamul_rca16_fa4_8_xor0 = s_csamul_rca16_and4_8 ^ s_csamul_rca16_fa5_7_xor1;
  assign s_csamul_rca16_fa4_8_and0 = s_csamul_rca16_and4_8 & s_csamul_rca16_fa5_7_xor1;
  assign s_csamul_rca16_fa4_8_xor1 = s_csamul_rca16_fa4_8_xor0 ^ s_csamul_rca16_fa4_7_or0;
  assign s_csamul_rca16_fa4_8_and1 = s_csamul_rca16_fa4_8_xor0 & s_csamul_rca16_fa4_7_or0;
  assign s_csamul_rca16_fa4_8_or0 = s_csamul_rca16_fa4_8_and0 | s_csamul_rca16_fa4_8_and1;
  assign s_csamul_rca16_and5_8 = a[5] & b[8];
  assign s_csamul_rca16_fa5_8_xor0 = s_csamul_rca16_and5_8 ^ s_csamul_rca16_fa6_7_xor1;
  assign s_csamul_rca16_fa5_8_and0 = s_csamul_rca16_and5_8 & s_csamul_rca16_fa6_7_xor1;
  assign s_csamul_rca16_fa5_8_xor1 = s_csamul_rca16_fa5_8_xor0 ^ s_csamul_rca16_fa5_7_or0;
  assign s_csamul_rca16_fa5_8_and1 = s_csamul_rca16_fa5_8_xor0 & s_csamul_rca16_fa5_7_or0;
  assign s_csamul_rca16_fa5_8_or0 = s_csamul_rca16_fa5_8_and0 | s_csamul_rca16_fa5_8_and1;
  assign s_csamul_rca16_and6_8 = a[6] & b[8];
  assign s_csamul_rca16_fa6_8_xor0 = s_csamul_rca16_and6_8 ^ s_csamul_rca16_fa7_7_xor1;
  assign s_csamul_rca16_fa6_8_and0 = s_csamul_rca16_and6_8 & s_csamul_rca16_fa7_7_xor1;
  assign s_csamul_rca16_fa6_8_xor1 = s_csamul_rca16_fa6_8_xor0 ^ s_csamul_rca16_fa6_7_or0;
  assign s_csamul_rca16_fa6_8_and1 = s_csamul_rca16_fa6_8_xor0 & s_csamul_rca16_fa6_7_or0;
  assign s_csamul_rca16_fa6_8_or0 = s_csamul_rca16_fa6_8_and0 | s_csamul_rca16_fa6_8_and1;
  assign s_csamul_rca16_and7_8 = a[7] & b[8];
  assign s_csamul_rca16_fa7_8_xor0 = s_csamul_rca16_and7_8 ^ s_csamul_rca16_fa8_7_xor1;
  assign s_csamul_rca16_fa7_8_and0 = s_csamul_rca16_and7_8 & s_csamul_rca16_fa8_7_xor1;
  assign s_csamul_rca16_fa7_8_xor1 = s_csamul_rca16_fa7_8_xor0 ^ s_csamul_rca16_fa7_7_or0;
  assign s_csamul_rca16_fa7_8_and1 = s_csamul_rca16_fa7_8_xor0 & s_csamul_rca16_fa7_7_or0;
  assign s_csamul_rca16_fa7_8_or0 = s_csamul_rca16_fa7_8_and0 | s_csamul_rca16_fa7_8_and1;
  assign s_csamul_rca16_and8_8 = a[8] & b[8];
  assign s_csamul_rca16_fa8_8_xor0 = s_csamul_rca16_and8_8 ^ s_csamul_rca16_fa9_7_xor1;
  assign s_csamul_rca16_fa8_8_and0 = s_csamul_rca16_and8_8 & s_csamul_rca16_fa9_7_xor1;
  assign s_csamul_rca16_fa8_8_xor1 = s_csamul_rca16_fa8_8_xor0 ^ s_csamul_rca16_fa8_7_or0;
  assign s_csamul_rca16_fa8_8_and1 = s_csamul_rca16_fa8_8_xor0 & s_csamul_rca16_fa8_7_or0;
  assign s_csamul_rca16_fa8_8_or0 = s_csamul_rca16_fa8_8_and0 | s_csamul_rca16_fa8_8_and1;
  assign s_csamul_rca16_and9_8 = a[9] & b[8];
  assign s_csamul_rca16_fa9_8_xor0 = s_csamul_rca16_and9_8 ^ s_csamul_rca16_fa10_7_xor1;
  assign s_csamul_rca16_fa9_8_and0 = s_csamul_rca16_and9_8 & s_csamul_rca16_fa10_7_xor1;
  assign s_csamul_rca16_fa9_8_xor1 = s_csamul_rca16_fa9_8_xor0 ^ s_csamul_rca16_fa9_7_or0;
  assign s_csamul_rca16_fa9_8_and1 = s_csamul_rca16_fa9_8_xor0 & s_csamul_rca16_fa9_7_or0;
  assign s_csamul_rca16_fa9_8_or0 = s_csamul_rca16_fa9_8_and0 | s_csamul_rca16_fa9_8_and1;
  assign s_csamul_rca16_and10_8 = a[10] & b[8];
  assign s_csamul_rca16_fa10_8_xor0 = s_csamul_rca16_and10_8 ^ s_csamul_rca16_fa11_7_xor1;
  assign s_csamul_rca16_fa10_8_and0 = s_csamul_rca16_and10_8 & s_csamul_rca16_fa11_7_xor1;
  assign s_csamul_rca16_fa10_8_xor1 = s_csamul_rca16_fa10_8_xor0 ^ s_csamul_rca16_fa10_7_or0;
  assign s_csamul_rca16_fa10_8_and1 = s_csamul_rca16_fa10_8_xor0 & s_csamul_rca16_fa10_7_or0;
  assign s_csamul_rca16_fa10_8_or0 = s_csamul_rca16_fa10_8_and0 | s_csamul_rca16_fa10_8_and1;
  assign s_csamul_rca16_and11_8 = a[11] & b[8];
  assign s_csamul_rca16_fa11_8_xor0 = s_csamul_rca16_and11_8 ^ s_csamul_rca16_fa12_7_xor1;
  assign s_csamul_rca16_fa11_8_and0 = s_csamul_rca16_and11_8 & s_csamul_rca16_fa12_7_xor1;
  assign s_csamul_rca16_fa11_8_xor1 = s_csamul_rca16_fa11_8_xor0 ^ s_csamul_rca16_fa11_7_or0;
  assign s_csamul_rca16_fa11_8_and1 = s_csamul_rca16_fa11_8_xor0 & s_csamul_rca16_fa11_7_or0;
  assign s_csamul_rca16_fa11_8_or0 = s_csamul_rca16_fa11_8_and0 | s_csamul_rca16_fa11_8_and1;
  assign s_csamul_rca16_and12_8 = a[12] & b[8];
  assign s_csamul_rca16_fa12_8_xor0 = s_csamul_rca16_and12_8 ^ s_csamul_rca16_fa13_7_xor1;
  assign s_csamul_rca16_fa12_8_and0 = s_csamul_rca16_and12_8 & s_csamul_rca16_fa13_7_xor1;
  assign s_csamul_rca16_fa12_8_xor1 = s_csamul_rca16_fa12_8_xor0 ^ s_csamul_rca16_fa12_7_or0;
  assign s_csamul_rca16_fa12_8_and1 = s_csamul_rca16_fa12_8_xor0 & s_csamul_rca16_fa12_7_or0;
  assign s_csamul_rca16_fa12_8_or0 = s_csamul_rca16_fa12_8_and0 | s_csamul_rca16_fa12_8_and1;
  assign s_csamul_rca16_and13_8 = a[13] & b[8];
  assign s_csamul_rca16_fa13_8_xor0 = s_csamul_rca16_and13_8 ^ s_csamul_rca16_fa14_7_xor1;
  assign s_csamul_rca16_fa13_8_and0 = s_csamul_rca16_and13_8 & s_csamul_rca16_fa14_7_xor1;
  assign s_csamul_rca16_fa13_8_xor1 = s_csamul_rca16_fa13_8_xor0 ^ s_csamul_rca16_fa13_7_or0;
  assign s_csamul_rca16_fa13_8_and1 = s_csamul_rca16_fa13_8_xor0 & s_csamul_rca16_fa13_7_or0;
  assign s_csamul_rca16_fa13_8_or0 = s_csamul_rca16_fa13_8_and0 | s_csamul_rca16_fa13_8_and1;
  assign s_csamul_rca16_and14_8 = a[14] & b[8];
  assign s_csamul_rca16_fa14_8_xor0 = s_csamul_rca16_and14_8 ^ s_csamul_rca16_ha15_7_xor0;
  assign s_csamul_rca16_fa14_8_and0 = s_csamul_rca16_and14_8 & s_csamul_rca16_ha15_7_xor0;
  assign s_csamul_rca16_fa14_8_xor1 = s_csamul_rca16_fa14_8_xor0 ^ s_csamul_rca16_fa14_7_or0;
  assign s_csamul_rca16_fa14_8_and1 = s_csamul_rca16_fa14_8_xor0 & s_csamul_rca16_fa14_7_or0;
  assign s_csamul_rca16_fa14_8_or0 = s_csamul_rca16_fa14_8_and0 | s_csamul_rca16_fa14_8_and1;
  assign s_csamul_rca16_nand15_8 = ~(a[15] & b[8]);
  assign s_csamul_rca16_ha15_8_xor0 = s_csamul_rca16_nand15_8 ^ s_csamul_rca16_ha15_7_and0;
  assign s_csamul_rca16_ha15_8_and0 = s_csamul_rca16_nand15_8 & s_csamul_rca16_ha15_7_and0;
  assign s_csamul_rca16_and0_9 = a[0] & b[9];
  assign s_csamul_rca16_fa0_9_xor0 = s_csamul_rca16_and0_9 ^ s_csamul_rca16_fa1_8_xor1;
  assign s_csamul_rca16_fa0_9_and0 = s_csamul_rca16_and0_9 & s_csamul_rca16_fa1_8_xor1;
  assign s_csamul_rca16_fa0_9_xor1 = s_csamul_rca16_fa0_9_xor0 ^ s_csamul_rca16_fa0_8_or0;
  assign s_csamul_rca16_fa0_9_and1 = s_csamul_rca16_fa0_9_xor0 & s_csamul_rca16_fa0_8_or0;
  assign s_csamul_rca16_fa0_9_or0 = s_csamul_rca16_fa0_9_and0 | s_csamul_rca16_fa0_9_and1;
  assign s_csamul_rca16_and1_9 = a[1] & b[9];
  assign s_csamul_rca16_fa1_9_xor0 = s_csamul_rca16_and1_9 ^ s_csamul_rca16_fa2_8_xor1;
  assign s_csamul_rca16_fa1_9_and0 = s_csamul_rca16_and1_9 & s_csamul_rca16_fa2_8_xor1;
  assign s_csamul_rca16_fa1_9_xor1 = s_csamul_rca16_fa1_9_xor0 ^ s_csamul_rca16_fa1_8_or0;
  assign s_csamul_rca16_fa1_9_and1 = s_csamul_rca16_fa1_9_xor0 & s_csamul_rca16_fa1_8_or0;
  assign s_csamul_rca16_fa1_9_or0 = s_csamul_rca16_fa1_9_and0 | s_csamul_rca16_fa1_9_and1;
  assign s_csamul_rca16_and2_9 = a[2] & b[9];
  assign s_csamul_rca16_fa2_9_xor0 = s_csamul_rca16_and2_9 ^ s_csamul_rca16_fa3_8_xor1;
  assign s_csamul_rca16_fa2_9_and0 = s_csamul_rca16_and2_9 & s_csamul_rca16_fa3_8_xor1;
  assign s_csamul_rca16_fa2_9_xor1 = s_csamul_rca16_fa2_9_xor0 ^ s_csamul_rca16_fa2_8_or0;
  assign s_csamul_rca16_fa2_9_and1 = s_csamul_rca16_fa2_9_xor0 & s_csamul_rca16_fa2_8_or0;
  assign s_csamul_rca16_fa2_9_or0 = s_csamul_rca16_fa2_9_and0 | s_csamul_rca16_fa2_9_and1;
  assign s_csamul_rca16_and3_9 = a[3] & b[9];
  assign s_csamul_rca16_fa3_9_xor0 = s_csamul_rca16_and3_9 ^ s_csamul_rca16_fa4_8_xor1;
  assign s_csamul_rca16_fa3_9_and0 = s_csamul_rca16_and3_9 & s_csamul_rca16_fa4_8_xor1;
  assign s_csamul_rca16_fa3_9_xor1 = s_csamul_rca16_fa3_9_xor0 ^ s_csamul_rca16_fa3_8_or0;
  assign s_csamul_rca16_fa3_9_and1 = s_csamul_rca16_fa3_9_xor0 & s_csamul_rca16_fa3_8_or0;
  assign s_csamul_rca16_fa3_9_or0 = s_csamul_rca16_fa3_9_and0 | s_csamul_rca16_fa3_9_and1;
  assign s_csamul_rca16_and4_9 = a[4] & b[9];
  assign s_csamul_rca16_fa4_9_xor0 = s_csamul_rca16_and4_9 ^ s_csamul_rca16_fa5_8_xor1;
  assign s_csamul_rca16_fa4_9_and0 = s_csamul_rca16_and4_9 & s_csamul_rca16_fa5_8_xor1;
  assign s_csamul_rca16_fa4_9_xor1 = s_csamul_rca16_fa4_9_xor0 ^ s_csamul_rca16_fa4_8_or0;
  assign s_csamul_rca16_fa4_9_and1 = s_csamul_rca16_fa4_9_xor0 & s_csamul_rca16_fa4_8_or0;
  assign s_csamul_rca16_fa4_9_or0 = s_csamul_rca16_fa4_9_and0 | s_csamul_rca16_fa4_9_and1;
  assign s_csamul_rca16_and5_9 = a[5] & b[9];
  assign s_csamul_rca16_fa5_9_xor0 = s_csamul_rca16_and5_9 ^ s_csamul_rca16_fa6_8_xor1;
  assign s_csamul_rca16_fa5_9_and0 = s_csamul_rca16_and5_9 & s_csamul_rca16_fa6_8_xor1;
  assign s_csamul_rca16_fa5_9_xor1 = s_csamul_rca16_fa5_9_xor0 ^ s_csamul_rca16_fa5_8_or0;
  assign s_csamul_rca16_fa5_9_and1 = s_csamul_rca16_fa5_9_xor0 & s_csamul_rca16_fa5_8_or0;
  assign s_csamul_rca16_fa5_9_or0 = s_csamul_rca16_fa5_9_and0 | s_csamul_rca16_fa5_9_and1;
  assign s_csamul_rca16_and6_9 = a[6] & b[9];
  assign s_csamul_rca16_fa6_9_xor0 = s_csamul_rca16_and6_9 ^ s_csamul_rca16_fa7_8_xor1;
  assign s_csamul_rca16_fa6_9_and0 = s_csamul_rca16_and6_9 & s_csamul_rca16_fa7_8_xor1;
  assign s_csamul_rca16_fa6_9_xor1 = s_csamul_rca16_fa6_9_xor0 ^ s_csamul_rca16_fa6_8_or0;
  assign s_csamul_rca16_fa6_9_and1 = s_csamul_rca16_fa6_9_xor0 & s_csamul_rca16_fa6_8_or0;
  assign s_csamul_rca16_fa6_9_or0 = s_csamul_rca16_fa6_9_and0 | s_csamul_rca16_fa6_9_and1;
  assign s_csamul_rca16_and7_9 = a[7] & b[9];
  assign s_csamul_rca16_fa7_9_xor0 = s_csamul_rca16_and7_9 ^ s_csamul_rca16_fa8_8_xor1;
  assign s_csamul_rca16_fa7_9_and0 = s_csamul_rca16_and7_9 & s_csamul_rca16_fa8_8_xor1;
  assign s_csamul_rca16_fa7_9_xor1 = s_csamul_rca16_fa7_9_xor0 ^ s_csamul_rca16_fa7_8_or0;
  assign s_csamul_rca16_fa7_9_and1 = s_csamul_rca16_fa7_9_xor0 & s_csamul_rca16_fa7_8_or0;
  assign s_csamul_rca16_fa7_9_or0 = s_csamul_rca16_fa7_9_and0 | s_csamul_rca16_fa7_9_and1;
  assign s_csamul_rca16_and8_9 = a[8] & b[9];
  assign s_csamul_rca16_fa8_9_xor0 = s_csamul_rca16_and8_9 ^ s_csamul_rca16_fa9_8_xor1;
  assign s_csamul_rca16_fa8_9_and0 = s_csamul_rca16_and8_9 & s_csamul_rca16_fa9_8_xor1;
  assign s_csamul_rca16_fa8_9_xor1 = s_csamul_rca16_fa8_9_xor0 ^ s_csamul_rca16_fa8_8_or0;
  assign s_csamul_rca16_fa8_9_and1 = s_csamul_rca16_fa8_9_xor0 & s_csamul_rca16_fa8_8_or0;
  assign s_csamul_rca16_fa8_9_or0 = s_csamul_rca16_fa8_9_and0 | s_csamul_rca16_fa8_9_and1;
  assign s_csamul_rca16_and9_9 = a[9] & b[9];
  assign s_csamul_rca16_fa9_9_xor0 = s_csamul_rca16_and9_9 ^ s_csamul_rca16_fa10_8_xor1;
  assign s_csamul_rca16_fa9_9_and0 = s_csamul_rca16_and9_9 & s_csamul_rca16_fa10_8_xor1;
  assign s_csamul_rca16_fa9_9_xor1 = s_csamul_rca16_fa9_9_xor0 ^ s_csamul_rca16_fa9_8_or0;
  assign s_csamul_rca16_fa9_9_and1 = s_csamul_rca16_fa9_9_xor0 & s_csamul_rca16_fa9_8_or0;
  assign s_csamul_rca16_fa9_9_or0 = s_csamul_rca16_fa9_9_and0 | s_csamul_rca16_fa9_9_and1;
  assign s_csamul_rca16_and10_9 = a[10] & b[9];
  assign s_csamul_rca16_fa10_9_xor0 = s_csamul_rca16_and10_9 ^ s_csamul_rca16_fa11_8_xor1;
  assign s_csamul_rca16_fa10_9_and0 = s_csamul_rca16_and10_9 & s_csamul_rca16_fa11_8_xor1;
  assign s_csamul_rca16_fa10_9_xor1 = s_csamul_rca16_fa10_9_xor0 ^ s_csamul_rca16_fa10_8_or0;
  assign s_csamul_rca16_fa10_9_and1 = s_csamul_rca16_fa10_9_xor0 & s_csamul_rca16_fa10_8_or0;
  assign s_csamul_rca16_fa10_9_or0 = s_csamul_rca16_fa10_9_and0 | s_csamul_rca16_fa10_9_and1;
  assign s_csamul_rca16_and11_9 = a[11] & b[9];
  assign s_csamul_rca16_fa11_9_xor0 = s_csamul_rca16_and11_9 ^ s_csamul_rca16_fa12_8_xor1;
  assign s_csamul_rca16_fa11_9_and0 = s_csamul_rca16_and11_9 & s_csamul_rca16_fa12_8_xor1;
  assign s_csamul_rca16_fa11_9_xor1 = s_csamul_rca16_fa11_9_xor0 ^ s_csamul_rca16_fa11_8_or0;
  assign s_csamul_rca16_fa11_9_and1 = s_csamul_rca16_fa11_9_xor0 & s_csamul_rca16_fa11_8_or0;
  assign s_csamul_rca16_fa11_9_or0 = s_csamul_rca16_fa11_9_and0 | s_csamul_rca16_fa11_9_and1;
  assign s_csamul_rca16_and12_9 = a[12] & b[9];
  assign s_csamul_rca16_fa12_9_xor0 = s_csamul_rca16_and12_9 ^ s_csamul_rca16_fa13_8_xor1;
  assign s_csamul_rca16_fa12_9_and0 = s_csamul_rca16_and12_9 & s_csamul_rca16_fa13_8_xor1;
  assign s_csamul_rca16_fa12_9_xor1 = s_csamul_rca16_fa12_9_xor0 ^ s_csamul_rca16_fa12_8_or0;
  assign s_csamul_rca16_fa12_9_and1 = s_csamul_rca16_fa12_9_xor0 & s_csamul_rca16_fa12_8_or0;
  assign s_csamul_rca16_fa12_9_or0 = s_csamul_rca16_fa12_9_and0 | s_csamul_rca16_fa12_9_and1;
  assign s_csamul_rca16_and13_9 = a[13] & b[9];
  assign s_csamul_rca16_fa13_9_xor0 = s_csamul_rca16_and13_9 ^ s_csamul_rca16_fa14_8_xor1;
  assign s_csamul_rca16_fa13_9_and0 = s_csamul_rca16_and13_9 & s_csamul_rca16_fa14_8_xor1;
  assign s_csamul_rca16_fa13_9_xor1 = s_csamul_rca16_fa13_9_xor0 ^ s_csamul_rca16_fa13_8_or0;
  assign s_csamul_rca16_fa13_9_and1 = s_csamul_rca16_fa13_9_xor0 & s_csamul_rca16_fa13_8_or0;
  assign s_csamul_rca16_fa13_9_or0 = s_csamul_rca16_fa13_9_and0 | s_csamul_rca16_fa13_9_and1;
  assign s_csamul_rca16_and14_9 = a[14] & b[9];
  assign s_csamul_rca16_fa14_9_xor0 = s_csamul_rca16_and14_9 ^ s_csamul_rca16_ha15_8_xor0;
  assign s_csamul_rca16_fa14_9_and0 = s_csamul_rca16_and14_9 & s_csamul_rca16_ha15_8_xor0;
  assign s_csamul_rca16_fa14_9_xor1 = s_csamul_rca16_fa14_9_xor0 ^ s_csamul_rca16_fa14_8_or0;
  assign s_csamul_rca16_fa14_9_and1 = s_csamul_rca16_fa14_9_xor0 & s_csamul_rca16_fa14_8_or0;
  assign s_csamul_rca16_fa14_9_or0 = s_csamul_rca16_fa14_9_and0 | s_csamul_rca16_fa14_9_and1;
  assign s_csamul_rca16_nand15_9 = ~(a[15] & b[9]);
  assign s_csamul_rca16_ha15_9_xor0 = s_csamul_rca16_nand15_9 ^ s_csamul_rca16_ha15_8_and0;
  assign s_csamul_rca16_ha15_9_and0 = s_csamul_rca16_nand15_9 & s_csamul_rca16_ha15_8_and0;
  assign s_csamul_rca16_and0_10 = a[0] & b[10];
  assign s_csamul_rca16_fa0_10_xor0 = s_csamul_rca16_and0_10 ^ s_csamul_rca16_fa1_9_xor1;
  assign s_csamul_rca16_fa0_10_and0 = s_csamul_rca16_and0_10 & s_csamul_rca16_fa1_9_xor1;
  assign s_csamul_rca16_fa0_10_xor1 = s_csamul_rca16_fa0_10_xor0 ^ s_csamul_rca16_fa0_9_or0;
  assign s_csamul_rca16_fa0_10_and1 = s_csamul_rca16_fa0_10_xor0 & s_csamul_rca16_fa0_9_or0;
  assign s_csamul_rca16_fa0_10_or0 = s_csamul_rca16_fa0_10_and0 | s_csamul_rca16_fa0_10_and1;
  assign s_csamul_rca16_and1_10 = a[1] & b[10];
  assign s_csamul_rca16_fa1_10_xor0 = s_csamul_rca16_and1_10 ^ s_csamul_rca16_fa2_9_xor1;
  assign s_csamul_rca16_fa1_10_and0 = s_csamul_rca16_and1_10 & s_csamul_rca16_fa2_9_xor1;
  assign s_csamul_rca16_fa1_10_xor1 = s_csamul_rca16_fa1_10_xor0 ^ s_csamul_rca16_fa1_9_or0;
  assign s_csamul_rca16_fa1_10_and1 = s_csamul_rca16_fa1_10_xor0 & s_csamul_rca16_fa1_9_or0;
  assign s_csamul_rca16_fa1_10_or0 = s_csamul_rca16_fa1_10_and0 | s_csamul_rca16_fa1_10_and1;
  assign s_csamul_rca16_and2_10 = a[2] & b[10];
  assign s_csamul_rca16_fa2_10_xor0 = s_csamul_rca16_and2_10 ^ s_csamul_rca16_fa3_9_xor1;
  assign s_csamul_rca16_fa2_10_and0 = s_csamul_rca16_and2_10 & s_csamul_rca16_fa3_9_xor1;
  assign s_csamul_rca16_fa2_10_xor1 = s_csamul_rca16_fa2_10_xor0 ^ s_csamul_rca16_fa2_9_or0;
  assign s_csamul_rca16_fa2_10_and1 = s_csamul_rca16_fa2_10_xor0 & s_csamul_rca16_fa2_9_or0;
  assign s_csamul_rca16_fa2_10_or0 = s_csamul_rca16_fa2_10_and0 | s_csamul_rca16_fa2_10_and1;
  assign s_csamul_rca16_and3_10 = a[3] & b[10];
  assign s_csamul_rca16_fa3_10_xor0 = s_csamul_rca16_and3_10 ^ s_csamul_rca16_fa4_9_xor1;
  assign s_csamul_rca16_fa3_10_and0 = s_csamul_rca16_and3_10 & s_csamul_rca16_fa4_9_xor1;
  assign s_csamul_rca16_fa3_10_xor1 = s_csamul_rca16_fa3_10_xor0 ^ s_csamul_rca16_fa3_9_or0;
  assign s_csamul_rca16_fa3_10_and1 = s_csamul_rca16_fa3_10_xor0 & s_csamul_rca16_fa3_9_or0;
  assign s_csamul_rca16_fa3_10_or0 = s_csamul_rca16_fa3_10_and0 | s_csamul_rca16_fa3_10_and1;
  assign s_csamul_rca16_and4_10 = a[4] & b[10];
  assign s_csamul_rca16_fa4_10_xor0 = s_csamul_rca16_and4_10 ^ s_csamul_rca16_fa5_9_xor1;
  assign s_csamul_rca16_fa4_10_and0 = s_csamul_rca16_and4_10 & s_csamul_rca16_fa5_9_xor1;
  assign s_csamul_rca16_fa4_10_xor1 = s_csamul_rca16_fa4_10_xor0 ^ s_csamul_rca16_fa4_9_or0;
  assign s_csamul_rca16_fa4_10_and1 = s_csamul_rca16_fa4_10_xor0 & s_csamul_rca16_fa4_9_or0;
  assign s_csamul_rca16_fa4_10_or0 = s_csamul_rca16_fa4_10_and0 | s_csamul_rca16_fa4_10_and1;
  assign s_csamul_rca16_and5_10 = a[5] & b[10];
  assign s_csamul_rca16_fa5_10_xor0 = s_csamul_rca16_and5_10 ^ s_csamul_rca16_fa6_9_xor1;
  assign s_csamul_rca16_fa5_10_and0 = s_csamul_rca16_and5_10 & s_csamul_rca16_fa6_9_xor1;
  assign s_csamul_rca16_fa5_10_xor1 = s_csamul_rca16_fa5_10_xor0 ^ s_csamul_rca16_fa5_9_or0;
  assign s_csamul_rca16_fa5_10_and1 = s_csamul_rca16_fa5_10_xor0 & s_csamul_rca16_fa5_9_or0;
  assign s_csamul_rca16_fa5_10_or0 = s_csamul_rca16_fa5_10_and0 | s_csamul_rca16_fa5_10_and1;
  assign s_csamul_rca16_and6_10 = a[6] & b[10];
  assign s_csamul_rca16_fa6_10_xor0 = s_csamul_rca16_and6_10 ^ s_csamul_rca16_fa7_9_xor1;
  assign s_csamul_rca16_fa6_10_and0 = s_csamul_rca16_and6_10 & s_csamul_rca16_fa7_9_xor1;
  assign s_csamul_rca16_fa6_10_xor1 = s_csamul_rca16_fa6_10_xor0 ^ s_csamul_rca16_fa6_9_or0;
  assign s_csamul_rca16_fa6_10_and1 = s_csamul_rca16_fa6_10_xor0 & s_csamul_rca16_fa6_9_or0;
  assign s_csamul_rca16_fa6_10_or0 = s_csamul_rca16_fa6_10_and0 | s_csamul_rca16_fa6_10_and1;
  assign s_csamul_rca16_and7_10 = a[7] & b[10];
  assign s_csamul_rca16_fa7_10_xor0 = s_csamul_rca16_and7_10 ^ s_csamul_rca16_fa8_9_xor1;
  assign s_csamul_rca16_fa7_10_and0 = s_csamul_rca16_and7_10 & s_csamul_rca16_fa8_9_xor1;
  assign s_csamul_rca16_fa7_10_xor1 = s_csamul_rca16_fa7_10_xor0 ^ s_csamul_rca16_fa7_9_or0;
  assign s_csamul_rca16_fa7_10_and1 = s_csamul_rca16_fa7_10_xor0 & s_csamul_rca16_fa7_9_or0;
  assign s_csamul_rca16_fa7_10_or0 = s_csamul_rca16_fa7_10_and0 | s_csamul_rca16_fa7_10_and1;
  assign s_csamul_rca16_and8_10 = a[8] & b[10];
  assign s_csamul_rca16_fa8_10_xor0 = s_csamul_rca16_and8_10 ^ s_csamul_rca16_fa9_9_xor1;
  assign s_csamul_rca16_fa8_10_and0 = s_csamul_rca16_and8_10 & s_csamul_rca16_fa9_9_xor1;
  assign s_csamul_rca16_fa8_10_xor1 = s_csamul_rca16_fa8_10_xor0 ^ s_csamul_rca16_fa8_9_or0;
  assign s_csamul_rca16_fa8_10_and1 = s_csamul_rca16_fa8_10_xor0 & s_csamul_rca16_fa8_9_or0;
  assign s_csamul_rca16_fa8_10_or0 = s_csamul_rca16_fa8_10_and0 | s_csamul_rca16_fa8_10_and1;
  assign s_csamul_rca16_and9_10 = a[9] & b[10];
  assign s_csamul_rca16_fa9_10_xor0 = s_csamul_rca16_and9_10 ^ s_csamul_rca16_fa10_9_xor1;
  assign s_csamul_rca16_fa9_10_and0 = s_csamul_rca16_and9_10 & s_csamul_rca16_fa10_9_xor1;
  assign s_csamul_rca16_fa9_10_xor1 = s_csamul_rca16_fa9_10_xor0 ^ s_csamul_rca16_fa9_9_or0;
  assign s_csamul_rca16_fa9_10_and1 = s_csamul_rca16_fa9_10_xor0 & s_csamul_rca16_fa9_9_or0;
  assign s_csamul_rca16_fa9_10_or0 = s_csamul_rca16_fa9_10_and0 | s_csamul_rca16_fa9_10_and1;
  assign s_csamul_rca16_and10_10 = a[10] & b[10];
  assign s_csamul_rca16_fa10_10_xor0 = s_csamul_rca16_and10_10 ^ s_csamul_rca16_fa11_9_xor1;
  assign s_csamul_rca16_fa10_10_and0 = s_csamul_rca16_and10_10 & s_csamul_rca16_fa11_9_xor1;
  assign s_csamul_rca16_fa10_10_xor1 = s_csamul_rca16_fa10_10_xor0 ^ s_csamul_rca16_fa10_9_or0;
  assign s_csamul_rca16_fa10_10_and1 = s_csamul_rca16_fa10_10_xor0 & s_csamul_rca16_fa10_9_or0;
  assign s_csamul_rca16_fa10_10_or0 = s_csamul_rca16_fa10_10_and0 | s_csamul_rca16_fa10_10_and1;
  assign s_csamul_rca16_and11_10 = a[11] & b[10];
  assign s_csamul_rca16_fa11_10_xor0 = s_csamul_rca16_and11_10 ^ s_csamul_rca16_fa12_9_xor1;
  assign s_csamul_rca16_fa11_10_and0 = s_csamul_rca16_and11_10 & s_csamul_rca16_fa12_9_xor1;
  assign s_csamul_rca16_fa11_10_xor1 = s_csamul_rca16_fa11_10_xor0 ^ s_csamul_rca16_fa11_9_or0;
  assign s_csamul_rca16_fa11_10_and1 = s_csamul_rca16_fa11_10_xor0 & s_csamul_rca16_fa11_9_or0;
  assign s_csamul_rca16_fa11_10_or0 = s_csamul_rca16_fa11_10_and0 | s_csamul_rca16_fa11_10_and1;
  assign s_csamul_rca16_and12_10 = a[12] & b[10];
  assign s_csamul_rca16_fa12_10_xor0 = s_csamul_rca16_and12_10 ^ s_csamul_rca16_fa13_9_xor1;
  assign s_csamul_rca16_fa12_10_and0 = s_csamul_rca16_and12_10 & s_csamul_rca16_fa13_9_xor1;
  assign s_csamul_rca16_fa12_10_xor1 = s_csamul_rca16_fa12_10_xor0 ^ s_csamul_rca16_fa12_9_or0;
  assign s_csamul_rca16_fa12_10_and1 = s_csamul_rca16_fa12_10_xor0 & s_csamul_rca16_fa12_9_or0;
  assign s_csamul_rca16_fa12_10_or0 = s_csamul_rca16_fa12_10_and0 | s_csamul_rca16_fa12_10_and1;
  assign s_csamul_rca16_and13_10 = a[13] & b[10];
  assign s_csamul_rca16_fa13_10_xor0 = s_csamul_rca16_and13_10 ^ s_csamul_rca16_fa14_9_xor1;
  assign s_csamul_rca16_fa13_10_and0 = s_csamul_rca16_and13_10 & s_csamul_rca16_fa14_9_xor1;
  assign s_csamul_rca16_fa13_10_xor1 = s_csamul_rca16_fa13_10_xor0 ^ s_csamul_rca16_fa13_9_or0;
  assign s_csamul_rca16_fa13_10_and1 = s_csamul_rca16_fa13_10_xor0 & s_csamul_rca16_fa13_9_or0;
  assign s_csamul_rca16_fa13_10_or0 = s_csamul_rca16_fa13_10_and0 | s_csamul_rca16_fa13_10_and1;
  assign s_csamul_rca16_and14_10 = a[14] & b[10];
  assign s_csamul_rca16_fa14_10_xor0 = s_csamul_rca16_and14_10 ^ s_csamul_rca16_ha15_9_xor0;
  assign s_csamul_rca16_fa14_10_and0 = s_csamul_rca16_and14_10 & s_csamul_rca16_ha15_9_xor0;
  assign s_csamul_rca16_fa14_10_xor1 = s_csamul_rca16_fa14_10_xor0 ^ s_csamul_rca16_fa14_9_or0;
  assign s_csamul_rca16_fa14_10_and1 = s_csamul_rca16_fa14_10_xor0 & s_csamul_rca16_fa14_9_or0;
  assign s_csamul_rca16_fa14_10_or0 = s_csamul_rca16_fa14_10_and0 | s_csamul_rca16_fa14_10_and1;
  assign s_csamul_rca16_nand15_10 = ~(a[15] & b[10]);
  assign s_csamul_rca16_ha15_10_xor0 = s_csamul_rca16_nand15_10 ^ s_csamul_rca16_ha15_9_and0;
  assign s_csamul_rca16_ha15_10_and0 = s_csamul_rca16_nand15_10 & s_csamul_rca16_ha15_9_and0;
  assign s_csamul_rca16_and0_11 = a[0] & b[11];
  assign s_csamul_rca16_fa0_11_xor0 = s_csamul_rca16_and0_11 ^ s_csamul_rca16_fa1_10_xor1;
  assign s_csamul_rca16_fa0_11_and0 = s_csamul_rca16_and0_11 & s_csamul_rca16_fa1_10_xor1;
  assign s_csamul_rca16_fa0_11_xor1 = s_csamul_rca16_fa0_11_xor0 ^ s_csamul_rca16_fa0_10_or0;
  assign s_csamul_rca16_fa0_11_and1 = s_csamul_rca16_fa0_11_xor0 & s_csamul_rca16_fa0_10_or0;
  assign s_csamul_rca16_fa0_11_or0 = s_csamul_rca16_fa0_11_and0 | s_csamul_rca16_fa0_11_and1;
  assign s_csamul_rca16_and1_11 = a[1] & b[11];
  assign s_csamul_rca16_fa1_11_xor0 = s_csamul_rca16_and1_11 ^ s_csamul_rca16_fa2_10_xor1;
  assign s_csamul_rca16_fa1_11_and0 = s_csamul_rca16_and1_11 & s_csamul_rca16_fa2_10_xor1;
  assign s_csamul_rca16_fa1_11_xor1 = s_csamul_rca16_fa1_11_xor0 ^ s_csamul_rca16_fa1_10_or0;
  assign s_csamul_rca16_fa1_11_and1 = s_csamul_rca16_fa1_11_xor0 & s_csamul_rca16_fa1_10_or0;
  assign s_csamul_rca16_fa1_11_or0 = s_csamul_rca16_fa1_11_and0 | s_csamul_rca16_fa1_11_and1;
  assign s_csamul_rca16_and2_11 = a[2] & b[11];
  assign s_csamul_rca16_fa2_11_xor0 = s_csamul_rca16_and2_11 ^ s_csamul_rca16_fa3_10_xor1;
  assign s_csamul_rca16_fa2_11_and0 = s_csamul_rca16_and2_11 & s_csamul_rca16_fa3_10_xor1;
  assign s_csamul_rca16_fa2_11_xor1 = s_csamul_rca16_fa2_11_xor0 ^ s_csamul_rca16_fa2_10_or0;
  assign s_csamul_rca16_fa2_11_and1 = s_csamul_rca16_fa2_11_xor0 & s_csamul_rca16_fa2_10_or0;
  assign s_csamul_rca16_fa2_11_or0 = s_csamul_rca16_fa2_11_and0 | s_csamul_rca16_fa2_11_and1;
  assign s_csamul_rca16_and3_11 = a[3] & b[11];
  assign s_csamul_rca16_fa3_11_xor0 = s_csamul_rca16_and3_11 ^ s_csamul_rca16_fa4_10_xor1;
  assign s_csamul_rca16_fa3_11_and0 = s_csamul_rca16_and3_11 & s_csamul_rca16_fa4_10_xor1;
  assign s_csamul_rca16_fa3_11_xor1 = s_csamul_rca16_fa3_11_xor0 ^ s_csamul_rca16_fa3_10_or0;
  assign s_csamul_rca16_fa3_11_and1 = s_csamul_rca16_fa3_11_xor0 & s_csamul_rca16_fa3_10_or0;
  assign s_csamul_rca16_fa3_11_or0 = s_csamul_rca16_fa3_11_and0 | s_csamul_rca16_fa3_11_and1;
  assign s_csamul_rca16_and4_11 = a[4] & b[11];
  assign s_csamul_rca16_fa4_11_xor0 = s_csamul_rca16_and4_11 ^ s_csamul_rca16_fa5_10_xor1;
  assign s_csamul_rca16_fa4_11_and0 = s_csamul_rca16_and4_11 & s_csamul_rca16_fa5_10_xor1;
  assign s_csamul_rca16_fa4_11_xor1 = s_csamul_rca16_fa4_11_xor0 ^ s_csamul_rca16_fa4_10_or0;
  assign s_csamul_rca16_fa4_11_and1 = s_csamul_rca16_fa4_11_xor0 & s_csamul_rca16_fa4_10_or0;
  assign s_csamul_rca16_fa4_11_or0 = s_csamul_rca16_fa4_11_and0 | s_csamul_rca16_fa4_11_and1;
  assign s_csamul_rca16_and5_11 = a[5] & b[11];
  assign s_csamul_rca16_fa5_11_xor0 = s_csamul_rca16_and5_11 ^ s_csamul_rca16_fa6_10_xor1;
  assign s_csamul_rca16_fa5_11_and0 = s_csamul_rca16_and5_11 & s_csamul_rca16_fa6_10_xor1;
  assign s_csamul_rca16_fa5_11_xor1 = s_csamul_rca16_fa5_11_xor0 ^ s_csamul_rca16_fa5_10_or0;
  assign s_csamul_rca16_fa5_11_and1 = s_csamul_rca16_fa5_11_xor0 & s_csamul_rca16_fa5_10_or0;
  assign s_csamul_rca16_fa5_11_or0 = s_csamul_rca16_fa5_11_and0 | s_csamul_rca16_fa5_11_and1;
  assign s_csamul_rca16_and6_11 = a[6] & b[11];
  assign s_csamul_rca16_fa6_11_xor0 = s_csamul_rca16_and6_11 ^ s_csamul_rca16_fa7_10_xor1;
  assign s_csamul_rca16_fa6_11_and0 = s_csamul_rca16_and6_11 & s_csamul_rca16_fa7_10_xor1;
  assign s_csamul_rca16_fa6_11_xor1 = s_csamul_rca16_fa6_11_xor0 ^ s_csamul_rca16_fa6_10_or0;
  assign s_csamul_rca16_fa6_11_and1 = s_csamul_rca16_fa6_11_xor0 & s_csamul_rca16_fa6_10_or0;
  assign s_csamul_rca16_fa6_11_or0 = s_csamul_rca16_fa6_11_and0 | s_csamul_rca16_fa6_11_and1;
  assign s_csamul_rca16_and7_11 = a[7] & b[11];
  assign s_csamul_rca16_fa7_11_xor0 = s_csamul_rca16_and7_11 ^ s_csamul_rca16_fa8_10_xor1;
  assign s_csamul_rca16_fa7_11_and0 = s_csamul_rca16_and7_11 & s_csamul_rca16_fa8_10_xor1;
  assign s_csamul_rca16_fa7_11_xor1 = s_csamul_rca16_fa7_11_xor0 ^ s_csamul_rca16_fa7_10_or0;
  assign s_csamul_rca16_fa7_11_and1 = s_csamul_rca16_fa7_11_xor0 & s_csamul_rca16_fa7_10_or0;
  assign s_csamul_rca16_fa7_11_or0 = s_csamul_rca16_fa7_11_and0 | s_csamul_rca16_fa7_11_and1;
  assign s_csamul_rca16_and8_11 = a[8] & b[11];
  assign s_csamul_rca16_fa8_11_xor0 = s_csamul_rca16_and8_11 ^ s_csamul_rca16_fa9_10_xor1;
  assign s_csamul_rca16_fa8_11_and0 = s_csamul_rca16_and8_11 & s_csamul_rca16_fa9_10_xor1;
  assign s_csamul_rca16_fa8_11_xor1 = s_csamul_rca16_fa8_11_xor0 ^ s_csamul_rca16_fa8_10_or0;
  assign s_csamul_rca16_fa8_11_and1 = s_csamul_rca16_fa8_11_xor0 & s_csamul_rca16_fa8_10_or0;
  assign s_csamul_rca16_fa8_11_or0 = s_csamul_rca16_fa8_11_and0 | s_csamul_rca16_fa8_11_and1;
  assign s_csamul_rca16_and9_11 = a[9] & b[11];
  assign s_csamul_rca16_fa9_11_xor0 = s_csamul_rca16_and9_11 ^ s_csamul_rca16_fa10_10_xor1;
  assign s_csamul_rca16_fa9_11_and0 = s_csamul_rca16_and9_11 & s_csamul_rca16_fa10_10_xor1;
  assign s_csamul_rca16_fa9_11_xor1 = s_csamul_rca16_fa9_11_xor0 ^ s_csamul_rca16_fa9_10_or0;
  assign s_csamul_rca16_fa9_11_and1 = s_csamul_rca16_fa9_11_xor0 & s_csamul_rca16_fa9_10_or0;
  assign s_csamul_rca16_fa9_11_or0 = s_csamul_rca16_fa9_11_and0 | s_csamul_rca16_fa9_11_and1;
  assign s_csamul_rca16_and10_11 = a[10] & b[11];
  assign s_csamul_rca16_fa10_11_xor0 = s_csamul_rca16_and10_11 ^ s_csamul_rca16_fa11_10_xor1;
  assign s_csamul_rca16_fa10_11_and0 = s_csamul_rca16_and10_11 & s_csamul_rca16_fa11_10_xor1;
  assign s_csamul_rca16_fa10_11_xor1 = s_csamul_rca16_fa10_11_xor0 ^ s_csamul_rca16_fa10_10_or0;
  assign s_csamul_rca16_fa10_11_and1 = s_csamul_rca16_fa10_11_xor0 & s_csamul_rca16_fa10_10_or0;
  assign s_csamul_rca16_fa10_11_or0 = s_csamul_rca16_fa10_11_and0 | s_csamul_rca16_fa10_11_and1;
  assign s_csamul_rca16_and11_11 = a[11] & b[11];
  assign s_csamul_rca16_fa11_11_xor0 = s_csamul_rca16_and11_11 ^ s_csamul_rca16_fa12_10_xor1;
  assign s_csamul_rca16_fa11_11_and0 = s_csamul_rca16_and11_11 & s_csamul_rca16_fa12_10_xor1;
  assign s_csamul_rca16_fa11_11_xor1 = s_csamul_rca16_fa11_11_xor0 ^ s_csamul_rca16_fa11_10_or0;
  assign s_csamul_rca16_fa11_11_and1 = s_csamul_rca16_fa11_11_xor0 & s_csamul_rca16_fa11_10_or0;
  assign s_csamul_rca16_fa11_11_or0 = s_csamul_rca16_fa11_11_and0 | s_csamul_rca16_fa11_11_and1;
  assign s_csamul_rca16_and12_11 = a[12] & b[11];
  assign s_csamul_rca16_fa12_11_xor0 = s_csamul_rca16_and12_11 ^ s_csamul_rca16_fa13_10_xor1;
  assign s_csamul_rca16_fa12_11_and0 = s_csamul_rca16_and12_11 & s_csamul_rca16_fa13_10_xor1;
  assign s_csamul_rca16_fa12_11_xor1 = s_csamul_rca16_fa12_11_xor0 ^ s_csamul_rca16_fa12_10_or0;
  assign s_csamul_rca16_fa12_11_and1 = s_csamul_rca16_fa12_11_xor0 & s_csamul_rca16_fa12_10_or0;
  assign s_csamul_rca16_fa12_11_or0 = s_csamul_rca16_fa12_11_and0 | s_csamul_rca16_fa12_11_and1;
  assign s_csamul_rca16_and13_11 = a[13] & b[11];
  assign s_csamul_rca16_fa13_11_xor0 = s_csamul_rca16_and13_11 ^ s_csamul_rca16_fa14_10_xor1;
  assign s_csamul_rca16_fa13_11_and0 = s_csamul_rca16_and13_11 & s_csamul_rca16_fa14_10_xor1;
  assign s_csamul_rca16_fa13_11_xor1 = s_csamul_rca16_fa13_11_xor0 ^ s_csamul_rca16_fa13_10_or0;
  assign s_csamul_rca16_fa13_11_and1 = s_csamul_rca16_fa13_11_xor0 & s_csamul_rca16_fa13_10_or0;
  assign s_csamul_rca16_fa13_11_or0 = s_csamul_rca16_fa13_11_and0 | s_csamul_rca16_fa13_11_and1;
  assign s_csamul_rca16_and14_11 = a[14] & b[11];
  assign s_csamul_rca16_fa14_11_xor0 = s_csamul_rca16_and14_11 ^ s_csamul_rca16_ha15_10_xor0;
  assign s_csamul_rca16_fa14_11_and0 = s_csamul_rca16_and14_11 & s_csamul_rca16_ha15_10_xor0;
  assign s_csamul_rca16_fa14_11_xor1 = s_csamul_rca16_fa14_11_xor0 ^ s_csamul_rca16_fa14_10_or0;
  assign s_csamul_rca16_fa14_11_and1 = s_csamul_rca16_fa14_11_xor0 & s_csamul_rca16_fa14_10_or0;
  assign s_csamul_rca16_fa14_11_or0 = s_csamul_rca16_fa14_11_and0 | s_csamul_rca16_fa14_11_and1;
  assign s_csamul_rca16_nand15_11 = ~(a[15] & b[11]);
  assign s_csamul_rca16_ha15_11_xor0 = s_csamul_rca16_nand15_11 ^ s_csamul_rca16_ha15_10_and0;
  assign s_csamul_rca16_ha15_11_and0 = s_csamul_rca16_nand15_11 & s_csamul_rca16_ha15_10_and0;
  assign s_csamul_rca16_and0_12 = a[0] & b[12];
  assign s_csamul_rca16_fa0_12_xor0 = s_csamul_rca16_and0_12 ^ s_csamul_rca16_fa1_11_xor1;
  assign s_csamul_rca16_fa0_12_and0 = s_csamul_rca16_and0_12 & s_csamul_rca16_fa1_11_xor1;
  assign s_csamul_rca16_fa0_12_xor1 = s_csamul_rca16_fa0_12_xor0 ^ s_csamul_rca16_fa0_11_or0;
  assign s_csamul_rca16_fa0_12_and1 = s_csamul_rca16_fa0_12_xor0 & s_csamul_rca16_fa0_11_or0;
  assign s_csamul_rca16_fa0_12_or0 = s_csamul_rca16_fa0_12_and0 | s_csamul_rca16_fa0_12_and1;
  assign s_csamul_rca16_and1_12 = a[1] & b[12];
  assign s_csamul_rca16_fa1_12_xor0 = s_csamul_rca16_and1_12 ^ s_csamul_rca16_fa2_11_xor1;
  assign s_csamul_rca16_fa1_12_and0 = s_csamul_rca16_and1_12 & s_csamul_rca16_fa2_11_xor1;
  assign s_csamul_rca16_fa1_12_xor1 = s_csamul_rca16_fa1_12_xor0 ^ s_csamul_rca16_fa1_11_or0;
  assign s_csamul_rca16_fa1_12_and1 = s_csamul_rca16_fa1_12_xor0 & s_csamul_rca16_fa1_11_or0;
  assign s_csamul_rca16_fa1_12_or0 = s_csamul_rca16_fa1_12_and0 | s_csamul_rca16_fa1_12_and1;
  assign s_csamul_rca16_and2_12 = a[2] & b[12];
  assign s_csamul_rca16_fa2_12_xor0 = s_csamul_rca16_and2_12 ^ s_csamul_rca16_fa3_11_xor1;
  assign s_csamul_rca16_fa2_12_and0 = s_csamul_rca16_and2_12 & s_csamul_rca16_fa3_11_xor1;
  assign s_csamul_rca16_fa2_12_xor1 = s_csamul_rca16_fa2_12_xor0 ^ s_csamul_rca16_fa2_11_or0;
  assign s_csamul_rca16_fa2_12_and1 = s_csamul_rca16_fa2_12_xor0 & s_csamul_rca16_fa2_11_or0;
  assign s_csamul_rca16_fa2_12_or0 = s_csamul_rca16_fa2_12_and0 | s_csamul_rca16_fa2_12_and1;
  assign s_csamul_rca16_and3_12 = a[3] & b[12];
  assign s_csamul_rca16_fa3_12_xor0 = s_csamul_rca16_and3_12 ^ s_csamul_rca16_fa4_11_xor1;
  assign s_csamul_rca16_fa3_12_and0 = s_csamul_rca16_and3_12 & s_csamul_rca16_fa4_11_xor1;
  assign s_csamul_rca16_fa3_12_xor1 = s_csamul_rca16_fa3_12_xor0 ^ s_csamul_rca16_fa3_11_or0;
  assign s_csamul_rca16_fa3_12_and1 = s_csamul_rca16_fa3_12_xor0 & s_csamul_rca16_fa3_11_or0;
  assign s_csamul_rca16_fa3_12_or0 = s_csamul_rca16_fa3_12_and0 | s_csamul_rca16_fa3_12_and1;
  assign s_csamul_rca16_and4_12 = a[4] & b[12];
  assign s_csamul_rca16_fa4_12_xor0 = s_csamul_rca16_and4_12 ^ s_csamul_rca16_fa5_11_xor1;
  assign s_csamul_rca16_fa4_12_and0 = s_csamul_rca16_and4_12 & s_csamul_rca16_fa5_11_xor1;
  assign s_csamul_rca16_fa4_12_xor1 = s_csamul_rca16_fa4_12_xor0 ^ s_csamul_rca16_fa4_11_or0;
  assign s_csamul_rca16_fa4_12_and1 = s_csamul_rca16_fa4_12_xor0 & s_csamul_rca16_fa4_11_or0;
  assign s_csamul_rca16_fa4_12_or0 = s_csamul_rca16_fa4_12_and0 | s_csamul_rca16_fa4_12_and1;
  assign s_csamul_rca16_and5_12 = a[5] & b[12];
  assign s_csamul_rca16_fa5_12_xor0 = s_csamul_rca16_and5_12 ^ s_csamul_rca16_fa6_11_xor1;
  assign s_csamul_rca16_fa5_12_and0 = s_csamul_rca16_and5_12 & s_csamul_rca16_fa6_11_xor1;
  assign s_csamul_rca16_fa5_12_xor1 = s_csamul_rca16_fa5_12_xor0 ^ s_csamul_rca16_fa5_11_or0;
  assign s_csamul_rca16_fa5_12_and1 = s_csamul_rca16_fa5_12_xor0 & s_csamul_rca16_fa5_11_or0;
  assign s_csamul_rca16_fa5_12_or0 = s_csamul_rca16_fa5_12_and0 | s_csamul_rca16_fa5_12_and1;
  assign s_csamul_rca16_and6_12 = a[6] & b[12];
  assign s_csamul_rca16_fa6_12_xor0 = s_csamul_rca16_and6_12 ^ s_csamul_rca16_fa7_11_xor1;
  assign s_csamul_rca16_fa6_12_and0 = s_csamul_rca16_and6_12 & s_csamul_rca16_fa7_11_xor1;
  assign s_csamul_rca16_fa6_12_xor1 = s_csamul_rca16_fa6_12_xor0 ^ s_csamul_rca16_fa6_11_or0;
  assign s_csamul_rca16_fa6_12_and1 = s_csamul_rca16_fa6_12_xor0 & s_csamul_rca16_fa6_11_or0;
  assign s_csamul_rca16_fa6_12_or0 = s_csamul_rca16_fa6_12_and0 | s_csamul_rca16_fa6_12_and1;
  assign s_csamul_rca16_and7_12 = a[7] & b[12];
  assign s_csamul_rca16_fa7_12_xor0 = s_csamul_rca16_and7_12 ^ s_csamul_rca16_fa8_11_xor1;
  assign s_csamul_rca16_fa7_12_and0 = s_csamul_rca16_and7_12 & s_csamul_rca16_fa8_11_xor1;
  assign s_csamul_rca16_fa7_12_xor1 = s_csamul_rca16_fa7_12_xor0 ^ s_csamul_rca16_fa7_11_or0;
  assign s_csamul_rca16_fa7_12_and1 = s_csamul_rca16_fa7_12_xor0 & s_csamul_rca16_fa7_11_or0;
  assign s_csamul_rca16_fa7_12_or0 = s_csamul_rca16_fa7_12_and0 | s_csamul_rca16_fa7_12_and1;
  assign s_csamul_rca16_and8_12 = a[8] & b[12];
  assign s_csamul_rca16_fa8_12_xor0 = s_csamul_rca16_and8_12 ^ s_csamul_rca16_fa9_11_xor1;
  assign s_csamul_rca16_fa8_12_and0 = s_csamul_rca16_and8_12 & s_csamul_rca16_fa9_11_xor1;
  assign s_csamul_rca16_fa8_12_xor1 = s_csamul_rca16_fa8_12_xor0 ^ s_csamul_rca16_fa8_11_or0;
  assign s_csamul_rca16_fa8_12_and1 = s_csamul_rca16_fa8_12_xor0 & s_csamul_rca16_fa8_11_or0;
  assign s_csamul_rca16_fa8_12_or0 = s_csamul_rca16_fa8_12_and0 | s_csamul_rca16_fa8_12_and1;
  assign s_csamul_rca16_and9_12 = a[9] & b[12];
  assign s_csamul_rca16_fa9_12_xor0 = s_csamul_rca16_and9_12 ^ s_csamul_rca16_fa10_11_xor1;
  assign s_csamul_rca16_fa9_12_and0 = s_csamul_rca16_and9_12 & s_csamul_rca16_fa10_11_xor1;
  assign s_csamul_rca16_fa9_12_xor1 = s_csamul_rca16_fa9_12_xor0 ^ s_csamul_rca16_fa9_11_or0;
  assign s_csamul_rca16_fa9_12_and1 = s_csamul_rca16_fa9_12_xor0 & s_csamul_rca16_fa9_11_or0;
  assign s_csamul_rca16_fa9_12_or0 = s_csamul_rca16_fa9_12_and0 | s_csamul_rca16_fa9_12_and1;
  assign s_csamul_rca16_and10_12 = a[10] & b[12];
  assign s_csamul_rca16_fa10_12_xor0 = s_csamul_rca16_and10_12 ^ s_csamul_rca16_fa11_11_xor1;
  assign s_csamul_rca16_fa10_12_and0 = s_csamul_rca16_and10_12 & s_csamul_rca16_fa11_11_xor1;
  assign s_csamul_rca16_fa10_12_xor1 = s_csamul_rca16_fa10_12_xor0 ^ s_csamul_rca16_fa10_11_or0;
  assign s_csamul_rca16_fa10_12_and1 = s_csamul_rca16_fa10_12_xor0 & s_csamul_rca16_fa10_11_or0;
  assign s_csamul_rca16_fa10_12_or0 = s_csamul_rca16_fa10_12_and0 | s_csamul_rca16_fa10_12_and1;
  assign s_csamul_rca16_and11_12 = a[11] & b[12];
  assign s_csamul_rca16_fa11_12_xor0 = s_csamul_rca16_and11_12 ^ s_csamul_rca16_fa12_11_xor1;
  assign s_csamul_rca16_fa11_12_and0 = s_csamul_rca16_and11_12 & s_csamul_rca16_fa12_11_xor1;
  assign s_csamul_rca16_fa11_12_xor1 = s_csamul_rca16_fa11_12_xor0 ^ s_csamul_rca16_fa11_11_or0;
  assign s_csamul_rca16_fa11_12_and1 = s_csamul_rca16_fa11_12_xor0 & s_csamul_rca16_fa11_11_or0;
  assign s_csamul_rca16_fa11_12_or0 = s_csamul_rca16_fa11_12_and0 | s_csamul_rca16_fa11_12_and1;
  assign s_csamul_rca16_and12_12 = a[12] & b[12];
  assign s_csamul_rca16_fa12_12_xor0 = s_csamul_rca16_and12_12 ^ s_csamul_rca16_fa13_11_xor1;
  assign s_csamul_rca16_fa12_12_and0 = s_csamul_rca16_and12_12 & s_csamul_rca16_fa13_11_xor1;
  assign s_csamul_rca16_fa12_12_xor1 = s_csamul_rca16_fa12_12_xor0 ^ s_csamul_rca16_fa12_11_or0;
  assign s_csamul_rca16_fa12_12_and1 = s_csamul_rca16_fa12_12_xor0 & s_csamul_rca16_fa12_11_or0;
  assign s_csamul_rca16_fa12_12_or0 = s_csamul_rca16_fa12_12_and0 | s_csamul_rca16_fa12_12_and1;
  assign s_csamul_rca16_and13_12 = a[13] & b[12];
  assign s_csamul_rca16_fa13_12_xor0 = s_csamul_rca16_and13_12 ^ s_csamul_rca16_fa14_11_xor1;
  assign s_csamul_rca16_fa13_12_and0 = s_csamul_rca16_and13_12 & s_csamul_rca16_fa14_11_xor1;
  assign s_csamul_rca16_fa13_12_xor1 = s_csamul_rca16_fa13_12_xor0 ^ s_csamul_rca16_fa13_11_or0;
  assign s_csamul_rca16_fa13_12_and1 = s_csamul_rca16_fa13_12_xor0 & s_csamul_rca16_fa13_11_or0;
  assign s_csamul_rca16_fa13_12_or0 = s_csamul_rca16_fa13_12_and0 | s_csamul_rca16_fa13_12_and1;
  assign s_csamul_rca16_and14_12 = a[14] & b[12];
  assign s_csamul_rca16_fa14_12_xor0 = s_csamul_rca16_and14_12 ^ s_csamul_rca16_ha15_11_xor0;
  assign s_csamul_rca16_fa14_12_and0 = s_csamul_rca16_and14_12 & s_csamul_rca16_ha15_11_xor0;
  assign s_csamul_rca16_fa14_12_xor1 = s_csamul_rca16_fa14_12_xor0 ^ s_csamul_rca16_fa14_11_or0;
  assign s_csamul_rca16_fa14_12_and1 = s_csamul_rca16_fa14_12_xor0 & s_csamul_rca16_fa14_11_or0;
  assign s_csamul_rca16_fa14_12_or0 = s_csamul_rca16_fa14_12_and0 | s_csamul_rca16_fa14_12_and1;
  assign s_csamul_rca16_nand15_12 = ~(a[15] & b[12]);
  assign s_csamul_rca16_ha15_12_xor0 = s_csamul_rca16_nand15_12 ^ s_csamul_rca16_ha15_11_and0;
  assign s_csamul_rca16_ha15_12_and0 = s_csamul_rca16_nand15_12 & s_csamul_rca16_ha15_11_and0;
  assign s_csamul_rca16_and0_13 = a[0] & b[13];
  assign s_csamul_rca16_fa0_13_xor0 = s_csamul_rca16_and0_13 ^ s_csamul_rca16_fa1_12_xor1;
  assign s_csamul_rca16_fa0_13_and0 = s_csamul_rca16_and0_13 & s_csamul_rca16_fa1_12_xor1;
  assign s_csamul_rca16_fa0_13_xor1 = s_csamul_rca16_fa0_13_xor0 ^ s_csamul_rca16_fa0_12_or0;
  assign s_csamul_rca16_fa0_13_and1 = s_csamul_rca16_fa0_13_xor0 & s_csamul_rca16_fa0_12_or0;
  assign s_csamul_rca16_fa0_13_or0 = s_csamul_rca16_fa0_13_and0 | s_csamul_rca16_fa0_13_and1;
  assign s_csamul_rca16_and1_13 = a[1] & b[13];
  assign s_csamul_rca16_fa1_13_xor0 = s_csamul_rca16_and1_13 ^ s_csamul_rca16_fa2_12_xor1;
  assign s_csamul_rca16_fa1_13_and0 = s_csamul_rca16_and1_13 & s_csamul_rca16_fa2_12_xor1;
  assign s_csamul_rca16_fa1_13_xor1 = s_csamul_rca16_fa1_13_xor0 ^ s_csamul_rca16_fa1_12_or0;
  assign s_csamul_rca16_fa1_13_and1 = s_csamul_rca16_fa1_13_xor0 & s_csamul_rca16_fa1_12_or0;
  assign s_csamul_rca16_fa1_13_or0 = s_csamul_rca16_fa1_13_and0 | s_csamul_rca16_fa1_13_and1;
  assign s_csamul_rca16_and2_13 = a[2] & b[13];
  assign s_csamul_rca16_fa2_13_xor0 = s_csamul_rca16_and2_13 ^ s_csamul_rca16_fa3_12_xor1;
  assign s_csamul_rca16_fa2_13_and0 = s_csamul_rca16_and2_13 & s_csamul_rca16_fa3_12_xor1;
  assign s_csamul_rca16_fa2_13_xor1 = s_csamul_rca16_fa2_13_xor0 ^ s_csamul_rca16_fa2_12_or0;
  assign s_csamul_rca16_fa2_13_and1 = s_csamul_rca16_fa2_13_xor0 & s_csamul_rca16_fa2_12_or0;
  assign s_csamul_rca16_fa2_13_or0 = s_csamul_rca16_fa2_13_and0 | s_csamul_rca16_fa2_13_and1;
  assign s_csamul_rca16_and3_13 = a[3] & b[13];
  assign s_csamul_rca16_fa3_13_xor0 = s_csamul_rca16_and3_13 ^ s_csamul_rca16_fa4_12_xor1;
  assign s_csamul_rca16_fa3_13_and0 = s_csamul_rca16_and3_13 & s_csamul_rca16_fa4_12_xor1;
  assign s_csamul_rca16_fa3_13_xor1 = s_csamul_rca16_fa3_13_xor0 ^ s_csamul_rca16_fa3_12_or0;
  assign s_csamul_rca16_fa3_13_and1 = s_csamul_rca16_fa3_13_xor0 & s_csamul_rca16_fa3_12_or0;
  assign s_csamul_rca16_fa3_13_or0 = s_csamul_rca16_fa3_13_and0 | s_csamul_rca16_fa3_13_and1;
  assign s_csamul_rca16_and4_13 = a[4] & b[13];
  assign s_csamul_rca16_fa4_13_xor0 = s_csamul_rca16_and4_13 ^ s_csamul_rca16_fa5_12_xor1;
  assign s_csamul_rca16_fa4_13_and0 = s_csamul_rca16_and4_13 & s_csamul_rca16_fa5_12_xor1;
  assign s_csamul_rca16_fa4_13_xor1 = s_csamul_rca16_fa4_13_xor0 ^ s_csamul_rca16_fa4_12_or0;
  assign s_csamul_rca16_fa4_13_and1 = s_csamul_rca16_fa4_13_xor0 & s_csamul_rca16_fa4_12_or0;
  assign s_csamul_rca16_fa4_13_or0 = s_csamul_rca16_fa4_13_and0 | s_csamul_rca16_fa4_13_and1;
  assign s_csamul_rca16_and5_13 = a[5] & b[13];
  assign s_csamul_rca16_fa5_13_xor0 = s_csamul_rca16_and5_13 ^ s_csamul_rca16_fa6_12_xor1;
  assign s_csamul_rca16_fa5_13_and0 = s_csamul_rca16_and5_13 & s_csamul_rca16_fa6_12_xor1;
  assign s_csamul_rca16_fa5_13_xor1 = s_csamul_rca16_fa5_13_xor0 ^ s_csamul_rca16_fa5_12_or0;
  assign s_csamul_rca16_fa5_13_and1 = s_csamul_rca16_fa5_13_xor0 & s_csamul_rca16_fa5_12_or0;
  assign s_csamul_rca16_fa5_13_or0 = s_csamul_rca16_fa5_13_and0 | s_csamul_rca16_fa5_13_and1;
  assign s_csamul_rca16_and6_13 = a[6] & b[13];
  assign s_csamul_rca16_fa6_13_xor0 = s_csamul_rca16_and6_13 ^ s_csamul_rca16_fa7_12_xor1;
  assign s_csamul_rca16_fa6_13_and0 = s_csamul_rca16_and6_13 & s_csamul_rca16_fa7_12_xor1;
  assign s_csamul_rca16_fa6_13_xor1 = s_csamul_rca16_fa6_13_xor0 ^ s_csamul_rca16_fa6_12_or0;
  assign s_csamul_rca16_fa6_13_and1 = s_csamul_rca16_fa6_13_xor0 & s_csamul_rca16_fa6_12_or0;
  assign s_csamul_rca16_fa6_13_or0 = s_csamul_rca16_fa6_13_and0 | s_csamul_rca16_fa6_13_and1;
  assign s_csamul_rca16_and7_13 = a[7] & b[13];
  assign s_csamul_rca16_fa7_13_xor0 = s_csamul_rca16_and7_13 ^ s_csamul_rca16_fa8_12_xor1;
  assign s_csamul_rca16_fa7_13_and0 = s_csamul_rca16_and7_13 & s_csamul_rca16_fa8_12_xor1;
  assign s_csamul_rca16_fa7_13_xor1 = s_csamul_rca16_fa7_13_xor0 ^ s_csamul_rca16_fa7_12_or0;
  assign s_csamul_rca16_fa7_13_and1 = s_csamul_rca16_fa7_13_xor0 & s_csamul_rca16_fa7_12_or0;
  assign s_csamul_rca16_fa7_13_or0 = s_csamul_rca16_fa7_13_and0 | s_csamul_rca16_fa7_13_and1;
  assign s_csamul_rca16_and8_13 = a[8] & b[13];
  assign s_csamul_rca16_fa8_13_xor0 = s_csamul_rca16_and8_13 ^ s_csamul_rca16_fa9_12_xor1;
  assign s_csamul_rca16_fa8_13_and0 = s_csamul_rca16_and8_13 & s_csamul_rca16_fa9_12_xor1;
  assign s_csamul_rca16_fa8_13_xor1 = s_csamul_rca16_fa8_13_xor0 ^ s_csamul_rca16_fa8_12_or0;
  assign s_csamul_rca16_fa8_13_and1 = s_csamul_rca16_fa8_13_xor0 & s_csamul_rca16_fa8_12_or0;
  assign s_csamul_rca16_fa8_13_or0 = s_csamul_rca16_fa8_13_and0 | s_csamul_rca16_fa8_13_and1;
  assign s_csamul_rca16_and9_13 = a[9] & b[13];
  assign s_csamul_rca16_fa9_13_xor0 = s_csamul_rca16_and9_13 ^ s_csamul_rca16_fa10_12_xor1;
  assign s_csamul_rca16_fa9_13_and0 = s_csamul_rca16_and9_13 & s_csamul_rca16_fa10_12_xor1;
  assign s_csamul_rca16_fa9_13_xor1 = s_csamul_rca16_fa9_13_xor0 ^ s_csamul_rca16_fa9_12_or0;
  assign s_csamul_rca16_fa9_13_and1 = s_csamul_rca16_fa9_13_xor0 & s_csamul_rca16_fa9_12_or0;
  assign s_csamul_rca16_fa9_13_or0 = s_csamul_rca16_fa9_13_and0 | s_csamul_rca16_fa9_13_and1;
  assign s_csamul_rca16_and10_13 = a[10] & b[13];
  assign s_csamul_rca16_fa10_13_xor0 = s_csamul_rca16_and10_13 ^ s_csamul_rca16_fa11_12_xor1;
  assign s_csamul_rca16_fa10_13_and0 = s_csamul_rca16_and10_13 & s_csamul_rca16_fa11_12_xor1;
  assign s_csamul_rca16_fa10_13_xor1 = s_csamul_rca16_fa10_13_xor0 ^ s_csamul_rca16_fa10_12_or0;
  assign s_csamul_rca16_fa10_13_and1 = s_csamul_rca16_fa10_13_xor0 & s_csamul_rca16_fa10_12_or0;
  assign s_csamul_rca16_fa10_13_or0 = s_csamul_rca16_fa10_13_and0 | s_csamul_rca16_fa10_13_and1;
  assign s_csamul_rca16_and11_13 = a[11] & b[13];
  assign s_csamul_rca16_fa11_13_xor0 = s_csamul_rca16_and11_13 ^ s_csamul_rca16_fa12_12_xor1;
  assign s_csamul_rca16_fa11_13_and0 = s_csamul_rca16_and11_13 & s_csamul_rca16_fa12_12_xor1;
  assign s_csamul_rca16_fa11_13_xor1 = s_csamul_rca16_fa11_13_xor0 ^ s_csamul_rca16_fa11_12_or0;
  assign s_csamul_rca16_fa11_13_and1 = s_csamul_rca16_fa11_13_xor0 & s_csamul_rca16_fa11_12_or0;
  assign s_csamul_rca16_fa11_13_or0 = s_csamul_rca16_fa11_13_and0 | s_csamul_rca16_fa11_13_and1;
  assign s_csamul_rca16_and12_13 = a[12] & b[13];
  assign s_csamul_rca16_fa12_13_xor0 = s_csamul_rca16_and12_13 ^ s_csamul_rca16_fa13_12_xor1;
  assign s_csamul_rca16_fa12_13_and0 = s_csamul_rca16_and12_13 & s_csamul_rca16_fa13_12_xor1;
  assign s_csamul_rca16_fa12_13_xor1 = s_csamul_rca16_fa12_13_xor0 ^ s_csamul_rca16_fa12_12_or0;
  assign s_csamul_rca16_fa12_13_and1 = s_csamul_rca16_fa12_13_xor0 & s_csamul_rca16_fa12_12_or0;
  assign s_csamul_rca16_fa12_13_or0 = s_csamul_rca16_fa12_13_and0 | s_csamul_rca16_fa12_13_and1;
  assign s_csamul_rca16_and13_13 = a[13] & b[13];
  assign s_csamul_rca16_fa13_13_xor0 = s_csamul_rca16_and13_13 ^ s_csamul_rca16_fa14_12_xor1;
  assign s_csamul_rca16_fa13_13_and0 = s_csamul_rca16_and13_13 & s_csamul_rca16_fa14_12_xor1;
  assign s_csamul_rca16_fa13_13_xor1 = s_csamul_rca16_fa13_13_xor0 ^ s_csamul_rca16_fa13_12_or0;
  assign s_csamul_rca16_fa13_13_and1 = s_csamul_rca16_fa13_13_xor0 & s_csamul_rca16_fa13_12_or0;
  assign s_csamul_rca16_fa13_13_or0 = s_csamul_rca16_fa13_13_and0 | s_csamul_rca16_fa13_13_and1;
  assign s_csamul_rca16_and14_13 = a[14] & b[13];
  assign s_csamul_rca16_fa14_13_xor0 = s_csamul_rca16_and14_13 ^ s_csamul_rca16_ha15_12_xor0;
  assign s_csamul_rca16_fa14_13_and0 = s_csamul_rca16_and14_13 & s_csamul_rca16_ha15_12_xor0;
  assign s_csamul_rca16_fa14_13_xor1 = s_csamul_rca16_fa14_13_xor0 ^ s_csamul_rca16_fa14_12_or0;
  assign s_csamul_rca16_fa14_13_and1 = s_csamul_rca16_fa14_13_xor0 & s_csamul_rca16_fa14_12_or0;
  assign s_csamul_rca16_fa14_13_or0 = s_csamul_rca16_fa14_13_and0 | s_csamul_rca16_fa14_13_and1;
  assign s_csamul_rca16_nand15_13 = ~(a[15] & b[13]);
  assign s_csamul_rca16_ha15_13_xor0 = s_csamul_rca16_nand15_13 ^ s_csamul_rca16_ha15_12_and0;
  assign s_csamul_rca16_ha15_13_and0 = s_csamul_rca16_nand15_13 & s_csamul_rca16_ha15_12_and0;
  assign s_csamul_rca16_and0_14 = a[0] & b[14];
  assign s_csamul_rca16_fa0_14_xor0 = s_csamul_rca16_and0_14 ^ s_csamul_rca16_fa1_13_xor1;
  assign s_csamul_rca16_fa0_14_and0 = s_csamul_rca16_and0_14 & s_csamul_rca16_fa1_13_xor1;
  assign s_csamul_rca16_fa0_14_xor1 = s_csamul_rca16_fa0_14_xor0 ^ s_csamul_rca16_fa0_13_or0;
  assign s_csamul_rca16_fa0_14_and1 = s_csamul_rca16_fa0_14_xor0 & s_csamul_rca16_fa0_13_or0;
  assign s_csamul_rca16_fa0_14_or0 = s_csamul_rca16_fa0_14_and0 | s_csamul_rca16_fa0_14_and1;
  assign s_csamul_rca16_and1_14 = a[1] & b[14];
  assign s_csamul_rca16_fa1_14_xor0 = s_csamul_rca16_and1_14 ^ s_csamul_rca16_fa2_13_xor1;
  assign s_csamul_rca16_fa1_14_and0 = s_csamul_rca16_and1_14 & s_csamul_rca16_fa2_13_xor1;
  assign s_csamul_rca16_fa1_14_xor1 = s_csamul_rca16_fa1_14_xor0 ^ s_csamul_rca16_fa1_13_or0;
  assign s_csamul_rca16_fa1_14_and1 = s_csamul_rca16_fa1_14_xor0 & s_csamul_rca16_fa1_13_or0;
  assign s_csamul_rca16_fa1_14_or0 = s_csamul_rca16_fa1_14_and0 | s_csamul_rca16_fa1_14_and1;
  assign s_csamul_rca16_and2_14 = a[2] & b[14];
  assign s_csamul_rca16_fa2_14_xor0 = s_csamul_rca16_and2_14 ^ s_csamul_rca16_fa3_13_xor1;
  assign s_csamul_rca16_fa2_14_and0 = s_csamul_rca16_and2_14 & s_csamul_rca16_fa3_13_xor1;
  assign s_csamul_rca16_fa2_14_xor1 = s_csamul_rca16_fa2_14_xor0 ^ s_csamul_rca16_fa2_13_or0;
  assign s_csamul_rca16_fa2_14_and1 = s_csamul_rca16_fa2_14_xor0 & s_csamul_rca16_fa2_13_or0;
  assign s_csamul_rca16_fa2_14_or0 = s_csamul_rca16_fa2_14_and0 | s_csamul_rca16_fa2_14_and1;
  assign s_csamul_rca16_and3_14 = a[3] & b[14];
  assign s_csamul_rca16_fa3_14_xor0 = s_csamul_rca16_and3_14 ^ s_csamul_rca16_fa4_13_xor1;
  assign s_csamul_rca16_fa3_14_and0 = s_csamul_rca16_and3_14 & s_csamul_rca16_fa4_13_xor1;
  assign s_csamul_rca16_fa3_14_xor1 = s_csamul_rca16_fa3_14_xor0 ^ s_csamul_rca16_fa3_13_or0;
  assign s_csamul_rca16_fa3_14_and1 = s_csamul_rca16_fa3_14_xor0 & s_csamul_rca16_fa3_13_or0;
  assign s_csamul_rca16_fa3_14_or0 = s_csamul_rca16_fa3_14_and0 | s_csamul_rca16_fa3_14_and1;
  assign s_csamul_rca16_and4_14 = a[4] & b[14];
  assign s_csamul_rca16_fa4_14_xor0 = s_csamul_rca16_and4_14 ^ s_csamul_rca16_fa5_13_xor1;
  assign s_csamul_rca16_fa4_14_and0 = s_csamul_rca16_and4_14 & s_csamul_rca16_fa5_13_xor1;
  assign s_csamul_rca16_fa4_14_xor1 = s_csamul_rca16_fa4_14_xor0 ^ s_csamul_rca16_fa4_13_or0;
  assign s_csamul_rca16_fa4_14_and1 = s_csamul_rca16_fa4_14_xor0 & s_csamul_rca16_fa4_13_or0;
  assign s_csamul_rca16_fa4_14_or0 = s_csamul_rca16_fa4_14_and0 | s_csamul_rca16_fa4_14_and1;
  assign s_csamul_rca16_and5_14 = a[5] & b[14];
  assign s_csamul_rca16_fa5_14_xor0 = s_csamul_rca16_and5_14 ^ s_csamul_rca16_fa6_13_xor1;
  assign s_csamul_rca16_fa5_14_and0 = s_csamul_rca16_and5_14 & s_csamul_rca16_fa6_13_xor1;
  assign s_csamul_rca16_fa5_14_xor1 = s_csamul_rca16_fa5_14_xor0 ^ s_csamul_rca16_fa5_13_or0;
  assign s_csamul_rca16_fa5_14_and1 = s_csamul_rca16_fa5_14_xor0 & s_csamul_rca16_fa5_13_or0;
  assign s_csamul_rca16_fa5_14_or0 = s_csamul_rca16_fa5_14_and0 | s_csamul_rca16_fa5_14_and1;
  assign s_csamul_rca16_and6_14 = a[6] & b[14];
  assign s_csamul_rca16_fa6_14_xor0 = s_csamul_rca16_and6_14 ^ s_csamul_rca16_fa7_13_xor1;
  assign s_csamul_rca16_fa6_14_and0 = s_csamul_rca16_and6_14 & s_csamul_rca16_fa7_13_xor1;
  assign s_csamul_rca16_fa6_14_xor1 = s_csamul_rca16_fa6_14_xor0 ^ s_csamul_rca16_fa6_13_or0;
  assign s_csamul_rca16_fa6_14_and1 = s_csamul_rca16_fa6_14_xor0 & s_csamul_rca16_fa6_13_or0;
  assign s_csamul_rca16_fa6_14_or0 = s_csamul_rca16_fa6_14_and0 | s_csamul_rca16_fa6_14_and1;
  assign s_csamul_rca16_and7_14 = a[7] & b[14];
  assign s_csamul_rca16_fa7_14_xor0 = s_csamul_rca16_and7_14 ^ s_csamul_rca16_fa8_13_xor1;
  assign s_csamul_rca16_fa7_14_and0 = s_csamul_rca16_and7_14 & s_csamul_rca16_fa8_13_xor1;
  assign s_csamul_rca16_fa7_14_xor1 = s_csamul_rca16_fa7_14_xor0 ^ s_csamul_rca16_fa7_13_or0;
  assign s_csamul_rca16_fa7_14_and1 = s_csamul_rca16_fa7_14_xor0 & s_csamul_rca16_fa7_13_or0;
  assign s_csamul_rca16_fa7_14_or0 = s_csamul_rca16_fa7_14_and0 | s_csamul_rca16_fa7_14_and1;
  assign s_csamul_rca16_and8_14 = a[8] & b[14];
  assign s_csamul_rca16_fa8_14_xor0 = s_csamul_rca16_and8_14 ^ s_csamul_rca16_fa9_13_xor1;
  assign s_csamul_rca16_fa8_14_and0 = s_csamul_rca16_and8_14 & s_csamul_rca16_fa9_13_xor1;
  assign s_csamul_rca16_fa8_14_xor1 = s_csamul_rca16_fa8_14_xor0 ^ s_csamul_rca16_fa8_13_or0;
  assign s_csamul_rca16_fa8_14_and1 = s_csamul_rca16_fa8_14_xor0 & s_csamul_rca16_fa8_13_or0;
  assign s_csamul_rca16_fa8_14_or0 = s_csamul_rca16_fa8_14_and0 | s_csamul_rca16_fa8_14_and1;
  assign s_csamul_rca16_and9_14 = a[9] & b[14];
  assign s_csamul_rca16_fa9_14_xor0 = s_csamul_rca16_and9_14 ^ s_csamul_rca16_fa10_13_xor1;
  assign s_csamul_rca16_fa9_14_and0 = s_csamul_rca16_and9_14 & s_csamul_rca16_fa10_13_xor1;
  assign s_csamul_rca16_fa9_14_xor1 = s_csamul_rca16_fa9_14_xor0 ^ s_csamul_rca16_fa9_13_or0;
  assign s_csamul_rca16_fa9_14_and1 = s_csamul_rca16_fa9_14_xor0 & s_csamul_rca16_fa9_13_or0;
  assign s_csamul_rca16_fa9_14_or0 = s_csamul_rca16_fa9_14_and0 | s_csamul_rca16_fa9_14_and1;
  assign s_csamul_rca16_and10_14 = a[10] & b[14];
  assign s_csamul_rca16_fa10_14_xor0 = s_csamul_rca16_and10_14 ^ s_csamul_rca16_fa11_13_xor1;
  assign s_csamul_rca16_fa10_14_and0 = s_csamul_rca16_and10_14 & s_csamul_rca16_fa11_13_xor1;
  assign s_csamul_rca16_fa10_14_xor1 = s_csamul_rca16_fa10_14_xor0 ^ s_csamul_rca16_fa10_13_or0;
  assign s_csamul_rca16_fa10_14_and1 = s_csamul_rca16_fa10_14_xor0 & s_csamul_rca16_fa10_13_or0;
  assign s_csamul_rca16_fa10_14_or0 = s_csamul_rca16_fa10_14_and0 | s_csamul_rca16_fa10_14_and1;
  assign s_csamul_rca16_and11_14 = a[11] & b[14];
  assign s_csamul_rca16_fa11_14_xor0 = s_csamul_rca16_and11_14 ^ s_csamul_rca16_fa12_13_xor1;
  assign s_csamul_rca16_fa11_14_and0 = s_csamul_rca16_and11_14 & s_csamul_rca16_fa12_13_xor1;
  assign s_csamul_rca16_fa11_14_xor1 = s_csamul_rca16_fa11_14_xor0 ^ s_csamul_rca16_fa11_13_or0;
  assign s_csamul_rca16_fa11_14_and1 = s_csamul_rca16_fa11_14_xor0 & s_csamul_rca16_fa11_13_or0;
  assign s_csamul_rca16_fa11_14_or0 = s_csamul_rca16_fa11_14_and0 | s_csamul_rca16_fa11_14_and1;
  assign s_csamul_rca16_and12_14 = a[12] & b[14];
  assign s_csamul_rca16_fa12_14_xor0 = s_csamul_rca16_and12_14 ^ s_csamul_rca16_fa13_13_xor1;
  assign s_csamul_rca16_fa12_14_and0 = s_csamul_rca16_and12_14 & s_csamul_rca16_fa13_13_xor1;
  assign s_csamul_rca16_fa12_14_xor1 = s_csamul_rca16_fa12_14_xor0 ^ s_csamul_rca16_fa12_13_or0;
  assign s_csamul_rca16_fa12_14_and1 = s_csamul_rca16_fa12_14_xor0 & s_csamul_rca16_fa12_13_or0;
  assign s_csamul_rca16_fa12_14_or0 = s_csamul_rca16_fa12_14_and0 | s_csamul_rca16_fa12_14_and1;
  assign s_csamul_rca16_and13_14 = a[13] & b[14];
  assign s_csamul_rca16_fa13_14_xor0 = s_csamul_rca16_and13_14 ^ s_csamul_rca16_fa14_13_xor1;
  assign s_csamul_rca16_fa13_14_and0 = s_csamul_rca16_and13_14 & s_csamul_rca16_fa14_13_xor1;
  assign s_csamul_rca16_fa13_14_xor1 = s_csamul_rca16_fa13_14_xor0 ^ s_csamul_rca16_fa13_13_or0;
  assign s_csamul_rca16_fa13_14_and1 = s_csamul_rca16_fa13_14_xor0 & s_csamul_rca16_fa13_13_or0;
  assign s_csamul_rca16_fa13_14_or0 = s_csamul_rca16_fa13_14_and0 | s_csamul_rca16_fa13_14_and1;
  assign s_csamul_rca16_and14_14 = a[14] & b[14];
  assign s_csamul_rca16_fa14_14_xor0 = s_csamul_rca16_and14_14 ^ s_csamul_rca16_ha15_13_xor0;
  assign s_csamul_rca16_fa14_14_and0 = s_csamul_rca16_and14_14 & s_csamul_rca16_ha15_13_xor0;
  assign s_csamul_rca16_fa14_14_xor1 = s_csamul_rca16_fa14_14_xor0 ^ s_csamul_rca16_fa14_13_or0;
  assign s_csamul_rca16_fa14_14_and1 = s_csamul_rca16_fa14_14_xor0 & s_csamul_rca16_fa14_13_or0;
  assign s_csamul_rca16_fa14_14_or0 = s_csamul_rca16_fa14_14_and0 | s_csamul_rca16_fa14_14_and1;
  assign s_csamul_rca16_nand15_14 = ~(a[15] & b[14]);
  assign s_csamul_rca16_ha15_14_xor0 = s_csamul_rca16_nand15_14 ^ s_csamul_rca16_ha15_13_and0;
  assign s_csamul_rca16_ha15_14_and0 = s_csamul_rca16_nand15_14 & s_csamul_rca16_ha15_13_and0;
  assign s_csamul_rca16_nand0_15 = ~(a[0] & b[15]);
  assign s_csamul_rca16_fa0_15_xor0 = s_csamul_rca16_nand0_15 ^ s_csamul_rca16_fa1_14_xor1;
  assign s_csamul_rca16_fa0_15_and0 = s_csamul_rca16_nand0_15 & s_csamul_rca16_fa1_14_xor1;
  assign s_csamul_rca16_fa0_15_xor1 = s_csamul_rca16_fa0_15_xor0 ^ s_csamul_rca16_fa0_14_or0;
  assign s_csamul_rca16_fa0_15_and1 = s_csamul_rca16_fa0_15_xor0 & s_csamul_rca16_fa0_14_or0;
  assign s_csamul_rca16_fa0_15_or0 = s_csamul_rca16_fa0_15_and0 | s_csamul_rca16_fa0_15_and1;
  assign s_csamul_rca16_nand1_15 = ~(a[1] & b[15]);
  assign s_csamul_rca16_fa1_15_xor0 = s_csamul_rca16_nand1_15 ^ s_csamul_rca16_fa2_14_xor1;
  assign s_csamul_rca16_fa1_15_and0 = s_csamul_rca16_nand1_15 & s_csamul_rca16_fa2_14_xor1;
  assign s_csamul_rca16_fa1_15_xor1 = s_csamul_rca16_fa1_15_xor0 ^ s_csamul_rca16_fa1_14_or0;
  assign s_csamul_rca16_fa1_15_and1 = s_csamul_rca16_fa1_15_xor0 & s_csamul_rca16_fa1_14_or0;
  assign s_csamul_rca16_fa1_15_or0 = s_csamul_rca16_fa1_15_and0 | s_csamul_rca16_fa1_15_and1;
  assign s_csamul_rca16_nand2_15 = ~(a[2] & b[15]);
  assign s_csamul_rca16_fa2_15_xor0 = s_csamul_rca16_nand2_15 ^ s_csamul_rca16_fa3_14_xor1;
  assign s_csamul_rca16_fa2_15_and0 = s_csamul_rca16_nand2_15 & s_csamul_rca16_fa3_14_xor1;
  assign s_csamul_rca16_fa2_15_xor1 = s_csamul_rca16_fa2_15_xor0 ^ s_csamul_rca16_fa2_14_or0;
  assign s_csamul_rca16_fa2_15_and1 = s_csamul_rca16_fa2_15_xor0 & s_csamul_rca16_fa2_14_or0;
  assign s_csamul_rca16_fa2_15_or0 = s_csamul_rca16_fa2_15_and0 | s_csamul_rca16_fa2_15_and1;
  assign s_csamul_rca16_nand3_15 = ~(a[3] & b[15]);
  assign s_csamul_rca16_fa3_15_xor0 = s_csamul_rca16_nand3_15 ^ s_csamul_rca16_fa4_14_xor1;
  assign s_csamul_rca16_fa3_15_and0 = s_csamul_rca16_nand3_15 & s_csamul_rca16_fa4_14_xor1;
  assign s_csamul_rca16_fa3_15_xor1 = s_csamul_rca16_fa3_15_xor0 ^ s_csamul_rca16_fa3_14_or0;
  assign s_csamul_rca16_fa3_15_and1 = s_csamul_rca16_fa3_15_xor0 & s_csamul_rca16_fa3_14_or0;
  assign s_csamul_rca16_fa3_15_or0 = s_csamul_rca16_fa3_15_and0 | s_csamul_rca16_fa3_15_and1;
  assign s_csamul_rca16_nand4_15 = ~(a[4] & b[15]);
  assign s_csamul_rca16_fa4_15_xor0 = s_csamul_rca16_nand4_15 ^ s_csamul_rca16_fa5_14_xor1;
  assign s_csamul_rca16_fa4_15_and0 = s_csamul_rca16_nand4_15 & s_csamul_rca16_fa5_14_xor1;
  assign s_csamul_rca16_fa4_15_xor1 = s_csamul_rca16_fa4_15_xor0 ^ s_csamul_rca16_fa4_14_or0;
  assign s_csamul_rca16_fa4_15_and1 = s_csamul_rca16_fa4_15_xor0 & s_csamul_rca16_fa4_14_or0;
  assign s_csamul_rca16_fa4_15_or0 = s_csamul_rca16_fa4_15_and0 | s_csamul_rca16_fa4_15_and1;
  assign s_csamul_rca16_nand5_15 = ~(a[5] & b[15]);
  assign s_csamul_rca16_fa5_15_xor0 = s_csamul_rca16_nand5_15 ^ s_csamul_rca16_fa6_14_xor1;
  assign s_csamul_rca16_fa5_15_and0 = s_csamul_rca16_nand5_15 & s_csamul_rca16_fa6_14_xor1;
  assign s_csamul_rca16_fa5_15_xor1 = s_csamul_rca16_fa5_15_xor0 ^ s_csamul_rca16_fa5_14_or0;
  assign s_csamul_rca16_fa5_15_and1 = s_csamul_rca16_fa5_15_xor0 & s_csamul_rca16_fa5_14_or0;
  assign s_csamul_rca16_fa5_15_or0 = s_csamul_rca16_fa5_15_and0 | s_csamul_rca16_fa5_15_and1;
  assign s_csamul_rca16_nand6_15 = ~(a[6] & b[15]);
  assign s_csamul_rca16_fa6_15_xor0 = s_csamul_rca16_nand6_15 ^ s_csamul_rca16_fa7_14_xor1;
  assign s_csamul_rca16_fa6_15_and0 = s_csamul_rca16_nand6_15 & s_csamul_rca16_fa7_14_xor1;
  assign s_csamul_rca16_fa6_15_xor1 = s_csamul_rca16_fa6_15_xor0 ^ s_csamul_rca16_fa6_14_or0;
  assign s_csamul_rca16_fa6_15_and1 = s_csamul_rca16_fa6_15_xor0 & s_csamul_rca16_fa6_14_or0;
  assign s_csamul_rca16_fa6_15_or0 = s_csamul_rca16_fa6_15_and0 | s_csamul_rca16_fa6_15_and1;
  assign s_csamul_rca16_nand7_15 = ~(a[7] & b[15]);
  assign s_csamul_rca16_fa7_15_xor0 = s_csamul_rca16_nand7_15 ^ s_csamul_rca16_fa8_14_xor1;
  assign s_csamul_rca16_fa7_15_and0 = s_csamul_rca16_nand7_15 & s_csamul_rca16_fa8_14_xor1;
  assign s_csamul_rca16_fa7_15_xor1 = s_csamul_rca16_fa7_15_xor0 ^ s_csamul_rca16_fa7_14_or0;
  assign s_csamul_rca16_fa7_15_and1 = s_csamul_rca16_fa7_15_xor0 & s_csamul_rca16_fa7_14_or0;
  assign s_csamul_rca16_fa7_15_or0 = s_csamul_rca16_fa7_15_and0 | s_csamul_rca16_fa7_15_and1;
  assign s_csamul_rca16_nand8_15 = ~(a[8] & b[15]);
  assign s_csamul_rca16_fa8_15_xor0 = s_csamul_rca16_nand8_15 ^ s_csamul_rca16_fa9_14_xor1;
  assign s_csamul_rca16_fa8_15_and0 = s_csamul_rca16_nand8_15 & s_csamul_rca16_fa9_14_xor1;
  assign s_csamul_rca16_fa8_15_xor1 = s_csamul_rca16_fa8_15_xor0 ^ s_csamul_rca16_fa8_14_or0;
  assign s_csamul_rca16_fa8_15_and1 = s_csamul_rca16_fa8_15_xor0 & s_csamul_rca16_fa8_14_or0;
  assign s_csamul_rca16_fa8_15_or0 = s_csamul_rca16_fa8_15_and0 | s_csamul_rca16_fa8_15_and1;
  assign s_csamul_rca16_nand9_15 = ~(a[9] & b[15]);
  assign s_csamul_rca16_fa9_15_xor0 = s_csamul_rca16_nand9_15 ^ s_csamul_rca16_fa10_14_xor1;
  assign s_csamul_rca16_fa9_15_and0 = s_csamul_rca16_nand9_15 & s_csamul_rca16_fa10_14_xor1;
  assign s_csamul_rca16_fa9_15_xor1 = s_csamul_rca16_fa9_15_xor0 ^ s_csamul_rca16_fa9_14_or0;
  assign s_csamul_rca16_fa9_15_and1 = s_csamul_rca16_fa9_15_xor0 & s_csamul_rca16_fa9_14_or0;
  assign s_csamul_rca16_fa9_15_or0 = s_csamul_rca16_fa9_15_and0 | s_csamul_rca16_fa9_15_and1;
  assign s_csamul_rca16_nand10_15 = ~(a[10] & b[15]);
  assign s_csamul_rca16_fa10_15_xor0 = s_csamul_rca16_nand10_15 ^ s_csamul_rca16_fa11_14_xor1;
  assign s_csamul_rca16_fa10_15_and0 = s_csamul_rca16_nand10_15 & s_csamul_rca16_fa11_14_xor1;
  assign s_csamul_rca16_fa10_15_xor1 = s_csamul_rca16_fa10_15_xor0 ^ s_csamul_rca16_fa10_14_or0;
  assign s_csamul_rca16_fa10_15_and1 = s_csamul_rca16_fa10_15_xor0 & s_csamul_rca16_fa10_14_or0;
  assign s_csamul_rca16_fa10_15_or0 = s_csamul_rca16_fa10_15_and0 | s_csamul_rca16_fa10_15_and1;
  assign s_csamul_rca16_nand11_15 = ~(a[11] & b[15]);
  assign s_csamul_rca16_fa11_15_xor0 = s_csamul_rca16_nand11_15 ^ s_csamul_rca16_fa12_14_xor1;
  assign s_csamul_rca16_fa11_15_and0 = s_csamul_rca16_nand11_15 & s_csamul_rca16_fa12_14_xor1;
  assign s_csamul_rca16_fa11_15_xor1 = s_csamul_rca16_fa11_15_xor0 ^ s_csamul_rca16_fa11_14_or0;
  assign s_csamul_rca16_fa11_15_and1 = s_csamul_rca16_fa11_15_xor0 & s_csamul_rca16_fa11_14_or0;
  assign s_csamul_rca16_fa11_15_or0 = s_csamul_rca16_fa11_15_and0 | s_csamul_rca16_fa11_15_and1;
  assign s_csamul_rca16_nand12_15 = ~(a[12] & b[15]);
  assign s_csamul_rca16_fa12_15_xor0 = s_csamul_rca16_nand12_15 ^ s_csamul_rca16_fa13_14_xor1;
  assign s_csamul_rca16_fa12_15_and0 = s_csamul_rca16_nand12_15 & s_csamul_rca16_fa13_14_xor1;
  assign s_csamul_rca16_fa12_15_xor1 = s_csamul_rca16_fa12_15_xor0 ^ s_csamul_rca16_fa12_14_or0;
  assign s_csamul_rca16_fa12_15_and1 = s_csamul_rca16_fa12_15_xor0 & s_csamul_rca16_fa12_14_or0;
  assign s_csamul_rca16_fa12_15_or0 = s_csamul_rca16_fa12_15_and0 | s_csamul_rca16_fa12_15_and1;
  assign s_csamul_rca16_nand13_15 = ~(a[13] & b[15]);
  assign s_csamul_rca16_fa13_15_xor0 = s_csamul_rca16_nand13_15 ^ s_csamul_rca16_fa14_14_xor1;
  assign s_csamul_rca16_fa13_15_and0 = s_csamul_rca16_nand13_15 & s_csamul_rca16_fa14_14_xor1;
  assign s_csamul_rca16_fa13_15_xor1 = s_csamul_rca16_fa13_15_xor0 ^ s_csamul_rca16_fa13_14_or0;
  assign s_csamul_rca16_fa13_15_and1 = s_csamul_rca16_fa13_15_xor0 & s_csamul_rca16_fa13_14_or0;
  assign s_csamul_rca16_fa13_15_or0 = s_csamul_rca16_fa13_15_and0 | s_csamul_rca16_fa13_15_and1;
  assign s_csamul_rca16_nand14_15 = ~(a[14] & b[15]);
  assign s_csamul_rca16_fa14_15_xor0 = s_csamul_rca16_nand14_15 ^ s_csamul_rca16_ha15_14_xor0;
  assign s_csamul_rca16_fa14_15_and0 = s_csamul_rca16_nand14_15 & s_csamul_rca16_ha15_14_xor0;
  assign s_csamul_rca16_fa14_15_xor1 = s_csamul_rca16_fa14_15_xor0 ^ s_csamul_rca16_fa14_14_or0;
  assign s_csamul_rca16_fa14_15_and1 = s_csamul_rca16_fa14_15_xor0 & s_csamul_rca16_fa14_14_or0;
  assign s_csamul_rca16_fa14_15_or0 = s_csamul_rca16_fa14_15_and0 | s_csamul_rca16_fa14_15_and1;
  assign s_csamul_rca16_and15_15 = a[15] & b[15];
  assign s_csamul_rca16_ha15_15_xor0 = s_csamul_rca16_and15_15 ^ s_csamul_rca16_ha15_14_and0;
  assign s_csamul_rca16_ha15_15_and0 = s_csamul_rca16_and15_15 & s_csamul_rca16_ha15_14_and0;
  assign s_csamul_rca16_u_rca16_ha_xor0 = s_csamul_rca16_fa1_15_xor1 ^ s_csamul_rca16_fa0_15_or0;
  assign s_csamul_rca16_u_rca16_ha_and0 = s_csamul_rca16_fa1_15_xor1 & s_csamul_rca16_fa0_15_or0;
  assign s_csamul_rca16_u_rca16_fa1_xor0 = s_csamul_rca16_fa2_15_xor1 ^ s_csamul_rca16_fa1_15_or0;
  assign s_csamul_rca16_u_rca16_fa1_and0 = s_csamul_rca16_fa2_15_xor1 & s_csamul_rca16_fa1_15_or0;
  assign s_csamul_rca16_u_rca16_fa1_xor1 = s_csamul_rca16_u_rca16_fa1_xor0 ^ s_csamul_rca16_u_rca16_ha_and0;
  assign s_csamul_rca16_u_rca16_fa1_and1 = s_csamul_rca16_u_rca16_fa1_xor0 & s_csamul_rca16_u_rca16_ha_and0;
  assign s_csamul_rca16_u_rca16_fa1_or0 = s_csamul_rca16_u_rca16_fa1_and0 | s_csamul_rca16_u_rca16_fa1_and1;
  assign s_csamul_rca16_u_rca16_fa2_xor0 = s_csamul_rca16_fa3_15_xor1 ^ s_csamul_rca16_fa2_15_or0;
  assign s_csamul_rca16_u_rca16_fa2_and0 = s_csamul_rca16_fa3_15_xor1 & s_csamul_rca16_fa2_15_or0;
  assign s_csamul_rca16_u_rca16_fa2_xor1 = s_csamul_rca16_u_rca16_fa2_xor0 ^ s_csamul_rca16_u_rca16_fa1_or0;
  assign s_csamul_rca16_u_rca16_fa2_and1 = s_csamul_rca16_u_rca16_fa2_xor0 & s_csamul_rca16_u_rca16_fa1_or0;
  assign s_csamul_rca16_u_rca16_fa2_or0 = s_csamul_rca16_u_rca16_fa2_and0 | s_csamul_rca16_u_rca16_fa2_and1;
  assign s_csamul_rca16_u_rca16_fa3_xor0 = s_csamul_rca16_fa4_15_xor1 ^ s_csamul_rca16_fa3_15_or0;
  assign s_csamul_rca16_u_rca16_fa3_and0 = s_csamul_rca16_fa4_15_xor1 & s_csamul_rca16_fa3_15_or0;
  assign s_csamul_rca16_u_rca16_fa3_xor1 = s_csamul_rca16_u_rca16_fa3_xor0 ^ s_csamul_rca16_u_rca16_fa2_or0;
  assign s_csamul_rca16_u_rca16_fa3_and1 = s_csamul_rca16_u_rca16_fa3_xor0 & s_csamul_rca16_u_rca16_fa2_or0;
  assign s_csamul_rca16_u_rca16_fa3_or0 = s_csamul_rca16_u_rca16_fa3_and0 | s_csamul_rca16_u_rca16_fa3_and1;
  assign s_csamul_rca16_u_rca16_fa4_xor0 = s_csamul_rca16_fa5_15_xor1 ^ s_csamul_rca16_fa4_15_or0;
  assign s_csamul_rca16_u_rca16_fa4_and0 = s_csamul_rca16_fa5_15_xor1 & s_csamul_rca16_fa4_15_or0;
  assign s_csamul_rca16_u_rca16_fa4_xor1 = s_csamul_rca16_u_rca16_fa4_xor0 ^ s_csamul_rca16_u_rca16_fa3_or0;
  assign s_csamul_rca16_u_rca16_fa4_and1 = s_csamul_rca16_u_rca16_fa4_xor0 & s_csamul_rca16_u_rca16_fa3_or0;
  assign s_csamul_rca16_u_rca16_fa4_or0 = s_csamul_rca16_u_rca16_fa4_and0 | s_csamul_rca16_u_rca16_fa4_and1;
  assign s_csamul_rca16_u_rca16_fa5_xor0 = s_csamul_rca16_fa6_15_xor1 ^ s_csamul_rca16_fa5_15_or0;
  assign s_csamul_rca16_u_rca16_fa5_and0 = s_csamul_rca16_fa6_15_xor1 & s_csamul_rca16_fa5_15_or0;
  assign s_csamul_rca16_u_rca16_fa5_xor1 = s_csamul_rca16_u_rca16_fa5_xor0 ^ s_csamul_rca16_u_rca16_fa4_or0;
  assign s_csamul_rca16_u_rca16_fa5_and1 = s_csamul_rca16_u_rca16_fa5_xor0 & s_csamul_rca16_u_rca16_fa4_or0;
  assign s_csamul_rca16_u_rca16_fa5_or0 = s_csamul_rca16_u_rca16_fa5_and0 | s_csamul_rca16_u_rca16_fa5_and1;
  assign s_csamul_rca16_u_rca16_fa6_xor0 = s_csamul_rca16_fa7_15_xor1 ^ s_csamul_rca16_fa6_15_or0;
  assign s_csamul_rca16_u_rca16_fa6_and0 = s_csamul_rca16_fa7_15_xor1 & s_csamul_rca16_fa6_15_or0;
  assign s_csamul_rca16_u_rca16_fa6_xor1 = s_csamul_rca16_u_rca16_fa6_xor0 ^ s_csamul_rca16_u_rca16_fa5_or0;
  assign s_csamul_rca16_u_rca16_fa6_and1 = s_csamul_rca16_u_rca16_fa6_xor0 & s_csamul_rca16_u_rca16_fa5_or0;
  assign s_csamul_rca16_u_rca16_fa6_or0 = s_csamul_rca16_u_rca16_fa6_and0 | s_csamul_rca16_u_rca16_fa6_and1;
  assign s_csamul_rca16_u_rca16_fa7_xor0 = s_csamul_rca16_fa8_15_xor1 ^ s_csamul_rca16_fa7_15_or0;
  assign s_csamul_rca16_u_rca16_fa7_and0 = s_csamul_rca16_fa8_15_xor1 & s_csamul_rca16_fa7_15_or0;
  assign s_csamul_rca16_u_rca16_fa7_xor1 = s_csamul_rca16_u_rca16_fa7_xor0 ^ s_csamul_rca16_u_rca16_fa6_or0;
  assign s_csamul_rca16_u_rca16_fa7_and1 = s_csamul_rca16_u_rca16_fa7_xor0 & s_csamul_rca16_u_rca16_fa6_or0;
  assign s_csamul_rca16_u_rca16_fa7_or0 = s_csamul_rca16_u_rca16_fa7_and0 | s_csamul_rca16_u_rca16_fa7_and1;
  assign s_csamul_rca16_u_rca16_fa8_xor0 = s_csamul_rca16_fa9_15_xor1 ^ s_csamul_rca16_fa8_15_or0;
  assign s_csamul_rca16_u_rca16_fa8_and0 = s_csamul_rca16_fa9_15_xor1 & s_csamul_rca16_fa8_15_or0;
  assign s_csamul_rca16_u_rca16_fa8_xor1 = s_csamul_rca16_u_rca16_fa8_xor0 ^ s_csamul_rca16_u_rca16_fa7_or0;
  assign s_csamul_rca16_u_rca16_fa8_and1 = s_csamul_rca16_u_rca16_fa8_xor0 & s_csamul_rca16_u_rca16_fa7_or0;
  assign s_csamul_rca16_u_rca16_fa8_or0 = s_csamul_rca16_u_rca16_fa8_and0 | s_csamul_rca16_u_rca16_fa8_and1;
  assign s_csamul_rca16_u_rca16_fa9_xor0 = s_csamul_rca16_fa10_15_xor1 ^ s_csamul_rca16_fa9_15_or0;
  assign s_csamul_rca16_u_rca16_fa9_and0 = s_csamul_rca16_fa10_15_xor1 & s_csamul_rca16_fa9_15_or0;
  assign s_csamul_rca16_u_rca16_fa9_xor1 = s_csamul_rca16_u_rca16_fa9_xor0 ^ s_csamul_rca16_u_rca16_fa8_or0;
  assign s_csamul_rca16_u_rca16_fa9_and1 = s_csamul_rca16_u_rca16_fa9_xor0 & s_csamul_rca16_u_rca16_fa8_or0;
  assign s_csamul_rca16_u_rca16_fa9_or0 = s_csamul_rca16_u_rca16_fa9_and0 | s_csamul_rca16_u_rca16_fa9_and1;
  assign s_csamul_rca16_u_rca16_fa10_xor0 = s_csamul_rca16_fa11_15_xor1 ^ s_csamul_rca16_fa10_15_or0;
  assign s_csamul_rca16_u_rca16_fa10_and0 = s_csamul_rca16_fa11_15_xor1 & s_csamul_rca16_fa10_15_or0;
  assign s_csamul_rca16_u_rca16_fa10_xor1 = s_csamul_rca16_u_rca16_fa10_xor0 ^ s_csamul_rca16_u_rca16_fa9_or0;
  assign s_csamul_rca16_u_rca16_fa10_and1 = s_csamul_rca16_u_rca16_fa10_xor0 & s_csamul_rca16_u_rca16_fa9_or0;
  assign s_csamul_rca16_u_rca16_fa10_or0 = s_csamul_rca16_u_rca16_fa10_and0 | s_csamul_rca16_u_rca16_fa10_and1;
  assign s_csamul_rca16_u_rca16_fa11_xor0 = s_csamul_rca16_fa12_15_xor1 ^ s_csamul_rca16_fa11_15_or0;
  assign s_csamul_rca16_u_rca16_fa11_and0 = s_csamul_rca16_fa12_15_xor1 & s_csamul_rca16_fa11_15_or0;
  assign s_csamul_rca16_u_rca16_fa11_xor1 = s_csamul_rca16_u_rca16_fa11_xor0 ^ s_csamul_rca16_u_rca16_fa10_or0;
  assign s_csamul_rca16_u_rca16_fa11_and1 = s_csamul_rca16_u_rca16_fa11_xor0 & s_csamul_rca16_u_rca16_fa10_or0;
  assign s_csamul_rca16_u_rca16_fa11_or0 = s_csamul_rca16_u_rca16_fa11_and0 | s_csamul_rca16_u_rca16_fa11_and1;
  assign s_csamul_rca16_u_rca16_fa12_xor0 = s_csamul_rca16_fa13_15_xor1 ^ s_csamul_rca16_fa12_15_or0;
  assign s_csamul_rca16_u_rca16_fa12_and0 = s_csamul_rca16_fa13_15_xor1 & s_csamul_rca16_fa12_15_or0;
  assign s_csamul_rca16_u_rca16_fa12_xor1 = s_csamul_rca16_u_rca16_fa12_xor0 ^ s_csamul_rca16_u_rca16_fa11_or0;
  assign s_csamul_rca16_u_rca16_fa12_and1 = s_csamul_rca16_u_rca16_fa12_xor0 & s_csamul_rca16_u_rca16_fa11_or0;
  assign s_csamul_rca16_u_rca16_fa12_or0 = s_csamul_rca16_u_rca16_fa12_and0 | s_csamul_rca16_u_rca16_fa12_and1;
  assign s_csamul_rca16_u_rca16_fa13_xor0 = s_csamul_rca16_fa14_15_xor1 ^ s_csamul_rca16_fa13_15_or0;
  assign s_csamul_rca16_u_rca16_fa13_and0 = s_csamul_rca16_fa14_15_xor1 & s_csamul_rca16_fa13_15_or0;
  assign s_csamul_rca16_u_rca16_fa13_xor1 = s_csamul_rca16_u_rca16_fa13_xor0 ^ s_csamul_rca16_u_rca16_fa12_or0;
  assign s_csamul_rca16_u_rca16_fa13_and1 = s_csamul_rca16_u_rca16_fa13_xor0 & s_csamul_rca16_u_rca16_fa12_or0;
  assign s_csamul_rca16_u_rca16_fa13_or0 = s_csamul_rca16_u_rca16_fa13_and0 | s_csamul_rca16_u_rca16_fa13_and1;
  assign s_csamul_rca16_u_rca16_fa14_xor0 = s_csamul_rca16_ha15_15_xor0 ^ s_csamul_rca16_fa14_15_or0;
  assign s_csamul_rca16_u_rca16_fa14_and0 = s_csamul_rca16_ha15_15_xor0 & s_csamul_rca16_fa14_15_or0;
  assign s_csamul_rca16_u_rca16_fa14_xor1 = s_csamul_rca16_u_rca16_fa14_xor0 ^ s_csamul_rca16_u_rca16_fa13_or0;
  assign s_csamul_rca16_u_rca16_fa14_and1 = s_csamul_rca16_u_rca16_fa14_xor0 & s_csamul_rca16_u_rca16_fa13_or0;
  assign s_csamul_rca16_u_rca16_fa14_or0 = s_csamul_rca16_u_rca16_fa14_and0 | s_csamul_rca16_u_rca16_fa14_and1;
  assign s_csamul_rca16_u_rca16_fa15_xor0 = ~s_csamul_rca16_ha15_15_and0;
  assign s_csamul_rca16_u_rca16_fa15_xor1 = s_csamul_rca16_u_rca16_fa15_xor0 ^ s_csamul_rca16_u_rca16_fa14_or0;
  assign s_csamul_rca16_u_rca16_fa15_and1 = s_csamul_rca16_u_rca16_fa15_xor0 & s_csamul_rca16_u_rca16_fa14_or0;
  assign s_csamul_rca16_u_rca16_fa15_or0 = s_csamul_rca16_ha15_15_and0 | s_csamul_rca16_u_rca16_fa15_and1;

  assign s_csamul_rca16_out[0] = s_csamul_rca16_and0_0;
  assign s_csamul_rca16_out[1] = s_csamul_rca16_ha0_1_xor0;
  assign s_csamul_rca16_out[2] = s_csamul_rca16_fa0_2_xor1;
  assign s_csamul_rca16_out[3] = s_csamul_rca16_fa0_3_xor1;
  assign s_csamul_rca16_out[4] = s_csamul_rca16_fa0_4_xor1;
  assign s_csamul_rca16_out[5] = s_csamul_rca16_fa0_5_xor1;
  assign s_csamul_rca16_out[6] = s_csamul_rca16_fa0_6_xor1;
  assign s_csamul_rca16_out[7] = s_csamul_rca16_fa0_7_xor1;
  assign s_csamul_rca16_out[8] = s_csamul_rca16_fa0_8_xor1;
  assign s_csamul_rca16_out[9] = s_csamul_rca16_fa0_9_xor1;
  assign s_csamul_rca16_out[10] = s_csamul_rca16_fa0_10_xor1;
  assign s_csamul_rca16_out[11] = s_csamul_rca16_fa0_11_xor1;
  assign s_csamul_rca16_out[12] = s_csamul_rca16_fa0_12_xor1;
  assign s_csamul_rca16_out[13] = s_csamul_rca16_fa0_13_xor1;
  assign s_csamul_rca16_out[14] = s_csamul_rca16_fa0_14_xor1;
  assign s_csamul_rca16_out[15] = s_csamul_rca16_fa0_15_xor1;
  assign s_csamul_rca16_out[16] = s_csamul_rca16_u_rca16_ha_xor0;
  assign s_csamul_rca16_out[17] = s_csamul_rca16_u_rca16_fa1_xor1;
  assign s_csamul_rca16_out[18] = s_csamul_rca16_u_rca16_fa2_xor1;
  assign s_csamul_rca16_out[19] = s_csamul_rca16_u_rca16_fa3_xor1;
  assign s_csamul_rca16_out[20] = s_csamul_rca16_u_rca16_fa4_xor1;
  assign s_csamul_rca16_out[21] = s_csamul_rca16_u_rca16_fa5_xor1;
  assign s_csamul_rca16_out[22] = s_csamul_rca16_u_rca16_fa6_xor1;
  assign s_csamul_rca16_out[23] = s_csamul_rca16_u_rca16_fa7_xor1;
  assign s_csamul_rca16_out[24] = s_csamul_rca16_u_rca16_fa8_xor1;
  assign s_csamul_rca16_out[25] = s_csamul_rca16_u_rca16_fa9_xor1;
  assign s_csamul_rca16_out[26] = s_csamul_rca16_u_rca16_fa10_xor1;
  assign s_csamul_rca16_out[27] = s_csamul_rca16_u_rca16_fa11_xor1;
  assign s_csamul_rca16_out[28] = s_csamul_rca16_u_rca16_fa12_xor1;
  assign s_csamul_rca16_out[29] = s_csamul_rca16_u_rca16_fa13_xor1;
  assign s_csamul_rca16_out[30] = s_csamul_rca16_u_rca16_fa14_xor1;
  assign s_csamul_rca16_out[31] = s_csamul_rca16_u_rca16_fa15_xor1;
endmodule