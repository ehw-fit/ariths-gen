module f_u_cla12(input [11:0] a, input [11:0] b, output [12:0] f_u_cla12_out);
  wire f_u_cla12_pg_logic0_or0;
  wire f_u_cla12_pg_logic0_and0;
  wire f_u_cla12_pg_logic0_xor0;
  wire f_u_cla12_pg_logic1_or0;
  wire f_u_cla12_pg_logic1_and0;
  wire f_u_cla12_pg_logic1_xor0;
  wire f_u_cla12_xor1;
  wire f_u_cla12_and0;
  wire f_u_cla12_or0;
  wire f_u_cla12_pg_logic2_or0;
  wire f_u_cla12_pg_logic2_and0;
  wire f_u_cla12_pg_logic2_xor0;
  wire f_u_cla12_xor2;
  wire f_u_cla12_and1;
  wire f_u_cla12_and2;
  wire f_u_cla12_and3;
  wire f_u_cla12_and4;
  wire f_u_cla12_or1;
  wire f_u_cla12_or2;
  wire f_u_cla12_pg_logic3_or0;
  wire f_u_cla12_pg_logic3_and0;
  wire f_u_cla12_pg_logic3_xor0;
  wire f_u_cla12_xor3;
  wire f_u_cla12_and5;
  wire f_u_cla12_and6;
  wire f_u_cla12_and7;
  wire f_u_cla12_and8;
  wire f_u_cla12_and9;
  wire f_u_cla12_and10;
  wire f_u_cla12_and11;
  wire f_u_cla12_or3;
  wire f_u_cla12_or4;
  wire f_u_cla12_or5;
  wire f_u_cla12_pg_logic4_or0;
  wire f_u_cla12_pg_logic4_and0;
  wire f_u_cla12_pg_logic4_xor0;
  wire f_u_cla12_xor4;
  wire f_u_cla12_and12;
  wire f_u_cla12_or6;
  wire f_u_cla12_pg_logic5_or0;
  wire f_u_cla12_pg_logic5_and0;
  wire f_u_cla12_pg_logic5_xor0;
  wire f_u_cla12_xor5;
  wire f_u_cla12_and13;
  wire f_u_cla12_and14;
  wire f_u_cla12_and15;
  wire f_u_cla12_or7;
  wire f_u_cla12_or8;
  wire f_u_cla12_pg_logic6_or0;
  wire f_u_cla12_pg_logic6_and0;
  wire f_u_cla12_pg_logic6_xor0;
  wire f_u_cla12_xor6;
  wire f_u_cla12_and16;
  wire f_u_cla12_and17;
  wire f_u_cla12_and18;
  wire f_u_cla12_and19;
  wire f_u_cla12_and20;
  wire f_u_cla12_and21;
  wire f_u_cla12_or9;
  wire f_u_cla12_or10;
  wire f_u_cla12_or11;
  wire f_u_cla12_pg_logic7_or0;
  wire f_u_cla12_pg_logic7_and0;
  wire f_u_cla12_pg_logic7_xor0;
  wire f_u_cla12_xor7;
  wire f_u_cla12_and22;
  wire f_u_cla12_and23;
  wire f_u_cla12_and24;
  wire f_u_cla12_and25;
  wire f_u_cla12_and26;
  wire f_u_cla12_and27;
  wire f_u_cla12_and28;
  wire f_u_cla12_and29;
  wire f_u_cla12_and30;
  wire f_u_cla12_and31;
  wire f_u_cla12_or12;
  wire f_u_cla12_or13;
  wire f_u_cla12_or14;
  wire f_u_cla12_or15;
  wire f_u_cla12_pg_logic8_or0;
  wire f_u_cla12_pg_logic8_and0;
  wire f_u_cla12_pg_logic8_xor0;
  wire f_u_cla12_xor8;
  wire f_u_cla12_and32;
  wire f_u_cla12_or16;
  wire f_u_cla12_pg_logic9_or0;
  wire f_u_cla12_pg_logic9_and0;
  wire f_u_cla12_pg_logic9_xor0;
  wire f_u_cla12_xor9;
  wire f_u_cla12_and33;
  wire f_u_cla12_and34;
  wire f_u_cla12_and35;
  wire f_u_cla12_or17;
  wire f_u_cla12_or18;
  wire f_u_cla12_pg_logic10_or0;
  wire f_u_cla12_pg_logic10_and0;
  wire f_u_cla12_pg_logic10_xor0;
  wire f_u_cla12_xor10;
  wire f_u_cla12_and36;
  wire f_u_cla12_and37;
  wire f_u_cla12_and38;
  wire f_u_cla12_and39;
  wire f_u_cla12_and40;
  wire f_u_cla12_and41;
  wire f_u_cla12_or19;
  wire f_u_cla12_or20;
  wire f_u_cla12_or21;
  wire f_u_cla12_pg_logic11_or0;
  wire f_u_cla12_pg_logic11_and0;
  wire f_u_cla12_pg_logic11_xor0;
  wire f_u_cla12_xor11;
  wire f_u_cla12_and42;
  wire f_u_cla12_and43;
  wire f_u_cla12_and44;
  wire f_u_cla12_and45;
  wire f_u_cla12_and46;
  wire f_u_cla12_and47;
  wire f_u_cla12_and48;
  wire f_u_cla12_and49;
  wire f_u_cla12_and50;
  wire f_u_cla12_and51;
  wire f_u_cla12_or22;
  wire f_u_cla12_or23;
  wire f_u_cla12_or24;
  wire f_u_cla12_or25;

  assign f_u_cla12_pg_logic0_or0 = a[0] | b[0];
  assign f_u_cla12_pg_logic0_and0 = a[0] & b[0];
  assign f_u_cla12_pg_logic0_xor0 = a[0] ^ b[0];
  assign f_u_cla12_pg_logic1_or0 = a[1] | b[1];
  assign f_u_cla12_pg_logic1_and0 = a[1] & b[1];
  assign f_u_cla12_pg_logic1_xor0 = a[1] ^ b[1];
  assign f_u_cla12_xor1 = f_u_cla12_pg_logic1_xor0 ^ f_u_cla12_pg_logic0_and0;
  assign f_u_cla12_and0 = f_u_cla12_pg_logic0_and0 & f_u_cla12_pg_logic1_or0;
  assign f_u_cla12_or0 = f_u_cla12_pg_logic1_and0 | f_u_cla12_and0;
  assign f_u_cla12_pg_logic2_or0 = a[2] | b[2];
  assign f_u_cla12_pg_logic2_and0 = a[2] & b[2];
  assign f_u_cla12_pg_logic2_xor0 = a[2] ^ b[2];
  assign f_u_cla12_xor2 = f_u_cla12_pg_logic2_xor0 ^ f_u_cla12_or0;
  assign f_u_cla12_and1 = f_u_cla12_pg_logic2_or0 & f_u_cla12_pg_logic0_or0;
  assign f_u_cla12_and2 = f_u_cla12_pg_logic0_and0 & f_u_cla12_pg_logic2_or0;
  assign f_u_cla12_and3 = f_u_cla12_and2 & f_u_cla12_pg_logic1_or0;
  assign f_u_cla12_and4 = f_u_cla12_pg_logic1_and0 & f_u_cla12_pg_logic2_or0;
  assign f_u_cla12_or1 = f_u_cla12_and3 | f_u_cla12_and4;
  assign f_u_cla12_or2 = f_u_cla12_pg_logic2_and0 | f_u_cla12_or1;
  assign f_u_cla12_pg_logic3_or0 = a[3] | b[3];
  assign f_u_cla12_pg_logic3_and0 = a[3] & b[3];
  assign f_u_cla12_pg_logic3_xor0 = a[3] ^ b[3];
  assign f_u_cla12_xor3 = f_u_cla12_pg_logic3_xor0 ^ f_u_cla12_or2;
  assign f_u_cla12_and5 = f_u_cla12_pg_logic3_or0 & f_u_cla12_pg_logic1_or0;
  assign f_u_cla12_and6 = f_u_cla12_pg_logic0_and0 & f_u_cla12_pg_logic2_or0;
  assign f_u_cla12_and7 = f_u_cla12_pg_logic3_or0 & f_u_cla12_pg_logic1_or0;
  assign f_u_cla12_and8 = f_u_cla12_and6 & f_u_cla12_and7;
  assign f_u_cla12_and9 = f_u_cla12_pg_logic1_and0 & f_u_cla12_pg_logic3_or0;
  assign f_u_cla12_and10 = f_u_cla12_and9 & f_u_cla12_pg_logic2_or0;
  assign f_u_cla12_and11 = f_u_cla12_pg_logic2_and0 & f_u_cla12_pg_logic3_or0;
  assign f_u_cla12_or3 = f_u_cla12_and8 | f_u_cla12_and11;
  assign f_u_cla12_or4 = f_u_cla12_and10 | f_u_cla12_or3;
  assign f_u_cla12_or5 = f_u_cla12_pg_logic3_and0 | f_u_cla12_or4;
  assign f_u_cla12_pg_logic4_or0 = a[4] | b[4];
  assign f_u_cla12_pg_logic4_and0 = a[4] & b[4];
  assign f_u_cla12_pg_logic4_xor0 = a[4] ^ b[4];
  assign f_u_cla12_xor4 = f_u_cla12_pg_logic4_xor0 ^ f_u_cla12_or5;
  assign f_u_cla12_and12 = f_u_cla12_or5 & f_u_cla12_pg_logic4_or0;
  assign f_u_cla12_or6 = f_u_cla12_pg_logic4_and0 | f_u_cla12_and12;
  assign f_u_cla12_pg_logic5_or0 = a[5] | b[5];
  assign f_u_cla12_pg_logic5_and0 = a[5] & b[5];
  assign f_u_cla12_pg_logic5_xor0 = a[5] ^ b[5];
  assign f_u_cla12_xor5 = f_u_cla12_pg_logic5_xor0 ^ f_u_cla12_or6;
  assign f_u_cla12_and13 = f_u_cla12_or5 & f_u_cla12_pg_logic5_or0;
  assign f_u_cla12_and14 = f_u_cla12_and13 & f_u_cla12_pg_logic4_or0;
  assign f_u_cla12_and15 = f_u_cla12_pg_logic4_and0 & f_u_cla12_pg_logic5_or0;
  assign f_u_cla12_or7 = f_u_cla12_and14 | f_u_cla12_and15;
  assign f_u_cla12_or8 = f_u_cla12_pg_logic5_and0 | f_u_cla12_or7;
  assign f_u_cla12_pg_logic6_or0 = a[6] | b[6];
  assign f_u_cla12_pg_logic6_and0 = a[6] & b[6];
  assign f_u_cla12_pg_logic6_xor0 = a[6] ^ b[6];
  assign f_u_cla12_xor6 = f_u_cla12_pg_logic6_xor0 ^ f_u_cla12_or8;
  assign f_u_cla12_and16 = f_u_cla12_or5 & f_u_cla12_pg_logic5_or0;
  assign f_u_cla12_and17 = f_u_cla12_pg_logic6_or0 & f_u_cla12_pg_logic4_or0;
  assign f_u_cla12_and18 = f_u_cla12_and16 & f_u_cla12_and17;
  assign f_u_cla12_and19 = f_u_cla12_pg_logic4_and0 & f_u_cla12_pg_logic6_or0;
  assign f_u_cla12_and20 = f_u_cla12_and19 & f_u_cla12_pg_logic5_or0;
  assign f_u_cla12_and21 = f_u_cla12_pg_logic5_and0 & f_u_cla12_pg_logic6_or0;
  assign f_u_cla12_or9 = f_u_cla12_and18 | f_u_cla12_and20;
  assign f_u_cla12_or10 = f_u_cla12_or9 | f_u_cla12_and21;
  assign f_u_cla12_or11 = f_u_cla12_pg_logic6_and0 | f_u_cla12_or10;
  assign f_u_cla12_pg_logic7_or0 = a[7] | b[7];
  assign f_u_cla12_pg_logic7_and0 = a[7] & b[7];
  assign f_u_cla12_pg_logic7_xor0 = a[7] ^ b[7];
  assign f_u_cla12_xor7 = f_u_cla12_pg_logic7_xor0 ^ f_u_cla12_or11;
  assign f_u_cla12_and22 = f_u_cla12_or5 & f_u_cla12_pg_logic6_or0;
  assign f_u_cla12_and23 = f_u_cla12_pg_logic7_or0 & f_u_cla12_pg_logic5_or0;
  assign f_u_cla12_and24 = f_u_cla12_and22 & f_u_cla12_and23;
  assign f_u_cla12_and25 = f_u_cla12_and24 & f_u_cla12_pg_logic4_or0;
  assign f_u_cla12_and26 = f_u_cla12_pg_logic4_and0 & f_u_cla12_pg_logic6_or0;
  assign f_u_cla12_and27 = f_u_cla12_pg_logic7_or0 & f_u_cla12_pg_logic5_or0;
  assign f_u_cla12_and28 = f_u_cla12_and26 & f_u_cla12_and27;
  assign f_u_cla12_and29 = f_u_cla12_pg_logic5_and0 & f_u_cla12_pg_logic7_or0;
  assign f_u_cla12_and30 = f_u_cla12_and29 & f_u_cla12_pg_logic6_or0;
  assign f_u_cla12_and31 = f_u_cla12_pg_logic6_and0 & f_u_cla12_pg_logic7_or0;
  assign f_u_cla12_or12 = f_u_cla12_and25 | f_u_cla12_and30;
  assign f_u_cla12_or13 = f_u_cla12_and28 | f_u_cla12_and31;
  assign f_u_cla12_or14 = f_u_cla12_or12 | f_u_cla12_or13;
  assign f_u_cla12_or15 = f_u_cla12_pg_logic7_and0 | f_u_cla12_or14;
  assign f_u_cla12_pg_logic8_or0 = a[8] | b[8];
  assign f_u_cla12_pg_logic8_and0 = a[8] & b[8];
  assign f_u_cla12_pg_logic8_xor0 = a[8] ^ b[8];
  assign f_u_cla12_xor8 = f_u_cla12_pg_logic8_xor0 ^ f_u_cla12_or15;
  assign f_u_cla12_and32 = f_u_cla12_or15 & f_u_cla12_pg_logic8_or0;
  assign f_u_cla12_or16 = f_u_cla12_pg_logic8_and0 | f_u_cla12_and32;
  assign f_u_cla12_pg_logic9_or0 = a[9] | b[9];
  assign f_u_cla12_pg_logic9_and0 = a[9] & b[9];
  assign f_u_cla12_pg_logic9_xor0 = a[9] ^ b[9];
  assign f_u_cla12_xor9 = f_u_cla12_pg_logic9_xor0 ^ f_u_cla12_or16;
  assign f_u_cla12_and33 = f_u_cla12_or15 & f_u_cla12_pg_logic9_or0;
  assign f_u_cla12_and34 = f_u_cla12_and33 & f_u_cla12_pg_logic8_or0;
  assign f_u_cla12_and35 = f_u_cla12_pg_logic8_and0 & f_u_cla12_pg_logic9_or0;
  assign f_u_cla12_or17 = f_u_cla12_and34 | f_u_cla12_and35;
  assign f_u_cla12_or18 = f_u_cla12_pg_logic9_and0 | f_u_cla12_or17;
  assign f_u_cla12_pg_logic10_or0 = a[10] | b[10];
  assign f_u_cla12_pg_logic10_and0 = a[10] & b[10];
  assign f_u_cla12_pg_logic10_xor0 = a[10] ^ b[10];
  assign f_u_cla12_xor10 = f_u_cla12_pg_logic10_xor0 ^ f_u_cla12_or18;
  assign f_u_cla12_and36 = f_u_cla12_or15 & f_u_cla12_pg_logic9_or0;
  assign f_u_cla12_and37 = f_u_cla12_pg_logic10_or0 & f_u_cla12_pg_logic8_or0;
  assign f_u_cla12_and38 = f_u_cla12_and36 & f_u_cla12_and37;
  assign f_u_cla12_and39 = f_u_cla12_pg_logic8_and0 & f_u_cla12_pg_logic10_or0;
  assign f_u_cla12_and40 = f_u_cla12_and39 & f_u_cla12_pg_logic9_or0;
  assign f_u_cla12_and41 = f_u_cla12_pg_logic9_and0 & f_u_cla12_pg_logic10_or0;
  assign f_u_cla12_or19 = f_u_cla12_and38 | f_u_cla12_and40;
  assign f_u_cla12_or20 = f_u_cla12_or19 | f_u_cla12_and41;
  assign f_u_cla12_or21 = f_u_cla12_pg_logic10_and0 | f_u_cla12_or20;
  assign f_u_cla12_pg_logic11_or0 = a[11] | b[11];
  assign f_u_cla12_pg_logic11_and0 = a[11] & b[11];
  assign f_u_cla12_pg_logic11_xor0 = a[11] ^ b[11];
  assign f_u_cla12_xor11 = f_u_cla12_pg_logic11_xor0 ^ f_u_cla12_or21;
  assign f_u_cla12_and42 = f_u_cla12_or15 & f_u_cla12_pg_logic10_or0;
  assign f_u_cla12_and43 = f_u_cla12_pg_logic11_or0 & f_u_cla12_pg_logic9_or0;
  assign f_u_cla12_and44 = f_u_cla12_and42 & f_u_cla12_and43;
  assign f_u_cla12_and45 = f_u_cla12_and44 & f_u_cla12_pg_logic8_or0;
  assign f_u_cla12_and46 = f_u_cla12_pg_logic8_and0 & f_u_cla12_pg_logic10_or0;
  assign f_u_cla12_and47 = f_u_cla12_pg_logic11_or0 & f_u_cla12_pg_logic9_or0;
  assign f_u_cla12_and48 = f_u_cla12_and46 & f_u_cla12_and47;
  assign f_u_cla12_and49 = f_u_cla12_pg_logic9_and0 & f_u_cla12_pg_logic11_or0;
  assign f_u_cla12_and50 = f_u_cla12_and49 & f_u_cla12_pg_logic10_or0;
  assign f_u_cla12_and51 = f_u_cla12_pg_logic10_and0 & f_u_cla12_pg_logic11_or0;
  assign f_u_cla12_or22 = f_u_cla12_and45 | f_u_cla12_and50;
  assign f_u_cla12_or23 = f_u_cla12_and48 | f_u_cla12_and51;
  assign f_u_cla12_or24 = f_u_cla12_or22 | f_u_cla12_or23;
  assign f_u_cla12_or25 = f_u_cla12_pg_logic11_and0 | f_u_cla12_or24;

  assign f_u_cla12_out[0] = f_u_cla12_pg_logic0_xor0;
  assign f_u_cla12_out[1] = f_u_cla12_xor1;
  assign f_u_cla12_out[2] = f_u_cla12_xor2;
  assign f_u_cla12_out[3] = f_u_cla12_xor3;
  assign f_u_cla12_out[4] = f_u_cla12_xor4;
  assign f_u_cla12_out[5] = f_u_cla12_xor5;
  assign f_u_cla12_out[6] = f_u_cla12_xor6;
  assign f_u_cla12_out[7] = f_u_cla12_xor7;
  assign f_u_cla12_out[8] = f_u_cla12_xor8;
  assign f_u_cla12_out[9] = f_u_cla12_xor9;
  assign f_u_cla12_out[10] = f_u_cla12_xor10;
  assign f_u_cla12_out[11] = f_u_cla12_xor11;
  assign f_u_cla12_out[12] = f_u_cla12_or25;
endmodule