module u_CSAwallace_cska8(input [7:0] a, input [7:0] b, output [15:0] u_CSAwallace_cska8_out);
  wire u_CSAwallace_cska8_and_0_0;
  wire u_CSAwallace_cska8_and_1_0;
  wire u_CSAwallace_cska8_and_2_0;
  wire u_CSAwallace_cska8_and_3_0;
  wire u_CSAwallace_cska8_and_4_0;
  wire u_CSAwallace_cska8_and_5_0;
  wire u_CSAwallace_cska8_and_6_0;
  wire u_CSAwallace_cska8_and_7_0;
  wire u_CSAwallace_cska8_and_0_1;
  wire u_CSAwallace_cska8_and_1_1;
  wire u_CSAwallace_cska8_and_2_1;
  wire u_CSAwallace_cska8_and_3_1;
  wire u_CSAwallace_cska8_and_4_1;
  wire u_CSAwallace_cska8_and_5_1;
  wire u_CSAwallace_cska8_and_6_1;
  wire u_CSAwallace_cska8_and_7_1;
  wire u_CSAwallace_cska8_and_0_2;
  wire u_CSAwallace_cska8_and_1_2;
  wire u_CSAwallace_cska8_and_2_2;
  wire u_CSAwallace_cska8_and_3_2;
  wire u_CSAwallace_cska8_and_4_2;
  wire u_CSAwallace_cska8_and_5_2;
  wire u_CSAwallace_cska8_and_6_2;
  wire u_CSAwallace_cska8_and_7_2;
  wire u_CSAwallace_cska8_and_0_3;
  wire u_CSAwallace_cska8_and_1_3;
  wire u_CSAwallace_cska8_and_2_3;
  wire u_CSAwallace_cska8_and_3_3;
  wire u_CSAwallace_cska8_and_4_3;
  wire u_CSAwallace_cska8_and_5_3;
  wire u_CSAwallace_cska8_and_6_3;
  wire u_CSAwallace_cska8_and_7_3;
  wire u_CSAwallace_cska8_and_0_4;
  wire u_CSAwallace_cska8_and_1_4;
  wire u_CSAwallace_cska8_and_2_4;
  wire u_CSAwallace_cska8_and_3_4;
  wire u_CSAwallace_cska8_and_4_4;
  wire u_CSAwallace_cska8_and_5_4;
  wire u_CSAwallace_cska8_and_6_4;
  wire u_CSAwallace_cska8_and_7_4;
  wire u_CSAwallace_cska8_and_0_5;
  wire u_CSAwallace_cska8_and_1_5;
  wire u_CSAwallace_cska8_and_2_5;
  wire u_CSAwallace_cska8_and_3_5;
  wire u_CSAwallace_cska8_and_4_5;
  wire u_CSAwallace_cska8_and_5_5;
  wire u_CSAwallace_cska8_and_6_5;
  wire u_CSAwallace_cska8_and_7_5;
  wire u_CSAwallace_cska8_and_0_6;
  wire u_CSAwallace_cska8_and_1_6;
  wire u_CSAwallace_cska8_and_2_6;
  wire u_CSAwallace_cska8_and_3_6;
  wire u_CSAwallace_cska8_and_4_6;
  wire u_CSAwallace_cska8_and_5_6;
  wire u_CSAwallace_cska8_and_6_6;
  wire u_CSAwallace_cska8_and_7_6;
  wire u_CSAwallace_cska8_and_0_7;
  wire u_CSAwallace_cska8_and_1_7;
  wire u_CSAwallace_cska8_and_2_7;
  wire u_CSAwallace_cska8_and_3_7;
  wire u_CSAwallace_cska8_and_4_7;
  wire u_CSAwallace_cska8_and_5_7;
  wire u_CSAwallace_cska8_and_6_7;
  wire u_CSAwallace_cska8_and_7_7;
  wire u_CSAwallace_cska8_csa0_csa_component_fa1_xor0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa1_and0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa2_xor0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa2_and0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa2_xor1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa2_and1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa2_or0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa3_xor0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa3_and0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa3_xor1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa3_and1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa3_or0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa4_xor0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa4_and0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa4_xor1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa4_and1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa4_or0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa5_xor0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa5_and0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa5_xor1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa5_and1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa5_or0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa6_xor0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa6_and0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa6_xor1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa6_and1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa6_or0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa7_xor0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa7_and0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa7_xor1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa7_and1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa7_or0;
  wire u_CSAwallace_cska8_csa0_csa_component_fa8_xor1;
  wire u_CSAwallace_cska8_csa0_csa_component_fa8_and1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa4_xor0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa4_and0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa5_xor0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa5_and0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa5_xor1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa5_and1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa5_or0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa6_xor0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa6_and0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa6_xor1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa6_and1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa6_or0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa7_xor0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa7_and0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa7_xor1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa7_and1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa7_or0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa8_xor0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa8_and0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa8_xor1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa8_and1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa8_or0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa9_xor0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa9_and0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa9_xor1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa9_and1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa9_or0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa10_xor0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa10_and0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa10_xor1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa10_and1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa10_or0;
  wire u_CSAwallace_cska8_csa1_csa_component_fa11_xor1;
  wire u_CSAwallace_cska8_csa1_csa_component_fa11_and1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa2_xor0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa2_and0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa3_xor0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa3_and0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa3_xor1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa3_and1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa3_or0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa4_xor0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa4_and0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa4_xor1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa4_and1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa4_or0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa5_xor0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa5_and0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa5_xor1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa5_and1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa5_or0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa6_xor0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa6_and0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa6_xor1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa6_and1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa6_or0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa7_xor0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa7_and0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa7_xor1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa7_and1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa7_or0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa8_xor0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa8_and0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa8_xor1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa8_and1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa8_or0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa9_xor0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa9_and0;
  wire u_CSAwallace_cska8_csa2_csa_component_fa9_xor1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa9_and1;
  wire u_CSAwallace_cska8_csa2_csa_component_fa9_or0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa6_xor0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa6_and0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa7_xor0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa7_and0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa7_xor1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa7_and1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa7_or0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa8_xor0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa8_and0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa8_xor1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa8_and1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa8_or0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa9_xor0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa9_and0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa9_xor1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa9_and1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa9_or0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa10_xor0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa10_and0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa10_xor1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa10_and1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa10_or0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa11_xor0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa11_and0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa11_xor1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa11_and1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa11_or0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa12_xor0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa12_and0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa12_xor1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa12_and1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa12_or0;
  wire u_CSAwallace_cska8_csa3_csa_component_fa13_xor1;
  wire u_CSAwallace_cska8_csa3_csa_component_fa13_and1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa3_xor0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa3_and0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa4_xor0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa4_and0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa5_xor0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa5_and0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa5_xor1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa5_and1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa5_or0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa6_xor0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa6_and0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa6_xor1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa6_and1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa6_or0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa7_xor0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa7_and0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa7_xor1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa7_and1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa7_or0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa8_xor0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa8_and0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa8_xor1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa8_and1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa8_or0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa9_xor0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa9_and0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa9_xor1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa9_and1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa9_or0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa10_xor0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa10_and0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa10_xor1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa10_and1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa10_or0;
  wire u_CSAwallace_cska8_csa4_csa_component_fa11_xor1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa11_and1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa12_xor1;
  wire u_CSAwallace_cska8_csa4_csa_component_fa12_and1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa4_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa4_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa5_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa5_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa6_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa6_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa7_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa7_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa7_xor1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa7_and1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa7_or0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa8_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa8_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa8_xor1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa8_and1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa8_or0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa9_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa9_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa9_xor1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa9_and1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa9_or0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa10_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa10_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa10_xor1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa10_and1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa10_or0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa11_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa11_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa11_xor1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa11_and1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa11_or0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa12_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa12_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa12_xor1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa12_and1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa12_or0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa13_xor0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa13_and0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa13_xor1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa13_and1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa13_or0;
  wire u_CSAwallace_cska8_csa5_csa_component_fa14_xor1;
  wire u_CSAwallace_cska8_csa5_csa_component_fa14_and1;
  wire u_CSAwallace_cska8_u_cska16_and_propagate00;
  wire u_CSAwallace_cska8_u_cska16_and_propagate01;
  wire u_CSAwallace_cska8_u_cska16_and_propagate02;
  wire u_CSAwallace_cska8_u_cska16_mux2to10_not0;
  wire u_CSAwallace_cska8_u_cska16_xor5;
  wire u_CSAwallace_cska8_u_cska16_fa4_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa4_and0;
  wire u_CSAwallace_cska8_u_cska16_xor6;
  wire u_CSAwallace_cska8_u_cska16_fa5_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa5_and0;
  wire u_CSAwallace_cska8_u_cska16_fa5_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa5_and1;
  wire u_CSAwallace_cska8_u_cska16_fa5_or0;
  wire u_CSAwallace_cska8_u_cska16_xor7;
  wire u_CSAwallace_cska8_u_cska16_fa6_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa6_and0;
  wire u_CSAwallace_cska8_u_cska16_fa6_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa6_and1;
  wire u_CSAwallace_cska8_u_cska16_fa6_or0;
  wire u_CSAwallace_cska8_u_cska16_and_propagate13;
  wire u_CSAwallace_cska8_u_cska16_and_propagate14;
  wire u_CSAwallace_cska8_u_cska16_and_propagate15;
  wire u_CSAwallace_cska8_u_cska16_mux2to11_not0;
  wire u_CSAwallace_cska8_u_cska16_mux2to11_and1;
  wire u_CSAwallace_cska8_u_cska16_xor8;
  wire u_CSAwallace_cska8_u_cska16_fa7_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa7_and0;
  wire u_CSAwallace_cska8_u_cska16_fa7_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa7_and1;
  wire u_CSAwallace_cska8_u_cska16_fa7_or0;
  wire u_CSAwallace_cska8_u_cska16_xor9;
  wire u_CSAwallace_cska8_u_cska16_fa8_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa8_and0;
  wire u_CSAwallace_cska8_u_cska16_fa8_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa8_and1;
  wire u_CSAwallace_cska8_u_cska16_fa8_or0;
  wire u_CSAwallace_cska8_u_cska16_xor10;
  wire u_CSAwallace_cska8_u_cska16_fa9_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa9_and0;
  wire u_CSAwallace_cska8_u_cska16_fa9_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa9_and1;
  wire u_CSAwallace_cska8_u_cska16_fa9_or0;
  wire u_CSAwallace_cska8_u_cska16_xor11;
  wire u_CSAwallace_cska8_u_cska16_fa10_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa10_and0;
  wire u_CSAwallace_cska8_u_cska16_fa10_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa10_and1;
  wire u_CSAwallace_cska8_u_cska16_fa10_or0;
  wire u_CSAwallace_cska8_u_cska16_and_propagate26;
  wire u_CSAwallace_cska8_u_cska16_and_propagate27;
  wire u_CSAwallace_cska8_u_cska16_and_propagate28;
  wire u_CSAwallace_cska8_u_cska16_mux2to12_and0;
  wire u_CSAwallace_cska8_u_cska16_mux2to12_not0;
  wire u_CSAwallace_cska8_u_cska16_mux2to12_and1;
  wire u_CSAwallace_cska8_u_cska16_mux2to12_xor0;
  wire u_CSAwallace_cska8_u_cska16_xor12;
  wire u_CSAwallace_cska8_u_cska16_fa11_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa11_and0;
  wire u_CSAwallace_cska8_u_cska16_fa11_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa11_and1;
  wire u_CSAwallace_cska8_u_cska16_fa11_or0;
  wire u_CSAwallace_cska8_u_cska16_xor13;
  wire u_CSAwallace_cska8_u_cska16_fa12_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa12_and0;
  wire u_CSAwallace_cska8_u_cska16_fa12_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa12_and1;
  wire u_CSAwallace_cska8_u_cska16_fa12_or0;
  wire u_CSAwallace_cska8_u_cska16_xor14;
  wire u_CSAwallace_cska8_u_cska16_fa13_xor0;
  wire u_CSAwallace_cska8_u_cska16_fa13_and0;
  wire u_CSAwallace_cska8_u_cska16_fa13_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa13_and1;
  wire u_CSAwallace_cska8_u_cska16_fa13_or0;
  wire u_CSAwallace_cska8_u_cska16_fa14_xor1;
  wire u_CSAwallace_cska8_u_cska16_fa14_and1;
  wire u_CSAwallace_cska8_u_cska16_and_propagate39;
  wire u_CSAwallace_cska8_u_cska16_and_propagate310;
  wire u_CSAwallace_cska8_u_cska16_and_propagate311;
  wire u_CSAwallace_cska8_u_cska16_mux2to13_and0;
  wire u_CSAwallace_cska8_u_cska16_mux2to13_not0;
  wire u_CSAwallace_cska8_u_cska16_mux2to13_and1;
  wire u_CSAwallace_cska8_u_cska16_mux2to13_xor0;

  assign u_CSAwallace_cska8_and_0_0 = a[0] & b[0];
  assign u_CSAwallace_cska8_and_1_0 = a[1] & b[0];
  assign u_CSAwallace_cska8_and_2_0 = a[2] & b[0];
  assign u_CSAwallace_cska8_and_3_0 = a[3] & b[0];
  assign u_CSAwallace_cska8_and_4_0 = a[4] & b[0];
  assign u_CSAwallace_cska8_and_5_0 = a[5] & b[0];
  assign u_CSAwallace_cska8_and_6_0 = a[6] & b[0];
  assign u_CSAwallace_cska8_and_7_0 = a[7] & b[0];
  assign u_CSAwallace_cska8_and_0_1 = a[0] & b[1];
  assign u_CSAwallace_cska8_and_1_1 = a[1] & b[1];
  assign u_CSAwallace_cska8_and_2_1 = a[2] & b[1];
  assign u_CSAwallace_cska8_and_3_1 = a[3] & b[1];
  assign u_CSAwallace_cska8_and_4_1 = a[4] & b[1];
  assign u_CSAwallace_cska8_and_5_1 = a[5] & b[1];
  assign u_CSAwallace_cska8_and_6_1 = a[6] & b[1];
  assign u_CSAwallace_cska8_and_7_1 = a[7] & b[1];
  assign u_CSAwallace_cska8_and_0_2 = a[0] & b[2];
  assign u_CSAwallace_cska8_and_1_2 = a[1] & b[2];
  assign u_CSAwallace_cska8_and_2_2 = a[2] & b[2];
  assign u_CSAwallace_cska8_and_3_2 = a[3] & b[2];
  assign u_CSAwallace_cska8_and_4_2 = a[4] & b[2];
  assign u_CSAwallace_cska8_and_5_2 = a[5] & b[2];
  assign u_CSAwallace_cska8_and_6_2 = a[6] & b[2];
  assign u_CSAwallace_cska8_and_7_2 = a[7] & b[2];
  assign u_CSAwallace_cska8_and_0_3 = a[0] & b[3];
  assign u_CSAwallace_cska8_and_1_3 = a[1] & b[3];
  assign u_CSAwallace_cska8_and_2_3 = a[2] & b[3];
  assign u_CSAwallace_cska8_and_3_3 = a[3] & b[3];
  assign u_CSAwallace_cska8_and_4_3 = a[4] & b[3];
  assign u_CSAwallace_cska8_and_5_3 = a[5] & b[3];
  assign u_CSAwallace_cska8_and_6_3 = a[6] & b[3];
  assign u_CSAwallace_cska8_and_7_3 = a[7] & b[3];
  assign u_CSAwallace_cska8_and_0_4 = a[0] & b[4];
  assign u_CSAwallace_cska8_and_1_4 = a[1] & b[4];
  assign u_CSAwallace_cska8_and_2_4 = a[2] & b[4];
  assign u_CSAwallace_cska8_and_3_4 = a[3] & b[4];
  assign u_CSAwallace_cska8_and_4_4 = a[4] & b[4];
  assign u_CSAwallace_cska8_and_5_4 = a[5] & b[4];
  assign u_CSAwallace_cska8_and_6_4 = a[6] & b[4];
  assign u_CSAwallace_cska8_and_7_4 = a[7] & b[4];
  assign u_CSAwallace_cska8_and_0_5 = a[0] & b[5];
  assign u_CSAwallace_cska8_and_1_5 = a[1] & b[5];
  assign u_CSAwallace_cska8_and_2_5 = a[2] & b[5];
  assign u_CSAwallace_cska8_and_3_5 = a[3] & b[5];
  assign u_CSAwallace_cska8_and_4_5 = a[4] & b[5];
  assign u_CSAwallace_cska8_and_5_5 = a[5] & b[5];
  assign u_CSAwallace_cska8_and_6_5 = a[6] & b[5];
  assign u_CSAwallace_cska8_and_7_5 = a[7] & b[5];
  assign u_CSAwallace_cska8_and_0_6 = a[0] & b[6];
  assign u_CSAwallace_cska8_and_1_6 = a[1] & b[6];
  assign u_CSAwallace_cska8_and_2_6 = a[2] & b[6];
  assign u_CSAwallace_cska8_and_3_6 = a[3] & b[6];
  assign u_CSAwallace_cska8_and_4_6 = a[4] & b[6];
  assign u_CSAwallace_cska8_and_5_6 = a[5] & b[6];
  assign u_CSAwallace_cska8_and_6_6 = a[6] & b[6];
  assign u_CSAwallace_cska8_and_7_6 = a[7] & b[6];
  assign u_CSAwallace_cska8_and_0_7 = a[0] & b[7];
  assign u_CSAwallace_cska8_and_1_7 = a[1] & b[7];
  assign u_CSAwallace_cska8_and_2_7 = a[2] & b[7];
  assign u_CSAwallace_cska8_and_3_7 = a[3] & b[7];
  assign u_CSAwallace_cska8_and_4_7 = a[4] & b[7];
  assign u_CSAwallace_cska8_and_5_7 = a[5] & b[7];
  assign u_CSAwallace_cska8_and_6_7 = a[6] & b[7];
  assign u_CSAwallace_cska8_and_7_7 = a[7] & b[7];
  assign u_CSAwallace_cska8_csa0_csa_component_fa1_xor0 = u_CSAwallace_cska8_and_1_0 ^ u_CSAwallace_cska8_and_0_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa1_and0 = u_CSAwallace_cska8_and_1_0 & u_CSAwallace_cska8_and_0_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa2_xor0 = u_CSAwallace_cska8_and_2_0 ^ u_CSAwallace_cska8_and_1_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa2_and0 = u_CSAwallace_cska8_and_2_0 & u_CSAwallace_cska8_and_1_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa2_xor1 = u_CSAwallace_cska8_csa0_csa_component_fa2_xor0 ^ u_CSAwallace_cska8_and_0_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa2_and1 = u_CSAwallace_cska8_csa0_csa_component_fa2_xor0 & u_CSAwallace_cska8_and_0_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa2_or0 = u_CSAwallace_cska8_csa0_csa_component_fa2_and0 | u_CSAwallace_cska8_csa0_csa_component_fa2_and1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa3_xor0 = u_CSAwallace_cska8_and_3_0 ^ u_CSAwallace_cska8_and_2_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa3_and0 = u_CSAwallace_cska8_and_3_0 & u_CSAwallace_cska8_and_2_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa3_xor1 = u_CSAwallace_cska8_csa0_csa_component_fa3_xor0 ^ u_CSAwallace_cska8_and_1_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa3_and1 = u_CSAwallace_cska8_csa0_csa_component_fa3_xor0 & u_CSAwallace_cska8_and_1_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa3_or0 = u_CSAwallace_cska8_csa0_csa_component_fa3_and0 | u_CSAwallace_cska8_csa0_csa_component_fa3_and1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa4_xor0 = u_CSAwallace_cska8_and_4_0 ^ u_CSAwallace_cska8_and_3_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa4_and0 = u_CSAwallace_cska8_and_4_0 & u_CSAwallace_cska8_and_3_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa4_xor1 = u_CSAwallace_cska8_csa0_csa_component_fa4_xor0 ^ u_CSAwallace_cska8_and_2_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa4_and1 = u_CSAwallace_cska8_csa0_csa_component_fa4_xor0 & u_CSAwallace_cska8_and_2_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa4_or0 = u_CSAwallace_cska8_csa0_csa_component_fa4_and0 | u_CSAwallace_cska8_csa0_csa_component_fa4_and1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa5_xor0 = u_CSAwallace_cska8_and_5_0 ^ u_CSAwallace_cska8_and_4_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa5_and0 = u_CSAwallace_cska8_and_5_0 & u_CSAwallace_cska8_and_4_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa5_xor1 = u_CSAwallace_cska8_csa0_csa_component_fa5_xor0 ^ u_CSAwallace_cska8_and_3_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa5_and1 = u_CSAwallace_cska8_csa0_csa_component_fa5_xor0 & u_CSAwallace_cska8_and_3_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa5_or0 = u_CSAwallace_cska8_csa0_csa_component_fa5_and0 | u_CSAwallace_cska8_csa0_csa_component_fa5_and1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa6_xor0 = u_CSAwallace_cska8_and_6_0 ^ u_CSAwallace_cska8_and_5_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa6_and0 = u_CSAwallace_cska8_and_6_0 & u_CSAwallace_cska8_and_5_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa6_xor1 = u_CSAwallace_cska8_csa0_csa_component_fa6_xor0 ^ u_CSAwallace_cska8_and_4_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa6_and1 = u_CSAwallace_cska8_csa0_csa_component_fa6_xor0 & u_CSAwallace_cska8_and_4_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa6_or0 = u_CSAwallace_cska8_csa0_csa_component_fa6_and0 | u_CSAwallace_cska8_csa0_csa_component_fa6_and1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa7_xor0 = u_CSAwallace_cska8_and_7_0 ^ u_CSAwallace_cska8_and_6_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa7_and0 = u_CSAwallace_cska8_and_7_0 & u_CSAwallace_cska8_and_6_1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa7_xor1 = u_CSAwallace_cska8_csa0_csa_component_fa7_xor0 ^ u_CSAwallace_cska8_and_5_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa7_and1 = u_CSAwallace_cska8_csa0_csa_component_fa7_xor0 & u_CSAwallace_cska8_and_5_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa7_or0 = u_CSAwallace_cska8_csa0_csa_component_fa7_and0 | u_CSAwallace_cska8_csa0_csa_component_fa7_and1;
  assign u_CSAwallace_cska8_csa0_csa_component_fa8_xor1 = u_CSAwallace_cska8_and_7_1 ^ u_CSAwallace_cska8_and_6_2;
  assign u_CSAwallace_cska8_csa0_csa_component_fa8_and1 = u_CSAwallace_cska8_and_7_1 & u_CSAwallace_cska8_and_6_2;
  assign u_CSAwallace_cska8_csa1_csa_component_fa4_xor0 = u_CSAwallace_cska8_and_1_3 ^ u_CSAwallace_cska8_and_0_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa4_and0 = u_CSAwallace_cska8_and_1_3 & u_CSAwallace_cska8_and_0_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa5_xor0 = u_CSAwallace_cska8_and_2_3 ^ u_CSAwallace_cska8_and_1_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa5_and0 = u_CSAwallace_cska8_and_2_3 & u_CSAwallace_cska8_and_1_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa5_xor1 = u_CSAwallace_cska8_csa1_csa_component_fa5_xor0 ^ u_CSAwallace_cska8_and_0_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa5_and1 = u_CSAwallace_cska8_csa1_csa_component_fa5_xor0 & u_CSAwallace_cska8_and_0_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa5_or0 = u_CSAwallace_cska8_csa1_csa_component_fa5_and0 | u_CSAwallace_cska8_csa1_csa_component_fa5_and1;
  assign u_CSAwallace_cska8_csa1_csa_component_fa6_xor0 = u_CSAwallace_cska8_and_3_3 ^ u_CSAwallace_cska8_and_2_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa6_and0 = u_CSAwallace_cska8_and_3_3 & u_CSAwallace_cska8_and_2_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa6_xor1 = u_CSAwallace_cska8_csa1_csa_component_fa6_xor0 ^ u_CSAwallace_cska8_and_1_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa6_and1 = u_CSAwallace_cska8_csa1_csa_component_fa6_xor0 & u_CSAwallace_cska8_and_1_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa6_or0 = u_CSAwallace_cska8_csa1_csa_component_fa6_and0 | u_CSAwallace_cska8_csa1_csa_component_fa6_and1;
  assign u_CSAwallace_cska8_csa1_csa_component_fa7_xor0 = u_CSAwallace_cska8_and_4_3 ^ u_CSAwallace_cska8_and_3_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa7_and0 = u_CSAwallace_cska8_and_4_3 & u_CSAwallace_cska8_and_3_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa7_xor1 = u_CSAwallace_cska8_csa1_csa_component_fa7_xor0 ^ u_CSAwallace_cska8_and_2_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa7_and1 = u_CSAwallace_cska8_csa1_csa_component_fa7_xor0 & u_CSAwallace_cska8_and_2_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa7_or0 = u_CSAwallace_cska8_csa1_csa_component_fa7_and0 | u_CSAwallace_cska8_csa1_csa_component_fa7_and1;
  assign u_CSAwallace_cska8_csa1_csa_component_fa8_xor0 = u_CSAwallace_cska8_and_5_3 ^ u_CSAwallace_cska8_and_4_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa8_and0 = u_CSAwallace_cska8_and_5_3 & u_CSAwallace_cska8_and_4_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa8_xor1 = u_CSAwallace_cska8_csa1_csa_component_fa8_xor0 ^ u_CSAwallace_cska8_and_3_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa8_and1 = u_CSAwallace_cska8_csa1_csa_component_fa8_xor0 & u_CSAwallace_cska8_and_3_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa8_or0 = u_CSAwallace_cska8_csa1_csa_component_fa8_and0 | u_CSAwallace_cska8_csa1_csa_component_fa8_and1;
  assign u_CSAwallace_cska8_csa1_csa_component_fa9_xor0 = u_CSAwallace_cska8_and_6_3 ^ u_CSAwallace_cska8_and_5_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa9_and0 = u_CSAwallace_cska8_and_6_3 & u_CSAwallace_cska8_and_5_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa9_xor1 = u_CSAwallace_cska8_csa1_csa_component_fa9_xor0 ^ u_CSAwallace_cska8_and_4_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa9_and1 = u_CSAwallace_cska8_csa1_csa_component_fa9_xor0 & u_CSAwallace_cska8_and_4_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa9_or0 = u_CSAwallace_cska8_csa1_csa_component_fa9_and0 | u_CSAwallace_cska8_csa1_csa_component_fa9_and1;
  assign u_CSAwallace_cska8_csa1_csa_component_fa10_xor0 = u_CSAwallace_cska8_and_7_3 ^ u_CSAwallace_cska8_and_6_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa10_and0 = u_CSAwallace_cska8_and_7_3 & u_CSAwallace_cska8_and_6_4;
  assign u_CSAwallace_cska8_csa1_csa_component_fa10_xor1 = u_CSAwallace_cska8_csa1_csa_component_fa10_xor0 ^ u_CSAwallace_cska8_and_5_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa10_and1 = u_CSAwallace_cska8_csa1_csa_component_fa10_xor0 & u_CSAwallace_cska8_and_5_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa10_or0 = u_CSAwallace_cska8_csa1_csa_component_fa10_and0 | u_CSAwallace_cska8_csa1_csa_component_fa10_and1;
  assign u_CSAwallace_cska8_csa1_csa_component_fa11_xor1 = u_CSAwallace_cska8_and_7_4 ^ u_CSAwallace_cska8_and_6_5;
  assign u_CSAwallace_cska8_csa1_csa_component_fa11_and1 = u_CSAwallace_cska8_and_7_4 & u_CSAwallace_cska8_and_6_5;
  assign u_CSAwallace_cska8_csa2_csa_component_fa2_xor0 = u_CSAwallace_cska8_csa0_csa_component_fa2_xor1 ^ u_CSAwallace_cska8_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa2_and0 = u_CSAwallace_cska8_csa0_csa_component_fa2_xor1 & u_CSAwallace_cska8_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa3_xor0 = u_CSAwallace_cska8_csa0_csa_component_fa3_xor1 ^ u_CSAwallace_cska8_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa3_and0 = u_CSAwallace_cska8_csa0_csa_component_fa3_xor1 & u_CSAwallace_cska8_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa3_xor1 = u_CSAwallace_cska8_csa2_csa_component_fa3_xor0 ^ u_CSAwallace_cska8_and_0_3;
  assign u_CSAwallace_cska8_csa2_csa_component_fa3_and1 = u_CSAwallace_cska8_csa2_csa_component_fa3_xor0 & u_CSAwallace_cska8_and_0_3;
  assign u_CSAwallace_cska8_csa2_csa_component_fa3_or0 = u_CSAwallace_cska8_csa2_csa_component_fa3_and0 | u_CSAwallace_cska8_csa2_csa_component_fa3_and1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa4_xor0 = u_CSAwallace_cska8_csa0_csa_component_fa4_xor1 ^ u_CSAwallace_cska8_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa4_and0 = u_CSAwallace_cska8_csa0_csa_component_fa4_xor1 & u_CSAwallace_cska8_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa4_xor1 = u_CSAwallace_cska8_csa2_csa_component_fa4_xor0 ^ u_CSAwallace_cska8_csa1_csa_component_fa4_xor0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa4_and1 = u_CSAwallace_cska8_csa2_csa_component_fa4_xor0 & u_CSAwallace_cska8_csa1_csa_component_fa4_xor0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa4_or0 = u_CSAwallace_cska8_csa2_csa_component_fa4_and0 | u_CSAwallace_cska8_csa2_csa_component_fa4_and1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa5_xor0 = u_CSAwallace_cska8_csa0_csa_component_fa5_xor1 ^ u_CSAwallace_cska8_csa0_csa_component_fa4_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa5_and0 = u_CSAwallace_cska8_csa0_csa_component_fa5_xor1 & u_CSAwallace_cska8_csa0_csa_component_fa4_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa5_xor1 = u_CSAwallace_cska8_csa2_csa_component_fa5_xor0 ^ u_CSAwallace_cska8_csa1_csa_component_fa5_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa5_and1 = u_CSAwallace_cska8_csa2_csa_component_fa5_xor0 & u_CSAwallace_cska8_csa1_csa_component_fa5_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa5_or0 = u_CSAwallace_cska8_csa2_csa_component_fa5_and0 | u_CSAwallace_cska8_csa2_csa_component_fa5_and1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa6_xor0 = u_CSAwallace_cska8_csa0_csa_component_fa6_xor1 ^ u_CSAwallace_cska8_csa0_csa_component_fa5_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa6_and0 = u_CSAwallace_cska8_csa0_csa_component_fa6_xor1 & u_CSAwallace_cska8_csa0_csa_component_fa5_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa6_xor1 = u_CSAwallace_cska8_csa2_csa_component_fa6_xor0 ^ u_CSAwallace_cska8_csa1_csa_component_fa6_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa6_and1 = u_CSAwallace_cska8_csa2_csa_component_fa6_xor0 & u_CSAwallace_cska8_csa1_csa_component_fa6_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa6_or0 = u_CSAwallace_cska8_csa2_csa_component_fa6_and0 | u_CSAwallace_cska8_csa2_csa_component_fa6_and1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa7_xor0 = u_CSAwallace_cska8_csa0_csa_component_fa7_xor1 ^ u_CSAwallace_cska8_csa0_csa_component_fa6_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa7_and0 = u_CSAwallace_cska8_csa0_csa_component_fa7_xor1 & u_CSAwallace_cska8_csa0_csa_component_fa6_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa7_xor1 = u_CSAwallace_cska8_csa2_csa_component_fa7_xor0 ^ u_CSAwallace_cska8_csa1_csa_component_fa7_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa7_and1 = u_CSAwallace_cska8_csa2_csa_component_fa7_xor0 & u_CSAwallace_cska8_csa1_csa_component_fa7_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa7_or0 = u_CSAwallace_cska8_csa2_csa_component_fa7_and0 | u_CSAwallace_cska8_csa2_csa_component_fa7_and1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa8_xor0 = u_CSAwallace_cska8_csa0_csa_component_fa8_xor1 ^ u_CSAwallace_cska8_csa0_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa8_and0 = u_CSAwallace_cska8_csa0_csa_component_fa8_xor1 & u_CSAwallace_cska8_csa0_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_csa2_csa_component_fa8_xor1 = u_CSAwallace_cska8_csa2_csa_component_fa8_xor0 ^ u_CSAwallace_cska8_csa1_csa_component_fa8_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa8_and1 = u_CSAwallace_cska8_csa2_csa_component_fa8_xor0 & u_CSAwallace_cska8_csa1_csa_component_fa8_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa8_or0 = u_CSAwallace_cska8_csa2_csa_component_fa8_and0 | u_CSAwallace_cska8_csa2_csa_component_fa8_and1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa9_xor0 = u_CSAwallace_cska8_and_7_2 ^ u_CSAwallace_cska8_csa0_csa_component_fa8_and1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa9_and0 = u_CSAwallace_cska8_and_7_2 & u_CSAwallace_cska8_csa0_csa_component_fa8_and1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa9_xor1 = u_CSAwallace_cska8_csa2_csa_component_fa9_xor0 ^ u_CSAwallace_cska8_csa1_csa_component_fa9_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa9_and1 = u_CSAwallace_cska8_csa2_csa_component_fa9_xor0 & u_CSAwallace_cska8_csa1_csa_component_fa9_xor1;
  assign u_CSAwallace_cska8_csa2_csa_component_fa9_or0 = u_CSAwallace_cska8_csa2_csa_component_fa9_and0 | u_CSAwallace_cska8_csa2_csa_component_fa9_and1;
  assign u_CSAwallace_cska8_csa3_csa_component_fa6_xor0 = u_CSAwallace_cska8_csa1_csa_component_fa5_or0 ^ u_CSAwallace_cska8_and_0_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa6_and0 = u_CSAwallace_cska8_csa1_csa_component_fa5_or0 & u_CSAwallace_cska8_and_0_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa7_xor0 = u_CSAwallace_cska8_csa1_csa_component_fa6_or0 ^ u_CSAwallace_cska8_and_1_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa7_and0 = u_CSAwallace_cska8_csa1_csa_component_fa6_or0 & u_CSAwallace_cska8_and_1_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa7_xor1 = u_CSAwallace_cska8_csa3_csa_component_fa7_xor0 ^ u_CSAwallace_cska8_and_0_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa7_and1 = u_CSAwallace_cska8_csa3_csa_component_fa7_xor0 & u_CSAwallace_cska8_and_0_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa7_or0 = u_CSAwallace_cska8_csa3_csa_component_fa7_and0 | u_CSAwallace_cska8_csa3_csa_component_fa7_and1;
  assign u_CSAwallace_cska8_csa3_csa_component_fa8_xor0 = u_CSAwallace_cska8_csa1_csa_component_fa7_or0 ^ u_CSAwallace_cska8_and_2_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa8_and0 = u_CSAwallace_cska8_csa1_csa_component_fa7_or0 & u_CSAwallace_cska8_and_2_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa8_xor1 = u_CSAwallace_cska8_csa3_csa_component_fa8_xor0 ^ u_CSAwallace_cska8_and_1_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa8_and1 = u_CSAwallace_cska8_csa3_csa_component_fa8_xor0 & u_CSAwallace_cska8_and_1_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa8_or0 = u_CSAwallace_cska8_csa3_csa_component_fa8_and0 | u_CSAwallace_cska8_csa3_csa_component_fa8_and1;
  assign u_CSAwallace_cska8_csa3_csa_component_fa9_xor0 = u_CSAwallace_cska8_csa1_csa_component_fa8_or0 ^ u_CSAwallace_cska8_and_3_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa9_and0 = u_CSAwallace_cska8_csa1_csa_component_fa8_or0 & u_CSAwallace_cska8_and_3_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa9_xor1 = u_CSAwallace_cska8_csa3_csa_component_fa9_xor0 ^ u_CSAwallace_cska8_and_2_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa9_and1 = u_CSAwallace_cska8_csa3_csa_component_fa9_xor0 & u_CSAwallace_cska8_and_2_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa9_or0 = u_CSAwallace_cska8_csa3_csa_component_fa9_and0 | u_CSAwallace_cska8_csa3_csa_component_fa9_and1;
  assign u_CSAwallace_cska8_csa3_csa_component_fa10_xor0 = u_CSAwallace_cska8_csa1_csa_component_fa9_or0 ^ u_CSAwallace_cska8_and_4_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa10_and0 = u_CSAwallace_cska8_csa1_csa_component_fa9_or0 & u_CSAwallace_cska8_and_4_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa10_xor1 = u_CSAwallace_cska8_csa3_csa_component_fa10_xor0 ^ u_CSAwallace_cska8_and_3_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa10_and1 = u_CSAwallace_cska8_csa3_csa_component_fa10_xor0 & u_CSAwallace_cska8_and_3_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa10_or0 = u_CSAwallace_cska8_csa3_csa_component_fa10_and0 | u_CSAwallace_cska8_csa3_csa_component_fa10_and1;
  assign u_CSAwallace_cska8_csa3_csa_component_fa11_xor0 = u_CSAwallace_cska8_csa1_csa_component_fa10_or0 ^ u_CSAwallace_cska8_and_5_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa11_and0 = u_CSAwallace_cska8_csa1_csa_component_fa10_or0 & u_CSAwallace_cska8_and_5_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa11_xor1 = u_CSAwallace_cska8_csa3_csa_component_fa11_xor0 ^ u_CSAwallace_cska8_and_4_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa11_and1 = u_CSAwallace_cska8_csa3_csa_component_fa11_xor0 & u_CSAwallace_cska8_and_4_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa11_or0 = u_CSAwallace_cska8_csa3_csa_component_fa11_and0 | u_CSAwallace_cska8_csa3_csa_component_fa11_and1;
  assign u_CSAwallace_cska8_csa3_csa_component_fa12_xor0 = u_CSAwallace_cska8_csa1_csa_component_fa11_and1 ^ u_CSAwallace_cska8_and_6_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa12_and0 = u_CSAwallace_cska8_csa1_csa_component_fa11_and1 & u_CSAwallace_cska8_and_6_6;
  assign u_CSAwallace_cska8_csa3_csa_component_fa12_xor1 = u_CSAwallace_cska8_csa3_csa_component_fa12_xor0 ^ u_CSAwallace_cska8_and_5_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa12_and1 = u_CSAwallace_cska8_csa3_csa_component_fa12_xor0 & u_CSAwallace_cska8_and_5_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa12_or0 = u_CSAwallace_cska8_csa3_csa_component_fa12_and0 | u_CSAwallace_cska8_csa3_csa_component_fa12_and1;
  assign u_CSAwallace_cska8_csa3_csa_component_fa13_xor1 = u_CSAwallace_cska8_and_7_6 ^ u_CSAwallace_cska8_and_6_7;
  assign u_CSAwallace_cska8_csa3_csa_component_fa13_and1 = u_CSAwallace_cska8_and_7_6 & u_CSAwallace_cska8_and_6_7;
  assign u_CSAwallace_cska8_csa4_csa_component_fa3_xor0 = u_CSAwallace_cska8_csa2_csa_component_fa3_xor1 ^ u_CSAwallace_cska8_csa2_csa_component_fa2_and0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa3_and0 = u_CSAwallace_cska8_csa2_csa_component_fa3_xor1 & u_CSAwallace_cska8_csa2_csa_component_fa2_and0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa4_xor0 = u_CSAwallace_cska8_csa2_csa_component_fa4_xor1 ^ u_CSAwallace_cska8_csa2_csa_component_fa3_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa4_and0 = u_CSAwallace_cska8_csa2_csa_component_fa4_xor1 & u_CSAwallace_cska8_csa2_csa_component_fa3_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa5_xor0 = u_CSAwallace_cska8_csa2_csa_component_fa5_xor1 ^ u_CSAwallace_cska8_csa2_csa_component_fa4_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa5_and0 = u_CSAwallace_cska8_csa2_csa_component_fa5_xor1 & u_CSAwallace_cska8_csa2_csa_component_fa4_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa5_xor1 = u_CSAwallace_cska8_csa4_csa_component_fa5_xor0 ^ u_CSAwallace_cska8_csa1_csa_component_fa4_and0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa5_and1 = u_CSAwallace_cska8_csa4_csa_component_fa5_xor0 & u_CSAwallace_cska8_csa1_csa_component_fa4_and0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa5_or0 = u_CSAwallace_cska8_csa4_csa_component_fa5_and0 | u_CSAwallace_cska8_csa4_csa_component_fa5_and1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa6_xor0 = u_CSAwallace_cska8_csa2_csa_component_fa6_xor1 ^ u_CSAwallace_cska8_csa2_csa_component_fa5_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa6_and0 = u_CSAwallace_cska8_csa2_csa_component_fa6_xor1 & u_CSAwallace_cska8_csa2_csa_component_fa5_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa6_xor1 = u_CSAwallace_cska8_csa4_csa_component_fa6_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa6_xor0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa6_and1 = u_CSAwallace_cska8_csa4_csa_component_fa6_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa6_xor0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa6_or0 = u_CSAwallace_cska8_csa4_csa_component_fa6_and0 | u_CSAwallace_cska8_csa4_csa_component_fa6_and1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa7_xor0 = u_CSAwallace_cska8_csa2_csa_component_fa7_xor1 ^ u_CSAwallace_cska8_csa2_csa_component_fa6_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa7_and0 = u_CSAwallace_cska8_csa2_csa_component_fa7_xor1 & u_CSAwallace_cska8_csa2_csa_component_fa6_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa7_xor1 = u_CSAwallace_cska8_csa4_csa_component_fa7_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa7_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa7_and1 = u_CSAwallace_cska8_csa4_csa_component_fa7_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa7_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa7_or0 = u_CSAwallace_cska8_csa4_csa_component_fa7_and0 | u_CSAwallace_cska8_csa4_csa_component_fa7_and1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa8_xor0 = u_CSAwallace_cska8_csa2_csa_component_fa8_xor1 ^ u_CSAwallace_cska8_csa2_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa8_and0 = u_CSAwallace_cska8_csa2_csa_component_fa8_xor1 & u_CSAwallace_cska8_csa2_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa8_xor1 = u_CSAwallace_cska8_csa4_csa_component_fa8_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa8_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa8_and1 = u_CSAwallace_cska8_csa4_csa_component_fa8_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa8_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa8_or0 = u_CSAwallace_cska8_csa4_csa_component_fa8_and0 | u_CSAwallace_cska8_csa4_csa_component_fa8_and1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa9_xor0 = u_CSAwallace_cska8_csa2_csa_component_fa9_xor1 ^ u_CSAwallace_cska8_csa2_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa9_and0 = u_CSAwallace_cska8_csa2_csa_component_fa9_xor1 & u_CSAwallace_cska8_csa2_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa9_xor1 = u_CSAwallace_cska8_csa4_csa_component_fa9_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa9_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa9_and1 = u_CSAwallace_cska8_csa4_csa_component_fa9_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa9_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa9_or0 = u_CSAwallace_cska8_csa4_csa_component_fa9_and0 | u_CSAwallace_cska8_csa4_csa_component_fa9_and1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa10_xor0 = u_CSAwallace_cska8_csa1_csa_component_fa10_xor1 ^ u_CSAwallace_cska8_csa2_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa10_and0 = u_CSAwallace_cska8_csa1_csa_component_fa10_xor1 & u_CSAwallace_cska8_csa2_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_csa4_csa_component_fa10_xor1 = u_CSAwallace_cska8_csa4_csa_component_fa10_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa10_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa10_and1 = u_CSAwallace_cska8_csa4_csa_component_fa10_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa10_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa10_or0 = u_CSAwallace_cska8_csa4_csa_component_fa10_and0 | u_CSAwallace_cska8_csa4_csa_component_fa10_and1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa11_xor1 = u_CSAwallace_cska8_csa1_csa_component_fa11_xor1 ^ u_CSAwallace_cska8_csa3_csa_component_fa11_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa11_and1 = u_CSAwallace_cska8_csa1_csa_component_fa11_xor1 & u_CSAwallace_cska8_csa3_csa_component_fa11_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa12_xor1 = u_CSAwallace_cska8_and_7_5 ^ u_CSAwallace_cska8_csa3_csa_component_fa12_xor1;
  assign u_CSAwallace_cska8_csa4_csa_component_fa12_and1 = u_CSAwallace_cska8_and_7_5 & u_CSAwallace_cska8_csa3_csa_component_fa12_xor1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa4_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa4_xor0 ^ u_CSAwallace_cska8_csa4_csa_component_fa3_and0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa4_and0 = u_CSAwallace_cska8_csa4_csa_component_fa4_xor0 & u_CSAwallace_cska8_csa4_csa_component_fa3_and0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa5_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa5_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa4_and0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa5_and0 = u_CSAwallace_cska8_csa4_csa_component_fa5_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa4_and0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa6_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa6_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa5_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa6_and0 = u_CSAwallace_cska8_csa4_csa_component_fa6_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa5_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa7_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa7_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa6_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa7_and0 = u_CSAwallace_cska8_csa4_csa_component_fa7_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa6_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa7_xor1 = u_CSAwallace_cska8_csa5_csa_component_fa7_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa6_and0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa7_and1 = u_CSAwallace_cska8_csa5_csa_component_fa7_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa6_and0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa7_or0 = u_CSAwallace_cska8_csa5_csa_component_fa7_and0 | u_CSAwallace_cska8_csa5_csa_component_fa7_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa8_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa8_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa8_and0 = u_CSAwallace_cska8_csa4_csa_component_fa8_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa8_xor1 = u_CSAwallace_cska8_csa5_csa_component_fa8_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa8_and1 = u_CSAwallace_cska8_csa5_csa_component_fa8_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa8_or0 = u_CSAwallace_cska8_csa5_csa_component_fa8_and0 | u_CSAwallace_cska8_csa5_csa_component_fa8_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa9_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa9_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa9_and0 = u_CSAwallace_cska8_csa4_csa_component_fa9_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa9_xor1 = u_CSAwallace_cska8_csa5_csa_component_fa9_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa9_and1 = u_CSAwallace_cska8_csa5_csa_component_fa9_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa9_or0 = u_CSAwallace_cska8_csa5_csa_component_fa9_and0 | u_CSAwallace_cska8_csa5_csa_component_fa9_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa10_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa10_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa10_and0 = u_CSAwallace_cska8_csa4_csa_component_fa10_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa10_xor1 = u_CSAwallace_cska8_csa5_csa_component_fa10_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa10_and1 = u_CSAwallace_cska8_csa5_csa_component_fa10_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa10_or0 = u_CSAwallace_cska8_csa5_csa_component_fa10_and0 | u_CSAwallace_cska8_csa5_csa_component_fa10_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa11_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa11_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa10_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa11_and0 = u_CSAwallace_cska8_csa4_csa_component_fa11_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa10_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa11_xor1 = u_CSAwallace_cska8_csa5_csa_component_fa11_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa10_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa11_and1 = u_CSAwallace_cska8_csa5_csa_component_fa11_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa10_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa11_or0 = u_CSAwallace_cska8_csa5_csa_component_fa11_and0 | u_CSAwallace_cska8_csa5_csa_component_fa11_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa12_xor0 = u_CSAwallace_cska8_csa4_csa_component_fa12_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa11_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa12_and0 = u_CSAwallace_cska8_csa4_csa_component_fa12_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa11_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa12_xor1 = u_CSAwallace_cska8_csa5_csa_component_fa12_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa11_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa12_and1 = u_CSAwallace_cska8_csa5_csa_component_fa12_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa11_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa12_or0 = u_CSAwallace_cska8_csa5_csa_component_fa12_and0 | u_CSAwallace_cska8_csa5_csa_component_fa12_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa13_xor0 = u_CSAwallace_cska8_csa3_csa_component_fa13_xor1 ^ u_CSAwallace_cska8_csa4_csa_component_fa12_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa13_and0 = u_CSAwallace_cska8_csa3_csa_component_fa13_xor1 & u_CSAwallace_cska8_csa4_csa_component_fa12_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa13_xor1 = u_CSAwallace_cska8_csa5_csa_component_fa13_xor0 ^ u_CSAwallace_cska8_csa3_csa_component_fa12_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa13_and1 = u_CSAwallace_cska8_csa5_csa_component_fa13_xor0 & u_CSAwallace_cska8_csa3_csa_component_fa12_or0;
  assign u_CSAwallace_cska8_csa5_csa_component_fa13_or0 = u_CSAwallace_cska8_csa5_csa_component_fa13_and0 | u_CSAwallace_cska8_csa5_csa_component_fa13_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa14_xor1 = u_CSAwallace_cska8_and_7_7 ^ u_CSAwallace_cska8_csa3_csa_component_fa13_and1;
  assign u_CSAwallace_cska8_csa5_csa_component_fa14_and1 = u_CSAwallace_cska8_and_7_7 & u_CSAwallace_cska8_csa3_csa_component_fa13_and1;
  assign u_CSAwallace_cska8_u_cska16_and_propagate00 = u_CSAwallace_cska8_and_0_0 & u_CSAwallace_cska8_csa2_csa_component_fa2_xor0;
  assign u_CSAwallace_cska8_u_cska16_and_propagate01 = u_CSAwallace_cska8_csa0_csa_component_fa1_xor0 & u_CSAwallace_cska8_csa4_csa_component_fa3_xor0;
  assign u_CSAwallace_cska8_u_cska16_and_propagate02 = u_CSAwallace_cska8_u_cska16_and_propagate00 & u_CSAwallace_cska8_u_cska16_and_propagate01;
  assign u_CSAwallace_cska8_u_cska16_mux2to10_not0 = ~u_CSAwallace_cska8_u_cska16_and_propagate02;
  assign u_CSAwallace_cska8_u_cska16_xor5 = u_CSAwallace_cska8_csa5_csa_component_fa5_xor0 ^ u_CSAwallace_cska8_csa5_csa_component_fa4_and0;
  assign u_CSAwallace_cska8_u_cska16_fa4_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa5_xor0 ^ u_CSAwallace_cska8_csa5_csa_component_fa4_and0;
  assign u_CSAwallace_cska8_u_cska16_fa4_and0 = u_CSAwallace_cska8_csa5_csa_component_fa5_xor0 & u_CSAwallace_cska8_csa5_csa_component_fa4_and0;
  assign u_CSAwallace_cska8_u_cska16_xor6 = u_CSAwallace_cska8_csa5_csa_component_fa6_xor0 ^ u_CSAwallace_cska8_csa5_csa_component_fa5_and0;
  assign u_CSAwallace_cska8_u_cska16_fa5_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa6_xor0 ^ u_CSAwallace_cska8_csa5_csa_component_fa5_and0;
  assign u_CSAwallace_cska8_u_cska16_fa5_and0 = u_CSAwallace_cska8_csa5_csa_component_fa6_xor0 & u_CSAwallace_cska8_csa5_csa_component_fa5_and0;
  assign u_CSAwallace_cska8_u_cska16_fa5_xor1 = u_CSAwallace_cska8_u_cska16_fa5_xor0 ^ u_CSAwallace_cska8_u_cska16_fa4_and0;
  assign u_CSAwallace_cska8_u_cska16_fa5_and1 = u_CSAwallace_cska8_u_cska16_fa5_xor0 & u_CSAwallace_cska8_u_cska16_fa4_and0;
  assign u_CSAwallace_cska8_u_cska16_fa5_or0 = u_CSAwallace_cska8_u_cska16_fa5_and0 | u_CSAwallace_cska8_u_cska16_fa5_and1;
  assign u_CSAwallace_cska8_u_cska16_xor7 = u_CSAwallace_cska8_csa5_csa_component_fa7_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa6_and0;
  assign u_CSAwallace_cska8_u_cska16_fa6_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa7_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa6_and0;
  assign u_CSAwallace_cska8_u_cska16_fa6_and0 = u_CSAwallace_cska8_csa5_csa_component_fa7_xor1 & u_CSAwallace_cska8_csa5_csa_component_fa6_and0;
  assign u_CSAwallace_cska8_u_cska16_fa6_xor1 = u_CSAwallace_cska8_u_cska16_fa6_xor0 ^ u_CSAwallace_cska8_u_cska16_fa5_or0;
  assign u_CSAwallace_cska8_u_cska16_fa6_and1 = u_CSAwallace_cska8_u_cska16_fa6_xor0 & u_CSAwallace_cska8_u_cska16_fa5_or0;
  assign u_CSAwallace_cska8_u_cska16_fa6_or0 = u_CSAwallace_cska8_u_cska16_fa6_and0 | u_CSAwallace_cska8_u_cska16_fa6_and1;
  assign u_CSAwallace_cska8_u_cska16_and_propagate13 = u_CSAwallace_cska8_csa5_csa_component_fa4_xor0 & u_CSAwallace_cska8_u_cska16_xor6;
  assign u_CSAwallace_cska8_u_cska16_and_propagate14 = u_CSAwallace_cska8_u_cska16_xor5 & u_CSAwallace_cska8_u_cska16_xor7;
  assign u_CSAwallace_cska8_u_cska16_and_propagate15 = u_CSAwallace_cska8_u_cska16_and_propagate13 & u_CSAwallace_cska8_u_cska16_and_propagate14;
  assign u_CSAwallace_cska8_u_cska16_mux2to11_not0 = ~u_CSAwallace_cska8_u_cska16_and_propagate15;
  assign u_CSAwallace_cska8_u_cska16_mux2to11_and1 = u_CSAwallace_cska8_u_cska16_fa6_or0 & u_CSAwallace_cska8_u_cska16_mux2to11_not0;
  assign u_CSAwallace_cska8_u_cska16_xor8 = u_CSAwallace_cska8_csa5_csa_component_fa8_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_u_cska16_fa7_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa8_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_u_cska16_fa7_and0 = u_CSAwallace_cska8_csa5_csa_component_fa8_xor1 & u_CSAwallace_cska8_csa5_csa_component_fa7_or0;
  assign u_CSAwallace_cska8_u_cska16_fa7_xor1 = u_CSAwallace_cska8_u_cska16_fa7_xor0 ^ u_CSAwallace_cska8_u_cska16_mux2to11_and1;
  assign u_CSAwallace_cska8_u_cska16_fa7_and1 = u_CSAwallace_cska8_u_cska16_fa7_xor0 & u_CSAwallace_cska8_u_cska16_mux2to11_and1;
  assign u_CSAwallace_cska8_u_cska16_fa7_or0 = u_CSAwallace_cska8_u_cska16_fa7_and0 | u_CSAwallace_cska8_u_cska16_fa7_and1;
  assign u_CSAwallace_cska8_u_cska16_xor9 = u_CSAwallace_cska8_csa5_csa_component_fa9_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_u_cska16_fa8_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa9_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_u_cska16_fa8_and0 = u_CSAwallace_cska8_csa5_csa_component_fa9_xor1 & u_CSAwallace_cska8_csa5_csa_component_fa8_or0;
  assign u_CSAwallace_cska8_u_cska16_fa8_xor1 = u_CSAwallace_cska8_u_cska16_fa8_xor0 ^ u_CSAwallace_cska8_u_cska16_fa7_or0;
  assign u_CSAwallace_cska8_u_cska16_fa8_and1 = u_CSAwallace_cska8_u_cska16_fa8_xor0 & u_CSAwallace_cska8_u_cska16_fa7_or0;
  assign u_CSAwallace_cska8_u_cska16_fa8_or0 = u_CSAwallace_cska8_u_cska16_fa8_and0 | u_CSAwallace_cska8_u_cska16_fa8_and1;
  assign u_CSAwallace_cska8_u_cska16_xor10 = u_CSAwallace_cska8_csa5_csa_component_fa10_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_u_cska16_fa9_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa10_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_u_cska16_fa9_and0 = u_CSAwallace_cska8_csa5_csa_component_fa10_xor1 & u_CSAwallace_cska8_csa5_csa_component_fa9_or0;
  assign u_CSAwallace_cska8_u_cska16_fa9_xor1 = u_CSAwallace_cska8_u_cska16_fa9_xor0 ^ u_CSAwallace_cska8_u_cska16_fa8_or0;
  assign u_CSAwallace_cska8_u_cska16_fa9_and1 = u_CSAwallace_cska8_u_cska16_fa9_xor0 & u_CSAwallace_cska8_u_cska16_fa8_or0;
  assign u_CSAwallace_cska8_u_cska16_fa9_or0 = u_CSAwallace_cska8_u_cska16_fa9_and0 | u_CSAwallace_cska8_u_cska16_fa9_and1;
  assign u_CSAwallace_cska8_u_cska16_xor11 = u_CSAwallace_cska8_csa5_csa_component_fa11_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa10_or0;
  assign u_CSAwallace_cska8_u_cska16_fa10_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa11_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa10_or0;
  assign u_CSAwallace_cska8_u_cska16_fa10_and0 = u_CSAwallace_cska8_csa5_csa_component_fa11_xor1 & u_CSAwallace_cska8_csa5_csa_component_fa10_or0;
  assign u_CSAwallace_cska8_u_cska16_fa10_xor1 = u_CSAwallace_cska8_u_cska16_fa10_xor0 ^ u_CSAwallace_cska8_u_cska16_fa9_or0;
  assign u_CSAwallace_cska8_u_cska16_fa10_and1 = u_CSAwallace_cska8_u_cska16_fa10_xor0 & u_CSAwallace_cska8_u_cska16_fa9_or0;
  assign u_CSAwallace_cska8_u_cska16_fa10_or0 = u_CSAwallace_cska8_u_cska16_fa10_and0 | u_CSAwallace_cska8_u_cska16_fa10_and1;
  assign u_CSAwallace_cska8_u_cska16_and_propagate26 = u_CSAwallace_cska8_u_cska16_xor8 & u_CSAwallace_cska8_u_cska16_xor10;
  assign u_CSAwallace_cska8_u_cska16_and_propagate27 = u_CSAwallace_cska8_u_cska16_xor9 & u_CSAwallace_cska8_u_cska16_xor11;
  assign u_CSAwallace_cska8_u_cska16_and_propagate28 = u_CSAwallace_cska8_u_cska16_and_propagate26 & u_CSAwallace_cska8_u_cska16_and_propagate27;
  assign u_CSAwallace_cska8_u_cska16_mux2to12_and0 = u_CSAwallace_cska8_u_cska16_mux2to11_and1 & u_CSAwallace_cska8_u_cska16_and_propagate28;
  assign u_CSAwallace_cska8_u_cska16_mux2to12_not0 = ~u_CSAwallace_cska8_u_cska16_and_propagate28;
  assign u_CSAwallace_cska8_u_cska16_mux2to12_and1 = u_CSAwallace_cska8_u_cska16_fa10_or0 & u_CSAwallace_cska8_u_cska16_mux2to12_not0;
  assign u_CSAwallace_cska8_u_cska16_mux2to12_xor0 = u_CSAwallace_cska8_u_cska16_mux2to12_and0 ^ u_CSAwallace_cska8_u_cska16_mux2to12_and1;
  assign u_CSAwallace_cska8_u_cska16_xor12 = u_CSAwallace_cska8_csa5_csa_component_fa12_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa11_or0;
  assign u_CSAwallace_cska8_u_cska16_fa11_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa12_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa11_or0;
  assign u_CSAwallace_cska8_u_cska16_fa11_and0 = u_CSAwallace_cska8_csa5_csa_component_fa12_xor1 & u_CSAwallace_cska8_csa5_csa_component_fa11_or0;
  assign u_CSAwallace_cska8_u_cska16_fa11_xor1 = u_CSAwallace_cska8_u_cska16_fa11_xor0 ^ u_CSAwallace_cska8_u_cska16_mux2to12_xor0;
  assign u_CSAwallace_cska8_u_cska16_fa11_and1 = u_CSAwallace_cska8_u_cska16_fa11_xor0 & u_CSAwallace_cska8_u_cska16_mux2to12_xor0;
  assign u_CSAwallace_cska8_u_cska16_fa11_or0 = u_CSAwallace_cska8_u_cska16_fa11_and0 | u_CSAwallace_cska8_u_cska16_fa11_and1;
  assign u_CSAwallace_cska8_u_cska16_xor13 = u_CSAwallace_cska8_csa5_csa_component_fa13_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa12_or0;
  assign u_CSAwallace_cska8_u_cska16_fa12_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa13_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa12_or0;
  assign u_CSAwallace_cska8_u_cska16_fa12_and0 = u_CSAwallace_cska8_csa5_csa_component_fa13_xor1 & u_CSAwallace_cska8_csa5_csa_component_fa12_or0;
  assign u_CSAwallace_cska8_u_cska16_fa12_xor1 = u_CSAwallace_cska8_u_cska16_fa12_xor0 ^ u_CSAwallace_cska8_u_cska16_fa11_or0;
  assign u_CSAwallace_cska8_u_cska16_fa12_and1 = u_CSAwallace_cska8_u_cska16_fa12_xor0 & u_CSAwallace_cska8_u_cska16_fa11_or0;
  assign u_CSAwallace_cska8_u_cska16_fa12_or0 = u_CSAwallace_cska8_u_cska16_fa12_and0 | u_CSAwallace_cska8_u_cska16_fa12_and1;
  assign u_CSAwallace_cska8_u_cska16_xor14 = u_CSAwallace_cska8_csa5_csa_component_fa14_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa13_or0;
  assign u_CSAwallace_cska8_u_cska16_fa13_xor0 = u_CSAwallace_cska8_csa5_csa_component_fa14_xor1 ^ u_CSAwallace_cska8_csa5_csa_component_fa13_or0;
  assign u_CSAwallace_cska8_u_cska16_fa13_and0 = u_CSAwallace_cska8_csa5_csa_component_fa14_xor1 & u_CSAwallace_cska8_csa5_csa_component_fa13_or0;
  assign u_CSAwallace_cska8_u_cska16_fa13_xor1 = u_CSAwallace_cska8_u_cska16_fa13_xor0 ^ u_CSAwallace_cska8_u_cska16_fa12_or0;
  assign u_CSAwallace_cska8_u_cska16_fa13_and1 = u_CSAwallace_cska8_u_cska16_fa13_xor0 & u_CSAwallace_cska8_u_cska16_fa12_or0;
  assign u_CSAwallace_cska8_u_cska16_fa13_or0 = u_CSAwallace_cska8_u_cska16_fa13_and0 | u_CSAwallace_cska8_u_cska16_fa13_and1;
  assign u_CSAwallace_cska8_u_cska16_fa14_xor1 = u_CSAwallace_cska8_csa5_csa_component_fa14_and1 ^ u_CSAwallace_cska8_u_cska16_fa13_or0;
  assign u_CSAwallace_cska8_u_cska16_fa14_and1 = u_CSAwallace_cska8_csa5_csa_component_fa14_and1 & u_CSAwallace_cska8_u_cska16_fa13_or0;
  assign u_CSAwallace_cska8_u_cska16_and_propagate39 = u_CSAwallace_cska8_u_cska16_xor12 & u_CSAwallace_cska8_u_cska16_xor14;
  assign u_CSAwallace_cska8_u_cska16_and_propagate310 = u_CSAwallace_cska8_u_cska16_xor13 & u_CSAwallace_cska8_csa5_csa_component_fa14_and1;
  assign u_CSAwallace_cska8_u_cska16_and_propagate311 = u_CSAwallace_cska8_u_cska16_and_propagate39 & u_CSAwallace_cska8_u_cska16_and_propagate310;
  assign u_CSAwallace_cska8_u_cska16_mux2to13_and0 = u_CSAwallace_cska8_u_cska16_mux2to12_xor0 & u_CSAwallace_cska8_u_cska16_and_propagate311;
  assign u_CSAwallace_cska8_u_cska16_mux2to13_not0 = ~u_CSAwallace_cska8_u_cska16_and_propagate311;
  assign u_CSAwallace_cska8_u_cska16_mux2to13_and1 = u_CSAwallace_cska8_u_cska16_fa14_and1 & u_CSAwallace_cska8_u_cska16_mux2to13_not0;
  assign u_CSAwallace_cska8_u_cska16_mux2to13_xor0 = u_CSAwallace_cska8_u_cska16_mux2to13_and0 ^ u_CSAwallace_cska8_u_cska16_mux2to13_and1;

  assign u_CSAwallace_cska8_out[0] = u_CSAwallace_cska8_and_0_0;
  assign u_CSAwallace_cska8_out[1] = u_CSAwallace_cska8_csa0_csa_component_fa1_xor0;
  assign u_CSAwallace_cska8_out[2] = u_CSAwallace_cska8_csa2_csa_component_fa2_xor0;
  assign u_CSAwallace_cska8_out[3] = u_CSAwallace_cska8_csa4_csa_component_fa3_xor0;
  assign u_CSAwallace_cska8_out[4] = u_CSAwallace_cska8_csa5_csa_component_fa4_xor0;
  assign u_CSAwallace_cska8_out[5] = u_CSAwallace_cska8_u_cska16_fa4_xor0;
  assign u_CSAwallace_cska8_out[6] = u_CSAwallace_cska8_u_cska16_fa5_xor1;
  assign u_CSAwallace_cska8_out[7] = u_CSAwallace_cska8_u_cska16_fa6_xor1;
  assign u_CSAwallace_cska8_out[8] = u_CSAwallace_cska8_u_cska16_fa7_xor1;
  assign u_CSAwallace_cska8_out[9] = u_CSAwallace_cska8_u_cska16_fa8_xor1;
  assign u_CSAwallace_cska8_out[10] = u_CSAwallace_cska8_u_cska16_fa9_xor1;
  assign u_CSAwallace_cska8_out[11] = u_CSAwallace_cska8_u_cska16_fa10_xor1;
  assign u_CSAwallace_cska8_out[12] = u_CSAwallace_cska8_u_cska16_fa11_xor1;
  assign u_CSAwallace_cska8_out[13] = u_CSAwallace_cska8_u_cska16_fa12_xor1;
  assign u_CSAwallace_cska8_out[14] = u_CSAwallace_cska8_u_cska16_fa13_xor1;
  assign u_CSAwallace_cska8_out[15] = u_CSAwallace_cska8_u_cska16_fa14_xor1;
endmodule