module u_CSAwallace_cla8(input [7:0] a, input [7:0] b, output [15:0] u_CSAwallace_cla8_out);
  wire u_CSAwallace_cla8_and_0_0;
  wire u_CSAwallace_cla8_and_1_0;
  wire u_CSAwallace_cla8_and_2_0;
  wire u_CSAwallace_cla8_and_3_0;
  wire u_CSAwallace_cla8_and_4_0;
  wire u_CSAwallace_cla8_and_5_0;
  wire u_CSAwallace_cla8_and_6_0;
  wire u_CSAwallace_cla8_and_7_0;
  wire u_CSAwallace_cla8_and_0_1;
  wire u_CSAwallace_cla8_and_1_1;
  wire u_CSAwallace_cla8_and_2_1;
  wire u_CSAwallace_cla8_and_3_1;
  wire u_CSAwallace_cla8_and_4_1;
  wire u_CSAwallace_cla8_and_5_1;
  wire u_CSAwallace_cla8_and_6_1;
  wire u_CSAwallace_cla8_and_7_1;
  wire u_CSAwallace_cla8_and_0_2;
  wire u_CSAwallace_cla8_and_1_2;
  wire u_CSAwallace_cla8_and_2_2;
  wire u_CSAwallace_cla8_and_3_2;
  wire u_CSAwallace_cla8_and_4_2;
  wire u_CSAwallace_cla8_and_5_2;
  wire u_CSAwallace_cla8_and_6_2;
  wire u_CSAwallace_cla8_and_7_2;
  wire u_CSAwallace_cla8_and_0_3;
  wire u_CSAwallace_cla8_and_1_3;
  wire u_CSAwallace_cla8_and_2_3;
  wire u_CSAwallace_cla8_and_3_3;
  wire u_CSAwallace_cla8_and_4_3;
  wire u_CSAwallace_cla8_and_5_3;
  wire u_CSAwallace_cla8_and_6_3;
  wire u_CSAwallace_cla8_and_7_3;
  wire u_CSAwallace_cla8_and_0_4;
  wire u_CSAwallace_cla8_and_1_4;
  wire u_CSAwallace_cla8_and_2_4;
  wire u_CSAwallace_cla8_and_3_4;
  wire u_CSAwallace_cla8_and_4_4;
  wire u_CSAwallace_cla8_and_5_4;
  wire u_CSAwallace_cla8_and_6_4;
  wire u_CSAwallace_cla8_and_7_4;
  wire u_CSAwallace_cla8_and_0_5;
  wire u_CSAwallace_cla8_and_1_5;
  wire u_CSAwallace_cla8_and_2_5;
  wire u_CSAwallace_cla8_and_3_5;
  wire u_CSAwallace_cla8_and_4_5;
  wire u_CSAwallace_cla8_and_5_5;
  wire u_CSAwallace_cla8_and_6_5;
  wire u_CSAwallace_cla8_and_7_5;
  wire u_CSAwallace_cla8_and_0_6;
  wire u_CSAwallace_cla8_and_1_6;
  wire u_CSAwallace_cla8_and_2_6;
  wire u_CSAwallace_cla8_and_3_6;
  wire u_CSAwallace_cla8_and_4_6;
  wire u_CSAwallace_cla8_and_5_6;
  wire u_CSAwallace_cla8_and_6_6;
  wire u_CSAwallace_cla8_and_7_6;
  wire u_CSAwallace_cla8_and_0_7;
  wire u_CSAwallace_cla8_and_1_7;
  wire u_CSAwallace_cla8_and_2_7;
  wire u_CSAwallace_cla8_and_3_7;
  wire u_CSAwallace_cla8_and_4_7;
  wire u_CSAwallace_cla8_and_5_7;
  wire u_CSAwallace_cla8_and_6_7;
  wire u_CSAwallace_cla8_and_7_7;
  wire u_CSAwallace_cla8_csa0_csa_component_fa1_xor0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa1_and0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa2_xor0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa2_and0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa2_xor1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa2_and1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa2_or0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa3_xor0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa3_and0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa3_xor1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa3_and1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa3_or0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa4_xor0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa4_and0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa4_xor1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa4_and1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa4_or0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa5_xor0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa5_and0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa5_xor1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa5_and1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa5_or0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa6_xor0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa6_and0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa6_xor1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa6_and1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa6_or0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa7_xor0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa7_and0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa7_xor1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa7_and1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa7_or0;
  wire u_CSAwallace_cla8_csa0_csa_component_fa8_xor1;
  wire u_CSAwallace_cla8_csa0_csa_component_fa8_and1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa4_xor0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa4_and0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa5_xor0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa5_and0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa5_xor1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa5_and1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa5_or0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa6_xor0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa6_and0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa6_xor1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa6_and1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa6_or0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa7_xor0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa7_and0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa7_xor1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa7_and1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa7_or0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa8_xor0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa8_and0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa8_xor1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa8_and1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa8_or0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa9_xor0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa9_and0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa9_xor1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa9_and1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa9_or0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa10_xor0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa10_and0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa10_xor1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa10_and1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa10_or0;
  wire u_CSAwallace_cla8_csa1_csa_component_fa11_xor1;
  wire u_CSAwallace_cla8_csa1_csa_component_fa11_and1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa2_xor0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa2_and0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa3_xor0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa3_and0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa3_xor1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa3_and1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa3_or0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa4_xor0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa4_and0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa4_xor1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa4_and1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa4_or0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa5_xor0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa5_and0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa5_xor1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa5_and1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa5_or0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa6_xor0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa6_and0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa6_xor1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa6_and1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa6_or0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa7_xor0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa7_and0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa7_xor1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa7_and1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa7_or0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa8_xor0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa8_and0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa8_xor1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa8_and1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa8_or0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa9_xor0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa9_and0;
  wire u_CSAwallace_cla8_csa2_csa_component_fa9_xor1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa9_and1;
  wire u_CSAwallace_cla8_csa2_csa_component_fa9_or0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa6_xor0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa6_and0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa7_xor0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa7_and0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa7_xor1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa7_and1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa7_or0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa8_xor0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa8_and0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa8_xor1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa8_and1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa8_or0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa9_xor0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa9_and0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa9_xor1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa9_and1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa9_or0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa10_xor0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa10_and0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa10_xor1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa10_and1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa10_or0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa11_xor0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa11_and0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa11_xor1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa11_and1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa11_or0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa12_xor0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa12_and0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa12_xor1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa12_and1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa12_or0;
  wire u_CSAwallace_cla8_csa3_csa_component_fa13_xor1;
  wire u_CSAwallace_cla8_csa3_csa_component_fa13_and1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa3_xor0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa3_and0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa4_xor0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa4_and0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa5_xor0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa5_and0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa5_xor1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa5_and1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa5_or0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa6_xor0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa6_and0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa6_xor1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa6_and1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa6_or0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa7_xor0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa7_and0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa7_xor1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa7_and1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa7_or0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa8_xor0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa8_and0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa8_xor1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa8_and1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa8_or0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa9_xor0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa9_and0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa9_xor1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa9_and1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa9_or0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa10_xor0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa10_and0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa10_xor1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa10_and1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa10_or0;
  wire u_CSAwallace_cla8_csa4_csa_component_fa11_xor1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa11_and1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa12_xor1;
  wire u_CSAwallace_cla8_csa4_csa_component_fa12_and1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa4_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa4_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa5_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa5_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa6_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa6_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa7_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa7_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa7_xor1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa7_and1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa7_or0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa8_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa8_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa8_xor1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa8_and1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa8_or0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa9_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa9_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa9_xor1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa9_and1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa9_or0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa10_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa10_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa10_xor1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa10_and1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa10_or0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa11_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa11_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa11_xor1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa11_and1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa11_or0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa12_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa12_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa12_xor1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa12_and1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa12_or0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa13_xor0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa13_and0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa13_xor1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa13_and1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa13_or0;
  wire u_CSAwallace_cla8_csa5_csa_component_fa14_xor1;
  wire u_CSAwallace_cla8_csa5_csa_component_fa14_and1;
  wire u_CSAwallace_cla8_u_cla16_and0;
  wire u_CSAwallace_cla8_u_cla16_and1;
  wire u_CSAwallace_cla8_u_cla16_and2;
  wire u_CSAwallace_cla8_u_cla16_pg_logic5_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic5_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic5_xor0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic6_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic6_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic6_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor6;
  wire u_CSAwallace_cla8_u_cla16_and3;
  wire u_CSAwallace_cla8_u_cla16_and4;
  wire u_CSAwallace_cla8_u_cla16_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic7_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic7_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic7_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor7;
  wire u_CSAwallace_cla8_u_cla16_and5;
  wire u_CSAwallace_cla8_u_cla16_and6;
  wire u_CSAwallace_cla8_u_cla16_and7;
  wire u_CSAwallace_cla8_u_cla16_and8;
  wire u_CSAwallace_cla8_u_cla16_and9;
  wire u_CSAwallace_cla8_u_cla16_or1;
  wire u_CSAwallace_cla8_u_cla16_or2;
  wire u_CSAwallace_cla8_u_cla16_pg_logic8_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic8_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic8_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor8;
  wire u_CSAwallace_cla8_u_cla16_and10;
  wire u_CSAwallace_cla8_u_cla16_or3;
  wire u_CSAwallace_cla8_u_cla16_pg_logic9_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic9_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic9_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor9;
  wire u_CSAwallace_cla8_u_cla16_and11;
  wire u_CSAwallace_cla8_u_cla16_and12;
  wire u_CSAwallace_cla8_u_cla16_and13;
  wire u_CSAwallace_cla8_u_cla16_or4;
  wire u_CSAwallace_cla8_u_cla16_or5;
  wire u_CSAwallace_cla8_u_cla16_pg_logic10_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic10_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic10_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor10;
  wire u_CSAwallace_cla8_u_cla16_and14;
  wire u_CSAwallace_cla8_u_cla16_and15;
  wire u_CSAwallace_cla8_u_cla16_and16;
  wire u_CSAwallace_cla8_u_cla16_and17;
  wire u_CSAwallace_cla8_u_cla16_and18;
  wire u_CSAwallace_cla8_u_cla16_and19;
  wire u_CSAwallace_cla8_u_cla16_or6;
  wire u_CSAwallace_cla8_u_cla16_or7;
  wire u_CSAwallace_cla8_u_cla16_or8;
  wire u_CSAwallace_cla8_u_cla16_pg_logic11_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic11_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic11_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor11;
  wire u_CSAwallace_cla8_u_cla16_and20;
  wire u_CSAwallace_cla8_u_cla16_and21;
  wire u_CSAwallace_cla8_u_cla16_and22;
  wire u_CSAwallace_cla8_u_cla16_and23;
  wire u_CSAwallace_cla8_u_cla16_and24;
  wire u_CSAwallace_cla8_u_cla16_and25;
  wire u_CSAwallace_cla8_u_cla16_and26;
  wire u_CSAwallace_cla8_u_cla16_and27;
  wire u_CSAwallace_cla8_u_cla16_and28;
  wire u_CSAwallace_cla8_u_cla16_and29;
  wire u_CSAwallace_cla8_u_cla16_or9;
  wire u_CSAwallace_cla8_u_cla16_or10;
  wire u_CSAwallace_cla8_u_cla16_or11;
  wire u_CSAwallace_cla8_u_cla16_or12;
  wire u_CSAwallace_cla8_u_cla16_pg_logic12_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic12_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic12_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor12;
  wire u_CSAwallace_cla8_u_cla16_and30;
  wire u_CSAwallace_cla8_u_cla16_or13;
  wire u_CSAwallace_cla8_u_cla16_pg_logic13_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic13_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic13_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor13;
  wire u_CSAwallace_cla8_u_cla16_and31;
  wire u_CSAwallace_cla8_u_cla16_and32;
  wire u_CSAwallace_cla8_u_cla16_and33;
  wire u_CSAwallace_cla8_u_cla16_or14;
  wire u_CSAwallace_cla8_u_cla16_or15;
  wire u_CSAwallace_cla8_u_cla16_pg_logic14_or0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic14_and0;
  wire u_CSAwallace_cla8_u_cla16_pg_logic14_xor0;
  wire u_CSAwallace_cla8_u_cla16_xor14;
  wire u_CSAwallace_cla8_u_cla16_and34;
  wire u_CSAwallace_cla8_u_cla16_and35;
  wire u_CSAwallace_cla8_u_cla16_and36;
  wire u_CSAwallace_cla8_u_cla16_and37;
  wire u_CSAwallace_cla8_u_cla16_and38;
  wire u_CSAwallace_cla8_u_cla16_and39;
  wire u_CSAwallace_cla8_u_cla16_or16;
  wire u_CSAwallace_cla8_u_cla16_or17;
  wire u_CSAwallace_cla8_u_cla16_or18;
  wire u_CSAwallace_cla8_u_cla16_xor15;
  wire u_CSAwallace_cla8_u_cla16_and40;
  wire u_CSAwallace_cla8_u_cla16_and41;
  wire u_CSAwallace_cla8_u_cla16_and42;
  wire u_CSAwallace_cla8_u_cla16_and43;
  wire u_CSAwallace_cla8_u_cla16_and44;
  wire u_CSAwallace_cla8_u_cla16_and45;
  wire u_CSAwallace_cla8_u_cla16_and46;
  wire u_CSAwallace_cla8_u_cla16_and47;
  wire u_CSAwallace_cla8_u_cla16_and48;
  wire u_CSAwallace_cla8_u_cla16_and49;
  wire u_CSAwallace_cla8_u_cla16_or19;
  wire u_CSAwallace_cla8_u_cla16_or20;
  wire u_CSAwallace_cla8_u_cla16_or21;

  assign u_CSAwallace_cla8_and_0_0 = a[0] & b[0];
  assign u_CSAwallace_cla8_and_1_0 = a[1] & b[0];
  assign u_CSAwallace_cla8_and_2_0 = a[2] & b[0];
  assign u_CSAwallace_cla8_and_3_0 = a[3] & b[0];
  assign u_CSAwallace_cla8_and_4_0 = a[4] & b[0];
  assign u_CSAwallace_cla8_and_5_0 = a[5] & b[0];
  assign u_CSAwallace_cla8_and_6_0 = a[6] & b[0];
  assign u_CSAwallace_cla8_and_7_0 = a[7] & b[0];
  assign u_CSAwallace_cla8_and_0_1 = a[0] & b[1];
  assign u_CSAwallace_cla8_and_1_1 = a[1] & b[1];
  assign u_CSAwallace_cla8_and_2_1 = a[2] & b[1];
  assign u_CSAwallace_cla8_and_3_1 = a[3] & b[1];
  assign u_CSAwallace_cla8_and_4_1 = a[4] & b[1];
  assign u_CSAwallace_cla8_and_5_1 = a[5] & b[1];
  assign u_CSAwallace_cla8_and_6_1 = a[6] & b[1];
  assign u_CSAwallace_cla8_and_7_1 = a[7] & b[1];
  assign u_CSAwallace_cla8_and_0_2 = a[0] & b[2];
  assign u_CSAwallace_cla8_and_1_2 = a[1] & b[2];
  assign u_CSAwallace_cla8_and_2_2 = a[2] & b[2];
  assign u_CSAwallace_cla8_and_3_2 = a[3] & b[2];
  assign u_CSAwallace_cla8_and_4_2 = a[4] & b[2];
  assign u_CSAwallace_cla8_and_5_2 = a[5] & b[2];
  assign u_CSAwallace_cla8_and_6_2 = a[6] & b[2];
  assign u_CSAwallace_cla8_and_7_2 = a[7] & b[2];
  assign u_CSAwallace_cla8_and_0_3 = a[0] & b[3];
  assign u_CSAwallace_cla8_and_1_3 = a[1] & b[3];
  assign u_CSAwallace_cla8_and_2_3 = a[2] & b[3];
  assign u_CSAwallace_cla8_and_3_3 = a[3] & b[3];
  assign u_CSAwallace_cla8_and_4_3 = a[4] & b[3];
  assign u_CSAwallace_cla8_and_5_3 = a[5] & b[3];
  assign u_CSAwallace_cla8_and_6_3 = a[6] & b[3];
  assign u_CSAwallace_cla8_and_7_3 = a[7] & b[3];
  assign u_CSAwallace_cla8_and_0_4 = a[0] & b[4];
  assign u_CSAwallace_cla8_and_1_4 = a[1] & b[4];
  assign u_CSAwallace_cla8_and_2_4 = a[2] & b[4];
  assign u_CSAwallace_cla8_and_3_4 = a[3] & b[4];
  assign u_CSAwallace_cla8_and_4_4 = a[4] & b[4];
  assign u_CSAwallace_cla8_and_5_4 = a[5] & b[4];
  assign u_CSAwallace_cla8_and_6_4 = a[6] & b[4];
  assign u_CSAwallace_cla8_and_7_4 = a[7] & b[4];
  assign u_CSAwallace_cla8_and_0_5 = a[0] & b[5];
  assign u_CSAwallace_cla8_and_1_5 = a[1] & b[5];
  assign u_CSAwallace_cla8_and_2_5 = a[2] & b[5];
  assign u_CSAwallace_cla8_and_3_5 = a[3] & b[5];
  assign u_CSAwallace_cla8_and_4_5 = a[4] & b[5];
  assign u_CSAwallace_cla8_and_5_5 = a[5] & b[5];
  assign u_CSAwallace_cla8_and_6_5 = a[6] & b[5];
  assign u_CSAwallace_cla8_and_7_5 = a[7] & b[5];
  assign u_CSAwallace_cla8_and_0_6 = a[0] & b[6];
  assign u_CSAwallace_cla8_and_1_6 = a[1] & b[6];
  assign u_CSAwallace_cla8_and_2_6 = a[2] & b[6];
  assign u_CSAwallace_cla8_and_3_6 = a[3] & b[6];
  assign u_CSAwallace_cla8_and_4_6 = a[4] & b[6];
  assign u_CSAwallace_cla8_and_5_6 = a[5] & b[6];
  assign u_CSAwallace_cla8_and_6_6 = a[6] & b[6];
  assign u_CSAwallace_cla8_and_7_6 = a[7] & b[6];
  assign u_CSAwallace_cla8_and_0_7 = a[0] & b[7];
  assign u_CSAwallace_cla8_and_1_7 = a[1] & b[7];
  assign u_CSAwallace_cla8_and_2_7 = a[2] & b[7];
  assign u_CSAwallace_cla8_and_3_7 = a[3] & b[7];
  assign u_CSAwallace_cla8_and_4_7 = a[4] & b[7];
  assign u_CSAwallace_cla8_and_5_7 = a[5] & b[7];
  assign u_CSAwallace_cla8_and_6_7 = a[6] & b[7];
  assign u_CSAwallace_cla8_and_7_7 = a[7] & b[7];
  assign u_CSAwallace_cla8_csa0_csa_component_fa1_xor0 = u_CSAwallace_cla8_and_1_0 ^ u_CSAwallace_cla8_and_0_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa1_and0 = u_CSAwallace_cla8_and_1_0 & u_CSAwallace_cla8_and_0_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa2_xor0 = u_CSAwallace_cla8_and_2_0 ^ u_CSAwallace_cla8_and_1_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa2_and0 = u_CSAwallace_cla8_and_2_0 & u_CSAwallace_cla8_and_1_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa2_xor1 = u_CSAwallace_cla8_csa0_csa_component_fa2_xor0 ^ u_CSAwallace_cla8_and_0_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa2_and1 = u_CSAwallace_cla8_csa0_csa_component_fa2_xor0 & u_CSAwallace_cla8_and_0_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa2_or0 = u_CSAwallace_cla8_csa0_csa_component_fa2_and0 | u_CSAwallace_cla8_csa0_csa_component_fa2_and1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa3_xor0 = u_CSAwallace_cla8_and_3_0 ^ u_CSAwallace_cla8_and_2_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa3_and0 = u_CSAwallace_cla8_and_3_0 & u_CSAwallace_cla8_and_2_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa3_xor1 = u_CSAwallace_cla8_csa0_csa_component_fa3_xor0 ^ u_CSAwallace_cla8_and_1_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa3_and1 = u_CSAwallace_cla8_csa0_csa_component_fa3_xor0 & u_CSAwallace_cla8_and_1_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa3_or0 = u_CSAwallace_cla8_csa0_csa_component_fa3_and0 | u_CSAwallace_cla8_csa0_csa_component_fa3_and1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa4_xor0 = u_CSAwallace_cla8_and_4_0 ^ u_CSAwallace_cla8_and_3_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa4_and0 = u_CSAwallace_cla8_and_4_0 & u_CSAwallace_cla8_and_3_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa4_xor1 = u_CSAwallace_cla8_csa0_csa_component_fa4_xor0 ^ u_CSAwallace_cla8_and_2_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa4_and1 = u_CSAwallace_cla8_csa0_csa_component_fa4_xor0 & u_CSAwallace_cla8_and_2_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa4_or0 = u_CSAwallace_cla8_csa0_csa_component_fa4_and0 | u_CSAwallace_cla8_csa0_csa_component_fa4_and1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa5_xor0 = u_CSAwallace_cla8_and_5_0 ^ u_CSAwallace_cla8_and_4_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa5_and0 = u_CSAwallace_cla8_and_5_0 & u_CSAwallace_cla8_and_4_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa5_xor1 = u_CSAwallace_cla8_csa0_csa_component_fa5_xor0 ^ u_CSAwallace_cla8_and_3_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa5_and1 = u_CSAwallace_cla8_csa0_csa_component_fa5_xor0 & u_CSAwallace_cla8_and_3_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa5_or0 = u_CSAwallace_cla8_csa0_csa_component_fa5_and0 | u_CSAwallace_cla8_csa0_csa_component_fa5_and1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa6_xor0 = u_CSAwallace_cla8_and_6_0 ^ u_CSAwallace_cla8_and_5_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa6_and0 = u_CSAwallace_cla8_and_6_0 & u_CSAwallace_cla8_and_5_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa6_xor1 = u_CSAwallace_cla8_csa0_csa_component_fa6_xor0 ^ u_CSAwallace_cla8_and_4_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa6_and1 = u_CSAwallace_cla8_csa0_csa_component_fa6_xor0 & u_CSAwallace_cla8_and_4_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa6_or0 = u_CSAwallace_cla8_csa0_csa_component_fa6_and0 | u_CSAwallace_cla8_csa0_csa_component_fa6_and1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa7_xor0 = u_CSAwallace_cla8_and_7_0 ^ u_CSAwallace_cla8_and_6_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa7_and0 = u_CSAwallace_cla8_and_7_0 & u_CSAwallace_cla8_and_6_1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa7_xor1 = u_CSAwallace_cla8_csa0_csa_component_fa7_xor0 ^ u_CSAwallace_cla8_and_5_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa7_and1 = u_CSAwallace_cla8_csa0_csa_component_fa7_xor0 & u_CSAwallace_cla8_and_5_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa7_or0 = u_CSAwallace_cla8_csa0_csa_component_fa7_and0 | u_CSAwallace_cla8_csa0_csa_component_fa7_and1;
  assign u_CSAwallace_cla8_csa0_csa_component_fa8_xor1 = u_CSAwallace_cla8_and_7_1 ^ u_CSAwallace_cla8_and_6_2;
  assign u_CSAwallace_cla8_csa0_csa_component_fa8_and1 = u_CSAwallace_cla8_and_7_1 & u_CSAwallace_cla8_and_6_2;
  assign u_CSAwallace_cla8_csa1_csa_component_fa4_xor0 = u_CSAwallace_cla8_and_1_3 ^ u_CSAwallace_cla8_and_0_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa4_and0 = u_CSAwallace_cla8_and_1_3 & u_CSAwallace_cla8_and_0_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa5_xor0 = u_CSAwallace_cla8_and_2_3 ^ u_CSAwallace_cla8_and_1_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa5_and0 = u_CSAwallace_cla8_and_2_3 & u_CSAwallace_cla8_and_1_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa5_xor1 = u_CSAwallace_cla8_csa1_csa_component_fa5_xor0 ^ u_CSAwallace_cla8_and_0_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa5_and1 = u_CSAwallace_cla8_csa1_csa_component_fa5_xor0 & u_CSAwallace_cla8_and_0_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa5_or0 = u_CSAwallace_cla8_csa1_csa_component_fa5_and0 | u_CSAwallace_cla8_csa1_csa_component_fa5_and1;
  assign u_CSAwallace_cla8_csa1_csa_component_fa6_xor0 = u_CSAwallace_cla8_and_3_3 ^ u_CSAwallace_cla8_and_2_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa6_and0 = u_CSAwallace_cla8_and_3_3 & u_CSAwallace_cla8_and_2_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa6_xor1 = u_CSAwallace_cla8_csa1_csa_component_fa6_xor0 ^ u_CSAwallace_cla8_and_1_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa6_and1 = u_CSAwallace_cla8_csa1_csa_component_fa6_xor0 & u_CSAwallace_cla8_and_1_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa6_or0 = u_CSAwallace_cla8_csa1_csa_component_fa6_and0 | u_CSAwallace_cla8_csa1_csa_component_fa6_and1;
  assign u_CSAwallace_cla8_csa1_csa_component_fa7_xor0 = u_CSAwallace_cla8_and_4_3 ^ u_CSAwallace_cla8_and_3_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa7_and0 = u_CSAwallace_cla8_and_4_3 & u_CSAwallace_cla8_and_3_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa7_xor1 = u_CSAwallace_cla8_csa1_csa_component_fa7_xor0 ^ u_CSAwallace_cla8_and_2_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa7_and1 = u_CSAwallace_cla8_csa1_csa_component_fa7_xor0 & u_CSAwallace_cla8_and_2_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa7_or0 = u_CSAwallace_cla8_csa1_csa_component_fa7_and0 | u_CSAwallace_cla8_csa1_csa_component_fa7_and1;
  assign u_CSAwallace_cla8_csa1_csa_component_fa8_xor0 = u_CSAwallace_cla8_and_5_3 ^ u_CSAwallace_cla8_and_4_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa8_and0 = u_CSAwallace_cla8_and_5_3 & u_CSAwallace_cla8_and_4_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa8_xor1 = u_CSAwallace_cla8_csa1_csa_component_fa8_xor0 ^ u_CSAwallace_cla8_and_3_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa8_and1 = u_CSAwallace_cla8_csa1_csa_component_fa8_xor0 & u_CSAwallace_cla8_and_3_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa8_or0 = u_CSAwallace_cla8_csa1_csa_component_fa8_and0 | u_CSAwallace_cla8_csa1_csa_component_fa8_and1;
  assign u_CSAwallace_cla8_csa1_csa_component_fa9_xor0 = u_CSAwallace_cla8_and_6_3 ^ u_CSAwallace_cla8_and_5_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa9_and0 = u_CSAwallace_cla8_and_6_3 & u_CSAwallace_cla8_and_5_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa9_xor1 = u_CSAwallace_cla8_csa1_csa_component_fa9_xor0 ^ u_CSAwallace_cla8_and_4_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa9_and1 = u_CSAwallace_cla8_csa1_csa_component_fa9_xor0 & u_CSAwallace_cla8_and_4_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa9_or0 = u_CSAwallace_cla8_csa1_csa_component_fa9_and0 | u_CSAwallace_cla8_csa1_csa_component_fa9_and1;
  assign u_CSAwallace_cla8_csa1_csa_component_fa10_xor0 = u_CSAwallace_cla8_and_7_3 ^ u_CSAwallace_cla8_and_6_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa10_and0 = u_CSAwallace_cla8_and_7_3 & u_CSAwallace_cla8_and_6_4;
  assign u_CSAwallace_cla8_csa1_csa_component_fa10_xor1 = u_CSAwallace_cla8_csa1_csa_component_fa10_xor0 ^ u_CSAwallace_cla8_and_5_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa10_and1 = u_CSAwallace_cla8_csa1_csa_component_fa10_xor0 & u_CSAwallace_cla8_and_5_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa10_or0 = u_CSAwallace_cla8_csa1_csa_component_fa10_and0 | u_CSAwallace_cla8_csa1_csa_component_fa10_and1;
  assign u_CSAwallace_cla8_csa1_csa_component_fa11_xor1 = u_CSAwallace_cla8_and_7_4 ^ u_CSAwallace_cla8_and_6_5;
  assign u_CSAwallace_cla8_csa1_csa_component_fa11_and1 = u_CSAwallace_cla8_and_7_4 & u_CSAwallace_cla8_and_6_5;
  assign u_CSAwallace_cla8_csa2_csa_component_fa2_xor0 = u_CSAwallace_cla8_csa0_csa_component_fa2_xor1 ^ u_CSAwallace_cla8_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa2_and0 = u_CSAwallace_cla8_csa0_csa_component_fa2_xor1 & u_CSAwallace_cla8_csa0_csa_component_fa1_and0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa3_xor0 = u_CSAwallace_cla8_csa0_csa_component_fa3_xor1 ^ u_CSAwallace_cla8_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa3_and0 = u_CSAwallace_cla8_csa0_csa_component_fa3_xor1 & u_CSAwallace_cla8_csa0_csa_component_fa2_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa3_xor1 = u_CSAwallace_cla8_csa2_csa_component_fa3_xor0 ^ u_CSAwallace_cla8_and_0_3;
  assign u_CSAwallace_cla8_csa2_csa_component_fa3_and1 = u_CSAwallace_cla8_csa2_csa_component_fa3_xor0 & u_CSAwallace_cla8_and_0_3;
  assign u_CSAwallace_cla8_csa2_csa_component_fa3_or0 = u_CSAwallace_cla8_csa2_csa_component_fa3_and0 | u_CSAwallace_cla8_csa2_csa_component_fa3_and1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa4_xor0 = u_CSAwallace_cla8_csa0_csa_component_fa4_xor1 ^ u_CSAwallace_cla8_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa4_and0 = u_CSAwallace_cla8_csa0_csa_component_fa4_xor1 & u_CSAwallace_cla8_csa0_csa_component_fa3_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa4_xor1 = u_CSAwallace_cla8_csa2_csa_component_fa4_xor0 ^ u_CSAwallace_cla8_csa1_csa_component_fa4_xor0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa4_and1 = u_CSAwallace_cla8_csa2_csa_component_fa4_xor0 & u_CSAwallace_cla8_csa1_csa_component_fa4_xor0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa4_or0 = u_CSAwallace_cla8_csa2_csa_component_fa4_and0 | u_CSAwallace_cla8_csa2_csa_component_fa4_and1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa5_xor0 = u_CSAwallace_cla8_csa0_csa_component_fa5_xor1 ^ u_CSAwallace_cla8_csa0_csa_component_fa4_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa5_and0 = u_CSAwallace_cla8_csa0_csa_component_fa5_xor1 & u_CSAwallace_cla8_csa0_csa_component_fa4_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa5_xor1 = u_CSAwallace_cla8_csa2_csa_component_fa5_xor0 ^ u_CSAwallace_cla8_csa1_csa_component_fa5_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa5_and1 = u_CSAwallace_cla8_csa2_csa_component_fa5_xor0 & u_CSAwallace_cla8_csa1_csa_component_fa5_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa5_or0 = u_CSAwallace_cla8_csa2_csa_component_fa5_and0 | u_CSAwallace_cla8_csa2_csa_component_fa5_and1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa6_xor0 = u_CSAwallace_cla8_csa0_csa_component_fa6_xor1 ^ u_CSAwallace_cla8_csa0_csa_component_fa5_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa6_and0 = u_CSAwallace_cla8_csa0_csa_component_fa6_xor1 & u_CSAwallace_cla8_csa0_csa_component_fa5_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa6_xor1 = u_CSAwallace_cla8_csa2_csa_component_fa6_xor0 ^ u_CSAwallace_cla8_csa1_csa_component_fa6_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa6_and1 = u_CSAwallace_cla8_csa2_csa_component_fa6_xor0 & u_CSAwallace_cla8_csa1_csa_component_fa6_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa6_or0 = u_CSAwallace_cla8_csa2_csa_component_fa6_and0 | u_CSAwallace_cla8_csa2_csa_component_fa6_and1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa7_xor0 = u_CSAwallace_cla8_csa0_csa_component_fa7_xor1 ^ u_CSAwallace_cla8_csa0_csa_component_fa6_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa7_and0 = u_CSAwallace_cla8_csa0_csa_component_fa7_xor1 & u_CSAwallace_cla8_csa0_csa_component_fa6_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa7_xor1 = u_CSAwallace_cla8_csa2_csa_component_fa7_xor0 ^ u_CSAwallace_cla8_csa1_csa_component_fa7_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa7_and1 = u_CSAwallace_cla8_csa2_csa_component_fa7_xor0 & u_CSAwallace_cla8_csa1_csa_component_fa7_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa7_or0 = u_CSAwallace_cla8_csa2_csa_component_fa7_and0 | u_CSAwallace_cla8_csa2_csa_component_fa7_and1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa8_xor0 = u_CSAwallace_cla8_csa0_csa_component_fa8_xor1 ^ u_CSAwallace_cla8_csa0_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa8_and0 = u_CSAwallace_cla8_csa0_csa_component_fa8_xor1 & u_CSAwallace_cla8_csa0_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_csa2_csa_component_fa8_xor1 = u_CSAwallace_cla8_csa2_csa_component_fa8_xor0 ^ u_CSAwallace_cla8_csa1_csa_component_fa8_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa8_and1 = u_CSAwallace_cla8_csa2_csa_component_fa8_xor0 & u_CSAwallace_cla8_csa1_csa_component_fa8_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa8_or0 = u_CSAwallace_cla8_csa2_csa_component_fa8_and0 | u_CSAwallace_cla8_csa2_csa_component_fa8_and1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa9_xor0 = u_CSAwallace_cla8_and_7_2 ^ u_CSAwallace_cla8_csa0_csa_component_fa8_and1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa9_and0 = u_CSAwallace_cla8_and_7_2 & u_CSAwallace_cla8_csa0_csa_component_fa8_and1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa9_xor1 = u_CSAwallace_cla8_csa2_csa_component_fa9_xor0 ^ u_CSAwallace_cla8_csa1_csa_component_fa9_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa9_and1 = u_CSAwallace_cla8_csa2_csa_component_fa9_xor0 & u_CSAwallace_cla8_csa1_csa_component_fa9_xor1;
  assign u_CSAwallace_cla8_csa2_csa_component_fa9_or0 = u_CSAwallace_cla8_csa2_csa_component_fa9_and0 | u_CSAwallace_cla8_csa2_csa_component_fa9_and1;
  assign u_CSAwallace_cla8_csa3_csa_component_fa6_xor0 = u_CSAwallace_cla8_csa1_csa_component_fa5_or0 ^ u_CSAwallace_cla8_and_0_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa6_and0 = u_CSAwallace_cla8_csa1_csa_component_fa5_or0 & u_CSAwallace_cla8_and_0_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa7_xor0 = u_CSAwallace_cla8_csa1_csa_component_fa6_or0 ^ u_CSAwallace_cla8_and_1_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa7_and0 = u_CSAwallace_cla8_csa1_csa_component_fa6_or0 & u_CSAwallace_cla8_and_1_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa7_xor1 = u_CSAwallace_cla8_csa3_csa_component_fa7_xor0 ^ u_CSAwallace_cla8_and_0_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa7_and1 = u_CSAwallace_cla8_csa3_csa_component_fa7_xor0 & u_CSAwallace_cla8_and_0_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa7_or0 = u_CSAwallace_cla8_csa3_csa_component_fa7_and0 | u_CSAwallace_cla8_csa3_csa_component_fa7_and1;
  assign u_CSAwallace_cla8_csa3_csa_component_fa8_xor0 = u_CSAwallace_cla8_csa1_csa_component_fa7_or0 ^ u_CSAwallace_cla8_and_2_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa8_and0 = u_CSAwallace_cla8_csa1_csa_component_fa7_or0 & u_CSAwallace_cla8_and_2_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa8_xor1 = u_CSAwallace_cla8_csa3_csa_component_fa8_xor0 ^ u_CSAwallace_cla8_and_1_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa8_and1 = u_CSAwallace_cla8_csa3_csa_component_fa8_xor0 & u_CSAwallace_cla8_and_1_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa8_or0 = u_CSAwallace_cla8_csa3_csa_component_fa8_and0 | u_CSAwallace_cla8_csa3_csa_component_fa8_and1;
  assign u_CSAwallace_cla8_csa3_csa_component_fa9_xor0 = u_CSAwallace_cla8_csa1_csa_component_fa8_or0 ^ u_CSAwallace_cla8_and_3_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa9_and0 = u_CSAwallace_cla8_csa1_csa_component_fa8_or0 & u_CSAwallace_cla8_and_3_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa9_xor1 = u_CSAwallace_cla8_csa3_csa_component_fa9_xor0 ^ u_CSAwallace_cla8_and_2_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa9_and1 = u_CSAwallace_cla8_csa3_csa_component_fa9_xor0 & u_CSAwallace_cla8_and_2_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa9_or0 = u_CSAwallace_cla8_csa3_csa_component_fa9_and0 | u_CSAwallace_cla8_csa3_csa_component_fa9_and1;
  assign u_CSAwallace_cla8_csa3_csa_component_fa10_xor0 = u_CSAwallace_cla8_csa1_csa_component_fa9_or0 ^ u_CSAwallace_cla8_and_4_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa10_and0 = u_CSAwallace_cla8_csa1_csa_component_fa9_or0 & u_CSAwallace_cla8_and_4_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa10_xor1 = u_CSAwallace_cla8_csa3_csa_component_fa10_xor0 ^ u_CSAwallace_cla8_and_3_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa10_and1 = u_CSAwallace_cla8_csa3_csa_component_fa10_xor0 & u_CSAwallace_cla8_and_3_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa10_or0 = u_CSAwallace_cla8_csa3_csa_component_fa10_and0 | u_CSAwallace_cla8_csa3_csa_component_fa10_and1;
  assign u_CSAwallace_cla8_csa3_csa_component_fa11_xor0 = u_CSAwallace_cla8_csa1_csa_component_fa10_or0 ^ u_CSAwallace_cla8_and_5_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa11_and0 = u_CSAwallace_cla8_csa1_csa_component_fa10_or0 & u_CSAwallace_cla8_and_5_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa11_xor1 = u_CSAwallace_cla8_csa3_csa_component_fa11_xor0 ^ u_CSAwallace_cla8_and_4_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa11_and1 = u_CSAwallace_cla8_csa3_csa_component_fa11_xor0 & u_CSAwallace_cla8_and_4_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa11_or0 = u_CSAwallace_cla8_csa3_csa_component_fa11_and0 | u_CSAwallace_cla8_csa3_csa_component_fa11_and1;
  assign u_CSAwallace_cla8_csa3_csa_component_fa12_xor0 = u_CSAwallace_cla8_csa1_csa_component_fa11_and1 ^ u_CSAwallace_cla8_and_6_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa12_and0 = u_CSAwallace_cla8_csa1_csa_component_fa11_and1 & u_CSAwallace_cla8_and_6_6;
  assign u_CSAwallace_cla8_csa3_csa_component_fa12_xor1 = u_CSAwallace_cla8_csa3_csa_component_fa12_xor0 ^ u_CSAwallace_cla8_and_5_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa12_and1 = u_CSAwallace_cla8_csa3_csa_component_fa12_xor0 & u_CSAwallace_cla8_and_5_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa12_or0 = u_CSAwallace_cla8_csa3_csa_component_fa12_and0 | u_CSAwallace_cla8_csa3_csa_component_fa12_and1;
  assign u_CSAwallace_cla8_csa3_csa_component_fa13_xor1 = u_CSAwallace_cla8_and_7_6 ^ u_CSAwallace_cla8_and_6_7;
  assign u_CSAwallace_cla8_csa3_csa_component_fa13_and1 = u_CSAwallace_cla8_and_7_6 & u_CSAwallace_cla8_and_6_7;
  assign u_CSAwallace_cla8_csa4_csa_component_fa3_xor0 = u_CSAwallace_cla8_csa2_csa_component_fa3_xor1 ^ u_CSAwallace_cla8_csa2_csa_component_fa2_and0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa3_and0 = u_CSAwallace_cla8_csa2_csa_component_fa3_xor1 & u_CSAwallace_cla8_csa2_csa_component_fa2_and0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa4_xor0 = u_CSAwallace_cla8_csa2_csa_component_fa4_xor1 ^ u_CSAwallace_cla8_csa2_csa_component_fa3_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa4_and0 = u_CSAwallace_cla8_csa2_csa_component_fa4_xor1 & u_CSAwallace_cla8_csa2_csa_component_fa3_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa5_xor0 = u_CSAwallace_cla8_csa2_csa_component_fa5_xor1 ^ u_CSAwallace_cla8_csa2_csa_component_fa4_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa5_and0 = u_CSAwallace_cla8_csa2_csa_component_fa5_xor1 & u_CSAwallace_cla8_csa2_csa_component_fa4_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa5_xor1 = u_CSAwallace_cla8_csa4_csa_component_fa5_xor0 ^ u_CSAwallace_cla8_csa1_csa_component_fa4_and0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa5_and1 = u_CSAwallace_cla8_csa4_csa_component_fa5_xor0 & u_CSAwallace_cla8_csa1_csa_component_fa4_and0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa5_or0 = u_CSAwallace_cla8_csa4_csa_component_fa5_and0 | u_CSAwallace_cla8_csa4_csa_component_fa5_and1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa6_xor0 = u_CSAwallace_cla8_csa2_csa_component_fa6_xor1 ^ u_CSAwallace_cla8_csa2_csa_component_fa5_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa6_and0 = u_CSAwallace_cla8_csa2_csa_component_fa6_xor1 & u_CSAwallace_cla8_csa2_csa_component_fa5_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa6_xor1 = u_CSAwallace_cla8_csa4_csa_component_fa6_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa6_xor0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa6_and1 = u_CSAwallace_cla8_csa4_csa_component_fa6_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa6_xor0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa6_or0 = u_CSAwallace_cla8_csa4_csa_component_fa6_and0 | u_CSAwallace_cla8_csa4_csa_component_fa6_and1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa7_xor0 = u_CSAwallace_cla8_csa2_csa_component_fa7_xor1 ^ u_CSAwallace_cla8_csa2_csa_component_fa6_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa7_and0 = u_CSAwallace_cla8_csa2_csa_component_fa7_xor1 & u_CSAwallace_cla8_csa2_csa_component_fa6_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa7_xor1 = u_CSAwallace_cla8_csa4_csa_component_fa7_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa7_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa7_and1 = u_CSAwallace_cla8_csa4_csa_component_fa7_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa7_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa7_or0 = u_CSAwallace_cla8_csa4_csa_component_fa7_and0 | u_CSAwallace_cla8_csa4_csa_component_fa7_and1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa8_xor0 = u_CSAwallace_cla8_csa2_csa_component_fa8_xor1 ^ u_CSAwallace_cla8_csa2_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa8_and0 = u_CSAwallace_cla8_csa2_csa_component_fa8_xor1 & u_CSAwallace_cla8_csa2_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa8_xor1 = u_CSAwallace_cla8_csa4_csa_component_fa8_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa8_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa8_and1 = u_CSAwallace_cla8_csa4_csa_component_fa8_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa8_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa8_or0 = u_CSAwallace_cla8_csa4_csa_component_fa8_and0 | u_CSAwallace_cla8_csa4_csa_component_fa8_and1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa9_xor0 = u_CSAwallace_cla8_csa2_csa_component_fa9_xor1 ^ u_CSAwallace_cla8_csa2_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa9_and0 = u_CSAwallace_cla8_csa2_csa_component_fa9_xor1 & u_CSAwallace_cla8_csa2_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa9_xor1 = u_CSAwallace_cla8_csa4_csa_component_fa9_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa9_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa9_and1 = u_CSAwallace_cla8_csa4_csa_component_fa9_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa9_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa9_or0 = u_CSAwallace_cla8_csa4_csa_component_fa9_and0 | u_CSAwallace_cla8_csa4_csa_component_fa9_and1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa10_xor0 = u_CSAwallace_cla8_csa1_csa_component_fa10_xor1 ^ u_CSAwallace_cla8_csa2_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa10_and0 = u_CSAwallace_cla8_csa1_csa_component_fa10_xor1 & u_CSAwallace_cla8_csa2_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_csa4_csa_component_fa10_xor1 = u_CSAwallace_cla8_csa4_csa_component_fa10_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa10_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa10_and1 = u_CSAwallace_cla8_csa4_csa_component_fa10_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa10_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa10_or0 = u_CSAwallace_cla8_csa4_csa_component_fa10_and0 | u_CSAwallace_cla8_csa4_csa_component_fa10_and1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa11_xor1 = u_CSAwallace_cla8_csa1_csa_component_fa11_xor1 ^ u_CSAwallace_cla8_csa3_csa_component_fa11_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa11_and1 = u_CSAwallace_cla8_csa1_csa_component_fa11_xor1 & u_CSAwallace_cla8_csa3_csa_component_fa11_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa12_xor1 = u_CSAwallace_cla8_and_7_5 ^ u_CSAwallace_cla8_csa3_csa_component_fa12_xor1;
  assign u_CSAwallace_cla8_csa4_csa_component_fa12_and1 = u_CSAwallace_cla8_and_7_5 & u_CSAwallace_cla8_csa3_csa_component_fa12_xor1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa4_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa4_xor0 ^ u_CSAwallace_cla8_csa4_csa_component_fa3_and0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa4_and0 = u_CSAwallace_cla8_csa4_csa_component_fa4_xor0 & u_CSAwallace_cla8_csa4_csa_component_fa3_and0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa5_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa5_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa4_and0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa5_and0 = u_CSAwallace_cla8_csa4_csa_component_fa5_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa4_and0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa6_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa6_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa5_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa6_and0 = u_CSAwallace_cla8_csa4_csa_component_fa6_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa5_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa7_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa7_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa6_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa7_and0 = u_CSAwallace_cla8_csa4_csa_component_fa7_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa6_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa7_xor1 = u_CSAwallace_cla8_csa5_csa_component_fa7_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa6_and0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa7_and1 = u_CSAwallace_cla8_csa5_csa_component_fa7_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa6_and0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa7_or0 = u_CSAwallace_cla8_csa5_csa_component_fa7_and0 | u_CSAwallace_cla8_csa5_csa_component_fa7_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa8_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa8_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa8_and0 = u_CSAwallace_cla8_csa4_csa_component_fa8_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa8_xor1 = u_CSAwallace_cla8_csa5_csa_component_fa8_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa8_and1 = u_CSAwallace_cla8_csa5_csa_component_fa8_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa8_or0 = u_CSAwallace_cla8_csa5_csa_component_fa8_and0 | u_CSAwallace_cla8_csa5_csa_component_fa8_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa9_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa9_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa9_and0 = u_CSAwallace_cla8_csa4_csa_component_fa9_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa9_xor1 = u_CSAwallace_cla8_csa5_csa_component_fa9_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa9_and1 = u_CSAwallace_cla8_csa5_csa_component_fa9_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa9_or0 = u_CSAwallace_cla8_csa5_csa_component_fa9_and0 | u_CSAwallace_cla8_csa5_csa_component_fa9_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa10_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa10_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa10_and0 = u_CSAwallace_cla8_csa4_csa_component_fa10_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa10_xor1 = u_CSAwallace_cla8_csa5_csa_component_fa10_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa10_and1 = u_CSAwallace_cla8_csa5_csa_component_fa10_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa10_or0 = u_CSAwallace_cla8_csa5_csa_component_fa10_and0 | u_CSAwallace_cla8_csa5_csa_component_fa10_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa11_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa11_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa10_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa11_and0 = u_CSAwallace_cla8_csa4_csa_component_fa11_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa10_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa11_xor1 = u_CSAwallace_cla8_csa5_csa_component_fa11_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa10_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa11_and1 = u_CSAwallace_cla8_csa5_csa_component_fa11_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa10_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa11_or0 = u_CSAwallace_cla8_csa5_csa_component_fa11_and0 | u_CSAwallace_cla8_csa5_csa_component_fa11_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa12_xor0 = u_CSAwallace_cla8_csa4_csa_component_fa12_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa11_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa12_and0 = u_CSAwallace_cla8_csa4_csa_component_fa12_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa11_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa12_xor1 = u_CSAwallace_cla8_csa5_csa_component_fa12_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa11_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa12_and1 = u_CSAwallace_cla8_csa5_csa_component_fa12_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa11_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa12_or0 = u_CSAwallace_cla8_csa5_csa_component_fa12_and0 | u_CSAwallace_cla8_csa5_csa_component_fa12_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa13_xor0 = u_CSAwallace_cla8_csa3_csa_component_fa13_xor1 ^ u_CSAwallace_cla8_csa4_csa_component_fa12_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa13_and0 = u_CSAwallace_cla8_csa3_csa_component_fa13_xor1 & u_CSAwallace_cla8_csa4_csa_component_fa12_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa13_xor1 = u_CSAwallace_cla8_csa5_csa_component_fa13_xor0 ^ u_CSAwallace_cla8_csa3_csa_component_fa12_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa13_and1 = u_CSAwallace_cla8_csa5_csa_component_fa13_xor0 & u_CSAwallace_cla8_csa3_csa_component_fa12_or0;
  assign u_CSAwallace_cla8_csa5_csa_component_fa13_or0 = u_CSAwallace_cla8_csa5_csa_component_fa13_and0 | u_CSAwallace_cla8_csa5_csa_component_fa13_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa14_xor1 = u_CSAwallace_cla8_and_7_7 ^ u_CSAwallace_cla8_csa3_csa_component_fa13_and1;
  assign u_CSAwallace_cla8_csa5_csa_component_fa14_and1 = u_CSAwallace_cla8_and_7_7 & u_CSAwallace_cla8_csa3_csa_component_fa13_and1;
  assign u_CSAwallace_cla8_u_cla16_and0 = u_CSAwallace_cla8_csa2_csa_component_fa2_xor0 & u_CSAwallace_cla8_and_0_0;
  assign u_CSAwallace_cla8_u_cla16_and1 = u_CSAwallace_cla8_csa4_csa_component_fa3_xor0 & u_CSAwallace_cla8_csa0_csa_component_fa1_xor0;
  assign u_CSAwallace_cla8_u_cla16_and2 = u_CSAwallace_cla8_csa4_csa_component_fa3_xor0 & u_CSAwallace_cla8_csa0_csa_component_fa1_xor0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic5_or0 = u_CSAwallace_cla8_csa5_csa_component_fa5_xor0 | u_CSAwallace_cla8_csa5_csa_component_fa4_and0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic5_and0 = u_CSAwallace_cla8_csa5_csa_component_fa5_xor0 & u_CSAwallace_cla8_csa5_csa_component_fa4_and0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic5_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa5_xor0 ^ u_CSAwallace_cla8_csa5_csa_component_fa4_and0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic6_or0 = u_CSAwallace_cla8_csa5_csa_component_fa6_xor0 | u_CSAwallace_cla8_csa5_csa_component_fa5_and0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic6_and0 = u_CSAwallace_cla8_csa5_csa_component_fa6_xor0 & u_CSAwallace_cla8_csa5_csa_component_fa5_and0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic6_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa6_xor0 ^ u_CSAwallace_cla8_csa5_csa_component_fa5_and0;
  assign u_CSAwallace_cla8_u_cla16_xor6 = u_CSAwallace_cla8_u_cla16_pg_logic6_xor0 ^ u_CSAwallace_cla8_u_cla16_pg_logic5_and0;
  assign u_CSAwallace_cla8_u_cla16_and3 = u_CSAwallace_cla8_u_cla16_pg_logic6_or0 & u_CSAwallace_cla8_csa5_csa_component_fa4_xor0;
  assign u_CSAwallace_cla8_u_cla16_and4 = u_CSAwallace_cla8_u_cla16_pg_logic5_and0 & u_CSAwallace_cla8_u_cla16_pg_logic6_or0;
  assign u_CSAwallace_cla8_u_cla16_or0 = u_CSAwallace_cla8_u_cla16_pg_logic6_and0 | u_CSAwallace_cla8_u_cla16_and4;
  assign u_CSAwallace_cla8_u_cla16_pg_logic7_or0 = u_CSAwallace_cla8_csa5_csa_component_fa7_xor1 | u_CSAwallace_cla8_csa5_csa_component_fa6_and0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic7_and0 = u_CSAwallace_cla8_csa5_csa_component_fa7_xor1 & u_CSAwallace_cla8_csa5_csa_component_fa6_and0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic7_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa7_xor1 ^ u_CSAwallace_cla8_csa5_csa_component_fa6_and0;
  assign u_CSAwallace_cla8_u_cla16_xor7 = u_CSAwallace_cla8_u_cla16_pg_logic7_xor0 ^ u_CSAwallace_cla8_u_cla16_or0;
  assign u_CSAwallace_cla8_u_cla16_and5 = u_CSAwallace_cla8_u_cla16_pg_logic7_or0 & u_CSAwallace_cla8_u_cla16_pg_logic5_or0;
  assign u_CSAwallace_cla8_u_cla16_and6 = u_CSAwallace_cla8_u_cla16_pg_logic7_or0 & u_CSAwallace_cla8_u_cla16_pg_logic5_or0;
  assign u_CSAwallace_cla8_u_cla16_and7 = u_CSAwallace_cla8_u_cla16_pg_logic5_and0 & u_CSAwallace_cla8_u_cla16_pg_logic7_or0;
  assign u_CSAwallace_cla8_u_cla16_and8 = u_CSAwallace_cla8_u_cla16_and7 & u_CSAwallace_cla8_u_cla16_pg_logic6_or0;
  assign u_CSAwallace_cla8_u_cla16_and9 = u_CSAwallace_cla8_u_cla16_pg_logic6_and0 & u_CSAwallace_cla8_u_cla16_pg_logic7_or0;
  assign u_CSAwallace_cla8_u_cla16_or1 = u_CSAwallace_cla8_u_cla16_and8 | u_CSAwallace_cla8_u_cla16_and9;
  assign u_CSAwallace_cla8_u_cla16_or2 = u_CSAwallace_cla8_u_cla16_pg_logic7_and0 | u_CSAwallace_cla8_u_cla16_or1;
  assign u_CSAwallace_cla8_u_cla16_pg_logic8_or0 = u_CSAwallace_cla8_csa5_csa_component_fa8_xor1 | u_CSAwallace_cla8_csa5_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic8_and0 = u_CSAwallace_cla8_csa5_csa_component_fa8_xor1 & u_CSAwallace_cla8_csa5_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic8_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa8_xor1 ^ u_CSAwallace_cla8_csa5_csa_component_fa7_or0;
  assign u_CSAwallace_cla8_u_cla16_xor8 = u_CSAwallace_cla8_u_cla16_pg_logic8_xor0 ^ u_CSAwallace_cla8_u_cla16_or2;
  assign u_CSAwallace_cla8_u_cla16_and10 = u_CSAwallace_cla8_u_cla16_or2 & u_CSAwallace_cla8_u_cla16_pg_logic8_or0;
  assign u_CSAwallace_cla8_u_cla16_or3 = u_CSAwallace_cla8_u_cla16_pg_logic8_and0 | u_CSAwallace_cla8_u_cla16_and10;
  assign u_CSAwallace_cla8_u_cla16_pg_logic9_or0 = u_CSAwallace_cla8_csa5_csa_component_fa9_xor1 | u_CSAwallace_cla8_csa5_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic9_and0 = u_CSAwallace_cla8_csa5_csa_component_fa9_xor1 & u_CSAwallace_cla8_csa5_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic9_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa9_xor1 ^ u_CSAwallace_cla8_csa5_csa_component_fa8_or0;
  assign u_CSAwallace_cla8_u_cla16_xor9 = u_CSAwallace_cla8_u_cla16_pg_logic9_xor0 ^ u_CSAwallace_cla8_u_cla16_or3;
  assign u_CSAwallace_cla8_u_cla16_and11 = u_CSAwallace_cla8_u_cla16_or2 & u_CSAwallace_cla8_u_cla16_pg_logic9_or0;
  assign u_CSAwallace_cla8_u_cla16_and12 = u_CSAwallace_cla8_u_cla16_and11 & u_CSAwallace_cla8_u_cla16_pg_logic8_or0;
  assign u_CSAwallace_cla8_u_cla16_and13 = u_CSAwallace_cla8_u_cla16_pg_logic8_and0 & u_CSAwallace_cla8_u_cla16_pg_logic9_or0;
  assign u_CSAwallace_cla8_u_cla16_or4 = u_CSAwallace_cla8_u_cla16_and12 | u_CSAwallace_cla8_u_cla16_and13;
  assign u_CSAwallace_cla8_u_cla16_or5 = u_CSAwallace_cla8_u_cla16_pg_logic9_and0 | u_CSAwallace_cla8_u_cla16_or4;
  assign u_CSAwallace_cla8_u_cla16_pg_logic10_or0 = u_CSAwallace_cla8_csa5_csa_component_fa10_xor1 | u_CSAwallace_cla8_csa5_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic10_and0 = u_CSAwallace_cla8_csa5_csa_component_fa10_xor1 & u_CSAwallace_cla8_csa5_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic10_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa10_xor1 ^ u_CSAwallace_cla8_csa5_csa_component_fa9_or0;
  assign u_CSAwallace_cla8_u_cla16_xor10 = u_CSAwallace_cla8_u_cla16_pg_logic10_xor0 ^ u_CSAwallace_cla8_u_cla16_or5;
  assign u_CSAwallace_cla8_u_cla16_and14 = u_CSAwallace_cla8_u_cla16_or2 & u_CSAwallace_cla8_u_cla16_pg_logic9_or0;
  assign u_CSAwallace_cla8_u_cla16_and15 = u_CSAwallace_cla8_u_cla16_pg_logic10_or0 & u_CSAwallace_cla8_u_cla16_pg_logic8_or0;
  assign u_CSAwallace_cla8_u_cla16_and16 = u_CSAwallace_cla8_u_cla16_and14 & u_CSAwallace_cla8_u_cla16_and15;
  assign u_CSAwallace_cla8_u_cla16_and17 = u_CSAwallace_cla8_u_cla16_pg_logic8_and0 & u_CSAwallace_cla8_u_cla16_pg_logic10_or0;
  assign u_CSAwallace_cla8_u_cla16_and18 = u_CSAwallace_cla8_u_cla16_and17 & u_CSAwallace_cla8_u_cla16_pg_logic9_or0;
  assign u_CSAwallace_cla8_u_cla16_and19 = u_CSAwallace_cla8_u_cla16_pg_logic9_and0 & u_CSAwallace_cla8_u_cla16_pg_logic10_or0;
  assign u_CSAwallace_cla8_u_cla16_or6 = u_CSAwallace_cla8_u_cla16_and16 | u_CSAwallace_cla8_u_cla16_and18;
  assign u_CSAwallace_cla8_u_cla16_or7 = u_CSAwallace_cla8_u_cla16_or6 | u_CSAwallace_cla8_u_cla16_and19;
  assign u_CSAwallace_cla8_u_cla16_or8 = u_CSAwallace_cla8_u_cla16_pg_logic10_and0 | u_CSAwallace_cla8_u_cla16_or7;
  assign u_CSAwallace_cla8_u_cla16_pg_logic11_or0 = u_CSAwallace_cla8_csa5_csa_component_fa11_xor1 | u_CSAwallace_cla8_csa5_csa_component_fa10_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic11_and0 = u_CSAwallace_cla8_csa5_csa_component_fa11_xor1 & u_CSAwallace_cla8_csa5_csa_component_fa10_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic11_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa11_xor1 ^ u_CSAwallace_cla8_csa5_csa_component_fa10_or0;
  assign u_CSAwallace_cla8_u_cla16_xor11 = u_CSAwallace_cla8_u_cla16_pg_logic11_xor0 ^ u_CSAwallace_cla8_u_cla16_or8;
  assign u_CSAwallace_cla8_u_cla16_and20 = u_CSAwallace_cla8_u_cla16_or2 & u_CSAwallace_cla8_u_cla16_pg_logic10_or0;
  assign u_CSAwallace_cla8_u_cla16_and21 = u_CSAwallace_cla8_u_cla16_pg_logic11_or0 & u_CSAwallace_cla8_u_cla16_pg_logic9_or0;
  assign u_CSAwallace_cla8_u_cla16_and22 = u_CSAwallace_cla8_u_cla16_and20 & u_CSAwallace_cla8_u_cla16_and21;
  assign u_CSAwallace_cla8_u_cla16_and23 = u_CSAwallace_cla8_u_cla16_and22 & u_CSAwallace_cla8_u_cla16_pg_logic8_or0;
  assign u_CSAwallace_cla8_u_cla16_and24 = u_CSAwallace_cla8_u_cla16_pg_logic8_and0 & u_CSAwallace_cla8_u_cla16_pg_logic10_or0;
  assign u_CSAwallace_cla8_u_cla16_and25 = u_CSAwallace_cla8_u_cla16_pg_logic11_or0 & u_CSAwallace_cla8_u_cla16_pg_logic9_or0;
  assign u_CSAwallace_cla8_u_cla16_and26 = u_CSAwallace_cla8_u_cla16_and24 & u_CSAwallace_cla8_u_cla16_and25;
  assign u_CSAwallace_cla8_u_cla16_and27 = u_CSAwallace_cla8_u_cla16_pg_logic9_and0 & u_CSAwallace_cla8_u_cla16_pg_logic11_or0;
  assign u_CSAwallace_cla8_u_cla16_and28 = u_CSAwallace_cla8_u_cla16_and27 & u_CSAwallace_cla8_u_cla16_pg_logic10_or0;
  assign u_CSAwallace_cla8_u_cla16_and29 = u_CSAwallace_cla8_u_cla16_pg_logic10_and0 & u_CSAwallace_cla8_u_cla16_pg_logic11_or0;
  assign u_CSAwallace_cla8_u_cla16_or9 = u_CSAwallace_cla8_u_cla16_and23 | u_CSAwallace_cla8_u_cla16_and28;
  assign u_CSAwallace_cla8_u_cla16_or10 = u_CSAwallace_cla8_u_cla16_and26 | u_CSAwallace_cla8_u_cla16_and29;
  assign u_CSAwallace_cla8_u_cla16_or11 = u_CSAwallace_cla8_u_cla16_or9 | u_CSAwallace_cla8_u_cla16_or10;
  assign u_CSAwallace_cla8_u_cla16_or12 = u_CSAwallace_cla8_u_cla16_pg_logic11_and0 | u_CSAwallace_cla8_u_cla16_or11;
  assign u_CSAwallace_cla8_u_cla16_pg_logic12_or0 = u_CSAwallace_cla8_csa5_csa_component_fa12_xor1 | u_CSAwallace_cla8_csa5_csa_component_fa11_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic12_and0 = u_CSAwallace_cla8_csa5_csa_component_fa12_xor1 & u_CSAwallace_cla8_csa5_csa_component_fa11_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic12_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa12_xor1 ^ u_CSAwallace_cla8_csa5_csa_component_fa11_or0;
  assign u_CSAwallace_cla8_u_cla16_xor12 = u_CSAwallace_cla8_u_cla16_pg_logic12_xor0 ^ u_CSAwallace_cla8_u_cla16_or12;
  assign u_CSAwallace_cla8_u_cla16_and30 = u_CSAwallace_cla8_u_cla16_or12 & u_CSAwallace_cla8_u_cla16_pg_logic12_or0;
  assign u_CSAwallace_cla8_u_cla16_or13 = u_CSAwallace_cla8_u_cla16_pg_logic12_and0 | u_CSAwallace_cla8_u_cla16_and30;
  assign u_CSAwallace_cla8_u_cla16_pg_logic13_or0 = u_CSAwallace_cla8_csa5_csa_component_fa13_xor1 | u_CSAwallace_cla8_csa5_csa_component_fa12_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic13_and0 = u_CSAwallace_cla8_csa5_csa_component_fa13_xor1 & u_CSAwallace_cla8_csa5_csa_component_fa12_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic13_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa13_xor1 ^ u_CSAwallace_cla8_csa5_csa_component_fa12_or0;
  assign u_CSAwallace_cla8_u_cla16_xor13 = u_CSAwallace_cla8_u_cla16_pg_logic13_xor0 ^ u_CSAwallace_cla8_u_cla16_or13;
  assign u_CSAwallace_cla8_u_cla16_and31 = u_CSAwallace_cla8_u_cla16_or12 & u_CSAwallace_cla8_u_cla16_pg_logic13_or0;
  assign u_CSAwallace_cla8_u_cla16_and32 = u_CSAwallace_cla8_u_cla16_and31 & u_CSAwallace_cla8_u_cla16_pg_logic12_or0;
  assign u_CSAwallace_cla8_u_cla16_and33 = u_CSAwallace_cla8_u_cla16_pg_logic12_and0 & u_CSAwallace_cla8_u_cla16_pg_logic13_or0;
  assign u_CSAwallace_cla8_u_cla16_or14 = u_CSAwallace_cla8_u_cla16_and32 | u_CSAwallace_cla8_u_cla16_and33;
  assign u_CSAwallace_cla8_u_cla16_or15 = u_CSAwallace_cla8_u_cla16_pg_logic13_and0 | u_CSAwallace_cla8_u_cla16_or14;
  assign u_CSAwallace_cla8_u_cla16_pg_logic14_or0 = u_CSAwallace_cla8_csa5_csa_component_fa14_xor1 | u_CSAwallace_cla8_csa5_csa_component_fa13_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic14_and0 = u_CSAwallace_cla8_csa5_csa_component_fa14_xor1 & u_CSAwallace_cla8_csa5_csa_component_fa13_or0;
  assign u_CSAwallace_cla8_u_cla16_pg_logic14_xor0 = u_CSAwallace_cla8_csa5_csa_component_fa14_xor1 ^ u_CSAwallace_cla8_csa5_csa_component_fa13_or0;
  assign u_CSAwallace_cla8_u_cla16_xor14 = u_CSAwallace_cla8_u_cla16_pg_logic14_xor0 ^ u_CSAwallace_cla8_u_cla16_or15;
  assign u_CSAwallace_cla8_u_cla16_and34 = u_CSAwallace_cla8_u_cla16_or12 & u_CSAwallace_cla8_u_cla16_pg_logic13_or0;
  assign u_CSAwallace_cla8_u_cla16_and35 = u_CSAwallace_cla8_u_cla16_pg_logic14_or0 & u_CSAwallace_cla8_u_cla16_pg_logic12_or0;
  assign u_CSAwallace_cla8_u_cla16_and36 = u_CSAwallace_cla8_u_cla16_and34 & u_CSAwallace_cla8_u_cla16_and35;
  assign u_CSAwallace_cla8_u_cla16_and37 = u_CSAwallace_cla8_u_cla16_pg_logic12_and0 & u_CSAwallace_cla8_u_cla16_pg_logic14_or0;
  assign u_CSAwallace_cla8_u_cla16_and38 = u_CSAwallace_cla8_u_cla16_and37 & u_CSAwallace_cla8_u_cla16_pg_logic13_or0;
  assign u_CSAwallace_cla8_u_cla16_and39 = u_CSAwallace_cla8_u_cla16_pg_logic13_and0 & u_CSAwallace_cla8_u_cla16_pg_logic14_or0;
  assign u_CSAwallace_cla8_u_cla16_or16 = u_CSAwallace_cla8_u_cla16_and36 | u_CSAwallace_cla8_u_cla16_and38;
  assign u_CSAwallace_cla8_u_cla16_or17 = u_CSAwallace_cla8_u_cla16_or16 | u_CSAwallace_cla8_u_cla16_and39;
  assign u_CSAwallace_cla8_u_cla16_or18 = u_CSAwallace_cla8_u_cla16_pg_logic14_and0 | u_CSAwallace_cla8_u_cla16_or17;
  assign u_CSAwallace_cla8_u_cla16_xor15 = u_CSAwallace_cla8_csa5_csa_component_fa14_and1 ^ u_CSAwallace_cla8_u_cla16_or18;
  assign u_CSAwallace_cla8_u_cla16_and40 = u_CSAwallace_cla8_u_cla16_or12 & u_CSAwallace_cla8_u_cla16_pg_logic14_or0;
  assign u_CSAwallace_cla8_u_cla16_and41 = u_CSAwallace_cla8_csa5_csa_component_fa14_and1 & u_CSAwallace_cla8_u_cla16_pg_logic13_or0;
  assign u_CSAwallace_cla8_u_cla16_and42 = u_CSAwallace_cla8_u_cla16_and40 & u_CSAwallace_cla8_u_cla16_and41;
  assign u_CSAwallace_cla8_u_cla16_and43 = u_CSAwallace_cla8_u_cla16_and42 & u_CSAwallace_cla8_u_cla16_pg_logic12_or0;
  assign u_CSAwallace_cla8_u_cla16_and44 = u_CSAwallace_cla8_u_cla16_pg_logic12_and0 & u_CSAwallace_cla8_u_cla16_pg_logic14_or0;
  assign u_CSAwallace_cla8_u_cla16_and45 = u_CSAwallace_cla8_csa5_csa_component_fa14_and1 & u_CSAwallace_cla8_u_cla16_pg_logic13_or0;
  assign u_CSAwallace_cla8_u_cla16_and46 = u_CSAwallace_cla8_u_cla16_and44 & u_CSAwallace_cla8_u_cla16_and45;
  assign u_CSAwallace_cla8_u_cla16_and47 = u_CSAwallace_cla8_u_cla16_pg_logic13_and0 & u_CSAwallace_cla8_csa5_csa_component_fa14_and1;
  assign u_CSAwallace_cla8_u_cla16_and48 = u_CSAwallace_cla8_u_cla16_and47 & u_CSAwallace_cla8_u_cla16_pg_logic14_or0;
  assign u_CSAwallace_cla8_u_cla16_and49 = u_CSAwallace_cla8_u_cla16_pg_logic14_and0 & u_CSAwallace_cla8_csa5_csa_component_fa14_and1;
  assign u_CSAwallace_cla8_u_cla16_or19 = u_CSAwallace_cla8_u_cla16_and43 | u_CSAwallace_cla8_u_cla16_and48;
  assign u_CSAwallace_cla8_u_cla16_or20 = u_CSAwallace_cla8_u_cla16_and46 | u_CSAwallace_cla8_u_cla16_and49;
  assign u_CSAwallace_cla8_u_cla16_or21 = u_CSAwallace_cla8_u_cla16_or19 | u_CSAwallace_cla8_u_cla16_or20;

  assign u_CSAwallace_cla8_out[0] = u_CSAwallace_cla8_and_0_0;
  assign u_CSAwallace_cla8_out[1] = u_CSAwallace_cla8_csa0_csa_component_fa1_xor0;
  assign u_CSAwallace_cla8_out[2] = u_CSAwallace_cla8_csa2_csa_component_fa2_xor0;
  assign u_CSAwallace_cla8_out[3] = u_CSAwallace_cla8_csa4_csa_component_fa3_xor0;
  assign u_CSAwallace_cla8_out[4] = u_CSAwallace_cla8_csa5_csa_component_fa4_xor0;
  assign u_CSAwallace_cla8_out[5] = u_CSAwallace_cla8_u_cla16_pg_logic5_xor0;
  assign u_CSAwallace_cla8_out[6] = u_CSAwallace_cla8_u_cla16_xor6;
  assign u_CSAwallace_cla8_out[7] = u_CSAwallace_cla8_u_cla16_xor7;
  assign u_CSAwallace_cla8_out[8] = u_CSAwallace_cla8_u_cla16_xor8;
  assign u_CSAwallace_cla8_out[9] = u_CSAwallace_cla8_u_cla16_xor9;
  assign u_CSAwallace_cla8_out[10] = u_CSAwallace_cla8_u_cla16_xor10;
  assign u_CSAwallace_cla8_out[11] = u_CSAwallace_cla8_u_cla16_xor11;
  assign u_CSAwallace_cla8_out[12] = u_CSAwallace_cla8_u_cla16_xor12;
  assign u_CSAwallace_cla8_out[13] = u_CSAwallace_cla8_u_cla16_xor13;
  assign u_CSAwallace_cla8_out[14] = u_CSAwallace_cla8_u_cla16_xor14;
  assign u_CSAwallace_cla8_out[15] = u_CSAwallace_cla8_u_cla16_xor15;
endmodule