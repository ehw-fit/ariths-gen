module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module nand_gate(input a, input b, output out);
  assign out = ~(a & b);
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module not_gate(input a, output out);
  assign out = ~a;
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module ha(input [0:0] a, input [0:0] b, output [0:0] ha_xor0, output [0:0] ha_and0);
  xor_gate xor_gate_ha_xor0(.a(a[0]), .b(b[0]), .out(ha_xor0));
  and_gate and_gate_ha_and0(.a(a[0]), .b(b[0]), .out(ha_and0));
endmodule

module csa_component14(input [13:0] a, input [13:0] b, input [13:0] c, output [29:0] csa_component14_out);
  wire [0:0] csa_component14_fa0_xor1;
  wire [0:0] csa_component14_fa0_or0;
  wire [0:0] csa_component14_fa1_xor1;
  wire [0:0] csa_component14_fa1_or0;
  wire [0:0] csa_component14_fa2_xor1;
  wire [0:0] csa_component14_fa2_or0;
  wire [0:0] csa_component14_fa3_xor1;
  wire [0:0] csa_component14_fa3_or0;
  wire [0:0] csa_component14_fa4_xor1;
  wire [0:0] csa_component14_fa4_or0;
  wire [0:0] csa_component14_fa5_xor1;
  wire [0:0] csa_component14_fa5_or0;
  wire [0:0] csa_component14_fa6_xor1;
  wire [0:0] csa_component14_fa6_or0;
  wire [0:0] csa_component14_fa7_xor1;
  wire [0:0] csa_component14_fa7_or0;
  wire [0:0] csa_component14_fa8_xor1;
  wire [0:0] csa_component14_fa8_or0;
  wire [0:0] csa_component14_fa9_xor1;
  wire [0:0] csa_component14_fa9_or0;
  wire [0:0] csa_component14_fa10_xor1;
  wire [0:0] csa_component14_fa10_or0;
  wire [0:0] csa_component14_fa11_xor1;
  wire [0:0] csa_component14_fa11_or0;
  wire [0:0] csa_component14_fa12_xor1;
  wire [0:0] csa_component14_fa12_or0;
  wire [0:0] csa_component14_fa13_xor1;
  wire [0:0] csa_component14_fa13_or0;

  fa fa_csa_component14_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component14_fa0_xor1), .fa_or0(csa_component14_fa0_or0));
  fa fa_csa_component14_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component14_fa1_xor1), .fa_or0(csa_component14_fa1_or0));
  fa fa_csa_component14_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component14_fa2_xor1), .fa_or0(csa_component14_fa2_or0));
  fa fa_csa_component14_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component14_fa3_xor1), .fa_or0(csa_component14_fa3_or0));
  fa fa_csa_component14_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component14_fa4_xor1), .fa_or0(csa_component14_fa4_or0));
  fa fa_csa_component14_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component14_fa5_xor1), .fa_or0(csa_component14_fa5_or0));
  fa fa_csa_component14_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component14_fa6_xor1), .fa_or0(csa_component14_fa6_or0));
  fa fa_csa_component14_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component14_fa7_xor1), .fa_or0(csa_component14_fa7_or0));
  fa fa_csa_component14_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component14_fa8_xor1), .fa_or0(csa_component14_fa8_or0));
  fa fa_csa_component14_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component14_fa9_xor1), .fa_or0(csa_component14_fa9_or0));
  fa fa_csa_component14_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component14_fa10_xor1), .fa_or0(csa_component14_fa10_or0));
  fa fa_csa_component14_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component14_fa11_xor1), .fa_or0(csa_component14_fa11_or0));
  fa fa_csa_component14_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component14_fa12_xor1), .fa_or0(csa_component14_fa12_or0));
  fa fa_csa_component14_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component14_fa13_xor1), .fa_or0(csa_component14_fa13_or0));

  assign csa_component14_out[0] = csa_component14_fa0_xor1[0];
  assign csa_component14_out[1] = csa_component14_fa1_xor1[0];
  assign csa_component14_out[2] = csa_component14_fa2_xor1[0];
  assign csa_component14_out[3] = csa_component14_fa3_xor1[0];
  assign csa_component14_out[4] = csa_component14_fa4_xor1[0];
  assign csa_component14_out[5] = csa_component14_fa5_xor1[0];
  assign csa_component14_out[6] = csa_component14_fa6_xor1[0];
  assign csa_component14_out[7] = csa_component14_fa7_xor1[0];
  assign csa_component14_out[8] = csa_component14_fa8_xor1[0];
  assign csa_component14_out[9] = csa_component14_fa9_xor1[0];
  assign csa_component14_out[10] = csa_component14_fa10_xor1[0];
  assign csa_component14_out[11] = csa_component14_fa11_xor1[0];
  assign csa_component14_out[12] = csa_component14_fa12_xor1[0];
  assign csa_component14_out[13] = csa_component14_fa13_xor1[0];
  assign csa_component14_out[14] = 1'b0;
  assign csa_component14_out[15] = 1'b0;
  assign csa_component14_out[16] = csa_component14_fa0_or0[0];
  assign csa_component14_out[17] = csa_component14_fa1_or0[0];
  assign csa_component14_out[18] = csa_component14_fa2_or0[0];
  assign csa_component14_out[19] = csa_component14_fa3_or0[0];
  assign csa_component14_out[20] = csa_component14_fa4_or0[0];
  assign csa_component14_out[21] = csa_component14_fa5_or0[0];
  assign csa_component14_out[22] = csa_component14_fa6_or0[0];
  assign csa_component14_out[23] = csa_component14_fa7_or0[0];
  assign csa_component14_out[24] = csa_component14_fa8_or0[0];
  assign csa_component14_out[25] = csa_component14_fa9_or0[0];
  assign csa_component14_out[26] = csa_component14_fa10_or0[0];
  assign csa_component14_out[27] = csa_component14_fa11_or0[0];
  assign csa_component14_out[28] = csa_component14_fa12_or0[0];
  assign csa_component14_out[29] = csa_component14_fa13_or0[0];
endmodule

module csa_component17(input [16:0] a, input [16:0] b, input [16:0] c, output [35:0] csa_component17_out);
  wire [0:0] csa_component17_fa0_xor1;
  wire [0:0] csa_component17_fa0_or0;
  wire [0:0] csa_component17_fa1_xor1;
  wire [0:0] csa_component17_fa1_or0;
  wire [0:0] csa_component17_fa2_xor1;
  wire [0:0] csa_component17_fa2_or0;
  wire [0:0] csa_component17_fa3_xor1;
  wire [0:0] csa_component17_fa3_or0;
  wire [0:0] csa_component17_fa4_xor1;
  wire [0:0] csa_component17_fa4_or0;
  wire [0:0] csa_component17_fa5_xor1;
  wire [0:0] csa_component17_fa5_or0;
  wire [0:0] csa_component17_fa6_xor1;
  wire [0:0] csa_component17_fa6_or0;
  wire [0:0] csa_component17_fa7_xor1;
  wire [0:0] csa_component17_fa7_or0;
  wire [0:0] csa_component17_fa8_xor1;
  wire [0:0] csa_component17_fa8_or0;
  wire [0:0] csa_component17_fa9_xor1;
  wire [0:0] csa_component17_fa9_or0;
  wire [0:0] csa_component17_fa10_xor1;
  wire [0:0] csa_component17_fa10_or0;
  wire [0:0] csa_component17_fa11_xor1;
  wire [0:0] csa_component17_fa11_or0;
  wire [0:0] csa_component17_fa12_xor1;
  wire [0:0] csa_component17_fa12_or0;
  wire [0:0] csa_component17_fa13_xor1;
  wire [0:0] csa_component17_fa13_or0;
  wire [0:0] csa_component17_fa14_xor1;
  wire [0:0] csa_component17_fa14_or0;
  wire [0:0] csa_component17_fa15_xor1;
  wire [0:0] csa_component17_fa15_or0;
  wire [0:0] csa_component17_fa16_xor1;
  wire [0:0] csa_component17_fa16_or0;

  fa fa_csa_component17_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component17_fa0_xor1), .fa_or0(csa_component17_fa0_or0));
  fa fa_csa_component17_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component17_fa1_xor1), .fa_or0(csa_component17_fa1_or0));
  fa fa_csa_component17_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component17_fa2_xor1), .fa_or0(csa_component17_fa2_or0));
  fa fa_csa_component17_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component17_fa3_xor1), .fa_or0(csa_component17_fa3_or0));
  fa fa_csa_component17_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component17_fa4_xor1), .fa_or0(csa_component17_fa4_or0));
  fa fa_csa_component17_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component17_fa5_xor1), .fa_or0(csa_component17_fa5_or0));
  fa fa_csa_component17_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component17_fa6_xor1), .fa_or0(csa_component17_fa6_or0));
  fa fa_csa_component17_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component17_fa7_xor1), .fa_or0(csa_component17_fa7_or0));
  fa fa_csa_component17_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component17_fa8_xor1), .fa_or0(csa_component17_fa8_or0));
  fa fa_csa_component17_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component17_fa9_xor1), .fa_or0(csa_component17_fa9_or0));
  fa fa_csa_component17_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component17_fa10_xor1), .fa_or0(csa_component17_fa10_or0));
  fa fa_csa_component17_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component17_fa11_xor1), .fa_or0(csa_component17_fa11_or0));
  fa fa_csa_component17_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component17_fa12_xor1), .fa_or0(csa_component17_fa12_or0));
  fa fa_csa_component17_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component17_fa13_xor1), .fa_or0(csa_component17_fa13_or0));
  fa fa_csa_component17_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component17_fa14_xor1), .fa_or0(csa_component17_fa14_or0));
  fa fa_csa_component17_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component17_fa15_xor1), .fa_or0(csa_component17_fa15_or0));
  fa fa_csa_component17_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component17_fa16_xor1), .fa_or0(csa_component17_fa16_or0));

  assign csa_component17_out[0] = csa_component17_fa0_xor1[0];
  assign csa_component17_out[1] = csa_component17_fa1_xor1[0];
  assign csa_component17_out[2] = csa_component17_fa2_xor1[0];
  assign csa_component17_out[3] = csa_component17_fa3_xor1[0];
  assign csa_component17_out[4] = csa_component17_fa4_xor1[0];
  assign csa_component17_out[5] = csa_component17_fa5_xor1[0];
  assign csa_component17_out[6] = csa_component17_fa6_xor1[0];
  assign csa_component17_out[7] = csa_component17_fa7_xor1[0];
  assign csa_component17_out[8] = csa_component17_fa8_xor1[0];
  assign csa_component17_out[9] = csa_component17_fa9_xor1[0];
  assign csa_component17_out[10] = csa_component17_fa10_xor1[0];
  assign csa_component17_out[11] = csa_component17_fa11_xor1[0];
  assign csa_component17_out[12] = csa_component17_fa12_xor1[0];
  assign csa_component17_out[13] = csa_component17_fa13_xor1[0];
  assign csa_component17_out[14] = csa_component17_fa14_xor1[0];
  assign csa_component17_out[15] = csa_component17_fa15_xor1[0];
  assign csa_component17_out[16] = csa_component17_fa16_xor1[0];
  assign csa_component17_out[17] = 1'b0;
  assign csa_component17_out[18] = 1'b0;
  assign csa_component17_out[19] = csa_component17_fa0_or0[0];
  assign csa_component17_out[20] = csa_component17_fa1_or0[0];
  assign csa_component17_out[21] = csa_component17_fa2_or0[0];
  assign csa_component17_out[22] = csa_component17_fa3_or0[0];
  assign csa_component17_out[23] = csa_component17_fa4_or0[0];
  assign csa_component17_out[24] = csa_component17_fa5_or0[0];
  assign csa_component17_out[25] = csa_component17_fa6_or0[0];
  assign csa_component17_out[26] = csa_component17_fa7_or0[0];
  assign csa_component17_out[27] = csa_component17_fa8_or0[0];
  assign csa_component17_out[28] = csa_component17_fa9_or0[0];
  assign csa_component17_out[29] = csa_component17_fa10_or0[0];
  assign csa_component17_out[30] = csa_component17_fa11_or0[0];
  assign csa_component17_out[31] = csa_component17_fa12_or0[0];
  assign csa_component17_out[32] = csa_component17_fa13_or0[0];
  assign csa_component17_out[33] = csa_component17_fa14_or0[0];
  assign csa_component17_out[34] = csa_component17_fa15_or0[0];
  assign csa_component17_out[35] = csa_component17_fa16_or0[0];
endmodule

module csa_component20(input [19:0] a, input [19:0] b, input [19:0] c, output [41:0] csa_component20_out);
  wire [0:0] csa_component20_fa0_xor1;
  wire [0:0] csa_component20_fa0_or0;
  wire [0:0] csa_component20_fa1_xor1;
  wire [0:0] csa_component20_fa1_or0;
  wire [0:0] csa_component20_fa2_xor1;
  wire [0:0] csa_component20_fa2_or0;
  wire [0:0] csa_component20_fa3_xor1;
  wire [0:0] csa_component20_fa3_or0;
  wire [0:0] csa_component20_fa4_xor1;
  wire [0:0] csa_component20_fa4_or0;
  wire [0:0] csa_component20_fa5_xor1;
  wire [0:0] csa_component20_fa5_or0;
  wire [0:0] csa_component20_fa6_xor1;
  wire [0:0] csa_component20_fa6_or0;
  wire [0:0] csa_component20_fa7_xor1;
  wire [0:0] csa_component20_fa7_or0;
  wire [0:0] csa_component20_fa8_xor1;
  wire [0:0] csa_component20_fa8_or0;
  wire [0:0] csa_component20_fa9_xor1;
  wire [0:0] csa_component20_fa9_or0;
  wire [0:0] csa_component20_fa10_xor1;
  wire [0:0] csa_component20_fa10_or0;
  wire [0:0] csa_component20_fa11_xor1;
  wire [0:0] csa_component20_fa11_or0;
  wire [0:0] csa_component20_fa12_xor1;
  wire [0:0] csa_component20_fa12_or0;
  wire [0:0] csa_component20_fa13_xor1;
  wire [0:0] csa_component20_fa13_or0;
  wire [0:0] csa_component20_fa14_xor1;
  wire [0:0] csa_component20_fa14_or0;
  wire [0:0] csa_component20_fa15_xor1;
  wire [0:0] csa_component20_fa15_or0;
  wire [0:0] csa_component20_fa16_xor1;
  wire [0:0] csa_component20_fa16_or0;
  wire [0:0] csa_component20_fa17_xor1;
  wire [0:0] csa_component20_fa17_or0;
  wire [0:0] csa_component20_fa18_xor1;
  wire [0:0] csa_component20_fa18_or0;
  wire [0:0] csa_component20_fa19_xor1;
  wire [0:0] csa_component20_fa19_or0;

  fa fa_csa_component20_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component20_fa0_xor1), .fa_or0(csa_component20_fa0_or0));
  fa fa_csa_component20_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component20_fa1_xor1), .fa_or0(csa_component20_fa1_or0));
  fa fa_csa_component20_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component20_fa2_xor1), .fa_or0(csa_component20_fa2_or0));
  fa fa_csa_component20_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component20_fa3_xor1), .fa_or0(csa_component20_fa3_or0));
  fa fa_csa_component20_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component20_fa4_xor1), .fa_or0(csa_component20_fa4_or0));
  fa fa_csa_component20_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component20_fa5_xor1), .fa_or0(csa_component20_fa5_or0));
  fa fa_csa_component20_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component20_fa6_xor1), .fa_or0(csa_component20_fa6_or0));
  fa fa_csa_component20_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component20_fa7_xor1), .fa_or0(csa_component20_fa7_or0));
  fa fa_csa_component20_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component20_fa8_xor1), .fa_or0(csa_component20_fa8_or0));
  fa fa_csa_component20_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component20_fa9_xor1), .fa_or0(csa_component20_fa9_or0));
  fa fa_csa_component20_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component20_fa10_xor1), .fa_or0(csa_component20_fa10_or0));
  fa fa_csa_component20_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component20_fa11_xor1), .fa_or0(csa_component20_fa11_or0));
  fa fa_csa_component20_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component20_fa12_xor1), .fa_or0(csa_component20_fa12_or0));
  fa fa_csa_component20_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component20_fa13_xor1), .fa_or0(csa_component20_fa13_or0));
  fa fa_csa_component20_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component20_fa14_xor1), .fa_or0(csa_component20_fa14_or0));
  fa fa_csa_component20_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component20_fa15_xor1), .fa_or0(csa_component20_fa15_or0));
  fa fa_csa_component20_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component20_fa16_xor1), .fa_or0(csa_component20_fa16_or0));
  fa fa_csa_component20_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component20_fa17_xor1), .fa_or0(csa_component20_fa17_or0));
  fa fa_csa_component20_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component20_fa18_xor1), .fa_or0(csa_component20_fa18_or0));
  fa fa_csa_component20_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component20_fa19_xor1), .fa_or0(csa_component20_fa19_or0));

  assign csa_component20_out[0] = csa_component20_fa0_xor1[0];
  assign csa_component20_out[1] = csa_component20_fa1_xor1[0];
  assign csa_component20_out[2] = csa_component20_fa2_xor1[0];
  assign csa_component20_out[3] = csa_component20_fa3_xor1[0];
  assign csa_component20_out[4] = csa_component20_fa4_xor1[0];
  assign csa_component20_out[5] = csa_component20_fa5_xor1[0];
  assign csa_component20_out[6] = csa_component20_fa6_xor1[0];
  assign csa_component20_out[7] = csa_component20_fa7_xor1[0];
  assign csa_component20_out[8] = csa_component20_fa8_xor1[0];
  assign csa_component20_out[9] = csa_component20_fa9_xor1[0];
  assign csa_component20_out[10] = csa_component20_fa10_xor1[0];
  assign csa_component20_out[11] = csa_component20_fa11_xor1[0];
  assign csa_component20_out[12] = csa_component20_fa12_xor1[0];
  assign csa_component20_out[13] = csa_component20_fa13_xor1[0];
  assign csa_component20_out[14] = csa_component20_fa14_xor1[0];
  assign csa_component20_out[15] = csa_component20_fa15_xor1[0];
  assign csa_component20_out[16] = csa_component20_fa16_xor1[0];
  assign csa_component20_out[17] = csa_component20_fa17_xor1[0];
  assign csa_component20_out[18] = csa_component20_fa18_xor1[0];
  assign csa_component20_out[19] = csa_component20_fa19_xor1[0];
  assign csa_component20_out[20] = 1'b0;
  assign csa_component20_out[21] = 1'b0;
  assign csa_component20_out[22] = csa_component20_fa0_or0[0];
  assign csa_component20_out[23] = csa_component20_fa1_or0[0];
  assign csa_component20_out[24] = csa_component20_fa2_or0[0];
  assign csa_component20_out[25] = csa_component20_fa3_or0[0];
  assign csa_component20_out[26] = csa_component20_fa4_or0[0];
  assign csa_component20_out[27] = csa_component20_fa5_or0[0];
  assign csa_component20_out[28] = csa_component20_fa6_or0[0];
  assign csa_component20_out[29] = csa_component20_fa7_or0[0];
  assign csa_component20_out[30] = csa_component20_fa8_or0[0];
  assign csa_component20_out[31] = csa_component20_fa9_or0[0];
  assign csa_component20_out[32] = csa_component20_fa10_or0[0];
  assign csa_component20_out[33] = csa_component20_fa11_or0[0];
  assign csa_component20_out[34] = csa_component20_fa12_or0[0];
  assign csa_component20_out[35] = csa_component20_fa13_or0[0];
  assign csa_component20_out[36] = csa_component20_fa14_or0[0];
  assign csa_component20_out[37] = csa_component20_fa15_or0[0];
  assign csa_component20_out[38] = csa_component20_fa16_or0[0];
  assign csa_component20_out[39] = csa_component20_fa17_or0[0];
  assign csa_component20_out[40] = csa_component20_fa18_or0[0];
  assign csa_component20_out[41] = csa_component20_fa19_or0[0];
endmodule

module csa_component23(input [22:0] a, input [22:0] b, input [22:0] c, output [47:0] csa_component23_out);
  wire [0:0] csa_component23_fa0_xor1;
  wire [0:0] csa_component23_fa0_or0;
  wire [0:0] csa_component23_fa1_xor1;
  wire [0:0] csa_component23_fa1_or0;
  wire [0:0] csa_component23_fa2_xor1;
  wire [0:0] csa_component23_fa2_or0;
  wire [0:0] csa_component23_fa3_xor1;
  wire [0:0] csa_component23_fa3_or0;
  wire [0:0] csa_component23_fa4_xor1;
  wire [0:0] csa_component23_fa4_or0;
  wire [0:0] csa_component23_fa5_xor1;
  wire [0:0] csa_component23_fa5_or0;
  wire [0:0] csa_component23_fa6_xor1;
  wire [0:0] csa_component23_fa6_or0;
  wire [0:0] csa_component23_fa7_xor1;
  wire [0:0] csa_component23_fa7_or0;
  wire [0:0] csa_component23_fa8_xor1;
  wire [0:0] csa_component23_fa8_or0;
  wire [0:0] csa_component23_fa9_xor1;
  wire [0:0] csa_component23_fa9_or0;
  wire [0:0] csa_component23_fa10_xor1;
  wire [0:0] csa_component23_fa10_or0;
  wire [0:0] csa_component23_fa11_xor1;
  wire [0:0] csa_component23_fa11_or0;
  wire [0:0] csa_component23_fa12_xor1;
  wire [0:0] csa_component23_fa12_or0;
  wire [0:0] csa_component23_fa13_xor1;
  wire [0:0] csa_component23_fa13_or0;
  wire [0:0] csa_component23_fa14_xor1;
  wire [0:0] csa_component23_fa14_or0;
  wire [0:0] csa_component23_fa15_xor1;
  wire [0:0] csa_component23_fa15_or0;
  wire [0:0] csa_component23_fa16_xor1;
  wire [0:0] csa_component23_fa16_or0;
  wire [0:0] csa_component23_fa17_xor1;
  wire [0:0] csa_component23_fa17_or0;
  wire [0:0] csa_component23_fa18_xor1;
  wire [0:0] csa_component23_fa18_or0;
  wire [0:0] csa_component23_fa19_xor1;
  wire [0:0] csa_component23_fa19_or0;
  wire [0:0] csa_component23_fa20_xor1;
  wire [0:0] csa_component23_fa20_or0;
  wire [0:0] csa_component23_fa21_xor1;
  wire [0:0] csa_component23_fa21_or0;
  wire [0:0] csa_component23_fa22_xor1;
  wire [0:0] csa_component23_fa22_or0;

  fa fa_csa_component23_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component23_fa0_xor1), .fa_or0(csa_component23_fa0_or0));
  fa fa_csa_component23_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component23_fa1_xor1), .fa_or0(csa_component23_fa1_or0));
  fa fa_csa_component23_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component23_fa2_xor1), .fa_or0(csa_component23_fa2_or0));
  fa fa_csa_component23_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component23_fa3_xor1), .fa_or0(csa_component23_fa3_or0));
  fa fa_csa_component23_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component23_fa4_xor1), .fa_or0(csa_component23_fa4_or0));
  fa fa_csa_component23_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component23_fa5_xor1), .fa_or0(csa_component23_fa5_or0));
  fa fa_csa_component23_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component23_fa6_xor1), .fa_or0(csa_component23_fa6_or0));
  fa fa_csa_component23_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component23_fa7_xor1), .fa_or0(csa_component23_fa7_or0));
  fa fa_csa_component23_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component23_fa8_xor1), .fa_or0(csa_component23_fa8_or0));
  fa fa_csa_component23_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component23_fa9_xor1), .fa_or0(csa_component23_fa9_or0));
  fa fa_csa_component23_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component23_fa10_xor1), .fa_or0(csa_component23_fa10_or0));
  fa fa_csa_component23_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component23_fa11_xor1), .fa_or0(csa_component23_fa11_or0));
  fa fa_csa_component23_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component23_fa12_xor1), .fa_or0(csa_component23_fa12_or0));
  fa fa_csa_component23_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component23_fa13_xor1), .fa_or0(csa_component23_fa13_or0));
  fa fa_csa_component23_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component23_fa14_xor1), .fa_or0(csa_component23_fa14_or0));
  fa fa_csa_component23_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component23_fa15_xor1), .fa_or0(csa_component23_fa15_or0));
  fa fa_csa_component23_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component23_fa16_xor1), .fa_or0(csa_component23_fa16_or0));
  fa fa_csa_component23_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component23_fa17_xor1), .fa_or0(csa_component23_fa17_or0));
  fa fa_csa_component23_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component23_fa18_xor1), .fa_or0(csa_component23_fa18_or0));
  fa fa_csa_component23_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component23_fa19_xor1), .fa_or0(csa_component23_fa19_or0));
  fa fa_csa_component23_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component23_fa20_xor1), .fa_or0(csa_component23_fa20_or0));
  fa fa_csa_component23_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component23_fa21_xor1), .fa_or0(csa_component23_fa21_or0));
  fa fa_csa_component23_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component23_fa22_xor1), .fa_or0(csa_component23_fa22_or0));

  assign csa_component23_out[0] = csa_component23_fa0_xor1[0];
  assign csa_component23_out[1] = csa_component23_fa1_xor1[0];
  assign csa_component23_out[2] = csa_component23_fa2_xor1[0];
  assign csa_component23_out[3] = csa_component23_fa3_xor1[0];
  assign csa_component23_out[4] = csa_component23_fa4_xor1[0];
  assign csa_component23_out[5] = csa_component23_fa5_xor1[0];
  assign csa_component23_out[6] = csa_component23_fa6_xor1[0];
  assign csa_component23_out[7] = csa_component23_fa7_xor1[0];
  assign csa_component23_out[8] = csa_component23_fa8_xor1[0];
  assign csa_component23_out[9] = csa_component23_fa9_xor1[0];
  assign csa_component23_out[10] = csa_component23_fa10_xor1[0];
  assign csa_component23_out[11] = csa_component23_fa11_xor1[0];
  assign csa_component23_out[12] = csa_component23_fa12_xor1[0];
  assign csa_component23_out[13] = csa_component23_fa13_xor1[0];
  assign csa_component23_out[14] = csa_component23_fa14_xor1[0];
  assign csa_component23_out[15] = csa_component23_fa15_xor1[0];
  assign csa_component23_out[16] = csa_component23_fa16_xor1[0];
  assign csa_component23_out[17] = csa_component23_fa17_xor1[0];
  assign csa_component23_out[18] = csa_component23_fa18_xor1[0];
  assign csa_component23_out[19] = csa_component23_fa19_xor1[0];
  assign csa_component23_out[20] = csa_component23_fa20_xor1[0];
  assign csa_component23_out[21] = csa_component23_fa21_xor1[0];
  assign csa_component23_out[22] = csa_component23_fa22_xor1[0];
  assign csa_component23_out[23] = 1'b0;
  assign csa_component23_out[24] = 1'b0;
  assign csa_component23_out[25] = csa_component23_fa0_or0[0];
  assign csa_component23_out[26] = csa_component23_fa1_or0[0];
  assign csa_component23_out[27] = csa_component23_fa2_or0[0];
  assign csa_component23_out[28] = csa_component23_fa3_or0[0];
  assign csa_component23_out[29] = csa_component23_fa4_or0[0];
  assign csa_component23_out[30] = csa_component23_fa5_or0[0];
  assign csa_component23_out[31] = csa_component23_fa6_or0[0];
  assign csa_component23_out[32] = csa_component23_fa7_or0[0];
  assign csa_component23_out[33] = csa_component23_fa8_or0[0];
  assign csa_component23_out[34] = csa_component23_fa9_or0[0];
  assign csa_component23_out[35] = csa_component23_fa10_or0[0];
  assign csa_component23_out[36] = csa_component23_fa11_or0[0];
  assign csa_component23_out[37] = csa_component23_fa12_or0[0];
  assign csa_component23_out[38] = csa_component23_fa13_or0[0];
  assign csa_component23_out[39] = csa_component23_fa14_or0[0];
  assign csa_component23_out[40] = csa_component23_fa15_or0[0];
  assign csa_component23_out[41] = csa_component23_fa16_or0[0];
  assign csa_component23_out[42] = csa_component23_fa17_or0[0];
  assign csa_component23_out[43] = csa_component23_fa18_or0[0];
  assign csa_component23_out[44] = csa_component23_fa19_or0[0];
  assign csa_component23_out[45] = csa_component23_fa20_or0[0];
  assign csa_component23_out[46] = csa_component23_fa21_or0[0];
  assign csa_component23_out[47] = csa_component23_fa22_or0[0];
endmodule

module csa_component18(input [17:0] a, input [17:0] b, input [17:0] c, output [37:0] csa_component18_out);
  wire [0:0] csa_component18_fa0_xor1;
  wire [0:0] csa_component18_fa0_or0;
  wire [0:0] csa_component18_fa1_xor1;
  wire [0:0] csa_component18_fa1_or0;
  wire [0:0] csa_component18_fa2_xor1;
  wire [0:0] csa_component18_fa2_or0;
  wire [0:0] csa_component18_fa3_xor1;
  wire [0:0] csa_component18_fa3_or0;
  wire [0:0] csa_component18_fa4_xor1;
  wire [0:0] csa_component18_fa4_or0;
  wire [0:0] csa_component18_fa5_xor1;
  wire [0:0] csa_component18_fa5_or0;
  wire [0:0] csa_component18_fa6_xor1;
  wire [0:0] csa_component18_fa6_or0;
  wire [0:0] csa_component18_fa7_xor1;
  wire [0:0] csa_component18_fa7_or0;
  wire [0:0] csa_component18_fa8_xor1;
  wire [0:0] csa_component18_fa8_or0;
  wire [0:0] csa_component18_fa9_xor1;
  wire [0:0] csa_component18_fa9_or0;
  wire [0:0] csa_component18_fa10_xor1;
  wire [0:0] csa_component18_fa10_or0;
  wire [0:0] csa_component18_fa11_xor1;
  wire [0:0] csa_component18_fa11_or0;
  wire [0:0] csa_component18_fa12_xor1;
  wire [0:0] csa_component18_fa12_or0;
  wire [0:0] csa_component18_fa13_xor1;
  wire [0:0] csa_component18_fa13_or0;
  wire [0:0] csa_component18_fa14_xor1;
  wire [0:0] csa_component18_fa14_or0;
  wire [0:0] csa_component18_fa15_xor1;
  wire [0:0] csa_component18_fa15_or0;
  wire [0:0] csa_component18_fa16_xor1;
  wire [0:0] csa_component18_fa16_or0;
  wire [0:0] csa_component18_fa17_xor1;
  wire [0:0] csa_component18_fa17_or0;

  fa fa_csa_component18_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component18_fa0_xor1), .fa_or0(csa_component18_fa0_or0));
  fa fa_csa_component18_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component18_fa1_xor1), .fa_or0(csa_component18_fa1_or0));
  fa fa_csa_component18_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component18_fa2_xor1), .fa_or0(csa_component18_fa2_or0));
  fa fa_csa_component18_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component18_fa3_xor1), .fa_or0(csa_component18_fa3_or0));
  fa fa_csa_component18_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component18_fa4_xor1), .fa_or0(csa_component18_fa4_or0));
  fa fa_csa_component18_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component18_fa5_xor1), .fa_or0(csa_component18_fa5_or0));
  fa fa_csa_component18_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component18_fa6_xor1), .fa_or0(csa_component18_fa6_or0));
  fa fa_csa_component18_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component18_fa7_xor1), .fa_or0(csa_component18_fa7_or0));
  fa fa_csa_component18_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component18_fa8_xor1), .fa_or0(csa_component18_fa8_or0));
  fa fa_csa_component18_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component18_fa9_xor1), .fa_or0(csa_component18_fa9_or0));
  fa fa_csa_component18_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component18_fa10_xor1), .fa_or0(csa_component18_fa10_or0));
  fa fa_csa_component18_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component18_fa11_xor1), .fa_or0(csa_component18_fa11_or0));
  fa fa_csa_component18_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component18_fa12_xor1), .fa_or0(csa_component18_fa12_or0));
  fa fa_csa_component18_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component18_fa13_xor1), .fa_or0(csa_component18_fa13_or0));
  fa fa_csa_component18_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component18_fa14_xor1), .fa_or0(csa_component18_fa14_or0));
  fa fa_csa_component18_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component18_fa15_xor1), .fa_or0(csa_component18_fa15_or0));
  fa fa_csa_component18_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component18_fa16_xor1), .fa_or0(csa_component18_fa16_or0));
  fa fa_csa_component18_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component18_fa17_xor1), .fa_or0(csa_component18_fa17_or0));

  assign csa_component18_out[0] = csa_component18_fa0_xor1[0];
  assign csa_component18_out[1] = csa_component18_fa1_xor1[0];
  assign csa_component18_out[2] = csa_component18_fa2_xor1[0];
  assign csa_component18_out[3] = csa_component18_fa3_xor1[0];
  assign csa_component18_out[4] = csa_component18_fa4_xor1[0];
  assign csa_component18_out[5] = csa_component18_fa5_xor1[0];
  assign csa_component18_out[6] = csa_component18_fa6_xor1[0];
  assign csa_component18_out[7] = csa_component18_fa7_xor1[0];
  assign csa_component18_out[8] = csa_component18_fa8_xor1[0];
  assign csa_component18_out[9] = csa_component18_fa9_xor1[0];
  assign csa_component18_out[10] = csa_component18_fa10_xor1[0];
  assign csa_component18_out[11] = csa_component18_fa11_xor1[0];
  assign csa_component18_out[12] = csa_component18_fa12_xor1[0];
  assign csa_component18_out[13] = csa_component18_fa13_xor1[0];
  assign csa_component18_out[14] = csa_component18_fa14_xor1[0];
  assign csa_component18_out[15] = csa_component18_fa15_xor1[0];
  assign csa_component18_out[16] = csa_component18_fa16_xor1[0];
  assign csa_component18_out[17] = csa_component18_fa17_xor1[0];
  assign csa_component18_out[18] = 1'b0;
  assign csa_component18_out[19] = 1'b0;
  assign csa_component18_out[20] = csa_component18_fa0_or0[0];
  assign csa_component18_out[21] = csa_component18_fa1_or0[0];
  assign csa_component18_out[22] = csa_component18_fa2_or0[0];
  assign csa_component18_out[23] = csa_component18_fa3_or0[0];
  assign csa_component18_out[24] = csa_component18_fa4_or0[0];
  assign csa_component18_out[25] = csa_component18_fa5_or0[0];
  assign csa_component18_out[26] = csa_component18_fa6_or0[0];
  assign csa_component18_out[27] = csa_component18_fa7_or0[0];
  assign csa_component18_out[28] = csa_component18_fa8_or0[0];
  assign csa_component18_out[29] = csa_component18_fa9_or0[0];
  assign csa_component18_out[30] = csa_component18_fa10_or0[0];
  assign csa_component18_out[31] = csa_component18_fa11_or0[0];
  assign csa_component18_out[32] = csa_component18_fa12_or0[0];
  assign csa_component18_out[33] = csa_component18_fa13_or0[0];
  assign csa_component18_out[34] = csa_component18_fa14_or0[0];
  assign csa_component18_out[35] = csa_component18_fa15_or0[0];
  assign csa_component18_out[36] = csa_component18_fa16_or0[0];
  assign csa_component18_out[37] = csa_component18_fa17_or0[0];
endmodule

module csa_component21(input [20:0] a, input [20:0] b, input [20:0] c, output [43:0] csa_component21_out);
  wire [0:0] csa_component21_fa0_xor1;
  wire [0:0] csa_component21_fa0_or0;
  wire [0:0] csa_component21_fa1_xor1;
  wire [0:0] csa_component21_fa1_or0;
  wire [0:0] csa_component21_fa2_xor1;
  wire [0:0] csa_component21_fa2_or0;
  wire [0:0] csa_component21_fa3_xor1;
  wire [0:0] csa_component21_fa3_or0;
  wire [0:0] csa_component21_fa4_xor1;
  wire [0:0] csa_component21_fa4_or0;
  wire [0:0] csa_component21_fa5_xor1;
  wire [0:0] csa_component21_fa5_or0;
  wire [0:0] csa_component21_fa6_xor1;
  wire [0:0] csa_component21_fa6_or0;
  wire [0:0] csa_component21_fa7_xor1;
  wire [0:0] csa_component21_fa7_or0;
  wire [0:0] csa_component21_fa8_xor1;
  wire [0:0] csa_component21_fa8_or0;
  wire [0:0] csa_component21_fa9_xor1;
  wire [0:0] csa_component21_fa9_or0;
  wire [0:0] csa_component21_fa10_xor1;
  wire [0:0] csa_component21_fa10_or0;
  wire [0:0] csa_component21_fa11_xor1;
  wire [0:0] csa_component21_fa11_or0;
  wire [0:0] csa_component21_fa12_xor1;
  wire [0:0] csa_component21_fa12_or0;
  wire [0:0] csa_component21_fa13_xor1;
  wire [0:0] csa_component21_fa13_or0;
  wire [0:0] csa_component21_fa14_xor1;
  wire [0:0] csa_component21_fa14_or0;
  wire [0:0] csa_component21_fa15_xor1;
  wire [0:0] csa_component21_fa15_or0;
  wire [0:0] csa_component21_fa16_xor1;
  wire [0:0] csa_component21_fa16_or0;
  wire [0:0] csa_component21_fa17_xor1;
  wire [0:0] csa_component21_fa17_or0;
  wire [0:0] csa_component21_fa18_xor1;
  wire [0:0] csa_component21_fa18_or0;
  wire [0:0] csa_component21_fa19_xor1;
  wire [0:0] csa_component21_fa19_or0;
  wire [0:0] csa_component21_fa20_xor1;
  wire [0:0] csa_component21_fa20_or0;

  fa fa_csa_component21_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component21_fa0_xor1), .fa_or0(csa_component21_fa0_or0));
  fa fa_csa_component21_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component21_fa1_xor1), .fa_or0(csa_component21_fa1_or0));
  fa fa_csa_component21_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component21_fa2_xor1), .fa_or0(csa_component21_fa2_or0));
  fa fa_csa_component21_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component21_fa3_xor1), .fa_or0(csa_component21_fa3_or0));
  fa fa_csa_component21_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component21_fa4_xor1), .fa_or0(csa_component21_fa4_or0));
  fa fa_csa_component21_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component21_fa5_xor1), .fa_or0(csa_component21_fa5_or0));
  fa fa_csa_component21_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component21_fa6_xor1), .fa_or0(csa_component21_fa6_or0));
  fa fa_csa_component21_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component21_fa7_xor1), .fa_or0(csa_component21_fa7_or0));
  fa fa_csa_component21_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component21_fa8_xor1), .fa_or0(csa_component21_fa8_or0));
  fa fa_csa_component21_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component21_fa9_xor1), .fa_or0(csa_component21_fa9_or0));
  fa fa_csa_component21_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component21_fa10_xor1), .fa_or0(csa_component21_fa10_or0));
  fa fa_csa_component21_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component21_fa11_xor1), .fa_or0(csa_component21_fa11_or0));
  fa fa_csa_component21_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component21_fa12_xor1), .fa_or0(csa_component21_fa12_or0));
  fa fa_csa_component21_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component21_fa13_xor1), .fa_or0(csa_component21_fa13_or0));
  fa fa_csa_component21_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component21_fa14_xor1), .fa_or0(csa_component21_fa14_or0));
  fa fa_csa_component21_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component21_fa15_xor1), .fa_or0(csa_component21_fa15_or0));
  fa fa_csa_component21_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component21_fa16_xor1), .fa_or0(csa_component21_fa16_or0));
  fa fa_csa_component21_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component21_fa17_xor1), .fa_or0(csa_component21_fa17_or0));
  fa fa_csa_component21_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component21_fa18_xor1), .fa_or0(csa_component21_fa18_or0));
  fa fa_csa_component21_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component21_fa19_xor1), .fa_or0(csa_component21_fa19_or0));
  fa fa_csa_component21_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component21_fa20_xor1), .fa_or0(csa_component21_fa20_or0));

  assign csa_component21_out[0] = csa_component21_fa0_xor1[0];
  assign csa_component21_out[1] = csa_component21_fa1_xor1[0];
  assign csa_component21_out[2] = csa_component21_fa2_xor1[0];
  assign csa_component21_out[3] = csa_component21_fa3_xor1[0];
  assign csa_component21_out[4] = csa_component21_fa4_xor1[0];
  assign csa_component21_out[5] = csa_component21_fa5_xor1[0];
  assign csa_component21_out[6] = csa_component21_fa6_xor1[0];
  assign csa_component21_out[7] = csa_component21_fa7_xor1[0];
  assign csa_component21_out[8] = csa_component21_fa8_xor1[0];
  assign csa_component21_out[9] = csa_component21_fa9_xor1[0];
  assign csa_component21_out[10] = csa_component21_fa10_xor1[0];
  assign csa_component21_out[11] = csa_component21_fa11_xor1[0];
  assign csa_component21_out[12] = csa_component21_fa12_xor1[0];
  assign csa_component21_out[13] = csa_component21_fa13_xor1[0];
  assign csa_component21_out[14] = csa_component21_fa14_xor1[0];
  assign csa_component21_out[15] = csa_component21_fa15_xor1[0];
  assign csa_component21_out[16] = csa_component21_fa16_xor1[0];
  assign csa_component21_out[17] = csa_component21_fa17_xor1[0];
  assign csa_component21_out[18] = csa_component21_fa18_xor1[0];
  assign csa_component21_out[19] = csa_component21_fa19_xor1[0];
  assign csa_component21_out[20] = csa_component21_fa20_xor1[0];
  assign csa_component21_out[21] = 1'b0;
  assign csa_component21_out[22] = 1'b0;
  assign csa_component21_out[23] = csa_component21_fa0_or0[0];
  assign csa_component21_out[24] = csa_component21_fa1_or0[0];
  assign csa_component21_out[25] = csa_component21_fa2_or0[0];
  assign csa_component21_out[26] = csa_component21_fa3_or0[0];
  assign csa_component21_out[27] = csa_component21_fa4_or0[0];
  assign csa_component21_out[28] = csa_component21_fa5_or0[0];
  assign csa_component21_out[29] = csa_component21_fa6_or0[0];
  assign csa_component21_out[30] = csa_component21_fa7_or0[0];
  assign csa_component21_out[31] = csa_component21_fa8_or0[0];
  assign csa_component21_out[32] = csa_component21_fa9_or0[0];
  assign csa_component21_out[33] = csa_component21_fa10_or0[0];
  assign csa_component21_out[34] = csa_component21_fa11_or0[0];
  assign csa_component21_out[35] = csa_component21_fa12_or0[0];
  assign csa_component21_out[36] = csa_component21_fa13_or0[0];
  assign csa_component21_out[37] = csa_component21_fa14_or0[0];
  assign csa_component21_out[38] = csa_component21_fa15_or0[0];
  assign csa_component21_out[39] = csa_component21_fa16_or0[0];
  assign csa_component21_out[40] = csa_component21_fa17_or0[0];
  assign csa_component21_out[41] = csa_component21_fa18_or0[0];
  assign csa_component21_out[42] = csa_component21_fa19_or0[0];
  assign csa_component21_out[43] = csa_component21_fa20_or0[0];
endmodule

module csa_component22(input [21:0] a, input [21:0] b, input [21:0] c, output [45:0] csa_component22_out);
  wire [0:0] csa_component22_fa0_xor1;
  wire [0:0] csa_component22_fa0_or0;
  wire [0:0] csa_component22_fa1_xor1;
  wire [0:0] csa_component22_fa1_or0;
  wire [0:0] csa_component22_fa2_xor1;
  wire [0:0] csa_component22_fa2_or0;
  wire [0:0] csa_component22_fa3_xor1;
  wire [0:0] csa_component22_fa3_or0;
  wire [0:0] csa_component22_fa4_xor1;
  wire [0:0] csa_component22_fa4_or0;
  wire [0:0] csa_component22_fa5_xor1;
  wire [0:0] csa_component22_fa5_or0;
  wire [0:0] csa_component22_fa6_xor1;
  wire [0:0] csa_component22_fa6_or0;
  wire [0:0] csa_component22_fa7_xor1;
  wire [0:0] csa_component22_fa7_or0;
  wire [0:0] csa_component22_fa8_xor1;
  wire [0:0] csa_component22_fa8_or0;
  wire [0:0] csa_component22_fa9_xor1;
  wire [0:0] csa_component22_fa9_or0;
  wire [0:0] csa_component22_fa10_xor1;
  wire [0:0] csa_component22_fa10_or0;
  wire [0:0] csa_component22_fa11_xor1;
  wire [0:0] csa_component22_fa11_or0;
  wire [0:0] csa_component22_fa12_xor1;
  wire [0:0] csa_component22_fa12_or0;
  wire [0:0] csa_component22_fa13_xor1;
  wire [0:0] csa_component22_fa13_or0;
  wire [0:0] csa_component22_fa14_xor1;
  wire [0:0] csa_component22_fa14_or0;
  wire [0:0] csa_component22_fa15_xor1;
  wire [0:0] csa_component22_fa15_or0;
  wire [0:0] csa_component22_fa16_xor1;
  wire [0:0] csa_component22_fa16_or0;
  wire [0:0] csa_component22_fa17_xor1;
  wire [0:0] csa_component22_fa17_or0;
  wire [0:0] csa_component22_fa18_xor1;
  wire [0:0] csa_component22_fa18_or0;
  wire [0:0] csa_component22_fa19_xor1;
  wire [0:0] csa_component22_fa19_or0;
  wire [0:0] csa_component22_fa20_xor1;
  wire [0:0] csa_component22_fa20_or0;
  wire [0:0] csa_component22_fa21_xor1;
  wire [0:0] csa_component22_fa21_or0;

  fa fa_csa_component22_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component22_fa0_xor1), .fa_or0(csa_component22_fa0_or0));
  fa fa_csa_component22_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component22_fa1_xor1), .fa_or0(csa_component22_fa1_or0));
  fa fa_csa_component22_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component22_fa2_xor1), .fa_or0(csa_component22_fa2_or0));
  fa fa_csa_component22_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component22_fa3_xor1), .fa_or0(csa_component22_fa3_or0));
  fa fa_csa_component22_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component22_fa4_xor1), .fa_or0(csa_component22_fa4_or0));
  fa fa_csa_component22_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component22_fa5_xor1), .fa_or0(csa_component22_fa5_or0));
  fa fa_csa_component22_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component22_fa6_xor1), .fa_or0(csa_component22_fa6_or0));
  fa fa_csa_component22_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component22_fa7_xor1), .fa_or0(csa_component22_fa7_or0));
  fa fa_csa_component22_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component22_fa8_xor1), .fa_or0(csa_component22_fa8_or0));
  fa fa_csa_component22_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component22_fa9_xor1), .fa_or0(csa_component22_fa9_or0));
  fa fa_csa_component22_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component22_fa10_xor1), .fa_or0(csa_component22_fa10_or0));
  fa fa_csa_component22_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component22_fa11_xor1), .fa_or0(csa_component22_fa11_or0));
  fa fa_csa_component22_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component22_fa12_xor1), .fa_or0(csa_component22_fa12_or0));
  fa fa_csa_component22_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component22_fa13_xor1), .fa_or0(csa_component22_fa13_or0));
  fa fa_csa_component22_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component22_fa14_xor1), .fa_or0(csa_component22_fa14_or0));
  fa fa_csa_component22_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component22_fa15_xor1), .fa_or0(csa_component22_fa15_or0));
  fa fa_csa_component22_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component22_fa16_xor1), .fa_or0(csa_component22_fa16_or0));
  fa fa_csa_component22_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component22_fa17_xor1), .fa_or0(csa_component22_fa17_or0));
  fa fa_csa_component22_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component22_fa18_xor1), .fa_or0(csa_component22_fa18_or0));
  fa fa_csa_component22_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component22_fa19_xor1), .fa_or0(csa_component22_fa19_or0));
  fa fa_csa_component22_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component22_fa20_xor1), .fa_or0(csa_component22_fa20_or0));
  fa fa_csa_component22_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component22_fa21_xor1), .fa_or0(csa_component22_fa21_or0));

  assign csa_component22_out[0] = csa_component22_fa0_xor1[0];
  assign csa_component22_out[1] = csa_component22_fa1_xor1[0];
  assign csa_component22_out[2] = csa_component22_fa2_xor1[0];
  assign csa_component22_out[3] = csa_component22_fa3_xor1[0];
  assign csa_component22_out[4] = csa_component22_fa4_xor1[0];
  assign csa_component22_out[5] = csa_component22_fa5_xor1[0];
  assign csa_component22_out[6] = csa_component22_fa6_xor1[0];
  assign csa_component22_out[7] = csa_component22_fa7_xor1[0];
  assign csa_component22_out[8] = csa_component22_fa8_xor1[0];
  assign csa_component22_out[9] = csa_component22_fa9_xor1[0];
  assign csa_component22_out[10] = csa_component22_fa10_xor1[0];
  assign csa_component22_out[11] = csa_component22_fa11_xor1[0];
  assign csa_component22_out[12] = csa_component22_fa12_xor1[0];
  assign csa_component22_out[13] = csa_component22_fa13_xor1[0];
  assign csa_component22_out[14] = csa_component22_fa14_xor1[0];
  assign csa_component22_out[15] = csa_component22_fa15_xor1[0];
  assign csa_component22_out[16] = csa_component22_fa16_xor1[0];
  assign csa_component22_out[17] = csa_component22_fa17_xor1[0];
  assign csa_component22_out[18] = csa_component22_fa18_xor1[0];
  assign csa_component22_out[19] = csa_component22_fa19_xor1[0];
  assign csa_component22_out[20] = csa_component22_fa20_xor1[0];
  assign csa_component22_out[21] = csa_component22_fa21_xor1[0];
  assign csa_component22_out[22] = 1'b0;
  assign csa_component22_out[23] = 1'b0;
  assign csa_component22_out[24] = csa_component22_fa0_or0[0];
  assign csa_component22_out[25] = csa_component22_fa1_or0[0];
  assign csa_component22_out[26] = csa_component22_fa2_or0[0];
  assign csa_component22_out[27] = csa_component22_fa3_or0[0];
  assign csa_component22_out[28] = csa_component22_fa4_or0[0];
  assign csa_component22_out[29] = csa_component22_fa5_or0[0];
  assign csa_component22_out[30] = csa_component22_fa6_or0[0];
  assign csa_component22_out[31] = csa_component22_fa7_or0[0];
  assign csa_component22_out[32] = csa_component22_fa8_or0[0];
  assign csa_component22_out[33] = csa_component22_fa9_or0[0];
  assign csa_component22_out[34] = csa_component22_fa10_or0[0];
  assign csa_component22_out[35] = csa_component22_fa11_or0[0];
  assign csa_component22_out[36] = csa_component22_fa12_or0[0];
  assign csa_component22_out[37] = csa_component22_fa13_or0[0];
  assign csa_component22_out[38] = csa_component22_fa14_or0[0];
  assign csa_component22_out[39] = csa_component22_fa15_or0[0];
  assign csa_component22_out[40] = csa_component22_fa16_or0[0];
  assign csa_component22_out[41] = csa_component22_fa17_or0[0];
  assign csa_component22_out[42] = csa_component22_fa18_or0[0];
  assign csa_component22_out[43] = csa_component22_fa19_or0[0];
  assign csa_component22_out[44] = csa_component22_fa20_or0[0];
  assign csa_component22_out[45] = csa_component22_fa21_or0[0];
endmodule

module csa_component24(input [23:0] a, input [23:0] b, input [23:0] c, output [49:0] csa_component24_out);
  wire [0:0] csa_component24_fa0_xor1;
  wire [0:0] csa_component24_fa0_or0;
  wire [0:0] csa_component24_fa1_xor1;
  wire [0:0] csa_component24_fa1_or0;
  wire [0:0] csa_component24_fa2_xor1;
  wire [0:0] csa_component24_fa2_or0;
  wire [0:0] csa_component24_fa3_xor1;
  wire [0:0] csa_component24_fa3_or0;
  wire [0:0] csa_component24_fa4_xor1;
  wire [0:0] csa_component24_fa4_or0;
  wire [0:0] csa_component24_fa5_xor1;
  wire [0:0] csa_component24_fa5_or0;
  wire [0:0] csa_component24_fa6_xor1;
  wire [0:0] csa_component24_fa6_or0;
  wire [0:0] csa_component24_fa7_xor1;
  wire [0:0] csa_component24_fa7_or0;
  wire [0:0] csa_component24_fa8_xor1;
  wire [0:0] csa_component24_fa8_or0;
  wire [0:0] csa_component24_fa9_xor1;
  wire [0:0] csa_component24_fa9_or0;
  wire [0:0] csa_component24_fa10_xor1;
  wire [0:0] csa_component24_fa10_or0;
  wire [0:0] csa_component24_fa11_xor1;
  wire [0:0] csa_component24_fa11_or0;
  wire [0:0] csa_component24_fa12_xor1;
  wire [0:0] csa_component24_fa12_or0;
  wire [0:0] csa_component24_fa13_xor1;
  wire [0:0] csa_component24_fa13_or0;
  wire [0:0] csa_component24_fa14_xor1;
  wire [0:0] csa_component24_fa14_or0;
  wire [0:0] csa_component24_fa15_xor1;
  wire [0:0] csa_component24_fa15_or0;
  wire [0:0] csa_component24_fa16_xor1;
  wire [0:0] csa_component24_fa16_or0;
  wire [0:0] csa_component24_fa17_xor1;
  wire [0:0] csa_component24_fa17_or0;
  wire [0:0] csa_component24_fa18_xor1;
  wire [0:0] csa_component24_fa18_or0;
  wire [0:0] csa_component24_fa19_xor1;
  wire [0:0] csa_component24_fa19_or0;
  wire [0:0] csa_component24_fa20_xor1;
  wire [0:0] csa_component24_fa20_or0;
  wire [0:0] csa_component24_fa21_xor1;
  wire [0:0] csa_component24_fa21_or0;
  wire [0:0] csa_component24_fa22_xor1;
  wire [0:0] csa_component24_fa22_or0;
  wire [0:0] csa_component24_fa23_xor1;
  wire [0:0] csa_component24_fa23_or0;

  fa fa_csa_component24_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component24_fa0_xor1), .fa_or0(csa_component24_fa0_or0));
  fa fa_csa_component24_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component24_fa1_xor1), .fa_or0(csa_component24_fa1_or0));
  fa fa_csa_component24_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component24_fa2_xor1), .fa_or0(csa_component24_fa2_or0));
  fa fa_csa_component24_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component24_fa3_xor1), .fa_or0(csa_component24_fa3_or0));
  fa fa_csa_component24_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component24_fa4_xor1), .fa_or0(csa_component24_fa4_or0));
  fa fa_csa_component24_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component24_fa5_xor1), .fa_or0(csa_component24_fa5_or0));
  fa fa_csa_component24_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component24_fa6_xor1), .fa_or0(csa_component24_fa6_or0));
  fa fa_csa_component24_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component24_fa7_xor1), .fa_or0(csa_component24_fa7_or0));
  fa fa_csa_component24_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component24_fa8_xor1), .fa_or0(csa_component24_fa8_or0));
  fa fa_csa_component24_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component24_fa9_xor1), .fa_or0(csa_component24_fa9_or0));
  fa fa_csa_component24_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component24_fa10_xor1), .fa_or0(csa_component24_fa10_or0));
  fa fa_csa_component24_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component24_fa11_xor1), .fa_or0(csa_component24_fa11_or0));
  fa fa_csa_component24_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component24_fa12_xor1), .fa_or0(csa_component24_fa12_or0));
  fa fa_csa_component24_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component24_fa13_xor1), .fa_or0(csa_component24_fa13_or0));
  fa fa_csa_component24_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component24_fa14_xor1), .fa_or0(csa_component24_fa14_or0));
  fa fa_csa_component24_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component24_fa15_xor1), .fa_or0(csa_component24_fa15_or0));
  fa fa_csa_component24_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component24_fa16_xor1), .fa_or0(csa_component24_fa16_or0));
  fa fa_csa_component24_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component24_fa17_xor1), .fa_or0(csa_component24_fa17_or0));
  fa fa_csa_component24_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component24_fa18_xor1), .fa_or0(csa_component24_fa18_or0));
  fa fa_csa_component24_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component24_fa19_xor1), .fa_or0(csa_component24_fa19_or0));
  fa fa_csa_component24_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component24_fa20_xor1), .fa_or0(csa_component24_fa20_or0));
  fa fa_csa_component24_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component24_fa21_xor1), .fa_or0(csa_component24_fa21_or0));
  fa fa_csa_component24_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component24_fa22_xor1), .fa_or0(csa_component24_fa22_or0));
  fa fa_csa_component24_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component24_fa23_xor1), .fa_or0(csa_component24_fa23_or0));

  assign csa_component24_out[0] = csa_component24_fa0_xor1[0];
  assign csa_component24_out[1] = csa_component24_fa1_xor1[0];
  assign csa_component24_out[2] = csa_component24_fa2_xor1[0];
  assign csa_component24_out[3] = csa_component24_fa3_xor1[0];
  assign csa_component24_out[4] = csa_component24_fa4_xor1[0];
  assign csa_component24_out[5] = csa_component24_fa5_xor1[0];
  assign csa_component24_out[6] = csa_component24_fa6_xor1[0];
  assign csa_component24_out[7] = csa_component24_fa7_xor1[0];
  assign csa_component24_out[8] = csa_component24_fa8_xor1[0];
  assign csa_component24_out[9] = csa_component24_fa9_xor1[0];
  assign csa_component24_out[10] = csa_component24_fa10_xor1[0];
  assign csa_component24_out[11] = csa_component24_fa11_xor1[0];
  assign csa_component24_out[12] = csa_component24_fa12_xor1[0];
  assign csa_component24_out[13] = csa_component24_fa13_xor1[0];
  assign csa_component24_out[14] = csa_component24_fa14_xor1[0];
  assign csa_component24_out[15] = csa_component24_fa15_xor1[0];
  assign csa_component24_out[16] = csa_component24_fa16_xor1[0];
  assign csa_component24_out[17] = csa_component24_fa17_xor1[0];
  assign csa_component24_out[18] = csa_component24_fa18_xor1[0];
  assign csa_component24_out[19] = csa_component24_fa19_xor1[0];
  assign csa_component24_out[20] = csa_component24_fa20_xor1[0];
  assign csa_component24_out[21] = csa_component24_fa21_xor1[0];
  assign csa_component24_out[22] = csa_component24_fa22_xor1[0];
  assign csa_component24_out[23] = csa_component24_fa23_xor1[0];
  assign csa_component24_out[24] = 1'b0;
  assign csa_component24_out[25] = 1'b0;
  assign csa_component24_out[26] = csa_component24_fa0_or0[0];
  assign csa_component24_out[27] = csa_component24_fa1_or0[0];
  assign csa_component24_out[28] = csa_component24_fa2_or0[0];
  assign csa_component24_out[29] = csa_component24_fa3_or0[0];
  assign csa_component24_out[30] = csa_component24_fa4_or0[0];
  assign csa_component24_out[31] = csa_component24_fa5_or0[0];
  assign csa_component24_out[32] = csa_component24_fa6_or0[0];
  assign csa_component24_out[33] = csa_component24_fa7_or0[0];
  assign csa_component24_out[34] = csa_component24_fa8_or0[0];
  assign csa_component24_out[35] = csa_component24_fa9_or0[0];
  assign csa_component24_out[36] = csa_component24_fa10_or0[0];
  assign csa_component24_out[37] = csa_component24_fa11_or0[0];
  assign csa_component24_out[38] = csa_component24_fa12_or0[0];
  assign csa_component24_out[39] = csa_component24_fa13_or0[0];
  assign csa_component24_out[40] = csa_component24_fa14_or0[0];
  assign csa_component24_out[41] = csa_component24_fa15_or0[0];
  assign csa_component24_out[42] = csa_component24_fa16_or0[0];
  assign csa_component24_out[43] = csa_component24_fa17_or0[0];
  assign csa_component24_out[44] = csa_component24_fa18_or0[0];
  assign csa_component24_out[45] = csa_component24_fa19_or0[0];
  assign csa_component24_out[46] = csa_component24_fa20_or0[0];
  assign csa_component24_out[47] = csa_component24_fa21_or0[0];
  assign csa_component24_out[48] = csa_component24_fa22_or0[0];
  assign csa_component24_out[49] = csa_component24_fa23_or0[0];
endmodule

module u_rca24(input [23:0] a, input [23:0] b, output [24:0] u_rca24_out);
  wire [0:0] u_rca24_ha_xor0;
  wire [0:0] u_rca24_ha_and0;
  wire [0:0] u_rca24_fa1_xor1;
  wire [0:0] u_rca24_fa1_or0;
  wire [0:0] u_rca24_fa2_xor1;
  wire [0:0] u_rca24_fa2_or0;
  wire [0:0] u_rca24_fa3_xor1;
  wire [0:0] u_rca24_fa3_or0;
  wire [0:0] u_rca24_fa4_xor1;
  wire [0:0] u_rca24_fa4_or0;
  wire [0:0] u_rca24_fa5_xor1;
  wire [0:0] u_rca24_fa5_or0;
  wire [0:0] u_rca24_fa6_xor1;
  wire [0:0] u_rca24_fa6_or0;
  wire [0:0] u_rca24_fa7_xor1;
  wire [0:0] u_rca24_fa7_or0;
  wire [0:0] u_rca24_fa8_xor1;
  wire [0:0] u_rca24_fa8_or0;
  wire [0:0] u_rca24_fa9_xor1;
  wire [0:0] u_rca24_fa9_or0;
  wire [0:0] u_rca24_fa10_xor1;
  wire [0:0] u_rca24_fa10_or0;
  wire [0:0] u_rca24_fa11_xor1;
  wire [0:0] u_rca24_fa11_or0;
  wire [0:0] u_rca24_fa12_xor1;
  wire [0:0] u_rca24_fa12_or0;
  wire [0:0] u_rca24_fa13_xor1;
  wire [0:0] u_rca24_fa13_or0;
  wire [0:0] u_rca24_fa14_xor1;
  wire [0:0] u_rca24_fa14_or0;
  wire [0:0] u_rca24_fa15_xor1;
  wire [0:0] u_rca24_fa15_or0;
  wire [0:0] u_rca24_fa16_xor1;
  wire [0:0] u_rca24_fa16_or0;
  wire [0:0] u_rca24_fa17_xor1;
  wire [0:0] u_rca24_fa17_or0;
  wire [0:0] u_rca24_fa18_xor1;
  wire [0:0] u_rca24_fa18_or0;
  wire [0:0] u_rca24_fa19_xor1;
  wire [0:0] u_rca24_fa19_or0;
  wire [0:0] u_rca24_fa20_xor1;
  wire [0:0] u_rca24_fa20_or0;
  wire [0:0] u_rca24_fa21_xor1;
  wire [0:0] u_rca24_fa21_or0;
  wire [0:0] u_rca24_fa22_xor1;
  wire [0:0] u_rca24_fa22_or0;
  wire [0:0] u_rca24_fa23_xor1;
  wire [0:0] u_rca24_fa23_or0;

  ha ha_u_rca24_ha_out(.a(a[0]), .b(b[0]), .ha_xor0(u_rca24_ha_xor0), .ha_and0(u_rca24_ha_and0));
  fa fa_u_rca24_fa1_out(.a(a[1]), .b(b[1]), .cin(u_rca24_ha_and0[0]), .fa_xor1(u_rca24_fa1_xor1), .fa_or0(u_rca24_fa1_or0));
  fa fa_u_rca24_fa2_out(.a(a[2]), .b(b[2]), .cin(u_rca24_fa1_or0[0]), .fa_xor1(u_rca24_fa2_xor1), .fa_or0(u_rca24_fa2_or0));
  fa fa_u_rca24_fa3_out(.a(a[3]), .b(b[3]), .cin(u_rca24_fa2_or0[0]), .fa_xor1(u_rca24_fa3_xor1), .fa_or0(u_rca24_fa3_or0));
  fa fa_u_rca24_fa4_out(.a(a[4]), .b(b[4]), .cin(u_rca24_fa3_or0[0]), .fa_xor1(u_rca24_fa4_xor1), .fa_or0(u_rca24_fa4_or0));
  fa fa_u_rca24_fa5_out(.a(a[5]), .b(b[5]), .cin(u_rca24_fa4_or0[0]), .fa_xor1(u_rca24_fa5_xor1), .fa_or0(u_rca24_fa5_or0));
  fa fa_u_rca24_fa6_out(.a(a[6]), .b(b[6]), .cin(u_rca24_fa5_or0[0]), .fa_xor1(u_rca24_fa6_xor1), .fa_or0(u_rca24_fa6_or0));
  fa fa_u_rca24_fa7_out(.a(a[7]), .b(b[7]), .cin(u_rca24_fa6_or0[0]), .fa_xor1(u_rca24_fa7_xor1), .fa_or0(u_rca24_fa7_or0));
  fa fa_u_rca24_fa8_out(.a(a[8]), .b(b[8]), .cin(u_rca24_fa7_or0[0]), .fa_xor1(u_rca24_fa8_xor1), .fa_or0(u_rca24_fa8_or0));
  fa fa_u_rca24_fa9_out(.a(a[9]), .b(b[9]), .cin(u_rca24_fa8_or0[0]), .fa_xor1(u_rca24_fa9_xor1), .fa_or0(u_rca24_fa9_or0));
  fa fa_u_rca24_fa10_out(.a(a[10]), .b(b[10]), .cin(u_rca24_fa9_or0[0]), .fa_xor1(u_rca24_fa10_xor1), .fa_or0(u_rca24_fa10_or0));
  fa fa_u_rca24_fa11_out(.a(a[11]), .b(b[11]), .cin(u_rca24_fa10_or0[0]), .fa_xor1(u_rca24_fa11_xor1), .fa_or0(u_rca24_fa11_or0));
  fa fa_u_rca24_fa12_out(.a(a[12]), .b(b[12]), .cin(u_rca24_fa11_or0[0]), .fa_xor1(u_rca24_fa12_xor1), .fa_or0(u_rca24_fa12_or0));
  fa fa_u_rca24_fa13_out(.a(a[13]), .b(b[13]), .cin(u_rca24_fa12_or0[0]), .fa_xor1(u_rca24_fa13_xor1), .fa_or0(u_rca24_fa13_or0));
  fa fa_u_rca24_fa14_out(.a(a[14]), .b(b[14]), .cin(u_rca24_fa13_or0[0]), .fa_xor1(u_rca24_fa14_xor1), .fa_or0(u_rca24_fa14_or0));
  fa fa_u_rca24_fa15_out(.a(a[15]), .b(b[15]), .cin(u_rca24_fa14_or0[0]), .fa_xor1(u_rca24_fa15_xor1), .fa_or0(u_rca24_fa15_or0));
  fa fa_u_rca24_fa16_out(.a(a[16]), .b(b[16]), .cin(u_rca24_fa15_or0[0]), .fa_xor1(u_rca24_fa16_xor1), .fa_or0(u_rca24_fa16_or0));
  fa fa_u_rca24_fa17_out(.a(a[17]), .b(b[17]), .cin(u_rca24_fa16_or0[0]), .fa_xor1(u_rca24_fa17_xor1), .fa_or0(u_rca24_fa17_or0));
  fa fa_u_rca24_fa18_out(.a(a[18]), .b(b[18]), .cin(u_rca24_fa17_or0[0]), .fa_xor1(u_rca24_fa18_xor1), .fa_or0(u_rca24_fa18_or0));
  fa fa_u_rca24_fa19_out(.a(a[19]), .b(b[19]), .cin(u_rca24_fa18_or0[0]), .fa_xor1(u_rca24_fa19_xor1), .fa_or0(u_rca24_fa19_or0));
  fa fa_u_rca24_fa20_out(.a(a[20]), .b(b[20]), .cin(u_rca24_fa19_or0[0]), .fa_xor1(u_rca24_fa20_xor1), .fa_or0(u_rca24_fa20_or0));
  fa fa_u_rca24_fa21_out(.a(a[21]), .b(b[21]), .cin(u_rca24_fa20_or0[0]), .fa_xor1(u_rca24_fa21_xor1), .fa_or0(u_rca24_fa21_or0));
  fa fa_u_rca24_fa22_out(.a(a[22]), .b(b[22]), .cin(u_rca24_fa21_or0[0]), .fa_xor1(u_rca24_fa22_xor1), .fa_or0(u_rca24_fa22_or0));
  fa fa_u_rca24_fa23_out(.a(a[23]), .b(b[23]), .cin(u_rca24_fa22_or0[0]), .fa_xor1(u_rca24_fa23_xor1), .fa_or0(u_rca24_fa23_or0));

  assign u_rca24_out[0] = u_rca24_ha_xor0[0];
  assign u_rca24_out[1] = u_rca24_fa1_xor1[0];
  assign u_rca24_out[2] = u_rca24_fa2_xor1[0];
  assign u_rca24_out[3] = u_rca24_fa3_xor1[0];
  assign u_rca24_out[4] = u_rca24_fa4_xor1[0];
  assign u_rca24_out[5] = u_rca24_fa5_xor1[0];
  assign u_rca24_out[6] = u_rca24_fa6_xor1[0];
  assign u_rca24_out[7] = u_rca24_fa7_xor1[0];
  assign u_rca24_out[8] = u_rca24_fa8_xor1[0];
  assign u_rca24_out[9] = u_rca24_fa9_xor1[0];
  assign u_rca24_out[10] = u_rca24_fa10_xor1[0];
  assign u_rca24_out[11] = u_rca24_fa11_xor1[0];
  assign u_rca24_out[12] = u_rca24_fa12_xor1[0];
  assign u_rca24_out[13] = u_rca24_fa13_xor1[0];
  assign u_rca24_out[14] = u_rca24_fa14_xor1[0];
  assign u_rca24_out[15] = u_rca24_fa15_xor1[0];
  assign u_rca24_out[16] = u_rca24_fa16_xor1[0];
  assign u_rca24_out[17] = u_rca24_fa17_xor1[0];
  assign u_rca24_out[18] = u_rca24_fa18_xor1[0];
  assign u_rca24_out[19] = u_rca24_fa19_xor1[0];
  assign u_rca24_out[20] = u_rca24_fa20_xor1[0];
  assign u_rca24_out[21] = u_rca24_fa21_xor1[0];
  assign u_rca24_out[22] = u_rca24_fa22_xor1[0];
  assign u_rca24_out[23] = u_rca24_fa23_xor1[0];
  assign u_rca24_out[24] = u_rca24_fa23_or0[0];
endmodule

module s_CSAwallace_rca12(input [11:0] a, input [11:0] b, output [23:0] s_CSAwallace_rca12_out);
  wire [0:0] s_CSAwallace_rca12_and_0_0;
  wire [0:0] s_CSAwallace_rca12_and_1_0;
  wire [0:0] s_CSAwallace_rca12_and_2_0;
  wire [0:0] s_CSAwallace_rca12_and_3_0;
  wire [0:0] s_CSAwallace_rca12_and_4_0;
  wire [0:0] s_CSAwallace_rca12_and_5_0;
  wire [0:0] s_CSAwallace_rca12_and_6_0;
  wire [0:0] s_CSAwallace_rca12_and_7_0;
  wire [0:0] s_CSAwallace_rca12_and_8_0;
  wire [0:0] s_CSAwallace_rca12_and_9_0;
  wire [0:0] s_CSAwallace_rca12_and_10_0;
  wire [0:0] s_CSAwallace_rca12_nand_11_0;
  wire [0:0] s_CSAwallace_rca12_and_0_1;
  wire [0:0] s_CSAwallace_rca12_and_1_1;
  wire [0:0] s_CSAwallace_rca12_and_2_1;
  wire [0:0] s_CSAwallace_rca12_and_3_1;
  wire [0:0] s_CSAwallace_rca12_and_4_1;
  wire [0:0] s_CSAwallace_rca12_and_5_1;
  wire [0:0] s_CSAwallace_rca12_and_6_1;
  wire [0:0] s_CSAwallace_rca12_and_7_1;
  wire [0:0] s_CSAwallace_rca12_and_8_1;
  wire [0:0] s_CSAwallace_rca12_and_9_1;
  wire [0:0] s_CSAwallace_rca12_and_10_1;
  wire [0:0] s_CSAwallace_rca12_nand_11_1;
  wire [0:0] s_CSAwallace_rca12_and_0_2;
  wire [0:0] s_CSAwallace_rca12_and_1_2;
  wire [0:0] s_CSAwallace_rca12_and_2_2;
  wire [0:0] s_CSAwallace_rca12_and_3_2;
  wire [0:0] s_CSAwallace_rca12_and_4_2;
  wire [0:0] s_CSAwallace_rca12_and_5_2;
  wire [0:0] s_CSAwallace_rca12_and_6_2;
  wire [0:0] s_CSAwallace_rca12_and_7_2;
  wire [0:0] s_CSAwallace_rca12_and_8_2;
  wire [0:0] s_CSAwallace_rca12_and_9_2;
  wire [0:0] s_CSAwallace_rca12_and_10_2;
  wire [0:0] s_CSAwallace_rca12_nand_11_2;
  wire [0:0] s_CSAwallace_rca12_and_0_3;
  wire [0:0] s_CSAwallace_rca12_and_1_3;
  wire [0:0] s_CSAwallace_rca12_and_2_3;
  wire [0:0] s_CSAwallace_rca12_and_3_3;
  wire [0:0] s_CSAwallace_rca12_and_4_3;
  wire [0:0] s_CSAwallace_rca12_and_5_3;
  wire [0:0] s_CSAwallace_rca12_and_6_3;
  wire [0:0] s_CSAwallace_rca12_and_7_3;
  wire [0:0] s_CSAwallace_rca12_and_8_3;
  wire [0:0] s_CSAwallace_rca12_and_9_3;
  wire [0:0] s_CSAwallace_rca12_and_10_3;
  wire [0:0] s_CSAwallace_rca12_nand_11_3;
  wire [0:0] s_CSAwallace_rca12_and_0_4;
  wire [0:0] s_CSAwallace_rca12_and_1_4;
  wire [0:0] s_CSAwallace_rca12_and_2_4;
  wire [0:0] s_CSAwallace_rca12_and_3_4;
  wire [0:0] s_CSAwallace_rca12_and_4_4;
  wire [0:0] s_CSAwallace_rca12_and_5_4;
  wire [0:0] s_CSAwallace_rca12_and_6_4;
  wire [0:0] s_CSAwallace_rca12_and_7_4;
  wire [0:0] s_CSAwallace_rca12_and_8_4;
  wire [0:0] s_CSAwallace_rca12_and_9_4;
  wire [0:0] s_CSAwallace_rca12_and_10_4;
  wire [0:0] s_CSAwallace_rca12_nand_11_4;
  wire [0:0] s_CSAwallace_rca12_and_0_5;
  wire [0:0] s_CSAwallace_rca12_and_1_5;
  wire [0:0] s_CSAwallace_rca12_and_2_5;
  wire [0:0] s_CSAwallace_rca12_and_3_5;
  wire [0:0] s_CSAwallace_rca12_and_4_5;
  wire [0:0] s_CSAwallace_rca12_and_5_5;
  wire [0:0] s_CSAwallace_rca12_and_6_5;
  wire [0:0] s_CSAwallace_rca12_and_7_5;
  wire [0:0] s_CSAwallace_rca12_and_8_5;
  wire [0:0] s_CSAwallace_rca12_and_9_5;
  wire [0:0] s_CSAwallace_rca12_and_10_5;
  wire [0:0] s_CSAwallace_rca12_nand_11_5;
  wire [0:0] s_CSAwallace_rca12_and_0_6;
  wire [0:0] s_CSAwallace_rca12_and_1_6;
  wire [0:0] s_CSAwallace_rca12_and_2_6;
  wire [0:0] s_CSAwallace_rca12_and_3_6;
  wire [0:0] s_CSAwallace_rca12_and_4_6;
  wire [0:0] s_CSAwallace_rca12_and_5_6;
  wire [0:0] s_CSAwallace_rca12_and_6_6;
  wire [0:0] s_CSAwallace_rca12_and_7_6;
  wire [0:0] s_CSAwallace_rca12_and_8_6;
  wire [0:0] s_CSAwallace_rca12_and_9_6;
  wire [0:0] s_CSAwallace_rca12_and_10_6;
  wire [0:0] s_CSAwallace_rca12_nand_11_6;
  wire [0:0] s_CSAwallace_rca12_and_0_7;
  wire [0:0] s_CSAwallace_rca12_and_1_7;
  wire [0:0] s_CSAwallace_rca12_and_2_7;
  wire [0:0] s_CSAwallace_rca12_and_3_7;
  wire [0:0] s_CSAwallace_rca12_and_4_7;
  wire [0:0] s_CSAwallace_rca12_and_5_7;
  wire [0:0] s_CSAwallace_rca12_and_6_7;
  wire [0:0] s_CSAwallace_rca12_and_7_7;
  wire [0:0] s_CSAwallace_rca12_and_8_7;
  wire [0:0] s_CSAwallace_rca12_and_9_7;
  wire [0:0] s_CSAwallace_rca12_and_10_7;
  wire [0:0] s_CSAwallace_rca12_nand_11_7;
  wire [0:0] s_CSAwallace_rca12_and_0_8;
  wire [0:0] s_CSAwallace_rca12_and_1_8;
  wire [0:0] s_CSAwallace_rca12_and_2_8;
  wire [0:0] s_CSAwallace_rca12_and_3_8;
  wire [0:0] s_CSAwallace_rca12_and_4_8;
  wire [0:0] s_CSAwallace_rca12_and_5_8;
  wire [0:0] s_CSAwallace_rca12_and_6_8;
  wire [0:0] s_CSAwallace_rca12_and_7_8;
  wire [0:0] s_CSAwallace_rca12_and_8_8;
  wire [0:0] s_CSAwallace_rca12_and_9_8;
  wire [0:0] s_CSAwallace_rca12_and_10_8;
  wire [0:0] s_CSAwallace_rca12_nand_11_8;
  wire [0:0] s_CSAwallace_rca12_and_0_9;
  wire [0:0] s_CSAwallace_rca12_and_1_9;
  wire [0:0] s_CSAwallace_rca12_and_2_9;
  wire [0:0] s_CSAwallace_rca12_and_3_9;
  wire [0:0] s_CSAwallace_rca12_and_4_9;
  wire [0:0] s_CSAwallace_rca12_and_5_9;
  wire [0:0] s_CSAwallace_rca12_and_6_9;
  wire [0:0] s_CSAwallace_rca12_and_7_9;
  wire [0:0] s_CSAwallace_rca12_and_8_9;
  wire [0:0] s_CSAwallace_rca12_and_9_9;
  wire [0:0] s_CSAwallace_rca12_and_10_9;
  wire [0:0] s_CSAwallace_rca12_nand_11_9;
  wire [0:0] s_CSAwallace_rca12_and_0_10;
  wire [0:0] s_CSAwallace_rca12_and_1_10;
  wire [0:0] s_CSAwallace_rca12_and_2_10;
  wire [0:0] s_CSAwallace_rca12_and_3_10;
  wire [0:0] s_CSAwallace_rca12_and_4_10;
  wire [0:0] s_CSAwallace_rca12_and_5_10;
  wire [0:0] s_CSAwallace_rca12_and_6_10;
  wire [0:0] s_CSAwallace_rca12_and_7_10;
  wire [0:0] s_CSAwallace_rca12_and_8_10;
  wire [0:0] s_CSAwallace_rca12_and_9_10;
  wire [0:0] s_CSAwallace_rca12_and_10_10;
  wire [0:0] s_CSAwallace_rca12_nand_11_10;
  wire [0:0] s_CSAwallace_rca12_nand_0_11;
  wire [0:0] s_CSAwallace_rca12_nand_1_11;
  wire [0:0] s_CSAwallace_rca12_nand_2_11;
  wire [0:0] s_CSAwallace_rca12_nand_3_11;
  wire [0:0] s_CSAwallace_rca12_nand_4_11;
  wire [0:0] s_CSAwallace_rca12_nand_5_11;
  wire [0:0] s_CSAwallace_rca12_nand_6_11;
  wire [0:0] s_CSAwallace_rca12_nand_7_11;
  wire [0:0] s_CSAwallace_rca12_nand_8_11;
  wire [0:0] s_CSAwallace_rca12_nand_9_11;
  wire [0:0] s_CSAwallace_rca12_nand_10_11;
  wire [0:0] s_CSAwallace_rca12_and_11_11;
  wire [13:0] s_CSAwallace_rca12_csa0_csa_component_pp_row0;
  wire [13:0] s_CSAwallace_rca12_csa0_csa_component_pp_row1;
  wire [13:0] s_CSAwallace_rca12_csa0_csa_component_pp_row2;
  wire [29:0] s_CSAwallace_rca12_csa0_csa_component_out;
  wire [16:0] s_CSAwallace_rca12_csa1_csa_component_pp_row3;
  wire [16:0] s_CSAwallace_rca12_csa1_csa_component_pp_row4;
  wire [16:0] s_CSAwallace_rca12_csa1_csa_component_pp_row5;
  wire [35:0] s_CSAwallace_rca12_csa1_csa_component_out;
  wire [19:0] s_CSAwallace_rca12_csa2_csa_component_pp_row6;
  wire [19:0] s_CSAwallace_rca12_csa2_csa_component_pp_row7;
  wire [19:0] s_CSAwallace_rca12_csa2_csa_component_pp_row8;
  wire [41:0] s_CSAwallace_rca12_csa2_csa_component_out;
  wire [22:0] s_CSAwallace_rca12_csa3_csa_component_pp_row9;
  wire [22:0] s_CSAwallace_rca12_csa3_csa_component_pp_row10;
  wire [22:0] s_CSAwallace_rca12_csa3_csa_component_pp_row11;
  wire [47:0] s_CSAwallace_rca12_csa3_csa_component_out;
  wire [17:0] s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1;
  wire [17:0] s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1;
  wire [17:0] s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2;
  wire [37:0] s_CSAwallace_rca12_csa4_csa_component_out;
  wire [20:0] s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2;
  wire [20:0] s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3;
  wire [20:0] s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3;
  wire [43:0] s_CSAwallace_rca12_csa5_csa_component_out;
  wire [21:0] s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5;
  wire [21:0] s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5;
  wire [21:0] s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6;
  wire [45:0] s_CSAwallace_rca12_csa6_csa_component_out;
  wire [23:0] s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6;
  wire [23:0] s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4;
  wire [23:0] s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4;
  wire [49:0] s_CSAwallace_rca12_csa7_csa_component_out;
  wire [23:0] s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7;
  wire [23:0] s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7;
  wire [23:0] s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8;
  wire [49:0] s_CSAwallace_rca12_csa8_csa_component_out;
  wire [23:0] s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9;
  wire [23:0] s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9;
  wire [23:0] s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8;
  wire [49:0] s_CSAwallace_rca12_csa9_csa_component_out;
  wire [23:0] s_CSAwallace_rca12_u_rca24_a;
  wire [23:0] s_CSAwallace_rca12_u_rca24_b;
  wire [24:0] s_CSAwallace_rca12_u_rca24_out;
  wire [0:0] s_CSAwallace_rca12_xor0;

  and_gate and_gate_s_CSAwallace_rca12_and_0_0(.a(a[0]), .b(b[0]), .out(s_CSAwallace_rca12_and_0_0));
  and_gate and_gate_s_CSAwallace_rca12_and_1_0(.a(a[1]), .b(b[0]), .out(s_CSAwallace_rca12_and_1_0));
  and_gate and_gate_s_CSAwallace_rca12_and_2_0(.a(a[2]), .b(b[0]), .out(s_CSAwallace_rca12_and_2_0));
  and_gate and_gate_s_CSAwallace_rca12_and_3_0(.a(a[3]), .b(b[0]), .out(s_CSAwallace_rca12_and_3_0));
  and_gate and_gate_s_CSAwallace_rca12_and_4_0(.a(a[4]), .b(b[0]), .out(s_CSAwallace_rca12_and_4_0));
  and_gate and_gate_s_CSAwallace_rca12_and_5_0(.a(a[5]), .b(b[0]), .out(s_CSAwallace_rca12_and_5_0));
  and_gate and_gate_s_CSAwallace_rca12_and_6_0(.a(a[6]), .b(b[0]), .out(s_CSAwallace_rca12_and_6_0));
  and_gate and_gate_s_CSAwallace_rca12_and_7_0(.a(a[7]), .b(b[0]), .out(s_CSAwallace_rca12_and_7_0));
  and_gate and_gate_s_CSAwallace_rca12_and_8_0(.a(a[8]), .b(b[0]), .out(s_CSAwallace_rca12_and_8_0));
  and_gate and_gate_s_CSAwallace_rca12_and_9_0(.a(a[9]), .b(b[0]), .out(s_CSAwallace_rca12_and_9_0));
  and_gate and_gate_s_CSAwallace_rca12_and_10_0(.a(a[10]), .b(b[0]), .out(s_CSAwallace_rca12_and_10_0));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_0(.a(a[11]), .b(b[0]), .out(s_CSAwallace_rca12_nand_11_0));
  and_gate and_gate_s_CSAwallace_rca12_and_0_1(.a(a[0]), .b(b[1]), .out(s_CSAwallace_rca12_and_0_1));
  and_gate and_gate_s_CSAwallace_rca12_and_1_1(.a(a[1]), .b(b[1]), .out(s_CSAwallace_rca12_and_1_1));
  and_gate and_gate_s_CSAwallace_rca12_and_2_1(.a(a[2]), .b(b[1]), .out(s_CSAwallace_rca12_and_2_1));
  and_gate and_gate_s_CSAwallace_rca12_and_3_1(.a(a[3]), .b(b[1]), .out(s_CSAwallace_rca12_and_3_1));
  and_gate and_gate_s_CSAwallace_rca12_and_4_1(.a(a[4]), .b(b[1]), .out(s_CSAwallace_rca12_and_4_1));
  and_gate and_gate_s_CSAwallace_rca12_and_5_1(.a(a[5]), .b(b[1]), .out(s_CSAwallace_rca12_and_5_1));
  and_gate and_gate_s_CSAwallace_rca12_and_6_1(.a(a[6]), .b(b[1]), .out(s_CSAwallace_rca12_and_6_1));
  and_gate and_gate_s_CSAwallace_rca12_and_7_1(.a(a[7]), .b(b[1]), .out(s_CSAwallace_rca12_and_7_1));
  and_gate and_gate_s_CSAwallace_rca12_and_8_1(.a(a[8]), .b(b[1]), .out(s_CSAwallace_rca12_and_8_1));
  and_gate and_gate_s_CSAwallace_rca12_and_9_1(.a(a[9]), .b(b[1]), .out(s_CSAwallace_rca12_and_9_1));
  and_gate and_gate_s_CSAwallace_rca12_and_10_1(.a(a[10]), .b(b[1]), .out(s_CSAwallace_rca12_and_10_1));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_1(.a(a[11]), .b(b[1]), .out(s_CSAwallace_rca12_nand_11_1));
  and_gate and_gate_s_CSAwallace_rca12_and_0_2(.a(a[0]), .b(b[2]), .out(s_CSAwallace_rca12_and_0_2));
  and_gate and_gate_s_CSAwallace_rca12_and_1_2(.a(a[1]), .b(b[2]), .out(s_CSAwallace_rca12_and_1_2));
  and_gate and_gate_s_CSAwallace_rca12_and_2_2(.a(a[2]), .b(b[2]), .out(s_CSAwallace_rca12_and_2_2));
  and_gate and_gate_s_CSAwallace_rca12_and_3_2(.a(a[3]), .b(b[2]), .out(s_CSAwallace_rca12_and_3_2));
  and_gate and_gate_s_CSAwallace_rca12_and_4_2(.a(a[4]), .b(b[2]), .out(s_CSAwallace_rca12_and_4_2));
  and_gate and_gate_s_CSAwallace_rca12_and_5_2(.a(a[5]), .b(b[2]), .out(s_CSAwallace_rca12_and_5_2));
  and_gate and_gate_s_CSAwallace_rca12_and_6_2(.a(a[6]), .b(b[2]), .out(s_CSAwallace_rca12_and_6_2));
  and_gate and_gate_s_CSAwallace_rca12_and_7_2(.a(a[7]), .b(b[2]), .out(s_CSAwallace_rca12_and_7_2));
  and_gate and_gate_s_CSAwallace_rca12_and_8_2(.a(a[8]), .b(b[2]), .out(s_CSAwallace_rca12_and_8_2));
  and_gate and_gate_s_CSAwallace_rca12_and_9_2(.a(a[9]), .b(b[2]), .out(s_CSAwallace_rca12_and_9_2));
  and_gate and_gate_s_CSAwallace_rca12_and_10_2(.a(a[10]), .b(b[2]), .out(s_CSAwallace_rca12_and_10_2));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_2(.a(a[11]), .b(b[2]), .out(s_CSAwallace_rca12_nand_11_2));
  and_gate and_gate_s_CSAwallace_rca12_and_0_3(.a(a[0]), .b(b[3]), .out(s_CSAwallace_rca12_and_0_3));
  and_gate and_gate_s_CSAwallace_rca12_and_1_3(.a(a[1]), .b(b[3]), .out(s_CSAwallace_rca12_and_1_3));
  and_gate and_gate_s_CSAwallace_rca12_and_2_3(.a(a[2]), .b(b[3]), .out(s_CSAwallace_rca12_and_2_3));
  and_gate and_gate_s_CSAwallace_rca12_and_3_3(.a(a[3]), .b(b[3]), .out(s_CSAwallace_rca12_and_3_3));
  and_gate and_gate_s_CSAwallace_rca12_and_4_3(.a(a[4]), .b(b[3]), .out(s_CSAwallace_rca12_and_4_3));
  and_gate and_gate_s_CSAwallace_rca12_and_5_3(.a(a[5]), .b(b[3]), .out(s_CSAwallace_rca12_and_5_3));
  and_gate and_gate_s_CSAwallace_rca12_and_6_3(.a(a[6]), .b(b[3]), .out(s_CSAwallace_rca12_and_6_3));
  and_gate and_gate_s_CSAwallace_rca12_and_7_3(.a(a[7]), .b(b[3]), .out(s_CSAwallace_rca12_and_7_3));
  and_gate and_gate_s_CSAwallace_rca12_and_8_3(.a(a[8]), .b(b[3]), .out(s_CSAwallace_rca12_and_8_3));
  and_gate and_gate_s_CSAwallace_rca12_and_9_3(.a(a[9]), .b(b[3]), .out(s_CSAwallace_rca12_and_9_3));
  and_gate and_gate_s_CSAwallace_rca12_and_10_3(.a(a[10]), .b(b[3]), .out(s_CSAwallace_rca12_and_10_3));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_3(.a(a[11]), .b(b[3]), .out(s_CSAwallace_rca12_nand_11_3));
  and_gate and_gate_s_CSAwallace_rca12_and_0_4(.a(a[0]), .b(b[4]), .out(s_CSAwallace_rca12_and_0_4));
  and_gate and_gate_s_CSAwallace_rca12_and_1_4(.a(a[1]), .b(b[4]), .out(s_CSAwallace_rca12_and_1_4));
  and_gate and_gate_s_CSAwallace_rca12_and_2_4(.a(a[2]), .b(b[4]), .out(s_CSAwallace_rca12_and_2_4));
  and_gate and_gate_s_CSAwallace_rca12_and_3_4(.a(a[3]), .b(b[4]), .out(s_CSAwallace_rca12_and_3_4));
  and_gate and_gate_s_CSAwallace_rca12_and_4_4(.a(a[4]), .b(b[4]), .out(s_CSAwallace_rca12_and_4_4));
  and_gate and_gate_s_CSAwallace_rca12_and_5_4(.a(a[5]), .b(b[4]), .out(s_CSAwallace_rca12_and_5_4));
  and_gate and_gate_s_CSAwallace_rca12_and_6_4(.a(a[6]), .b(b[4]), .out(s_CSAwallace_rca12_and_6_4));
  and_gate and_gate_s_CSAwallace_rca12_and_7_4(.a(a[7]), .b(b[4]), .out(s_CSAwallace_rca12_and_7_4));
  and_gate and_gate_s_CSAwallace_rca12_and_8_4(.a(a[8]), .b(b[4]), .out(s_CSAwallace_rca12_and_8_4));
  and_gate and_gate_s_CSAwallace_rca12_and_9_4(.a(a[9]), .b(b[4]), .out(s_CSAwallace_rca12_and_9_4));
  and_gate and_gate_s_CSAwallace_rca12_and_10_4(.a(a[10]), .b(b[4]), .out(s_CSAwallace_rca12_and_10_4));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_4(.a(a[11]), .b(b[4]), .out(s_CSAwallace_rca12_nand_11_4));
  and_gate and_gate_s_CSAwallace_rca12_and_0_5(.a(a[0]), .b(b[5]), .out(s_CSAwallace_rca12_and_0_5));
  and_gate and_gate_s_CSAwallace_rca12_and_1_5(.a(a[1]), .b(b[5]), .out(s_CSAwallace_rca12_and_1_5));
  and_gate and_gate_s_CSAwallace_rca12_and_2_5(.a(a[2]), .b(b[5]), .out(s_CSAwallace_rca12_and_2_5));
  and_gate and_gate_s_CSAwallace_rca12_and_3_5(.a(a[3]), .b(b[5]), .out(s_CSAwallace_rca12_and_3_5));
  and_gate and_gate_s_CSAwallace_rca12_and_4_5(.a(a[4]), .b(b[5]), .out(s_CSAwallace_rca12_and_4_5));
  and_gate and_gate_s_CSAwallace_rca12_and_5_5(.a(a[5]), .b(b[5]), .out(s_CSAwallace_rca12_and_5_5));
  and_gate and_gate_s_CSAwallace_rca12_and_6_5(.a(a[6]), .b(b[5]), .out(s_CSAwallace_rca12_and_6_5));
  and_gate and_gate_s_CSAwallace_rca12_and_7_5(.a(a[7]), .b(b[5]), .out(s_CSAwallace_rca12_and_7_5));
  and_gate and_gate_s_CSAwallace_rca12_and_8_5(.a(a[8]), .b(b[5]), .out(s_CSAwallace_rca12_and_8_5));
  and_gate and_gate_s_CSAwallace_rca12_and_9_5(.a(a[9]), .b(b[5]), .out(s_CSAwallace_rca12_and_9_5));
  and_gate and_gate_s_CSAwallace_rca12_and_10_5(.a(a[10]), .b(b[5]), .out(s_CSAwallace_rca12_and_10_5));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_5(.a(a[11]), .b(b[5]), .out(s_CSAwallace_rca12_nand_11_5));
  and_gate and_gate_s_CSAwallace_rca12_and_0_6(.a(a[0]), .b(b[6]), .out(s_CSAwallace_rca12_and_0_6));
  and_gate and_gate_s_CSAwallace_rca12_and_1_6(.a(a[1]), .b(b[6]), .out(s_CSAwallace_rca12_and_1_6));
  and_gate and_gate_s_CSAwallace_rca12_and_2_6(.a(a[2]), .b(b[6]), .out(s_CSAwallace_rca12_and_2_6));
  and_gate and_gate_s_CSAwallace_rca12_and_3_6(.a(a[3]), .b(b[6]), .out(s_CSAwallace_rca12_and_3_6));
  and_gate and_gate_s_CSAwallace_rca12_and_4_6(.a(a[4]), .b(b[6]), .out(s_CSAwallace_rca12_and_4_6));
  and_gate and_gate_s_CSAwallace_rca12_and_5_6(.a(a[5]), .b(b[6]), .out(s_CSAwallace_rca12_and_5_6));
  and_gate and_gate_s_CSAwallace_rca12_and_6_6(.a(a[6]), .b(b[6]), .out(s_CSAwallace_rca12_and_6_6));
  and_gate and_gate_s_CSAwallace_rca12_and_7_6(.a(a[7]), .b(b[6]), .out(s_CSAwallace_rca12_and_7_6));
  and_gate and_gate_s_CSAwallace_rca12_and_8_6(.a(a[8]), .b(b[6]), .out(s_CSAwallace_rca12_and_8_6));
  and_gate and_gate_s_CSAwallace_rca12_and_9_6(.a(a[9]), .b(b[6]), .out(s_CSAwallace_rca12_and_9_6));
  and_gate and_gate_s_CSAwallace_rca12_and_10_6(.a(a[10]), .b(b[6]), .out(s_CSAwallace_rca12_and_10_6));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_6(.a(a[11]), .b(b[6]), .out(s_CSAwallace_rca12_nand_11_6));
  and_gate and_gate_s_CSAwallace_rca12_and_0_7(.a(a[0]), .b(b[7]), .out(s_CSAwallace_rca12_and_0_7));
  and_gate and_gate_s_CSAwallace_rca12_and_1_7(.a(a[1]), .b(b[7]), .out(s_CSAwallace_rca12_and_1_7));
  and_gate and_gate_s_CSAwallace_rca12_and_2_7(.a(a[2]), .b(b[7]), .out(s_CSAwallace_rca12_and_2_7));
  and_gate and_gate_s_CSAwallace_rca12_and_3_7(.a(a[3]), .b(b[7]), .out(s_CSAwallace_rca12_and_3_7));
  and_gate and_gate_s_CSAwallace_rca12_and_4_7(.a(a[4]), .b(b[7]), .out(s_CSAwallace_rca12_and_4_7));
  and_gate and_gate_s_CSAwallace_rca12_and_5_7(.a(a[5]), .b(b[7]), .out(s_CSAwallace_rca12_and_5_7));
  and_gate and_gate_s_CSAwallace_rca12_and_6_7(.a(a[6]), .b(b[7]), .out(s_CSAwallace_rca12_and_6_7));
  and_gate and_gate_s_CSAwallace_rca12_and_7_7(.a(a[7]), .b(b[7]), .out(s_CSAwallace_rca12_and_7_7));
  and_gate and_gate_s_CSAwallace_rca12_and_8_7(.a(a[8]), .b(b[7]), .out(s_CSAwallace_rca12_and_8_7));
  and_gate and_gate_s_CSAwallace_rca12_and_9_7(.a(a[9]), .b(b[7]), .out(s_CSAwallace_rca12_and_9_7));
  and_gate and_gate_s_CSAwallace_rca12_and_10_7(.a(a[10]), .b(b[7]), .out(s_CSAwallace_rca12_and_10_7));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_7(.a(a[11]), .b(b[7]), .out(s_CSAwallace_rca12_nand_11_7));
  and_gate and_gate_s_CSAwallace_rca12_and_0_8(.a(a[0]), .b(b[8]), .out(s_CSAwallace_rca12_and_0_8));
  and_gate and_gate_s_CSAwallace_rca12_and_1_8(.a(a[1]), .b(b[8]), .out(s_CSAwallace_rca12_and_1_8));
  and_gate and_gate_s_CSAwallace_rca12_and_2_8(.a(a[2]), .b(b[8]), .out(s_CSAwallace_rca12_and_2_8));
  and_gate and_gate_s_CSAwallace_rca12_and_3_8(.a(a[3]), .b(b[8]), .out(s_CSAwallace_rca12_and_3_8));
  and_gate and_gate_s_CSAwallace_rca12_and_4_8(.a(a[4]), .b(b[8]), .out(s_CSAwallace_rca12_and_4_8));
  and_gate and_gate_s_CSAwallace_rca12_and_5_8(.a(a[5]), .b(b[8]), .out(s_CSAwallace_rca12_and_5_8));
  and_gate and_gate_s_CSAwallace_rca12_and_6_8(.a(a[6]), .b(b[8]), .out(s_CSAwallace_rca12_and_6_8));
  and_gate and_gate_s_CSAwallace_rca12_and_7_8(.a(a[7]), .b(b[8]), .out(s_CSAwallace_rca12_and_7_8));
  and_gate and_gate_s_CSAwallace_rca12_and_8_8(.a(a[8]), .b(b[8]), .out(s_CSAwallace_rca12_and_8_8));
  and_gate and_gate_s_CSAwallace_rca12_and_9_8(.a(a[9]), .b(b[8]), .out(s_CSAwallace_rca12_and_9_8));
  and_gate and_gate_s_CSAwallace_rca12_and_10_8(.a(a[10]), .b(b[8]), .out(s_CSAwallace_rca12_and_10_8));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_8(.a(a[11]), .b(b[8]), .out(s_CSAwallace_rca12_nand_11_8));
  and_gate and_gate_s_CSAwallace_rca12_and_0_9(.a(a[0]), .b(b[9]), .out(s_CSAwallace_rca12_and_0_9));
  and_gate and_gate_s_CSAwallace_rca12_and_1_9(.a(a[1]), .b(b[9]), .out(s_CSAwallace_rca12_and_1_9));
  and_gate and_gate_s_CSAwallace_rca12_and_2_9(.a(a[2]), .b(b[9]), .out(s_CSAwallace_rca12_and_2_9));
  and_gate and_gate_s_CSAwallace_rca12_and_3_9(.a(a[3]), .b(b[9]), .out(s_CSAwallace_rca12_and_3_9));
  and_gate and_gate_s_CSAwallace_rca12_and_4_9(.a(a[4]), .b(b[9]), .out(s_CSAwallace_rca12_and_4_9));
  and_gate and_gate_s_CSAwallace_rca12_and_5_9(.a(a[5]), .b(b[9]), .out(s_CSAwallace_rca12_and_5_9));
  and_gate and_gate_s_CSAwallace_rca12_and_6_9(.a(a[6]), .b(b[9]), .out(s_CSAwallace_rca12_and_6_9));
  and_gate and_gate_s_CSAwallace_rca12_and_7_9(.a(a[7]), .b(b[9]), .out(s_CSAwallace_rca12_and_7_9));
  and_gate and_gate_s_CSAwallace_rca12_and_8_9(.a(a[8]), .b(b[9]), .out(s_CSAwallace_rca12_and_8_9));
  and_gate and_gate_s_CSAwallace_rca12_and_9_9(.a(a[9]), .b(b[9]), .out(s_CSAwallace_rca12_and_9_9));
  and_gate and_gate_s_CSAwallace_rca12_and_10_9(.a(a[10]), .b(b[9]), .out(s_CSAwallace_rca12_and_10_9));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_9(.a(a[11]), .b(b[9]), .out(s_CSAwallace_rca12_nand_11_9));
  and_gate and_gate_s_CSAwallace_rca12_and_0_10(.a(a[0]), .b(b[10]), .out(s_CSAwallace_rca12_and_0_10));
  and_gate and_gate_s_CSAwallace_rca12_and_1_10(.a(a[1]), .b(b[10]), .out(s_CSAwallace_rca12_and_1_10));
  and_gate and_gate_s_CSAwallace_rca12_and_2_10(.a(a[2]), .b(b[10]), .out(s_CSAwallace_rca12_and_2_10));
  and_gate and_gate_s_CSAwallace_rca12_and_3_10(.a(a[3]), .b(b[10]), .out(s_CSAwallace_rca12_and_3_10));
  and_gate and_gate_s_CSAwallace_rca12_and_4_10(.a(a[4]), .b(b[10]), .out(s_CSAwallace_rca12_and_4_10));
  and_gate and_gate_s_CSAwallace_rca12_and_5_10(.a(a[5]), .b(b[10]), .out(s_CSAwallace_rca12_and_5_10));
  and_gate and_gate_s_CSAwallace_rca12_and_6_10(.a(a[6]), .b(b[10]), .out(s_CSAwallace_rca12_and_6_10));
  and_gate and_gate_s_CSAwallace_rca12_and_7_10(.a(a[7]), .b(b[10]), .out(s_CSAwallace_rca12_and_7_10));
  and_gate and_gate_s_CSAwallace_rca12_and_8_10(.a(a[8]), .b(b[10]), .out(s_CSAwallace_rca12_and_8_10));
  and_gate and_gate_s_CSAwallace_rca12_and_9_10(.a(a[9]), .b(b[10]), .out(s_CSAwallace_rca12_and_9_10));
  and_gate and_gate_s_CSAwallace_rca12_and_10_10(.a(a[10]), .b(b[10]), .out(s_CSAwallace_rca12_and_10_10));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_11_10(.a(a[11]), .b(b[10]), .out(s_CSAwallace_rca12_nand_11_10));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_0_11(.a(a[0]), .b(b[11]), .out(s_CSAwallace_rca12_nand_0_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_1_11(.a(a[1]), .b(b[11]), .out(s_CSAwallace_rca12_nand_1_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_2_11(.a(a[2]), .b(b[11]), .out(s_CSAwallace_rca12_nand_2_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_3_11(.a(a[3]), .b(b[11]), .out(s_CSAwallace_rca12_nand_3_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_4_11(.a(a[4]), .b(b[11]), .out(s_CSAwallace_rca12_nand_4_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_5_11(.a(a[5]), .b(b[11]), .out(s_CSAwallace_rca12_nand_5_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_6_11(.a(a[6]), .b(b[11]), .out(s_CSAwallace_rca12_nand_6_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_7_11(.a(a[7]), .b(b[11]), .out(s_CSAwallace_rca12_nand_7_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_8_11(.a(a[8]), .b(b[11]), .out(s_CSAwallace_rca12_nand_8_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_9_11(.a(a[9]), .b(b[11]), .out(s_CSAwallace_rca12_nand_9_11));
  nand_gate nand_gate_s_CSAwallace_rca12_nand_10_11(.a(a[10]), .b(b[11]), .out(s_CSAwallace_rca12_nand_10_11));
  and_gate and_gate_s_CSAwallace_rca12_and_11_11(.a(a[11]), .b(b[11]), .out(s_CSAwallace_rca12_and_11_11));
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[0] = s_CSAwallace_rca12_and_0_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[1] = s_CSAwallace_rca12_and_1_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[2] = s_CSAwallace_rca12_and_2_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[3] = s_CSAwallace_rca12_and_3_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[4] = s_CSAwallace_rca12_and_4_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[5] = s_CSAwallace_rca12_and_5_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[6] = s_CSAwallace_rca12_and_6_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[7] = s_CSAwallace_rca12_and_7_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[8] = s_CSAwallace_rca12_and_8_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[9] = s_CSAwallace_rca12_and_9_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[10] = s_CSAwallace_rca12_and_10_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[11] = s_CSAwallace_rca12_nand_11_0[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[12] = 1'b1;
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row0[13] = 1'b1;
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[0] = 1'b0;
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[1] = s_CSAwallace_rca12_and_0_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[2] = s_CSAwallace_rca12_and_1_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[3] = s_CSAwallace_rca12_and_2_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[4] = s_CSAwallace_rca12_and_3_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[5] = s_CSAwallace_rca12_and_4_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[6] = s_CSAwallace_rca12_and_5_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[7] = s_CSAwallace_rca12_and_6_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[8] = s_CSAwallace_rca12_and_7_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[9] = s_CSAwallace_rca12_and_8_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[10] = s_CSAwallace_rca12_and_9_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[11] = s_CSAwallace_rca12_and_10_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[12] = s_CSAwallace_rca12_nand_11_1[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row1[13] = 1'b1;
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[0] = 1'b0;
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[1] = 1'b0;
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[2] = s_CSAwallace_rca12_and_0_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[3] = s_CSAwallace_rca12_and_1_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[4] = s_CSAwallace_rca12_and_2_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[5] = s_CSAwallace_rca12_and_3_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[6] = s_CSAwallace_rca12_and_4_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[7] = s_CSAwallace_rca12_and_5_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[8] = s_CSAwallace_rca12_and_6_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[9] = s_CSAwallace_rca12_and_7_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[10] = s_CSAwallace_rca12_and_8_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[11] = s_CSAwallace_rca12_and_9_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[12] = s_CSAwallace_rca12_and_10_2[0];
  assign s_CSAwallace_rca12_csa0_csa_component_pp_row2[13] = s_CSAwallace_rca12_nand_11_2[0];
  csa_component14 csa_component14_s_CSAwallace_rca12_csa0_csa_component_out(.a(s_CSAwallace_rca12_csa0_csa_component_pp_row0), .b(s_CSAwallace_rca12_csa0_csa_component_pp_row1), .c(s_CSAwallace_rca12_csa0_csa_component_pp_row2), .csa_component14_out(s_CSAwallace_rca12_csa0_csa_component_out));
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[0] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[1] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[2] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[3] = s_CSAwallace_rca12_and_0_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[4] = s_CSAwallace_rca12_and_1_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[5] = s_CSAwallace_rca12_and_2_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[6] = s_CSAwallace_rca12_and_3_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[7] = s_CSAwallace_rca12_and_4_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[8] = s_CSAwallace_rca12_and_5_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[9] = s_CSAwallace_rca12_and_6_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[10] = s_CSAwallace_rca12_and_7_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[11] = s_CSAwallace_rca12_and_8_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[12] = s_CSAwallace_rca12_and_9_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[13] = s_CSAwallace_rca12_and_10_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[14] = s_CSAwallace_rca12_nand_11_3[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[15] = 1'b1;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row3[16] = 1'b1;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[0] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[1] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[2] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[3] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[4] = s_CSAwallace_rca12_and_0_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[5] = s_CSAwallace_rca12_and_1_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[6] = s_CSAwallace_rca12_and_2_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[7] = s_CSAwallace_rca12_and_3_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[8] = s_CSAwallace_rca12_and_4_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[9] = s_CSAwallace_rca12_and_5_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[10] = s_CSAwallace_rca12_and_6_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[11] = s_CSAwallace_rca12_and_7_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[12] = s_CSAwallace_rca12_and_8_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[13] = s_CSAwallace_rca12_and_9_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[14] = s_CSAwallace_rca12_and_10_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[15] = s_CSAwallace_rca12_nand_11_4[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row4[16] = 1'b1;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[0] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[1] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[2] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[3] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[4] = 1'b0;
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[5] = s_CSAwallace_rca12_and_0_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[6] = s_CSAwallace_rca12_and_1_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[7] = s_CSAwallace_rca12_and_2_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[8] = s_CSAwallace_rca12_and_3_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[9] = s_CSAwallace_rca12_and_4_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[10] = s_CSAwallace_rca12_and_5_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[11] = s_CSAwallace_rca12_and_6_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[12] = s_CSAwallace_rca12_and_7_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[13] = s_CSAwallace_rca12_and_8_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[14] = s_CSAwallace_rca12_and_9_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[15] = s_CSAwallace_rca12_and_10_5[0];
  assign s_CSAwallace_rca12_csa1_csa_component_pp_row5[16] = s_CSAwallace_rca12_nand_11_5[0];
  csa_component17 csa_component17_s_CSAwallace_rca12_csa1_csa_component_out(.a(s_CSAwallace_rca12_csa1_csa_component_pp_row3), .b(s_CSAwallace_rca12_csa1_csa_component_pp_row4), .c(s_CSAwallace_rca12_csa1_csa_component_pp_row5), .csa_component17_out(s_CSAwallace_rca12_csa1_csa_component_out));
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[0] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[1] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[2] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[3] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[4] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[5] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[6] = s_CSAwallace_rca12_and_0_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[7] = s_CSAwallace_rca12_and_1_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[8] = s_CSAwallace_rca12_and_2_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[9] = s_CSAwallace_rca12_and_3_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[10] = s_CSAwallace_rca12_and_4_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[11] = s_CSAwallace_rca12_and_5_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[12] = s_CSAwallace_rca12_and_6_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[13] = s_CSAwallace_rca12_and_7_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[14] = s_CSAwallace_rca12_and_8_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[15] = s_CSAwallace_rca12_and_9_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[16] = s_CSAwallace_rca12_and_10_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[17] = s_CSAwallace_rca12_nand_11_6[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[18] = 1'b1;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row6[19] = 1'b1;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[0] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[1] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[2] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[3] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[4] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[5] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[6] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[7] = s_CSAwallace_rca12_and_0_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[8] = s_CSAwallace_rca12_and_1_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[9] = s_CSAwallace_rca12_and_2_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[10] = s_CSAwallace_rca12_and_3_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[11] = s_CSAwallace_rca12_and_4_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[12] = s_CSAwallace_rca12_and_5_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[13] = s_CSAwallace_rca12_and_6_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[14] = s_CSAwallace_rca12_and_7_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[15] = s_CSAwallace_rca12_and_8_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[16] = s_CSAwallace_rca12_and_9_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[17] = s_CSAwallace_rca12_and_10_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[18] = s_CSAwallace_rca12_nand_11_7[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row7[19] = 1'b1;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[0] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[1] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[2] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[3] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[4] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[5] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[6] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[7] = 1'b0;
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[8] = s_CSAwallace_rca12_and_0_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[9] = s_CSAwallace_rca12_and_1_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[10] = s_CSAwallace_rca12_and_2_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[11] = s_CSAwallace_rca12_and_3_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[12] = s_CSAwallace_rca12_and_4_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[13] = s_CSAwallace_rca12_and_5_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[14] = s_CSAwallace_rca12_and_6_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[15] = s_CSAwallace_rca12_and_7_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[16] = s_CSAwallace_rca12_and_8_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[17] = s_CSAwallace_rca12_and_9_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[18] = s_CSAwallace_rca12_and_10_8[0];
  assign s_CSAwallace_rca12_csa2_csa_component_pp_row8[19] = s_CSAwallace_rca12_nand_11_8[0];
  csa_component20 csa_component20_s_CSAwallace_rca12_csa2_csa_component_out(.a(s_CSAwallace_rca12_csa2_csa_component_pp_row6), .b(s_CSAwallace_rca12_csa2_csa_component_pp_row7), .c(s_CSAwallace_rca12_csa2_csa_component_pp_row8), .csa_component20_out(s_CSAwallace_rca12_csa2_csa_component_out));
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[0] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[1] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[2] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[3] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[4] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[5] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[6] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[7] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[8] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[9] = s_CSAwallace_rca12_and_0_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[10] = s_CSAwallace_rca12_and_1_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[11] = s_CSAwallace_rca12_and_2_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[12] = s_CSAwallace_rca12_and_3_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[13] = s_CSAwallace_rca12_and_4_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[14] = s_CSAwallace_rca12_and_5_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[15] = s_CSAwallace_rca12_and_6_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[16] = s_CSAwallace_rca12_and_7_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[17] = s_CSAwallace_rca12_and_8_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[18] = s_CSAwallace_rca12_and_9_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[19] = s_CSAwallace_rca12_and_10_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[20] = s_CSAwallace_rca12_nand_11_9[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[21] = 1'b1;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row9[22] = 1'b1;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[0] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[1] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[2] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[3] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[4] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[5] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[6] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[7] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[8] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[9] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[10] = s_CSAwallace_rca12_and_0_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[11] = s_CSAwallace_rca12_and_1_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[12] = s_CSAwallace_rca12_and_2_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[13] = s_CSAwallace_rca12_and_3_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[14] = s_CSAwallace_rca12_and_4_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[15] = s_CSAwallace_rca12_and_5_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[16] = s_CSAwallace_rca12_and_6_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[17] = s_CSAwallace_rca12_and_7_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[18] = s_CSAwallace_rca12_and_8_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[19] = s_CSAwallace_rca12_and_9_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[20] = s_CSAwallace_rca12_and_10_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[21] = s_CSAwallace_rca12_nand_11_10[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row10[22] = 1'b1;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[0] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[1] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[2] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[3] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[4] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[5] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[6] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[7] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[8] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[9] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[10] = 1'b0;
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[11] = s_CSAwallace_rca12_nand_0_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[12] = s_CSAwallace_rca12_nand_1_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[13] = s_CSAwallace_rca12_nand_2_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[14] = s_CSAwallace_rca12_nand_3_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[15] = s_CSAwallace_rca12_nand_4_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[16] = s_CSAwallace_rca12_nand_5_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[17] = s_CSAwallace_rca12_nand_6_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[18] = s_CSAwallace_rca12_nand_7_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[19] = s_CSAwallace_rca12_nand_8_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[20] = s_CSAwallace_rca12_nand_9_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[21] = s_CSAwallace_rca12_nand_10_11[0];
  assign s_CSAwallace_rca12_csa3_csa_component_pp_row11[22] = s_CSAwallace_rca12_and_11_11[0];
  csa_component23 csa_component23_s_CSAwallace_rca12_csa3_csa_component_out(.a(s_CSAwallace_rca12_csa3_csa_component_pp_row9), .b(s_CSAwallace_rca12_csa3_csa_component_pp_row10), .c(s_CSAwallace_rca12_csa3_csa_component_pp_row11), .csa_component23_out(s_CSAwallace_rca12_csa3_csa_component_out));
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[0] = s_CSAwallace_rca12_csa0_csa_component_out[0];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[1] = s_CSAwallace_rca12_csa0_csa_component_out[1];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[2] = s_CSAwallace_rca12_csa0_csa_component_out[2];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[3] = s_CSAwallace_rca12_csa0_csa_component_out[3];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[4] = s_CSAwallace_rca12_csa0_csa_component_out[4];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[5] = s_CSAwallace_rca12_csa0_csa_component_out[5];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[6] = s_CSAwallace_rca12_csa0_csa_component_out[6];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[7] = s_CSAwallace_rca12_csa0_csa_component_out[7];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[8] = s_CSAwallace_rca12_csa0_csa_component_out[8];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[9] = s_CSAwallace_rca12_csa0_csa_component_out[9];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[10] = s_CSAwallace_rca12_csa0_csa_component_out[10];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[11] = s_CSAwallace_rca12_csa0_csa_component_out[11];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[12] = s_CSAwallace_rca12_csa0_csa_component_out[12];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[13] = s_CSAwallace_rca12_csa0_csa_component_out[13];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[14] = 1'b1;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[15] = 1'b1;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[16] = 1'b1;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1[17] = 1'b1;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[0] = 1'b0;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[1] = 1'b0;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[2] = s_CSAwallace_rca12_csa0_csa_component_out[17];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[3] = s_CSAwallace_rca12_csa0_csa_component_out[18];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[4] = s_CSAwallace_rca12_csa0_csa_component_out[19];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[5] = s_CSAwallace_rca12_csa0_csa_component_out[20];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[6] = s_CSAwallace_rca12_csa0_csa_component_out[21];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[7] = s_CSAwallace_rca12_csa0_csa_component_out[22];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[8] = s_CSAwallace_rca12_csa0_csa_component_out[23];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[9] = s_CSAwallace_rca12_csa0_csa_component_out[24];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[10] = s_CSAwallace_rca12_csa0_csa_component_out[25];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[11] = s_CSAwallace_rca12_csa0_csa_component_out[26];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[12] = s_CSAwallace_rca12_csa0_csa_component_out[27];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[13] = s_CSAwallace_rca12_csa0_csa_component_out[28];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[14] = 1'b1;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[15] = 1'b1;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[16] = 1'b1;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1[17] = 1'b1;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[0] = 1'b0;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[1] = 1'b0;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[2] = 1'b0;
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[3] = s_CSAwallace_rca12_csa1_csa_component_out[3];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[4] = s_CSAwallace_rca12_csa1_csa_component_out[4];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[5] = s_CSAwallace_rca12_csa1_csa_component_out[5];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[6] = s_CSAwallace_rca12_csa1_csa_component_out[6];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[7] = s_CSAwallace_rca12_csa1_csa_component_out[7];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[8] = s_CSAwallace_rca12_csa1_csa_component_out[8];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[9] = s_CSAwallace_rca12_csa1_csa_component_out[9];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[10] = s_CSAwallace_rca12_csa1_csa_component_out[10];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[11] = s_CSAwallace_rca12_csa1_csa_component_out[11];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[12] = s_CSAwallace_rca12_csa1_csa_component_out[12];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[13] = s_CSAwallace_rca12_csa1_csa_component_out[13];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[14] = s_CSAwallace_rca12_csa1_csa_component_out[14];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[15] = s_CSAwallace_rca12_csa1_csa_component_out[15];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[16] = s_CSAwallace_rca12_csa1_csa_component_out[16];
  assign s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2[17] = 1'b1;
  csa_component18 csa_component18_s_CSAwallace_rca12_csa4_csa_component_out(.a(s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s1), .b(s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_c1), .c(s_CSAwallace_rca12_csa4_csa_component_s_CSAwallace_rca12_csa_s2), .csa_component18_out(s_CSAwallace_rca12_csa4_csa_component_out));
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[0] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[1] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[2] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[3] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[4] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[5] = s_CSAwallace_rca12_csa1_csa_component_out[23];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[6] = s_CSAwallace_rca12_csa1_csa_component_out[24];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[7] = s_CSAwallace_rca12_csa1_csa_component_out[25];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[8] = s_CSAwallace_rca12_csa1_csa_component_out[26];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[9] = s_CSAwallace_rca12_csa1_csa_component_out[27];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[10] = s_CSAwallace_rca12_csa1_csa_component_out[28];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[11] = s_CSAwallace_rca12_csa1_csa_component_out[29];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[12] = s_CSAwallace_rca12_csa1_csa_component_out[30];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[13] = s_CSAwallace_rca12_csa1_csa_component_out[31];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[14] = s_CSAwallace_rca12_csa1_csa_component_out[32];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[15] = s_CSAwallace_rca12_csa1_csa_component_out[33];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[16] = s_CSAwallace_rca12_csa1_csa_component_out[34];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[17] = 1'b1;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[18] = 1'b1;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[19] = 1'b1;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2[20] = 1'b1;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[0] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[1] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[2] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[3] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[4] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[5] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[6] = s_CSAwallace_rca12_csa2_csa_component_out[6];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[7] = s_CSAwallace_rca12_csa2_csa_component_out[7];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[8] = s_CSAwallace_rca12_csa2_csa_component_out[8];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[9] = s_CSAwallace_rca12_csa2_csa_component_out[9];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[10] = s_CSAwallace_rca12_csa2_csa_component_out[10];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[11] = s_CSAwallace_rca12_csa2_csa_component_out[11];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[12] = s_CSAwallace_rca12_csa2_csa_component_out[12];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[13] = s_CSAwallace_rca12_csa2_csa_component_out[13];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[14] = s_CSAwallace_rca12_csa2_csa_component_out[14];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[15] = s_CSAwallace_rca12_csa2_csa_component_out[15];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[16] = s_CSAwallace_rca12_csa2_csa_component_out[16];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[17] = s_CSAwallace_rca12_csa2_csa_component_out[17];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[18] = s_CSAwallace_rca12_csa2_csa_component_out[18];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[19] = s_CSAwallace_rca12_csa2_csa_component_out[19];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3[20] = 1'b1;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[0] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[1] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[2] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[3] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[4] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[5] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[6] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[7] = 1'b0;
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[8] = s_CSAwallace_rca12_csa2_csa_component_out[29];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[9] = s_CSAwallace_rca12_csa2_csa_component_out[30];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[10] = s_CSAwallace_rca12_csa2_csa_component_out[31];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[11] = s_CSAwallace_rca12_csa2_csa_component_out[32];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[12] = s_CSAwallace_rca12_csa2_csa_component_out[33];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[13] = s_CSAwallace_rca12_csa2_csa_component_out[34];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[14] = s_CSAwallace_rca12_csa2_csa_component_out[35];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[15] = s_CSAwallace_rca12_csa2_csa_component_out[36];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[16] = s_CSAwallace_rca12_csa2_csa_component_out[37];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[17] = s_CSAwallace_rca12_csa2_csa_component_out[38];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[18] = s_CSAwallace_rca12_csa2_csa_component_out[39];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[19] = s_CSAwallace_rca12_csa2_csa_component_out[40];
  assign s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3[20] = 1'b1;
  csa_component21 csa_component21_s_CSAwallace_rca12_csa5_csa_component_out(.a(s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c2), .b(s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_s3), .c(s_CSAwallace_rca12_csa5_csa_component_s_CSAwallace_rca12_csa_c3), .csa_component21_out(s_CSAwallace_rca12_csa5_csa_component_out));
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[0] = s_CSAwallace_rca12_csa4_csa_component_out[0];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[1] = s_CSAwallace_rca12_csa4_csa_component_out[1];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[2] = s_CSAwallace_rca12_csa4_csa_component_out[2];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[3] = s_CSAwallace_rca12_csa4_csa_component_out[3];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[4] = s_CSAwallace_rca12_csa4_csa_component_out[4];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[5] = s_CSAwallace_rca12_csa4_csa_component_out[5];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[6] = s_CSAwallace_rca12_csa4_csa_component_out[6];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[7] = s_CSAwallace_rca12_csa4_csa_component_out[7];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[8] = s_CSAwallace_rca12_csa4_csa_component_out[8];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[9] = s_CSAwallace_rca12_csa4_csa_component_out[9];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[10] = s_CSAwallace_rca12_csa4_csa_component_out[10];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[11] = s_CSAwallace_rca12_csa4_csa_component_out[11];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[12] = s_CSAwallace_rca12_csa4_csa_component_out[12];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[13] = s_CSAwallace_rca12_csa4_csa_component_out[13];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[14] = s_CSAwallace_rca12_csa4_csa_component_out[14];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[15] = s_CSAwallace_rca12_csa4_csa_component_out[15];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[16] = s_CSAwallace_rca12_csa4_csa_component_out[16];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[17] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[18] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[19] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[20] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5[21] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[0] = 1'b0;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[1] = 1'b0;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[2] = 1'b0;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[3] = s_CSAwallace_rca12_csa4_csa_component_out[22];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[4] = s_CSAwallace_rca12_csa4_csa_component_out[23];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[5] = s_CSAwallace_rca12_csa4_csa_component_out[24];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[6] = s_CSAwallace_rca12_csa4_csa_component_out[25];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[7] = s_CSAwallace_rca12_csa4_csa_component_out[26];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[8] = s_CSAwallace_rca12_csa4_csa_component_out[27];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[9] = s_CSAwallace_rca12_csa4_csa_component_out[28];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[10] = s_CSAwallace_rca12_csa4_csa_component_out[29];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[11] = s_CSAwallace_rca12_csa4_csa_component_out[30];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[12] = s_CSAwallace_rca12_csa4_csa_component_out[31];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[13] = s_CSAwallace_rca12_csa4_csa_component_out[32];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[14] = s_CSAwallace_rca12_csa4_csa_component_out[33];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[15] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[16] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[17] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[18] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[19] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[20] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5[21] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[0] = 1'b0;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[1] = 1'b0;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[2] = 1'b0;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[3] = 1'b0;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[4] = 1'b0;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[5] = s_CSAwallace_rca12_csa5_csa_component_out[5];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[6] = s_CSAwallace_rca12_csa5_csa_component_out[6];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[7] = s_CSAwallace_rca12_csa5_csa_component_out[7];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[8] = s_CSAwallace_rca12_csa5_csa_component_out[8];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[9] = s_CSAwallace_rca12_csa5_csa_component_out[9];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[10] = s_CSAwallace_rca12_csa5_csa_component_out[10];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[11] = s_CSAwallace_rca12_csa5_csa_component_out[11];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[12] = s_CSAwallace_rca12_csa5_csa_component_out[12];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[13] = s_CSAwallace_rca12_csa5_csa_component_out[13];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[14] = s_CSAwallace_rca12_csa5_csa_component_out[14];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[15] = s_CSAwallace_rca12_csa5_csa_component_out[15];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[16] = s_CSAwallace_rca12_csa5_csa_component_out[16];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[17] = s_CSAwallace_rca12_csa5_csa_component_out[17];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[18] = s_CSAwallace_rca12_csa5_csa_component_out[18];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[19] = s_CSAwallace_rca12_csa5_csa_component_out[19];
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[20] = 1'b1;
  assign s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6[21] = 1'b1;
  csa_component22 csa_component22_s_CSAwallace_rca12_csa6_csa_component_out(.a(s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s5), .b(s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_c5), .c(s_CSAwallace_rca12_csa6_csa_component_s_CSAwallace_rca12_csa_s6), .csa_component22_out(s_CSAwallace_rca12_csa6_csa_component_out));
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[0] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[1] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[2] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[3] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[4] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[5] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[6] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[7] = s_CSAwallace_rca12_csa5_csa_component_out[29];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[8] = s_CSAwallace_rca12_csa5_csa_component_out[30];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[9] = s_CSAwallace_rca12_csa5_csa_component_out[31];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[10] = s_CSAwallace_rca12_csa5_csa_component_out[32];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[11] = s_CSAwallace_rca12_csa5_csa_component_out[33];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[12] = s_CSAwallace_rca12_csa5_csa_component_out[34];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[13] = s_CSAwallace_rca12_csa5_csa_component_out[35];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[14] = s_CSAwallace_rca12_csa5_csa_component_out[36];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[15] = s_CSAwallace_rca12_csa5_csa_component_out[37];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[16] = s_CSAwallace_rca12_csa5_csa_component_out[38];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[17] = s_CSAwallace_rca12_csa5_csa_component_out[39];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[18] = s_CSAwallace_rca12_csa5_csa_component_out[40];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[19] = s_CSAwallace_rca12_csa5_csa_component_out[41];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[20] = s_CSAwallace_rca12_csa5_csa_component_out[42];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[21] = 1'b1;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[22] = 1'b1;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6[23] = 1'b1;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[0] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[1] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[2] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[3] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[4] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[5] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[6] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[7] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[8] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[9] = s_CSAwallace_rca12_csa3_csa_component_out[9];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[10] = s_CSAwallace_rca12_csa3_csa_component_out[10];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[11] = s_CSAwallace_rca12_csa3_csa_component_out[11];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[12] = s_CSAwallace_rca12_csa3_csa_component_out[12];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[13] = s_CSAwallace_rca12_csa3_csa_component_out[13];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[14] = s_CSAwallace_rca12_csa3_csa_component_out[14];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[15] = s_CSAwallace_rca12_csa3_csa_component_out[15];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[16] = s_CSAwallace_rca12_csa3_csa_component_out[16];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[17] = s_CSAwallace_rca12_csa3_csa_component_out[17];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[18] = s_CSAwallace_rca12_csa3_csa_component_out[18];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[19] = s_CSAwallace_rca12_csa3_csa_component_out[19];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[20] = s_CSAwallace_rca12_csa3_csa_component_out[20];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[21] = s_CSAwallace_rca12_csa3_csa_component_out[21];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[22] = s_CSAwallace_rca12_csa3_csa_component_out[22];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4[23] = 1'b1;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[0] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[1] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[2] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[3] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[4] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[5] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[6] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[7] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[8] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[9] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[10] = 1'b0;
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[11] = s_CSAwallace_rca12_csa3_csa_component_out[35];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[12] = s_CSAwallace_rca12_csa3_csa_component_out[36];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[13] = s_CSAwallace_rca12_csa3_csa_component_out[37];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[14] = s_CSAwallace_rca12_csa3_csa_component_out[38];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[15] = s_CSAwallace_rca12_csa3_csa_component_out[39];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[16] = s_CSAwallace_rca12_csa3_csa_component_out[40];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[17] = s_CSAwallace_rca12_csa3_csa_component_out[41];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[18] = s_CSAwallace_rca12_csa3_csa_component_out[42];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[19] = s_CSAwallace_rca12_csa3_csa_component_out[43];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[20] = s_CSAwallace_rca12_csa3_csa_component_out[44];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[21] = s_CSAwallace_rca12_csa3_csa_component_out[45];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[22] = s_CSAwallace_rca12_csa3_csa_component_out[46];
  assign s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4[23] = 1'b1;
  csa_component24 csa_component24_s_CSAwallace_rca12_csa7_csa_component_out(.a(s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c6), .b(s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_s4), .c(s_CSAwallace_rca12_csa7_csa_component_s_CSAwallace_rca12_csa_c4), .csa_component24_out(s_CSAwallace_rca12_csa7_csa_component_out));
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[0] = s_CSAwallace_rca12_csa6_csa_component_out[0];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[1] = s_CSAwallace_rca12_csa6_csa_component_out[1];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[2] = s_CSAwallace_rca12_csa6_csa_component_out[2];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[3] = s_CSAwallace_rca12_csa6_csa_component_out[3];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[4] = s_CSAwallace_rca12_csa6_csa_component_out[4];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[5] = s_CSAwallace_rca12_csa6_csa_component_out[5];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[6] = s_CSAwallace_rca12_csa6_csa_component_out[6];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[7] = s_CSAwallace_rca12_csa6_csa_component_out[7];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[8] = s_CSAwallace_rca12_csa6_csa_component_out[8];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[9] = s_CSAwallace_rca12_csa6_csa_component_out[9];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[10] = s_CSAwallace_rca12_csa6_csa_component_out[10];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[11] = s_CSAwallace_rca12_csa6_csa_component_out[11];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[12] = s_CSAwallace_rca12_csa6_csa_component_out[12];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[13] = s_CSAwallace_rca12_csa6_csa_component_out[13];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[14] = s_CSAwallace_rca12_csa6_csa_component_out[14];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[15] = s_CSAwallace_rca12_csa6_csa_component_out[15];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[16] = s_CSAwallace_rca12_csa6_csa_component_out[16];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[17] = s_CSAwallace_rca12_csa6_csa_component_out[17];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[18] = s_CSAwallace_rca12_csa6_csa_component_out[18];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[19] = s_CSAwallace_rca12_csa6_csa_component_out[19];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[20] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[21] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[22] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7[23] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[0] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[1] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[2] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[3] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[4] = s_CSAwallace_rca12_csa6_csa_component_out[27];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[5] = s_CSAwallace_rca12_csa6_csa_component_out[28];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[6] = s_CSAwallace_rca12_csa6_csa_component_out[29];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[7] = s_CSAwallace_rca12_csa6_csa_component_out[30];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[8] = s_CSAwallace_rca12_csa6_csa_component_out[31];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[9] = s_CSAwallace_rca12_csa6_csa_component_out[32];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[10] = s_CSAwallace_rca12_csa6_csa_component_out[33];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[11] = s_CSAwallace_rca12_csa6_csa_component_out[34];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[12] = s_CSAwallace_rca12_csa6_csa_component_out[35];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[13] = s_CSAwallace_rca12_csa6_csa_component_out[36];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[14] = s_CSAwallace_rca12_csa6_csa_component_out[37];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[15] = s_CSAwallace_rca12_csa6_csa_component_out[38];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[16] = s_CSAwallace_rca12_csa6_csa_component_out[39];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[17] = s_CSAwallace_rca12_csa6_csa_component_out[40];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[18] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[19] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[20] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[21] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[22] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7[23] = 1'b1;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[0] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[1] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[2] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[3] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[4] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[5] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[6] = 1'b0;
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[7] = s_CSAwallace_rca12_csa7_csa_component_out[7];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[8] = s_CSAwallace_rca12_csa7_csa_component_out[8];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[9] = s_CSAwallace_rca12_csa7_csa_component_out[9];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[10] = s_CSAwallace_rca12_csa7_csa_component_out[10];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[11] = s_CSAwallace_rca12_csa7_csa_component_out[11];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[12] = s_CSAwallace_rca12_csa7_csa_component_out[12];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[13] = s_CSAwallace_rca12_csa7_csa_component_out[13];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[14] = s_CSAwallace_rca12_csa7_csa_component_out[14];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[15] = s_CSAwallace_rca12_csa7_csa_component_out[15];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[16] = s_CSAwallace_rca12_csa7_csa_component_out[16];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[17] = s_CSAwallace_rca12_csa7_csa_component_out[17];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[18] = s_CSAwallace_rca12_csa7_csa_component_out[18];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[19] = s_CSAwallace_rca12_csa7_csa_component_out[19];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[20] = s_CSAwallace_rca12_csa7_csa_component_out[20];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[21] = s_CSAwallace_rca12_csa7_csa_component_out[21];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[22] = s_CSAwallace_rca12_csa7_csa_component_out[22];
  assign s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8[23] = 1'b1;
  csa_component24 csa_component24_s_CSAwallace_rca12_csa8_csa_component_out(.a(s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s7), .b(s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_c7), .c(s_CSAwallace_rca12_csa8_csa_component_s_CSAwallace_rca12_csa_s8), .csa_component24_out(s_CSAwallace_rca12_csa8_csa_component_out));
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[0] = s_CSAwallace_rca12_csa8_csa_component_out[0];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[1] = s_CSAwallace_rca12_csa8_csa_component_out[1];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[2] = s_CSAwallace_rca12_csa8_csa_component_out[2];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[3] = s_CSAwallace_rca12_csa8_csa_component_out[3];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[4] = s_CSAwallace_rca12_csa8_csa_component_out[4];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[5] = s_CSAwallace_rca12_csa8_csa_component_out[5];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[6] = s_CSAwallace_rca12_csa8_csa_component_out[6];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[7] = s_CSAwallace_rca12_csa8_csa_component_out[7];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[8] = s_CSAwallace_rca12_csa8_csa_component_out[8];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[9] = s_CSAwallace_rca12_csa8_csa_component_out[9];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[10] = s_CSAwallace_rca12_csa8_csa_component_out[10];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[11] = s_CSAwallace_rca12_csa8_csa_component_out[11];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[12] = s_CSAwallace_rca12_csa8_csa_component_out[12];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[13] = s_CSAwallace_rca12_csa8_csa_component_out[13];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[14] = s_CSAwallace_rca12_csa8_csa_component_out[14];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[15] = s_CSAwallace_rca12_csa8_csa_component_out[15];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[16] = s_CSAwallace_rca12_csa8_csa_component_out[16];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[17] = s_CSAwallace_rca12_csa8_csa_component_out[17];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[18] = s_CSAwallace_rca12_csa8_csa_component_out[18];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[19] = s_CSAwallace_rca12_csa8_csa_component_out[19];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[20] = s_CSAwallace_rca12_csa8_csa_component_out[20];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[21] = s_CSAwallace_rca12_csa8_csa_component_out[21];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[22] = s_CSAwallace_rca12_csa8_csa_component_out[22];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9[23] = 1'b1;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[0] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[1] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[2] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[3] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[4] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[5] = s_CSAwallace_rca12_csa8_csa_component_out[30];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[6] = s_CSAwallace_rca12_csa8_csa_component_out[31];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[7] = s_CSAwallace_rca12_csa8_csa_component_out[32];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[8] = s_CSAwallace_rca12_csa8_csa_component_out[33];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[9] = s_CSAwallace_rca12_csa8_csa_component_out[34];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[10] = s_CSAwallace_rca12_csa8_csa_component_out[35];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[11] = s_CSAwallace_rca12_csa8_csa_component_out[36];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[12] = s_CSAwallace_rca12_csa8_csa_component_out[37];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[13] = s_CSAwallace_rca12_csa8_csa_component_out[38];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[14] = s_CSAwallace_rca12_csa8_csa_component_out[39];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[15] = s_CSAwallace_rca12_csa8_csa_component_out[40];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[16] = s_CSAwallace_rca12_csa8_csa_component_out[41];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[17] = s_CSAwallace_rca12_csa8_csa_component_out[42];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[18] = s_CSAwallace_rca12_csa8_csa_component_out[43];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[19] = s_CSAwallace_rca12_csa8_csa_component_out[44];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[20] = s_CSAwallace_rca12_csa8_csa_component_out[45];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[21] = 1'b1;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[22] = 1'b1;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9[23] = 1'b1;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[0] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[1] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[2] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[3] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[4] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[5] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[6] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[7] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[8] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[9] = 1'b0;
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[10] = s_CSAwallace_rca12_csa7_csa_component_out[35];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[11] = s_CSAwallace_rca12_csa7_csa_component_out[36];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[12] = s_CSAwallace_rca12_csa7_csa_component_out[37];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[13] = s_CSAwallace_rca12_csa7_csa_component_out[38];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[14] = s_CSAwallace_rca12_csa7_csa_component_out[39];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[15] = s_CSAwallace_rca12_csa7_csa_component_out[40];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[16] = s_CSAwallace_rca12_csa7_csa_component_out[41];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[17] = s_CSAwallace_rca12_csa7_csa_component_out[42];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[18] = s_CSAwallace_rca12_csa7_csa_component_out[43];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[19] = s_CSAwallace_rca12_csa7_csa_component_out[44];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[20] = s_CSAwallace_rca12_csa7_csa_component_out[45];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[21] = s_CSAwallace_rca12_csa7_csa_component_out[46];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[22] = s_CSAwallace_rca12_csa7_csa_component_out[47];
  assign s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8[23] = s_CSAwallace_rca12_csa7_csa_component_out[48];
  csa_component24 csa_component24_s_CSAwallace_rca12_csa9_csa_component_out(.a(s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_s9), .b(s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c9), .c(s_CSAwallace_rca12_csa9_csa_component_s_CSAwallace_rca12_csa_c8), .csa_component24_out(s_CSAwallace_rca12_csa9_csa_component_out));
  assign s_CSAwallace_rca12_u_rca24_a[0] = s_CSAwallace_rca12_csa9_csa_component_out[0];
  assign s_CSAwallace_rca12_u_rca24_a[1] = s_CSAwallace_rca12_csa9_csa_component_out[1];
  assign s_CSAwallace_rca12_u_rca24_a[2] = s_CSAwallace_rca12_csa9_csa_component_out[2];
  assign s_CSAwallace_rca12_u_rca24_a[3] = s_CSAwallace_rca12_csa9_csa_component_out[3];
  assign s_CSAwallace_rca12_u_rca24_a[4] = s_CSAwallace_rca12_csa9_csa_component_out[4];
  assign s_CSAwallace_rca12_u_rca24_a[5] = s_CSAwallace_rca12_csa9_csa_component_out[5];
  assign s_CSAwallace_rca12_u_rca24_a[6] = s_CSAwallace_rca12_csa9_csa_component_out[6];
  assign s_CSAwallace_rca12_u_rca24_a[7] = s_CSAwallace_rca12_csa9_csa_component_out[7];
  assign s_CSAwallace_rca12_u_rca24_a[8] = s_CSAwallace_rca12_csa9_csa_component_out[8];
  assign s_CSAwallace_rca12_u_rca24_a[9] = s_CSAwallace_rca12_csa9_csa_component_out[9];
  assign s_CSAwallace_rca12_u_rca24_a[10] = s_CSAwallace_rca12_csa9_csa_component_out[10];
  assign s_CSAwallace_rca12_u_rca24_a[11] = s_CSAwallace_rca12_csa9_csa_component_out[11];
  assign s_CSAwallace_rca12_u_rca24_a[12] = s_CSAwallace_rca12_csa9_csa_component_out[12];
  assign s_CSAwallace_rca12_u_rca24_a[13] = s_CSAwallace_rca12_csa9_csa_component_out[13];
  assign s_CSAwallace_rca12_u_rca24_a[14] = s_CSAwallace_rca12_csa9_csa_component_out[14];
  assign s_CSAwallace_rca12_u_rca24_a[15] = s_CSAwallace_rca12_csa9_csa_component_out[15];
  assign s_CSAwallace_rca12_u_rca24_a[16] = s_CSAwallace_rca12_csa9_csa_component_out[16];
  assign s_CSAwallace_rca12_u_rca24_a[17] = s_CSAwallace_rca12_csa9_csa_component_out[17];
  assign s_CSAwallace_rca12_u_rca24_a[18] = s_CSAwallace_rca12_csa9_csa_component_out[18];
  assign s_CSAwallace_rca12_u_rca24_a[19] = s_CSAwallace_rca12_csa9_csa_component_out[19];
  assign s_CSAwallace_rca12_u_rca24_a[20] = s_CSAwallace_rca12_csa9_csa_component_out[20];
  assign s_CSAwallace_rca12_u_rca24_a[21] = s_CSAwallace_rca12_csa9_csa_component_out[21];
  assign s_CSAwallace_rca12_u_rca24_a[22] = s_CSAwallace_rca12_csa9_csa_component_out[22];
  assign s_CSAwallace_rca12_u_rca24_a[23] = s_CSAwallace_rca12_csa9_csa_component_out[23];
  assign s_CSAwallace_rca12_u_rca24_b[0] = 1'b0;
  assign s_CSAwallace_rca12_u_rca24_b[1] = 1'b0;
  assign s_CSAwallace_rca12_u_rca24_b[2] = 1'b0;
  assign s_CSAwallace_rca12_u_rca24_b[3] = 1'b0;
  assign s_CSAwallace_rca12_u_rca24_b[4] = 1'b0;
  assign s_CSAwallace_rca12_u_rca24_b[5] = 1'b0;
  assign s_CSAwallace_rca12_u_rca24_b[6] = s_CSAwallace_rca12_csa9_csa_component_out[31];
  assign s_CSAwallace_rca12_u_rca24_b[7] = s_CSAwallace_rca12_csa9_csa_component_out[32];
  assign s_CSAwallace_rca12_u_rca24_b[8] = s_CSAwallace_rca12_csa9_csa_component_out[33];
  assign s_CSAwallace_rca12_u_rca24_b[9] = s_CSAwallace_rca12_csa9_csa_component_out[34];
  assign s_CSAwallace_rca12_u_rca24_b[10] = s_CSAwallace_rca12_csa9_csa_component_out[35];
  assign s_CSAwallace_rca12_u_rca24_b[11] = s_CSAwallace_rca12_csa9_csa_component_out[36];
  assign s_CSAwallace_rca12_u_rca24_b[12] = s_CSAwallace_rca12_csa9_csa_component_out[37];
  assign s_CSAwallace_rca12_u_rca24_b[13] = s_CSAwallace_rca12_csa9_csa_component_out[38];
  assign s_CSAwallace_rca12_u_rca24_b[14] = s_CSAwallace_rca12_csa9_csa_component_out[39];
  assign s_CSAwallace_rca12_u_rca24_b[15] = s_CSAwallace_rca12_csa9_csa_component_out[40];
  assign s_CSAwallace_rca12_u_rca24_b[16] = s_CSAwallace_rca12_csa9_csa_component_out[41];
  assign s_CSAwallace_rca12_u_rca24_b[17] = s_CSAwallace_rca12_csa9_csa_component_out[42];
  assign s_CSAwallace_rca12_u_rca24_b[18] = s_CSAwallace_rca12_csa9_csa_component_out[43];
  assign s_CSAwallace_rca12_u_rca24_b[19] = s_CSAwallace_rca12_csa9_csa_component_out[44];
  assign s_CSAwallace_rca12_u_rca24_b[20] = s_CSAwallace_rca12_csa9_csa_component_out[45];
  assign s_CSAwallace_rca12_u_rca24_b[21] = s_CSAwallace_rca12_csa9_csa_component_out[46];
  assign s_CSAwallace_rca12_u_rca24_b[22] = s_CSAwallace_rca12_csa9_csa_component_out[47];
  assign s_CSAwallace_rca12_u_rca24_b[23] = s_CSAwallace_rca12_csa9_csa_component_out[48];
  u_rca24 u_rca24_s_CSAwallace_rca12_u_rca24_out(.a(s_CSAwallace_rca12_u_rca24_a), .b(s_CSAwallace_rca12_u_rca24_b), .u_rca24_out(s_CSAwallace_rca12_u_rca24_out));
  not_gate not_gate_s_CSAwallace_rca12_xor0(.a(s_CSAwallace_rca12_u_rca24_out[23]), .out(s_CSAwallace_rca12_xor0));

  assign s_CSAwallace_rca12_out[0] = s_CSAwallace_rca12_u_rca24_out[0];
  assign s_CSAwallace_rca12_out[1] = s_CSAwallace_rca12_u_rca24_out[1];
  assign s_CSAwallace_rca12_out[2] = s_CSAwallace_rca12_u_rca24_out[2];
  assign s_CSAwallace_rca12_out[3] = s_CSAwallace_rca12_u_rca24_out[3];
  assign s_CSAwallace_rca12_out[4] = s_CSAwallace_rca12_u_rca24_out[4];
  assign s_CSAwallace_rca12_out[5] = s_CSAwallace_rca12_u_rca24_out[5];
  assign s_CSAwallace_rca12_out[6] = s_CSAwallace_rca12_u_rca24_out[6];
  assign s_CSAwallace_rca12_out[7] = s_CSAwallace_rca12_u_rca24_out[7];
  assign s_CSAwallace_rca12_out[8] = s_CSAwallace_rca12_u_rca24_out[8];
  assign s_CSAwallace_rca12_out[9] = s_CSAwallace_rca12_u_rca24_out[9];
  assign s_CSAwallace_rca12_out[10] = s_CSAwallace_rca12_u_rca24_out[10];
  assign s_CSAwallace_rca12_out[11] = s_CSAwallace_rca12_u_rca24_out[11];
  assign s_CSAwallace_rca12_out[12] = s_CSAwallace_rca12_u_rca24_out[12];
  assign s_CSAwallace_rca12_out[13] = s_CSAwallace_rca12_u_rca24_out[13];
  assign s_CSAwallace_rca12_out[14] = s_CSAwallace_rca12_u_rca24_out[14];
  assign s_CSAwallace_rca12_out[15] = s_CSAwallace_rca12_u_rca24_out[15];
  assign s_CSAwallace_rca12_out[16] = s_CSAwallace_rca12_u_rca24_out[16];
  assign s_CSAwallace_rca12_out[17] = s_CSAwallace_rca12_u_rca24_out[17];
  assign s_CSAwallace_rca12_out[18] = s_CSAwallace_rca12_u_rca24_out[18];
  assign s_CSAwallace_rca12_out[19] = s_CSAwallace_rca12_u_rca24_out[19];
  assign s_CSAwallace_rca12_out[20] = s_CSAwallace_rca12_u_rca24_out[20];
  assign s_CSAwallace_rca12_out[21] = s_CSAwallace_rca12_u_rca24_out[21];
  assign s_CSAwallace_rca12_out[22] = s_CSAwallace_rca12_u_rca24_out[22];
  assign s_CSAwallace_rca12_out[23] = s_CSAwallace_rca12_xor0[0];
endmodule