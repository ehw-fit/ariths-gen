module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(a[0], b[0], pg_logic_or0);
  and_gate and_gate_pg_logic_and0(a[0], b[0], pg_logic_and0);
  xor_gate xor_gate_pg_logic_xor0(a[0], b[0], pg_logic_xor0);
endmodule

module h_s_cla24(input [23:0] a, input [23:0] b, output [24:0] h_s_cla24_out);
  wire [0:0] h_s_cla24_pg_logic0_or0;
  wire [0:0] h_s_cla24_pg_logic0_and0;
  wire [0:0] h_s_cla24_pg_logic0_xor0;
  wire [0:0] h_s_cla24_pg_logic1_or0;
  wire [0:0] h_s_cla24_pg_logic1_and0;
  wire [0:0] h_s_cla24_pg_logic1_xor0;
  wire [0:0] h_s_cla24_xor1;
  wire [0:0] h_s_cla24_and0;
  wire [0:0] h_s_cla24_or0;
  wire [0:0] h_s_cla24_pg_logic2_or0;
  wire [0:0] h_s_cla24_pg_logic2_and0;
  wire [0:0] h_s_cla24_pg_logic2_xor0;
  wire [0:0] h_s_cla24_xor2;
  wire [0:0] h_s_cla24_and1;
  wire [0:0] h_s_cla24_and2;
  wire [0:0] h_s_cla24_and3;
  wire [0:0] h_s_cla24_and4;
  wire [0:0] h_s_cla24_or1;
  wire [0:0] h_s_cla24_or2;
  wire [0:0] h_s_cla24_pg_logic3_or0;
  wire [0:0] h_s_cla24_pg_logic3_and0;
  wire [0:0] h_s_cla24_pg_logic3_xor0;
  wire [0:0] h_s_cla24_xor3;
  wire [0:0] h_s_cla24_and5;
  wire [0:0] h_s_cla24_and6;
  wire [0:0] h_s_cla24_and7;
  wire [0:0] h_s_cla24_and8;
  wire [0:0] h_s_cla24_and9;
  wire [0:0] h_s_cla24_and10;
  wire [0:0] h_s_cla24_and11;
  wire [0:0] h_s_cla24_or3;
  wire [0:0] h_s_cla24_or4;
  wire [0:0] h_s_cla24_or5;
  wire [0:0] h_s_cla24_pg_logic4_or0;
  wire [0:0] h_s_cla24_pg_logic4_and0;
  wire [0:0] h_s_cla24_pg_logic4_xor0;
  wire [0:0] h_s_cla24_xor4;
  wire [0:0] h_s_cla24_and12;
  wire [0:0] h_s_cla24_or6;
  wire [0:0] h_s_cla24_pg_logic5_or0;
  wire [0:0] h_s_cla24_pg_logic5_and0;
  wire [0:0] h_s_cla24_pg_logic5_xor0;
  wire [0:0] h_s_cla24_xor5;
  wire [0:0] h_s_cla24_and13;
  wire [0:0] h_s_cla24_and14;
  wire [0:0] h_s_cla24_and15;
  wire [0:0] h_s_cla24_or7;
  wire [0:0] h_s_cla24_or8;
  wire [0:0] h_s_cla24_pg_logic6_or0;
  wire [0:0] h_s_cla24_pg_logic6_and0;
  wire [0:0] h_s_cla24_pg_logic6_xor0;
  wire [0:0] h_s_cla24_xor6;
  wire [0:0] h_s_cla24_and16;
  wire [0:0] h_s_cla24_and17;
  wire [0:0] h_s_cla24_and18;
  wire [0:0] h_s_cla24_and19;
  wire [0:0] h_s_cla24_and20;
  wire [0:0] h_s_cla24_and21;
  wire [0:0] h_s_cla24_or9;
  wire [0:0] h_s_cla24_or10;
  wire [0:0] h_s_cla24_or11;
  wire [0:0] h_s_cla24_pg_logic7_or0;
  wire [0:0] h_s_cla24_pg_logic7_and0;
  wire [0:0] h_s_cla24_pg_logic7_xor0;
  wire [0:0] h_s_cla24_xor7;
  wire [0:0] h_s_cla24_and22;
  wire [0:0] h_s_cla24_and23;
  wire [0:0] h_s_cla24_and24;
  wire [0:0] h_s_cla24_and25;
  wire [0:0] h_s_cla24_and26;
  wire [0:0] h_s_cla24_and27;
  wire [0:0] h_s_cla24_and28;
  wire [0:0] h_s_cla24_and29;
  wire [0:0] h_s_cla24_and30;
  wire [0:0] h_s_cla24_and31;
  wire [0:0] h_s_cla24_or12;
  wire [0:0] h_s_cla24_or13;
  wire [0:0] h_s_cla24_or14;
  wire [0:0] h_s_cla24_or15;
  wire [0:0] h_s_cla24_pg_logic8_or0;
  wire [0:0] h_s_cla24_pg_logic8_and0;
  wire [0:0] h_s_cla24_pg_logic8_xor0;
  wire [0:0] h_s_cla24_xor8;
  wire [0:0] h_s_cla24_and32;
  wire [0:0] h_s_cla24_or16;
  wire [0:0] h_s_cla24_pg_logic9_or0;
  wire [0:0] h_s_cla24_pg_logic9_and0;
  wire [0:0] h_s_cla24_pg_logic9_xor0;
  wire [0:0] h_s_cla24_xor9;
  wire [0:0] h_s_cla24_and33;
  wire [0:0] h_s_cla24_and34;
  wire [0:0] h_s_cla24_and35;
  wire [0:0] h_s_cla24_or17;
  wire [0:0] h_s_cla24_or18;
  wire [0:0] h_s_cla24_pg_logic10_or0;
  wire [0:0] h_s_cla24_pg_logic10_and0;
  wire [0:0] h_s_cla24_pg_logic10_xor0;
  wire [0:0] h_s_cla24_xor10;
  wire [0:0] h_s_cla24_and36;
  wire [0:0] h_s_cla24_and37;
  wire [0:0] h_s_cla24_and38;
  wire [0:0] h_s_cla24_and39;
  wire [0:0] h_s_cla24_and40;
  wire [0:0] h_s_cla24_and41;
  wire [0:0] h_s_cla24_or19;
  wire [0:0] h_s_cla24_or20;
  wire [0:0] h_s_cla24_or21;
  wire [0:0] h_s_cla24_pg_logic11_or0;
  wire [0:0] h_s_cla24_pg_logic11_and0;
  wire [0:0] h_s_cla24_pg_logic11_xor0;
  wire [0:0] h_s_cla24_xor11;
  wire [0:0] h_s_cla24_and42;
  wire [0:0] h_s_cla24_and43;
  wire [0:0] h_s_cla24_and44;
  wire [0:0] h_s_cla24_and45;
  wire [0:0] h_s_cla24_and46;
  wire [0:0] h_s_cla24_and47;
  wire [0:0] h_s_cla24_and48;
  wire [0:0] h_s_cla24_and49;
  wire [0:0] h_s_cla24_and50;
  wire [0:0] h_s_cla24_and51;
  wire [0:0] h_s_cla24_or22;
  wire [0:0] h_s_cla24_or23;
  wire [0:0] h_s_cla24_or24;
  wire [0:0] h_s_cla24_or25;
  wire [0:0] h_s_cla24_pg_logic12_or0;
  wire [0:0] h_s_cla24_pg_logic12_and0;
  wire [0:0] h_s_cla24_pg_logic12_xor0;
  wire [0:0] h_s_cla24_xor12;
  wire [0:0] h_s_cla24_and52;
  wire [0:0] h_s_cla24_or26;
  wire [0:0] h_s_cla24_pg_logic13_or0;
  wire [0:0] h_s_cla24_pg_logic13_and0;
  wire [0:0] h_s_cla24_pg_logic13_xor0;
  wire [0:0] h_s_cla24_xor13;
  wire [0:0] h_s_cla24_and53;
  wire [0:0] h_s_cla24_and54;
  wire [0:0] h_s_cla24_and55;
  wire [0:0] h_s_cla24_or27;
  wire [0:0] h_s_cla24_or28;
  wire [0:0] h_s_cla24_pg_logic14_or0;
  wire [0:0] h_s_cla24_pg_logic14_and0;
  wire [0:0] h_s_cla24_pg_logic14_xor0;
  wire [0:0] h_s_cla24_xor14;
  wire [0:0] h_s_cla24_and56;
  wire [0:0] h_s_cla24_and57;
  wire [0:0] h_s_cla24_and58;
  wire [0:0] h_s_cla24_and59;
  wire [0:0] h_s_cla24_and60;
  wire [0:0] h_s_cla24_and61;
  wire [0:0] h_s_cla24_or29;
  wire [0:0] h_s_cla24_or30;
  wire [0:0] h_s_cla24_or31;
  wire [0:0] h_s_cla24_pg_logic15_or0;
  wire [0:0] h_s_cla24_pg_logic15_and0;
  wire [0:0] h_s_cla24_pg_logic15_xor0;
  wire [0:0] h_s_cla24_xor15;
  wire [0:0] h_s_cla24_and62;
  wire [0:0] h_s_cla24_and63;
  wire [0:0] h_s_cla24_and64;
  wire [0:0] h_s_cla24_and65;
  wire [0:0] h_s_cla24_and66;
  wire [0:0] h_s_cla24_and67;
  wire [0:0] h_s_cla24_and68;
  wire [0:0] h_s_cla24_and69;
  wire [0:0] h_s_cla24_and70;
  wire [0:0] h_s_cla24_and71;
  wire [0:0] h_s_cla24_or32;
  wire [0:0] h_s_cla24_or33;
  wire [0:0] h_s_cla24_or34;
  wire [0:0] h_s_cla24_or35;
  wire [0:0] h_s_cla24_pg_logic16_or0;
  wire [0:0] h_s_cla24_pg_logic16_and0;
  wire [0:0] h_s_cla24_pg_logic16_xor0;
  wire [0:0] h_s_cla24_xor16;
  wire [0:0] h_s_cla24_and72;
  wire [0:0] h_s_cla24_or36;
  wire [0:0] h_s_cla24_pg_logic17_or0;
  wire [0:0] h_s_cla24_pg_logic17_and0;
  wire [0:0] h_s_cla24_pg_logic17_xor0;
  wire [0:0] h_s_cla24_xor17;
  wire [0:0] h_s_cla24_and73;
  wire [0:0] h_s_cla24_and74;
  wire [0:0] h_s_cla24_and75;
  wire [0:0] h_s_cla24_or37;
  wire [0:0] h_s_cla24_or38;
  wire [0:0] h_s_cla24_pg_logic18_or0;
  wire [0:0] h_s_cla24_pg_logic18_and0;
  wire [0:0] h_s_cla24_pg_logic18_xor0;
  wire [0:0] h_s_cla24_xor18;
  wire [0:0] h_s_cla24_and76;
  wire [0:0] h_s_cla24_and77;
  wire [0:0] h_s_cla24_and78;
  wire [0:0] h_s_cla24_and79;
  wire [0:0] h_s_cla24_and80;
  wire [0:0] h_s_cla24_and81;
  wire [0:0] h_s_cla24_or39;
  wire [0:0] h_s_cla24_or40;
  wire [0:0] h_s_cla24_or41;
  wire [0:0] h_s_cla24_pg_logic19_or0;
  wire [0:0] h_s_cla24_pg_logic19_and0;
  wire [0:0] h_s_cla24_pg_logic19_xor0;
  wire [0:0] h_s_cla24_xor19;
  wire [0:0] h_s_cla24_and82;
  wire [0:0] h_s_cla24_and83;
  wire [0:0] h_s_cla24_and84;
  wire [0:0] h_s_cla24_and85;
  wire [0:0] h_s_cla24_and86;
  wire [0:0] h_s_cla24_and87;
  wire [0:0] h_s_cla24_and88;
  wire [0:0] h_s_cla24_and89;
  wire [0:0] h_s_cla24_and90;
  wire [0:0] h_s_cla24_and91;
  wire [0:0] h_s_cla24_or42;
  wire [0:0] h_s_cla24_or43;
  wire [0:0] h_s_cla24_or44;
  wire [0:0] h_s_cla24_or45;
  wire [0:0] h_s_cla24_pg_logic20_or0;
  wire [0:0] h_s_cla24_pg_logic20_and0;
  wire [0:0] h_s_cla24_pg_logic20_xor0;
  wire [0:0] h_s_cla24_xor20;
  wire [0:0] h_s_cla24_and92;
  wire [0:0] h_s_cla24_or46;
  wire [0:0] h_s_cla24_pg_logic21_or0;
  wire [0:0] h_s_cla24_pg_logic21_and0;
  wire [0:0] h_s_cla24_pg_logic21_xor0;
  wire [0:0] h_s_cla24_xor21;
  wire [0:0] h_s_cla24_and93;
  wire [0:0] h_s_cla24_and94;
  wire [0:0] h_s_cla24_and95;
  wire [0:0] h_s_cla24_or47;
  wire [0:0] h_s_cla24_or48;
  wire [0:0] h_s_cla24_pg_logic22_or0;
  wire [0:0] h_s_cla24_pg_logic22_and0;
  wire [0:0] h_s_cla24_pg_logic22_xor0;
  wire [0:0] h_s_cla24_xor22;
  wire [0:0] h_s_cla24_and96;
  wire [0:0] h_s_cla24_and97;
  wire [0:0] h_s_cla24_and98;
  wire [0:0] h_s_cla24_and99;
  wire [0:0] h_s_cla24_and100;
  wire [0:0] h_s_cla24_and101;
  wire [0:0] h_s_cla24_or49;
  wire [0:0] h_s_cla24_or50;
  wire [0:0] h_s_cla24_or51;
  wire [0:0] h_s_cla24_pg_logic23_or0;
  wire [0:0] h_s_cla24_pg_logic23_and0;
  wire [0:0] h_s_cla24_pg_logic23_xor0;
  wire [0:0] h_s_cla24_xor23;
  wire [0:0] h_s_cla24_and102;
  wire [0:0] h_s_cla24_and103;
  wire [0:0] h_s_cla24_and104;
  wire [0:0] h_s_cla24_and105;
  wire [0:0] h_s_cla24_and106;
  wire [0:0] h_s_cla24_and107;
  wire [0:0] h_s_cla24_and108;
  wire [0:0] h_s_cla24_and109;
  wire [0:0] h_s_cla24_and110;
  wire [0:0] h_s_cla24_and111;
  wire [0:0] h_s_cla24_or52;
  wire [0:0] h_s_cla24_or53;
  wire [0:0] h_s_cla24_or54;
  wire [0:0] h_s_cla24_or55;
  wire [0:0] h_s_cla24_xor24;
  wire [0:0] h_s_cla24_xor25;

  pg_logic pg_logic_h_s_cla24_pg_logic0_out(a[0], b[0], h_s_cla24_pg_logic0_or0, h_s_cla24_pg_logic0_and0, h_s_cla24_pg_logic0_xor0);
  pg_logic pg_logic_h_s_cla24_pg_logic1_out(a[1], b[1], h_s_cla24_pg_logic1_or0, h_s_cla24_pg_logic1_and0, h_s_cla24_pg_logic1_xor0);
  xor_gate xor_gate_h_s_cla24_xor1(h_s_cla24_pg_logic1_xor0[0], h_s_cla24_pg_logic0_and0[0], h_s_cla24_xor1);
  and_gate and_gate_h_s_cla24_and0(h_s_cla24_pg_logic0_and0[0], h_s_cla24_pg_logic1_or0[0], h_s_cla24_and0);
  or_gate or_gate_h_s_cla24_or0(h_s_cla24_pg_logic1_and0[0], h_s_cla24_and0[0], h_s_cla24_or0);
  pg_logic pg_logic_h_s_cla24_pg_logic2_out(a[2], b[2], h_s_cla24_pg_logic2_or0, h_s_cla24_pg_logic2_and0, h_s_cla24_pg_logic2_xor0);
  xor_gate xor_gate_h_s_cla24_xor2(h_s_cla24_pg_logic2_xor0[0], h_s_cla24_or0[0], h_s_cla24_xor2);
  and_gate and_gate_h_s_cla24_and1(h_s_cla24_pg_logic2_or0[0], h_s_cla24_pg_logic0_or0[0], h_s_cla24_and1);
  and_gate and_gate_h_s_cla24_and2(h_s_cla24_pg_logic0_and0[0], h_s_cla24_pg_logic2_or0[0], h_s_cla24_and2);
  and_gate and_gate_h_s_cla24_and3(h_s_cla24_and2[0], h_s_cla24_pg_logic1_or0[0], h_s_cla24_and3);
  and_gate and_gate_h_s_cla24_and4(h_s_cla24_pg_logic1_and0[0], h_s_cla24_pg_logic2_or0[0], h_s_cla24_and4);
  or_gate or_gate_h_s_cla24_or1(h_s_cla24_and3[0], h_s_cla24_and4[0], h_s_cla24_or1);
  or_gate or_gate_h_s_cla24_or2(h_s_cla24_pg_logic2_and0[0], h_s_cla24_or1[0], h_s_cla24_or2);
  pg_logic pg_logic_h_s_cla24_pg_logic3_out(a[3], b[3], h_s_cla24_pg_logic3_or0, h_s_cla24_pg_logic3_and0, h_s_cla24_pg_logic3_xor0);
  xor_gate xor_gate_h_s_cla24_xor3(h_s_cla24_pg_logic3_xor0[0], h_s_cla24_or2[0], h_s_cla24_xor3);
  and_gate and_gate_h_s_cla24_and5(h_s_cla24_pg_logic3_or0[0], h_s_cla24_pg_logic1_or0[0], h_s_cla24_and5);
  and_gate and_gate_h_s_cla24_and6(h_s_cla24_pg_logic0_and0[0], h_s_cla24_pg_logic2_or0[0], h_s_cla24_and6);
  and_gate and_gate_h_s_cla24_and7(h_s_cla24_pg_logic3_or0[0], h_s_cla24_pg_logic1_or0[0], h_s_cla24_and7);
  and_gate and_gate_h_s_cla24_and8(h_s_cla24_and6[0], h_s_cla24_and7[0], h_s_cla24_and8);
  and_gate and_gate_h_s_cla24_and9(h_s_cla24_pg_logic1_and0[0], h_s_cla24_pg_logic3_or0[0], h_s_cla24_and9);
  and_gate and_gate_h_s_cla24_and10(h_s_cla24_and9[0], h_s_cla24_pg_logic2_or0[0], h_s_cla24_and10);
  and_gate and_gate_h_s_cla24_and11(h_s_cla24_pg_logic2_and0[0], h_s_cla24_pg_logic3_or0[0], h_s_cla24_and11);
  or_gate or_gate_h_s_cla24_or3(h_s_cla24_and8[0], h_s_cla24_and11[0], h_s_cla24_or3);
  or_gate or_gate_h_s_cla24_or4(h_s_cla24_and10[0], h_s_cla24_or3[0], h_s_cla24_or4);
  or_gate or_gate_h_s_cla24_or5(h_s_cla24_pg_logic3_and0[0], h_s_cla24_or4[0], h_s_cla24_or5);
  pg_logic pg_logic_h_s_cla24_pg_logic4_out(a[4], b[4], h_s_cla24_pg_logic4_or0, h_s_cla24_pg_logic4_and0, h_s_cla24_pg_logic4_xor0);
  xor_gate xor_gate_h_s_cla24_xor4(h_s_cla24_pg_logic4_xor0[0], h_s_cla24_or5[0], h_s_cla24_xor4);
  and_gate and_gate_h_s_cla24_and12(h_s_cla24_or5[0], h_s_cla24_pg_logic4_or0[0], h_s_cla24_and12);
  or_gate or_gate_h_s_cla24_or6(h_s_cla24_pg_logic4_and0[0], h_s_cla24_and12[0], h_s_cla24_or6);
  pg_logic pg_logic_h_s_cla24_pg_logic5_out(a[5], b[5], h_s_cla24_pg_logic5_or0, h_s_cla24_pg_logic5_and0, h_s_cla24_pg_logic5_xor0);
  xor_gate xor_gate_h_s_cla24_xor5(h_s_cla24_pg_logic5_xor0[0], h_s_cla24_or6[0], h_s_cla24_xor5);
  and_gate and_gate_h_s_cla24_and13(h_s_cla24_or5[0], h_s_cla24_pg_logic5_or0[0], h_s_cla24_and13);
  and_gate and_gate_h_s_cla24_and14(h_s_cla24_and13[0], h_s_cla24_pg_logic4_or0[0], h_s_cla24_and14);
  and_gate and_gate_h_s_cla24_and15(h_s_cla24_pg_logic4_and0[0], h_s_cla24_pg_logic5_or0[0], h_s_cla24_and15);
  or_gate or_gate_h_s_cla24_or7(h_s_cla24_and14[0], h_s_cla24_and15[0], h_s_cla24_or7);
  or_gate or_gate_h_s_cla24_or8(h_s_cla24_pg_logic5_and0[0], h_s_cla24_or7[0], h_s_cla24_or8);
  pg_logic pg_logic_h_s_cla24_pg_logic6_out(a[6], b[6], h_s_cla24_pg_logic6_or0, h_s_cla24_pg_logic6_and0, h_s_cla24_pg_logic6_xor0);
  xor_gate xor_gate_h_s_cla24_xor6(h_s_cla24_pg_logic6_xor0[0], h_s_cla24_or8[0], h_s_cla24_xor6);
  and_gate and_gate_h_s_cla24_and16(h_s_cla24_or5[0], h_s_cla24_pg_logic5_or0[0], h_s_cla24_and16);
  and_gate and_gate_h_s_cla24_and17(h_s_cla24_pg_logic6_or0[0], h_s_cla24_pg_logic4_or0[0], h_s_cla24_and17);
  and_gate and_gate_h_s_cla24_and18(h_s_cla24_and16[0], h_s_cla24_and17[0], h_s_cla24_and18);
  and_gate and_gate_h_s_cla24_and19(h_s_cla24_pg_logic4_and0[0], h_s_cla24_pg_logic6_or0[0], h_s_cla24_and19);
  and_gate and_gate_h_s_cla24_and20(h_s_cla24_and19[0], h_s_cla24_pg_logic5_or0[0], h_s_cla24_and20);
  and_gate and_gate_h_s_cla24_and21(h_s_cla24_pg_logic5_and0[0], h_s_cla24_pg_logic6_or0[0], h_s_cla24_and21);
  or_gate or_gate_h_s_cla24_or9(h_s_cla24_and18[0], h_s_cla24_and20[0], h_s_cla24_or9);
  or_gate or_gate_h_s_cla24_or10(h_s_cla24_or9[0], h_s_cla24_and21[0], h_s_cla24_or10);
  or_gate or_gate_h_s_cla24_or11(h_s_cla24_pg_logic6_and0[0], h_s_cla24_or10[0], h_s_cla24_or11);
  pg_logic pg_logic_h_s_cla24_pg_logic7_out(a[7], b[7], h_s_cla24_pg_logic7_or0, h_s_cla24_pg_logic7_and0, h_s_cla24_pg_logic7_xor0);
  xor_gate xor_gate_h_s_cla24_xor7(h_s_cla24_pg_logic7_xor0[0], h_s_cla24_or11[0], h_s_cla24_xor7);
  and_gate and_gate_h_s_cla24_and22(h_s_cla24_or5[0], h_s_cla24_pg_logic6_or0[0], h_s_cla24_and22);
  and_gate and_gate_h_s_cla24_and23(h_s_cla24_pg_logic7_or0[0], h_s_cla24_pg_logic5_or0[0], h_s_cla24_and23);
  and_gate and_gate_h_s_cla24_and24(h_s_cla24_and22[0], h_s_cla24_and23[0], h_s_cla24_and24);
  and_gate and_gate_h_s_cla24_and25(h_s_cla24_and24[0], h_s_cla24_pg_logic4_or0[0], h_s_cla24_and25);
  and_gate and_gate_h_s_cla24_and26(h_s_cla24_pg_logic4_and0[0], h_s_cla24_pg_logic6_or0[0], h_s_cla24_and26);
  and_gate and_gate_h_s_cla24_and27(h_s_cla24_pg_logic7_or0[0], h_s_cla24_pg_logic5_or0[0], h_s_cla24_and27);
  and_gate and_gate_h_s_cla24_and28(h_s_cla24_and26[0], h_s_cla24_and27[0], h_s_cla24_and28);
  and_gate and_gate_h_s_cla24_and29(h_s_cla24_pg_logic5_and0[0], h_s_cla24_pg_logic7_or0[0], h_s_cla24_and29);
  and_gate and_gate_h_s_cla24_and30(h_s_cla24_and29[0], h_s_cla24_pg_logic6_or0[0], h_s_cla24_and30);
  and_gate and_gate_h_s_cla24_and31(h_s_cla24_pg_logic6_and0[0], h_s_cla24_pg_logic7_or0[0], h_s_cla24_and31);
  or_gate or_gate_h_s_cla24_or12(h_s_cla24_and25[0], h_s_cla24_and30[0], h_s_cla24_or12);
  or_gate or_gate_h_s_cla24_or13(h_s_cla24_and28[0], h_s_cla24_and31[0], h_s_cla24_or13);
  or_gate or_gate_h_s_cla24_or14(h_s_cla24_or12[0], h_s_cla24_or13[0], h_s_cla24_or14);
  or_gate or_gate_h_s_cla24_or15(h_s_cla24_pg_logic7_and0[0], h_s_cla24_or14[0], h_s_cla24_or15);
  pg_logic pg_logic_h_s_cla24_pg_logic8_out(a[8], b[8], h_s_cla24_pg_logic8_or0, h_s_cla24_pg_logic8_and0, h_s_cla24_pg_logic8_xor0);
  xor_gate xor_gate_h_s_cla24_xor8(h_s_cla24_pg_logic8_xor0[0], h_s_cla24_or15[0], h_s_cla24_xor8);
  and_gate and_gate_h_s_cla24_and32(h_s_cla24_or15[0], h_s_cla24_pg_logic8_or0[0], h_s_cla24_and32);
  or_gate or_gate_h_s_cla24_or16(h_s_cla24_pg_logic8_and0[0], h_s_cla24_and32[0], h_s_cla24_or16);
  pg_logic pg_logic_h_s_cla24_pg_logic9_out(a[9], b[9], h_s_cla24_pg_logic9_or0, h_s_cla24_pg_logic9_and0, h_s_cla24_pg_logic9_xor0);
  xor_gate xor_gate_h_s_cla24_xor9(h_s_cla24_pg_logic9_xor0[0], h_s_cla24_or16[0], h_s_cla24_xor9);
  and_gate and_gate_h_s_cla24_and33(h_s_cla24_or15[0], h_s_cla24_pg_logic9_or0[0], h_s_cla24_and33);
  and_gate and_gate_h_s_cla24_and34(h_s_cla24_and33[0], h_s_cla24_pg_logic8_or0[0], h_s_cla24_and34);
  and_gate and_gate_h_s_cla24_and35(h_s_cla24_pg_logic8_and0[0], h_s_cla24_pg_logic9_or0[0], h_s_cla24_and35);
  or_gate or_gate_h_s_cla24_or17(h_s_cla24_and34[0], h_s_cla24_and35[0], h_s_cla24_or17);
  or_gate or_gate_h_s_cla24_or18(h_s_cla24_pg_logic9_and0[0], h_s_cla24_or17[0], h_s_cla24_or18);
  pg_logic pg_logic_h_s_cla24_pg_logic10_out(a[10], b[10], h_s_cla24_pg_logic10_or0, h_s_cla24_pg_logic10_and0, h_s_cla24_pg_logic10_xor0);
  xor_gate xor_gate_h_s_cla24_xor10(h_s_cla24_pg_logic10_xor0[0], h_s_cla24_or18[0], h_s_cla24_xor10);
  and_gate and_gate_h_s_cla24_and36(h_s_cla24_or15[0], h_s_cla24_pg_logic9_or0[0], h_s_cla24_and36);
  and_gate and_gate_h_s_cla24_and37(h_s_cla24_pg_logic10_or0[0], h_s_cla24_pg_logic8_or0[0], h_s_cla24_and37);
  and_gate and_gate_h_s_cla24_and38(h_s_cla24_and36[0], h_s_cla24_and37[0], h_s_cla24_and38);
  and_gate and_gate_h_s_cla24_and39(h_s_cla24_pg_logic8_and0[0], h_s_cla24_pg_logic10_or0[0], h_s_cla24_and39);
  and_gate and_gate_h_s_cla24_and40(h_s_cla24_and39[0], h_s_cla24_pg_logic9_or0[0], h_s_cla24_and40);
  and_gate and_gate_h_s_cla24_and41(h_s_cla24_pg_logic9_and0[0], h_s_cla24_pg_logic10_or0[0], h_s_cla24_and41);
  or_gate or_gate_h_s_cla24_or19(h_s_cla24_and38[0], h_s_cla24_and40[0], h_s_cla24_or19);
  or_gate or_gate_h_s_cla24_or20(h_s_cla24_or19[0], h_s_cla24_and41[0], h_s_cla24_or20);
  or_gate or_gate_h_s_cla24_or21(h_s_cla24_pg_logic10_and0[0], h_s_cla24_or20[0], h_s_cla24_or21);
  pg_logic pg_logic_h_s_cla24_pg_logic11_out(a[11], b[11], h_s_cla24_pg_logic11_or0, h_s_cla24_pg_logic11_and0, h_s_cla24_pg_logic11_xor0);
  xor_gate xor_gate_h_s_cla24_xor11(h_s_cla24_pg_logic11_xor0[0], h_s_cla24_or21[0], h_s_cla24_xor11);
  and_gate and_gate_h_s_cla24_and42(h_s_cla24_or15[0], h_s_cla24_pg_logic10_or0[0], h_s_cla24_and42);
  and_gate and_gate_h_s_cla24_and43(h_s_cla24_pg_logic11_or0[0], h_s_cla24_pg_logic9_or0[0], h_s_cla24_and43);
  and_gate and_gate_h_s_cla24_and44(h_s_cla24_and42[0], h_s_cla24_and43[0], h_s_cla24_and44);
  and_gate and_gate_h_s_cla24_and45(h_s_cla24_and44[0], h_s_cla24_pg_logic8_or0[0], h_s_cla24_and45);
  and_gate and_gate_h_s_cla24_and46(h_s_cla24_pg_logic8_and0[0], h_s_cla24_pg_logic10_or0[0], h_s_cla24_and46);
  and_gate and_gate_h_s_cla24_and47(h_s_cla24_pg_logic11_or0[0], h_s_cla24_pg_logic9_or0[0], h_s_cla24_and47);
  and_gate and_gate_h_s_cla24_and48(h_s_cla24_and46[0], h_s_cla24_and47[0], h_s_cla24_and48);
  and_gate and_gate_h_s_cla24_and49(h_s_cla24_pg_logic9_and0[0], h_s_cla24_pg_logic11_or0[0], h_s_cla24_and49);
  and_gate and_gate_h_s_cla24_and50(h_s_cla24_and49[0], h_s_cla24_pg_logic10_or0[0], h_s_cla24_and50);
  and_gate and_gate_h_s_cla24_and51(h_s_cla24_pg_logic10_and0[0], h_s_cla24_pg_logic11_or0[0], h_s_cla24_and51);
  or_gate or_gate_h_s_cla24_or22(h_s_cla24_and45[0], h_s_cla24_and50[0], h_s_cla24_or22);
  or_gate or_gate_h_s_cla24_or23(h_s_cla24_and48[0], h_s_cla24_and51[0], h_s_cla24_or23);
  or_gate or_gate_h_s_cla24_or24(h_s_cla24_or22[0], h_s_cla24_or23[0], h_s_cla24_or24);
  or_gate or_gate_h_s_cla24_or25(h_s_cla24_pg_logic11_and0[0], h_s_cla24_or24[0], h_s_cla24_or25);
  pg_logic pg_logic_h_s_cla24_pg_logic12_out(a[12], b[12], h_s_cla24_pg_logic12_or0, h_s_cla24_pg_logic12_and0, h_s_cla24_pg_logic12_xor0);
  xor_gate xor_gate_h_s_cla24_xor12(h_s_cla24_pg_logic12_xor0[0], h_s_cla24_or25[0], h_s_cla24_xor12);
  and_gate and_gate_h_s_cla24_and52(h_s_cla24_or25[0], h_s_cla24_pg_logic12_or0[0], h_s_cla24_and52);
  or_gate or_gate_h_s_cla24_or26(h_s_cla24_pg_logic12_and0[0], h_s_cla24_and52[0], h_s_cla24_or26);
  pg_logic pg_logic_h_s_cla24_pg_logic13_out(a[13], b[13], h_s_cla24_pg_logic13_or0, h_s_cla24_pg_logic13_and0, h_s_cla24_pg_logic13_xor0);
  xor_gate xor_gate_h_s_cla24_xor13(h_s_cla24_pg_logic13_xor0[0], h_s_cla24_or26[0], h_s_cla24_xor13);
  and_gate and_gate_h_s_cla24_and53(h_s_cla24_or25[0], h_s_cla24_pg_logic13_or0[0], h_s_cla24_and53);
  and_gate and_gate_h_s_cla24_and54(h_s_cla24_and53[0], h_s_cla24_pg_logic12_or0[0], h_s_cla24_and54);
  and_gate and_gate_h_s_cla24_and55(h_s_cla24_pg_logic12_and0[0], h_s_cla24_pg_logic13_or0[0], h_s_cla24_and55);
  or_gate or_gate_h_s_cla24_or27(h_s_cla24_and54[0], h_s_cla24_and55[0], h_s_cla24_or27);
  or_gate or_gate_h_s_cla24_or28(h_s_cla24_pg_logic13_and0[0], h_s_cla24_or27[0], h_s_cla24_or28);
  pg_logic pg_logic_h_s_cla24_pg_logic14_out(a[14], b[14], h_s_cla24_pg_logic14_or0, h_s_cla24_pg_logic14_and0, h_s_cla24_pg_logic14_xor0);
  xor_gate xor_gate_h_s_cla24_xor14(h_s_cla24_pg_logic14_xor0[0], h_s_cla24_or28[0], h_s_cla24_xor14);
  and_gate and_gate_h_s_cla24_and56(h_s_cla24_or25[0], h_s_cla24_pg_logic13_or0[0], h_s_cla24_and56);
  and_gate and_gate_h_s_cla24_and57(h_s_cla24_pg_logic14_or0[0], h_s_cla24_pg_logic12_or0[0], h_s_cla24_and57);
  and_gate and_gate_h_s_cla24_and58(h_s_cla24_and56[0], h_s_cla24_and57[0], h_s_cla24_and58);
  and_gate and_gate_h_s_cla24_and59(h_s_cla24_pg_logic12_and0[0], h_s_cla24_pg_logic14_or0[0], h_s_cla24_and59);
  and_gate and_gate_h_s_cla24_and60(h_s_cla24_and59[0], h_s_cla24_pg_logic13_or0[0], h_s_cla24_and60);
  and_gate and_gate_h_s_cla24_and61(h_s_cla24_pg_logic13_and0[0], h_s_cla24_pg_logic14_or0[0], h_s_cla24_and61);
  or_gate or_gate_h_s_cla24_or29(h_s_cla24_and58[0], h_s_cla24_and60[0], h_s_cla24_or29);
  or_gate or_gate_h_s_cla24_or30(h_s_cla24_or29[0], h_s_cla24_and61[0], h_s_cla24_or30);
  or_gate or_gate_h_s_cla24_or31(h_s_cla24_pg_logic14_and0[0], h_s_cla24_or30[0], h_s_cla24_or31);
  pg_logic pg_logic_h_s_cla24_pg_logic15_out(a[15], b[15], h_s_cla24_pg_logic15_or0, h_s_cla24_pg_logic15_and0, h_s_cla24_pg_logic15_xor0);
  xor_gate xor_gate_h_s_cla24_xor15(h_s_cla24_pg_logic15_xor0[0], h_s_cla24_or31[0], h_s_cla24_xor15);
  and_gate and_gate_h_s_cla24_and62(h_s_cla24_or25[0], h_s_cla24_pg_logic14_or0[0], h_s_cla24_and62);
  and_gate and_gate_h_s_cla24_and63(h_s_cla24_pg_logic15_or0[0], h_s_cla24_pg_logic13_or0[0], h_s_cla24_and63);
  and_gate and_gate_h_s_cla24_and64(h_s_cla24_and62[0], h_s_cla24_and63[0], h_s_cla24_and64);
  and_gate and_gate_h_s_cla24_and65(h_s_cla24_and64[0], h_s_cla24_pg_logic12_or0[0], h_s_cla24_and65);
  and_gate and_gate_h_s_cla24_and66(h_s_cla24_pg_logic12_and0[0], h_s_cla24_pg_logic14_or0[0], h_s_cla24_and66);
  and_gate and_gate_h_s_cla24_and67(h_s_cla24_pg_logic15_or0[0], h_s_cla24_pg_logic13_or0[0], h_s_cla24_and67);
  and_gate and_gate_h_s_cla24_and68(h_s_cla24_and66[0], h_s_cla24_and67[0], h_s_cla24_and68);
  and_gate and_gate_h_s_cla24_and69(h_s_cla24_pg_logic13_and0[0], h_s_cla24_pg_logic15_or0[0], h_s_cla24_and69);
  and_gate and_gate_h_s_cla24_and70(h_s_cla24_and69[0], h_s_cla24_pg_logic14_or0[0], h_s_cla24_and70);
  and_gate and_gate_h_s_cla24_and71(h_s_cla24_pg_logic14_and0[0], h_s_cla24_pg_logic15_or0[0], h_s_cla24_and71);
  or_gate or_gate_h_s_cla24_or32(h_s_cla24_and65[0], h_s_cla24_and70[0], h_s_cla24_or32);
  or_gate or_gate_h_s_cla24_or33(h_s_cla24_and68[0], h_s_cla24_and71[0], h_s_cla24_or33);
  or_gate or_gate_h_s_cla24_or34(h_s_cla24_or32[0], h_s_cla24_or33[0], h_s_cla24_or34);
  or_gate or_gate_h_s_cla24_or35(h_s_cla24_pg_logic15_and0[0], h_s_cla24_or34[0], h_s_cla24_or35);
  pg_logic pg_logic_h_s_cla24_pg_logic16_out(a[16], b[16], h_s_cla24_pg_logic16_or0, h_s_cla24_pg_logic16_and0, h_s_cla24_pg_logic16_xor0);
  xor_gate xor_gate_h_s_cla24_xor16(h_s_cla24_pg_logic16_xor0[0], h_s_cla24_or35[0], h_s_cla24_xor16);
  and_gate and_gate_h_s_cla24_and72(h_s_cla24_or35[0], h_s_cla24_pg_logic16_or0[0], h_s_cla24_and72);
  or_gate or_gate_h_s_cla24_or36(h_s_cla24_pg_logic16_and0[0], h_s_cla24_and72[0], h_s_cla24_or36);
  pg_logic pg_logic_h_s_cla24_pg_logic17_out(a[17], b[17], h_s_cla24_pg_logic17_or0, h_s_cla24_pg_logic17_and0, h_s_cla24_pg_logic17_xor0);
  xor_gate xor_gate_h_s_cla24_xor17(h_s_cla24_pg_logic17_xor0[0], h_s_cla24_or36[0], h_s_cla24_xor17);
  and_gate and_gate_h_s_cla24_and73(h_s_cla24_or35[0], h_s_cla24_pg_logic17_or0[0], h_s_cla24_and73);
  and_gate and_gate_h_s_cla24_and74(h_s_cla24_and73[0], h_s_cla24_pg_logic16_or0[0], h_s_cla24_and74);
  and_gate and_gate_h_s_cla24_and75(h_s_cla24_pg_logic16_and0[0], h_s_cla24_pg_logic17_or0[0], h_s_cla24_and75);
  or_gate or_gate_h_s_cla24_or37(h_s_cla24_and74[0], h_s_cla24_and75[0], h_s_cla24_or37);
  or_gate or_gate_h_s_cla24_or38(h_s_cla24_pg_logic17_and0[0], h_s_cla24_or37[0], h_s_cla24_or38);
  pg_logic pg_logic_h_s_cla24_pg_logic18_out(a[18], b[18], h_s_cla24_pg_logic18_or0, h_s_cla24_pg_logic18_and0, h_s_cla24_pg_logic18_xor0);
  xor_gate xor_gate_h_s_cla24_xor18(h_s_cla24_pg_logic18_xor0[0], h_s_cla24_or38[0], h_s_cla24_xor18);
  and_gate and_gate_h_s_cla24_and76(h_s_cla24_or35[0], h_s_cla24_pg_logic17_or0[0], h_s_cla24_and76);
  and_gate and_gate_h_s_cla24_and77(h_s_cla24_pg_logic18_or0[0], h_s_cla24_pg_logic16_or0[0], h_s_cla24_and77);
  and_gate and_gate_h_s_cla24_and78(h_s_cla24_and76[0], h_s_cla24_and77[0], h_s_cla24_and78);
  and_gate and_gate_h_s_cla24_and79(h_s_cla24_pg_logic16_and0[0], h_s_cla24_pg_logic18_or0[0], h_s_cla24_and79);
  and_gate and_gate_h_s_cla24_and80(h_s_cla24_and79[0], h_s_cla24_pg_logic17_or0[0], h_s_cla24_and80);
  and_gate and_gate_h_s_cla24_and81(h_s_cla24_pg_logic17_and0[0], h_s_cla24_pg_logic18_or0[0], h_s_cla24_and81);
  or_gate or_gate_h_s_cla24_or39(h_s_cla24_and78[0], h_s_cla24_and80[0], h_s_cla24_or39);
  or_gate or_gate_h_s_cla24_or40(h_s_cla24_or39[0], h_s_cla24_and81[0], h_s_cla24_or40);
  or_gate or_gate_h_s_cla24_or41(h_s_cla24_pg_logic18_and0[0], h_s_cla24_or40[0], h_s_cla24_or41);
  pg_logic pg_logic_h_s_cla24_pg_logic19_out(a[19], b[19], h_s_cla24_pg_logic19_or0, h_s_cla24_pg_logic19_and0, h_s_cla24_pg_logic19_xor0);
  xor_gate xor_gate_h_s_cla24_xor19(h_s_cla24_pg_logic19_xor0[0], h_s_cla24_or41[0], h_s_cla24_xor19);
  and_gate and_gate_h_s_cla24_and82(h_s_cla24_or35[0], h_s_cla24_pg_logic18_or0[0], h_s_cla24_and82);
  and_gate and_gate_h_s_cla24_and83(h_s_cla24_pg_logic19_or0[0], h_s_cla24_pg_logic17_or0[0], h_s_cla24_and83);
  and_gate and_gate_h_s_cla24_and84(h_s_cla24_and82[0], h_s_cla24_and83[0], h_s_cla24_and84);
  and_gate and_gate_h_s_cla24_and85(h_s_cla24_and84[0], h_s_cla24_pg_logic16_or0[0], h_s_cla24_and85);
  and_gate and_gate_h_s_cla24_and86(h_s_cla24_pg_logic16_and0[0], h_s_cla24_pg_logic18_or0[0], h_s_cla24_and86);
  and_gate and_gate_h_s_cla24_and87(h_s_cla24_pg_logic19_or0[0], h_s_cla24_pg_logic17_or0[0], h_s_cla24_and87);
  and_gate and_gate_h_s_cla24_and88(h_s_cla24_and86[0], h_s_cla24_and87[0], h_s_cla24_and88);
  and_gate and_gate_h_s_cla24_and89(h_s_cla24_pg_logic17_and0[0], h_s_cla24_pg_logic19_or0[0], h_s_cla24_and89);
  and_gate and_gate_h_s_cla24_and90(h_s_cla24_and89[0], h_s_cla24_pg_logic18_or0[0], h_s_cla24_and90);
  and_gate and_gate_h_s_cla24_and91(h_s_cla24_pg_logic18_and0[0], h_s_cla24_pg_logic19_or0[0], h_s_cla24_and91);
  or_gate or_gate_h_s_cla24_or42(h_s_cla24_and85[0], h_s_cla24_and90[0], h_s_cla24_or42);
  or_gate or_gate_h_s_cla24_or43(h_s_cla24_and88[0], h_s_cla24_and91[0], h_s_cla24_or43);
  or_gate or_gate_h_s_cla24_or44(h_s_cla24_or42[0], h_s_cla24_or43[0], h_s_cla24_or44);
  or_gate or_gate_h_s_cla24_or45(h_s_cla24_pg_logic19_and0[0], h_s_cla24_or44[0], h_s_cla24_or45);
  pg_logic pg_logic_h_s_cla24_pg_logic20_out(a[20], b[20], h_s_cla24_pg_logic20_or0, h_s_cla24_pg_logic20_and0, h_s_cla24_pg_logic20_xor0);
  xor_gate xor_gate_h_s_cla24_xor20(h_s_cla24_pg_logic20_xor0[0], h_s_cla24_or45[0], h_s_cla24_xor20);
  and_gate and_gate_h_s_cla24_and92(h_s_cla24_or45[0], h_s_cla24_pg_logic20_or0[0], h_s_cla24_and92);
  or_gate or_gate_h_s_cla24_or46(h_s_cla24_pg_logic20_and0[0], h_s_cla24_and92[0], h_s_cla24_or46);
  pg_logic pg_logic_h_s_cla24_pg_logic21_out(a[21], b[21], h_s_cla24_pg_logic21_or0, h_s_cla24_pg_logic21_and0, h_s_cla24_pg_logic21_xor0);
  xor_gate xor_gate_h_s_cla24_xor21(h_s_cla24_pg_logic21_xor0[0], h_s_cla24_or46[0], h_s_cla24_xor21);
  and_gate and_gate_h_s_cla24_and93(h_s_cla24_or45[0], h_s_cla24_pg_logic21_or0[0], h_s_cla24_and93);
  and_gate and_gate_h_s_cla24_and94(h_s_cla24_and93[0], h_s_cla24_pg_logic20_or0[0], h_s_cla24_and94);
  and_gate and_gate_h_s_cla24_and95(h_s_cla24_pg_logic20_and0[0], h_s_cla24_pg_logic21_or0[0], h_s_cla24_and95);
  or_gate or_gate_h_s_cla24_or47(h_s_cla24_and94[0], h_s_cla24_and95[0], h_s_cla24_or47);
  or_gate or_gate_h_s_cla24_or48(h_s_cla24_pg_logic21_and0[0], h_s_cla24_or47[0], h_s_cla24_or48);
  pg_logic pg_logic_h_s_cla24_pg_logic22_out(a[22], b[22], h_s_cla24_pg_logic22_or0, h_s_cla24_pg_logic22_and0, h_s_cla24_pg_logic22_xor0);
  xor_gate xor_gate_h_s_cla24_xor22(h_s_cla24_pg_logic22_xor0[0], h_s_cla24_or48[0], h_s_cla24_xor22);
  and_gate and_gate_h_s_cla24_and96(h_s_cla24_or45[0], h_s_cla24_pg_logic21_or0[0], h_s_cla24_and96);
  and_gate and_gate_h_s_cla24_and97(h_s_cla24_pg_logic22_or0[0], h_s_cla24_pg_logic20_or0[0], h_s_cla24_and97);
  and_gate and_gate_h_s_cla24_and98(h_s_cla24_and96[0], h_s_cla24_and97[0], h_s_cla24_and98);
  and_gate and_gate_h_s_cla24_and99(h_s_cla24_pg_logic20_and0[0], h_s_cla24_pg_logic22_or0[0], h_s_cla24_and99);
  and_gate and_gate_h_s_cla24_and100(h_s_cla24_and99[0], h_s_cla24_pg_logic21_or0[0], h_s_cla24_and100);
  and_gate and_gate_h_s_cla24_and101(h_s_cla24_pg_logic21_and0[0], h_s_cla24_pg_logic22_or0[0], h_s_cla24_and101);
  or_gate or_gate_h_s_cla24_or49(h_s_cla24_and98[0], h_s_cla24_and100[0], h_s_cla24_or49);
  or_gate or_gate_h_s_cla24_or50(h_s_cla24_or49[0], h_s_cla24_and101[0], h_s_cla24_or50);
  or_gate or_gate_h_s_cla24_or51(h_s_cla24_pg_logic22_and0[0], h_s_cla24_or50[0], h_s_cla24_or51);
  pg_logic pg_logic_h_s_cla24_pg_logic23_out(a[23], b[23], h_s_cla24_pg_logic23_or0, h_s_cla24_pg_logic23_and0, h_s_cla24_pg_logic23_xor0);
  xor_gate xor_gate_h_s_cla24_xor23(h_s_cla24_pg_logic23_xor0[0], h_s_cla24_or51[0], h_s_cla24_xor23);
  and_gate and_gate_h_s_cla24_and102(h_s_cla24_or45[0], h_s_cla24_pg_logic22_or0[0], h_s_cla24_and102);
  and_gate and_gate_h_s_cla24_and103(h_s_cla24_pg_logic23_or0[0], h_s_cla24_pg_logic21_or0[0], h_s_cla24_and103);
  and_gate and_gate_h_s_cla24_and104(h_s_cla24_and102[0], h_s_cla24_and103[0], h_s_cla24_and104);
  and_gate and_gate_h_s_cla24_and105(h_s_cla24_and104[0], h_s_cla24_pg_logic20_or0[0], h_s_cla24_and105);
  and_gate and_gate_h_s_cla24_and106(h_s_cla24_pg_logic20_and0[0], h_s_cla24_pg_logic22_or0[0], h_s_cla24_and106);
  and_gate and_gate_h_s_cla24_and107(h_s_cla24_pg_logic23_or0[0], h_s_cla24_pg_logic21_or0[0], h_s_cla24_and107);
  and_gate and_gate_h_s_cla24_and108(h_s_cla24_and106[0], h_s_cla24_and107[0], h_s_cla24_and108);
  and_gate and_gate_h_s_cla24_and109(h_s_cla24_pg_logic21_and0[0], h_s_cla24_pg_logic23_or0[0], h_s_cla24_and109);
  and_gate and_gate_h_s_cla24_and110(h_s_cla24_and109[0], h_s_cla24_pg_logic22_or0[0], h_s_cla24_and110);
  and_gate and_gate_h_s_cla24_and111(h_s_cla24_pg_logic22_and0[0], h_s_cla24_pg_logic23_or0[0], h_s_cla24_and111);
  or_gate or_gate_h_s_cla24_or52(h_s_cla24_and105[0], h_s_cla24_and110[0], h_s_cla24_or52);
  or_gate or_gate_h_s_cla24_or53(h_s_cla24_and108[0], h_s_cla24_and111[0], h_s_cla24_or53);
  or_gate or_gate_h_s_cla24_or54(h_s_cla24_or52[0], h_s_cla24_or53[0], h_s_cla24_or54);
  or_gate or_gate_h_s_cla24_or55(h_s_cla24_pg_logic23_and0[0], h_s_cla24_or54[0], h_s_cla24_or55);
  xor_gate xor_gate_h_s_cla24_xor24(a[23], b[23], h_s_cla24_xor24);
  xor_gate xor_gate_h_s_cla24_xor25(h_s_cla24_xor24[0], h_s_cla24_or55[0], h_s_cla24_xor25);

  assign h_s_cla24_out[0] = h_s_cla24_pg_logic0_xor0[0];
  assign h_s_cla24_out[1] = h_s_cla24_xor1[0];
  assign h_s_cla24_out[2] = h_s_cla24_xor2[0];
  assign h_s_cla24_out[3] = h_s_cla24_xor3[0];
  assign h_s_cla24_out[4] = h_s_cla24_xor4[0];
  assign h_s_cla24_out[5] = h_s_cla24_xor5[0];
  assign h_s_cla24_out[6] = h_s_cla24_xor6[0];
  assign h_s_cla24_out[7] = h_s_cla24_xor7[0];
  assign h_s_cla24_out[8] = h_s_cla24_xor8[0];
  assign h_s_cla24_out[9] = h_s_cla24_xor9[0];
  assign h_s_cla24_out[10] = h_s_cla24_xor10[0];
  assign h_s_cla24_out[11] = h_s_cla24_xor11[0];
  assign h_s_cla24_out[12] = h_s_cla24_xor12[0];
  assign h_s_cla24_out[13] = h_s_cla24_xor13[0];
  assign h_s_cla24_out[14] = h_s_cla24_xor14[0];
  assign h_s_cla24_out[15] = h_s_cla24_xor15[0];
  assign h_s_cla24_out[16] = h_s_cla24_xor16[0];
  assign h_s_cla24_out[17] = h_s_cla24_xor17[0];
  assign h_s_cla24_out[18] = h_s_cla24_xor18[0];
  assign h_s_cla24_out[19] = h_s_cla24_xor19[0];
  assign h_s_cla24_out[20] = h_s_cla24_xor20[0];
  assign h_s_cla24_out[21] = h_s_cla24_xor21[0];
  assign h_s_cla24_out[22] = h_s_cla24_xor22[0];
  assign h_s_cla24_out[23] = h_s_cla24_xor23[0];
  assign h_s_cla24_out[24] = h_s_cla24_xor25[0];
endmodule