module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module nand_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a & _b);
endmodule

module constant_wire_value_1(input a, input b, output constant_wire_1);
  wire constant_wire_value_1_a;
  wire constant_wire_value_1_b;

  assign constant_wire_value_1_a = a;
  assign constant_wire_value_1_b = b;

  xor_gate xor_gate_constant_wire_value_1_y0(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y0);
  xnor_gate xnor_gate_constant_wire_value_1_y1(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y1);
  or_gate or_gate_constant_wire_1(constant_wire_value_1_y0, constant_wire_value_1_y1, constant_wire_1);
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_cin;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module u_rca(input [13:0] a, input [13:0] b, output [14:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire u_rca_ha_y0;
  wire u_rca_ha_y1;
  wire u_rca_fa1_y2;
  wire u_rca_fa1_y4;
  wire u_rca_fa2_y2;
  wire u_rca_fa2_y4;
  wire u_rca_fa3_y2;
  wire u_rca_fa3_y4;
  wire u_rca_fa4_y2;
  wire u_rca_fa4_y4;
  wire u_rca_fa5_y2;
  wire u_rca_fa5_y4;
  wire u_rca_fa6_y2;
  wire u_rca_fa6_y4;
  wire u_rca_fa7_y2;
  wire u_rca_fa7_y4;
  wire u_rca_fa8_y2;
  wire u_rca_fa8_y4;
  wire u_rca_fa9_y2;
  wire u_rca_fa9_y4;
  wire u_rca_fa10_y2;
  wire u_rca_fa10_y4;
  wire u_rca_fa11_y2;
  wire u_rca_fa11_y4;
  wire u_rca_fa12_y2;
  wire u_rca_fa12_y4;
  wire u_rca_fa13_y2;
  wire u_rca_fa13_y4;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  ha ha_u_rca_ha_y0(a_0, b_0, u_rca_ha_y0, u_rca_ha_y1);
  fa fa_u_rca_fa1_y2(a_1, b_1, u_rca_ha_y1, u_rca_fa1_y2, u_rca_fa1_y4);
  fa fa_u_rca_fa2_y2(a_2, b_2, u_rca_fa1_y4, u_rca_fa2_y2, u_rca_fa2_y4);
  fa fa_u_rca_fa3_y2(a_3, b_3, u_rca_fa2_y4, u_rca_fa3_y2, u_rca_fa3_y4);
  fa fa_u_rca_fa4_y2(a_4, b_4, u_rca_fa3_y4, u_rca_fa4_y2, u_rca_fa4_y4);
  fa fa_u_rca_fa5_y2(a_5, b_5, u_rca_fa4_y4, u_rca_fa5_y2, u_rca_fa5_y4);
  fa fa_u_rca_fa6_y2(a_6, b_6, u_rca_fa5_y4, u_rca_fa6_y2, u_rca_fa6_y4);
  fa fa_u_rca_fa7_y2(a_7, b_7, u_rca_fa6_y4, u_rca_fa7_y2, u_rca_fa7_y4);
  fa fa_u_rca_fa8_y2(a_8, b_8, u_rca_fa7_y4, u_rca_fa8_y2, u_rca_fa8_y4);
  fa fa_u_rca_fa9_y2(a_9, b_9, u_rca_fa8_y4, u_rca_fa9_y2, u_rca_fa9_y4);
  fa fa_u_rca_fa10_y2(a_10, b_10, u_rca_fa9_y4, u_rca_fa10_y2, u_rca_fa10_y4);
  fa fa_u_rca_fa11_y2(a_11, b_11, u_rca_fa10_y4, u_rca_fa11_y2, u_rca_fa11_y4);
  fa fa_u_rca_fa12_y2(a_12, b_12, u_rca_fa11_y4, u_rca_fa12_y2, u_rca_fa12_y4);
  fa fa_u_rca_fa13_y2(a_13, b_13, u_rca_fa12_y4, u_rca_fa13_y2, u_rca_fa13_y4);

  assign out[0] = u_rca_ha_y0;
  assign out[1] = u_rca_fa1_y2;
  assign out[2] = u_rca_fa2_y2;
  assign out[3] = u_rca_fa3_y2;
  assign out[4] = u_rca_fa4_y2;
  assign out[5] = u_rca_fa5_y2;
  assign out[6] = u_rca_fa6_y2;
  assign out[7] = u_rca_fa7_y2;
  assign out[8] = u_rca_fa8_y2;
  assign out[9] = u_rca_fa9_y2;
  assign out[10] = u_rca_fa10_y2;
  assign out[11] = u_rca_fa11_y2;
  assign out[12] = u_rca_fa12_y2;
  assign out[13] = u_rca_fa13_y2;
  assign out[14] = u_rca_fa13_y4;
endmodule

module h_s_dadda_rca8(input [7:0] a, input [7:0] b, output [15:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire constant_wire_1;
  wire h_s_dadda_rca8_and_6_0_y0;
  wire h_s_dadda_rca8_and_5_1_y0;
  wire h_s_dadda_rca8_ha0_y0;
  wire h_s_dadda_rca8_ha0_y1;
  wire h_s_dadda_rca8_nand_7_0_y0;
  wire h_s_dadda_rca8_and_6_1_y0;
  wire h_s_dadda_rca8_fa0_y2;
  wire h_s_dadda_rca8_fa0_y4;
  wire h_s_dadda_rca8_and_5_2_y0;
  wire h_s_dadda_rca8_and_4_3_y0;
  wire h_s_dadda_rca8_ha1_y0;
  wire h_s_dadda_rca8_ha1_y1;
  wire h_s_dadda_rca8_fa1_y2;
  wire h_s_dadda_rca8_fa1_y4;
  wire h_s_dadda_rca8_nand_7_1_y0;
  wire h_s_dadda_rca8_and_6_2_y0;
  wire h_s_dadda_rca8_and_5_3_y0;
  wire h_s_dadda_rca8_fa2_y2;
  wire h_s_dadda_rca8_fa2_y4;
  wire h_s_dadda_rca8_nand_7_2_y0;
  wire h_s_dadda_rca8_fa3_y2;
  wire h_s_dadda_rca8_fa3_y4;
  wire h_s_dadda_rca8_and_3_0_y0;
  wire h_s_dadda_rca8_and_2_1_y0;
  wire h_s_dadda_rca8_ha2_y0;
  wire h_s_dadda_rca8_ha2_y1;
  wire h_s_dadda_rca8_and_4_0_y0;
  wire h_s_dadda_rca8_and_3_1_y0;
  wire h_s_dadda_rca8_fa4_y2;
  wire h_s_dadda_rca8_fa4_y4;
  wire h_s_dadda_rca8_and_2_2_y0;
  wire h_s_dadda_rca8_and_1_3_y0;
  wire h_s_dadda_rca8_ha3_y0;
  wire h_s_dadda_rca8_ha3_y1;
  wire h_s_dadda_rca8_and_5_0_y0;
  wire h_s_dadda_rca8_fa5_y2;
  wire h_s_dadda_rca8_fa5_y4;
  wire h_s_dadda_rca8_and_4_1_y0;
  wire h_s_dadda_rca8_and_3_2_y0;
  wire h_s_dadda_rca8_and_2_3_y0;
  wire h_s_dadda_rca8_fa6_y2;
  wire h_s_dadda_rca8_fa6_y4;
  wire h_s_dadda_rca8_and_1_4_y0;
  wire h_s_dadda_rca8_and_0_5_y0;
  wire h_s_dadda_rca8_ha4_y0;
  wire h_s_dadda_rca8_ha4_y1;
  wire h_s_dadda_rca8_fa7_y2;
  wire h_s_dadda_rca8_fa7_y4;
  wire h_s_dadda_rca8_and_4_2_y0;
  wire h_s_dadda_rca8_and_3_3_y0;
  wire h_s_dadda_rca8_and_2_4_y0;
  wire h_s_dadda_rca8_fa8_y2;
  wire h_s_dadda_rca8_fa8_y4;
  wire h_s_dadda_rca8_and_1_5_y0;
  wire h_s_dadda_rca8_and_0_6_y0;
  wire h_s_dadda_rca8_fa9_y2;
  wire h_s_dadda_rca8_fa9_y4;
  wire h_s_dadda_rca8_fa10_y2;
  wire h_s_dadda_rca8_fa10_y4;
  wire h_s_dadda_rca8_and_3_4_y0;
  wire h_s_dadda_rca8_and_2_5_y0;
  wire h_s_dadda_rca8_and_1_6_y0;
  wire h_s_dadda_rca8_fa11_y2;
  wire h_s_dadda_rca8_fa11_y4;
  wire h_s_dadda_rca8_nand_0_7_y0;
  wire h_s_dadda_rca8_fa12_y2;
  wire h_s_dadda_rca8_fa12_y4;
  wire h_s_dadda_rca8_fa13_y2;
  wire h_s_dadda_rca8_fa13_y4;
  wire h_s_dadda_rca8_and_4_4_y0;
  wire h_s_dadda_rca8_and_3_5_y0;
  wire h_s_dadda_rca8_and_2_6_y0;
  wire h_s_dadda_rca8_fa14_y2;
  wire h_s_dadda_rca8_fa14_y4;
  wire h_s_dadda_rca8_nand_1_7_y0;
  wire h_s_dadda_rca8_fa15_y2;
  wire h_s_dadda_rca8_fa15_y4;
  wire h_s_dadda_rca8_fa16_y2;
  wire h_s_dadda_rca8_fa16_y4;
  wire h_s_dadda_rca8_and_6_3_y0;
  wire h_s_dadda_rca8_and_5_4_y0;
  wire h_s_dadda_rca8_and_4_5_y0;
  wire h_s_dadda_rca8_fa17_y2;
  wire h_s_dadda_rca8_fa17_y4;
  wire h_s_dadda_rca8_and_3_6_y0;
  wire h_s_dadda_rca8_nand_2_7_y0;
  wire h_s_dadda_rca8_fa18_y2;
  wire h_s_dadda_rca8_fa18_y4;
  wire h_s_dadda_rca8_fa19_y2;
  wire h_s_dadda_rca8_fa19_y4;
  wire h_s_dadda_rca8_nand_7_3_y0;
  wire h_s_dadda_rca8_and_6_4_y0;
  wire h_s_dadda_rca8_fa20_y2;
  wire h_s_dadda_rca8_fa20_y4;
  wire h_s_dadda_rca8_and_5_5_y0;
  wire h_s_dadda_rca8_and_4_6_y0;
  wire h_s_dadda_rca8_nand_3_7_y0;
  wire h_s_dadda_rca8_fa21_y2;
  wire h_s_dadda_rca8_fa21_y4;
  wire h_s_dadda_rca8_fa22_y2;
  wire h_s_dadda_rca8_fa22_y4;
  wire h_s_dadda_rca8_nand_7_4_y0;
  wire h_s_dadda_rca8_and_6_5_y0;
  wire h_s_dadda_rca8_and_5_6_y0;
  wire h_s_dadda_rca8_fa23_y2;
  wire h_s_dadda_rca8_fa23_y4;
  wire h_s_dadda_rca8_nand_7_5_y0;
  wire h_s_dadda_rca8_fa24_y2;
  wire h_s_dadda_rca8_fa24_y4;
  wire h_s_dadda_rca8_and_2_0_y0;
  wire h_s_dadda_rca8_and_1_1_y0;
  wire h_s_dadda_rca8_ha5_y0;
  wire h_s_dadda_rca8_ha5_y1;
  wire h_s_dadda_rca8_and_1_2_y0;
  wire h_s_dadda_rca8_and_0_3_y0;
  wire h_s_dadda_rca8_fa25_y2;
  wire h_s_dadda_rca8_fa25_y4;
  wire h_s_dadda_rca8_and_0_4_y0;
  wire h_s_dadda_rca8_fa26_y2;
  wire h_s_dadda_rca8_fa26_y4;
  wire h_s_dadda_rca8_fa27_y2;
  wire h_s_dadda_rca8_fa27_y4;
  wire h_s_dadda_rca8_fa28_y2;
  wire h_s_dadda_rca8_fa28_y4;
  wire h_s_dadda_rca8_fa29_y2;
  wire h_s_dadda_rca8_fa29_y4;
  wire h_s_dadda_rca8_fa30_y2;
  wire h_s_dadda_rca8_fa30_y4;
  wire h_s_dadda_rca8_fa31_y2;
  wire h_s_dadda_rca8_fa31_y4;
  wire h_s_dadda_rca8_fa32_y2;
  wire h_s_dadda_rca8_fa32_y4;
  wire h_s_dadda_rca8_nand_4_7_y0;
  wire h_s_dadda_rca8_fa33_y2;
  wire h_s_dadda_rca8_fa33_y4;
  wire h_s_dadda_rca8_and_6_6_y0;
  wire h_s_dadda_rca8_nand_5_7_y0;
  wire h_s_dadda_rca8_fa34_y2;
  wire h_s_dadda_rca8_fa34_y4;
  wire h_s_dadda_rca8_nand_7_6_y0;
  wire h_s_dadda_rca8_fa35_y2;
  wire h_s_dadda_rca8_fa35_y4;
  wire h_s_dadda_rca8_and_0_0_y0;
  wire h_s_dadda_rca8_and_1_0_y0;
  wire h_s_dadda_rca8_and_0_2_y0;
  wire h_s_dadda_rca8_nand_6_7_y0;
  wire h_s_dadda_rca8_and_0_1_y0;
  wire h_s_dadda_rca8_and_7_7_y0;
  wire [13:0] h_s_dadda_rca8_u_rca_u_rca_a;
  wire [13:0] h_s_dadda_rca8_u_rca_u_rca_b;
  wire [14:0] h_s_dadda_rca8_u_rca_out;
  wire h_s_dadda_rca8_u_rca_ha_y0;
  wire h_s_dadda_rca8_u_rca_fa1_y2;
  wire h_s_dadda_rca8_u_rca_fa2_y2;
  wire h_s_dadda_rca8_u_rca_fa3_y2;
  wire h_s_dadda_rca8_u_rca_fa4_y2;
  wire h_s_dadda_rca8_u_rca_fa5_y2;
  wire h_s_dadda_rca8_u_rca_fa6_y2;
  wire h_s_dadda_rca8_u_rca_fa7_y2;
  wire h_s_dadda_rca8_u_rca_fa8_y2;
  wire h_s_dadda_rca8_u_rca_fa9_y2;
  wire h_s_dadda_rca8_u_rca_fa10_y2;
  wire h_s_dadda_rca8_u_rca_fa11_y2;
  wire h_s_dadda_rca8_u_rca_fa12_y2;
  wire h_s_dadda_rca8_u_rca_fa13_y2;
  wire h_s_dadda_rca8_u_rca_fa13_y4;
  wire h_s_dadda_rca8_xor0_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  constant_wire_value_1 constant_wire_value_1_constant_wire_1(a_0, b_0, constant_wire_1);
  and_gate and_gate_h_s_dadda_rca8_and_6_0_y0(a_6, b_0, h_s_dadda_rca8_and_6_0_y0);
  and_gate and_gate_h_s_dadda_rca8_and_5_1_y0(a_5, b_1, h_s_dadda_rca8_and_5_1_y0);
  ha ha_h_s_dadda_rca8_ha0_y0(h_s_dadda_rca8_and_6_0_y0, h_s_dadda_rca8_and_5_1_y0, h_s_dadda_rca8_ha0_y0, h_s_dadda_rca8_ha0_y1);
  nand_gate nand_gate_h_s_dadda_rca8_nand_7_0_y0(a_7, b_0, h_s_dadda_rca8_nand_7_0_y0);
  and_gate and_gate_h_s_dadda_rca8_and_6_1_y0(a_6, b_1, h_s_dadda_rca8_and_6_1_y0);
  fa fa_h_s_dadda_rca8_fa0_y2(h_s_dadda_rca8_ha0_y1, h_s_dadda_rca8_nand_7_0_y0, h_s_dadda_rca8_and_6_1_y0, h_s_dadda_rca8_fa0_y2, h_s_dadda_rca8_fa0_y4);
  and_gate and_gate_h_s_dadda_rca8_and_5_2_y0(a_5, b_2, h_s_dadda_rca8_and_5_2_y0);
  and_gate and_gate_h_s_dadda_rca8_and_4_3_y0(a_4, b_3, h_s_dadda_rca8_and_4_3_y0);
  ha ha_h_s_dadda_rca8_ha1_y0(h_s_dadda_rca8_and_5_2_y0, h_s_dadda_rca8_and_4_3_y0, h_s_dadda_rca8_ha1_y0, h_s_dadda_rca8_ha1_y1);
  fa fa_h_s_dadda_rca8_fa1_y2(h_s_dadda_rca8_ha1_y1, h_s_dadda_rca8_fa0_y4, constant_wire_1, h_s_dadda_rca8_fa1_y2, h_s_dadda_rca8_fa1_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_7_1_y0(a_7, b_1, h_s_dadda_rca8_nand_7_1_y0);
  and_gate and_gate_h_s_dadda_rca8_and_6_2_y0(a_6, b_2, h_s_dadda_rca8_and_6_2_y0);
  and_gate and_gate_h_s_dadda_rca8_and_5_3_y0(a_5, b_3, h_s_dadda_rca8_and_5_3_y0);
  fa fa_h_s_dadda_rca8_fa2_y2(h_s_dadda_rca8_nand_7_1_y0, h_s_dadda_rca8_and_6_2_y0, h_s_dadda_rca8_and_5_3_y0, h_s_dadda_rca8_fa2_y2, h_s_dadda_rca8_fa2_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_7_2_y0(a_7, b_2, h_s_dadda_rca8_nand_7_2_y0);
  fa fa_h_s_dadda_rca8_fa3_y2(h_s_dadda_rca8_fa2_y4, h_s_dadda_rca8_fa1_y4, h_s_dadda_rca8_nand_7_2_y0, h_s_dadda_rca8_fa3_y2, h_s_dadda_rca8_fa3_y4);
  and_gate and_gate_h_s_dadda_rca8_and_3_0_y0(a_3, b_0, h_s_dadda_rca8_and_3_0_y0);
  and_gate and_gate_h_s_dadda_rca8_and_2_1_y0(a_2, b_1, h_s_dadda_rca8_and_2_1_y0);
  ha ha_h_s_dadda_rca8_ha2_y0(h_s_dadda_rca8_and_3_0_y0, h_s_dadda_rca8_and_2_1_y0, h_s_dadda_rca8_ha2_y0, h_s_dadda_rca8_ha2_y1);
  and_gate and_gate_h_s_dadda_rca8_and_4_0_y0(a_4, b_0, h_s_dadda_rca8_and_4_0_y0);
  and_gate and_gate_h_s_dadda_rca8_and_3_1_y0(a_3, b_1, h_s_dadda_rca8_and_3_1_y0);
  fa fa_h_s_dadda_rca8_fa4_y2(h_s_dadda_rca8_ha2_y1, h_s_dadda_rca8_and_4_0_y0, h_s_dadda_rca8_and_3_1_y0, h_s_dadda_rca8_fa4_y2, h_s_dadda_rca8_fa4_y4);
  and_gate and_gate_h_s_dadda_rca8_and_2_2_y0(a_2, b_2, h_s_dadda_rca8_and_2_2_y0);
  and_gate and_gate_h_s_dadda_rca8_and_1_3_y0(a_1, b_3, h_s_dadda_rca8_and_1_3_y0);
  ha ha_h_s_dadda_rca8_ha3_y0(h_s_dadda_rca8_and_2_2_y0, h_s_dadda_rca8_and_1_3_y0, h_s_dadda_rca8_ha3_y0, h_s_dadda_rca8_ha3_y1);
  and_gate and_gate_h_s_dadda_rca8_and_5_0_y0(a_5, b_0, h_s_dadda_rca8_and_5_0_y0);
  fa fa_h_s_dadda_rca8_fa5_y2(h_s_dadda_rca8_ha3_y1, h_s_dadda_rca8_fa4_y4, h_s_dadda_rca8_and_5_0_y0, h_s_dadda_rca8_fa5_y2, h_s_dadda_rca8_fa5_y4);
  and_gate and_gate_h_s_dadda_rca8_and_4_1_y0(a_4, b_1, h_s_dadda_rca8_and_4_1_y0);
  and_gate and_gate_h_s_dadda_rca8_and_3_2_y0(a_3, b_2, h_s_dadda_rca8_and_3_2_y0);
  and_gate and_gate_h_s_dadda_rca8_and_2_3_y0(a_2, b_3, h_s_dadda_rca8_and_2_3_y0);
  fa fa_h_s_dadda_rca8_fa6_y2(h_s_dadda_rca8_and_4_1_y0, h_s_dadda_rca8_and_3_2_y0, h_s_dadda_rca8_and_2_3_y0, h_s_dadda_rca8_fa6_y2, h_s_dadda_rca8_fa6_y4);
  and_gate and_gate_h_s_dadda_rca8_and_1_4_y0(a_1, b_4, h_s_dadda_rca8_and_1_4_y0);
  and_gate and_gate_h_s_dadda_rca8_and_0_5_y0(a_0, b_5, h_s_dadda_rca8_and_0_5_y0);
  ha ha_h_s_dadda_rca8_ha4_y0(h_s_dadda_rca8_and_1_4_y0, h_s_dadda_rca8_and_0_5_y0, h_s_dadda_rca8_ha4_y0, h_s_dadda_rca8_ha4_y1);
  fa fa_h_s_dadda_rca8_fa7_y2(h_s_dadda_rca8_ha4_y1, h_s_dadda_rca8_fa6_y4, h_s_dadda_rca8_fa5_y4, h_s_dadda_rca8_fa7_y2, h_s_dadda_rca8_fa7_y4);
  and_gate and_gate_h_s_dadda_rca8_and_4_2_y0(a_4, b_2, h_s_dadda_rca8_and_4_2_y0);
  and_gate and_gate_h_s_dadda_rca8_and_3_3_y0(a_3, b_3, h_s_dadda_rca8_and_3_3_y0);
  and_gate and_gate_h_s_dadda_rca8_and_2_4_y0(a_2, b_4, h_s_dadda_rca8_and_2_4_y0);
  fa fa_h_s_dadda_rca8_fa8_y2(h_s_dadda_rca8_and_4_2_y0, h_s_dadda_rca8_and_3_3_y0, h_s_dadda_rca8_and_2_4_y0, h_s_dadda_rca8_fa8_y2, h_s_dadda_rca8_fa8_y4);
  and_gate and_gate_h_s_dadda_rca8_and_1_5_y0(a_1, b_5, h_s_dadda_rca8_and_1_5_y0);
  and_gate and_gate_h_s_dadda_rca8_and_0_6_y0(a_0, b_6, h_s_dadda_rca8_and_0_6_y0);
  fa fa_h_s_dadda_rca8_fa9_y2(h_s_dadda_rca8_and_1_5_y0, h_s_dadda_rca8_and_0_6_y0, h_s_dadda_rca8_ha0_y0, h_s_dadda_rca8_fa9_y2, h_s_dadda_rca8_fa9_y4);
  fa fa_h_s_dadda_rca8_fa10_y2(h_s_dadda_rca8_fa9_y4, h_s_dadda_rca8_fa8_y4, h_s_dadda_rca8_fa7_y4, h_s_dadda_rca8_fa10_y2, h_s_dadda_rca8_fa10_y4);
  and_gate and_gate_h_s_dadda_rca8_and_3_4_y0(a_3, b_4, h_s_dadda_rca8_and_3_4_y0);
  and_gate and_gate_h_s_dadda_rca8_and_2_5_y0(a_2, b_5, h_s_dadda_rca8_and_2_5_y0);
  and_gate and_gate_h_s_dadda_rca8_and_1_6_y0(a_1, b_6, h_s_dadda_rca8_and_1_6_y0);
  fa fa_h_s_dadda_rca8_fa11_y2(h_s_dadda_rca8_and_3_4_y0, h_s_dadda_rca8_and_2_5_y0, h_s_dadda_rca8_and_1_6_y0, h_s_dadda_rca8_fa11_y2, h_s_dadda_rca8_fa11_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_0_7_y0(a_0, b_7, h_s_dadda_rca8_nand_0_7_y0);
  fa fa_h_s_dadda_rca8_fa12_y2(h_s_dadda_rca8_nand_0_7_y0, h_s_dadda_rca8_fa0_y2, h_s_dadda_rca8_ha1_y0, h_s_dadda_rca8_fa12_y2, h_s_dadda_rca8_fa12_y4);
  fa fa_h_s_dadda_rca8_fa13_y2(h_s_dadda_rca8_fa12_y4, h_s_dadda_rca8_fa11_y4, h_s_dadda_rca8_fa10_y4, h_s_dadda_rca8_fa13_y2, h_s_dadda_rca8_fa13_y4);
  and_gate and_gate_h_s_dadda_rca8_and_4_4_y0(a_4, b_4, h_s_dadda_rca8_and_4_4_y0);
  and_gate and_gate_h_s_dadda_rca8_and_3_5_y0(a_3, b_5, h_s_dadda_rca8_and_3_5_y0);
  and_gate and_gate_h_s_dadda_rca8_and_2_6_y0(a_2, b_6, h_s_dadda_rca8_and_2_6_y0);
  fa fa_h_s_dadda_rca8_fa14_y2(h_s_dadda_rca8_and_4_4_y0, h_s_dadda_rca8_and_3_5_y0, h_s_dadda_rca8_and_2_6_y0, h_s_dadda_rca8_fa14_y2, h_s_dadda_rca8_fa14_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_1_7_y0(a_1, b_7, h_s_dadda_rca8_nand_1_7_y0);
  fa fa_h_s_dadda_rca8_fa15_y2(h_s_dadda_rca8_nand_1_7_y0, h_s_dadda_rca8_fa1_y2, h_s_dadda_rca8_fa2_y2, h_s_dadda_rca8_fa15_y2, h_s_dadda_rca8_fa15_y4);
  fa fa_h_s_dadda_rca8_fa16_y2(h_s_dadda_rca8_fa15_y4, h_s_dadda_rca8_fa14_y4, h_s_dadda_rca8_fa13_y4, h_s_dadda_rca8_fa16_y2, h_s_dadda_rca8_fa16_y4);
  and_gate and_gate_h_s_dadda_rca8_and_6_3_y0(a_6, b_3, h_s_dadda_rca8_and_6_3_y0);
  and_gate and_gate_h_s_dadda_rca8_and_5_4_y0(a_5, b_4, h_s_dadda_rca8_and_5_4_y0);
  and_gate and_gate_h_s_dadda_rca8_and_4_5_y0(a_4, b_5, h_s_dadda_rca8_and_4_5_y0);
  fa fa_h_s_dadda_rca8_fa17_y2(h_s_dadda_rca8_and_6_3_y0, h_s_dadda_rca8_and_5_4_y0, h_s_dadda_rca8_and_4_5_y0, h_s_dadda_rca8_fa17_y2, h_s_dadda_rca8_fa17_y4);
  and_gate and_gate_h_s_dadda_rca8_and_3_6_y0(a_3, b_6, h_s_dadda_rca8_and_3_6_y0);
  nand_gate nand_gate_h_s_dadda_rca8_nand_2_7_y0(a_2, b_7, h_s_dadda_rca8_nand_2_7_y0);
  fa fa_h_s_dadda_rca8_fa18_y2(h_s_dadda_rca8_and_3_6_y0, h_s_dadda_rca8_nand_2_7_y0, h_s_dadda_rca8_fa3_y2, h_s_dadda_rca8_fa18_y2, h_s_dadda_rca8_fa18_y4);
  fa fa_h_s_dadda_rca8_fa19_y2(h_s_dadda_rca8_fa18_y4, h_s_dadda_rca8_fa17_y4, h_s_dadda_rca8_fa16_y4, h_s_dadda_rca8_fa19_y2, h_s_dadda_rca8_fa19_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_7_3_y0(a_7, b_3, h_s_dadda_rca8_nand_7_3_y0);
  and_gate and_gate_h_s_dadda_rca8_and_6_4_y0(a_6, b_4, h_s_dadda_rca8_and_6_4_y0);
  fa fa_h_s_dadda_rca8_fa20_y2(h_s_dadda_rca8_fa3_y4, h_s_dadda_rca8_nand_7_3_y0, h_s_dadda_rca8_and_6_4_y0, h_s_dadda_rca8_fa20_y2, h_s_dadda_rca8_fa20_y4);
  and_gate and_gate_h_s_dadda_rca8_and_5_5_y0(a_5, b_5, h_s_dadda_rca8_and_5_5_y0);
  and_gate and_gate_h_s_dadda_rca8_and_4_6_y0(a_4, b_6, h_s_dadda_rca8_and_4_6_y0);
  nand_gate nand_gate_h_s_dadda_rca8_nand_3_7_y0(a_3, b_7, h_s_dadda_rca8_nand_3_7_y0);
  fa fa_h_s_dadda_rca8_fa21_y2(h_s_dadda_rca8_and_5_5_y0, h_s_dadda_rca8_and_4_6_y0, h_s_dadda_rca8_nand_3_7_y0, h_s_dadda_rca8_fa21_y2, h_s_dadda_rca8_fa21_y4);
  fa fa_h_s_dadda_rca8_fa22_y2(h_s_dadda_rca8_fa21_y4, h_s_dadda_rca8_fa20_y4, h_s_dadda_rca8_fa19_y4, h_s_dadda_rca8_fa22_y2, h_s_dadda_rca8_fa22_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_7_4_y0(a_7, b_4, h_s_dadda_rca8_nand_7_4_y0);
  and_gate and_gate_h_s_dadda_rca8_and_6_5_y0(a_6, b_5, h_s_dadda_rca8_and_6_5_y0);
  and_gate and_gate_h_s_dadda_rca8_and_5_6_y0(a_5, b_6, h_s_dadda_rca8_and_5_6_y0);
  fa fa_h_s_dadda_rca8_fa23_y2(h_s_dadda_rca8_nand_7_4_y0, h_s_dadda_rca8_and_6_5_y0, h_s_dadda_rca8_and_5_6_y0, h_s_dadda_rca8_fa23_y2, h_s_dadda_rca8_fa23_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_7_5_y0(a_7, b_5, h_s_dadda_rca8_nand_7_5_y0);
  fa fa_h_s_dadda_rca8_fa24_y2(h_s_dadda_rca8_fa23_y4, h_s_dadda_rca8_fa22_y4, h_s_dadda_rca8_nand_7_5_y0, h_s_dadda_rca8_fa24_y2, h_s_dadda_rca8_fa24_y4);
  and_gate and_gate_h_s_dadda_rca8_and_2_0_y0(a_2, b_0, h_s_dadda_rca8_and_2_0_y0);
  and_gate and_gate_h_s_dadda_rca8_and_1_1_y0(a_1, b_1, h_s_dadda_rca8_and_1_1_y0);
  ha ha_h_s_dadda_rca8_ha5_y0(h_s_dadda_rca8_and_2_0_y0, h_s_dadda_rca8_and_1_1_y0, h_s_dadda_rca8_ha5_y0, h_s_dadda_rca8_ha5_y1);
  and_gate and_gate_h_s_dadda_rca8_and_1_2_y0(a_1, b_2, h_s_dadda_rca8_and_1_2_y0);
  and_gate and_gate_h_s_dadda_rca8_and_0_3_y0(a_0, b_3, h_s_dadda_rca8_and_0_3_y0);
  fa fa_h_s_dadda_rca8_fa25_y2(h_s_dadda_rca8_ha5_y1, h_s_dadda_rca8_and_1_2_y0, h_s_dadda_rca8_and_0_3_y0, h_s_dadda_rca8_fa25_y2, h_s_dadda_rca8_fa25_y4);
  and_gate and_gate_h_s_dadda_rca8_and_0_4_y0(a_0, b_4, h_s_dadda_rca8_and_0_4_y0);
  fa fa_h_s_dadda_rca8_fa26_y2(h_s_dadda_rca8_fa25_y4, h_s_dadda_rca8_and_0_4_y0, h_s_dadda_rca8_fa4_y2, h_s_dadda_rca8_fa26_y2, h_s_dadda_rca8_fa26_y4);
  fa fa_h_s_dadda_rca8_fa27_y2(h_s_dadda_rca8_fa26_y4, h_s_dadda_rca8_fa5_y2, h_s_dadda_rca8_fa6_y2, h_s_dadda_rca8_fa27_y2, h_s_dadda_rca8_fa27_y4);
  fa fa_h_s_dadda_rca8_fa28_y2(h_s_dadda_rca8_fa27_y4, h_s_dadda_rca8_fa7_y2, h_s_dadda_rca8_fa8_y2, h_s_dadda_rca8_fa28_y2, h_s_dadda_rca8_fa28_y4);
  fa fa_h_s_dadda_rca8_fa29_y2(h_s_dadda_rca8_fa28_y4, h_s_dadda_rca8_fa10_y2, h_s_dadda_rca8_fa11_y2, h_s_dadda_rca8_fa29_y2, h_s_dadda_rca8_fa29_y4);
  fa fa_h_s_dadda_rca8_fa30_y2(h_s_dadda_rca8_fa29_y4, h_s_dadda_rca8_fa13_y2, h_s_dadda_rca8_fa14_y2, h_s_dadda_rca8_fa30_y2, h_s_dadda_rca8_fa30_y4);
  fa fa_h_s_dadda_rca8_fa31_y2(h_s_dadda_rca8_fa30_y4, h_s_dadda_rca8_fa16_y2, h_s_dadda_rca8_fa17_y2, h_s_dadda_rca8_fa31_y2, h_s_dadda_rca8_fa31_y4);
  fa fa_h_s_dadda_rca8_fa32_y2(h_s_dadda_rca8_fa31_y4, h_s_dadda_rca8_fa19_y2, h_s_dadda_rca8_fa20_y2, h_s_dadda_rca8_fa32_y2, h_s_dadda_rca8_fa32_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_4_7_y0(a_4, b_7, h_s_dadda_rca8_nand_4_7_y0);
  fa fa_h_s_dadda_rca8_fa33_y2(h_s_dadda_rca8_fa32_y4, h_s_dadda_rca8_nand_4_7_y0, h_s_dadda_rca8_fa22_y2, h_s_dadda_rca8_fa33_y2, h_s_dadda_rca8_fa33_y4);
  and_gate and_gate_h_s_dadda_rca8_and_6_6_y0(a_6, b_6, h_s_dadda_rca8_and_6_6_y0);
  nand_gate nand_gate_h_s_dadda_rca8_nand_5_7_y0(a_5, b_7, h_s_dadda_rca8_nand_5_7_y0);
  fa fa_h_s_dadda_rca8_fa34_y2(h_s_dadda_rca8_fa33_y4, h_s_dadda_rca8_and_6_6_y0, h_s_dadda_rca8_nand_5_7_y0, h_s_dadda_rca8_fa34_y2, h_s_dadda_rca8_fa34_y4);
  nand_gate nand_gate_h_s_dadda_rca8_nand_7_6_y0(a_7, b_6, h_s_dadda_rca8_nand_7_6_y0);
  fa fa_h_s_dadda_rca8_fa35_y2(h_s_dadda_rca8_fa34_y4, h_s_dadda_rca8_fa24_y4, h_s_dadda_rca8_nand_7_6_y0, h_s_dadda_rca8_fa35_y2, h_s_dadda_rca8_fa35_y4);
  and_gate and_gate_h_s_dadda_rca8_and_0_0_y0(a_0, b_0, h_s_dadda_rca8_and_0_0_y0);
  and_gate and_gate_h_s_dadda_rca8_and_1_0_y0(a_1, b_0, h_s_dadda_rca8_and_1_0_y0);
  and_gate and_gate_h_s_dadda_rca8_and_0_2_y0(a_0, b_2, h_s_dadda_rca8_and_0_2_y0);
  nand_gate nand_gate_h_s_dadda_rca8_nand_6_7_y0(a_6, b_7, h_s_dadda_rca8_nand_6_7_y0);
  and_gate and_gate_h_s_dadda_rca8_and_0_1_y0(a_0, b_1, h_s_dadda_rca8_and_0_1_y0);
  and_gate and_gate_h_s_dadda_rca8_and_7_7_y0(a_7, b_7, h_s_dadda_rca8_and_7_7_y0);
  assign h_s_dadda_rca8_u_rca_u_rca_a[0] = h_s_dadda_rca8_and_1_0_y0;
  assign h_s_dadda_rca8_u_rca_u_rca_a[1] = h_s_dadda_rca8_and_0_2_y0;
  assign h_s_dadda_rca8_u_rca_u_rca_a[2] = h_s_dadda_rca8_ha2_y0;
  assign h_s_dadda_rca8_u_rca_u_rca_a[3] = h_s_dadda_rca8_ha3_y0;
  assign h_s_dadda_rca8_u_rca_u_rca_a[4] = h_s_dadda_rca8_ha4_y0;
  assign h_s_dadda_rca8_u_rca_u_rca_a[5] = h_s_dadda_rca8_fa9_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_a[6] = h_s_dadda_rca8_fa12_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_a[7] = h_s_dadda_rca8_fa15_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_a[8] = h_s_dadda_rca8_fa18_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_a[9] = h_s_dadda_rca8_fa21_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_a[10] = h_s_dadda_rca8_fa23_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_a[11] = h_s_dadda_rca8_fa24_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_a[12] = h_s_dadda_rca8_nand_6_7_y0;
  assign h_s_dadda_rca8_u_rca_u_rca_a[13] = h_s_dadda_rca8_fa35_y4;
  assign h_s_dadda_rca8_u_rca_u_rca_b[0] = h_s_dadda_rca8_and_0_1_y0;
  assign h_s_dadda_rca8_u_rca_u_rca_b[1] = h_s_dadda_rca8_ha5_y0;
  assign h_s_dadda_rca8_u_rca_u_rca_b[2] = h_s_dadda_rca8_fa25_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[3] = h_s_dadda_rca8_fa26_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[4] = h_s_dadda_rca8_fa27_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[5] = h_s_dadda_rca8_fa28_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[6] = h_s_dadda_rca8_fa29_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[7] = h_s_dadda_rca8_fa30_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[8] = h_s_dadda_rca8_fa31_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[9] = h_s_dadda_rca8_fa32_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[10] = h_s_dadda_rca8_fa33_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[11] = h_s_dadda_rca8_fa34_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[12] = h_s_dadda_rca8_fa35_y2;
  assign h_s_dadda_rca8_u_rca_u_rca_b[13] = h_s_dadda_rca8_and_7_7_y0;
  u_rca u_rca_out(h_s_dadda_rca8_u_rca_u_rca_a, h_s_dadda_rca8_u_rca_u_rca_b, h_s_dadda_rca8_u_rca_out);
  assign h_s_dadda_rca8_u_rca_ha_y0 = h_s_dadda_rca8_u_rca_out[0];
  assign h_s_dadda_rca8_u_rca_fa1_y2 = h_s_dadda_rca8_u_rca_out[1];
  assign h_s_dadda_rca8_u_rca_fa2_y2 = h_s_dadda_rca8_u_rca_out[2];
  assign h_s_dadda_rca8_u_rca_fa3_y2 = h_s_dadda_rca8_u_rca_out[3];
  assign h_s_dadda_rca8_u_rca_fa4_y2 = h_s_dadda_rca8_u_rca_out[4];
  assign h_s_dadda_rca8_u_rca_fa5_y2 = h_s_dadda_rca8_u_rca_out[5];
  assign h_s_dadda_rca8_u_rca_fa6_y2 = h_s_dadda_rca8_u_rca_out[6];
  assign h_s_dadda_rca8_u_rca_fa7_y2 = h_s_dadda_rca8_u_rca_out[7];
  assign h_s_dadda_rca8_u_rca_fa8_y2 = h_s_dadda_rca8_u_rca_out[8];
  assign h_s_dadda_rca8_u_rca_fa9_y2 = h_s_dadda_rca8_u_rca_out[9];
  assign h_s_dadda_rca8_u_rca_fa10_y2 = h_s_dadda_rca8_u_rca_out[10];
  assign h_s_dadda_rca8_u_rca_fa11_y2 = h_s_dadda_rca8_u_rca_out[11];
  assign h_s_dadda_rca8_u_rca_fa12_y2 = h_s_dadda_rca8_u_rca_out[12];
  assign h_s_dadda_rca8_u_rca_fa13_y2 = h_s_dadda_rca8_u_rca_out[13];
  assign h_s_dadda_rca8_u_rca_fa13_y4 = h_s_dadda_rca8_u_rca_out[14];
  xor_gate xor_gate_h_s_dadda_rca8_xor0_y0(constant_wire_1, h_s_dadda_rca8_u_rca_fa13_y4, h_s_dadda_rca8_xor0_y0);

  assign out[0] = h_s_dadda_rca8_and_0_0_y0;
  assign out[1] = h_s_dadda_rca8_u_rca_ha_y0;
  assign out[2] = h_s_dadda_rca8_u_rca_fa1_y2;
  assign out[3] = h_s_dadda_rca8_u_rca_fa2_y2;
  assign out[4] = h_s_dadda_rca8_u_rca_fa3_y2;
  assign out[5] = h_s_dadda_rca8_u_rca_fa4_y2;
  assign out[6] = h_s_dadda_rca8_u_rca_fa5_y2;
  assign out[7] = h_s_dadda_rca8_u_rca_fa6_y2;
  assign out[8] = h_s_dadda_rca8_u_rca_fa7_y2;
  assign out[9] = h_s_dadda_rca8_u_rca_fa8_y2;
  assign out[10] = h_s_dadda_rca8_u_rca_fa9_y2;
  assign out[11] = h_s_dadda_rca8_u_rca_fa10_y2;
  assign out[12] = h_s_dadda_rca8_u_rca_fa11_y2;
  assign out[13] = h_s_dadda_rca8_u_rca_fa12_y2;
  assign out[14] = h_s_dadda_rca8_u_rca_fa13_y2;
  assign out[15] = h_s_dadda_rca8_xor0_y0;
endmodule