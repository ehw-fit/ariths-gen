module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module nand_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a & _b);
endmodule

module nor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a | _b);
endmodule

module constant_wire_value_1(input a, input b, output constant_wire_1);
  wire constant_wire_value_1_a;
  wire constant_wire_value_1_b;

  assign constant_wire_value_1_a = a;
  assign constant_wire_value_1_b = b;

  xor_gate xor_gate_constant_wire_value_1_y0(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y0);
  xnor_gate xnor_gate_constant_wire_value_1_y1(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y1);
  or_gate or_gate_constant_wire_1(constant_wire_value_1_y0, constant_wire_value_1_y1, constant_wire_1);
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_cin;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module constant_wire_value_0(input a, input b, output constant_wire_0);
  wire constant_wire_value_0_a;
  wire constant_wire_value_0_b;

  assign constant_wire_value_0_a = a;
  assign constant_wire_value_0_b = b;

  xor_gate xor_gate_constant_wire_value_0_y0(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y0);
  xnor_gate xnor_gate_constant_wire_value_0_y1(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y1);
  nor_gate nor_gate_constant_wire_0(constant_wire_value_0_y0, constant_wire_value_0_y1, constant_wire_0);
endmodule

module fa_cla(input a, input b, input cin, output fa_cla_y0, output fa_cla_y1, output fa_cla_y2);
  wire fa_cla_a;
  wire fa_cla_b;
  wire fa_cla_cin;

  assign fa_cla_a = a;
  assign fa_cla_b = b;
  assign fa_cla_cin = cin;

  xor_gate xor_gate_fa_cla_y0(fa_cla_a, fa_cla_b, fa_cla_y0);
  and_gate and_gate_fa_cla_y1(fa_cla_a, fa_cla_b, fa_cla_y1);
  xor_gate xor_gate_fa_cla_y2(fa_cla_y0, fa_cla_cin, fa_cla_y2);
endmodule

module u_pg_rca(input [21:0] a, input [21:0] b, output [22:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire constant_wire_0;
  wire u_pg_rca_fa0_y0;
  wire u_pg_rca_fa0_y1;
  wire u_pg_rca_fa0_y2;
  wire u_pg_rca_and0_y0;
  wire u_pg_rca_or0_y0;
  wire u_pg_rca_fa1_y0;
  wire u_pg_rca_fa1_y1;
  wire u_pg_rca_fa1_y2;
  wire u_pg_rca_and1_y0;
  wire u_pg_rca_or1_y0;
  wire u_pg_rca_fa2_y0;
  wire u_pg_rca_fa2_y1;
  wire u_pg_rca_fa2_y2;
  wire u_pg_rca_and2_y0;
  wire u_pg_rca_or2_y0;
  wire u_pg_rca_fa3_y0;
  wire u_pg_rca_fa3_y1;
  wire u_pg_rca_fa3_y2;
  wire u_pg_rca_and3_y0;
  wire u_pg_rca_or3_y0;
  wire u_pg_rca_fa4_y0;
  wire u_pg_rca_fa4_y1;
  wire u_pg_rca_fa4_y2;
  wire u_pg_rca_and4_y0;
  wire u_pg_rca_or4_y0;
  wire u_pg_rca_fa5_y0;
  wire u_pg_rca_fa5_y1;
  wire u_pg_rca_fa5_y2;
  wire u_pg_rca_and5_y0;
  wire u_pg_rca_or5_y0;
  wire u_pg_rca_fa6_y0;
  wire u_pg_rca_fa6_y1;
  wire u_pg_rca_fa6_y2;
  wire u_pg_rca_and6_y0;
  wire u_pg_rca_or6_y0;
  wire u_pg_rca_fa7_y0;
  wire u_pg_rca_fa7_y1;
  wire u_pg_rca_fa7_y2;
  wire u_pg_rca_and7_y0;
  wire u_pg_rca_or7_y0;
  wire u_pg_rca_fa8_y0;
  wire u_pg_rca_fa8_y1;
  wire u_pg_rca_fa8_y2;
  wire u_pg_rca_and8_y0;
  wire u_pg_rca_or8_y0;
  wire u_pg_rca_fa9_y0;
  wire u_pg_rca_fa9_y1;
  wire u_pg_rca_fa9_y2;
  wire u_pg_rca_and9_y0;
  wire u_pg_rca_or9_y0;
  wire u_pg_rca_fa10_y0;
  wire u_pg_rca_fa10_y1;
  wire u_pg_rca_fa10_y2;
  wire u_pg_rca_and10_y0;
  wire u_pg_rca_or10_y0;
  wire u_pg_rca_fa11_y0;
  wire u_pg_rca_fa11_y1;
  wire u_pg_rca_fa11_y2;
  wire u_pg_rca_and11_y0;
  wire u_pg_rca_or11_y0;
  wire u_pg_rca_fa12_y0;
  wire u_pg_rca_fa12_y1;
  wire u_pg_rca_fa12_y2;
  wire u_pg_rca_and12_y0;
  wire u_pg_rca_or12_y0;
  wire u_pg_rca_fa13_y0;
  wire u_pg_rca_fa13_y1;
  wire u_pg_rca_fa13_y2;
  wire u_pg_rca_and13_y0;
  wire u_pg_rca_or13_y0;
  wire u_pg_rca_fa14_y0;
  wire u_pg_rca_fa14_y1;
  wire u_pg_rca_fa14_y2;
  wire u_pg_rca_and14_y0;
  wire u_pg_rca_or14_y0;
  wire u_pg_rca_fa15_y0;
  wire u_pg_rca_fa15_y1;
  wire u_pg_rca_fa15_y2;
  wire u_pg_rca_and15_y0;
  wire u_pg_rca_or15_y0;
  wire u_pg_rca_fa16_y0;
  wire u_pg_rca_fa16_y1;
  wire u_pg_rca_fa16_y2;
  wire u_pg_rca_and16_y0;
  wire u_pg_rca_or16_y0;
  wire u_pg_rca_fa17_y0;
  wire u_pg_rca_fa17_y1;
  wire u_pg_rca_fa17_y2;
  wire u_pg_rca_and17_y0;
  wire u_pg_rca_or17_y0;
  wire u_pg_rca_fa18_y0;
  wire u_pg_rca_fa18_y1;
  wire u_pg_rca_fa18_y2;
  wire u_pg_rca_and18_y0;
  wire u_pg_rca_or18_y0;
  wire u_pg_rca_fa19_y0;
  wire u_pg_rca_fa19_y1;
  wire u_pg_rca_fa19_y2;
  wire u_pg_rca_and19_y0;
  wire u_pg_rca_or19_y0;
  wire u_pg_rca_fa20_y0;
  wire u_pg_rca_fa20_y1;
  wire u_pg_rca_fa20_y2;
  wire u_pg_rca_and20_y0;
  wire u_pg_rca_or20_y0;
  wire u_pg_rca_fa21_y0;
  wire u_pg_rca_fa21_y1;
  wire u_pg_rca_fa21_y2;
  wire u_pg_rca_and21_y0;
  wire u_pg_rca_or21_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  constant_wire_value_0 constant_wire_value_0_constant_wire_0(a_0, b_0, constant_wire_0);
  fa_cla fa_cla_u_pg_rca_fa0_y0(a_0, b_0, constant_wire_0, u_pg_rca_fa0_y0, u_pg_rca_fa0_y1, u_pg_rca_fa0_y2);
  and_gate and_gate_u_pg_rca_and0_y0(constant_wire_0, u_pg_rca_fa0_y0, u_pg_rca_and0_y0);
  or_gate or_gate_u_pg_rca_or0_y0(u_pg_rca_and0_y0, u_pg_rca_fa0_y1, u_pg_rca_or0_y0);
  fa_cla fa_cla_u_pg_rca_fa1_y0(a_1, b_1, u_pg_rca_or0_y0, u_pg_rca_fa1_y0, u_pg_rca_fa1_y1, u_pg_rca_fa1_y2);
  and_gate and_gate_u_pg_rca_and1_y0(u_pg_rca_or0_y0, u_pg_rca_fa1_y0, u_pg_rca_and1_y0);
  or_gate or_gate_u_pg_rca_or1_y0(u_pg_rca_and1_y0, u_pg_rca_fa1_y1, u_pg_rca_or1_y0);
  fa_cla fa_cla_u_pg_rca_fa2_y0(a_2, b_2, u_pg_rca_or1_y0, u_pg_rca_fa2_y0, u_pg_rca_fa2_y1, u_pg_rca_fa2_y2);
  and_gate and_gate_u_pg_rca_and2_y0(u_pg_rca_or1_y0, u_pg_rca_fa2_y0, u_pg_rca_and2_y0);
  or_gate or_gate_u_pg_rca_or2_y0(u_pg_rca_and2_y0, u_pg_rca_fa2_y1, u_pg_rca_or2_y0);
  fa_cla fa_cla_u_pg_rca_fa3_y0(a_3, b_3, u_pg_rca_or2_y0, u_pg_rca_fa3_y0, u_pg_rca_fa3_y1, u_pg_rca_fa3_y2);
  and_gate and_gate_u_pg_rca_and3_y0(u_pg_rca_or2_y0, u_pg_rca_fa3_y0, u_pg_rca_and3_y0);
  or_gate or_gate_u_pg_rca_or3_y0(u_pg_rca_and3_y0, u_pg_rca_fa3_y1, u_pg_rca_or3_y0);
  fa_cla fa_cla_u_pg_rca_fa4_y0(a_4, b_4, u_pg_rca_or3_y0, u_pg_rca_fa4_y0, u_pg_rca_fa4_y1, u_pg_rca_fa4_y2);
  and_gate and_gate_u_pg_rca_and4_y0(u_pg_rca_or3_y0, u_pg_rca_fa4_y0, u_pg_rca_and4_y0);
  or_gate or_gate_u_pg_rca_or4_y0(u_pg_rca_and4_y0, u_pg_rca_fa4_y1, u_pg_rca_or4_y0);
  fa_cla fa_cla_u_pg_rca_fa5_y0(a_5, b_5, u_pg_rca_or4_y0, u_pg_rca_fa5_y0, u_pg_rca_fa5_y1, u_pg_rca_fa5_y2);
  and_gate and_gate_u_pg_rca_and5_y0(u_pg_rca_or4_y0, u_pg_rca_fa5_y0, u_pg_rca_and5_y0);
  or_gate or_gate_u_pg_rca_or5_y0(u_pg_rca_and5_y0, u_pg_rca_fa5_y1, u_pg_rca_or5_y0);
  fa_cla fa_cla_u_pg_rca_fa6_y0(a_6, b_6, u_pg_rca_or5_y0, u_pg_rca_fa6_y0, u_pg_rca_fa6_y1, u_pg_rca_fa6_y2);
  and_gate and_gate_u_pg_rca_and6_y0(u_pg_rca_or5_y0, u_pg_rca_fa6_y0, u_pg_rca_and6_y0);
  or_gate or_gate_u_pg_rca_or6_y0(u_pg_rca_and6_y0, u_pg_rca_fa6_y1, u_pg_rca_or6_y0);
  fa_cla fa_cla_u_pg_rca_fa7_y0(a_7, b_7, u_pg_rca_or6_y0, u_pg_rca_fa7_y0, u_pg_rca_fa7_y1, u_pg_rca_fa7_y2);
  and_gate and_gate_u_pg_rca_and7_y0(u_pg_rca_or6_y0, u_pg_rca_fa7_y0, u_pg_rca_and7_y0);
  or_gate or_gate_u_pg_rca_or7_y0(u_pg_rca_and7_y0, u_pg_rca_fa7_y1, u_pg_rca_or7_y0);
  fa_cla fa_cla_u_pg_rca_fa8_y0(a_8, b_8, u_pg_rca_or7_y0, u_pg_rca_fa8_y0, u_pg_rca_fa8_y1, u_pg_rca_fa8_y2);
  and_gate and_gate_u_pg_rca_and8_y0(u_pg_rca_or7_y0, u_pg_rca_fa8_y0, u_pg_rca_and8_y0);
  or_gate or_gate_u_pg_rca_or8_y0(u_pg_rca_and8_y0, u_pg_rca_fa8_y1, u_pg_rca_or8_y0);
  fa_cla fa_cla_u_pg_rca_fa9_y0(a_9, b_9, u_pg_rca_or8_y0, u_pg_rca_fa9_y0, u_pg_rca_fa9_y1, u_pg_rca_fa9_y2);
  and_gate and_gate_u_pg_rca_and9_y0(u_pg_rca_or8_y0, u_pg_rca_fa9_y0, u_pg_rca_and9_y0);
  or_gate or_gate_u_pg_rca_or9_y0(u_pg_rca_and9_y0, u_pg_rca_fa9_y1, u_pg_rca_or9_y0);
  fa_cla fa_cla_u_pg_rca_fa10_y0(a_10, b_10, u_pg_rca_or9_y0, u_pg_rca_fa10_y0, u_pg_rca_fa10_y1, u_pg_rca_fa10_y2);
  and_gate and_gate_u_pg_rca_and10_y0(u_pg_rca_or9_y0, u_pg_rca_fa10_y0, u_pg_rca_and10_y0);
  or_gate or_gate_u_pg_rca_or10_y0(u_pg_rca_and10_y0, u_pg_rca_fa10_y1, u_pg_rca_or10_y0);
  fa_cla fa_cla_u_pg_rca_fa11_y0(a_11, b_11, u_pg_rca_or10_y0, u_pg_rca_fa11_y0, u_pg_rca_fa11_y1, u_pg_rca_fa11_y2);
  and_gate and_gate_u_pg_rca_and11_y0(u_pg_rca_or10_y0, u_pg_rca_fa11_y0, u_pg_rca_and11_y0);
  or_gate or_gate_u_pg_rca_or11_y0(u_pg_rca_and11_y0, u_pg_rca_fa11_y1, u_pg_rca_or11_y0);
  fa_cla fa_cla_u_pg_rca_fa12_y0(a_12, b_12, u_pg_rca_or11_y0, u_pg_rca_fa12_y0, u_pg_rca_fa12_y1, u_pg_rca_fa12_y2);
  and_gate and_gate_u_pg_rca_and12_y0(u_pg_rca_or11_y0, u_pg_rca_fa12_y0, u_pg_rca_and12_y0);
  or_gate or_gate_u_pg_rca_or12_y0(u_pg_rca_and12_y0, u_pg_rca_fa12_y1, u_pg_rca_or12_y0);
  fa_cla fa_cla_u_pg_rca_fa13_y0(a_13, b_13, u_pg_rca_or12_y0, u_pg_rca_fa13_y0, u_pg_rca_fa13_y1, u_pg_rca_fa13_y2);
  and_gate and_gate_u_pg_rca_and13_y0(u_pg_rca_or12_y0, u_pg_rca_fa13_y0, u_pg_rca_and13_y0);
  or_gate or_gate_u_pg_rca_or13_y0(u_pg_rca_and13_y0, u_pg_rca_fa13_y1, u_pg_rca_or13_y0);
  fa_cla fa_cla_u_pg_rca_fa14_y0(a_14, b_14, u_pg_rca_or13_y0, u_pg_rca_fa14_y0, u_pg_rca_fa14_y1, u_pg_rca_fa14_y2);
  and_gate and_gate_u_pg_rca_and14_y0(u_pg_rca_or13_y0, u_pg_rca_fa14_y0, u_pg_rca_and14_y0);
  or_gate or_gate_u_pg_rca_or14_y0(u_pg_rca_and14_y0, u_pg_rca_fa14_y1, u_pg_rca_or14_y0);
  fa_cla fa_cla_u_pg_rca_fa15_y0(a_15, b_15, u_pg_rca_or14_y0, u_pg_rca_fa15_y0, u_pg_rca_fa15_y1, u_pg_rca_fa15_y2);
  and_gate and_gate_u_pg_rca_and15_y0(u_pg_rca_or14_y0, u_pg_rca_fa15_y0, u_pg_rca_and15_y0);
  or_gate or_gate_u_pg_rca_or15_y0(u_pg_rca_and15_y0, u_pg_rca_fa15_y1, u_pg_rca_or15_y0);
  fa_cla fa_cla_u_pg_rca_fa16_y0(a_16, b_16, u_pg_rca_or15_y0, u_pg_rca_fa16_y0, u_pg_rca_fa16_y1, u_pg_rca_fa16_y2);
  and_gate and_gate_u_pg_rca_and16_y0(u_pg_rca_or15_y0, u_pg_rca_fa16_y0, u_pg_rca_and16_y0);
  or_gate or_gate_u_pg_rca_or16_y0(u_pg_rca_and16_y0, u_pg_rca_fa16_y1, u_pg_rca_or16_y0);
  fa_cla fa_cla_u_pg_rca_fa17_y0(a_17, b_17, u_pg_rca_or16_y0, u_pg_rca_fa17_y0, u_pg_rca_fa17_y1, u_pg_rca_fa17_y2);
  and_gate and_gate_u_pg_rca_and17_y0(u_pg_rca_or16_y0, u_pg_rca_fa17_y0, u_pg_rca_and17_y0);
  or_gate or_gate_u_pg_rca_or17_y0(u_pg_rca_and17_y0, u_pg_rca_fa17_y1, u_pg_rca_or17_y0);
  fa_cla fa_cla_u_pg_rca_fa18_y0(a_18, b_18, u_pg_rca_or17_y0, u_pg_rca_fa18_y0, u_pg_rca_fa18_y1, u_pg_rca_fa18_y2);
  and_gate and_gate_u_pg_rca_and18_y0(u_pg_rca_or17_y0, u_pg_rca_fa18_y0, u_pg_rca_and18_y0);
  or_gate or_gate_u_pg_rca_or18_y0(u_pg_rca_and18_y0, u_pg_rca_fa18_y1, u_pg_rca_or18_y0);
  fa_cla fa_cla_u_pg_rca_fa19_y0(a_19, b_19, u_pg_rca_or18_y0, u_pg_rca_fa19_y0, u_pg_rca_fa19_y1, u_pg_rca_fa19_y2);
  and_gate and_gate_u_pg_rca_and19_y0(u_pg_rca_or18_y0, u_pg_rca_fa19_y0, u_pg_rca_and19_y0);
  or_gate or_gate_u_pg_rca_or19_y0(u_pg_rca_and19_y0, u_pg_rca_fa19_y1, u_pg_rca_or19_y0);
  fa_cla fa_cla_u_pg_rca_fa20_y0(a_20, b_20, u_pg_rca_or19_y0, u_pg_rca_fa20_y0, u_pg_rca_fa20_y1, u_pg_rca_fa20_y2);
  and_gate and_gate_u_pg_rca_and20_y0(u_pg_rca_or19_y0, u_pg_rca_fa20_y0, u_pg_rca_and20_y0);
  or_gate or_gate_u_pg_rca_or20_y0(u_pg_rca_and20_y0, u_pg_rca_fa20_y1, u_pg_rca_or20_y0);
  fa_cla fa_cla_u_pg_rca_fa21_y0(a_21, b_21, u_pg_rca_or20_y0, u_pg_rca_fa21_y0, u_pg_rca_fa21_y1, u_pg_rca_fa21_y2);
  and_gate and_gate_u_pg_rca_and21_y0(u_pg_rca_or20_y0, u_pg_rca_fa21_y0, u_pg_rca_and21_y0);
  or_gate or_gate_u_pg_rca_or21_y0(u_pg_rca_and21_y0, u_pg_rca_fa21_y1, u_pg_rca_or21_y0);

  assign out[0] = u_pg_rca_fa0_y2;
  assign out[1] = u_pg_rca_fa1_y2;
  assign out[2] = u_pg_rca_fa2_y2;
  assign out[3] = u_pg_rca_fa3_y2;
  assign out[4] = u_pg_rca_fa4_y2;
  assign out[5] = u_pg_rca_fa5_y2;
  assign out[6] = u_pg_rca_fa6_y2;
  assign out[7] = u_pg_rca_fa7_y2;
  assign out[8] = u_pg_rca_fa8_y2;
  assign out[9] = u_pg_rca_fa9_y2;
  assign out[10] = u_pg_rca_fa10_y2;
  assign out[11] = u_pg_rca_fa11_y2;
  assign out[12] = u_pg_rca_fa12_y2;
  assign out[13] = u_pg_rca_fa13_y2;
  assign out[14] = u_pg_rca_fa14_y2;
  assign out[15] = u_pg_rca_fa15_y2;
  assign out[16] = u_pg_rca_fa16_y2;
  assign out[17] = u_pg_rca_fa17_y2;
  assign out[18] = u_pg_rca_fa18_y2;
  assign out[19] = u_pg_rca_fa19_y2;
  assign out[20] = u_pg_rca_fa20_y2;
  assign out[21] = u_pg_rca_fa21_y2;
  assign out[22] = u_pg_rca_or21_y0;
endmodule

module h_s_dadda_pg_rca12(input [11:0] a, input [11:0] b, output [23:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire constant_wire_1;
  wire h_s_dadda_pg_rca12_and_9_0_y0;
  wire h_s_dadda_pg_rca12_and_8_1_y0;
  wire h_s_dadda_pg_rca12_ha0_y0;
  wire h_s_dadda_pg_rca12_ha0_y1;
  wire h_s_dadda_pg_rca12_and_10_0_y0;
  wire h_s_dadda_pg_rca12_and_9_1_y0;
  wire h_s_dadda_pg_rca12_fa0_y2;
  wire h_s_dadda_pg_rca12_fa0_y4;
  wire h_s_dadda_pg_rca12_and_8_2_y0;
  wire h_s_dadda_pg_rca12_and_7_3_y0;
  wire h_s_dadda_pg_rca12_ha1_y0;
  wire h_s_dadda_pg_rca12_ha1_y1;
  wire h_s_dadda_pg_rca12_nand_11_0_y0;
  wire h_s_dadda_pg_rca12_fa1_y2;
  wire h_s_dadda_pg_rca12_fa1_y4;
  wire h_s_dadda_pg_rca12_and_10_1_y0;
  wire h_s_dadda_pg_rca12_and_9_2_y0;
  wire h_s_dadda_pg_rca12_and_8_3_y0;
  wire h_s_dadda_pg_rca12_fa2_y2;
  wire h_s_dadda_pg_rca12_fa2_y4;
  wire h_s_dadda_pg_rca12_and_7_4_y0;
  wire h_s_dadda_pg_rca12_and_6_5_y0;
  wire h_s_dadda_pg_rca12_ha2_y0;
  wire h_s_dadda_pg_rca12_ha2_y1;
  wire h_s_dadda_pg_rca12_fa3_y2;
  wire h_s_dadda_pg_rca12_fa3_y4;
  wire h_s_dadda_pg_rca12_nand_11_1_y0;
  wire h_s_dadda_pg_rca12_and_10_2_y0;
  wire h_s_dadda_pg_rca12_fa4_y2;
  wire h_s_dadda_pg_rca12_fa4_y4;
  wire h_s_dadda_pg_rca12_and_9_3_y0;
  wire h_s_dadda_pg_rca12_and_8_4_y0;
  wire h_s_dadda_pg_rca12_and_7_5_y0;
  wire h_s_dadda_pg_rca12_fa5_y2;
  wire h_s_dadda_pg_rca12_fa5_y4;
  wire h_s_dadda_pg_rca12_fa6_y2;
  wire h_s_dadda_pg_rca12_fa6_y4;
  wire h_s_dadda_pg_rca12_nand_11_2_y0;
  wire h_s_dadda_pg_rca12_and_10_3_y0;
  wire h_s_dadda_pg_rca12_and_9_4_y0;
  wire h_s_dadda_pg_rca12_fa7_y2;
  wire h_s_dadda_pg_rca12_fa7_y4;
  wire h_s_dadda_pg_rca12_nand_11_3_y0;
  wire h_s_dadda_pg_rca12_fa8_y2;
  wire h_s_dadda_pg_rca12_fa8_y4;
  wire h_s_dadda_pg_rca12_and_4_0_y0;
  wire h_s_dadda_pg_rca12_and_3_1_y0;
  wire h_s_dadda_pg_rca12_ha3_y0;
  wire h_s_dadda_pg_rca12_ha3_y1;
  wire h_s_dadda_pg_rca12_and_5_0_y0;
  wire h_s_dadda_pg_rca12_and_4_1_y0;
  wire h_s_dadda_pg_rca12_fa9_y2;
  wire h_s_dadda_pg_rca12_fa9_y4;
  wire h_s_dadda_pg_rca12_and_3_2_y0;
  wire h_s_dadda_pg_rca12_and_2_3_y0;
  wire h_s_dadda_pg_rca12_ha4_y0;
  wire h_s_dadda_pg_rca12_ha4_y1;
  wire h_s_dadda_pg_rca12_and_6_0_y0;
  wire h_s_dadda_pg_rca12_fa10_y2;
  wire h_s_dadda_pg_rca12_fa10_y4;
  wire h_s_dadda_pg_rca12_and_5_1_y0;
  wire h_s_dadda_pg_rca12_and_4_2_y0;
  wire h_s_dadda_pg_rca12_and_3_3_y0;
  wire h_s_dadda_pg_rca12_fa11_y2;
  wire h_s_dadda_pg_rca12_fa11_y4;
  wire h_s_dadda_pg_rca12_and_2_4_y0;
  wire h_s_dadda_pg_rca12_and_1_5_y0;
  wire h_s_dadda_pg_rca12_ha5_y0;
  wire h_s_dadda_pg_rca12_ha5_y1;
  wire h_s_dadda_pg_rca12_fa12_y2;
  wire h_s_dadda_pg_rca12_fa12_y4;
  wire h_s_dadda_pg_rca12_and_7_0_y0;
  wire h_s_dadda_pg_rca12_and_6_1_y0;
  wire h_s_dadda_pg_rca12_and_5_2_y0;
  wire h_s_dadda_pg_rca12_fa13_y2;
  wire h_s_dadda_pg_rca12_fa13_y4;
  wire h_s_dadda_pg_rca12_and_4_3_y0;
  wire h_s_dadda_pg_rca12_and_3_4_y0;
  wire h_s_dadda_pg_rca12_and_2_5_y0;
  wire h_s_dadda_pg_rca12_fa14_y2;
  wire h_s_dadda_pg_rca12_fa14_y4;
  wire h_s_dadda_pg_rca12_and_1_6_y0;
  wire h_s_dadda_pg_rca12_and_0_7_y0;
  wire h_s_dadda_pg_rca12_ha6_y0;
  wire h_s_dadda_pg_rca12_ha6_y1;
  wire h_s_dadda_pg_rca12_fa15_y2;
  wire h_s_dadda_pg_rca12_fa15_y4;
  wire h_s_dadda_pg_rca12_and_8_0_y0;
  wire h_s_dadda_pg_rca12_and_7_1_y0;
  wire h_s_dadda_pg_rca12_fa16_y2;
  wire h_s_dadda_pg_rca12_fa16_y4;
  wire h_s_dadda_pg_rca12_and_6_2_y0;
  wire h_s_dadda_pg_rca12_and_5_3_y0;
  wire h_s_dadda_pg_rca12_and_4_4_y0;
  wire h_s_dadda_pg_rca12_fa17_y2;
  wire h_s_dadda_pg_rca12_fa17_y4;
  wire h_s_dadda_pg_rca12_and_3_5_y0;
  wire h_s_dadda_pg_rca12_and_2_6_y0;
  wire h_s_dadda_pg_rca12_and_1_7_y0;
  wire h_s_dadda_pg_rca12_fa18_y2;
  wire h_s_dadda_pg_rca12_fa18_y4;
  wire h_s_dadda_pg_rca12_and_0_8_y0;
  wire h_s_dadda_pg_rca12_ha7_y0;
  wire h_s_dadda_pg_rca12_ha7_y1;
  wire h_s_dadda_pg_rca12_fa19_y2;
  wire h_s_dadda_pg_rca12_fa19_y4;
  wire h_s_dadda_pg_rca12_and_7_2_y0;
  wire h_s_dadda_pg_rca12_fa20_y2;
  wire h_s_dadda_pg_rca12_fa20_y4;
  wire h_s_dadda_pg_rca12_and_6_3_y0;
  wire h_s_dadda_pg_rca12_and_5_4_y0;
  wire h_s_dadda_pg_rca12_and_4_5_y0;
  wire h_s_dadda_pg_rca12_fa21_y2;
  wire h_s_dadda_pg_rca12_fa21_y4;
  wire h_s_dadda_pg_rca12_and_3_6_y0;
  wire h_s_dadda_pg_rca12_and_2_7_y0;
  wire h_s_dadda_pg_rca12_and_1_8_y0;
  wire h_s_dadda_pg_rca12_fa22_y2;
  wire h_s_dadda_pg_rca12_fa22_y4;
  wire h_s_dadda_pg_rca12_and_0_9_y0;
  wire h_s_dadda_pg_rca12_fa23_y2;
  wire h_s_dadda_pg_rca12_fa23_y4;
  wire h_s_dadda_pg_rca12_fa24_y2;
  wire h_s_dadda_pg_rca12_fa24_y4;
  wire h_s_dadda_pg_rca12_and_6_4_y0;
  wire h_s_dadda_pg_rca12_fa25_y2;
  wire h_s_dadda_pg_rca12_fa25_y4;
  wire h_s_dadda_pg_rca12_and_5_5_y0;
  wire h_s_dadda_pg_rca12_and_4_6_y0;
  wire h_s_dadda_pg_rca12_and_3_7_y0;
  wire h_s_dadda_pg_rca12_fa26_y2;
  wire h_s_dadda_pg_rca12_fa26_y4;
  wire h_s_dadda_pg_rca12_and_2_8_y0;
  wire h_s_dadda_pg_rca12_and_1_9_y0;
  wire h_s_dadda_pg_rca12_and_0_10_y0;
  wire h_s_dadda_pg_rca12_fa27_y2;
  wire h_s_dadda_pg_rca12_fa27_y4;
  wire h_s_dadda_pg_rca12_fa28_y2;
  wire h_s_dadda_pg_rca12_fa28_y4;
  wire h_s_dadda_pg_rca12_fa29_y2;
  wire h_s_dadda_pg_rca12_fa29_y4;
  wire h_s_dadda_pg_rca12_and_5_6_y0;
  wire h_s_dadda_pg_rca12_fa30_y2;
  wire h_s_dadda_pg_rca12_fa30_y4;
  wire h_s_dadda_pg_rca12_and_4_7_y0;
  wire h_s_dadda_pg_rca12_and_3_8_y0;
  wire h_s_dadda_pg_rca12_and_2_9_y0;
  wire h_s_dadda_pg_rca12_fa31_y2;
  wire h_s_dadda_pg_rca12_fa31_y4;
  wire h_s_dadda_pg_rca12_and_1_10_y0;
  wire h_s_dadda_pg_rca12_nand_0_11_y0;
  wire h_s_dadda_pg_rca12_fa32_y2;
  wire h_s_dadda_pg_rca12_fa32_y4;
  wire h_s_dadda_pg_rca12_fa33_y2;
  wire h_s_dadda_pg_rca12_fa33_y4;
  wire h_s_dadda_pg_rca12_fa34_y2;
  wire h_s_dadda_pg_rca12_fa34_y4;
  wire h_s_dadda_pg_rca12_and_6_6_y0;
  wire h_s_dadda_pg_rca12_fa35_y2;
  wire h_s_dadda_pg_rca12_fa35_y4;
  wire h_s_dadda_pg_rca12_and_5_7_y0;
  wire h_s_dadda_pg_rca12_and_4_8_y0;
  wire h_s_dadda_pg_rca12_and_3_9_y0;
  wire h_s_dadda_pg_rca12_fa36_y2;
  wire h_s_dadda_pg_rca12_fa36_y4;
  wire h_s_dadda_pg_rca12_and_2_10_y0;
  wire h_s_dadda_pg_rca12_nand_1_11_y0;
  wire h_s_dadda_pg_rca12_fa37_y2;
  wire h_s_dadda_pg_rca12_fa37_y4;
  wire h_s_dadda_pg_rca12_fa38_y2;
  wire h_s_dadda_pg_rca12_fa38_y4;
  wire h_s_dadda_pg_rca12_fa39_y2;
  wire h_s_dadda_pg_rca12_fa39_y4;
  wire h_s_dadda_pg_rca12_and_8_5_y0;
  wire h_s_dadda_pg_rca12_fa40_y2;
  wire h_s_dadda_pg_rca12_fa40_y4;
  wire h_s_dadda_pg_rca12_and_7_6_y0;
  wire h_s_dadda_pg_rca12_and_6_7_y0;
  wire h_s_dadda_pg_rca12_and_5_8_y0;
  wire h_s_dadda_pg_rca12_fa41_y2;
  wire h_s_dadda_pg_rca12_fa41_y4;
  wire h_s_dadda_pg_rca12_and_4_9_y0;
  wire h_s_dadda_pg_rca12_and_3_10_y0;
  wire h_s_dadda_pg_rca12_nand_2_11_y0;
  wire h_s_dadda_pg_rca12_fa42_y2;
  wire h_s_dadda_pg_rca12_fa42_y4;
  wire h_s_dadda_pg_rca12_fa43_y2;
  wire h_s_dadda_pg_rca12_fa43_y4;
  wire h_s_dadda_pg_rca12_fa44_y2;
  wire h_s_dadda_pg_rca12_fa44_y4;
  wire h_s_dadda_pg_rca12_and_10_4_y0;
  wire h_s_dadda_pg_rca12_fa45_y2;
  wire h_s_dadda_pg_rca12_fa45_y4;
  wire h_s_dadda_pg_rca12_and_9_5_y0;
  wire h_s_dadda_pg_rca12_and_8_6_y0;
  wire h_s_dadda_pg_rca12_and_7_7_y0;
  wire h_s_dadda_pg_rca12_fa46_y2;
  wire h_s_dadda_pg_rca12_fa46_y4;
  wire h_s_dadda_pg_rca12_and_6_8_y0;
  wire h_s_dadda_pg_rca12_and_5_9_y0;
  wire h_s_dadda_pg_rca12_and_4_10_y0;
  wire h_s_dadda_pg_rca12_fa47_y2;
  wire h_s_dadda_pg_rca12_fa47_y4;
  wire h_s_dadda_pg_rca12_nand_3_11_y0;
  wire h_s_dadda_pg_rca12_fa48_y2;
  wire h_s_dadda_pg_rca12_fa48_y4;
  wire h_s_dadda_pg_rca12_fa49_y2;
  wire h_s_dadda_pg_rca12_fa49_y4;
  wire h_s_dadda_pg_rca12_fa50_y2;
  wire h_s_dadda_pg_rca12_fa50_y4;
  wire h_s_dadda_pg_rca12_nand_11_4_y0;
  wire h_s_dadda_pg_rca12_and_10_5_y0;
  wire h_s_dadda_pg_rca12_and_9_6_y0;
  wire h_s_dadda_pg_rca12_fa51_y2;
  wire h_s_dadda_pg_rca12_fa51_y4;
  wire h_s_dadda_pg_rca12_and_8_7_y0;
  wire h_s_dadda_pg_rca12_and_7_8_y0;
  wire h_s_dadda_pg_rca12_and_6_9_y0;
  wire h_s_dadda_pg_rca12_fa52_y2;
  wire h_s_dadda_pg_rca12_fa52_y4;
  wire h_s_dadda_pg_rca12_and_5_10_y0;
  wire h_s_dadda_pg_rca12_nand_4_11_y0;
  wire h_s_dadda_pg_rca12_fa53_y2;
  wire h_s_dadda_pg_rca12_fa53_y4;
  wire h_s_dadda_pg_rca12_fa54_y2;
  wire h_s_dadda_pg_rca12_fa54_y4;
  wire h_s_dadda_pg_rca12_nand_11_5_y0;
  wire h_s_dadda_pg_rca12_fa55_y2;
  wire h_s_dadda_pg_rca12_fa55_y4;
  wire h_s_dadda_pg_rca12_and_10_6_y0;
  wire h_s_dadda_pg_rca12_and_9_7_y0;
  wire h_s_dadda_pg_rca12_and_8_8_y0;
  wire h_s_dadda_pg_rca12_fa56_y2;
  wire h_s_dadda_pg_rca12_fa56_y4;
  wire h_s_dadda_pg_rca12_and_7_9_y0;
  wire h_s_dadda_pg_rca12_and_6_10_y0;
  wire h_s_dadda_pg_rca12_nand_5_11_y0;
  wire h_s_dadda_pg_rca12_fa57_y2;
  wire h_s_dadda_pg_rca12_fa57_y4;
  wire h_s_dadda_pg_rca12_fa58_y2;
  wire h_s_dadda_pg_rca12_fa58_y4;
  wire h_s_dadda_pg_rca12_nand_11_6_y0;
  wire h_s_dadda_pg_rca12_and_10_7_y0;
  wire h_s_dadda_pg_rca12_fa59_y2;
  wire h_s_dadda_pg_rca12_fa59_y4;
  wire h_s_dadda_pg_rca12_and_9_8_y0;
  wire h_s_dadda_pg_rca12_and_8_9_y0;
  wire h_s_dadda_pg_rca12_and_7_10_y0;
  wire h_s_dadda_pg_rca12_fa60_y2;
  wire h_s_dadda_pg_rca12_fa60_y4;
  wire h_s_dadda_pg_rca12_fa61_y2;
  wire h_s_dadda_pg_rca12_fa61_y4;
  wire h_s_dadda_pg_rca12_nand_11_7_y0;
  wire h_s_dadda_pg_rca12_and_10_8_y0;
  wire h_s_dadda_pg_rca12_and_9_9_y0;
  wire h_s_dadda_pg_rca12_fa62_y2;
  wire h_s_dadda_pg_rca12_fa62_y4;
  wire h_s_dadda_pg_rca12_nand_11_8_y0;
  wire h_s_dadda_pg_rca12_fa63_y2;
  wire h_s_dadda_pg_rca12_fa63_y4;
  wire h_s_dadda_pg_rca12_and_3_0_y0;
  wire h_s_dadda_pg_rca12_and_2_1_y0;
  wire h_s_dadda_pg_rca12_ha8_y0;
  wire h_s_dadda_pg_rca12_ha8_y1;
  wire h_s_dadda_pg_rca12_and_2_2_y0;
  wire h_s_dadda_pg_rca12_and_1_3_y0;
  wire h_s_dadda_pg_rca12_fa64_y2;
  wire h_s_dadda_pg_rca12_fa64_y4;
  wire h_s_dadda_pg_rca12_and_1_4_y0;
  wire h_s_dadda_pg_rca12_and_0_5_y0;
  wire h_s_dadda_pg_rca12_fa65_y2;
  wire h_s_dadda_pg_rca12_fa65_y4;
  wire h_s_dadda_pg_rca12_and_0_6_y0;
  wire h_s_dadda_pg_rca12_fa66_y2;
  wire h_s_dadda_pg_rca12_fa66_y4;
  wire h_s_dadda_pg_rca12_fa67_y2;
  wire h_s_dadda_pg_rca12_fa67_y4;
  wire h_s_dadda_pg_rca12_fa68_y2;
  wire h_s_dadda_pg_rca12_fa68_y4;
  wire h_s_dadda_pg_rca12_fa69_y2;
  wire h_s_dadda_pg_rca12_fa69_y4;
  wire h_s_dadda_pg_rca12_fa70_y2;
  wire h_s_dadda_pg_rca12_fa70_y4;
  wire h_s_dadda_pg_rca12_fa71_y2;
  wire h_s_dadda_pg_rca12_fa71_y4;
  wire h_s_dadda_pg_rca12_fa72_y2;
  wire h_s_dadda_pg_rca12_fa72_y4;
  wire h_s_dadda_pg_rca12_fa73_y2;
  wire h_s_dadda_pg_rca12_fa73_y4;
  wire h_s_dadda_pg_rca12_fa74_y2;
  wire h_s_dadda_pg_rca12_fa74_y4;
  wire h_s_dadda_pg_rca12_fa75_y2;
  wire h_s_dadda_pg_rca12_fa75_y4;
  wire h_s_dadda_pg_rca12_fa76_y2;
  wire h_s_dadda_pg_rca12_fa76_y4;
  wire h_s_dadda_pg_rca12_nand_6_11_y0;
  wire h_s_dadda_pg_rca12_fa77_y2;
  wire h_s_dadda_pg_rca12_fa77_y4;
  wire h_s_dadda_pg_rca12_and_8_10_y0;
  wire h_s_dadda_pg_rca12_nand_7_11_y0;
  wire h_s_dadda_pg_rca12_fa78_y2;
  wire h_s_dadda_pg_rca12_fa78_y4;
  wire h_s_dadda_pg_rca12_and_10_9_y0;
  wire h_s_dadda_pg_rca12_and_9_10_y0;
  wire h_s_dadda_pg_rca12_fa79_y2;
  wire h_s_dadda_pg_rca12_fa79_y4;
  wire h_s_dadda_pg_rca12_nand_11_9_y0;
  wire h_s_dadda_pg_rca12_fa80_y2;
  wire h_s_dadda_pg_rca12_fa80_y4;
  wire h_s_dadda_pg_rca12_and_2_0_y0;
  wire h_s_dadda_pg_rca12_and_1_1_y0;
  wire h_s_dadda_pg_rca12_ha9_y0;
  wire h_s_dadda_pg_rca12_ha9_y1;
  wire h_s_dadda_pg_rca12_and_1_2_y0;
  wire h_s_dadda_pg_rca12_and_0_3_y0;
  wire h_s_dadda_pg_rca12_fa81_y2;
  wire h_s_dadda_pg_rca12_fa81_y4;
  wire h_s_dadda_pg_rca12_and_0_4_y0;
  wire h_s_dadda_pg_rca12_fa82_y2;
  wire h_s_dadda_pg_rca12_fa82_y4;
  wire h_s_dadda_pg_rca12_fa83_y2;
  wire h_s_dadda_pg_rca12_fa83_y4;
  wire h_s_dadda_pg_rca12_fa84_y2;
  wire h_s_dadda_pg_rca12_fa84_y4;
  wire h_s_dadda_pg_rca12_fa85_y2;
  wire h_s_dadda_pg_rca12_fa85_y4;
  wire h_s_dadda_pg_rca12_fa86_y2;
  wire h_s_dadda_pg_rca12_fa86_y4;
  wire h_s_dadda_pg_rca12_fa87_y2;
  wire h_s_dadda_pg_rca12_fa87_y4;
  wire h_s_dadda_pg_rca12_fa88_y2;
  wire h_s_dadda_pg_rca12_fa88_y4;
  wire h_s_dadda_pg_rca12_fa89_y2;
  wire h_s_dadda_pg_rca12_fa89_y4;
  wire h_s_dadda_pg_rca12_fa90_y2;
  wire h_s_dadda_pg_rca12_fa90_y4;
  wire h_s_dadda_pg_rca12_fa91_y2;
  wire h_s_dadda_pg_rca12_fa91_y4;
  wire h_s_dadda_pg_rca12_fa92_y2;
  wire h_s_dadda_pg_rca12_fa92_y4;
  wire h_s_dadda_pg_rca12_fa93_y2;
  wire h_s_dadda_pg_rca12_fa93_y4;
  wire h_s_dadda_pg_rca12_fa94_y2;
  wire h_s_dadda_pg_rca12_fa94_y4;
  wire h_s_dadda_pg_rca12_fa95_y2;
  wire h_s_dadda_pg_rca12_fa95_y4;
  wire h_s_dadda_pg_rca12_fa96_y2;
  wire h_s_dadda_pg_rca12_fa96_y4;
  wire h_s_dadda_pg_rca12_nand_8_11_y0;
  wire h_s_dadda_pg_rca12_fa97_y2;
  wire h_s_dadda_pg_rca12_fa97_y4;
  wire h_s_dadda_pg_rca12_and_10_10_y0;
  wire h_s_dadda_pg_rca12_nand_9_11_y0;
  wire h_s_dadda_pg_rca12_fa98_y2;
  wire h_s_dadda_pg_rca12_fa98_y4;
  wire h_s_dadda_pg_rca12_nand_11_10_y0;
  wire h_s_dadda_pg_rca12_fa99_y2;
  wire h_s_dadda_pg_rca12_fa99_y4;
  wire h_s_dadda_pg_rca12_and_0_0_y0;
  wire h_s_dadda_pg_rca12_and_1_0_y0;
  wire h_s_dadda_pg_rca12_and_0_2_y0;
  wire h_s_dadda_pg_rca12_nand_10_11_y0;
  wire h_s_dadda_pg_rca12_and_0_1_y0;
  wire h_s_dadda_pg_rca12_and_11_11_y0;
  wire [21:0] h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a;
  wire [21:0] h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b;
  wire [22:0] h_s_dadda_pg_rca12_u_pg_rca_out;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa0_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa1_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa2_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa3_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa4_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa5_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa6_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa7_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa8_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa9_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa10_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa11_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa12_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa13_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa14_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa15_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa16_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa17_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa18_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa19_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa20_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_fa21_y2;
  wire h_s_dadda_pg_rca12_u_pg_rca_or21_y0;
  wire h_s_dadda_pg_rca12_xor0_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  constant_wire_value_1 constant_wire_value_1_constant_wire_1(a_0, b_0, constant_wire_1);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_0_y0(a_9, b_0, h_s_dadda_pg_rca12_and_9_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_1_y0(a_8, b_1, h_s_dadda_pg_rca12_and_8_1_y0);
  ha ha_h_s_dadda_pg_rca12_ha0_y0(h_s_dadda_pg_rca12_and_9_0_y0, h_s_dadda_pg_rca12_and_8_1_y0, h_s_dadda_pg_rca12_ha0_y0, h_s_dadda_pg_rca12_ha0_y1);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_0_y0(a_10, b_0, h_s_dadda_pg_rca12_and_10_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_1_y0(a_9, b_1, h_s_dadda_pg_rca12_and_9_1_y0);
  fa fa_h_s_dadda_pg_rca12_fa0_y2(h_s_dadda_pg_rca12_ha0_y1, h_s_dadda_pg_rca12_and_10_0_y0, h_s_dadda_pg_rca12_and_9_1_y0, h_s_dadda_pg_rca12_fa0_y2, h_s_dadda_pg_rca12_fa0_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_2_y0(a_8, b_2, h_s_dadda_pg_rca12_and_8_2_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_3_y0(a_7, b_3, h_s_dadda_pg_rca12_and_7_3_y0);
  ha ha_h_s_dadda_pg_rca12_ha1_y0(h_s_dadda_pg_rca12_and_8_2_y0, h_s_dadda_pg_rca12_and_7_3_y0, h_s_dadda_pg_rca12_ha1_y0, h_s_dadda_pg_rca12_ha1_y1);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_0_y0(a_11, b_0, h_s_dadda_pg_rca12_nand_11_0_y0);
  fa fa_h_s_dadda_pg_rca12_fa1_y2(h_s_dadda_pg_rca12_ha1_y1, h_s_dadda_pg_rca12_fa0_y4, h_s_dadda_pg_rca12_nand_11_0_y0, h_s_dadda_pg_rca12_fa1_y2, h_s_dadda_pg_rca12_fa1_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_1_y0(a_10, b_1, h_s_dadda_pg_rca12_and_10_1_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_2_y0(a_9, b_2, h_s_dadda_pg_rca12_and_9_2_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_3_y0(a_8, b_3, h_s_dadda_pg_rca12_and_8_3_y0);
  fa fa_h_s_dadda_pg_rca12_fa2_y2(h_s_dadda_pg_rca12_and_10_1_y0, h_s_dadda_pg_rca12_and_9_2_y0, h_s_dadda_pg_rca12_and_8_3_y0, h_s_dadda_pg_rca12_fa2_y2, h_s_dadda_pg_rca12_fa2_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_4_y0(a_7, b_4, h_s_dadda_pg_rca12_and_7_4_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_5_y0(a_6, b_5, h_s_dadda_pg_rca12_and_6_5_y0);
  ha ha_h_s_dadda_pg_rca12_ha2_y0(h_s_dadda_pg_rca12_and_7_4_y0, h_s_dadda_pg_rca12_and_6_5_y0, h_s_dadda_pg_rca12_ha2_y0, h_s_dadda_pg_rca12_ha2_y1);
  fa fa_h_s_dadda_pg_rca12_fa3_y2(h_s_dadda_pg_rca12_ha2_y1, h_s_dadda_pg_rca12_fa2_y4, h_s_dadda_pg_rca12_fa1_y4, h_s_dadda_pg_rca12_fa3_y2, h_s_dadda_pg_rca12_fa3_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_1_y0(a_11, b_1, h_s_dadda_pg_rca12_nand_11_1_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_2_y0(a_10, b_2, h_s_dadda_pg_rca12_and_10_2_y0);
  fa fa_h_s_dadda_pg_rca12_fa4_y2(constant_wire_1, h_s_dadda_pg_rca12_nand_11_1_y0, h_s_dadda_pg_rca12_and_10_2_y0, h_s_dadda_pg_rca12_fa4_y2, h_s_dadda_pg_rca12_fa4_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_3_y0(a_9, b_3, h_s_dadda_pg_rca12_and_9_3_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_4_y0(a_8, b_4, h_s_dadda_pg_rca12_and_8_4_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_5_y0(a_7, b_5, h_s_dadda_pg_rca12_and_7_5_y0);
  fa fa_h_s_dadda_pg_rca12_fa5_y2(h_s_dadda_pg_rca12_and_9_3_y0, h_s_dadda_pg_rca12_and_8_4_y0, h_s_dadda_pg_rca12_and_7_5_y0, h_s_dadda_pg_rca12_fa5_y2, h_s_dadda_pg_rca12_fa5_y4);
  fa fa_h_s_dadda_pg_rca12_fa6_y2(h_s_dadda_pg_rca12_fa5_y4, h_s_dadda_pg_rca12_fa4_y4, h_s_dadda_pg_rca12_fa3_y4, h_s_dadda_pg_rca12_fa6_y2, h_s_dadda_pg_rca12_fa6_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_2_y0(a_11, b_2, h_s_dadda_pg_rca12_nand_11_2_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_3_y0(a_10, b_3, h_s_dadda_pg_rca12_and_10_3_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_4_y0(a_9, b_4, h_s_dadda_pg_rca12_and_9_4_y0);
  fa fa_h_s_dadda_pg_rca12_fa7_y2(h_s_dadda_pg_rca12_nand_11_2_y0, h_s_dadda_pg_rca12_and_10_3_y0, h_s_dadda_pg_rca12_and_9_4_y0, h_s_dadda_pg_rca12_fa7_y2, h_s_dadda_pg_rca12_fa7_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_3_y0(a_11, b_3, h_s_dadda_pg_rca12_nand_11_3_y0);
  fa fa_h_s_dadda_pg_rca12_fa8_y2(h_s_dadda_pg_rca12_fa7_y4, h_s_dadda_pg_rca12_fa6_y4, h_s_dadda_pg_rca12_nand_11_3_y0, h_s_dadda_pg_rca12_fa8_y2, h_s_dadda_pg_rca12_fa8_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_0_y0(a_4, b_0, h_s_dadda_pg_rca12_and_4_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_1_y0(a_3, b_1, h_s_dadda_pg_rca12_and_3_1_y0);
  ha ha_h_s_dadda_pg_rca12_ha3_y0(h_s_dadda_pg_rca12_and_4_0_y0, h_s_dadda_pg_rca12_and_3_1_y0, h_s_dadda_pg_rca12_ha3_y0, h_s_dadda_pg_rca12_ha3_y1);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_0_y0(a_5, b_0, h_s_dadda_pg_rca12_and_5_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_1_y0(a_4, b_1, h_s_dadda_pg_rca12_and_4_1_y0);
  fa fa_h_s_dadda_pg_rca12_fa9_y2(h_s_dadda_pg_rca12_ha3_y1, h_s_dadda_pg_rca12_and_5_0_y0, h_s_dadda_pg_rca12_and_4_1_y0, h_s_dadda_pg_rca12_fa9_y2, h_s_dadda_pg_rca12_fa9_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_2_y0(a_3, b_2, h_s_dadda_pg_rca12_and_3_2_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_3_y0(a_2, b_3, h_s_dadda_pg_rca12_and_2_3_y0);
  ha ha_h_s_dadda_pg_rca12_ha4_y0(h_s_dadda_pg_rca12_and_3_2_y0, h_s_dadda_pg_rca12_and_2_3_y0, h_s_dadda_pg_rca12_ha4_y0, h_s_dadda_pg_rca12_ha4_y1);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_0_y0(a_6, b_0, h_s_dadda_pg_rca12_and_6_0_y0);
  fa fa_h_s_dadda_pg_rca12_fa10_y2(h_s_dadda_pg_rca12_ha4_y1, h_s_dadda_pg_rca12_fa9_y4, h_s_dadda_pg_rca12_and_6_0_y0, h_s_dadda_pg_rca12_fa10_y2, h_s_dadda_pg_rca12_fa10_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_1_y0(a_5, b_1, h_s_dadda_pg_rca12_and_5_1_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_2_y0(a_4, b_2, h_s_dadda_pg_rca12_and_4_2_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_3_y0(a_3, b_3, h_s_dadda_pg_rca12_and_3_3_y0);
  fa fa_h_s_dadda_pg_rca12_fa11_y2(h_s_dadda_pg_rca12_and_5_1_y0, h_s_dadda_pg_rca12_and_4_2_y0, h_s_dadda_pg_rca12_and_3_3_y0, h_s_dadda_pg_rca12_fa11_y2, h_s_dadda_pg_rca12_fa11_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_4_y0(a_2, b_4, h_s_dadda_pg_rca12_and_2_4_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_5_y0(a_1, b_5, h_s_dadda_pg_rca12_and_1_5_y0);
  ha ha_h_s_dadda_pg_rca12_ha5_y0(h_s_dadda_pg_rca12_and_2_4_y0, h_s_dadda_pg_rca12_and_1_5_y0, h_s_dadda_pg_rca12_ha5_y0, h_s_dadda_pg_rca12_ha5_y1);
  fa fa_h_s_dadda_pg_rca12_fa12_y2(h_s_dadda_pg_rca12_ha5_y1, h_s_dadda_pg_rca12_fa11_y4, h_s_dadda_pg_rca12_fa10_y4, h_s_dadda_pg_rca12_fa12_y2, h_s_dadda_pg_rca12_fa12_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_0_y0(a_7, b_0, h_s_dadda_pg_rca12_and_7_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_1_y0(a_6, b_1, h_s_dadda_pg_rca12_and_6_1_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_2_y0(a_5, b_2, h_s_dadda_pg_rca12_and_5_2_y0);
  fa fa_h_s_dadda_pg_rca12_fa13_y2(h_s_dadda_pg_rca12_and_7_0_y0, h_s_dadda_pg_rca12_and_6_1_y0, h_s_dadda_pg_rca12_and_5_2_y0, h_s_dadda_pg_rca12_fa13_y2, h_s_dadda_pg_rca12_fa13_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_3_y0(a_4, b_3, h_s_dadda_pg_rca12_and_4_3_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_4_y0(a_3, b_4, h_s_dadda_pg_rca12_and_3_4_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_5_y0(a_2, b_5, h_s_dadda_pg_rca12_and_2_5_y0);
  fa fa_h_s_dadda_pg_rca12_fa14_y2(h_s_dadda_pg_rca12_and_4_3_y0, h_s_dadda_pg_rca12_and_3_4_y0, h_s_dadda_pg_rca12_and_2_5_y0, h_s_dadda_pg_rca12_fa14_y2, h_s_dadda_pg_rca12_fa14_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_6_y0(a_1, b_6, h_s_dadda_pg_rca12_and_1_6_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_7_y0(a_0, b_7, h_s_dadda_pg_rca12_and_0_7_y0);
  ha ha_h_s_dadda_pg_rca12_ha6_y0(h_s_dadda_pg_rca12_and_1_6_y0, h_s_dadda_pg_rca12_and_0_7_y0, h_s_dadda_pg_rca12_ha6_y0, h_s_dadda_pg_rca12_ha6_y1);
  fa fa_h_s_dadda_pg_rca12_fa15_y2(h_s_dadda_pg_rca12_ha6_y1, h_s_dadda_pg_rca12_fa14_y4, h_s_dadda_pg_rca12_fa13_y4, h_s_dadda_pg_rca12_fa15_y2, h_s_dadda_pg_rca12_fa15_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_0_y0(a_8, b_0, h_s_dadda_pg_rca12_and_8_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_1_y0(a_7, b_1, h_s_dadda_pg_rca12_and_7_1_y0);
  fa fa_h_s_dadda_pg_rca12_fa16_y2(h_s_dadda_pg_rca12_fa12_y4, h_s_dadda_pg_rca12_and_8_0_y0, h_s_dadda_pg_rca12_and_7_1_y0, h_s_dadda_pg_rca12_fa16_y2, h_s_dadda_pg_rca12_fa16_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_2_y0(a_6, b_2, h_s_dadda_pg_rca12_and_6_2_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_3_y0(a_5, b_3, h_s_dadda_pg_rca12_and_5_3_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_4_y0(a_4, b_4, h_s_dadda_pg_rca12_and_4_4_y0);
  fa fa_h_s_dadda_pg_rca12_fa17_y2(h_s_dadda_pg_rca12_and_6_2_y0, h_s_dadda_pg_rca12_and_5_3_y0, h_s_dadda_pg_rca12_and_4_4_y0, h_s_dadda_pg_rca12_fa17_y2, h_s_dadda_pg_rca12_fa17_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_5_y0(a_3, b_5, h_s_dadda_pg_rca12_and_3_5_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_6_y0(a_2, b_6, h_s_dadda_pg_rca12_and_2_6_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_7_y0(a_1, b_7, h_s_dadda_pg_rca12_and_1_7_y0);
  fa fa_h_s_dadda_pg_rca12_fa18_y2(h_s_dadda_pg_rca12_and_3_5_y0, h_s_dadda_pg_rca12_and_2_6_y0, h_s_dadda_pg_rca12_and_1_7_y0, h_s_dadda_pg_rca12_fa18_y2, h_s_dadda_pg_rca12_fa18_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_8_y0(a_0, b_8, h_s_dadda_pg_rca12_and_0_8_y0);
  ha ha_h_s_dadda_pg_rca12_ha7_y0(h_s_dadda_pg_rca12_and_0_8_y0, h_s_dadda_pg_rca12_fa15_y2, h_s_dadda_pg_rca12_ha7_y0, h_s_dadda_pg_rca12_ha7_y1);
  fa fa_h_s_dadda_pg_rca12_fa19_y2(h_s_dadda_pg_rca12_ha7_y1, h_s_dadda_pg_rca12_fa18_y4, h_s_dadda_pg_rca12_fa17_y4, h_s_dadda_pg_rca12_fa19_y2, h_s_dadda_pg_rca12_fa19_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_2_y0(a_7, b_2, h_s_dadda_pg_rca12_and_7_2_y0);
  fa fa_h_s_dadda_pg_rca12_fa20_y2(h_s_dadda_pg_rca12_fa16_y4, h_s_dadda_pg_rca12_fa15_y4, h_s_dadda_pg_rca12_and_7_2_y0, h_s_dadda_pg_rca12_fa20_y2, h_s_dadda_pg_rca12_fa20_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_3_y0(a_6, b_3, h_s_dadda_pg_rca12_and_6_3_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_4_y0(a_5, b_4, h_s_dadda_pg_rca12_and_5_4_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_5_y0(a_4, b_5, h_s_dadda_pg_rca12_and_4_5_y0);
  fa fa_h_s_dadda_pg_rca12_fa21_y2(h_s_dadda_pg_rca12_and_6_3_y0, h_s_dadda_pg_rca12_and_5_4_y0, h_s_dadda_pg_rca12_and_4_5_y0, h_s_dadda_pg_rca12_fa21_y2, h_s_dadda_pg_rca12_fa21_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_6_y0(a_3, b_6, h_s_dadda_pg_rca12_and_3_6_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_7_y0(a_2, b_7, h_s_dadda_pg_rca12_and_2_7_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_8_y0(a_1, b_8, h_s_dadda_pg_rca12_and_1_8_y0);
  fa fa_h_s_dadda_pg_rca12_fa22_y2(h_s_dadda_pg_rca12_and_3_6_y0, h_s_dadda_pg_rca12_and_2_7_y0, h_s_dadda_pg_rca12_and_1_8_y0, h_s_dadda_pg_rca12_fa22_y2, h_s_dadda_pg_rca12_fa22_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_9_y0(a_0, b_9, h_s_dadda_pg_rca12_and_0_9_y0);
  fa fa_h_s_dadda_pg_rca12_fa23_y2(h_s_dadda_pg_rca12_and_0_9_y0, h_s_dadda_pg_rca12_ha0_y0, h_s_dadda_pg_rca12_fa19_y2, h_s_dadda_pg_rca12_fa23_y2, h_s_dadda_pg_rca12_fa23_y4);
  fa fa_h_s_dadda_pg_rca12_fa24_y2(h_s_dadda_pg_rca12_fa23_y4, h_s_dadda_pg_rca12_fa22_y4, h_s_dadda_pg_rca12_fa21_y4, h_s_dadda_pg_rca12_fa24_y2, h_s_dadda_pg_rca12_fa24_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_4_y0(a_6, b_4, h_s_dadda_pg_rca12_and_6_4_y0);
  fa fa_h_s_dadda_pg_rca12_fa25_y2(h_s_dadda_pg_rca12_fa20_y4, h_s_dadda_pg_rca12_fa19_y4, h_s_dadda_pg_rca12_and_6_4_y0, h_s_dadda_pg_rca12_fa25_y2, h_s_dadda_pg_rca12_fa25_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_5_y0(a_5, b_5, h_s_dadda_pg_rca12_and_5_5_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_6_y0(a_4, b_6, h_s_dadda_pg_rca12_and_4_6_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_7_y0(a_3, b_7, h_s_dadda_pg_rca12_and_3_7_y0);
  fa fa_h_s_dadda_pg_rca12_fa26_y2(h_s_dadda_pg_rca12_and_5_5_y0, h_s_dadda_pg_rca12_and_4_6_y0, h_s_dadda_pg_rca12_and_3_7_y0, h_s_dadda_pg_rca12_fa26_y2, h_s_dadda_pg_rca12_fa26_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_8_y0(a_2, b_8, h_s_dadda_pg_rca12_and_2_8_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_9_y0(a_1, b_9, h_s_dadda_pg_rca12_and_1_9_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_10_y0(a_0, b_10, h_s_dadda_pg_rca12_and_0_10_y0);
  fa fa_h_s_dadda_pg_rca12_fa27_y2(h_s_dadda_pg_rca12_and_2_8_y0, h_s_dadda_pg_rca12_and_1_9_y0, h_s_dadda_pg_rca12_and_0_10_y0, h_s_dadda_pg_rca12_fa27_y2, h_s_dadda_pg_rca12_fa27_y4);
  fa fa_h_s_dadda_pg_rca12_fa28_y2(h_s_dadda_pg_rca12_fa0_y2, h_s_dadda_pg_rca12_ha1_y0, h_s_dadda_pg_rca12_fa24_y2, h_s_dadda_pg_rca12_fa28_y2, h_s_dadda_pg_rca12_fa28_y4);
  fa fa_h_s_dadda_pg_rca12_fa29_y2(h_s_dadda_pg_rca12_fa28_y4, h_s_dadda_pg_rca12_fa27_y4, h_s_dadda_pg_rca12_fa26_y4, h_s_dadda_pg_rca12_fa29_y2, h_s_dadda_pg_rca12_fa29_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_6_y0(a_5, b_6, h_s_dadda_pg_rca12_and_5_6_y0);
  fa fa_h_s_dadda_pg_rca12_fa30_y2(h_s_dadda_pg_rca12_fa25_y4, h_s_dadda_pg_rca12_fa24_y4, h_s_dadda_pg_rca12_and_5_6_y0, h_s_dadda_pg_rca12_fa30_y2, h_s_dadda_pg_rca12_fa30_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_7_y0(a_4, b_7, h_s_dadda_pg_rca12_and_4_7_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_8_y0(a_3, b_8, h_s_dadda_pg_rca12_and_3_8_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_9_y0(a_2, b_9, h_s_dadda_pg_rca12_and_2_9_y0);
  fa fa_h_s_dadda_pg_rca12_fa31_y2(h_s_dadda_pg_rca12_and_4_7_y0, h_s_dadda_pg_rca12_and_3_8_y0, h_s_dadda_pg_rca12_and_2_9_y0, h_s_dadda_pg_rca12_fa31_y2, h_s_dadda_pg_rca12_fa31_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_10_y0(a_1, b_10, h_s_dadda_pg_rca12_and_1_10_y0);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_0_11_y0(a_0, b_11, h_s_dadda_pg_rca12_nand_0_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa32_y2(h_s_dadda_pg_rca12_and_1_10_y0, h_s_dadda_pg_rca12_nand_0_11_y0, h_s_dadda_pg_rca12_fa1_y2, h_s_dadda_pg_rca12_fa32_y2, h_s_dadda_pg_rca12_fa32_y4);
  fa fa_h_s_dadda_pg_rca12_fa33_y2(h_s_dadda_pg_rca12_fa2_y2, h_s_dadda_pg_rca12_ha2_y0, h_s_dadda_pg_rca12_fa29_y2, h_s_dadda_pg_rca12_fa33_y2, h_s_dadda_pg_rca12_fa33_y4);
  fa fa_h_s_dadda_pg_rca12_fa34_y2(h_s_dadda_pg_rca12_fa33_y4, h_s_dadda_pg_rca12_fa32_y4, h_s_dadda_pg_rca12_fa31_y4, h_s_dadda_pg_rca12_fa34_y2, h_s_dadda_pg_rca12_fa34_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_6_y0(a_6, b_6, h_s_dadda_pg_rca12_and_6_6_y0);
  fa fa_h_s_dadda_pg_rca12_fa35_y2(h_s_dadda_pg_rca12_fa30_y4, h_s_dadda_pg_rca12_fa29_y4, h_s_dadda_pg_rca12_and_6_6_y0, h_s_dadda_pg_rca12_fa35_y2, h_s_dadda_pg_rca12_fa35_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_7_y0(a_5, b_7, h_s_dadda_pg_rca12_and_5_7_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_8_y0(a_4, b_8, h_s_dadda_pg_rca12_and_4_8_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_9_y0(a_3, b_9, h_s_dadda_pg_rca12_and_3_9_y0);
  fa fa_h_s_dadda_pg_rca12_fa36_y2(h_s_dadda_pg_rca12_and_5_7_y0, h_s_dadda_pg_rca12_and_4_8_y0, h_s_dadda_pg_rca12_and_3_9_y0, h_s_dadda_pg_rca12_fa36_y2, h_s_dadda_pg_rca12_fa36_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_10_y0(a_2, b_10, h_s_dadda_pg_rca12_and_2_10_y0);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_1_11_y0(a_1, b_11, h_s_dadda_pg_rca12_nand_1_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa37_y2(h_s_dadda_pg_rca12_and_2_10_y0, h_s_dadda_pg_rca12_nand_1_11_y0, h_s_dadda_pg_rca12_fa3_y2, h_s_dadda_pg_rca12_fa37_y2, h_s_dadda_pg_rca12_fa37_y4);
  fa fa_h_s_dadda_pg_rca12_fa38_y2(h_s_dadda_pg_rca12_fa4_y2, h_s_dadda_pg_rca12_fa5_y2, h_s_dadda_pg_rca12_fa34_y2, h_s_dadda_pg_rca12_fa38_y2, h_s_dadda_pg_rca12_fa38_y4);
  fa fa_h_s_dadda_pg_rca12_fa39_y2(h_s_dadda_pg_rca12_fa38_y4, h_s_dadda_pg_rca12_fa37_y4, h_s_dadda_pg_rca12_fa36_y4, h_s_dadda_pg_rca12_fa39_y2, h_s_dadda_pg_rca12_fa39_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_5_y0(a_8, b_5, h_s_dadda_pg_rca12_and_8_5_y0);
  fa fa_h_s_dadda_pg_rca12_fa40_y2(h_s_dadda_pg_rca12_fa35_y4, h_s_dadda_pg_rca12_fa34_y4, h_s_dadda_pg_rca12_and_8_5_y0, h_s_dadda_pg_rca12_fa40_y2, h_s_dadda_pg_rca12_fa40_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_6_y0(a_7, b_6, h_s_dadda_pg_rca12_and_7_6_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_7_y0(a_6, b_7, h_s_dadda_pg_rca12_and_6_7_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_8_y0(a_5, b_8, h_s_dadda_pg_rca12_and_5_8_y0);
  fa fa_h_s_dadda_pg_rca12_fa41_y2(h_s_dadda_pg_rca12_and_7_6_y0, h_s_dadda_pg_rca12_and_6_7_y0, h_s_dadda_pg_rca12_and_5_8_y0, h_s_dadda_pg_rca12_fa41_y2, h_s_dadda_pg_rca12_fa41_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_9_y0(a_4, b_9, h_s_dadda_pg_rca12_and_4_9_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_10_y0(a_3, b_10, h_s_dadda_pg_rca12_and_3_10_y0);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_2_11_y0(a_2, b_11, h_s_dadda_pg_rca12_nand_2_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa42_y2(h_s_dadda_pg_rca12_and_4_9_y0, h_s_dadda_pg_rca12_and_3_10_y0, h_s_dadda_pg_rca12_nand_2_11_y0, h_s_dadda_pg_rca12_fa42_y2, h_s_dadda_pg_rca12_fa42_y4);
  fa fa_h_s_dadda_pg_rca12_fa43_y2(h_s_dadda_pg_rca12_fa6_y2, h_s_dadda_pg_rca12_fa7_y2, h_s_dadda_pg_rca12_fa39_y2, h_s_dadda_pg_rca12_fa43_y2, h_s_dadda_pg_rca12_fa43_y4);
  fa fa_h_s_dadda_pg_rca12_fa44_y2(h_s_dadda_pg_rca12_fa43_y4, h_s_dadda_pg_rca12_fa42_y4, h_s_dadda_pg_rca12_fa41_y4, h_s_dadda_pg_rca12_fa44_y2, h_s_dadda_pg_rca12_fa44_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_4_y0(a_10, b_4, h_s_dadda_pg_rca12_and_10_4_y0);
  fa fa_h_s_dadda_pg_rca12_fa45_y2(h_s_dadda_pg_rca12_fa40_y4, h_s_dadda_pg_rca12_fa39_y4, h_s_dadda_pg_rca12_and_10_4_y0, h_s_dadda_pg_rca12_fa45_y2, h_s_dadda_pg_rca12_fa45_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_5_y0(a_9, b_5, h_s_dadda_pg_rca12_and_9_5_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_6_y0(a_8, b_6, h_s_dadda_pg_rca12_and_8_6_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_7_y0(a_7, b_7, h_s_dadda_pg_rca12_and_7_7_y0);
  fa fa_h_s_dadda_pg_rca12_fa46_y2(h_s_dadda_pg_rca12_and_9_5_y0, h_s_dadda_pg_rca12_and_8_6_y0, h_s_dadda_pg_rca12_and_7_7_y0, h_s_dadda_pg_rca12_fa46_y2, h_s_dadda_pg_rca12_fa46_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_8_y0(a_6, b_8, h_s_dadda_pg_rca12_and_6_8_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_9_y0(a_5, b_9, h_s_dadda_pg_rca12_and_5_9_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_4_10_y0(a_4, b_10, h_s_dadda_pg_rca12_and_4_10_y0);
  fa fa_h_s_dadda_pg_rca12_fa47_y2(h_s_dadda_pg_rca12_and_6_8_y0, h_s_dadda_pg_rca12_and_5_9_y0, h_s_dadda_pg_rca12_and_4_10_y0, h_s_dadda_pg_rca12_fa47_y2, h_s_dadda_pg_rca12_fa47_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_3_11_y0(a_3, b_11, h_s_dadda_pg_rca12_nand_3_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa48_y2(h_s_dadda_pg_rca12_nand_3_11_y0, h_s_dadda_pg_rca12_fa8_y2, h_s_dadda_pg_rca12_fa44_y2, h_s_dadda_pg_rca12_fa48_y2, h_s_dadda_pg_rca12_fa48_y4);
  fa fa_h_s_dadda_pg_rca12_fa49_y2(h_s_dadda_pg_rca12_fa48_y4, h_s_dadda_pg_rca12_fa47_y4, h_s_dadda_pg_rca12_fa46_y4, h_s_dadda_pg_rca12_fa49_y2, h_s_dadda_pg_rca12_fa49_y4);
  fa fa_h_s_dadda_pg_rca12_fa50_y2(h_s_dadda_pg_rca12_fa45_y4, h_s_dadda_pg_rca12_fa44_y4, h_s_dadda_pg_rca12_fa8_y4, h_s_dadda_pg_rca12_fa50_y2, h_s_dadda_pg_rca12_fa50_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_4_y0(a_11, b_4, h_s_dadda_pg_rca12_nand_11_4_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_5_y0(a_10, b_5, h_s_dadda_pg_rca12_and_10_5_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_6_y0(a_9, b_6, h_s_dadda_pg_rca12_and_9_6_y0);
  fa fa_h_s_dadda_pg_rca12_fa51_y2(h_s_dadda_pg_rca12_nand_11_4_y0, h_s_dadda_pg_rca12_and_10_5_y0, h_s_dadda_pg_rca12_and_9_6_y0, h_s_dadda_pg_rca12_fa51_y2, h_s_dadda_pg_rca12_fa51_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_7_y0(a_8, b_7, h_s_dadda_pg_rca12_and_8_7_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_8_y0(a_7, b_8, h_s_dadda_pg_rca12_and_7_8_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_9_y0(a_6, b_9, h_s_dadda_pg_rca12_and_6_9_y0);
  fa fa_h_s_dadda_pg_rca12_fa52_y2(h_s_dadda_pg_rca12_and_8_7_y0, h_s_dadda_pg_rca12_and_7_8_y0, h_s_dadda_pg_rca12_and_6_9_y0, h_s_dadda_pg_rca12_fa52_y2, h_s_dadda_pg_rca12_fa52_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_5_10_y0(a_5, b_10, h_s_dadda_pg_rca12_and_5_10_y0);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_4_11_y0(a_4, b_11, h_s_dadda_pg_rca12_nand_4_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa53_y2(h_s_dadda_pg_rca12_and_5_10_y0, h_s_dadda_pg_rca12_nand_4_11_y0, h_s_dadda_pg_rca12_fa49_y2, h_s_dadda_pg_rca12_fa53_y2, h_s_dadda_pg_rca12_fa53_y4);
  fa fa_h_s_dadda_pg_rca12_fa54_y2(h_s_dadda_pg_rca12_fa53_y4, h_s_dadda_pg_rca12_fa52_y4, h_s_dadda_pg_rca12_fa51_y4, h_s_dadda_pg_rca12_fa54_y2, h_s_dadda_pg_rca12_fa54_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_5_y0(a_11, b_5, h_s_dadda_pg_rca12_nand_11_5_y0);
  fa fa_h_s_dadda_pg_rca12_fa55_y2(h_s_dadda_pg_rca12_fa50_y4, h_s_dadda_pg_rca12_fa49_y4, h_s_dadda_pg_rca12_nand_11_5_y0, h_s_dadda_pg_rca12_fa55_y2, h_s_dadda_pg_rca12_fa55_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_6_y0(a_10, b_6, h_s_dadda_pg_rca12_and_10_6_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_7_y0(a_9, b_7, h_s_dadda_pg_rca12_and_9_7_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_8_y0(a_8, b_8, h_s_dadda_pg_rca12_and_8_8_y0);
  fa fa_h_s_dadda_pg_rca12_fa56_y2(h_s_dadda_pg_rca12_and_10_6_y0, h_s_dadda_pg_rca12_and_9_7_y0, h_s_dadda_pg_rca12_and_8_8_y0, h_s_dadda_pg_rca12_fa56_y2, h_s_dadda_pg_rca12_fa56_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_9_y0(a_7, b_9, h_s_dadda_pg_rca12_and_7_9_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_6_10_y0(a_6, b_10, h_s_dadda_pg_rca12_and_6_10_y0);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_5_11_y0(a_5, b_11, h_s_dadda_pg_rca12_nand_5_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa57_y2(h_s_dadda_pg_rca12_and_7_9_y0, h_s_dadda_pg_rca12_and_6_10_y0, h_s_dadda_pg_rca12_nand_5_11_y0, h_s_dadda_pg_rca12_fa57_y2, h_s_dadda_pg_rca12_fa57_y4);
  fa fa_h_s_dadda_pg_rca12_fa58_y2(h_s_dadda_pg_rca12_fa57_y4, h_s_dadda_pg_rca12_fa56_y4, h_s_dadda_pg_rca12_fa55_y4, h_s_dadda_pg_rca12_fa58_y2, h_s_dadda_pg_rca12_fa58_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_6_y0(a_11, b_6, h_s_dadda_pg_rca12_nand_11_6_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_7_y0(a_10, b_7, h_s_dadda_pg_rca12_and_10_7_y0);
  fa fa_h_s_dadda_pg_rca12_fa59_y2(h_s_dadda_pg_rca12_fa54_y4, h_s_dadda_pg_rca12_nand_11_6_y0, h_s_dadda_pg_rca12_and_10_7_y0, h_s_dadda_pg_rca12_fa59_y2, h_s_dadda_pg_rca12_fa59_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_8_y0(a_9, b_8, h_s_dadda_pg_rca12_and_9_8_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_9_y0(a_8, b_9, h_s_dadda_pg_rca12_and_8_9_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_7_10_y0(a_7, b_10, h_s_dadda_pg_rca12_and_7_10_y0);
  fa fa_h_s_dadda_pg_rca12_fa60_y2(h_s_dadda_pg_rca12_and_9_8_y0, h_s_dadda_pg_rca12_and_8_9_y0, h_s_dadda_pg_rca12_and_7_10_y0, h_s_dadda_pg_rca12_fa60_y2, h_s_dadda_pg_rca12_fa60_y4);
  fa fa_h_s_dadda_pg_rca12_fa61_y2(h_s_dadda_pg_rca12_fa60_y4, h_s_dadda_pg_rca12_fa59_y4, h_s_dadda_pg_rca12_fa58_y4, h_s_dadda_pg_rca12_fa61_y2, h_s_dadda_pg_rca12_fa61_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_7_y0(a_11, b_7, h_s_dadda_pg_rca12_nand_11_7_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_8_y0(a_10, b_8, h_s_dadda_pg_rca12_and_10_8_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_9_y0(a_9, b_9, h_s_dadda_pg_rca12_and_9_9_y0);
  fa fa_h_s_dadda_pg_rca12_fa62_y2(h_s_dadda_pg_rca12_nand_11_7_y0, h_s_dadda_pg_rca12_and_10_8_y0, h_s_dadda_pg_rca12_and_9_9_y0, h_s_dadda_pg_rca12_fa62_y2, h_s_dadda_pg_rca12_fa62_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_8_y0(a_11, b_8, h_s_dadda_pg_rca12_nand_11_8_y0);
  fa fa_h_s_dadda_pg_rca12_fa63_y2(h_s_dadda_pg_rca12_fa62_y4, h_s_dadda_pg_rca12_fa61_y4, h_s_dadda_pg_rca12_nand_11_8_y0, h_s_dadda_pg_rca12_fa63_y2, h_s_dadda_pg_rca12_fa63_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_3_0_y0(a_3, b_0, h_s_dadda_pg_rca12_and_3_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_1_y0(a_2, b_1, h_s_dadda_pg_rca12_and_2_1_y0);
  ha ha_h_s_dadda_pg_rca12_ha8_y0(h_s_dadda_pg_rca12_and_3_0_y0, h_s_dadda_pg_rca12_and_2_1_y0, h_s_dadda_pg_rca12_ha8_y0, h_s_dadda_pg_rca12_ha8_y1);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_2_y0(a_2, b_2, h_s_dadda_pg_rca12_and_2_2_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_3_y0(a_1, b_3, h_s_dadda_pg_rca12_and_1_3_y0);
  fa fa_h_s_dadda_pg_rca12_fa64_y2(h_s_dadda_pg_rca12_ha8_y1, h_s_dadda_pg_rca12_and_2_2_y0, h_s_dadda_pg_rca12_and_1_3_y0, h_s_dadda_pg_rca12_fa64_y2, h_s_dadda_pg_rca12_fa64_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_4_y0(a_1, b_4, h_s_dadda_pg_rca12_and_1_4_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_5_y0(a_0, b_5, h_s_dadda_pg_rca12_and_0_5_y0);
  fa fa_h_s_dadda_pg_rca12_fa65_y2(h_s_dadda_pg_rca12_fa64_y4, h_s_dadda_pg_rca12_and_1_4_y0, h_s_dadda_pg_rca12_and_0_5_y0, h_s_dadda_pg_rca12_fa65_y2, h_s_dadda_pg_rca12_fa65_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_6_y0(a_0, b_6, h_s_dadda_pg_rca12_and_0_6_y0);
  fa fa_h_s_dadda_pg_rca12_fa66_y2(h_s_dadda_pg_rca12_fa65_y4, h_s_dadda_pg_rca12_and_0_6_y0, h_s_dadda_pg_rca12_fa10_y2, h_s_dadda_pg_rca12_fa66_y2, h_s_dadda_pg_rca12_fa66_y4);
  fa fa_h_s_dadda_pg_rca12_fa67_y2(h_s_dadda_pg_rca12_fa66_y4, h_s_dadda_pg_rca12_fa12_y2, h_s_dadda_pg_rca12_fa13_y2, h_s_dadda_pg_rca12_fa67_y2, h_s_dadda_pg_rca12_fa67_y4);
  fa fa_h_s_dadda_pg_rca12_fa68_y2(h_s_dadda_pg_rca12_fa67_y4, h_s_dadda_pg_rca12_fa16_y2, h_s_dadda_pg_rca12_fa17_y2, h_s_dadda_pg_rca12_fa68_y2, h_s_dadda_pg_rca12_fa68_y4);
  fa fa_h_s_dadda_pg_rca12_fa69_y2(h_s_dadda_pg_rca12_fa68_y4, h_s_dadda_pg_rca12_fa20_y2, h_s_dadda_pg_rca12_fa21_y2, h_s_dadda_pg_rca12_fa69_y2, h_s_dadda_pg_rca12_fa69_y4);
  fa fa_h_s_dadda_pg_rca12_fa70_y2(h_s_dadda_pg_rca12_fa69_y4, h_s_dadda_pg_rca12_fa25_y2, h_s_dadda_pg_rca12_fa26_y2, h_s_dadda_pg_rca12_fa70_y2, h_s_dadda_pg_rca12_fa70_y4);
  fa fa_h_s_dadda_pg_rca12_fa71_y2(h_s_dadda_pg_rca12_fa70_y4, h_s_dadda_pg_rca12_fa30_y2, h_s_dadda_pg_rca12_fa31_y2, h_s_dadda_pg_rca12_fa71_y2, h_s_dadda_pg_rca12_fa71_y4);
  fa fa_h_s_dadda_pg_rca12_fa72_y2(h_s_dadda_pg_rca12_fa71_y4, h_s_dadda_pg_rca12_fa35_y2, h_s_dadda_pg_rca12_fa36_y2, h_s_dadda_pg_rca12_fa72_y2, h_s_dadda_pg_rca12_fa72_y4);
  fa fa_h_s_dadda_pg_rca12_fa73_y2(h_s_dadda_pg_rca12_fa72_y4, h_s_dadda_pg_rca12_fa40_y2, h_s_dadda_pg_rca12_fa41_y2, h_s_dadda_pg_rca12_fa73_y2, h_s_dadda_pg_rca12_fa73_y4);
  fa fa_h_s_dadda_pg_rca12_fa74_y2(h_s_dadda_pg_rca12_fa73_y4, h_s_dadda_pg_rca12_fa45_y2, h_s_dadda_pg_rca12_fa46_y2, h_s_dadda_pg_rca12_fa74_y2, h_s_dadda_pg_rca12_fa74_y4);
  fa fa_h_s_dadda_pg_rca12_fa75_y2(h_s_dadda_pg_rca12_fa74_y4, h_s_dadda_pg_rca12_fa50_y2, h_s_dadda_pg_rca12_fa51_y2, h_s_dadda_pg_rca12_fa75_y2, h_s_dadda_pg_rca12_fa75_y4);
  fa fa_h_s_dadda_pg_rca12_fa76_y2(h_s_dadda_pg_rca12_fa75_y4, h_s_dadda_pg_rca12_fa54_y2, h_s_dadda_pg_rca12_fa55_y2, h_s_dadda_pg_rca12_fa76_y2, h_s_dadda_pg_rca12_fa76_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_6_11_y0(a_6, b_11, h_s_dadda_pg_rca12_nand_6_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa77_y2(h_s_dadda_pg_rca12_fa76_y4, h_s_dadda_pg_rca12_nand_6_11_y0, h_s_dadda_pg_rca12_fa58_y2, h_s_dadda_pg_rca12_fa77_y2, h_s_dadda_pg_rca12_fa77_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_8_10_y0(a_8, b_10, h_s_dadda_pg_rca12_and_8_10_y0);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_7_11_y0(a_7, b_11, h_s_dadda_pg_rca12_nand_7_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa78_y2(h_s_dadda_pg_rca12_fa77_y4, h_s_dadda_pg_rca12_and_8_10_y0, h_s_dadda_pg_rca12_nand_7_11_y0, h_s_dadda_pg_rca12_fa78_y2, h_s_dadda_pg_rca12_fa78_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_9_y0(a_10, b_9, h_s_dadda_pg_rca12_and_10_9_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_9_10_y0(a_9, b_10, h_s_dadda_pg_rca12_and_9_10_y0);
  fa fa_h_s_dadda_pg_rca12_fa79_y2(h_s_dadda_pg_rca12_fa78_y4, h_s_dadda_pg_rca12_and_10_9_y0, h_s_dadda_pg_rca12_and_9_10_y0, h_s_dadda_pg_rca12_fa79_y2, h_s_dadda_pg_rca12_fa79_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_9_y0(a_11, b_9, h_s_dadda_pg_rca12_nand_11_9_y0);
  fa fa_h_s_dadda_pg_rca12_fa80_y2(h_s_dadda_pg_rca12_fa79_y4, h_s_dadda_pg_rca12_fa63_y4, h_s_dadda_pg_rca12_nand_11_9_y0, h_s_dadda_pg_rca12_fa80_y2, h_s_dadda_pg_rca12_fa80_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_2_0_y0(a_2, b_0, h_s_dadda_pg_rca12_and_2_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_1_y0(a_1, b_1, h_s_dadda_pg_rca12_and_1_1_y0);
  ha ha_h_s_dadda_pg_rca12_ha9_y0(h_s_dadda_pg_rca12_and_2_0_y0, h_s_dadda_pg_rca12_and_1_1_y0, h_s_dadda_pg_rca12_ha9_y0, h_s_dadda_pg_rca12_ha9_y1);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_2_y0(a_1, b_2, h_s_dadda_pg_rca12_and_1_2_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_3_y0(a_0, b_3, h_s_dadda_pg_rca12_and_0_3_y0);
  fa fa_h_s_dadda_pg_rca12_fa81_y2(h_s_dadda_pg_rca12_ha9_y1, h_s_dadda_pg_rca12_and_1_2_y0, h_s_dadda_pg_rca12_and_0_3_y0, h_s_dadda_pg_rca12_fa81_y2, h_s_dadda_pg_rca12_fa81_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_4_y0(a_0, b_4, h_s_dadda_pg_rca12_and_0_4_y0);
  fa fa_h_s_dadda_pg_rca12_fa82_y2(h_s_dadda_pg_rca12_fa81_y4, h_s_dadda_pg_rca12_and_0_4_y0, h_s_dadda_pg_rca12_ha3_y0, h_s_dadda_pg_rca12_fa82_y2, h_s_dadda_pg_rca12_fa82_y4);
  fa fa_h_s_dadda_pg_rca12_fa83_y2(h_s_dadda_pg_rca12_fa82_y4, h_s_dadda_pg_rca12_fa9_y2, h_s_dadda_pg_rca12_ha4_y0, h_s_dadda_pg_rca12_fa83_y2, h_s_dadda_pg_rca12_fa83_y4);
  fa fa_h_s_dadda_pg_rca12_fa84_y2(h_s_dadda_pg_rca12_fa83_y4, h_s_dadda_pg_rca12_fa11_y2, h_s_dadda_pg_rca12_ha5_y0, h_s_dadda_pg_rca12_fa84_y2, h_s_dadda_pg_rca12_fa84_y4);
  fa fa_h_s_dadda_pg_rca12_fa85_y2(h_s_dadda_pg_rca12_fa84_y4, h_s_dadda_pg_rca12_fa14_y2, h_s_dadda_pg_rca12_ha6_y0, h_s_dadda_pg_rca12_fa85_y2, h_s_dadda_pg_rca12_fa85_y4);
  fa fa_h_s_dadda_pg_rca12_fa86_y2(h_s_dadda_pg_rca12_fa85_y4, h_s_dadda_pg_rca12_fa18_y2, h_s_dadda_pg_rca12_ha7_y0, h_s_dadda_pg_rca12_fa86_y2, h_s_dadda_pg_rca12_fa86_y4);
  fa fa_h_s_dadda_pg_rca12_fa87_y2(h_s_dadda_pg_rca12_fa86_y4, h_s_dadda_pg_rca12_fa22_y2, h_s_dadda_pg_rca12_fa23_y2, h_s_dadda_pg_rca12_fa87_y2, h_s_dadda_pg_rca12_fa87_y4);
  fa fa_h_s_dadda_pg_rca12_fa88_y2(h_s_dadda_pg_rca12_fa87_y4, h_s_dadda_pg_rca12_fa27_y2, h_s_dadda_pg_rca12_fa28_y2, h_s_dadda_pg_rca12_fa88_y2, h_s_dadda_pg_rca12_fa88_y4);
  fa fa_h_s_dadda_pg_rca12_fa89_y2(h_s_dadda_pg_rca12_fa88_y4, h_s_dadda_pg_rca12_fa32_y2, h_s_dadda_pg_rca12_fa33_y2, h_s_dadda_pg_rca12_fa89_y2, h_s_dadda_pg_rca12_fa89_y4);
  fa fa_h_s_dadda_pg_rca12_fa90_y2(h_s_dadda_pg_rca12_fa89_y4, h_s_dadda_pg_rca12_fa37_y2, h_s_dadda_pg_rca12_fa38_y2, h_s_dadda_pg_rca12_fa90_y2, h_s_dadda_pg_rca12_fa90_y4);
  fa fa_h_s_dadda_pg_rca12_fa91_y2(h_s_dadda_pg_rca12_fa90_y4, h_s_dadda_pg_rca12_fa42_y2, h_s_dadda_pg_rca12_fa43_y2, h_s_dadda_pg_rca12_fa91_y2, h_s_dadda_pg_rca12_fa91_y4);
  fa fa_h_s_dadda_pg_rca12_fa92_y2(h_s_dadda_pg_rca12_fa91_y4, h_s_dadda_pg_rca12_fa47_y2, h_s_dadda_pg_rca12_fa48_y2, h_s_dadda_pg_rca12_fa92_y2, h_s_dadda_pg_rca12_fa92_y4);
  fa fa_h_s_dadda_pg_rca12_fa93_y2(h_s_dadda_pg_rca12_fa92_y4, h_s_dadda_pg_rca12_fa52_y2, h_s_dadda_pg_rca12_fa53_y2, h_s_dadda_pg_rca12_fa93_y2, h_s_dadda_pg_rca12_fa93_y4);
  fa fa_h_s_dadda_pg_rca12_fa94_y2(h_s_dadda_pg_rca12_fa93_y4, h_s_dadda_pg_rca12_fa56_y2, h_s_dadda_pg_rca12_fa57_y2, h_s_dadda_pg_rca12_fa94_y2, h_s_dadda_pg_rca12_fa94_y4);
  fa fa_h_s_dadda_pg_rca12_fa95_y2(h_s_dadda_pg_rca12_fa94_y4, h_s_dadda_pg_rca12_fa59_y2, h_s_dadda_pg_rca12_fa60_y2, h_s_dadda_pg_rca12_fa95_y2, h_s_dadda_pg_rca12_fa95_y4);
  fa fa_h_s_dadda_pg_rca12_fa96_y2(h_s_dadda_pg_rca12_fa95_y4, h_s_dadda_pg_rca12_fa61_y2, h_s_dadda_pg_rca12_fa62_y2, h_s_dadda_pg_rca12_fa96_y2, h_s_dadda_pg_rca12_fa96_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_8_11_y0(a_8, b_11, h_s_dadda_pg_rca12_nand_8_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa97_y2(h_s_dadda_pg_rca12_fa96_y4, h_s_dadda_pg_rca12_nand_8_11_y0, h_s_dadda_pg_rca12_fa63_y2, h_s_dadda_pg_rca12_fa97_y2, h_s_dadda_pg_rca12_fa97_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_10_10_y0(a_10, b_10, h_s_dadda_pg_rca12_and_10_10_y0);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_9_11_y0(a_9, b_11, h_s_dadda_pg_rca12_nand_9_11_y0);
  fa fa_h_s_dadda_pg_rca12_fa98_y2(h_s_dadda_pg_rca12_fa97_y4, h_s_dadda_pg_rca12_and_10_10_y0, h_s_dadda_pg_rca12_nand_9_11_y0, h_s_dadda_pg_rca12_fa98_y2, h_s_dadda_pg_rca12_fa98_y4);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_11_10_y0(a_11, b_10, h_s_dadda_pg_rca12_nand_11_10_y0);
  fa fa_h_s_dadda_pg_rca12_fa99_y2(h_s_dadda_pg_rca12_fa98_y4, h_s_dadda_pg_rca12_fa80_y4, h_s_dadda_pg_rca12_nand_11_10_y0, h_s_dadda_pg_rca12_fa99_y2, h_s_dadda_pg_rca12_fa99_y4);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_0_y0(a_0, b_0, h_s_dadda_pg_rca12_and_0_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_1_0_y0(a_1, b_0, h_s_dadda_pg_rca12_and_1_0_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_2_y0(a_0, b_2, h_s_dadda_pg_rca12_and_0_2_y0);
  nand_gate nand_gate_h_s_dadda_pg_rca12_nand_10_11_y0(a_10, b_11, h_s_dadda_pg_rca12_nand_10_11_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_0_1_y0(a_0, b_1, h_s_dadda_pg_rca12_and_0_1_y0);
  and_gate and_gate_h_s_dadda_pg_rca12_and_11_11_y0(a_11, b_11, h_s_dadda_pg_rca12_and_11_11_y0);
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[0] = h_s_dadda_pg_rca12_and_1_0_y0;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[1] = h_s_dadda_pg_rca12_and_0_2_y0;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[2] = h_s_dadda_pg_rca12_ha8_y0;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[3] = h_s_dadda_pg_rca12_fa64_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[4] = h_s_dadda_pg_rca12_fa65_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[5] = h_s_dadda_pg_rca12_fa66_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[6] = h_s_dadda_pg_rca12_fa67_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[7] = h_s_dadda_pg_rca12_fa68_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[8] = h_s_dadda_pg_rca12_fa69_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[9] = h_s_dadda_pg_rca12_fa70_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[10] = h_s_dadda_pg_rca12_fa71_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[11] = h_s_dadda_pg_rca12_fa72_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[12] = h_s_dadda_pg_rca12_fa73_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[13] = h_s_dadda_pg_rca12_fa74_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[14] = h_s_dadda_pg_rca12_fa75_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[15] = h_s_dadda_pg_rca12_fa76_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[16] = h_s_dadda_pg_rca12_fa77_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[17] = h_s_dadda_pg_rca12_fa78_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[18] = h_s_dadda_pg_rca12_fa79_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[19] = h_s_dadda_pg_rca12_fa80_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[20] = h_s_dadda_pg_rca12_nand_10_11_y0;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a[21] = h_s_dadda_pg_rca12_fa99_y4;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[0] = h_s_dadda_pg_rca12_and_0_1_y0;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[1] = h_s_dadda_pg_rca12_ha9_y0;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[2] = h_s_dadda_pg_rca12_fa81_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[3] = h_s_dadda_pg_rca12_fa82_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[4] = h_s_dadda_pg_rca12_fa83_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[5] = h_s_dadda_pg_rca12_fa84_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[6] = h_s_dadda_pg_rca12_fa85_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[7] = h_s_dadda_pg_rca12_fa86_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[8] = h_s_dadda_pg_rca12_fa87_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[9] = h_s_dadda_pg_rca12_fa88_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[10] = h_s_dadda_pg_rca12_fa89_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[11] = h_s_dadda_pg_rca12_fa90_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[12] = h_s_dadda_pg_rca12_fa91_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[13] = h_s_dadda_pg_rca12_fa92_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[14] = h_s_dadda_pg_rca12_fa93_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[15] = h_s_dadda_pg_rca12_fa94_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[16] = h_s_dadda_pg_rca12_fa95_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[17] = h_s_dadda_pg_rca12_fa96_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[18] = h_s_dadda_pg_rca12_fa97_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[19] = h_s_dadda_pg_rca12_fa98_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[20] = h_s_dadda_pg_rca12_fa99_y2;
  assign h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b[21] = h_s_dadda_pg_rca12_and_11_11_y0;
  u_pg_rca u_pg_rca_out(h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_a, h_s_dadda_pg_rca12_u_pg_rca_u_pg_rca_b, h_s_dadda_pg_rca12_u_pg_rca_out);
  assign h_s_dadda_pg_rca12_u_pg_rca_fa0_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[0];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa1_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[1];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa2_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[2];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa3_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[3];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa4_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[4];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa5_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[5];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa6_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[6];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa7_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[7];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa8_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[8];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa9_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[9];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa10_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[10];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa11_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[11];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa12_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[12];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa13_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[13];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa14_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[14];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa15_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[15];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa16_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[16];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa17_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[17];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa18_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[18];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa19_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[19];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa20_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[20];
  assign h_s_dadda_pg_rca12_u_pg_rca_fa21_y2 = h_s_dadda_pg_rca12_u_pg_rca_out[21];
  assign h_s_dadda_pg_rca12_u_pg_rca_or21_y0 = h_s_dadda_pg_rca12_u_pg_rca_out[22];
  xor_gate xor_gate_h_s_dadda_pg_rca12_xor0_y0(constant_wire_1, h_s_dadda_pg_rca12_u_pg_rca_or21_y0, h_s_dadda_pg_rca12_xor0_y0);

  assign out[0] = h_s_dadda_pg_rca12_and_0_0_y0;
  assign out[1] = h_s_dadda_pg_rca12_u_pg_rca_fa0_y2;
  assign out[2] = h_s_dadda_pg_rca12_u_pg_rca_fa1_y2;
  assign out[3] = h_s_dadda_pg_rca12_u_pg_rca_fa2_y2;
  assign out[4] = h_s_dadda_pg_rca12_u_pg_rca_fa3_y2;
  assign out[5] = h_s_dadda_pg_rca12_u_pg_rca_fa4_y2;
  assign out[6] = h_s_dadda_pg_rca12_u_pg_rca_fa5_y2;
  assign out[7] = h_s_dadda_pg_rca12_u_pg_rca_fa6_y2;
  assign out[8] = h_s_dadda_pg_rca12_u_pg_rca_fa7_y2;
  assign out[9] = h_s_dadda_pg_rca12_u_pg_rca_fa8_y2;
  assign out[10] = h_s_dadda_pg_rca12_u_pg_rca_fa9_y2;
  assign out[11] = h_s_dadda_pg_rca12_u_pg_rca_fa10_y2;
  assign out[12] = h_s_dadda_pg_rca12_u_pg_rca_fa11_y2;
  assign out[13] = h_s_dadda_pg_rca12_u_pg_rca_fa12_y2;
  assign out[14] = h_s_dadda_pg_rca12_u_pg_rca_fa13_y2;
  assign out[15] = h_s_dadda_pg_rca12_u_pg_rca_fa14_y2;
  assign out[16] = h_s_dadda_pg_rca12_u_pg_rca_fa15_y2;
  assign out[17] = h_s_dadda_pg_rca12_u_pg_rca_fa16_y2;
  assign out[18] = h_s_dadda_pg_rca12_u_pg_rca_fa17_y2;
  assign out[19] = h_s_dadda_pg_rca12_u_pg_rca_fa18_y2;
  assign out[20] = h_s_dadda_pg_rca12_u_pg_rca_fa19_y2;
  assign out[21] = h_s_dadda_pg_rca12_u_pg_rca_fa20_y2;
  assign out[22] = h_s_dadda_pg_rca12_u_pg_rca_fa21_y2;
  assign out[23] = h_s_dadda_pg_rca12_xor0_y0;
endmodule