module f_u_cla12(input [11:0] a, input [11:0] b, output [12:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire constant_wire_value_0_a_0;
  wire constant_wire_value_0_b_0;
  wire constant_wire_value_0_y0;
  wire constant_wire_value_0_y1;
  wire constant_wire_0;
  wire f_u_cla12_pg_logic0_a_0;
  wire f_u_cla12_pg_logic0_b_0;
  wire f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_pg_logic0_y2;
  wire f_u_cla12_xor0_f_u_cla12_pg_logic0_y2;
  wire f_u_cla12_xor0_constant_wire_0;
  wire f_u_cla12_xor0_y0;
  wire f_u_cla12_and0_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and0_constant_wire_0;
  wire f_u_cla12_and0_y0;
  wire f_u_cla12_or0_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_or0_f_u_cla12_and0_y0;
  wire f_u_cla12_or0_y0;
  wire f_u_cla12_pg_logic1_a_1;
  wire f_u_cla12_pg_logic1_b_1;
  wire f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_pg_logic1_y2;
  wire f_u_cla12_xor1_f_u_cla12_pg_logic1_y2;
  wire f_u_cla12_xor1_f_u_cla12_or0_y0;
  wire f_u_cla12_xor1_y0;
  wire f_u_cla12_and1_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and1_constant_wire_0;
  wire f_u_cla12_and1_y0;
  wire f_u_cla12_and2_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and2_constant_wire_0;
  wire f_u_cla12_and2_y0;
  wire f_u_cla12_and3_f_u_cla12_and2_y0;
  wire f_u_cla12_and3_f_u_cla12_and1_y0;
  wire f_u_cla12_and3_y0;
  wire f_u_cla12_and4_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and4_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and4_y0;
  wire f_u_cla12_or1_f_u_cla12_and4_y0;
  wire f_u_cla12_or1_f_u_cla12_and3_y0;
  wire f_u_cla12_or1_y0;
  wire f_u_cla12_or2_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_or2_f_u_cla12_or1_y0;
  wire f_u_cla12_or2_y0;
  wire f_u_cla12_pg_logic2_a_2;
  wire f_u_cla12_pg_logic2_b_2;
  wire f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_pg_logic2_y2;
  wire f_u_cla12_xor2_f_u_cla12_pg_logic2_y2;
  wire f_u_cla12_xor2_f_u_cla12_or2_y0;
  wire f_u_cla12_xor2_y0;
  wire f_u_cla12_and5_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and5_constant_wire_0;
  wire f_u_cla12_and5_y0;
  wire f_u_cla12_and6_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and6_constant_wire_0;
  wire f_u_cla12_and6_y0;
  wire f_u_cla12_and7_f_u_cla12_and6_y0;
  wire f_u_cla12_and7_f_u_cla12_and5_y0;
  wire f_u_cla12_and7_y0;
  wire f_u_cla12_and8_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and8_constant_wire_0;
  wire f_u_cla12_and8_y0;
  wire f_u_cla12_and9_f_u_cla12_and8_y0;
  wire f_u_cla12_and9_f_u_cla12_and7_y0;
  wire f_u_cla12_and9_y0;
  wire f_u_cla12_and10_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and10_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and10_y0;
  wire f_u_cla12_and11_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and11_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and11_y0;
  wire f_u_cla12_and12_f_u_cla12_and11_y0;
  wire f_u_cla12_and12_f_u_cla12_and10_y0;
  wire f_u_cla12_and12_y0;
  wire f_u_cla12_and13_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and13_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and13_y0;
  wire f_u_cla12_or3_f_u_cla12_and13_y0;
  wire f_u_cla12_or3_f_u_cla12_and9_y0;
  wire f_u_cla12_or3_y0;
  wire f_u_cla12_or4_f_u_cla12_or3_y0;
  wire f_u_cla12_or4_f_u_cla12_and12_y0;
  wire f_u_cla12_or4_y0;
  wire f_u_cla12_or5_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_or5_f_u_cla12_or4_y0;
  wire f_u_cla12_or5_y0;
  wire f_u_cla12_pg_logic3_a_3;
  wire f_u_cla12_pg_logic3_b_3;
  wire f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_pg_logic3_y2;
  wire f_u_cla12_xor3_f_u_cla12_pg_logic3_y2;
  wire f_u_cla12_xor3_f_u_cla12_or5_y0;
  wire f_u_cla12_xor3_y0;
  wire f_u_cla12_and14_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and14_constant_wire_0;
  wire f_u_cla12_and14_y0;
  wire f_u_cla12_and15_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and15_constant_wire_0;
  wire f_u_cla12_and15_y0;
  wire f_u_cla12_and16_f_u_cla12_and15_y0;
  wire f_u_cla12_and16_f_u_cla12_and14_y0;
  wire f_u_cla12_and16_y0;
  wire f_u_cla12_and17_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and17_constant_wire_0;
  wire f_u_cla12_and17_y0;
  wire f_u_cla12_and18_f_u_cla12_and17_y0;
  wire f_u_cla12_and18_f_u_cla12_and16_y0;
  wire f_u_cla12_and18_y0;
  wire f_u_cla12_and19_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and19_constant_wire_0;
  wire f_u_cla12_and19_y0;
  wire f_u_cla12_and20_f_u_cla12_and19_y0;
  wire f_u_cla12_and20_f_u_cla12_and18_y0;
  wire f_u_cla12_and20_y0;
  wire f_u_cla12_and21_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and21_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and21_y0;
  wire f_u_cla12_and22_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and22_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and22_y0;
  wire f_u_cla12_and23_f_u_cla12_and22_y0;
  wire f_u_cla12_and23_f_u_cla12_and21_y0;
  wire f_u_cla12_and23_y0;
  wire f_u_cla12_and24_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and24_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and24_y0;
  wire f_u_cla12_and25_f_u_cla12_and24_y0;
  wire f_u_cla12_and25_f_u_cla12_and23_y0;
  wire f_u_cla12_and25_y0;
  wire f_u_cla12_and26_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and26_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and26_y0;
  wire f_u_cla12_and27_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and27_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and27_y0;
  wire f_u_cla12_and28_f_u_cla12_and27_y0;
  wire f_u_cla12_and28_f_u_cla12_and26_y0;
  wire f_u_cla12_and28_y0;
  wire f_u_cla12_and29_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and29_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and29_y0;
  wire f_u_cla12_or6_f_u_cla12_and29_y0;
  wire f_u_cla12_or6_f_u_cla12_and20_y0;
  wire f_u_cla12_or6_y0;
  wire f_u_cla12_or7_f_u_cla12_or6_y0;
  wire f_u_cla12_or7_f_u_cla12_and25_y0;
  wire f_u_cla12_or7_y0;
  wire f_u_cla12_or8_f_u_cla12_or7_y0;
  wire f_u_cla12_or8_f_u_cla12_and28_y0;
  wire f_u_cla12_or8_y0;
  wire f_u_cla12_or9_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_or9_f_u_cla12_or8_y0;
  wire f_u_cla12_or9_y0;
  wire f_u_cla12_pg_logic4_a_4;
  wire f_u_cla12_pg_logic4_b_4;
  wire f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_pg_logic4_y2;
  wire f_u_cla12_xor4_f_u_cla12_pg_logic4_y2;
  wire f_u_cla12_xor4_f_u_cla12_or9_y0;
  wire f_u_cla12_xor4_y0;
  wire f_u_cla12_and30_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and30_constant_wire_0;
  wire f_u_cla12_and30_y0;
  wire f_u_cla12_and31_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and31_constant_wire_0;
  wire f_u_cla12_and31_y0;
  wire f_u_cla12_and32_f_u_cla12_and31_y0;
  wire f_u_cla12_and32_f_u_cla12_and30_y0;
  wire f_u_cla12_and32_y0;
  wire f_u_cla12_and33_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and33_constant_wire_0;
  wire f_u_cla12_and33_y0;
  wire f_u_cla12_and34_f_u_cla12_and33_y0;
  wire f_u_cla12_and34_f_u_cla12_and32_y0;
  wire f_u_cla12_and34_y0;
  wire f_u_cla12_and35_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and35_constant_wire_0;
  wire f_u_cla12_and35_y0;
  wire f_u_cla12_and36_f_u_cla12_and35_y0;
  wire f_u_cla12_and36_f_u_cla12_and34_y0;
  wire f_u_cla12_and36_y0;
  wire f_u_cla12_and37_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and37_constant_wire_0;
  wire f_u_cla12_and37_y0;
  wire f_u_cla12_and38_f_u_cla12_and37_y0;
  wire f_u_cla12_and38_f_u_cla12_and36_y0;
  wire f_u_cla12_and38_y0;
  wire f_u_cla12_and39_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and39_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and39_y0;
  wire f_u_cla12_and40_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and40_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and40_y0;
  wire f_u_cla12_and41_f_u_cla12_and40_y0;
  wire f_u_cla12_and41_f_u_cla12_and39_y0;
  wire f_u_cla12_and41_y0;
  wire f_u_cla12_and42_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and42_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and42_y0;
  wire f_u_cla12_and43_f_u_cla12_and42_y0;
  wire f_u_cla12_and43_f_u_cla12_and41_y0;
  wire f_u_cla12_and43_y0;
  wire f_u_cla12_and44_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and44_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and44_y0;
  wire f_u_cla12_and45_f_u_cla12_and44_y0;
  wire f_u_cla12_and45_f_u_cla12_and43_y0;
  wire f_u_cla12_and45_y0;
  wire f_u_cla12_and46_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and46_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and46_y0;
  wire f_u_cla12_and47_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and47_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and47_y0;
  wire f_u_cla12_and48_f_u_cla12_and47_y0;
  wire f_u_cla12_and48_f_u_cla12_and46_y0;
  wire f_u_cla12_and48_y0;
  wire f_u_cla12_and49_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and49_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and49_y0;
  wire f_u_cla12_and50_f_u_cla12_and49_y0;
  wire f_u_cla12_and50_f_u_cla12_and48_y0;
  wire f_u_cla12_and50_y0;
  wire f_u_cla12_and51_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and51_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and51_y0;
  wire f_u_cla12_and52_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and52_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and52_y0;
  wire f_u_cla12_and53_f_u_cla12_and52_y0;
  wire f_u_cla12_and53_f_u_cla12_and51_y0;
  wire f_u_cla12_and53_y0;
  wire f_u_cla12_and54_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and54_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and54_y0;
  wire f_u_cla12_or10_f_u_cla12_and54_y0;
  wire f_u_cla12_or10_f_u_cla12_and38_y0;
  wire f_u_cla12_or10_y0;
  wire f_u_cla12_or11_f_u_cla12_or10_y0;
  wire f_u_cla12_or11_f_u_cla12_and45_y0;
  wire f_u_cla12_or11_y0;
  wire f_u_cla12_or12_f_u_cla12_or11_y0;
  wire f_u_cla12_or12_f_u_cla12_and50_y0;
  wire f_u_cla12_or12_y0;
  wire f_u_cla12_or13_f_u_cla12_or12_y0;
  wire f_u_cla12_or13_f_u_cla12_and53_y0;
  wire f_u_cla12_or13_y0;
  wire f_u_cla12_or14_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_or14_f_u_cla12_or13_y0;
  wire f_u_cla12_or14_y0;
  wire f_u_cla12_pg_logic5_a_5;
  wire f_u_cla12_pg_logic5_b_5;
  wire f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_pg_logic5_y2;
  wire f_u_cla12_xor5_f_u_cla12_pg_logic5_y2;
  wire f_u_cla12_xor5_f_u_cla12_or14_y0;
  wire f_u_cla12_xor5_y0;
  wire f_u_cla12_and55_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and55_constant_wire_0;
  wire f_u_cla12_and55_y0;
  wire f_u_cla12_and56_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and56_constant_wire_0;
  wire f_u_cla12_and56_y0;
  wire f_u_cla12_and57_f_u_cla12_and56_y0;
  wire f_u_cla12_and57_f_u_cla12_and55_y0;
  wire f_u_cla12_and57_y0;
  wire f_u_cla12_and58_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and58_constant_wire_0;
  wire f_u_cla12_and58_y0;
  wire f_u_cla12_and59_f_u_cla12_and58_y0;
  wire f_u_cla12_and59_f_u_cla12_and57_y0;
  wire f_u_cla12_and59_y0;
  wire f_u_cla12_and60_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and60_constant_wire_0;
  wire f_u_cla12_and60_y0;
  wire f_u_cla12_and61_f_u_cla12_and60_y0;
  wire f_u_cla12_and61_f_u_cla12_and59_y0;
  wire f_u_cla12_and61_y0;
  wire f_u_cla12_and62_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and62_constant_wire_0;
  wire f_u_cla12_and62_y0;
  wire f_u_cla12_and63_f_u_cla12_and62_y0;
  wire f_u_cla12_and63_f_u_cla12_and61_y0;
  wire f_u_cla12_and63_y0;
  wire f_u_cla12_and64_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and64_constant_wire_0;
  wire f_u_cla12_and64_y0;
  wire f_u_cla12_and65_f_u_cla12_and64_y0;
  wire f_u_cla12_and65_f_u_cla12_and63_y0;
  wire f_u_cla12_and65_y0;
  wire f_u_cla12_and66_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and66_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and66_y0;
  wire f_u_cla12_and67_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and67_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and67_y0;
  wire f_u_cla12_and68_f_u_cla12_and67_y0;
  wire f_u_cla12_and68_f_u_cla12_and66_y0;
  wire f_u_cla12_and68_y0;
  wire f_u_cla12_and69_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and69_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and69_y0;
  wire f_u_cla12_and70_f_u_cla12_and69_y0;
  wire f_u_cla12_and70_f_u_cla12_and68_y0;
  wire f_u_cla12_and70_y0;
  wire f_u_cla12_and71_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and71_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and71_y0;
  wire f_u_cla12_and72_f_u_cla12_and71_y0;
  wire f_u_cla12_and72_f_u_cla12_and70_y0;
  wire f_u_cla12_and72_y0;
  wire f_u_cla12_and73_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and73_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and73_y0;
  wire f_u_cla12_and74_f_u_cla12_and73_y0;
  wire f_u_cla12_and74_f_u_cla12_and72_y0;
  wire f_u_cla12_and74_y0;
  wire f_u_cla12_and75_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and75_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and75_y0;
  wire f_u_cla12_and76_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and76_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and76_y0;
  wire f_u_cla12_and77_f_u_cla12_and76_y0;
  wire f_u_cla12_and77_f_u_cla12_and75_y0;
  wire f_u_cla12_and77_y0;
  wire f_u_cla12_and78_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and78_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and78_y0;
  wire f_u_cla12_and79_f_u_cla12_and78_y0;
  wire f_u_cla12_and79_f_u_cla12_and77_y0;
  wire f_u_cla12_and79_y0;
  wire f_u_cla12_and80_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and80_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and80_y0;
  wire f_u_cla12_and81_f_u_cla12_and80_y0;
  wire f_u_cla12_and81_f_u_cla12_and79_y0;
  wire f_u_cla12_and81_y0;
  wire f_u_cla12_and82_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and82_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and82_y0;
  wire f_u_cla12_and83_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and83_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and83_y0;
  wire f_u_cla12_and84_f_u_cla12_and83_y0;
  wire f_u_cla12_and84_f_u_cla12_and82_y0;
  wire f_u_cla12_and84_y0;
  wire f_u_cla12_and85_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and85_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and85_y0;
  wire f_u_cla12_and86_f_u_cla12_and85_y0;
  wire f_u_cla12_and86_f_u_cla12_and84_y0;
  wire f_u_cla12_and86_y0;
  wire f_u_cla12_and87_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and87_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and87_y0;
  wire f_u_cla12_and88_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and88_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and88_y0;
  wire f_u_cla12_and89_f_u_cla12_and88_y0;
  wire f_u_cla12_and89_f_u_cla12_and87_y0;
  wire f_u_cla12_and89_y0;
  wire f_u_cla12_and90_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and90_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and90_y0;
  wire f_u_cla12_or15_f_u_cla12_and90_y0;
  wire f_u_cla12_or15_f_u_cla12_and65_y0;
  wire f_u_cla12_or15_y0;
  wire f_u_cla12_or16_f_u_cla12_or15_y0;
  wire f_u_cla12_or16_f_u_cla12_and74_y0;
  wire f_u_cla12_or16_y0;
  wire f_u_cla12_or17_f_u_cla12_or16_y0;
  wire f_u_cla12_or17_f_u_cla12_and81_y0;
  wire f_u_cla12_or17_y0;
  wire f_u_cla12_or18_f_u_cla12_or17_y0;
  wire f_u_cla12_or18_f_u_cla12_and86_y0;
  wire f_u_cla12_or18_y0;
  wire f_u_cla12_or19_f_u_cla12_or18_y0;
  wire f_u_cla12_or19_f_u_cla12_and89_y0;
  wire f_u_cla12_or19_y0;
  wire f_u_cla12_or20_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_or20_f_u_cla12_or19_y0;
  wire f_u_cla12_or20_y0;
  wire f_u_cla12_pg_logic6_a_6;
  wire f_u_cla12_pg_logic6_b_6;
  wire f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_pg_logic6_y2;
  wire f_u_cla12_xor6_f_u_cla12_pg_logic6_y2;
  wire f_u_cla12_xor6_f_u_cla12_or20_y0;
  wire f_u_cla12_xor6_y0;
  wire f_u_cla12_and91_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and91_constant_wire_0;
  wire f_u_cla12_and91_y0;
  wire f_u_cla12_and92_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and92_constant_wire_0;
  wire f_u_cla12_and92_y0;
  wire f_u_cla12_and93_f_u_cla12_and92_y0;
  wire f_u_cla12_and93_f_u_cla12_and91_y0;
  wire f_u_cla12_and93_y0;
  wire f_u_cla12_and94_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and94_constant_wire_0;
  wire f_u_cla12_and94_y0;
  wire f_u_cla12_and95_f_u_cla12_and94_y0;
  wire f_u_cla12_and95_f_u_cla12_and93_y0;
  wire f_u_cla12_and95_y0;
  wire f_u_cla12_and96_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and96_constant_wire_0;
  wire f_u_cla12_and96_y0;
  wire f_u_cla12_and97_f_u_cla12_and96_y0;
  wire f_u_cla12_and97_f_u_cla12_and95_y0;
  wire f_u_cla12_and97_y0;
  wire f_u_cla12_and98_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and98_constant_wire_0;
  wire f_u_cla12_and98_y0;
  wire f_u_cla12_and99_f_u_cla12_and98_y0;
  wire f_u_cla12_and99_f_u_cla12_and97_y0;
  wire f_u_cla12_and99_y0;
  wire f_u_cla12_and100_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and100_constant_wire_0;
  wire f_u_cla12_and100_y0;
  wire f_u_cla12_and101_f_u_cla12_and100_y0;
  wire f_u_cla12_and101_f_u_cla12_and99_y0;
  wire f_u_cla12_and101_y0;
  wire f_u_cla12_and102_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and102_constant_wire_0;
  wire f_u_cla12_and102_y0;
  wire f_u_cla12_and103_f_u_cla12_and102_y0;
  wire f_u_cla12_and103_f_u_cla12_and101_y0;
  wire f_u_cla12_and103_y0;
  wire f_u_cla12_and104_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and104_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and104_y0;
  wire f_u_cla12_and105_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and105_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and105_y0;
  wire f_u_cla12_and106_f_u_cla12_and105_y0;
  wire f_u_cla12_and106_f_u_cla12_and104_y0;
  wire f_u_cla12_and106_y0;
  wire f_u_cla12_and107_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and107_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and107_y0;
  wire f_u_cla12_and108_f_u_cla12_and107_y0;
  wire f_u_cla12_and108_f_u_cla12_and106_y0;
  wire f_u_cla12_and108_y0;
  wire f_u_cla12_and109_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and109_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and109_y0;
  wire f_u_cla12_and110_f_u_cla12_and109_y0;
  wire f_u_cla12_and110_f_u_cla12_and108_y0;
  wire f_u_cla12_and110_y0;
  wire f_u_cla12_and111_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and111_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and111_y0;
  wire f_u_cla12_and112_f_u_cla12_and111_y0;
  wire f_u_cla12_and112_f_u_cla12_and110_y0;
  wire f_u_cla12_and112_y0;
  wire f_u_cla12_and113_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and113_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and113_y0;
  wire f_u_cla12_and114_f_u_cla12_and113_y0;
  wire f_u_cla12_and114_f_u_cla12_and112_y0;
  wire f_u_cla12_and114_y0;
  wire f_u_cla12_and115_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and115_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and115_y0;
  wire f_u_cla12_and116_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and116_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and116_y0;
  wire f_u_cla12_and117_f_u_cla12_and116_y0;
  wire f_u_cla12_and117_f_u_cla12_and115_y0;
  wire f_u_cla12_and117_y0;
  wire f_u_cla12_and118_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and118_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and118_y0;
  wire f_u_cla12_and119_f_u_cla12_and118_y0;
  wire f_u_cla12_and119_f_u_cla12_and117_y0;
  wire f_u_cla12_and119_y0;
  wire f_u_cla12_and120_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and120_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and120_y0;
  wire f_u_cla12_and121_f_u_cla12_and120_y0;
  wire f_u_cla12_and121_f_u_cla12_and119_y0;
  wire f_u_cla12_and121_y0;
  wire f_u_cla12_and122_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and122_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and122_y0;
  wire f_u_cla12_and123_f_u_cla12_and122_y0;
  wire f_u_cla12_and123_f_u_cla12_and121_y0;
  wire f_u_cla12_and123_y0;
  wire f_u_cla12_and124_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and124_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and124_y0;
  wire f_u_cla12_and125_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and125_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and125_y0;
  wire f_u_cla12_and126_f_u_cla12_and125_y0;
  wire f_u_cla12_and126_f_u_cla12_and124_y0;
  wire f_u_cla12_and126_y0;
  wire f_u_cla12_and127_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and127_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and127_y0;
  wire f_u_cla12_and128_f_u_cla12_and127_y0;
  wire f_u_cla12_and128_f_u_cla12_and126_y0;
  wire f_u_cla12_and128_y0;
  wire f_u_cla12_and129_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and129_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and129_y0;
  wire f_u_cla12_and130_f_u_cla12_and129_y0;
  wire f_u_cla12_and130_f_u_cla12_and128_y0;
  wire f_u_cla12_and130_y0;
  wire f_u_cla12_and131_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and131_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and131_y0;
  wire f_u_cla12_and132_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and132_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and132_y0;
  wire f_u_cla12_and133_f_u_cla12_and132_y0;
  wire f_u_cla12_and133_f_u_cla12_and131_y0;
  wire f_u_cla12_and133_y0;
  wire f_u_cla12_and134_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and134_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and134_y0;
  wire f_u_cla12_and135_f_u_cla12_and134_y0;
  wire f_u_cla12_and135_f_u_cla12_and133_y0;
  wire f_u_cla12_and135_y0;
  wire f_u_cla12_and136_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and136_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and136_y0;
  wire f_u_cla12_and137_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and137_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and137_y0;
  wire f_u_cla12_and138_f_u_cla12_and137_y0;
  wire f_u_cla12_and138_f_u_cla12_and136_y0;
  wire f_u_cla12_and138_y0;
  wire f_u_cla12_and139_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and139_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and139_y0;
  wire f_u_cla12_or21_f_u_cla12_and139_y0;
  wire f_u_cla12_or21_f_u_cla12_and103_y0;
  wire f_u_cla12_or21_y0;
  wire f_u_cla12_or22_f_u_cla12_or21_y0;
  wire f_u_cla12_or22_f_u_cla12_and114_y0;
  wire f_u_cla12_or22_y0;
  wire f_u_cla12_or23_f_u_cla12_or22_y0;
  wire f_u_cla12_or23_f_u_cla12_and123_y0;
  wire f_u_cla12_or23_y0;
  wire f_u_cla12_or24_f_u_cla12_or23_y0;
  wire f_u_cla12_or24_f_u_cla12_and130_y0;
  wire f_u_cla12_or24_y0;
  wire f_u_cla12_or25_f_u_cla12_or24_y0;
  wire f_u_cla12_or25_f_u_cla12_and135_y0;
  wire f_u_cla12_or25_y0;
  wire f_u_cla12_or26_f_u_cla12_or25_y0;
  wire f_u_cla12_or26_f_u_cla12_and138_y0;
  wire f_u_cla12_or26_y0;
  wire f_u_cla12_or27_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_or27_f_u_cla12_or26_y0;
  wire f_u_cla12_or27_y0;
  wire f_u_cla12_pg_logic7_a_7;
  wire f_u_cla12_pg_logic7_b_7;
  wire f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_pg_logic7_y2;
  wire f_u_cla12_xor7_f_u_cla12_pg_logic7_y2;
  wire f_u_cla12_xor7_f_u_cla12_or27_y0;
  wire f_u_cla12_xor7_y0;
  wire f_u_cla12_and140_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and140_constant_wire_0;
  wire f_u_cla12_and140_y0;
  wire f_u_cla12_and141_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and141_constant_wire_0;
  wire f_u_cla12_and141_y0;
  wire f_u_cla12_and142_f_u_cla12_and141_y0;
  wire f_u_cla12_and142_f_u_cla12_and140_y0;
  wire f_u_cla12_and142_y0;
  wire f_u_cla12_and143_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and143_constant_wire_0;
  wire f_u_cla12_and143_y0;
  wire f_u_cla12_and144_f_u_cla12_and143_y0;
  wire f_u_cla12_and144_f_u_cla12_and142_y0;
  wire f_u_cla12_and144_y0;
  wire f_u_cla12_and145_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and145_constant_wire_0;
  wire f_u_cla12_and145_y0;
  wire f_u_cla12_and146_f_u_cla12_and145_y0;
  wire f_u_cla12_and146_f_u_cla12_and144_y0;
  wire f_u_cla12_and146_y0;
  wire f_u_cla12_and147_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and147_constant_wire_0;
  wire f_u_cla12_and147_y0;
  wire f_u_cla12_and148_f_u_cla12_and147_y0;
  wire f_u_cla12_and148_f_u_cla12_and146_y0;
  wire f_u_cla12_and148_y0;
  wire f_u_cla12_and149_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and149_constant_wire_0;
  wire f_u_cla12_and149_y0;
  wire f_u_cla12_and150_f_u_cla12_and149_y0;
  wire f_u_cla12_and150_f_u_cla12_and148_y0;
  wire f_u_cla12_and150_y0;
  wire f_u_cla12_and151_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and151_constant_wire_0;
  wire f_u_cla12_and151_y0;
  wire f_u_cla12_and152_f_u_cla12_and151_y0;
  wire f_u_cla12_and152_f_u_cla12_and150_y0;
  wire f_u_cla12_and152_y0;
  wire f_u_cla12_and153_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and153_constant_wire_0;
  wire f_u_cla12_and153_y0;
  wire f_u_cla12_and154_f_u_cla12_and153_y0;
  wire f_u_cla12_and154_f_u_cla12_and152_y0;
  wire f_u_cla12_and154_y0;
  wire f_u_cla12_and155_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and155_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and155_y0;
  wire f_u_cla12_and156_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and156_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and156_y0;
  wire f_u_cla12_and157_f_u_cla12_and156_y0;
  wire f_u_cla12_and157_f_u_cla12_and155_y0;
  wire f_u_cla12_and157_y0;
  wire f_u_cla12_and158_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and158_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and158_y0;
  wire f_u_cla12_and159_f_u_cla12_and158_y0;
  wire f_u_cla12_and159_f_u_cla12_and157_y0;
  wire f_u_cla12_and159_y0;
  wire f_u_cla12_and160_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and160_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and160_y0;
  wire f_u_cla12_and161_f_u_cla12_and160_y0;
  wire f_u_cla12_and161_f_u_cla12_and159_y0;
  wire f_u_cla12_and161_y0;
  wire f_u_cla12_and162_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and162_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and162_y0;
  wire f_u_cla12_and163_f_u_cla12_and162_y0;
  wire f_u_cla12_and163_f_u_cla12_and161_y0;
  wire f_u_cla12_and163_y0;
  wire f_u_cla12_and164_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and164_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and164_y0;
  wire f_u_cla12_and165_f_u_cla12_and164_y0;
  wire f_u_cla12_and165_f_u_cla12_and163_y0;
  wire f_u_cla12_and165_y0;
  wire f_u_cla12_and166_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and166_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and166_y0;
  wire f_u_cla12_and167_f_u_cla12_and166_y0;
  wire f_u_cla12_and167_f_u_cla12_and165_y0;
  wire f_u_cla12_and167_y0;
  wire f_u_cla12_and168_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and168_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and168_y0;
  wire f_u_cla12_and169_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and169_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and169_y0;
  wire f_u_cla12_and170_f_u_cla12_and169_y0;
  wire f_u_cla12_and170_f_u_cla12_and168_y0;
  wire f_u_cla12_and170_y0;
  wire f_u_cla12_and171_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and171_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and171_y0;
  wire f_u_cla12_and172_f_u_cla12_and171_y0;
  wire f_u_cla12_and172_f_u_cla12_and170_y0;
  wire f_u_cla12_and172_y0;
  wire f_u_cla12_and173_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and173_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and173_y0;
  wire f_u_cla12_and174_f_u_cla12_and173_y0;
  wire f_u_cla12_and174_f_u_cla12_and172_y0;
  wire f_u_cla12_and174_y0;
  wire f_u_cla12_and175_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and175_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and175_y0;
  wire f_u_cla12_and176_f_u_cla12_and175_y0;
  wire f_u_cla12_and176_f_u_cla12_and174_y0;
  wire f_u_cla12_and176_y0;
  wire f_u_cla12_and177_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and177_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and177_y0;
  wire f_u_cla12_and178_f_u_cla12_and177_y0;
  wire f_u_cla12_and178_f_u_cla12_and176_y0;
  wire f_u_cla12_and178_y0;
  wire f_u_cla12_and179_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and179_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and179_y0;
  wire f_u_cla12_and180_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and180_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and180_y0;
  wire f_u_cla12_and181_f_u_cla12_and180_y0;
  wire f_u_cla12_and181_f_u_cla12_and179_y0;
  wire f_u_cla12_and181_y0;
  wire f_u_cla12_and182_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and182_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and182_y0;
  wire f_u_cla12_and183_f_u_cla12_and182_y0;
  wire f_u_cla12_and183_f_u_cla12_and181_y0;
  wire f_u_cla12_and183_y0;
  wire f_u_cla12_and184_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and184_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and184_y0;
  wire f_u_cla12_and185_f_u_cla12_and184_y0;
  wire f_u_cla12_and185_f_u_cla12_and183_y0;
  wire f_u_cla12_and185_y0;
  wire f_u_cla12_and186_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and186_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and186_y0;
  wire f_u_cla12_and187_f_u_cla12_and186_y0;
  wire f_u_cla12_and187_f_u_cla12_and185_y0;
  wire f_u_cla12_and187_y0;
  wire f_u_cla12_and188_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and188_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and188_y0;
  wire f_u_cla12_and189_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and189_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and189_y0;
  wire f_u_cla12_and190_f_u_cla12_and189_y0;
  wire f_u_cla12_and190_f_u_cla12_and188_y0;
  wire f_u_cla12_and190_y0;
  wire f_u_cla12_and191_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and191_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and191_y0;
  wire f_u_cla12_and192_f_u_cla12_and191_y0;
  wire f_u_cla12_and192_f_u_cla12_and190_y0;
  wire f_u_cla12_and192_y0;
  wire f_u_cla12_and193_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and193_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and193_y0;
  wire f_u_cla12_and194_f_u_cla12_and193_y0;
  wire f_u_cla12_and194_f_u_cla12_and192_y0;
  wire f_u_cla12_and194_y0;
  wire f_u_cla12_and195_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and195_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and195_y0;
  wire f_u_cla12_and196_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and196_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and196_y0;
  wire f_u_cla12_and197_f_u_cla12_and196_y0;
  wire f_u_cla12_and197_f_u_cla12_and195_y0;
  wire f_u_cla12_and197_y0;
  wire f_u_cla12_and198_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and198_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and198_y0;
  wire f_u_cla12_and199_f_u_cla12_and198_y0;
  wire f_u_cla12_and199_f_u_cla12_and197_y0;
  wire f_u_cla12_and199_y0;
  wire f_u_cla12_and200_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and200_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and200_y0;
  wire f_u_cla12_and201_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and201_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and201_y0;
  wire f_u_cla12_and202_f_u_cla12_and201_y0;
  wire f_u_cla12_and202_f_u_cla12_and200_y0;
  wire f_u_cla12_and202_y0;
  wire f_u_cla12_and203_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and203_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and203_y0;
  wire f_u_cla12_or28_f_u_cla12_and203_y0;
  wire f_u_cla12_or28_f_u_cla12_and154_y0;
  wire f_u_cla12_or28_y0;
  wire f_u_cla12_or29_f_u_cla12_or28_y0;
  wire f_u_cla12_or29_f_u_cla12_and167_y0;
  wire f_u_cla12_or29_y0;
  wire f_u_cla12_or30_f_u_cla12_or29_y0;
  wire f_u_cla12_or30_f_u_cla12_and178_y0;
  wire f_u_cla12_or30_y0;
  wire f_u_cla12_or31_f_u_cla12_or30_y0;
  wire f_u_cla12_or31_f_u_cla12_and187_y0;
  wire f_u_cla12_or31_y0;
  wire f_u_cla12_or32_f_u_cla12_or31_y0;
  wire f_u_cla12_or32_f_u_cla12_and194_y0;
  wire f_u_cla12_or32_y0;
  wire f_u_cla12_or33_f_u_cla12_or32_y0;
  wire f_u_cla12_or33_f_u_cla12_and199_y0;
  wire f_u_cla12_or33_y0;
  wire f_u_cla12_or34_f_u_cla12_or33_y0;
  wire f_u_cla12_or34_f_u_cla12_and202_y0;
  wire f_u_cla12_or34_y0;
  wire f_u_cla12_or35_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_or35_f_u_cla12_or34_y0;
  wire f_u_cla12_or35_y0;
  wire f_u_cla12_pg_logic8_a_8;
  wire f_u_cla12_pg_logic8_b_8;
  wire f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_pg_logic8_y1;
  wire f_u_cla12_pg_logic8_y2;
  wire f_u_cla12_xor8_f_u_cla12_pg_logic8_y2;
  wire f_u_cla12_xor8_f_u_cla12_or35_y0;
  wire f_u_cla12_xor8_y0;
  wire f_u_cla12_and204_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and204_constant_wire_0;
  wire f_u_cla12_and204_y0;
  wire f_u_cla12_and205_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and205_constant_wire_0;
  wire f_u_cla12_and205_y0;
  wire f_u_cla12_and206_f_u_cla12_and205_y0;
  wire f_u_cla12_and206_f_u_cla12_and204_y0;
  wire f_u_cla12_and206_y0;
  wire f_u_cla12_and207_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and207_constant_wire_0;
  wire f_u_cla12_and207_y0;
  wire f_u_cla12_and208_f_u_cla12_and207_y0;
  wire f_u_cla12_and208_f_u_cla12_and206_y0;
  wire f_u_cla12_and208_y0;
  wire f_u_cla12_and209_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and209_constant_wire_0;
  wire f_u_cla12_and209_y0;
  wire f_u_cla12_and210_f_u_cla12_and209_y0;
  wire f_u_cla12_and210_f_u_cla12_and208_y0;
  wire f_u_cla12_and210_y0;
  wire f_u_cla12_and211_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and211_constant_wire_0;
  wire f_u_cla12_and211_y0;
  wire f_u_cla12_and212_f_u_cla12_and211_y0;
  wire f_u_cla12_and212_f_u_cla12_and210_y0;
  wire f_u_cla12_and212_y0;
  wire f_u_cla12_and213_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and213_constant_wire_0;
  wire f_u_cla12_and213_y0;
  wire f_u_cla12_and214_f_u_cla12_and213_y0;
  wire f_u_cla12_and214_f_u_cla12_and212_y0;
  wire f_u_cla12_and214_y0;
  wire f_u_cla12_and215_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and215_constant_wire_0;
  wire f_u_cla12_and215_y0;
  wire f_u_cla12_and216_f_u_cla12_and215_y0;
  wire f_u_cla12_and216_f_u_cla12_and214_y0;
  wire f_u_cla12_and216_y0;
  wire f_u_cla12_and217_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and217_constant_wire_0;
  wire f_u_cla12_and217_y0;
  wire f_u_cla12_and218_f_u_cla12_and217_y0;
  wire f_u_cla12_and218_f_u_cla12_and216_y0;
  wire f_u_cla12_and218_y0;
  wire f_u_cla12_and219_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and219_constant_wire_0;
  wire f_u_cla12_and219_y0;
  wire f_u_cla12_and220_f_u_cla12_and219_y0;
  wire f_u_cla12_and220_f_u_cla12_and218_y0;
  wire f_u_cla12_and220_y0;
  wire f_u_cla12_and221_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and221_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and221_y0;
  wire f_u_cla12_and222_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and222_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and222_y0;
  wire f_u_cla12_and223_f_u_cla12_and222_y0;
  wire f_u_cla12_and223_f_u_cla12_and221_y0;
  wire f_u_cla12_and223_y0;
  wire f_u_cla12_and224_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and224_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and224_y0;
  wire f_u_cla12_and225_f_u_cla12_and224_y0;
  wire f_u_cla12_and225_f_u_cla12_and223_y0;
  wire f_u_cla12_and225_y0;
  wire f_u_cla12_and226_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and226_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and226_y0;
  wire f_u_cla12_and227_f_u_cla12_and226_y0;
  wire f_u_cla12_and227_f_u_cla12_and225_y0;
  wire f_u_cla12_and227_y0;
  wire f_u_cla12_and228_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and228_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and228_y0;
  wire f_u_cla12_and229_f_u_cla12_and228_y0;
  wire f_u_cla12_and229_f_u_cla12_and227_y0;
  wire f_u_cla12_and229_y0;
  wire f_u_cla12_and230_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and230_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and230_y0;
  wire f_u_cla12_and231_f_u_cla12_and230_y0;
  wire f_u_cla12_and231_f_u_cla12_and229_y0;
  wire f_u_cla12_and231_y0;
  wire f_u_cla12_and232_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and232_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and232_y0;
  wire f_u_cla12_and233_f_u_cla12_and232_y0;
  wire f_u_cla12_and233_f_u_cla12_and231_y0;
  wire f_u_cla12_and233_y0;
  wire f_u_cla12_and234_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and234_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and234_y0;
  wire f_u_cla12_and235_f_u_cla12_and234_y0;
  wire f_u_cla12_and235_f_u_cla12_and233_y0;
  wire f_u_cla12_and235_y0;
  wire f_u_cla12_and236_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and236_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and236_y0;
  wire f_u_cla12_and237_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and237_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and237_y0;
  wire f_u_cla12_and238_f_u_cla12_and237_y0;
  wire f_u_cla12_and238_f_u_cla12_and236_y0;
  wire f_u_cla12_and238_y0;
  wire f_u_cla12_and239_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and239_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and239_y0;
  wire f_u_cla12_and240_f_u_cla12_and239_y0;
  wire f_u_cla12_and240_f_u_cla12_and238_y0;
  wire f_u_cla12_and240_y0;
  wire f_u_cla12_and241_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and241_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and241_y0;
  wire f_u_cla12_and242_f_u_cla12_and241_y0;
  wire f_u_cla12_and242_f_u_cla12_and240_y0;
  wire f_u_cla12_and242_y0;
  wire f_u_cla12_and243_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and243_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and243_y0;
  wire f_u_cla12_and244_f_u_cla12_and243_y0;
  wire f_u_cla12_and244_f_u_cla12_and242_y0;
  wire f_u_cla12_and244_y0;
  wire f_u_cla12_and245_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and245_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and245_y0;
  wire f_u_cla12_and246_f_u_cla12_and245_y0;
  wire f_u_cla12_and246_f_u_cla12_and244_y0;
  wire f_u_cla12_and246_y0;
  wire f_u_cla12_and247_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and247_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and247_y0;
  wire f_u_cla12_and248_f_u_cla12_and247_y0;
  wire f_u_cla12_and248_f_u_cla12_and246_y0;
  wire f_u_cla12_and248_y0;
  wire f_u_cla12_and249_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and249_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and249_y0;
  wire f_u_cla12_and250_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and250_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and250_y0;
  wire f_u_cla12_and251_f_u_cla12_and250_y0;
  wire f_u_cla12_and251_f_u_cla12_and249_y0;
  wire f_u_cla12_and251_y0;
  wire f_u_cla12_and252_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and252_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and252_y0;
  wire f_u_cla12_and253_f_u_cla12_and252_y0;
  wire f_u_cla12_and253_f_u_cla12_and251_y0;
  wire f_u_cla12_and253_y0;
  wire f_u_cla12_and254_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and254_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and254_y0;
  wire f_u_cla12_and255_f_u_cla12_and254_y0;
  wire f_u_cla12_and255_f_u_cla12_and253_y0;
  wire f_u_cla12_and255_y0;
  wire f_u_cla12_and256_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and256_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and256_y0;
  wire f_u_cla12_and257_f_u_cla12_and256_y0;
  wire f_u_cla12_and257_f_u_cla12_and255_y0;
  wire f_u_cla12_and257_y0;
  wire f_u_cla12_and258_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and258_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and258_y0;
  wire f_u_cla12_and259_f_u_cla12_and258_y0;
  wire f_u_cla12_and259_f_u_cla12_and257_y0;
  wire f_u_cla12_and259_y0;
  wire f_u_cla12_and260_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and260_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and260_y0;
  wire f_u_cla12_and261_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and261_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and261_y0;
  wire f_u_cla12_and262_f_u_cla12_and261_y0;
  wire f_u_cla12_and262_f_u_cla12_and260_y0;
  wire f_u_cla12_and262_y0;
  wire f_u_cla12_and263_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and263_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and263_y0;
  wire f_u_cla12_and264_f_u_cla12_and263_y0;
  wire f_u_cla12_and264_f_u_cla12_and262_y0;
  wire f_u_cla12_and264_y0;
  wire f_u_cla12_and265_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and265_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and265_y0;
  wire f_u_cla12_and266_f_u_cla12_and265_y0;
  wire f_u_cla12_and266_f_u_cla12_and264_y0;
  wire f_u_cla12_and266_y0;
  wire f_u_cla12_and267_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and267_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and267_y0;
  wire f_u_cla12_and268_f_u_cla12_and267_y0;
  wire f_u_cla12_and268_f_u_cla12_and266_y0;
  wire f_u_cla12_and268_y0;
  wire f_u_cla12_and269_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and269_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and269_y0;
  wire f_u_cla12_and270_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and270_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and270_y0;
  wire f_u_cla12_and271_f_u_cla12_and270_y0;
  wire f_u_cla12_and271_f_u_cla12_and269_y0;
  wire f_u_cla12_and271_y0;
  wire f_u_cla12_and272_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and272_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and272_y0;
  wire f_u_cla12_and273_f_u_cla12_and272_y0;
  wire f_u_cla12_and273_f_u_cla12_and271_y0;
  wire f_u_cla12_and273_y0;
  wire f_u_cla12_and274_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and274_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and274_y0;
  wire f_u_cla12_and275_f_u_cla12_and274_y0;
  wire f_u_cla12_and275_f_u_cla12_and273_y0;
  wire f_u_cla12_and275_y0;
  wire f_u_cla12_and276_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and276_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and276_y0;
  wire f_u_cla12_and277_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and277_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and277_y0;
  wire f_u_cla12_and278_f_u_cla12_and277_y0;
  wire f_u_cla12_and278_f_u_cla12_and276_y0;
  wire f_u_cla12_and278_y0;
  wire f_u_cla12_and279_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and279_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and279_y0;
  wire f_u_cla12_and280_f_u_cla12_and279_y0;
  wire f_u_cla12_and280_f_u_cla12_and278_y0;
  wire f_u_cla12_and280_y0;
  wire f_u_cla12_and281_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and281_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and281_y0;
  wire f_u_cla12_and282_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and282_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and282_y0;
  wire f_u_cla12_and283_f_u_cla12_and282_y0;
  wire f_u_cla12_and283_f_u_cla12_and281_y0;
  wire f_u_cla12_and283_y0;
  wire f_u_cla12_and284_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and284_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and284_y0;
  wire f_u_cla12_or36_f_u_cla12_and284_y0;
  wire f_u_cla12_or36_f_u_cla12_and220_y0;
  wire f_u_cla12_or36_y0;
  wire f_u_cla12_or37_f_u_cla12_or36_y0;
  wire f_u_cla12_or37_f_u_cla12_and235_y0;
  wire f_u_cla12_or37_y0;
  wire f_u_cla12_or38_f_u_cla12_or37_y0;
  wire f_u_cla12_or38_f_u_cla12_and248_y0;
  wire f_u_cla12_or38_y0;
  wire f_u_cla12_or39_f_u_cla12_or38_y0;
  wire f_u_cla12_or39_f_u_cla12_and259_y0;
  wire f_u_cla12_or39_y0;
  wire f_u_cla12_or40_f_u_cla12_or39_y0;
  wire f_u_cla12_or40_f_u_cla12_and268_y0;
  wire f_u_cla12_or40_y0;
  wire f_u_cla12_or41_f_u_cla12_or40_y0;
  wire f_u_cla12_or41_f_u_cla12_and275_y0;
  wire f_u_cla12_or41_y0;
  wire f_u_cla12_or42_f_u_cla12_or41_y0;
  wire f_u_cla12_or42_f_u_cla12_and280_y0;
  wire f_u_cla12_or42_y0;
  wire f_u_cla12_or43_f_u_cla12_or42_y0;
  wire f_u_cla12_or43_f_u_cla12_and283_y0;
  wire f_u_cla12_or43_y0;
  wire f_u_cla12_or44_f_u_cla12_pg_logic8_y1;
  wire f_u_cla12_or44_f_u_cla12_or43_y0;
  wire f_u_cla12_or44_y0;
  wire f_u_cla12_pg_logic9_a_9;
  wire f_u_cla12_pg_logic9_b_9;
  wire f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_pg_logic9_y1;
  wire f_u_cla12_pg_logic9_y2;
  wire f_u_cla12_xor9_f_u_cla12_pg_logic9_y2;
  wire f_u_cla12_xor9_f_u_cla12_or44_y0;
  wire f_u_cla12_xor9_y0;
  wire f_u_cla12_and285_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and285_constant_wire_0;
  wire f_u_cla12_and285_y0;
  wire f_u_cla12_and286_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and286_constant_wire_0;
  wire f_u_cla12_and286_y0;
  wire f_u_cla12_and287_f_u_cla12_and286_y0;
  wire f_u_cla12_and287_f_u_cla12_and285_y0;
  wire f_u_cla12_and287_y0;
  wire f_u_cla12_and288_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and288_constant_wire_0;
  wire f_u_cla12_and288_y0;
  wire f_u_cla12_and289_f_u_cla12_and288_y0;
  wire f_u_cla12_and289_f_u_cla12_and287_y0;
  wire f_u_cla12_and289_y0;
  wire f_u_cla12_and290_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and290_constant_wire_0;
  wire f_u_cla12_and290_y0;
  wire f_u_cla12_and291_f_u_cla12_and290_y0;
  wire f_u_cla12_and291_f_u_cla12_and289_y0;
  wire f_u_cla12_and291_y0;
  wire f_u_cla12_and292_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and292_constant_wire_0;
  wire f_u_cla12_and292_y0;
  wire f_u_cla12_and293_f_u_cla12_and292_y0;
  wire f_u_cla12_and293_f_u_cla12_and291_y0;
  wire f_u_cla12_and293_y0;
  wire f_u_cla12_and294_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and294_constant_wire_0;
  wire f_u_cla12_and294_y0;
  wire f_u_cla12_and295_f_u_cla12_and294_y0;
  wire f_u_cla12_and295_f_u_cla12_and293_y0;
  wire f_u_cla12_and295_y0;
  wire f_u_cla12_and296_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and296_constant_wire_0;
  wire f_u_cla12_and296_y0;
  wire f_u_cla12_and297_f_u_cla12_and296_y0;
  wire f_u_cla12_and297_f_u_cla12_and295_y0;
  wire f_u_cla12_and297_y0;
  wire f_u_cla12_and298_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and298_constant_wire_0;
  wire f_u_cla12_and298_y0;
  wire f_u_cla12_and299_f_u_cla12_and298_y0;
  wire f_u_cla12_and299_f_u_cla12_and297_y0;
  wire f_u_cla12_and299_y0;
  wire f_u_cla12_and300_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and300_constant_wire_0;
  wire f_u_cla12_and300_y0;
  wire f_u_cla12_and301_f_u_cla12_and300_y0;
  wire f_u_cla12_and301_f_u_cla12_and299_y0;
  wire f_u_cla12_and301_y0;
  wire f_u_cla12_and302_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and302_constant_wire_0;
  wire f_u_cla12_and302_y0;
  wire f_u_cla12_and303_f_u_cla12_and302_y0;
  wire f_u_cla12_and303_f_u_cla12_and301_y0;
  wire f_u_cla12_and303_y0;
  wire f_u_cla12_and304_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and304_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and304_y0;
  wire f_u_cla12_and305_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and305_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and305_y0;
  wire f_u_cla12_and306_f_u_cla12_and305_y0;
  wire f_u_cla12_and306_f_u_cla12_and304_y0;
  wire f_u_cla12_and306_y0;
  wire f_u_cla12_and307_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and307_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and307_y0;
  wire f_u_cla12_and308_f_u_cla12_and307_y0;
  wire f_u_cla12_and308_f_u_cla12_and306_y0;
  wire f_u_cla12_and308_y0;
  wire f_u_cla12_and309_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and309_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and309_y0;
  wire f_u_cla12_and310_f_u_cla12_and309_y0;
  wire f_u_cla12_and310_f_u_cla12_and308_y0;
  wire f_u_cla12_and310_y0;
  wire f_u_cla12_and311_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and311_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and311_y0;
  wire f_u_cla12_and312_f_u_cla12_and311_y0;
  wire f_u_cla12_and312_f_u_cla12_and310_y0;
  wire f_u_cla12_and312_y0;
  wire f_u_cla12_and313_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and313_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and313_y0;
  wire f_u_cla12_and314_f_u_cla12_and313_y0;
  wire f_u_cla12_and314_f_u_cla12_and312_y0;
  wire f_u_cla12_and314_y0;
  wire f_u_cla12_and315_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and315_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and315_y0;
  wire f_u_cla12_and316_f_u_cla12_and315_y0;
  wire f_u_cla12_and316_f_u_cla12_and314_y0;
  wire f_u_cla12_and316_y0;
  wire f_u_cla12_and317_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and317_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and317_y0;
  wire f_u_cla12_and318_f_u_cla12_and317_y0;
  wire f_u_cla12_and318_f_u_cla12_and316_y0;
  wire f_u_cla12_and318_y0;
  wire f_u_cla12_and319_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and319_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and319_y0;
  wire f_u_cla12_and320_f_u_cla12_and319_y0;
  wire f_u_cla12_and320_f_u_cla12_and318_y0;
  wire f_u_cla12_and320_y0;
  wire f_u_cla12_and321_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and321_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and321_y0;
  wire f_u_cla12_and322_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and322_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and322_y0;
  wire f_u_cla12_and323_f_u_cla12_and322_y0;
  wire f_u_cla12_and323_f_u_cla12_and321_y0;
  wire f_u_cla12_and323_y0;
  wire f_u_cla12_and324_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and324_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and324_y0;
  wire f_u_cla12_and325_f_u_cla12_and324_y0;
  wire f_u_cla12_and325_f_u_cla12_and323_y0;
  wire f_u_cla12_and325_y0;
  wire f_u_cla12_and326_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and326_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and326_y0;
  wire f_u_cla12_and327_f_u_cla12_and326_y0;
  wire f_u_cla12_and327_f_u_cla12_and325_y0;
  wire f_u_cla12_and327_y0;
  wire f_u_cla12_and328_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and328_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and328_y0;
  wire f_u_cla12_and329_f_u_cla12_and328_y0;
  wire f_u_cla12_and329_f_u_cla12_and327_y0;
  wire f_u_cla12_and329_y0;
  wire f_u_cla12_and330_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and330_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and330_y0;
  wire f_u_cla12_and331_f_u_cla12_and330_y0;
  wire f_u_cla12_and331_f_u_cla12_and329_y0;
  wire f_u_cla12_and331_y0;
  wire f_u_cla12_and332_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and332_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and332_y0;
  wire f_u_cla12_and333_f_u_cla12_and332_y0;
  wire f_u_cla12_and333_f_u_cla12_and331_y0;
  wire f_u_cla12_and333_y0;
  wire f_u_cla12_and334_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and334_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and334_y0;
  wire f_u_cla12_and335_f_u_cla12_and334_y0;
  wire f_u_cla12_and335_f_u_cla12_and333_y0;
  wire f_u_cla12_and335_y0;
  wire f_u_cla12_and336_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and336_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and336_y0;
  wire f_u_cla12_and337_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and337_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and337_y0;
  wire f_u_cla12_and338_f_u_cla12_and337_y0;
  wire f_u_cla12_and338_f_u_cla12_and336_y0;
  wire f_u_cla12_and338_y0;
  wire f_u_cla12_and339_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and339_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and339_y0;
  wire f_u_cla12_and340_f_u_cla12_and339_y0;
  wire f_u_cla12_and340_f_u_cla12_and338_y0;
  wire f_u_cla12_and340_y0;
  wire f_u_cla12_and341_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and341_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and341_y0;
  wire f_u_cla12_and342_f_u_cla12_and341_y0;
  wire f_u_cla12_and342_f_u_cla12_and340_y0;
  wire f_u_cla12_and342_y0;
  wire f_u_cla12_and343_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and343_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and343_y0;
  wire f_u_cla12_and344_f_u_cla12_and343_y0;
  wire f_u_cla12_and344_f_u_cla12_and342_y0;
  wire f_u_cla12_and344_y0;
  wire f_u_cla12_and345_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and345_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and345_y0;
  wire f_u_cla12_and346_f_u_cla12_and345_y0;
  wire f_u_cla12_and346_f_u_cla12_and344_y0;
  wire f_u_cla12_and346_y0;
  wire f_u_cla12_and347_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and347_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and347_y0;
  wire f_u_cla12_and348_f_u_cla12_and347_y0;
  wire f_u_cla12_and348_f_u_cla12_and346_y0;
  wire f_u_cla12_and348_y0;
  wire f_u_cla12_and349_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and349_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and349_y0;
  wire f_u_cla12_and350_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and350_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and350_y0;
  wire f_u_cla12_and351_f_u_cla12_and350_y0;
  wire f_u_cla12_and351_f_u_cla12_and349_y0;
  wire f_u_cla12_and351_y0;
  wire f_u_cla12_and352_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and352_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and352_y0;
  wire f_u_cla12_and353_f_u_cla12_and352_y0;
  wire f_u_cla12_and353_f_u_cla12_and351_y0;
  wire f_u_cla12_and353_y0;
  wire f_u_cla12_and354_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and354_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and354_y0;
  wire f_u_cla12_and355_f_u_cla12_and354_y0;
  wire f_u_cla12_and355_f_u_cla12_and353_y0;
  wire f_u_cla12_and355_y0;
  wire f_u_cla12_and356_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and356_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and356_y0;
  wire f_u_cla12_and357_f_u_cla12_and356_y0;
  wire f_u_cla12_and357_f_u_cla12_and355_y0;
  wire f_u_cla12_and357_y0;
  wire f_u_cla12_and358_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and358_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and358_y0;
  wire f_u_cla12_and359_f_u_cla12_and358_y0;
  wire f_u_cla12_and359_f_u_cla12_and357_y0;
  wire f_u_cla12_and359_y0;
  wire f_u_cla12_and360_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and360_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and360_y0;
  wire f_u_cla12_and361_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and361_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and361_y0;
  wire f_u_cla12_and362_f_u_cla12_and361_y0;
  wire f_u_cla12_and362_f_u_cla12_and360_y0;
  wire f_u_cla12_and362_y0;
  wire f_u_cla12_and363_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and363_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and363_y0;
  wire f_u_cla12_and364_f_u_cla12_and363_y0;
  wire f_u_cla12_and364_f_u_cla12_and362_y0;
  wire f_u_cla12_and364_y0;
  wire f_u_cla12_and365_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and365_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and365_y0;
  wire f_u_cla12_and366_f_u_cla12_and365_y0;
  wire f_u_cla12_and366_f_u_cla12_and364_y0;
  wire f_u_cla12_and366_y0;
  wire f_u_cla12_and367_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and367_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and367_y0;
  wire f_u_cla12_and368_f_u_cla12_and367_y0;
  wire f_u_cla12_and368_f_u_cla12_and366_y0;
  wire f_u_cla12_and368_y0;
  wire f_u_cla12_and369_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and369_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and369_y0;
  wire f_u_cla12_and370_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and370_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and370_y0;
  wire f_u_cla12_and371_f_u_cla12_and370_y0;
  wire f_u_cla12_and371_f_u_cla12_and369_y0;
  wire f_u_cla12_and371_y0;
  wire f_u_cla12_and372_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and372_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and372_y0;
  wire f_u_cla12_and373_f_u_cla12_and372_y0;
  wire f_u_cla12_and373_f_u_cla12_and371_y0;
  wire f_u_cla12_and373_y0;
  wire f_u_cla12_and374_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and374_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and374_y0;
  wire f_u_cla12_and375_f_u_cla12_and374_y0;
  wire f_u_cla12_and375_f_u_cla12_and373_y0;
  wire f_u_cla12_and375_y0;
  wire f_u_cla12_and376_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and376_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and376_y0;
  wire f_u_cla12_and377_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and377_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and377_y0;
  wire f_u_cla12_and378_f_u_cla12_and377_y0;
  wire f_u_cla12_and378_f_u_cla12_and376_y0;
  wire f_u_cla12_and378_y0;
  wire f_u_cla12_and379_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and379_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and379_y0;
  wire f_u_cla12_and380_f_u_cla12_and379_y0;
  wire f_u_cla12_and380_f_u_cla12_and378_y0;
  wire f_u_cla12_and380_y0;
  wire f_u_cla12_and381_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and381_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and381_y0;
  wire f_u_cla12_and382_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and382_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and382_y0;
  wire f_u_cla12_and383_f_u_cla12_and382_y0;
  wire f_u_cla12_and383_f_u_cla12_and381_y0;
  wire f_u_cla12_and383_y0;
  wire f_u_cla12_and384_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and384_f_u_cla12_pg_logic8_y1;
  wire f_u_cla12_and384_y0;
  wire f_u_cla12_or45_f_u_cla12_and384_y0;
  wire f_u_cla12_or45_f_u_cla12_and303_y0;
  wire f_u_cla12_or45_y0;
  wire f_u_cla12_or46_f_u_cla12_or45_y0;
  wire f_u_cla12_or46_f_u_cla12_and320_y0;
  wire f_u_cla12_or46_y0;
  wire f_u_cla12_or47_f_u_cla12_or46_y0;
  wire f_u_cla12_or47_f_u_cla12_and335_y0;
  wire f_u_cla12_or47_y0;
  wire f_u_cla12_or48_f_u_cla12_or47_y0;
  wire f_u_cla12_or48_f_u_cla12_and348_y0;
  wire f_u_cla12_or48_y0;
  wire f_u_cla12_or49_f_u_cla12_or48_y0;
  wire f_u_cla12_or49_f_u_cla12_and359_y0;
  wire f_u_cla12_or49_y0;
  wire f_u_cla12_or50_f_u_cla12_or49_y0;
  wire f_u_cla12_or50_f_u_cla12_and368_y0;
  wire f_u_cla12_or50_y0;
  wire f_u_cla12_or51_f_u_cla12_or50_y0;
  wire f_u_cla12_or51_f_u_cla12_and375_y0;
  wire f_u_cla12_or51_y0;
  wire f_u_cla12_or52_f_u_cla12_or51_y0;
  wire f_u_cla12_or52_f_u_cla12_and380_y0;
  wire f_u_cla12_or52_y0;
  wire f_u_cla12_or53_f_u_cla12_or52_y0;
  wire f_u_cla12_or53_f_u_cla12_and383_y0;
  wire f_u_cla12_or53_y0;
  wire f_u_cla12_or54_f_u_cla12_pg_logic9_y1;
  wire f_u_cla12_or54_f_u_cla12_or53_y0;
  wire f_u_cla12_or54_y0;
  wire f_u_cla12_pg_logic10_a_10;
  wire f_u_cla12_pg_logic10_b_10;
  wire f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_pg_logic10_y1;
  wire f_u_cla12_pg_logic10_y2;
  wire f_u_cla12_xor10_f_u_cla12_pg_logic10_y2;
  wire f_u_cla12_xor10_f_u_cla12_or54_y0;
  wire f_u_cla12_xor10_y0;
  wire f_u_cla12_and385_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and385_constant_wire_0;
  wire f_u_cla12_and385_y0;
  wire f_u_cla12_and386_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and386_constant_wire_0;
  wire f_u_cla12_and386_y0;
  wire f_u_cla12_and387_f_u_cla12_and386_y0;
  wire f_u_cla12_and387_f_u_cla12_and385_y0;
  wire f_u_cla12_and387_y0;
  wire f_u_cla12_and388_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and388_constant_wire_0;
  wire f_u_cla12_and388_y0;
  wire f_u_cla12_and389_f_u_cla12_and388_y0;
  wire f_u_cla12_and389_f_u_cla12_and387_y0;
  wire f_u_cla12_and389_y0;
  wire f_u_cla12_and390_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and390_constant_wire_0;
  wire f_u_cla12_and390_y0;
  wire f_u_cla12_and391_f_u_cla12_and390_y0;
  wire f_u_cla12_and391_f_u_cla12_and389_y0;
  wire f_u_cla12_and391_y0;
  wire f_u_cla12_and392_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and392_constant_wire_0;
  wire f_u_cla12_and392_y0;
  wire f_u_cla12_and393_f_u_cla12_and392_y0;
  wire f_u_cla12_and393_f_u_cla12_and391_y0;
  wire f_u_cla12_and393_y0;
  wire f_u_cla12_and394_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and394_constant_wire_0;
  wire f_u_cla12_and394_y0;
  wire f_u_cla12_and395_f_u_cla12_and394_y0;
  wire f_u_cla12_and395_f_u_cla12_and393_y0;
  wire f_u_cla12_and395_y0;
  wire f_u_cla12_and396_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and396_constant_wire_0;
  wire f_u_cla12_and396_y0;
  wire f_u_cla12_and397_f_u_cla12_and396_y0;
  wire f_u_cla12_and397_f_u_cla12_and395_y0;
  wire f_u_cla12_and397_y0;
  wire f_u_cla12_and398_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and398_constant_wire_0;
  wire f_u_cla12_and398_y0;
  wire f_u_cla12_and399_f_u_cla12_and398_y0;
  wire f_u_cla12_and399_f_u_cla12_and397_y0;
  wire f_u_cla12_and399_y0;
  wire f_u_cla12_and400_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and400_constant_wire_0;
  wire f_u_cla12_and400_y0;
  wire f_u_cla12_and401_f_u_cla12_and400_y0;
  wire f_u_cla12_and401_f_u_cla12_and399_y0;
  wire f_u_cla12_and401_y0;
  wire f_u_cla12_and402_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and402_constant_wire_0;
  wire f_u_cla12_and402_y0;
  wire f_u_cla12_and403_f_u_cla12_and402_y0;
  wire f_u_cla12_and403_f_u_cla12_and401_y0;
  wire f_u_cla12_and403_y0;
  wire f_u_cla12_and404_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and404_constant_wire_0;
  wire f_u_cla12_and404_y0;
  wire f_u_cla12_and405_f_u_cla12_and404_y0;
  wire f_u_cla12_and405_f_u_cla12_and403_y0;
  wire f_u_cla12_and405_y0;
  wire f_u_cla12_and406_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and406_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and406_y0;
  wire f_u_cla12_and407_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and407_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and407_y0;
  wire f_u_cla12_and408_f_u_cla12_and407_y0;
  wire f_u_cla12_and408_f_u_cla12_and406_y0;
  wire f_u_cla12_and408_y0;
  wire f_u_cla12_and409_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and409_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and409_y0;
  wire f_u_cla12_and410_f_u_cla12_and409_y0;
  wire f_u_cla12_and410_f_u_cla12_and408_y0;
  wire f_u_cla12_and410_y0;
  wire f_u_cla12_and411_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and411_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and411_y0;
  wire f_u_cla12_and412_f_u_cla12_and411_y0;
  wire f_u_cla12_and412_f_u_cla12_and410_y0;
  wire f_u_cla12_and412_y0;
  wire f_u_cla12_and413_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and413_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and413_y0;
  wire f_u_cla12_and414_f_u_cla12_and413_y0;
  wire f_u_cla12_and414_f_u_cla12_and412_y0;
  wire f_u_cla12_and414_y0;
  wire f_u_cla12_and415_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and415_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and415_y0;
  wire f_u_cla12_and416_f_u_cla12_and415_y0;
  wire f_u_cla12_and416_f_u_cla12_and414_y0;
  wire f_u_cla12_and416_y0;
  wire f_u_cla12_and417_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and417_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and417_y0;
  wire f_u_cla12_and418_f_u_cla12_and417_y0;
  wire f_u_cla12_and418_f_u_cla12_and416_y0;
  wire f_u_cla12_and418_y0;
  wire f_u_cla12_and419_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and419_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and419_y0;
  wire f_u_cla12_and420_f_u_cla12_and419_y0;
  wire f_u_cla12_and420_f_u_cla12_and418_y0;
  wire f_u_cla12_and420_y0;
  wire f_u_cla12_and421_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and421_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and421_y0;
  wire f_u_cla12_and422_f_u_cla12_and421_y0;
  wire f_u_cla12_and422_f_u_cla12_and420_y0;
  wire f_u_cla12_and422_y0;
  wire f_u_cla12_and423_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and423_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and423_y0;
  wire f_u_cla12_and424_f_u_cla12_and423_y0;
  wire f_u_cla12_and424_f_u_cla12_and422_y0;
  wire f_u_cla12_and424_y0;
  wire f_u_cla12_and425_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and425_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and425_y0;
  wire f_u_cla12_and426_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and426_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and426_y0;
  wire f_u_cla12_and427_f_u_cla12_and426_y0;
  wire f_u_cla12_and427_f_u_cla12_and425_y0;
  wire f_u_cla12_and427_y0;
  wire f_u_cla12_and428_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and428_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and428_y0;
  wire f_u_cla12_and429_f_u_cla12_and428_y0;
  wire f_u_cla12_and429_f_u_cla12_and427_y0;
  wire f_u_cla12_and429_y0;
  wire f_u_cla12_and430_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and430_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and430_y0;
  wire f_u_cla12_and431_f_u_cla12_and430_y0;
  wire f_u_cla12_and431_f_u_cla12_and429_y0;
  wire f_u_cla12_and431_y0;
  wire f_u_cla12_and432_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and432_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and432_y0;
  wire f_u_cla12_and433_f_u_cla12_and432_y0;
  wire f_u_cla12_and433_f_u_cla12_and431_y0;
  wire f_u_cla12_and433_y0;
  wire f_u_cla12_and434_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and434_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and434_y0;
  wire f_u_cla12_and435_f_u_cla12_and434_y0;
  wire f_u_cla12_and435_f_u_cla12_and433_y0;
  wire f_u_cla12_and435_y0;
  wire f_u_cla12_and436_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and436_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and436_y0;
  wire f_u_cla12_and437_f_u_cla12_and436_y0;
  wire f_u_cla12_and437_f_u_cla12_and435_y0;
  wire f_u_cla12_and437_y0;
  wire f_u_cla12_and438_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and438_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and438_y0;
  wire f_u_cla12_and439_f_u_cla12_and438_y0;
  wire f_u_cla12_and439_f_u_cla12_and437_y0;
  wire f_u_cla12_and439_y0;
  wire f_u_cla12_and440_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and440_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and440_y0;
  wire f_u_cla12_and441_f_u_cla12_and440_y0;
  wire f_u_cla12_and441_f_u_cla12_and439_y0;
  wire f_u_cla12_and441_y0;
  wire f_u_cla12_and442_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and442_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and442_y0;
  wire f_u_cla12_and443_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and443_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and443_y0;
  wire f_u_cla12_and444_f_u_cla12_and443_y0;
  wire f_u_cla12_and444_f_u_cla12_and442_y0;
  wire f_u_cla12_and444_y0;
  wire f_u_cla12_and445_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and445_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and445_y0;
  wire f_u_cla12_and446_f_u_cla12_and445_y0;
  wire f_u_cla12_and446_f_u_cla12_and444_y0;
  wire f_u_cla12_and446_y0;
  wire f_u_cla12_and447_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and447_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and447_y0;
  wire f_u_cla12_and448_f_u_cla12_and447_y0;
  wire f_u_cla12_and448_f_u_cla12_and446_y0;
  wire f_u_cla12_and448_y0;
  wire f_u_cla12_and449_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and449_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and449_y0;
  wire f_u_cla12_and450_f_u_cla12_and449_y0;
  wire f_u_cla12_and450_f_u_cla12_and448_y0;
  wire f_u_cla12_and450_y0;
  wire f_u_cla12_and451_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and451_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and451_y0;
  wire f_u_cla12_and452_f_u_cla12_and451_y0;
  wire f_u_cla12_and452_f_u_cla12_and450_y0;
  wire f_u_cla12_and452_y0;
  wire f_u_cla12_and453_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and453_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and453_y0;
  wire f_u_cla12_and454_f_u_cla12_and453_y0;
  wire f_u_cla12_and454_f_u_cla12_and452_y0;
  wire f_u_cla12_and454_y0;
  wire f_u_cla12_and455_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and455_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and455_y0;
  wire f_u_cla12_and456_f_u_cla12_and455_y0;
  wire f_u_cla12_and456_f_u_cla12_and454_y0;
  wire f_u_cla12_and456_y0;
  wire f_u_cla12_and457_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and457_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and457_y0;
  wire f_u_cla12_and458_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and458_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and458_y0;
  wire f_u_cla12_and459_f_u_cla12_and458_y0;
  wire f_u_cla12_and459_f_u_cla12_and457_y0;
  wire f_u_cla12_and459_y0;
  wire f_u_cla12_and460_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and460_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and460_y0;
  wire f_u_cla12_and461_f_u_cla12_and460_y0;
  wire f_u_cla12_and461_f_u_cla12_and459_y0;
  wire f_u_cla12_and461_y0;
  wire f_u_cla12_and462_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and462_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and462_y0;
  wire f_u_cla12_and463_f_u_cla12_and462_y0;
  wire f_u_cla12_and463_f_u_cla12_and461_y0;
  wire f_u_cla12_and463_y0;
  wire f_u_cla12_and464_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and464_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and464_y0;
  wire f_u_cla12_and465_f_u_cla12_and464_y0;
  wire f_u_cla12_and465_f_u_cla12_and463_y0;
  wire f_u_cla12_and465_y0;
  wire f_u_cla12_and466_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and466_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and466_y0;
  wire f_u_cla12_and467_f_u_cla12_and466_y0;
  wire f_u_cla12_and467_f_u_cla12_and465_y0;
  wire f_u_cla12_and467_y0;
  wire f_u_cla12_and468_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and468_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and468_y0;
  wire f_u_cla12_and469_f_u_cla12_and468_y0;
  wire f_u_cla12_and469_f_u_cla12_and467_y0;
  wire f_u_cla12_and469_y0;
  wire f_u_cla12_and470_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and470_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and470_y0;
  wire f_u_cla12_and471_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and471_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and471_y0;
  wire f_u_cla12_and472_f_u_cla12_and471_y0;
  wire f_u_cla12_and472_f_u_cla12_and470_y0;
  wire f_u_cla12_and472_y0;
  wire f_u_cla12_and473_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and473_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and473_y0;
  wire f_u_cla12_and474_f_u_cla12_and473_y0;
  wire f_u_cla12_and474_f_u_cla12_and472_y0;
  wire f_u_cla12_and474_y0;
  wire f_u_cla12_and475_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and475_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and475_y0;
  wire f_u_cla12_and476_f_u_cla12_and475_y0;
  wire f_u_cla12_and476_f_u_cla12_and474_y0;
  wire f_u_cla12_and476_y0;
  wire f_u_cla12_and477_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and477_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and477_y0;
  wire f_u_cla12_and478_f_u_cla12_and477_y0;
  wire f_u_cla12_and478_f_u_cla12_and476_y0;
  wire f_u_cla12_and478_y0;
  wire f_u_cla12_and479_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and479_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and479_y0;
  wire f_u_cla12_and480_f_u_cla12_and479_y0;
  wire f_u_cla12_and480_f_u_cla12_and478_y0;
  wire f_u_cla12_and480_y0;
  wire f_u_cla12_and481_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and481_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and481_y0;
  wire f_u_cla12_and482_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and482_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and482_y0;
  wire f_u_cla12_and483_f_u_cla12_and482_y0;
  wire f_u_cla12_and483_f_u_cla12_and481_y0;
  wire f_u_cla12_and483_y0;
  wire f_u_cla12_and484_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and484_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and484_y0;
  wire f_u_cla12_and485_f_u_cla12_and484_y0;
  wire f_u_cla12_and485_f_u_cla12_and483_y0;
  wire f_u_cla12_and485_y0;
  wire f_u_cla12_and486_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and486_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and486_y0;
  wire f_u_cla12_and487_f_u_cla12_and486_y0;
  wire f_u_cla12_and487_f_u_cla12_and485_y0;
  wire f_u_cla12_and487_y0;
  wire f_u_cla12_and488_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and488_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and488_y0;
  wire f_u_cla12_and489_f_u_cla12_and488_y0;
  wire f_u_cla12_and489_f_u_cla12_and487_y0;
  wire f_u_cla12_and489_y0;
  wire f_u_cla12_and490_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and490_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and490_y0;
  wire f_u_cla12_and491_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and491_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and491_y0;
  wire f_u_cla12_and492_f_u_cla12_and491_y0;
  wire f_u_cla12_and492_f_u_cla12_and490_y0;
  wire f_u_cla12_and492_y0;
  wire f_u_cla12_and493_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and493_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and493_y0;
  wire f_u_cla12_and494_f_u_cla12_and493_y0;
  wire f_u_cla12_and494_f_u_cla12_and492_y0;
  wire f_u_cla12_and494_y0;
  wire f_u_cla12_and495_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and495_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and495_y0;
  wire f_u_cla12_and496_f_u_cla12_and495_y0;
  wire f_u_cla12_and496_f_u_cla12_and494_y0;
  wire f_u_cla12_and496_y0;
  wire f_u_cla12_and497_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and497_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and497_y0;
  wire f_u_cla12_and498_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and498_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and498_y0;
  wire f_u_cla12_and499_f_u_cla12_and498_y0;
  wire f_u_cla12_and499_f_u_cla12_and497_y0;
  wire f_u_cla12_and499_y0;
  wire f_u_cla12_and500_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and500_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and500_y0;
  wire f_u_cla12_and501_f_u_cla12_and500_y0;
  wire f_u_cla12_and501_f_u_cla12_and499_y0;
  wire f_u_cla12_and501_y0;
  wire f_u_cla12_and502_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and502_f_u_cla12_pg_logic8_y1;
  wire f_u_cla12_and502_y0;
  wire f_u_cla12_and503_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and503_f_u_cla12_pg_logic8_y1;
  wire f_u_cla12_and503_y0;
  wire f_u_cla12_and504_f_u_cla12_and503_y0;
  wire f_u_cla12_and504_f_u_cla12_and502_y0;
  wire f_u_cla12_and504_y0;
  wire f_u_cla12_and505_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and505_f_u_cla12_pg_logic9_y1;
  wire f_u_cla12_and505_y0;
  wire f_u_cla12_or55_f_u_cla12_and505_y0;
  wire f_u_cla12_or55_f_u_cla12_and405_y0;
  wire f_u_cla12_or55_y0;
  wire f_u_cla12_or56_f_u_cla12_or55_y0;
  wire f_u_cla12_or56_f_u_cla12_and424_y0;
  wire f_u_cla12_or56_y0;
  wire f_u_cla12_or57_f_u_cla12_or56_y0;
  wire f_u_cla12_or57_f_u_cla12_and441_y0;
  wire f_u_cla12_or57_y0;
  wire f_u_cla12_or58_f_u_cla12_or57_y0;
  wire f_u_cla12_or58_f_u_cla12_and456_y0;
  wire f_u_cla12_or58_y0;
  wire f_u_cla12_or59_f_u_cla12_or58_y0;
  wire f_u_cla12_or59_f_u_cla12_and469_y0;
  wire f_u_cla12_or59_y0;
  wire f_u_cla12_or60_f_u_cla12_or59_y0;
  wire f_u_cla12_or60_f_u_cla12_and480_y0;
  wire f_u_cla12_or60_y0;
  wire f_u_cla12_or61_f_u_cla12_or60_y0;
  wire f_u_cla12_or61_f_u_cla12_and489_y0;
  wire f_u_cla12_or61_y0;
  wire f_u_cla12_or62_f_u_cla12_or61_y0;
  wire f_u_cla12_or62_f_u_cla12_and496_y0;
  wire f_u_cla12_or62_y0;
  wire f_u_cla12_or63_f_u_cla12_or62_y0;
  wire f_u_cla12_or63_f_u_cla12_and501_y0;
  wire f_u_cla12_or63_y0;
  wire f_u_cla12_or64_f_u_cla12_or63_y0;
  wire f_u_cla12_or64_f_u_cla12_and504_y0;
  wire f_u_cla12_or64_y0;
  wire f_u_cla12_or65_f_u_cla12_pg_logic10_y1;
  wire f_u_cla12_or65_f_u_cla12_or64_y0;
  wire f_u_cla12_or65_y0;
  wire f_u_cla12_pg_logic11_a_11;
  wire f_u_cla12_pg_logic11_b_11;
  wire f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_pg_logic11_y1;
  wire f_u_cla12_pg_logic11_y2;
  wire f_u_cla12_xor11_f_u_cla12_pg_logic11_y2;
  wire f_u_cla12_xor11_f_u_cla12_or65_y0;
  wire f_u_cla12_xor11_y0;
  wire f_u_cla12_and506_f_u_cla12_pg_logic0_y0;
  wire f_u_cla12_and506_constant_wire_0;
  wire f_u_cla12_and506_y0;
  wire f_u_cla12_and507_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and507_constant_wire_0;
  wire f_u_cla12_and507_y0;
  wire f_u_cla12_and508_f_u_cla12_and507_y0;
  wire f_u_cla12_and508_f_u_cla12_and506_y0;
  wire f_u_cla12_and508_y0;
  wire f_u_cla12_and509_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and509_constant_wire_0;
  wire f_u_cla12_and509_y0;
  wire f_u_cla12_and510_f_u_cla12_and509_y0;
  wire f_u_cla12_and510_f_u_cla12_and508_y0;
  wire f_u_cla12_and510_y0;
  wire f_u_cla12_and511_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and511_constant_wire_0;
  wire f_u_cla12_and511_y0;
  wire f_u_cla12_and512_f_u_cla12_and511_y0;
  wire f_u_cla12_and512_f_u_cla12_and510_y0;
  wire f_u_cla12_and512_y0;
  wire f_u_cla12_and513_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and513_constant_wire_0;
  wire f_u_cla12_and513_y0;
  wire f_u_cla12_and514_f_u_cla12_and513_y0;
  wire f_u_cla12_and514_f_u_cla12_and512_y0;
  wire f_u_cla12_and514_y0;
  wire f_u_cla12_and515_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and515_constant_wire_0;
  wire f_u_cla12_and515_y0;
  wire f_u_cla12_and516_f_u_cla12_and515_y0;
  wire f_u_cla12_and516_f_u_cla12_and514_y0;
  wire f_u_cla12_and516_y0;
  wire f_u_cla12_and517_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and517_constant_wire_0;
  wire f_u_cla12_and517_y0;
  wire f_u_cla12_and518_f_u_cla12_and517_y0;
  wire f_u_cla12_and518_f_u_cla12_and516_y0;
  wire f_u_cla12_and518_y0;
  wire f_u_cla12_and519_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and519_constant_wire_0;
  wire f_u_cla12_and519_y0;
  wire f_u_cla12_and520_f_u_cla12_and519_y0;
  wire f_u_cla12_and520_f_u_cla12_and518_y0;
  wire f_u_cla12_and520_y0;
  wire f_u_cla12_and521_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and521_constant_wire_0;
  wire f_u_cla12_and521_y0;
  wire f_u_cla12_and522_f_u_cla12_and521_y0;
  wire f_u_cla12_and522_f_u_cla12_and520_y0;
  wire f_u_cla12_and522_y0;
  wire f_u_cla12_and523_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and523_constant_wire_0;
  wire f_u_cla12_and523_y0;
  wire f_u_cla12_and524_f_u_cla12_and523_y0;
  wire f_u_cla12_and524_f_u_cla12_and522_y0;
  wire f_u_cla12_and524_y0;
  wire f_u_cla12_and525_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and525_constant_wire_0;
  wire f_u_cla12_and525_y0;
  wire f_u_cla12_and526_f_u_cla12_and525_y0;
  wire f_u_cla12_and526_f_u_cla12_and524_y0;
  wire f_u_cla12_and526_y0;
  wire f_u_cla12_and527_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and527_constant_wire_0;
  wire f_u_cla12_and527_y0;
  wire f_u_cla12_and528_f_u_cla12_and527_y0;
  wire f_u_cla12_and528_f_u_cla12_and526_y0;
  wire f_u_cla12_and528_y0;
  wire f_u_cla12_and529_f_u_cla12_pg_logic1_y0;
  wire f_u_cla12_and529_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and529_y0;
  wire f_u_cla12_and530_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and530_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and530_y0;
  wire f_u_cla12_and531_f_u_cla12_and530_y0;
  wire f_u_cla12_and531_f_u_cla12_and529_y0;
  wire f_u_cla12_and531_y0;
  wire f_u_cla12_and532_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and532_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and532_y0;
  wire f_u_cla12_and533_f_u_cla12_and532_y0;
  wire f_u_cla12_and533_f_u_cla12_and531_y0;
  wire f_u_cla12_and533_y0;
  wire f_u_cla12_and534_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and534_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and534_y0;
  wire f_u_cla12_and535_f_u_cla12_and534_y0;
  wire f_u_cla12_and535_f_u_cla12_and533_y0;
  wire f_u_cla12_and535_y0;
  wire f_u_cla12_and536_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and536_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and536_y0;
  wire f_u_cla12_and537_f_u_cla12_and536_y0;
  wire f_u_cla12_and537_f_u_cla12_and535_y0;
  wire f_u_cla12_and537_y0;
  wire f_u_cla12_and538_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and538_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and538_y0;
  wire f_u_cla12_and539_f_u_cla12_and538_y0;
  wire f_u_cla12_and539_f_u_cla12_and537_y0;
  wire f_u_cla12_and539_y0;
  wire f_u_cla12_and540_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and540_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and540_y0;
  wire f_u_cla12_and541_f_u_cla12_and540_y0;
  wire f_u_cla12_and541_f_u_cla12_and539_y0;
  wire f_u_cla12_and541_y0;
  wire f_u_cla12_and542_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and542_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and542_y0;
  wire f_u_cla12_and543_f_u_cla12_and542_y0;
  wire f_u_cla12_and543_f_u_cla12_and541_y0;
  wire f_u_cla12_and543_y0;
  wire f_u_cla12_and544_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and544_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and544_y0;
  wire f_u_cla12_and545_f_u_cla12_and544_y0;
  wire f_u_cla12_and545_f_u_cla12_and543_y0;
  wire f_u_cla12_and545_y0;
  wire f_u_cla12_and546_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and546_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and546_y0;
  wire f_u_cla12_and547_f_u_cla12_and546_y0;
  wire f_u_cla12_and547_f_u_cla12_and545_y0;
  wire f_u_cla12_and547_y0;
  wire f_u_cla12_and548_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and548_f_u_cla12_pg_logic0_y1;
  wire f_u_cla12_and548_y0;
  wire f_u_cla12_and549_f_u_cla12_and548_y0;
  wire f_u_cla12_and549_f_u_cla12_and547_y0;
  wire f_u_cla12_and549_y0;
  wire f_u_cla12_and550_f_u_cla12_pg_logic2_y0;
  wire f_u_cla12_and550_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and550_y0;
  wire f_u_cla12_and551_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and551_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and551_y0;
  wire f_u_cla12_and552_f_u_cla12_and551_y0;
  wire f_u_cla12_and552_f_u_cla12_and550_y0;
  wire f_u_cla12_and552_y0;
  wire f_u_cla12_and553_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and553_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and553_y0;
  wire f_u_cla12_and554_f_u_cla12_and553_y0;
  wire f_u_cla12_and554_f_u_cla12_and552_y0;
  wire f_u_cla12_and554_y0;
  wire f_u_cla12_and555_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and555_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and555_y0;
  wire f_u_cla12_and556_f_u_cla12_and555_y0;
  wire f_u_cla12_and556_f_u_cla12_and554_y0;
  wire f_u_cla12_and556_y0;
  wire f_u_cla12_and557_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and557_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and557_y0;
  wire f_u_cla12_and558_f_u_cla12_and557_y0;
  wire f_u_cla12_and558_f_u_cla12_and556_y0;
  wire f_u_cla12_and558_y0;
  wire f_u_cla12_and559_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and559_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and559_y0;
  wire f_u_cla12_and560_f_u_cla12_and559_y0;
  wire f_u_cla12_and560_f_u_cla12_and558_y0;
  wire f_u_cla12_and560_y0;
  wire f_u_cla12_and561_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and561_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and561_y0;
  wire f_u_cla12_and562_f_u_cla12_and561_y0;
  wire f_u_cla12_and562_f_u_cla12_and560_y0;
  wire f_u_cla12_and562_y0;
  wire f_u_cla12_and563_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and563_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and563_y0;
  wire f_u_cla12_and564_f_u_cla12_and563_y0;
  wire f_u_cla12_and564_f_u_cla12_and562_y0;
  wire f_u_cla12_and564_y0;
  wire f_u_cla12_and565_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and565_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and565_y0;
  wire f_u_cla12_and566_f_u_cla12_and565_y0;
  wire f_u_cla12_and566_f_u_cla12_and564_y0;
  wire f_u_cla12_and566_y0;
  wire f_u_cla12_and567_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and567_f_u_cla12_pg_logic1_y1;
  wire f_u_cla12_and567_y0;
  wire f_u_cla12_and568_f_u_cla12_and567_y0;
  wire f_u_cla12_and568_f_u_cla12_and566_y0;
  wire f_u_cla12_and568_y0;
  wire f_u_cla12_and569_f_u_cla12_pg_logic3_y0;
  wire f_u_cla12_and569_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and569_y0;
  wire f_u_cla12_and570_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and570_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and570_y0;
  wire f_u_cla12_and571_f_u_cla12_and570_y0;
  wire f_u_cla12_and571_f_u_cla12_and569_y0;
  wire f_u_cla12_and571_y0;
  wire f_u_cla12_and572_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and572_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and572_y0;
  wire f_u_cla12_and573_f_u_cla12_and572_y0;
  wire f_u_cla12_and573_f_u_cla12_and571_y0;
  wire f_u_cla12_and573_y0;
  wire f_u_cla12_and574_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and574_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and574_y0;
  wire f_u_cla12_and575_f_u_cla12_and574_y0;
  wire f_u_cla12_and575_f_u_cla12_and573_y0;
  wire f_u_cla12_and575_y0;
  wire f_u_cla12_and576_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and576_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and576_y0;
  wire f_u_cla12_and577_f_u_cla12_and576_y0;
  wire f_u_cla12_and577_f_u_cla12_and575_y0;
  wire f_u_cla12_and577_y0;
  wire f_u_cla12_and578_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and578_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and578_y0;
  wire f_u_cla12_and579_f_u_cla12_and578_y0;
  wire f_u_cla12_and579_f_u_cla12_and577_y0;
  wire f_u_cla12_and579_y0;
  wire f_u_cla12_and580_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and580_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and580_y0;
  wire f_u_cla12_and581_f_u_cla12_and580_y0;
  wire f_u_cla12_and581_f_u_cla12_and579_y0;
  wire f_u_cla12_and581_y0;
  wire f_u_cla12_and582_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and582_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and582_y0;
  wire f_u_cla12_and583_f_u_cla12_and582_y0;
  wire f_u_cla12_and583_f_u_cla12_and581_y0;
  wire f_u_cla12_and583_y0;
  wire f_u_cla12_and584_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and584_f_u_cla12_pg_logic2_y1;
  wire f_u_cla12_and584_y0;
  wire f_u_cla12_and585_f_u_cla12_and584_y0;
  wire f_u_cla12_and585_f_u_cla12_and583_y0;
  wire f_u_cla12_and585_y0;
  wire f_u_cla12_and586_f_u_cla12_pg_logic4_y0;
  wire f_u_cla12_and586_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and586_y0;
  wire f_u_cla12_and587_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and587_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and587_y0;
  wire f_u_cla12_and588_f_u_cla12_and587_y0;
  wire f_u_cla12_and588_f_u_cla12_and586_y0;
  wire f_u_cla12_and588_y0;
  wire f_u_cla12_and589_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and589_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and589_y0;
  wire f_u_cla12_and590_f_u_cla12_and589_y0;
  wire f_u_cla12_and590_f_u_cla12_and588_y0;
  wire f_u_cla12_and590_y0;
  wire f_u_cla12_and591_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and591_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and591_y0;
  wire f_u_cla12_and592_f_u_cla12_and591_y0;
  wire f_u_cla12_and592_f_u_cla12_and590_y0;
  wire f_u_cla12_and592_y0;
  wire f_u_cla12_and593_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and593_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and593_y0;
  wire f_u_cla12_and594_f_u_cla12_and593_y0;
  wire f_u_cla12_and594_f_u_cla12_and592_y0;
  wire f_u_cla12_and594_y0;
  wire f_u_cla12_and595_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and595_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and595_y0;
  wire f_u_cla12_and596_f_u_cla12_and595_y0;
  wire f_u_cla12_and596_f_u_cla12_and594_y0;
  wire f_u_cla12_and596_y0;
  wire f_u_cla12_and597_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and597_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and597_y0;
  wire f_u_cla12_and598_f_u_cla12_and597_y0;
  wire f_u_cla12_and598_f_u_cla12_and596_y0;
  wire f_u_cla12_and598_y0;
  wire f_u_cla12_and599_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and599_f_u_cla12_pg_logic3_y1;
  wire f_u_cla12_and599_y0;
  wire f_u_cla12_and600_f_u_cla12_and599_y0;
  wire f_u_cla12_and600_f_u_cla12_and598_y0;
  wire f_u_cla12_and600_y0;
  wire f_u_cla12_and601_f_u_cla12_pg_logic5_y0;
  wire f_u_cla12_and601_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and601_y0;
  wire f_u_cla12_and602_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and602_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and602_y0;
  wire f_u_cla12_and603_f_u_cla12_and602_y0;
  wire f_u_cla12_and603_f_u_cla12_and601_y0;
  wire f_u_cla12_and603_y0;
  wire f_u_cla12_and604_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and604_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and604_y0;
  wire f_u_cla12_and605_f_u_cla12_and604_y0;
  wire f_u_cla12_and605_f_u_cla12_and603_y0;
  wire f_u_cla12_and605_y0;
  wire f_u_cla12_and606_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and606_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and606_y0;
  wire f_u_cla12_and607_f_u_cla12_and606_y0;
  wire f_u_cla12_and607_f_u_cla12_and605_y0;
  wire f_u_cla12_and607_y0;
  wire f_u_cla12_and608_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and608_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and608_y0;
  wire f_u_cla12_and609_f_u_cla12_and608_y0;
  wire f_u_cla12_and609_f_u_cla12_and607_y0;
  wire f_u_cla12_and609_y0;
  wire f_u_cla12_and610_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and610_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and610_y0;
  wire f_u_cla12_and611_f_u_cla12_and610_y0;
  wire f_u_cla12_and611_f_u_cla12_and609_y0;
  wire f_u_cla12_and611_y0;
  wire f_u_cla12_and612_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and612_f_u_cla12_pg_logic4_y1;
  wire f_u_cla12_and612_y0;
  wire f_u_cla12_and613_f_u_cla12_and612_y0;
  wire f_u_cla12_and613_f_u_cla12_and611_y0;
  wire f_u_cla12_and613_y0;
  wire f_u_cla12_and614_f_u_cla12_pg_logic6_y0;
  wire f_u_cla12_and614_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and614_y0;
  wire f_u_cla12_and615_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and615_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and615_y0;
  wire f_u_cla12_and616_f_u_cla12_and615_y0;
  wire f_u_cla12_and616_f_u_cla12_and614_y0;
  wire f_u_cla12_and616_y0;
  wire f_u_cla12_and617_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and617_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and617_y0;
  wire f_u_cla12_and618_f_u_cla12_and617_y0;
  wire f_u_cla12_and618_f_u_cla12_and616_y0;
  wire f_u_cla12_and618_y0;
  wire f_u_cla12_and619_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and619_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and619_y0;
  wire f_u_cla12_and620_f_u_cla12_and619_y0;
  wire f_u_cla12_and620_f_u_cla12_and618_y0;
  wire f_u_cla12_and620_y0;
  wire f_u_cla12_and621_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and621_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and621_y0;
  wire f_u_cla12_and622_f_u_cla12_and621_y0;
  wire f_u_cla12_and622_f_u_cla12_and620_y0;
  wire f_u_cla12_and622_y0;
  wire f_u_cla12_and623_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and623_f_u_cla12_pg_logic5_y1;
  wire f_u_cla12_and623_y0;
  wire f_u_cla12_and624_f_u_cla12_and623_y0;
  wire f_u_cla12_and624_f_u_cla12_and622_y0;
  wire f_u_cla12_and624_y0;
  wire f_u_cla12_and625_f_u_cla12_pg_logic7_y0;
  wire f_u_cla12_and625_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and625_y0;
  wire f_u_cla12_and626_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and626_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and626_y0;
  wire f_u_cla12_and627_f_u_cla12_and626_y0;
  wire f_u_cla12_and627_f_u_cla12_and625_y0;
  wire f_u_cla12_and627_y0;
  wire f_u_cla12_and628_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and628_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and628_y0;
  wire f_u_cla12_and629_f_u_cla12_and628_y0;
  wire f_u_cla12_and629_f_u_cla12_and627_y0;
  wire f_u_cla12_and629_y0;
  wire f_u_cla12_and630_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and630_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and630_y0;
  wire f_u_cla12_and631_f_u_cla12_and630_y0;
  wire f_u_cla12_and631_f_u_cla12_and629_y0;
  wire f_u_cla12_and631_y0;
  wire f_u_cla12_and632_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and632_f_u_cla12_pg_logic6_y1;
  wire f_u_cla12_and632_y0;
  wire f_u_cla12_and633_f_u_cla12_and632_y0;
  wire f_u_cla12_and633_f_u_cla12_and631_y0;
  wire f_u_cla12_and633_y0;
  wire f_u_cla12_and634_f_u_cla12_pg_logic8_y0;
  wire f_u_cla12_and634_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and634_y0;
  wire f_u_cla12_and635_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and635_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and635_y0;
  wire f_u_cla12_and636_f_u_cla12_and635_y0;
  wire f_u_cla12_and636_f_u_cla12_and634_y0;
  wire f_u_cla12_and636_y0;
  wire f_u_cla12_and637_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and637_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and637_y0;
  wire f_u_cla12_and638_f_u_cla12_and637_y0;
  wire f_u_cla12_and638_f_u_cla12_and636_y0;
  wire f_u_cla12_and638_y0;
  wire f_u_cla12_and639_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and639_f_u_cla12_pg_logic7_y1;
  wire f_u_cla12_and639_y0;
  wire f_u_cla12_and640_f_u_cla12_and639_y0;
  wire f_u_cla12_and640_f_u_cla12_and638_y0;
  wire f_u_cla12_and640_y0;
  wire f_u_cla12_and641_f_u_cla12_pg_logic9_y0;
  wire f_u_cla12_and641_f_u_cla12_pg_logic8_y1;
  wire f_u_cla12_and641_y0;
  wire f_u_cla12_and642_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and642_f_u_cla12_pg_logic8_y1;
  wire f_u_cla12_and642_y0;
  wire f_u_cla12_and643_f_u_cla12_and642_y0;
  wire f_u_cla12_and643_f_u_cla12_and641_y0;
  wire f_u_cla12_and643_y0;
  wire f_u_cla12_and644_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and644_f_u_cla12_pg_logic8_y1;
  wire f_u_cla12_and644_y0;
  wire f_u_cla12_and645_f_u_cla12_and644_y0;
  wire f_u_cla12_and645_f_u_cla12_and643_y0;
  wire f_u_cla12_and645_y0;
  wire f_u_cla12_and646_f_u_cla12_pg_logic10_y0;
  wire f_u_cla12_and646_f_u_cla12_pg_logic9_y1;
  wire f_u_cla12_and646_y0;
  wire f_u_cla12_and647_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and647_f_u_cla12_pg_logic9_y1;
  wire f_u_cla12_and647_y0;
  wire f_u_cla12_and648_f_u_cla12_and647_y0;
  wire f_u_cla12_and648_f_u_cla12_and646_y0;
  wire f_u_cla12_and648_y0;
  wire f_u_cla12_and649_f_u_cla12_pg_logic11_y0;
  wire f_u_cla12_and649_f_u_cla12_pg_logic10_y1;
  wire f_u_cla12_and649_y0;
  wire f_u_cla12_or66_f_u_cla12_and649_y0;
  wire f_u_cla12_or66_f_u_cla12_and528_y0;
  wire f_u_cla12_or66_y0;
  wire f_u_cla12_or67_f_u_cla12_or66_y0;
  wire f_u_cla12_or67_f_u_cla12_and549_y0;
  wire f_u_cla12_or67_y0;
  wire f_u_cla12_or68_f_u_cla12_or67_y0;
  wire f_u_cla12_or68_f_u_cla12_and568_y0;
  wire f_u_cla12_or68_y0;
  wire f_u_cla12_or69_f_u_cla12_or68_y0;
  wire f_u_cla12_or69_f_u_cla12_and585_y0;
  wire f_u_cla12_or69_y0;
  wire f_u_cla12_or70_f_u_cla12_or69_y0;
  wire f_u_cla12_or70_f_u_cla12_and600_y0;
  wire f_u_cla12_or70_y0;
  wire f_u_cla12_or71_f_u_cla12_or70_y0;
  wire f_u_cla12_or71_f_u_cla12_and613_y0;
  wire f_u_cla12_or71_y0;
  wire f_u_cla12_or72_f_u_cla12_or71_y0;
  wire f_u_cla12_or72_f_u_cla12_and624_y0;
  wire f_u_cla12_or72_y0;
  wire f_u_cla12_or73_f_u_cla12_or72_y0;
  wire f_u_cla12_or73_f_u_cla12_and633_y0;
  wire f_u_cla12_or73_y0;
  wire f_u_cla12_or74_f_u_cla12_or73_y0;
  wire f_u_cla12_or74_f_u_cla12_and640_y0;
  wire f_u_cla12_or74_y0;
  wire f_u_cla12_or75_f_u_cla12_or74_y0;
  wire f_u_cla12_or75_f_u_cla12_and645_y0;
  wire f_u_cla12_or75_y0;
  wire f_u_cla12_or76_f_u_cla12_or75_y0;
  wire f_u_cla12_or76_f_u_cla12_and648_y0;
  wire f_u_cla12_or76_y0;
  wire f_u_cla12_or77_f_u_cla12_pg_logic11_y1;
  wire f_u_cla12_or77_f_u_cla12_or76_y0;
  wire f_u_cla12_or77_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign constant_wire_value_0_a_0 = a_0;
  assign constant_wire_value_0_b_0 = b_0;
  assign constant_wire_value_0_y0 = constant_wire_value_0_a_0 ^ constant_wire_value_0_b_0;
  assign constant_wire_value_0_y1 = ~(constant_wire_value_0_a_0 ^ constant_wire_value_0_b_0);
  assign constant_wire_0 = ~(constant_wire_value_0_y0 | constant_wire_value_0_y1);
  assign f_u_cla12_pg_logic0_a_0 = a_0;
  assign f_u_cla12_pg_logic0_b_0 = b_0;
  assign f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_a_0 | f_u_cla12_pg_logic0_b_0;
  assign f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_a_0 & f_u_cla12_pg_logic0_b_0;
  assign f_u_cla12_pg_logic0_y2 = f_u_cla12_pg_logic0_a_0 ^ f_u_cla12_pg_logic0_b_0;
  assign f_u_cla12_xor0_f_u_cla12_pg_logic0_y2 = f_u_cla12_pg_logic0_y2;
  assign f_u_cla12_xor0_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_xor0_y0 = f_u_cla12_xor0_f_u_cla12_pg_logic0_y2 ^ f_u_cla12_xor0_constant_wire_0;
  assign f_u_cla12_and0_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and0_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and0_y0 = f_u_cla12_and0_f_u_cla12_pg_logic0_y0 & f_u_cla12_and0_constant_wire_0;
  assign f_u_cla12_or0_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_or0_f_u_cla12_and0_y0 = f_u_cla12_and0_y0;
  assign f_u_cla12_or0_y0 = f_u_cla12_or0_f_u_cla12_pg_logic0_y1 | f_u_cla12_or0_f_u_cla12_and0_y0;
  assign f_u_cla12_pg_logic1_a_1 = a_1;
  assign f_u_cla12_pg_logic1_b_1 = b_1;
  assign f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_a_1 | f_u_cla12_pg_logic1_b_1;
  assign f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_a_1 & f_u_cla12_pg_logic1_b_1;
  assign f_u_cla12_pg_logic1_y2 = f_u_cla12_pg_logic1_a_1 ^ f_u_cla12_pg_logic1_b_1;
  assign f_u_cla12_xor1_f_u_cla12_pg_logic1_y2 = f_u_cla12_pg_logic1_y2;
  assign f_u_cla12_xor1_f_u_cla12_or0_y0 = f_u_cla12_or0_y0;
  assign f_u_cla12_xor1_y0 = f_u_cla12_xor1_f_u_cla12_pg_logic1_y2 ^ f_u_cla12_xor1_f_u_cla12_or0_y0;
  assign f_u_cla12_and1_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and1_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and1_y0 = f_u_cla12_and1_f_u_cla12_pg_logic0_y0 & f_u_cla12_and1_constant_wire_0;
  assign f_u_cla12_and2_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and2_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and2_y0 = f_u_cla12_and2_f_u_cla12_pg_logic1_y0 & f_u_cla12_and2_constant_wire_0;
  assign f_u_cla12_and3_f_u_cla12_and2_y0 = f_u_cla12_and2_y0;
  assign f_u_cla12_and3_f_u_cla12_and1_y0 = f_u_cla12_and1_y0;
  assign f_u_cla12_and3_y0 = f_u_cla12_and3_f_u_cla12_and2_y0 & f_u_cla12_and3_f_u_cla12_and1_y0;
  assign f_u_cla12_and4_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and4_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and4_y0 = f_u_cla12_and4_f_u_cla12_pg_logic1_y0 & f_u_cla12_and4_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_or1_f_u_cla12_and4_y0 = f_u_cla12_and4_y0;
  assign f_u_cla12_or1_f_u_cla12_and3_y0 = f_u_cla12_and3_y0;
  assign f_u_cla12_or1_y0 = f_u_cla12_or1_f_u_cla12_and4_y0 | f_u_cla12_or1_f_u_cla12_and3_y0;
  assign f_u_cla12_or2_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_or2_f_u_cla12_or1_y0 = f_u_cla12_or1_y0;
  assign f_u_cla12_or2_y0 = f_u_cla12_or2_f_u_cla12_pg_logic1_y1 | f_u_cla12_or2_f_u_cla12_or1_y0;
  assign f_u_cla12_pg_logic2_a_2 = a_2;
  assign f_u_cla12_pg_logic2_b_2 = b_2;
  assign f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_a_2 | f_u_cla12_pg_logic2_b_2;
  assign f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_a_2 & f_u_cla12_pg_logic2_b_2;
  assign f_u_cla12_pg_logic2_y2 = f_u_cla12_pg_logic2_a_2 ^ f_u_cla12_pg_logic2_b_2;
  assign f_u_cla12_xor2_f_u_cla12_pg_logic2_y2 = f_u_cla12_pg_logic2_y2;
  assign f_u_cla12_xor2_f_u_cla12_or2_y0 = f_u_cla12_or2_y0;
  assign f_u_cla12_xor2_y0 = f_u_cla12_xor2_f_u_cla12_pg_logic2_y2 ^ f_u_cla12_xor2_f_u_cla12_or2_y0;
  assign f_u_cla12_and5_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and5_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and5_y0 = f_u_cla12_and5_f_u_cla12_pg_logic0_y0 & f_u_cla12_and5_constant_wire_0;
  assign f_u_cla12_and6_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and6_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and6_y0 = f_u_cla12_and6_f_u_cla12_pg_logic1_y0 & f_u_cla12_and6_constant_wire_0;
  assign f_u_cla12_and7_f_u_cla12_and6_y0 = f_u_cla12_and6_y0;
  assign f_u_cla12_and7_f_u_cla12_and5_y0 = f_u_cla12_and5_y0;
  assign f_u_cla12_and7_y0 = f_u_cla12_and7_f_u_cla12_and6_y0 & f_u_cla12_and7_f_u_cla12_and5_y0;
  assign f_u_cla12_and8_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and8_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and8_y0 = f_u_cla12_and8_f_u_cla12_pg_logic2_y0 & f_u_cla12_and8_constant_wire_0;
  assign f_u_cla12_and9_f_u_cla12_and8_y0 = f_u_cla12_and8_y0;
  assign f_u_cla12_and9_f_u_cla12_and7_y0 = f_u_cla12_and7_y0;
  assign f_u_cla12_and9_y0 = f_u_cla12_and9_f_u_cla12_and8_y0 & f_u_cla12_and9_f_u_cla12_and7_y0;
  assign f_u_cla12_and10_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and10_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and10_y0 = f_u_cla12_and10_f_u_cla12_pg_logic1_y0 & f_u_cla12_and10_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and11_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and11_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and11_y0 = f_u_cla12_and11_f_u_cla12_pg_logic2_y0 & f_u_cla12_and11_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and12_f_u_cla12_and11_y0 = f_u_cla12_and11_y0;
  assign f_u_cla12_and12_f_u_cla12_and10_y0 = f_u_cla12_and10_y0;
  assign f_u_cla12_and12_y0 = f_u_cla12_and12_f_u_cla12_and11_y0 & f_u_cla12_and12_f_u_cla12_and10_y0;
  assign f_u_cla12_and13_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and13_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and13_y0 = f_u_cla12_and13_f_u_cla12_pg_logic2_y0 & f_u_cla12_and13_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_or3_f_u_cla12_and13_y0 = f_u_cla12_and13_y0;
  assign f_u_cla12_or3_f_u_cla12_and9_y0 = f_u_cla12_and9_y0;
  assign f_u_cla12_or3_y0 = f_u_cla12_or3_f_u_cla12_and13_y0 | f_u_cla12_or3_f_u_cla12_and9_y0;
  assign f_u_cla12_or4_f_u_cla12_or3_y0 = f_u_cla12_or3_y0;
  assign f_u_cla12_or4_f_u_cla12_and12_y0 = f_u_cla12_and12_y0;
  assign f_u_cla12_or4_y0 = f_u_cla12_or4_f_u_cla12_or3_y0 | f_u_cla12_or4_f_u_cla12_and12_y0;
  assign f_u_cla12_or5_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_or5_f_u_cla12_or4_y0 = f_u_cla12_or4_y0;
  assign f_u_cla12_or5_y0 = f_u_cla12_or5_f_u_cla12_pg_logic2_y1 | f_u_cla12_or5_f_u_cla12_or4_y0;
  assign f_u_cla12_pg_logic3_a_3 = a_3;
  assign f_u_cla12_pg_logic3_b_3 = b_3;
  assign f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_a_3 | f_u_cla12_pg_logic3_b_3;
  assign f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_a_3 & f_u_cla12_pg_logic3_b_3;
  assign f_u_cla12_pg_logic3_y2 = f_u_cla12_pg_logic3_a_3 ^ f_u_cla12_pg_logic3_b_3;
  assign f_u_cla12_xor3_f_u_cla12_pg_logic3_y2 = f_u_cla12_pg_logic3_y2;
  assign f_u_cla12_xor3_f_u_cla12_or5_y0 = f_u_cla12_or5_y0;
  assign f_u_cla12_xor3_y0 = f_u_cla12_xor3_f_u_cla12_pg_logic3_y2 ^ f_u_cla12_xor3_f_u_cla12_or5_y0;
  assign f_u_cla12_and14_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and14_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and14_y0 = f_u_cla12_and14_f_u_cla12_pg_logic0_y0 & f_u_cla12_and14_constant_wire_0;
  assign f_u_cla12_and15_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and15_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and15_y0 = f_u_cla12_and15_f_u_cla12_pg_logic1_y0 & f_u_cla12_and15_constant_wire_0;
  assign f_u_cla12_and16_f_u_cla12_and15_y0 = f_u_cla12_and15_y0;
  assign f_u_cla12_and16_f_u_cla12_and14_y0 = f_u_cla12_and14_y0;
  assign f_u_cla12_and16_y0 = f_u_cla12_and16_f_u_cla12_and15_y0 & f_u_cla12_and16_f_u_cla12_and14_y0;
  assign f_u_cla12_and17_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and17_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and17_y0 = f_u_cla12_and17_f_u_cla12_pg_logic2_y0 & f_u_cla12_and17_constant_wire_0;
  assign f_u_cla12_and18_f_u_cla12_and17_y0 = f_u_cla12_and17_y0;
  assign f_u_cla12_and18_f_u_cla12_and16_y0 = f_u_cla12_and16_y0;
  assign f_u_cla12_and18_y0 = f_u_cla12_and18_f_u_cla12_and17_y0 & f_u_cla12_and18_f_u_cla12_and16_y0;
  assign f_u_cla12_and19_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and19_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and19_y0 = f_u_cla12_and19_f_u_cla12_pg_logic3_y0 & f_u_cla12_and19_constant_wire_0;
  assign f_u_cla12_and20_f_u_cla12_and19_y0 = f_u_cla12_and19_y0;
  assign f_u_cla12_and20_f_u_cla12_and18_y0 = f_u_cla12_and18_y0;
  assign f_u_cla12_and20_y0 = f_u_cla12_and20_f_u_cla12_and19_y0 & f_u_cla12_and20_f_u_cla12_and18_y0;
  assign f_u_cla12_and21_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and21_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and21_y0 = f_u_cla12_and21_f_u_cla12_pg_logic1_y0 & f_u_cla12_and21_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and22_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and22_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and22_y0 = f_u_cla12_and22_f_u_cla12_pg_logic2_y0 & f_u_cla12_and22_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and23_f_u_cla12_and22_y0 = f_u_cla12_and22_y0;
  assign f_u_cla12_and23_f_u_cla12_and21_y0 = f_u_cla12_and21_y0;
  assign f_u_cla12_and23_y0 = f_u_cla12_and23_f_u_cla12_and22_y0 & f_u_cla12_and23_f_u_cla12_and21_y0;
  assign f_u_cla12_and24_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and24_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and24_y0 = f_u_cla12_and24_f_u_cla12_pg_logic3_y0 & f_u_cla12_and24_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and25_f_u_cla12_and24_y0 = f_u_cla12_and24_y0;
  assign f_u_cla12_and25_f_u_cla12_and23_y0 = f_u_cla12_and23_y0;
  assign f_u_cla12_and25_y0 = f_u_cla12_and25_f_u_cla12_and24_y0 & f_u_cla12_and25_f_u_cla12_and23_y0;
  assign f_u_cla12_and26_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and26_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and26_y0 = f_u_cla12_and26_f_u_cla12_pg_logic2_y0 & f_u_cla12_and26_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and27_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and27_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and27_y0 = f_u_cla12_and27_f_u_cla12_pg_logic3_y0 & f_u_cla12_and27_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and28_f_u_cla12_and27_y0 = f_u_cla12_and27_y0;
  assign f_u_cla12_and28_f_u_cla12_and26_y0 = f_u_cla12_and26_y0;
  assign f_u_cla12_and28_y0 = f_u_cla12_and28_f_u_cla12_and27_y0 & f_u_cla12_and28_f_u_cla12_and26_y0;
  assign f_u_cla12_and29_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and29_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and29_y0 = f_u_cla12_and29_f_u_cla12_pg_logic3_y0 & f_u_cla12_and29_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_or6_f_u_cla12_and29_y0 = f_u_cla12_and29_y0;
  assign f_u_cla12_or6_f_u_cla12_and20_y0 = f_u_cla12_and20_y0;
  assign f_u_cla12_or6_y0 = f_u_cla12_or6_f_u_cla12_and29_y0 | f_u_cla12_or6_f_u_cla12_and20_y0;
  assign f_u_cla12_or7_f_u_cla12_or6_y0 = f_u_cla12_or6_y0;
  assign f_u_cla12_or7_f_u_cla12_and25_y0 = f_u_cla12_and25_y0;
  assign f_u_cla12_or7_y0 = f_u_cla12_or7_f_u_cla12_or6_y0 | f_u_cla12_or7_f_u_cla12_and25_y0;
  assign f_u_cla12_or8_f_u_cla12_or7_y0 = f_u_cla12_or7_y0;
  assign f_u_cla12_or8_f_u_cla12_and28_y0 = f_u_cla12_and28_y0;
  assign f_u_cla12_or8_y0 = f_u_cla12_or8_f_u_cla12_or7_y0 | f_u_cla12_or8_f_u_cla12_and28_y0;
  assign f_u_cla12_or9_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_or9_f_u_cla12_or8_y0 = f_u_cla12_or8_y0;
  assign f_u_cla12_or9_y0 = f_u_cla12_or9_f_u_cla12_pg_logic3_y1 | f_u_cla12_or9_f_u_cla12_or8_y0;
  assign f_u_cla12_pg_logic4_a_4 = a_4;
  assign f_u_cla12_pg_logic4_b_4 = b_4;
  assign f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_a_4 | f_u_cla12_pg_logic4_b_4;
  assign f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_a_4 & f_u_cla12_pg_logic4_b_4;
  assign f_u_cla12_pg_logic4_y2 = f_u_cla12_pg_logic4_a_4 ^ f_u_cla12_pg_logic4_b_4;
  assign f_u_cla12_xor4_f_u_cla12_pg_logic4_y2 = f_u_cla12_pg_logic4_y2;
  assign f_u_cla12_xor4_f_u_cla12_or9_y0 = f_u_cla12_or9_y0;
  assign f_u_cla12_xor4_y0 = f_u_cla12_xor4_f_u_cla12_pg_logic4_y2 ^ f_u_cla12_xor4_f_u_cla12_or9_y0;
  assign f_u_cla12_and30_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and30_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and30_y0 = f_u_cla12_and30_f_u_cla12_pg_logic0_y0 & f_u_cla12_and30_constant_wire_0;
  assign f_u_cla12_and31_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and31_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and31_y0 = f_u_cla12_and31_f_u_cla12_pg_logic1_y0 & f_u_cla12_and31_constant_wire_0;
  assign f_u_cla12_and32_f_u_cla12_and31_y0 = f_u_cla12_and31_y0;
  assign f_u_cla12_and32_f_u_cla12_and30_y0 = f_u_cla12_and30_y0;
  assign f_u_cla12_and32_y0 = f_u_cla12_and32_f_u_cla12_and31_y0 & f_u_cla12_and32_f_u_cla12_and30_y0;
  assign f_u_cla12_and33_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and33_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and33_y0 = f_u_cla12_and33_f_u_cla12_pg_logic2_y0 & f_u_cla12_and33_constant_wire_0;
  assign f_u_cla12_and34_f_u_cla12_and33_y0 = f_u_cla12_and33_y0;
  assign f_u_cla12_and34_f_u_cla12_and32_y0 = f_u_cla12_and32_y0;
  assign f_u_cla12_and34_y0 = f_u_cla12_and34_f_u_cla12_and33_y0 & f_u_cla12_and34_f_u_cla12_and32_y0;
  assign f_u_cla12_and35_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and35_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and35_y0 = f_u_cla12_and35_f_u_cla12_pg_logic3_y0 & f_u_cla12_and35_constant_wire_0;
  assign f_u_cla12_and36_f_u_cla12_and35_y0 = f_u_cla12_and35_y0;
  assign f_u_cla12_and36_f_u_cla12_and34_y0 = f_u_cla12_and34_y0;
  assign f_u_cla12_and36_y0 = f_u_cla12_and36_f_u_cla12_and35_y0 & f_u_cla12_and36_f_u_cla12_and34_y0;
  assign f_u_cla12_and37_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and37_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and37_y0 = f_u_cla12_and37_f_u_cla12_pg_logic4_y0 & f_u_cla12_and37_constant_wire_0;
  assign f_u_cla12_and38_f_u_cla12_and37_y0 = f_u_cla12_and37_y0;
  assign f_u_cla12_and38_f_u_cla12_and36_y0 = f_u_cla12_and36_y0;
  assign f_u_cla12_and38_y0 = f_u_cla12_and38_f_u_cla12_and37_y0 & f_u_cla12_and38_f_u_cla12_and36_y0;
  assign f_u_cla12_and39_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and39_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and39_y0 = f_u_cla12_and39_f_u_cla12_pg_logic1_y0 & f_u_cla12_and39_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and40_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and40_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and40_y0 = f_u_cla12_and40_f_u_cla12_pg_logic2_y0 & f_u_cla12_and40_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and41_f_u_cla12_and40_y0 = f_u_cla12_and40_y0;
  assign f_u_cla12_and41_f_u_cla12_and39_y0 = f_u_cla12_and39_y0;
  assign f_u_cla12_and41_y0 = f_u_cla12_and41_f_u_cla12_and40_y0 & f_u_cla12_and41_f_u_cla12_and39_y0;
  assign f_u_cla12_and42_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and42_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and42_y0 = f_u_cla12_and42_f_u_cla12_pg_logic3_y0 & f_u_cla12_and42_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and43_f_u_cla12_and42_y0 = f_u_cla12_and42_y0;
  assign f_u_cla12_and43_f_u_cla12_and41_y0 = f_u_cla12_and41_y0;
  assign f_u_cla12_and43_y0 = f_u_cla12_and43_f_u_cla12_and42_y0 & f_u_cla12_and43_f_u_cla12_and41_y0;
  assign f_u_cla12_and44_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and44_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and44_y0 = f_u_cla12_and44_f_u_cla12_pg_logic4_y0 & f_u_cla12_and44_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and45_f_u_cla12_and44_y0 = f_u_cla12_and44_y0;
  assign f_u_cla12_and45_f_u_cla12_and43_y0 = f_u_cla12_and43_y0;
  assign f_u_cla12_and45_y0 = f_u_cla12_and45_f_u_cla12_and44_y0 & f_u_cla12_and45_f_u_cla12_and43_y0;
  assign f_u_cla12_and46_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and46_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and46_y0 = f_u_cla12_and46_f_u_cla12_pg_logic2_y0 & f_u_cla12_and46_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and47_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and47_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and47_y0 = f_u_cla12_and47_f_u_cla12_pg_logic3_y0 & f_u_cla12_and47_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and48_f_u_cla12_and47_y0 = f_u_cla12_and47_y0;
  assign f_u_cla12_and48_f_u_cla12_and46_y0 = f_u_cla12_and46_y0;
  assign f_u_cla12_and48_y0 = f_u_cla12_and48_f_u_cla12_and47_y0 & f_u_cla12_and48_f_u_cla12_and46_y0;
  assign f_u_cla12_and49_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and49_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and49_y0 = f_u_cla12_and49_f_u_cla12_pg_logic4_y0 & f_u_cla12_and49_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and50_f_u_cla12_and49_y0 = f_u_cla12_and49_y0;
  assign f_u_cla12_and50_f_u_cla12_and48_y0 = f_u_cla12_and48_y0;
  assign f_u_cla12_and50_y0 = f_u_cla12_and50_f_u_cla12_and49_y0 & f_u_cla12_and50_f_u_cla12_and48_y0;
  assign f_u_cla12_and51_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and51_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and51_y0 = f_u_cla12_and51_f_u_cla12_pg_logic3_y0 & f_u_cla12_and51_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and52_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and52_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and52_y0 = f_u_cla12_and52_f_u_cla12_pg_logic4_y0 & f_u_cla12_and52_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and53_f_u_cla12_and52_y0 = f_u_cla12_and52_y0;
  assign f_u_cla12_and53_f_u_cla12_and51_y0 = f_u_cla12_and51_y0;
  assign f_u_cla12_and53_y0 = f_u_cla12_and53_f_u_cla12_and52_y0 & f_u_cla12_and53_f_u_cla12_and51_y0;
  assign f_u_cla12_and54_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and54_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and54_y0 = f_u_cla12_and54_f_u_cla12_pg_logic4_y0 & f_u_cla12_and54_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_or10_f_u_cla12_and54_y0 = f_u_cla12_and54_y0;
  assign f_u_cla12_or10_f_u_cla12_and38_y0 = f_u_cla12_and38_y0;
  assign f_u_cla12_or10_y0 = f_u_cla12_or10_f_u_cla12_and54_y0 | f_u_cla12_or10_f_u_cla12_and38_y0;
  assign f_u_cla12_or11_f_u_cla12_or10_y0 = f_u_cla12_or10_y0;
  assign f_u_cla12_or11_f_u_cla12_and45_y0 = f_u_cla12_and45_y0;
  assign f_u_cla12_or11_y0 = f_u_cla12_or11_f_u_cla12_or10_y0 | f_u_cla12_or11_f_u_cla12_and45_y0;
  assign f_u_cla12_or12_f_u_cla12_or11_y0 = f_u_cla12_or11_y0;
  assign f_u_cla12_or12_f_u_cla12_and50_y0 = f_u_cla12_and50_y0;
  assign f_u_cla12_or12_y0 = f_u_cla12_or12_f_u_cla12_or11_y0 | f_u_cla12_or12_f_u_cla12_and50_y0;
  assign f_u_cla12_or13_f_u_cla12_or12_y0 = f_u_cla12_or12_y0;
  assign f_u_cla12_or13_f_u_cla12_and53_y0 = f_u_cla12_and53_y0;
  assign f_u_cla12_or13_y0 = f_u_cla12_or13_f_u_cla12_or12_y0 | f_u_cla12_or13_f_u_cla12_and53_y0;
  assign f_u_cla12_or14_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_or14_f_u_cla12_or13_y0 = f_u_cla12_or13_y0;
  assign f_u_cla12_or14_y0 = f_u_cla12_or14_f_u_cla12_pg_logic4_y1 | f_u_cla12_or14_f_u_cla12_or13_y0;
  assign f_u_cla12_pg_logic5_a_5 = a_5;
  assign f_u_cla12_pg_logic5_b_5 = b_5;
  assign f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_a_5 | f_u_cla12_pg_logic5_b_5;
  assign f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_a_5 & f_u_cla12_pg_logic5_b_5;
  assign f_u_cla12_pg_logic5_y2 = f_u_cla12_pg_logic5_a_5 ^ f_u_cla12_pg_logic5_b_5;
  assign f_u_cla12_xor5_f_u_cla12_pg_logic5_y2 = f_u_cla12_pg_logic5_y2;
  assign f_u_cla12_xor5_f_u_cla12_or14_y0 = f_u_cla12_or14_y0;
  assign f_u_cla12_xor5_y0 = f_u_cla12_xor5_f_u_cla12_pg_logic5_y2 ^ f_u_cla12_xor5_f_u_cla12_or14_y0;
  assign f_u_cla12_and55_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and55_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and55_y0 = f_u_cla12_and55_f_u_cla12_pg_logic0_y0 & f_u_cla12_and55_constant_wire_0;
  assign f_u_cla12_and56_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and56_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and56_y0 = f_u_cla12_and56_f_u_cla12_pg_logic1_y0 & f_u_cla12_and56_constant_wire_0;
  assign f_u_cla12_and57_f_u_cla12_and56_y0 = f_u_cla12_and56_y0;
  assign f_u_cla12_and57_f_u_cla12_and55_y0 = f_u_cla12_and55_y0;
  assign f_u_cla12_and57_y0 = f_u_cla12_and57_f_u_cla12_and56_y0 & f_u_cla12_and57_f_u_cla12_and55_y0;
  assign f_u_cla12_and58_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and58_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and58_y0 = f_u_cla12_and58_f_u_cla12_pg_logic2_y0 & f_u_cla12_and58_constant_wire_0;
  assign f_u_cla12_and59_f_u_cla12_and58_y0 = f_u_cla12_and58_y0;
  assign f_u_cla12_and59_f_u_cla12_and57_y0 = f_u_cla12_and57_y0;
  assign f_u_cla12_and59_y0 = f_u_cla12_and59_f_u_cla12_and58_y0 & f_u_cla12_and59_f_u_cla12_and57_y0;
  assign f_u_cla12_and60_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and60_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and60_y0 = f_u_cla12_and60_f_u_cla12_pg_logic3_y0 & f_u_cla12_and60_constant_wire_0;
  assign f_u_cla12_and61_f_u_cla12_and60_y0 = f_u_cla12_and60_y0;
  assign f_u_cla12_and61_f_u_cla12_and59_y0 = f_u_cla12_and59_y0;
  assign f_u_cla12_and61_y0 = f_u_cla12_and61_f_u_cla12_and60_y0 & f_u_cla12_and61_f_u_cla12_and59_y0;
  assign f_u_cla12_and62_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and62_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and62_y0 = f_u_cla12_and62_f_u_cla12_pg_logic4_y0 & f_u_cla12_and62_constant_wire_0;
  assign f_u_cla12_and63_f_u_cla12_and62_y0 = f_u_cla12_and62_y0;
  assign f_u_cla12_and63_f_u_cla12_and61_y0 = f_u_cla12_and61_y0;
  assign f_u_cla12_and63_y0 = f_u_cla12_and63_f_u_cla12_and62_y0 & f_u_cla12_and63_f_u_cla12_and61_y0;
  assign f_u_cla12_and64_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and64_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and64_y0 = f_u_cla12_and64_f_u_cla12_pg_logic5_y0 & f_u_cla12_and64_constant_wire_0;
  assign f_u_cla12_and65_f_u_cla12_and64_y0 = f_u_cla12_and64_y0;
  assign f_u_cla12_and65_f_u_cla12_and63_y0 = f_u_cla12_and63_y0;
  assign f_u_cla12_and65_y0 = f_u_cla12_and65_f_u_cla12_and64_y0 & f_u_cla12_and65_f_u_cla12_and63_y0;
  assign f_u_cla12_and66_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and66_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and66_y0 = f_u_cla12_and66_f_u_cla12_pg_logic1_y0 & f_u_cla12_and66_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and67_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and67_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and67_y0 = f_u_cla12_and67_f_u_cla12_pg_logic2_y0 & f_u_cla12_and67_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and68_f_u_cla12_and67_y0 = f_u_cla12_and67_y0;
  assign f_u_cla12_and68_f_u_cla12_and66_y0 = f_u_cla12_and66_y0;
  assign f_u_cla12_and68_y0 = f_u_cla12_and68_f_u_cla12_and67_y0 & f_u_cla12_and68_f_u_cla12_and66_y0;
  assign f_u_cla12_and69_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and69_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and69_y0 = f_u_cla12_and69_f_u_cla12_pg_logic3_y0 & f_u_cla12_and69_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and70_f_u_cla12_and69_y0 = f_u_cla12_and69_y0;
  assign f_u_cla12_and70_f_u_cla12_and68_y0 = f_u_cla12_and68_y0;
  assign f_u_cla12_and70_y0 = f_u_cla12_and70_f_u_cla12_and69_y0 & f_u_cla12_and70_f_u_cla12_and68_y0;
  assign f_u_cla12_and71_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and71_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and71_y0 = f_u_cla12_and71_f_u_cla12_pg_logic4_y0 & f_u_cla12_and71_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and72_f_u_cla12_and71_y0 = f_u_cla12_and71_y0;
  assign f_u_cla12_and72_f_u_cla12_and70_y0 = f_u_cla12_and70_y0;
  assign f_u_cla12_and72_y0 = f_u_cla12_and72_f_u_cla12_and71_y0 & f_u_cla12_and72_f_u_cla12_and70_y0;
  assign f_u_cla12_and73_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and73_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and73_y0 = f_u_cla12_and73_f_u_cla12_pg_logic5_y0 & f_u_cla12_and73_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and74_f_u_cla12_and73_y0 = f_u_cla12_and73_y0;
  assign f_u_cla12_and74_f_u_cla12_and72_y0 = f_u_cla12_and72_y0;
  assign f_u_cla12_and74_y0 = f_u_cla12_and74_f_u_cla12_and73_y0 & f_u_cla12_and74_f_u_cla12_and72_y0;
  assign f_u_cla12_and75_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and75_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and75_y0 = f_u_cla12_and75_f_u_cla12_pg_logic2_y0 & f_u_cla12_and75_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and76_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and76_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and76_y0 = f_u_cla12_and76_f_u_cla12_pg_logic3_y0 & f_u_cla12_and76_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and77_f_u_cla12_and76_y0 = f_u_cla12_and76_y0;
  assign f_u_cla12_and77_f_u_cla12_and75_y0 = f_u_cla12_and75_y0;
  assign f_u_cla12_and77_y0 = f_u_cla12_and77_f_u_cla12_and76_y0 & f_u_cla12_and77_f_u_cla12_and75_y0;
  assign f_u_cla12_and78_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and78_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and78_y0 = f_u_cla12_and78_f_u_cla12_pg_logic4_y0 & f_u_cla12_and78_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and79_f_u_cla12_and78_y0 = f_u_cla12_and78_y0;
  assign f_u_cla12_and79_f_u_cla12_and77_y0 = f_u_cla12_and77_y0;
  assign f_u_cla12_and79_y0 = f_u_cla12_and79_f_u_cla12_and78_y0 & f_u_cla12_and79_f_u_cla12_and77_y0;
  assign f_u_cla12_and80_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and80_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and80_y0 = f_u_cla12_and80_f_u_cla12_pg_logic5_y0 & f_u_cla12_and80_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and81_f_u_cla12_and80_y0 = f_u_cla12_and80_y0;
  assign f_u_cla12_and81_f_u_cla12_and79_y0 = f_u_cla12_and79_y0;
  assign f_u_cla12_and81_y0 = f_u_cla12_and81_f_u_cla12_and80_y0 & f_u_cla12_and81_f_u_cla12_and79_y0;
  assign f_u_cla12_and82_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and82_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and82_y0 = f_u_cla12_and82_f_u_cla12_pg_logic3_y0 & f_u_cla12_and82_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and83_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and83_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and83_y0 = f_u_cla12_and83_f_u_cla12_pg_logic4_y0 & f_u_cla12_and83_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and84_f_u_cla12_and83_y0 = f_u_cla12_and83_y0;
  assign f_u_cla12_and84_f_u_cla12_and82_y0 = f_u_cla12_and82_y0;
  assign f_u_cla12_and84_y0 = f_u_cla12_and84_f_u_cla12_and83_y0 & f_u_cla12_and84_f_u_cla12_and82_y0;
  assign f_u_cla12_and85_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and85_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and85_y0 = f_u_cla12_and85_f_u_cla12_pg_logic5_y0 & f_u_cla12_and85_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and86_f_u_cla12_and85_y0 = f_u_cla12_and85_y0;
  assign f_u_cla12_and86_f_u_cla12_and84_y0 = f_u_cla12_and84_y0;
  assign f_u_cla12_and86_y0 = f_u_cla12_and86_f_u_cla12_and85_y0 & f_u_cla12_and86_f_u_cla12_and84_y0;
  assign f_u_cla12_and87_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and87_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and87_y0 = f_u_cla12_and87_f_u_cla12_pg_logic4_y0 & f_u_cla12_and87_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and88_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and88_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and88_y0 = f_u_cla12_and88_f_u_cla12_pg_logic5_y0 & f_u_cla12_and88_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and89_f_u_cla12_and88_y0 = f_u_cla12_and88_y0;
  assign f_u_cla12_and89_f_u_cla12_and87_y0 = f_u_cla12_and87_y0;
  assign f_u_cla12_and89_y0 = f_u_cla12_and89_f_u_cla12_and88_y0 & f_u_cla12_and89_f_u_cla12_and87_y0;
  assign f_u_cla12_and90_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and90_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and90_y0 = f_u_cla12_and90_f_u_cla12_pg_logic5_y0 & f_u_cla12_and90_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_or15_f_u_cla12_and90_y0 = f_u_cla12_and90_y0;
  assign f_u_cla12_or15_f_u_cla12_and65_y0 = f_u_cla12_and65_y0;
  assign f_u_cla12_or15_y0 = f_u_cla12_or15_f_u_cla12_and90_y0 | f_u_cla12_or15_f_u_cla12_and65_y0;
  assign f_u_cla12_or16_f_u_cla12_or15_y0 = f_u_cla12_or15_y0;
  assign f_u_cla12_or16_f_u_cla12_and74_y0 = f_u_cla12_and74_y0;
  assign f_u_cla12_or16_y0 = f_u_cla12_or16_f_u_cla12_or15_y0 | f_u_cla12_or16_f_u_cla12_and74_y0;
  assign f_u_cla12_or17_f_u_cla12_or16_y0 = f_u_cla12_or16_y0;
  assign f_u_cla12_or17_f_u_cla12_and81_y0 = f_u_cla12_and81_y0;
  assign f_u_cla12_or17_y0 = f_u_cla12_or17_f_u_cla12_or16_y0 | f_u_cla12_or17_f_u_cla12_and81_y0;
  assign f_u_cla12_or18_f_u_cla12_or17_y0 = f_u_cla12_or17_y0;
  assign f_u_cla12_or18_f_u_cla12_and86_y0 = f_u_cla12_and86_y0;
  assign f_u_cla12_or18_y0 = f_u_cla12_or18_f_u_cla12_or17_y0 | f_u_cla12_or18_f_u_cla12_and86_y0;
  assign f_u_cla12_or19_f_u_cla12_or18_y0 = f_u_cla12_or18_y0;
  assign f_u_cla12_or19_f_u_cla12_and89_y0 = f_u_cla12_and89_y0;
  assign f_u_cla12_or19_y0 = f_u_cla12_or19_f_u_cla12_or18_y0 | f_u_cla12_or19_f_u_cla12_and89_y0;
  assign f_u_cla12_or20_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_or20_f_u_cla12_or19_y0 = f_u_cla12_or19_y0;
  assign f_u_cla12_or20_y0 = f_u_cla12_or20_f_u_cla12_pg_logic5_y1 | f_u_cla12_or20_f_u_cla12_or19_y0;
  assign f_u_cla12_pg_logic6_a_6 = a_6;
  assign f_u_cla12_pg_logic6_b_6 = b_6;
  assign f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_a_6 | f_u_cla12_pg_logic6_b_6;
  assign f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_a_6 & f_u_cla12_pg_logic6_b_6;
  assign f_u_cla12_pg_logic6_y2 = f_u_cla12_pg_logic6_a_6 ^ f_u_cla12_pg_logic6_b_6;
  assign f_u_cla12_xor6_f_u_cla12_pg_logic6_y2 = f_u_cla12_pg_logic6_y2;
  assign f_u_cla12_xor6_f_u_cla12_or20_y0 = f_u_cla12_or20_y0;
  assign f_u_cla12_xor6_y0 = f_u_cla12_xor6_f_u_cla12_pg_logic6_y2 ^ f_u_cla12_xor6_f_u_cla12_or20_y0;
  assign f_u_cla12_and91_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and91_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and91_y0 = f_u_cla12_and91_f_u_cla12_pg_logic0_y0 & f_u_cla12_and91_constant_wire_0;
  assign f_u_cla12_and92_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and92_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and92_y0 = f_u_cla12_and92_f_u_cla12_pg_logic1_y0 & f_u_cla12_and92_constant_wire_0;
  assign f_u_cla12_and93_f_u_cla12_and92_y0 = f_u_cla12_and92_y0;
  assign f_u_cla12_and93_f_u_cla12_and91_y0 = f_u_cla12_and91_y0;
  assign f_u_cla12_and93_y0 = f_u_cla12_and93_f_u_cla12_and92_y0 & f_u_cla12_and93_f_u_cla12_and91_y0;
  assign f_u_cla12_and94_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and94_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and94_y0 = f_u_cla12_and94_f_u_cla12_pg_logic2_y0 & f_u_cla12_and94_constant_wire_0;
  assign f_u_cla12_and95_f_u_cla12_and94_y0 = f_u_cla12_and94_y0;
  assign f_u_cla12_and95_f_u_cla12_and93_y0 = f_u_cla12_and93_y0;
  assign f_u_cla12_and95_y0 = f_u_cla12_and95_f_u_cla12_and94_y0 & f_u_cla12_and95_f_u_cla12_and93_y0;
  assign f_u_cla12_and96_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and96_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and96_y0 = f_u_cla12_and96_f_u_cla12_pg_logic3_y0 & f_u_cla12_and96_constant_wire_0;
  assign f_u_cla12_and97_f_u_cla12_and96_y0 = f_u_cla12_and96_y0;
  assign f_u_cla12_and97_f_u_cla12_and95_y0 = f_u_cla12_and95_y0;
  assign f_u_cla12_and97_y0 = f_u_cla12_and97_f_u_cla12_and96_y0 & f_u_cla12_and97_f_u_cla12_and95_y0;
  assign f_u_cla12_and98_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and98_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and98_y0 = f_u_cla12_and98_f_u_cla12_pg_logic4_y0 & f_u_cla12_and98_constant_wire_0;
  assign f_u_cla12_and99_f_u_cla12_and98_y0 = f_u_cla12_and98_y0;
  assign f_u_cla12_and99_f_u_cla12_and97_y0 = f_u_cla12_and97_y0;
  assign f_u_cla12_and99_y0 = f_u_cla12_and99_f_u_cla12_and98_y0 & f_u_cla12_and99_f_u_cla12_and97_y0;
  assign f_u_cla12_and100_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and100_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and100_y0 = f_u_cla12_and100_f_u_cla12_pg_logic5_y0 & f_u_cla12_and100_constant_wire_0;
  assign f_u_cla12_and101_f_u_cla12_and100_y0 = f_u_cla12_and100_y0;
  assign f_u_cla12_and101_f_u_cla12_and99_y0 = f_u_cla12_and99_y0;
  assign f_u_cla12_and101_y0 = f_u_cla12_and101_f_u_cla12_and100_y0 & f_u_cla12_and101_f_u_cla12_and99_y0;
  assign f_u_cla12_and102_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and102_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and102_y0 = f_u_cla12_and102_f_u_cla12_pg_logic6_y0 & f_u_cla12_and102_constant_wire_0;
  assign f_u_cla12_and103_f_u_cla12_and102_y0 = f_u_cla12_and102_y0;
  assign f_u_cla12_and103_f_u_cla12_and101_y0 = f_u_cla12_and101_y0;
  assign f_u_cla12_and103_y0 = f_u_cla12_and103_f_u_cla12_and102_y0 & f_u_cla12_and103_f_u_cla12_and101_y0;
  assign f_u_cla12_and104_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and104_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and104_y0 = f_u_cla12_and104_f_u_cla12_pg_logic1_y0 & f_u_cla12_and104_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and105_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and105_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and105_y0 = f_u_cla12_and105_f_u_cla12_pg_logic2_y0 & f_u_cla12_and105_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and106_f_u_cla12_and105_y0 = f_u_cla12_and105_y0;
  assign f_u_cla12_and106_f_u_cla12_and104_y0 = f_u_cla12_and104_y0;
  assign f_u_cla12_and106_y0 = f_u_cla12_and106_f_u_cla12_and105_y0 & f_u_cla12_and106_f_u_cla12_and104_y0;
  assign f_u_cla12_and107_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and107_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and107_y0 = f_u_cla12_and107_f_u_cla12_pg_logic3_y0 & f_u_cla12_and107_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and108_f_u_cla12_and107_y0 = f_u_cla12_and107_y0;
  assign f_u_cla12_and108_f_u_cla12_and106_y0 = f_u_cla12_and106_y0;
  assign f_u_cla12_and108_y0 = f_u_cla12_and108_f_u_cla12_and107_y0 & f_u_cla12_and108_f_u_cla12_and106_y0;
  assign f_u_cla12_and109_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and109_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and109_y0 = f_u_cla12_and109_f_u_cla12_pg_logic4_y0 & f_u_cla12_and109_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and110_f_u_cla12_and109_y0 = f_u_cla12_and109_y0;
  assign f_u_cla12_and110_f_u_cla12_and108_y0 = f_u_cla12_and108_y0;
  assign f_u_cla12_and110_y0 = f_u_cla12_and110_f_u_cla12_and109_y0 & f_u_cla12_and110_f_u_cla12_and108_y0;
  assign f_u_cla12_and111_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and111_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and111_y0 = f_u_cla12_and111_f_u_cla12_pg_logic5_y0 & f_u_cla12_and111_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and112_f_u_cla12_and111_y0 = f_u_cla12_and111_y0;
  assign f_u_cla12_and112_f_u_cla12_and110_y0 = f_u_cla12_and110_y0;
  assign f_u_cla12_and112_y0 = f_u_cla12_and112_f_u_cla12_and111_y0 & f_u_cla12_and112_f_u_cla12_and110_y0;
  assign f_u_cla12_and113_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and113_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and113_y0 = f_u_cla12_and113_f_u_cla12_pg_logic6_y0 & f_u_cla12_and113_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and114_f_u_cla12_and113_y0 = f_u_cla12_and113_y0;
  assign f_u_cla12_and114_f_u_cla12_and112_y0 = f_u_cla12_and112_y0;
  assign f_u_cla12_and114_y0 = f_u_cla12_and114_f_u_cla12_and113_y0 & f_u_cla12_and114_f_u_cla12_and112_y0;
  assign f_u_cla12_and115_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and115_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and115_y0 = f_u_cla12_and115_f_u_cla12_pg_logic2_y0 & f_u_cla12_and115_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and116_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and116_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and116_y0 = f_u_cla12_and116_f_u_cla12_pg_logic3_y0 & f_u_cla12_and116_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and117_f_u_cla12_and116_y0 = f_u_cla12_and116_y0;
  assign f_u_cla12_and117_f_u_cla12_and115_y0 = f_u_cla12_and115_y0;
  assign f_u_cla12_and117_y0 = f_u_cla12_and117_f_u_cla12_and116_y0 & f_u_cla12_and117_f_u_cla12_and115_y0;
  assign f_u_cla12_and118_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and118_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and118_y0 = f_u_cla12_and118_f_u_cla12_pg_logic4_y0 & f_u_cla12_and118_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and119_f_u_cla12_and118_y0 = f_u_cla12_and118_y0;
  assign f_u_cla12_and119_f_u_cla12_and117_y0 = f_u_cla12_and117_y0;
  assign f_u_cla12_and119_y0 = f_u_cla12_and119_f_u_cla12_and118_y0 & f_u_cla12_and119_f_u_cla12_and117_y0;
  assign f_u_cla12_and120_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and120_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and120_y0 = f_u_cla12_and120_f_u_cla12_pg_logic5_y0 & f_u_cla12_and120_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and121_f_u_cla12_and120_y0 = f_u_cla12_and120_y0;
  assign f_u_cla12_and121_f_u_cla12_and119_y0 = f_u_cla12_and119_y0;
  assign f_u_cla12_and121_y0 = f_u_cla12_and121_f_u_cla12_and120_y0 & f_u_cla12_and121_f_u_cla12_and119_y0;
  assign f_u_cla12_and122_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and122_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and122_y0 = f_u_cla12_and122_f_u_cla12_pg_logic6_y0 & f_u_cla12_and122_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and123_f_u_cla12_and122_y0 = f_u_cla12_and122_y0;
  assign f_u_cla12_and123_f_u_cla12_and121_y0 = f_u_cla12_and121_y0;
  assign f_u_cla12_and123_y0 = f_u_cla12_and123_f_u_cla12_and122_y0 & f_u_cla12_and123_f_u_cla12_and121_y0;
  assign f_u_cla12_and124_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and124_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and124_y0 = f_u_cla12_and124_f_u_cla12_pg_logic3_y0 & f_u_cla12_and124_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and125_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and125_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and125_y0 = f_u_cla12_and125_f_u_cla12_pg_logic4_y0 & f_u_cla12_and125_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and126_f_u_cla12_and125_y0 = f_u_cla12_and125_y0;
  assign f_u_cla12_and126_f_u_cla12_and124_y0 = f_u_cla12_and124_y0;
  assign f_u_cla12_and126_y0 = f_u_cla12_and126_f_u_cla12_and125_y0 & f_u_cla12_and126_f_u_cla12_and124_y0;
  assign f_u_cla12_and127_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and127_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and127_y0 = f_u_cla12_and127_f_u_cla12_pg_logic5_y0 & f_u_cla12_and127_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and128_f_u_cla12_and127_y0 = f_u_cla12_and127_y0;
  assign f_u_cla12_and128_f_u_cla12_and126_y0 = f_u_cla12_and126_y0;
  assign f_u_cla12_and128_y0 = f_u_cla12_and128_f_u_cla12_and127_y0 & f_u_cla12_and128_f_u_cla12_and126_y0;
  assign f_u_cla12_and129_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and129_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and129_y0 = f_u_cla12_and129_f_u_cla12_pg_logic6_y0 & f_u_cla12_and129_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and130_f_u_cla12_and129_y0 = f_u_cla12_and129_y0;
  assign f_u_cla12_and130_f_u_cla12_and128_y0 = f_u_cla12_and128_y0;
  assign f_u_cla12_and130_y0 = f_u_cla12_and130_f_u_cla12_and129_y0 & f_u_cla12_and130_f_u_cla12_and128_y0;
  assign f_u_cla12_and131_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and131_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and131_y0 = f_u_cla12_and131_f_u_cla12_pg_logic4_y0 & f_u_cla12_and131_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and132_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and132_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and132_y0 = f_u_cla12_and132_f_u_cla12_pg_logic5_y0 & f_u_cla12_and132_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and133_f_u_cla12_and132_y0 = f_u_cla12_and132_y0;
  assign f_u_cla12_and133_f_u_cla12_and131_y0 = f_u_cla12_and131_y0;
  assign f_u_cla12_and133_y0 = f_u_cla12_and133_f_u_cla12_and132_y0 & f_u_cla12_and133_f_u_cla12_and131_y0;
  assign f_u_cla12_and134_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and134_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and134_y0 = f_u_cla12_and134_f_u_cla12_pg_logic6_y0 & f_u_cla12_and134_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and135_f_u_cla12_and134_y0 = f_u_cla12_and134_y0;
  assign f_u_cla12_and135_f_u_cla12_and133_y0 = f_u_cla12_and133_y0;
  assign f_u_cla12_and135_y0 = f_u_cla12_and135_f_u_cla12_and134_y0 & f_u_cla12_and135_f_u_cla12_and133_y0;
  assign f_u_cla12_and136_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and136_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and136_y0 = f_u_cla12_and136_f_u_cla12_pg_logic5_y0 & f_u_cla12_and136_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and137_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and137_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and137_y0 = f_u_cla12_and137_f_u_cla12_pg_logic6_y0 & f_u_cla12_and137_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and138_f_u_cla12_and137_y0 = f_u_cla12_and137_y0;
  assign f_u_cla12_and138_f_u_cla12_and136_y0 = f_u_cla12_and136_y0;
  assign f_u_cla12_and138_y0 = f_u_cla12_and138_f_u_cla12_and137_y0 & f_u_cla12_and138_f_u_cla12_and136_y0;
  assign f_u_cla12_and139_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and139_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and139_y0 = f_u_cla12_and139_f_u_cla12_pg_logic6_y0 & f_u_cla12_and139_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_or21_f_u_cla12_and139_y0 = f_u_cla12_and139_y0;
  assign f_u_cla12_or21_f_u_cla12_and103_y0 = f_u_cla12_and103_y0;
  assign f_u_cla12_or21_y0 = f_u_cla12_or21_f_u_cla12_and139_y0 | f_u_cla12_or21_f_u_cla12_and103_y0;
  assign f_u_cla12_or22_f_u_cla12_or21_y0 = f_u_cla12_or21_y0;
  assign f_u_cla12_or22_f_u_cla12_and114_y0 = f_u_cla12_and114_y0;
  assign f_u_cla12_or22_y0 = f_u_cla12_or22_f_u_cla12_or21_y0 | f_u_cla12_or22_f_u_cla12_and114_y0;
  assign f_u_cla12_or23_f_u_cla12_or22_y0 = f_u_cla12_or22_y0;
  assign f_u_cla12_or23_f_u_cla12_and123_y0 = f_u_cla12_and123_y0;
  assign f_u_cla12_or23_y0 = f_u_cla12_or23_f_u_cla12_or22_y0 | f_u_cla12_or23_f_u_cla12_and123_y0;
  assign f_u_cla12_or24_f_u_cla12_or23_y0 = f_u_cla12_or23_y0;
  assign f_u_cla12_or24_f_u_cla12_and130_y0 = f_u_cla12_and130_y0;
  assign f_u_cla12_or24_y0 = f_u_cla12_or24_f_u_cla12_or23_y0 | f_u_cla12_or24_f_u_cla12_and130_y0;
  assign f_u_cla12_or25_f_u_cla12_or24_y0 = f_u_cla12_or24_y0;
  assign f_u_cla12_or25_f_u_cla12_and135_y0 = f_u_cla12_and135_y0;
  assign f_u_cla12_or25_y0 = f_u_cla12_or25_f_u_cla12_or24_y0 | f_u_cla12_or25_f_u_cla12_and135_y0;
  assign f_u_cla12_or26_f_u_cla12_or25_y0 = f_u_cla12_or25_y0;
  assign f_u_cla12_or26_f_u_cla12_and138_y0 = f_u_cla12_and138_y0;
  assign f_u_cla12_or26_y0 = f_u_cla12_or26_f_u_cla12_or25_y0 | f_u_cla12_or26_f_u_cla12_and138_y0;
  assign f_u_cla12_or27_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_or27_f_u_cla12_or26_y0 = f_u_cla12_or26_y0;
  assign f_u_cla12_or27_y0 = f_u_cla12_or27_f_u_cla12_pg_logic6_y1 | f_u_cla12_or27_f_u_cla12_or26_y0;
  assign f_u_cla12_pg_logic7_a_7 = a_7;
  assign f_u_cla12_pg_logic7_b_7 = b_7;
  assign f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_a_7 | f_u_cla12_pg_logic7_b_7;
  assign f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_a_7 & f_u_cla12_pg_logic7_b_7;
  assign f_u_cla12_pg_logic7_y2 = f_u_cla12_pg_logic7_a_7 ^ f_u_cla12_pg_logic7_b_7;
  assign f_u_cla12_xor7_f_u_cla12_pg_logic7_y2 = f_u_cla12_pg_logic7_y2;
  assign f_u_cla12_xor7_f_u_cla12_or27_y0 = f_u_cla12_or27_y0;
  assign f_u_cla12_xor7_y0 = f_u_cla12_xor7_f_u_cla12_pg_logic7_y2 ^ f_u_cla12_xor7_f_u_cla12_or27_y0;
  assign f_u_cla12_and140_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and140_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and140_y0 = f_u_cla12_and140_f_u_cla12_pg_logic0_y0 & f_u_cla12_and140_constant_wire_0;
  assign f_u_cla12_and141_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and141_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and141_y0 = f_u_cla12_and141_f_u_cla12_pg_logic1_y0 & f_u_cla12_and141_constant_wire_0;
  assign f_u_cla12_and142_f_u_cla12_and141_y0 = f_u_cla12_and141_y0;
  assign f_u_cla12_and142_f_u_cla12_and140_y0 = f_u_cla12_and140_y0;
  assign f_u_cla12_and142_y0 = f_u_cla12_and142_f_u_cla12_and141_y0 & f_u_cla12_and142_f_u_cla12_and140_y0;
  assign f_u_cla12_and143_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and143_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and143_y0 = f_u_cla12_and143_f_u_cla12_pg_logic2_y0 & f_u_cla12_and143_constant_wire_0;
  assign f_u_cla12_and144_f_u_cla12_and143_y0 = f_u_cla12_and143_y0;
  assign f_u_cla12_and144_f_u_cla12_and142_y0 = f_u_cla12_and142_y0;
  assign f_u_cla12_and144_y0 = f_u_cla12_and144_f_u_cla12_and143_y0 & f_u_cla12_and144_f_u_cla12_and142_y0;
  assign f_u_cla12_and145_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and145_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and145_y0 = f_u_cla12_and145_f_u_cla12_pg_logic3_y0 & f_u_cla12_and145_constant_wire_0;
  assign f_u_cla12_and146_f_u_cla12_and145_y0 = f_u_cla12_and145_y0;
  assign f_u_cla12_and146_f_u_cla12_and144_y0 = f_u_cla12_and144_y0;
  assign f_u_cla12_and146_y0 = f_u_cla12_and146_f_u_cla12_and145_y0 & f_u_cla12_and146_f_u_cla12_and144_y0;
  assign f_u_cla12_and147_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and147_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and147_y0 = f_u_cla12_and147_f_u_cla12_pg_logic4_y0 & f_u_cla12_and147_constant_wire_0;
  assign f_u_cla12_and148_f_u_cla12_and147_y0 = f_u_cla12_and147_y0;
  assign f_u_cla12_and148_f_u_cla12_and146_y0 = f_u_cla12_and146_y0;
  assign f_u_cla12_and148_y0 = f_u_cla12_and148_f_u_cla12_and147_y0 & f_u_cla12_and148_f_u_cla12_and146_y0;
  assign f_u_cla12_and149_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and149_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and149_y0 = f_u_cla12_and149_f_u_cla12_pg_logic5_y0 & f_u_cla12_and149_constant_wire_0;
  assign f_u_cla12_and150_f_u_cla12_and149_y0 = f_u_cla12_and149_y0;
  assign f_u_cla12_and150_f_u_cla12_and148_y0 = f_u_cla12_and148_y0;
  assign f_u_cla12_and150_y0 = f_u_cla12_and150_f_u_cla12_and149_y0 & f_u_cla12_and150_f_u_cla12_and148_y0;
  assign f_u_cla12_and151_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and151_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and151_y0 = f_u_cla12_and151_f_u_cla12_pg_logic6_y0 & f_u_cla12_and151_constant_wire_0;
  assign f_u_cla12_and152_f_u_cla12_and151_y0 = f_u_cla12_and151_y0;
  assign f_u_cla12_and152_f_u_cla12_and150_y0 = f_u_cla12_and150_y0;
  assign f_u_cla12_and152_y0 = f_u_cla12_and152_f_u_cla12_and151_y0 & f_u_cla12_and152_f_u_cla12_and150_y0;
  assign f_u_cla12_and153_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and153_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and153_y0 = f_u_cla12_and153_f_u_cla12_pg_logic7_y0 & f_u_cla12_and153_constant_wire_0;
  assign f_u_cla12_and154_f_u_cla12_and153_y0 = f_u_cla12_and153_y0;
  assign f_u_cla12_and154_f_u_cla12_and152_y0 = f_u_cla12_and152_y0;
  assign f_u_cla12_and154_y0 = f_u_cla12_and154_f_u_cla12_and153_y0 & f_u_cla12_and154_f_u_cla12_and152_y0;
  assign f_u_cla12_and155_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and155_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and155_y0 = f_u_cla12_and155_f_u_cla12_pg_logic1_y0 & f_u_cla12_and155_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and156_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and156_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and156_y0 = f_u_cla12_and156_f_u_cla12_pg_logic2_y0 & f_u_cla12_and156_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and157_f_u_cla12_and156_y0 = f_u_cla12_and156_y0;
  assign f_u_cla12_and157_f_u_cla12_and155_y0 = f_u_cla12_and155_y0;
  assign f_u_cla12_and157_y0 = f_u_cla12_and157_f_u_cla12_and156_y0 & f_u_cla12_and157_f_u_cla12_and155_y0;
  assign f_u_cla12_and158_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and158_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and158_y0 = f_u_cla12_and158_f_u_cla12_pg_logic3_y0 & f_u_cla12_and158_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and159_f_u_cla12_and158_y0 = f_u_cla12_and158_y0;
  assign f_u_cla12_and159_f_u_cla12_and157_y0 = f_u_cla12_and157_y0;
  assign f_u_cla12_and159_y0 = f_u_cla12_and159_f_u_cla12_and158_y0 & f_u_cla12_and159_f_u_cla12_and157_y0;
  assign f_u_cla12_and160_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and160_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and160_y0 = f_u_cla12_and160_f_u_cla12_pg_logic4_y0 & f_u_cla12_and160_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and161_f_u_cla12_and160_y0 = f_u_cla12_and160_y0;
  assign f_u_cla12_and161_f_u_cla12_and159_y0 = f_u_cla12_and159_y0;
  assign f_u_cla12_and161_y0 = f_u_cla12_and161_f_u_cla12_and160_y0 & f_u_cla12_and161_f_u_cla12_and159_y0;
  assign f_u_cla12_and162_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and162_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and162_y0 = f_u_cla12_and162_f_u_cla12_pg_logic5_y0 & f_u_cla12_and162_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and163_f_u_cla12_and162_y0 = f_u_cla12_and162_y0;
  assign f_u_cla12_and163_f_u_cla12_and161_y0 = f_u_cla12_and161_y0;
  assign f_u_cla12_and163_y0 = f_u_cla12_and163_f_u_cla12_and162_y0 & f_u_cla12_and163_f_u_cla12_and161_y0;
  assign f_u_cla12_and164_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and164_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and164_y0 = f_u_cla12_and164_f_u_cla12_pg_logic6_y0 & f_u_cla12_and164_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and165_f_u_cla12_and164_y0 = f_u_cla12_and164_y0;
  assign f_u_cla12_and165_f_u_cla12_and163_y0 = f_u_cla12_and163_y0;
  assign f_u_cla12_and165_y0 = f_u_cla12_and165_f_u_cla12_and164_y0 & f_u_cla12_and165_f_u_cla12_and163_y0;
  assign f_u_cla12_and166_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and166_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and166_y0 = f_u_cla12_and166_f_u_cla12_pg_logic7_y0 & f_u_cla12_and166_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and167_f_u_cla12_and166_y0 = f_u_cla12_and166_y0;
  assign f_u_cla12_and167_f_u_cla12_and165_y0 = f_u_cla12_and165_y0;
  assign f_u_cla12_and167_y0 = f_u_cla12_and167_f_u_cla12_and166_y0 & f_u_cla12_and167_f_u_cla12_and165_y0;
  assign f_u_cla12_and168_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and168_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and168_y0 = f_u_cla12_and168_f_u_cla12_pg_logic2_y0 & f_u_cla12_and168_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and169_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and169_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and169_y0 = f_u_cla12_and169_f_u_cla12_pg_logic3_y0 & f_u_cla12_and169_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and170_f_u_cla12_and169_y0 = f_u_cla12_and169_y0;
  assign f_u_cla12_and170_f_u_cla12_and168_y0 = f_u_cla12_and168_y0;
  assign f_u_cla12_and170_y0 = f_u_cla12_and170_f_u_cla12_and169_y0 & f_u_cla12_and170_f_u_cla12_and168_y0;
  assign f_u_cla12_and171_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and171_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and171_y0 = f_u_cla12_and171_f_u_cla12_pg_logic4_y0 & f_u_cla12_and171_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and172_f_u_cla12_and171_y0 = f_u_cla12_and171_y0;
  assign f_u_cla12_and172_f_u_cla12_and170_y0 = f_u_cla12_and170_y0;
  assign f_u_cla12_and172_y0 = f_u_cla12_and172_f_u_cla12_and171_y0 & f_u_cla12_and172_f_u_cla12_and170_y0;
  assign f_u_cla12_and173_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and173_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and173_y0 = f_u_cla12_and173_f_u_cla12_pg_logic5_y0 & f_u_cla12_and173_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and174_f_u_cla12_and173_y0 = f_u_cla12_and173_y0;
  assign f_u_cla12_and174_f_u_cla12_and172_y0 = f_u_cla12_and172_y0;
  assign f_u_cla12_and174_y0 = f_u_cla12_and174_f_u_cla12_and173_y0 & f_u_cla12_and174_f_u_cla12_and172_y0;
  assign f_u_cla12_and175_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and175_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and175_y0 = f_u_cla12_and175_f_u_cla12_pg_logic6_y0 & f_u_cla12_and175_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and176_f_u_cla12_and175_y0 = f_u_cla12_and175_y0;
  assign f_u_cla12_and176_f_u_cla12_and174_y0 = f_u_cla12_and174_y0;
  assign f_u_cla12_and176_y0 = f_u_cla12_and176_f_u_cla12_and175_y0 & f_u_cla12_and176_f_u_cla12_and174_y0;
  assign f_u_cla12_and177_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and177_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and177_y0 = f_u_cla12_and177_f_u_cla12_pg_logic7_y0 & f_u_cla12_and177_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and178_f_u_cla12_and177_y0 = f_u_cla12_and177_y0;
  assign f_u_cla12_and178_f_u_cla12_and176_y0 = f_u_cla12_and176_y0;
  assign f_u_cla12_and178_y0 = f_u_cla12_and178_f_u_cla12_and177_y0 & f_u_cla12_and178_f_u_cla12_and176_y0;
  assign f_u_cla12_and179_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and179_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and179_y0 = f_u_cla12_and179_f_u_cla12_pg_logic3_y0 & f_u_cla12_and179_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and180_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and180_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and180_y0 = f_u_cla12_and180_f_u_cla12_pg_logic4_y0 & f_u_cla12_and180_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and181_f_u_cla12_and180_y0 = f_u_cla12_and180_y0;
  assign f_u_cla12_and181_f_u_cla12_and179_y0 = f_u_cla12_and179_y0;
  assign f_u_cla12_and181_y0 = f_u_cla12_and181_f_u_cla12_and180_y0 & f_u_cla12_and181_f_u_cla12_and179_y0;
  assign f_u_cla12_and182_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and182_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and182_y0 = f_u_cla12_and182_f_u_cla12_pg_logic5_y0 & f_u_cla12_and182_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and183_f_u_cla12_and182_y0 = f_u_cla12_and182_y0;
  assign f_u_cla12_and183_f_u_cla12_and181_y0 = f_u_cla12_and181_y0;
  assign f_u_cla12_and183_y0 = f_u_cla12_and183_f_u_cla12_and182_y0 & f_u_cla12_and183_f_u_cla12_and181_y0;
  assign f_u_cla12_and184_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and184_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and184_y0 = f_u_cla12_and184_f_u_cla12_pg_logic6_y0 & f_u_cla12_and184_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and185_f_u_cla12_and184_y0 = f_u_cla12_and184_y0;
  assign f_u_cla12_and185_f_u_cla12_and183_y0 = f_u_cla12_and183_y0;
  assign f_u_cla12_and185_y0 = f_u_cla12_and185_f_u_cla12_and184_y0 & f_u_cla12_and185_f_u_cla12_and183_y0;
  assign f_u_cla12_and186_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and186_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and186_y0 = f_u_cla12_and186_f_u_cla12_pg_logic7_y0 & f_u_cla12_and186_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and187_f_u_cla12_and186_y0 = f_u_cla12_and186_y0;
  assign f_u_cla12_and187_f_u_cla12_and185_y0 = f_u_cla12_and185_y0;
  assign f_u_cla12_and187_y0 = f_u_cla12_and187_f_u_cla12_and186_y0 & f_u_cla12_and187_f_u_cla12_and185_y0;
  assign f_u_cla12_and188_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and188_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and188_y0 = f_u_cla12_and188_f_u_cla12_pg_logic4_y0 & f_u_cla12_and188_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and189_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and189_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and189_y0 = f_u_cla12_and189_f_u_cla12_pg_logic5_y0 & f_u_cla12_and189_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and190_f_u_cla12_and189_y0 = f_u_cla12_and189_y0;
  assign f_u_cla12_and190_f_u_cla12_and188_y0 = f_u_cla12_and188_y0;
  assign f_u_cla12_and190_y0 = f_u_cla12_and190_f_u_cla12_and189_y0 & f_u_cla12_and190_f_u_cla12_and188_y0;
  assign f_u_cla12_and191_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and191_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and191_y0 = f_u_cla12_and191_f_u_cla12_pg_logic6_y0 & f_u_cla12_and191_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and192_f_u_cla12_and191_y0 = f_u_cla12_and191_y0;
  assign f_u_cla12_and192_f_u_cla12_and190_y0 = f_u_cla12_and190_y0;
  assign f_u_cla12_and192_y0 = f_u_cla12_and192_f_u_cla12_and191_y0 & f_u_cla12_and192_f_u_cla12_and190_y0;
  assign f_u_cla12_and193_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and193_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and193_y0 = f_u_cla12_and193_f_u_cla12_pg_logic7_y0 & f_u_cla12_and193_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and194_f_u_cla12_and193_y0 = f_u_cla12_and193_y0;
  assign f_u_cla12_and194_f_u_cla12_and192_y0 = f_u_cla12_and192_y0;
  assign f_u_cla12_and194_y0 = f_u_cla12_and194_f_u_cla12_and193_y0 & f_u_cla12_and194_f_u_cla12_and192_y0;
  assign f_u_cla12_and195_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and195_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and195_y0 = f_u_cla12_and195_f_u_cla12_pg_logic5_y0 & f_u_cla12_and195_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and196_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and196_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and196_y0 = f_u_cla12_and196_f_u_cla12_pg_logic6_y0 & f_u_cla12_and196_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and197_f_u_cla12_and196_y0 = f_u_cla12_and196_y0;
  assign f_u_cla12_and197_f_u_cla12_and195_y0 = f_u_cla12_and195_y0;
  assign f_u_cla12_and197_y0 = f_u_cla12_and197_f_u_cla12_and196_y0 & f_u_cla12_and197_f_u_cla12_and195_y0;
  assign f_u_cla12_and198_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and198_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and198_y0 = f_u_cla12_and198_f_u_cla12_pg_logic7_y0 & f_u_cla12_and198_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and199_f_u_cla12_and198_y0 = f_u_cla12_and198_y0;
  assign f_u_cla12_and199_f_u_cla12_and197_y0 = f_u_cla12_and197_y0;
  assign f_u_cla12_and199_y0 = f_u_cla12_and199_f_u_cla12_and198_y0 & f_u_cla12_and199_f_u_cla12_and197_y0;
  assign f_u_cla12_and200_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and200_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and200_y0 = f_u_cla12_and200_f_u_cla12_pg_logic6_y0 & f_u_cla12_and200_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and201_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and201_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and201_y0 = f_u_cla12_and201_f_u_cla12_pg_logic7_y0 & f_u_cla12_and201_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and202_f_u_cla12_and201_y0 = f_u_cla12_and201_y0;
  assign f_u_cla12_and202_f_u_cla12_and200_y0 = f_u_cla12_and200_y0;
  assign f_u_cla12_and202_y0 = f_u_cla12_and202_f_u_cla12_and201_y0 & f_u_cla12_and202_f_u_cla12_and200_y0;
  assign f_u_cla12_and203_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and203_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and203_y0 = f_u_cla12_and203_f_u_cla12_pg_logic7_y0 & f_u_cla12_and203_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_or28_f_u_cla12_and203_y0 = f_u_cla12_and203_y0;
  assign f_u_cla12_or28_f_u_cla12_and154_y0 = f_u_cla12_and154_y0;
  assign f_u_cla12_or28_y0 = f_u_cla12_or28_f_u_cla12_and203_y0 | f_u_cla12_or28_f_u_cla12_and154_y0;
  assign f_u_cla12_or29_f_u_cla12_or28_y0 = f_u_cla12_or28_y0;
  assign f_u_cla12_or29_f_u_cla12_and167_y0 = f_u_cla12_and167_y0;
  assign f_u_cla12_or29_y0 = f_u_cla12_or29_f_u_cla12_or28_y0 | f_u_cla12_or29_f_u_cla12_and167_y0;
  assign f_u_cla12_or30_f_u_cla12_or29_y0 = f_u_cla12_or29_y0;
  assign f_u_cla12_or30_f_u_cla12_and178_y0 = f_u_cla12_and178_y0;
  assign f_u_cla12_or30_y0 = f_u_cla12_or30_f_u_cla12_or29_y0 | f_u_cla12_or30_f_u_cla12_and178_y0;
  assign f_u_cla12_or31_f_u_cla12_or30_y0 = f_u_cla12_or30_y0;
  assign f_u_cla12_or31_f_u_cla12_and187_y0 = f_u_cla12_and187_y0;
  assign f_u_cla12_or31_y0 = f_u_cla12_or31_f_u_cla12_or30_y0 | f_u_cla12_or31_f_u_cla12_and187_y0;
  assign f_u_cla12_or32_f_u_cla12_or31_y0 = f_u_cla12_or31_y0;
  assign f_u_cla12_or32_f_u_cla12_and194_y0 = f_u_cla12_and194_y0;
  assign f_u_cla12_or32_y0 = f_u_cla12_or32_f_u_cla12_or31_y0 | f_u_cla12_or32_f_u_cla12_and194_y0;
  assign f_u_cla12_or33_f_u_cla12_or32_y0 = f_u_cla12_or32_y0;
  assign f_u_cla12_or33_f_u_cla12_and199_y0 = f_u_cla12_and199_y0;
  assign f_u_cla12_or33_y0 = f_u_cla12_or33_f_u_cla12_or32_y0 | f_u_cla12_or33_f_u_cla12_and199_y0;
  assign f_u_cla12_or34_f_u_cla12_or33_y0 = f_u_cla12_or33_y0;
  assign f_u_cla12_or34_f_u_cla12_and202_y0 = f_u_cla12_and202_y0;
  assign f_u_cla12_or34_y0 = f_u_cla12_or34_f_u_cla12_or33_y0 | f_u_cla12_or34_f_u_cla12_and202_y0;
  assign f_u_cla12_or35_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_or35_f_u_cla12_or34_y0 = f_u_cla12_or34_y0;
  assign f_u_cla12_or35_y0 = f_u_cla12_or35_f_u_cla12_pg_logic7_y1 | f_u_cla12_or35_f_u_cla12_or34_y0;
  assign f_u_cla12_pg_logic8_a_8 = a_8;
  assign f_u_cla12_pg_logic8_b_8 = b_8;
  assign f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_a_8 | f_u_cla12_pg_logic8_b_8;
  assign f_u_cla12_pg_logic8_y1 = f_u_cla12_pg_logic8_a_8 & f_u_cla12_pg_logic8_b_8;
  assign f_u_cla12_pg_logic8_y2 = f_u_cla12_pg_logic8_a_8 ^ f_u_cla12_pg_logic8_b_8;
  assign f_u_cla12_xor8_f_u_cla12_pg_logic8_y2 = f_u_cla12_pg_logic8_y2;
  assign f_u_cla12_xor8_f_u_cla12_or35_y0 = f_u_cla12_or35_y0;
  assign f_u_cla12_xor8_y0 = f_u_cla12_xor8_f_u_cla12_pg_logic8_y2 ^ f_u_cla12_xor8_f_u_cla12_or35_y0;
  assign f_u_cla12_and204_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and204_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and204_y0 = f_u_cla12_and204_f_u_cla12_pg_logic0_y0 & f_u_cla12_and204_constant_wire_0;
  assign f_u_cla12_and205_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and205_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and205_y0 = f_u_cla12_and205_f_u_cla12_pg_logic1_y0 & f_u_cla12_and205_constant_wire_0;
  assign f_u_cla12_and206_f_u_cla12_and205_y0 = f_u_cla12_and205_y0;
  assign f_u_cla12_and206_f_u_cla12_and204_y0 = f_u_cla12_and204_y0;
  assign f_u_cla12_and206_y0 = f_u_cla12_and206_f_u_cla12_and205_y0 & f_u_cla12_and206_f_u_cla12_and204_y0;
  assign f_u_cla12_and207_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and207_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and207_y0 = f_u_cla12_and207_f_u_cla12_pg_logic2_y0 & f_u_cla12_and207_constant_wire_0;
  assign f_u_cla12_and208_f_u_cla12_and207_y0 = f_u_cla12_and207_y0;
  assign f_u_cla12_and208_f_u_cla12_and206_y0 = f_u_cla12_and206_y0;
  assign f_u_cla12_and208_y0 = f_u_cla12_and208_f_u_cla12_and207_y0 & f_u_cla12_and208_f_u_cla12_and206_y0;
  assign f_u_cla12_and209_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and209_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and209_y0 = f_u_cla12_and209_f_u_cla12_pg_logic3_y0 & f_u_cla12_and209_constant_wire_0;
  assign f_u_cla12_and210_f_u_cla12_and209_y0 = f_u_cla12_and209_y0;
  assign f_u_cla12_and210_f_u_cla12_and208_y0 = f_u_cla12_and208_y0;
  assign f_u_cla12_and210_y0 = f_u_cla12_and210_f_u_cla12_and209_y0 & f_u_cla12_and210_f_u_cla12_and208_y0;
  assign f_u_cla12_and211_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and211_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and211_y0 = f_u_cla12_and211_f_u_cla12_pg_logic4_y0 & f_u_cla12_and211_constant_wire_0;
  assign f_u_cla12_and212_f_u_cla12_and211_y0 = f_u_cla12_and211_y0;
  assign f_u_cla12_and212_f_u_cla12_and210_y0 = f_u_cla12_and210_y0;
  assign f_u_cla12_and212_y0 = f_u_cla12_and212_f_u_cla12_and211_y0 & f_u_cla12_and212_f_u_cla12_and210_y0;
  assign f_u_cla12_and213_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and213_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and213_y0 = f_u_cla12_and213_f_u_cla12_pg_logic5_y0 & f_u_cla12_and213_constant_wire_0;
  assign f_u_cla12_and214_f_u_cla12_and213_y0 = f_u_cla12_and213_y0;
  assign f_u_cla12_and214_f_u_cla12_and212_y0 = f_u_cla12_and212_y0;
  assign f_u_cla12_and214_y0 = f_u_cla12_and214_f_u_cla12_and213_y0 & f_u_cla12_and214_f_u_cla12_and212_y0;
  assign f_u_cla12_and215_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and215_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and215_y0 = f_u_cla12_and215_f_u_cla12_pg_logic6_y0 & f_u_cla12_and215_constant_wire_0;
  assign f_u_cla12_and216_f_u_cla12_and215_y0 = f_u_cla12_and215_y0;
  assign f_u_cla12_and216_f_u_cla12_and214_y0 = f_u_cla12_and214_y0;
  assign f_u_cla12_and216_y0 = f_u_cla12_and216_f_u_cla12_and215_y0 & f_u_cla12_and216_f_u_cla12_and214_y0;
  assign f_u_cla12_and217_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and217_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and217_y0 = f_u_cla12_and217_f_u_cla12_pg_logic7_y0 & f_u_cla12_and217_constant_wire_0;
  assign f_u_cla12_and218_f_u_cla12_and217_y0 = f_u_cla12_and217_y0;
  assign f_u_cla12_and218_f_u_cla12_and216_y0 = f_u_cla12_and216_y0;
  assign f_u_cla12_and218_y0 = f_u_cla12_and218_f_u_cla12_and217_y0 & f_u_cla12_and218_f_u_cla12_and216_y0;
  assign f_u_cla12_and219_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and219_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and219_y0 = f_u_cla12_and219_f_u_cla12_pg_logic8_y0 & f_u_cla12_and219_constant_wire_0;
  assign f_u_cla12_and220_f_u_cla12_and219_y0 = f_u_cla12_and219_y0;
  assign f_u_cla12_and220_f_u_cla12_and218_y0 = f_u_cla12_and218_y0;
  assign f_u_cla12_and220_y0 = f_u_cla12_and220_f_u_cla12_and219_y0 & f_u_cla12_and220_f_u_cla12_and218_y0;
  assign f_u_cla12_and221_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and221_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and221_y0 = f_u_cla12_and221_f_u_cla12_pg_logic1_y0 & f_u_cla12_and221_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and222_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and222_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and222_y0 = f_u_cla12_and222_f_u_cla12_pg_logic2_y0 & f_u_cla12_and222_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and223_f_u_cla12_and222_y0 = f_u_cla12_and222_y0;
  assign f_u_cla12_and223_f_u_cla12_and221_y0 = f_u_cla12_and221_y0;
  assign f_u_cla12_and223_y0 = f_u_cla12_and223_f_u_cla12_and222_y0 & f_u_cla12_and223_f_u_cla12_and221_y0;
  assign f_u_cla12_and224_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and224_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and224_y0 = f_u_cla12_and224_f_u_cla12_pg_logic3_y0 & f_u_cla12_and224_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and225_f_u_cla12_and224_y0 = f_u_cla12_and224_y0;
  assign f_u_cla12_and225_f_u_cla12_and223_y0 = f_u_cla12_and223_y0;
  assign f_u_cla12_and225_y0 = f_u_cla12_and225_f_u_cla12_and224_y0 & f_u_cla12_and225_f_u_cla12_and223_y0;
  assign f_u_cla12_and226_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and226_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and226_y0 = f_u_cla12_and226_f_u_cla12_pg_logic4_y0 & f_u_cla12_and226_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and227_f_u_cla12_and226_y0 = f_u_cla12_and226_y0;
  assign f_u_cla12_and227_f_u_cla12_and225_y0 = f_u_cla12_and225_y0;
  assign f_u_cla12_and227_y0 = f_u_cla12_and227_f_u_cla12_and226_y0 & f_u_cla12_and227_f_u_cla12_and225_y0;
  assign f_u_cla12_and228_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and228_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and228_y0 = f_u_cla12_and228_f_u_cla12_pg_logic5_y0 & f_u_cla12_and228_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and229_f_u_cla12_and228_y0 = f_u_cla12_and228_y0;
  assign f_u_cla12_and229_f_u_cla12_and227_y0 = f_u_cla12_and227_y0;
  assign f_u_cla12_and229_y0 = f_u_cla12_and229_f_u_cla12_and228_y0 & f_u_cla12_and229_f_u_cla12_and227_y0;
  assign f_u_cla12_and230_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and230_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and230_y0 = f_u_cla12_and230_f_u_cla12_pg_logic6_y0 & f_u_cla12_and230_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and231_f_u_cla12_and230_y0 = f_u_cla12_and230_y0;
  assign f_u_cla12_and231_f_u_cla12_and229_y0 = f_u_cla12_and229_y0;
  assign f_u_cla12_and231_y0 = f_u_cla12_and231_f_u_cla12_and230_y0 & f_u_cla12_and231_f_u_cla12_and229_y0;
  assign f_u_cla12_and232_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and232_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and232_y0 = f_u_cla12_and232_f_u_cla12_pg_logic7_y0 & f_u_cla12_and232_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and233_f_u_cla12_and232_y0 = f_u_cla12_and232_y0;
  assign f_u_cla12_and233_f_u_cla12_and231_y0 = f_u_cla12_and231_y0;
  assign f_u_cla12_and233_y0 = f_u_cla12_and233_f_u_cla12_and232_y0 & f_u_cla12_and233_f_u_cla12_and231_y0;
  assign f_u_cla12_and234_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and234_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and234_y0 = f_u_cla12_and234_f_u_cla12_pg_logic8_y0 & f_u_cla12_and234_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and235_f_u_cla12_and234_y0 = f_u_cla12_and234_y0;
  assign f_u_cla12_and235_f_u_cla12_and233_y0 = f_u_cla12_and233_y0;
  assign f_u_cla12_and235_y0 = f_u_cla12_and235_f_u_cla12_and234_y0 & f_u_cla12_and235_f_u_cla12_and233_y0;
  assign f_u_cla12_and236_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and236_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and236_y0 = f_u_cla12_and236_f_u_cla12_pg_logic2_y0 & f_u_cla12_and236_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and237_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and237_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and237_y0 = f_u_cla12_and237_f_u_cla12_pg_logic3_y0 & f_u_cla12_and237_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and238_f_u_cla12_and237_y0 = f_u_cla12_and237_y0;
  assign f_u_cla12_and238_f_u_cla12_and236_y0 = f_u_cla12_and236_y0;
  assign f_u_cla12_and238_y0 = f_u_cla12_and238_f_u_cla12_and237_y0 & f_u_cla12_and238_f_u_cla12_and236_y0;
  assign f_u_cla12_and239_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and239_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and239_y0 = f_u_cla12_and239_f_u_cla12_pg_logic4_y0 & f_u_cla12_and239_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and240_f_u_cla12_and239_y0 = f_u_cla12_and239_y0;
  assign f_u_cla12_and240_f_u_cla12_and238_y0 = f_u_cla12_and238_y0;
  assign f_u_cla12_and240_y0 = f_u_cla12_and240_f_u_cla12_and239_y0 & f_u_cla12_and240_f_u_cla12_and238_y0;
  assign f_u_cla12_and241_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and241_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and241_y0 = f_u_cla12_and241_f_u_cla12_pg_logic5_y0 & f_u_cla12_and241_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and242_f_u_cla12_and241_y0 = f_u_cla12_and241_y0;
  assign f_u_cla12_and242_f_u_cla12_and240_y0 = f_u_cla12_and240_y0;
  assign f_u_cla12_and242_y0 = f_u_cla12_and242_f_u_cla12_and241_y0 & f_u_cla12_and242_f_u_cla12_and240_y0;
  assign f_u_cla12_and243_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and243_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and243_y0 = f_u_cla12_and243_f_u_cla12_pg_logic6_y0 & f_u_cla12_and243_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and244_f_u_cla12_and243_y0 = f_u_cla12_and243_y0;
  assign f_u_cla12_and244_f_u_cla12_and242_y0 = f_u_cla12_and242_y0;
  assign f_u_cla12_and244_y0 = f_u_cla12_and244_f_u_cla12_and243_y0 & f_u_cla12_and244_f_u_cla12_and242_y0;
  assign f_u_cla12_and245_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and245_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and245_y0 = f_u_cla12_and245_f_u_cla12_pg_logic7_y0 & f_u_cla12_and245_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and246_f_u_cla12_and245_y0 = f_u_cla12_and245_y0;
  assign f_u_cla12_and246_f_u_cla12_and244_y0 = f_u_cla12_and244_y0;
  assign f_u_cla12_and246_y0 = f_u_cla12_and246_f_u_cla12_and245_y0 & f_u_cla12_and246_f_u_cla12_and244_y0;
  assign f_u_cla12_and247_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and247_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and247_y0 = f_u_cla12_and247_f_u_cla12_pg_logic8_y0 & f_u_cla12_and247_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and248_f_u_cla12_and247_y0 = f_u_cla12_and247_y0;
  assign f_u_cla12_and248_f_u_cla12_and246_y0 = f_u_cla12_and246_y0;
  assign f_u_cla12_and248_y0 = f_u_cla12_and248_f_u_cla12_and247_y0 & f_u_cla12_and248_f_u_cla12_and246_y0;
  assign f_u_cla12_and249_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and249_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and249_y0 = f_u_cla12_and249_f_u_cla12_pg_logic3_y0 & f_u_cla12_and249_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and250_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and250_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and250_y0 = f_u_cla12_and250_f_u_cla12_pg_logic4_y0 & f_u_cla12_and250_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and251_f_u_cla12_and250_y0 = f_u_cla12_and250_y0;
  assign f_u_cla12_and251_f_u_cla12_and249_y0 = f_u_cla12_and249_y0;
  assign f_u_cla12_and251_y0 = f_u_cla12_and251_f_u_cla12_and250_y0 & f_u_cla12_and251_f_u_cla12_and249_y0;
  assign f_u_cla12_and252_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and252_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and252_y0 = f_u_cla12_and252_f_u_cla12_pg_logic5_y0 & f_u_cla12_and252_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and253_f_u_cla12_and252_y0 = f_u_cla12_and252_y0;
  assign f_u_cla12_and253_f_u_cla12_and251_y0 = f_u_cla12_and251_y0;
  assign f_u_cla12_and253_y0 = f_u_cla12_and253_f_u_cla12_and252_y0 & f_u_cla12_and253_f_u_cla12_and251_y0;
  assign f_u_cla12_and254_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and254_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and254_y0 = f_u_cla12_and254_f_u_cla12_pg_logic6_y0 & f_u_cla12_and254_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and255_f_u_cla12_and254_y0 = f_u_cla12_and254_y0;
  assign f_u_cla12_and255_f_u_cla12_and253_y0 = f_u_cla12_and253_y0;
  assign f_u_cla12_and255_y0 = f_u_cla12_and255_f_u_cla12_and254_y0 & f_u_cla12_and255_f_u_cla12_and253_y0;
  assign f_u_cla12_and256_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and256_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and256_y0 = f_u_cla12_and256_f_u_cla12_pg_logic7_y0 & f_u_cla12_and256_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and257_f_u_cla12_and256_y0 = f_u_cla12_and256_y0;
  assign f_u_cla12_and257_f_u_cla12_and255_y0 = f_u_cla12_and255_y0;
  assign f_u_cla12_and257_y0 = f_u_cla12_and257_f_u_cla12_and256_y0 & f_u_cla12_and257_f_u_cla12_and255_y0;
  assign f_u_cla12_and258_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and258_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and258_y0 = f_u_cla12_and258_f_u_cla12_pg_logic8_y0 & f_u_cla12_and258_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and259_f_u_cla12_and258_y0 = f_u_cla12_and258_y0;
  assign f_u_cla12_and259_f_u_cla12_and257_y0 = f_u_cla12_and257_y0;
  assign f_u_cla12_and259_y0 = f_u_cla12_and259_f_u_cla12_and258_y0 & f_u_cla12_and259_f_u_cla12_and257_y0;
  assign f_u_cla12_and260_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and260_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and260_y0 = f_u_cla12_and260_f_u_cla12_pg_logic4_y0 & f_u_cla12_and260_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and261_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and261_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and261_y0 = f_u_cla12_and261_f_u_cla12_pg_logic5_y0 & f_u_cla12_and261_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and262_f_u_cla12_and261_y0 = f_u_cla12_and261_y0;
  assign f_u_cla12_and262_f_u_cla12_and260_y0 = f_u_cla12_and260_y0;
  assign f_u_cla12_and262_y0 = f_u_cla12_and262_f_u_cla12_and261_y0 & f_u_cla12_and262_f_u_cla12_and260_y0;
  assign f_u_cla12_and263_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and263_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and263_y0 = f_u_cla12_and263_f_u_cla12_pg_logic6_y0 & f_u_cla12_and263_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and264_f_u_cla12_and263_y0 = f_u_cla12_and263_y0;
  assign f_u_cla12_and264_f_u_cla12_and262_y0 = f_u_cla12_and262_y0;
  assign f_u_cla12_and264_y0 = f_u_cla12_and264_f_u_cla12_and263_y0 & f_u_cla12_and264_f_u_cla12_and262_y0;
  assign f_u_cla12_and265_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and265_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and265_y0 = f_u_cla12_and265_f_u_cla12_pg_logic7_y0 & f_u_cla12_and265_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and266_f_u_cla12_and265_y0 = f_u_cla12_and265_y0;
  assign f_u_cla12_and266_f_u_cla12_and264_y0 = f_u_cla12_and264_y0;
  assign f_u_cla12_and266_y0 = f_u_cla12_and266_f_u_cla12_and265_y0 & f_u_cla12_and266_f_u_cla12_and264_y0;
  assign f_u_cla12_and267_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and267_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and267_y0 = f_u_cla12_and267_f_u_cla12_pg_logic8_y0 & f_u_cla12_and267_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and268_f_u_cla12_and267_y0 = f_u_cla12_and267_y0;
  assign f_u_cla12_and268_f_u_cla12_and266_y0 = f_u_cla12_and266_y0;
  assign f_u_cla12_and268_y0 = f_u_cla12_and268_f_u_cla12_and267_y0 & f_u_cla12_and268_f_u_cla12_and266_y0;
  assign f_u_cla12_and269_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and269_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and269_y0 = f_u_cla12_and269_f_u_cla12_pg_logic5_y0 & f_u_cla12_and269_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and270_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and270_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and270_y0 = f_u_cla12_and270_f_u_cla12_pg_logic6_y0 & f_u_cla12_and270_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and271_f_u_cla12_and270_y0 = f_u_cla12_and270_y0;
  assign f_u_cla12_and271_f_u_cla12_and269_y0 = f_u_cla12_and269_y0;
  assign f_u_cla12_and271_y0 = f_u_cla12_and271_f_u_cla12_and270_y0 & f_u_cla12_and271_f_u_cla12_and269_y0;
  assign f_u_cla12_and272_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and272_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and272_y0 = f_u_cla12_and272_f_u_cla12_pg_logic7_y0 & f_u_cla12_and272_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and273_f_u_cla12_and272_y0 = f_u_cla12_and272_y0;
  assign f_u_cla12_and273_f_u_cla12_and271_y0 = f_u_cla12_and271_y0;
  assign f_u_cla12_and273_y0 = f_u_cla12_and273_f_u_cla12_and272_y0 & f_u_cla12_and273_f_u_cla12_and271_y0;
  assign f_u_cla12_and274_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and274_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and274_y0 = f_u_cla12_and274_f_u_cla12_pg_logic8_y0 & f_u_cla12_and274_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and275_f_u_cla12_and274_y0 = f_u_cla12_and274_y0;
  assign f_u_cla12_and275_f_u_cla12_and273_y0 = f_u_cla12_and273_y0;
  assign f_u_cla12_and275_y0 = f_u_cla12_and275_f_u_cla12_and274_y0 & f_u_cla12_and275_f_u_cla12_and273_y0;
  assign f_u_cla12_and276_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and276_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and276_y0 = f_u_cla12_and276_f_u_cla12_pg_logic6_y0 & f_u_cla12_and276_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and277_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and277_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and277_y0 = f_u_cla12_and277_f_u_cla12_pg_logic7_y0 & f_u_cla12_and277_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and278_f_u_cla12_and277_y0 = f_u_cla12_and277_y0;
  assign f_u_cla12_and278_f_u_cla12_and276_y0 = f_u_cla12_and276_y0;
  assign f_u_cla12_and278_y0 = f_u_cla12_and278_f_u_cla12_and277_y0 & f_u_cla12_and278_f_u_cla12_and276_y0;
  assign f_u_cla12_and279_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and279_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and279_y0 = f_u_cla12_and279_f_u_cla12_pg_logic8_y0 & f_u_cla12_and279_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and280_f_u_cla12_and279_y0 = f_u_cla12_and279_y0;
  assign f_u_cla12_and280_f_u_cla12_and278_y0 = f_u_cla12_and278_y0;
  assign f_u_cla12_and280_y0 = f_u_cla12_and280_f_u_cla12_and279_y0 & f_u_cla12_and280_f_u_cla12_and278_y0;
  assign f_u_cla12_and281_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and281_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and281_y0 = f_u_cla12_and281_f_u_cla12_pg_logic7_y0 & f_u_cla12_and281_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and282_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and282_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and282_y0 = f_u_cla12_and282_f_u_cla12_pg_logic8_y0 & f_u_cla12_and282_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and283_f_u_cla12_and282_y0 = f_u_cla12_and282_y0;
  assign f_u_cla12_and283_f_u_cla12_and281_y0 = f_u_cla12_and281_y0;
  assign f_u_cla12_and283_y0 = f_u_cla12_and283_f_u_cla12_and282_y0 & f_u_cla12_and283_f_u_cla12_and281_y0;
  assign f_u_cla12_and284_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and284_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and284_y0 = f_u_cla12_and284_f_u_cla12_pg_logic8_y0 & f_u_cla12_and284_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_or36_f_u_cla12_and284_y0 = f_u_cla12_and284_y0;
  assign f_u_cla12_or36_f_u_cla12_and220_y0 = f_u_cla12_and220_y0;
  assign f_u_cla12_or36_y0 = f_u_cla12_or36_f_u_cla12_and284_y0 | f_u_cla12_or36_f_u_cla12_and220_y0;
  assign f_u_cla12_or37_f_u_cla12_or36_y0 = f_u_cla12_or36_y0;
  assign f_u_cla12_or37_f_u_cla12_and235_y0 = f_u_cla12_and235_y0;
  assign f_u_cla12_or37_y0 = f_u_cla12_or37_f_u_cla12_or36_y0 | f_u_cla12_or37_f_u_cla12_and235_y0;
  assign f_u_cla12_or38_f_u_cla12_or37_y0 = f_u_cla12_or37_y0;
  assign f_u_cla12_or38_f_u_cla12_and248_y0 = f_u_cla12_and248_y0;
  assign f_u_cla12_or38_y0 = f_u_cla12_or38_f_u_cla12_or37_y0 | f_u_cla12_or38_f_u_cla12_and248_y0;
  assign f_u_cla12_or39_f_u_cla12_or38_y0 = f_u_cla12_or38_y0;
  assign f_u_cla12_or39_f_u_cla12_and259_y0 = f_u_cla12_and259_y0;
  assign f_u_cla12_or39_y0 = f_u_cla12_or39_f_u_cla12_or38_y0 | f_u_cla12_or39_f_u_cla12_and259_y0;
  assign f_u_cla12_or40_f_u_cla12_or39_y0 = f_u_cla12_or39_y0;
  assign f_u_cla12_or40_f_u_cla12_and268_y0 = f_u_cla12_and268_y0;
  assign f_u_cla12_or40_y0 = f_u_cla12_or40_f_u_cla12_or39_y0 | f_u_cla12_or40_f_u_cla12_and268_y0;
  assign f_u_cla12_or41_f_u_cla12_or40_y0 = f_u_cla12_or40_y0;
  assign f_u_cla12_or41_f_u_cla12_and275_y0 = f_u_cla12_and275_y0;
  assign f_u_cla12_or41_y0 = f_u_cla12_or41_f_u_cla12_or40_y0 | f_u_cla12_or41_f_u_cla12_and275_y0;
  assign f_u_cla12_or42_f_u_cla12_or41_y0 = f_u_cla12_or41_y0;
  assign f_u_cla12_or42_f_u_cla12_and280_y0 = f_u_cla12_and280_y0;
  assign f_u_cla12_or42_y0 = f_u_cla12_or42_f_u_cla12_or41_y0 | f_u_cla12_or42_f_u_cla12_and280_y0;
  assign f_u_cla12_or43_f_u_cla12_or42_y0 = f_u_cla12_or42_y0;
  assign f_u_cla12_or43_f_u_cla12_and283_y0 = f_u_cla12_and283_y0;
  assign f_u_cla12_or43_y0 = f_u_cla12_or43_f_u_cla12_or42_y0 | f_u_cla12_or43_f_u_cla12_and283_y0;
  assign f_u_cla12_or44_f_u_cla12_pg_logic8_y1 = f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_or44_f_u_cla12_or43_y0 = f_u_cla12_or43_y0;
  assign f_u_cla12_or44_y0 = f_u_cla12_or44_f_u_cla12_pg_logic8_y1 | f_u_cla12_or44_f_u_cla12_or43_y0;
  assign f_u_cla12_pg_logic9_a_9 = a_9;
  assign f_u_cla12_pg_logic9_b_9 = b_9;
  assign f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_a_9 | f_u_cla12_pg_logic9_b_9;
  assign f_u_cla12_pg_logic9_y1 = f_u_cla12_pg_logic9_a_9 & f_u_cla12_pg_logic9_b_9;
  assign f_u_cla12_pg_logic9_y2 = f_u_cla12_pg_logic9_a_9 ^ f_u_cla12_pg_logic9_b_9;
  assign f_u_cla12_xor9_f_u_cla12_pg_logic9_y2 = f_u_cla12_pg_logic9_y2;
  assign f_u_cla12_xor9_f_u_cla12_or44_y0 = f_u_cla12_or44_y0;
  assign f_u_cla12_xor9_y0 = f_u_cla12_xor9_f_u_cla12_pg_logic9_y2 ^ f_u_cla12_xor9_f_u_cla12_or44_y0;
  assign f_u_cla12_and285_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and285_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and285_y0 = f_u_cla12_and285_f_u_cla12_pg_logic0_y0 & f_u_cla12_and285_constant_wire_0;
  assign f_u_cla12_and286_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and286_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and286_y0 = f_u_cla12_and286_f_u_cla12_pg_logic1_y0 & f_u_cla12_and286_constant_wire_0;
  assign f_u_cla12_and287_f_u_cla12_and286_y0 = f_u_cla12_and286_y0;
  assign f_u_cla12_and287_f_u_cla12_and285_y0 = f_u_cla12_and285_y0;
  assign f_u_cla12_and287_y0 = f_u_cla12_and287_f_u_cla12_and286_y0 & f_u_cla12_and287_f_u_cla12_and285_y0;
  assign f_u_cla12_and288_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and288_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and288_y0 = f_u_cla12_and288_f_u_cla12_pg_logic2_y0 & f_u_cla12_and288_constant_wire_0;
  assign f_u_cla12_and289_f_u_cla12_and288_y0 = f_u_cla12_and288_y0;
  assign f_u_cla12_and289_f_u_cla12_and287_y0 = f_u_cla12_and287_y0;
  assign f_u_cla12_and289_y0 = f_u_cla12_and289_f_u_cla12_and288_y0 & f_u_cla12_and289_f_u_cla12_and287_y0;
  assign f_u_cla12_and290_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and290_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and290_y0 = f_u_cla12_and290_f_u_cla12_pg_logic3_y0 & f_u_cla12_and290_constant_wire_0;
  assign f_u_cla12_and291_f_u_cla12_and290_y0 = f_u_cla12_and290_y0;
  assign f_u_cla12_and291_f_u_cla12_and289_y0 = f_u_cla12_and289_y0;
  assign f_u_cla12_and291_y0 = f_u_cla12_and291_f_u_cla12_and290_y0 & f_u_cla12_and291_f_u_cla12_and289_y0;
  assign f_u_cla12_and292_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and292_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and292_y0 = f_u_cla12_and292_f_u_cla12_pg_logic4_y0 & f_u_cla12_and292_constant_wire_0;
  assign f_u_cla12_and293_f_u_cla12_and292_y0 = f_u_cla12_and292_y0;
  assign f_u_cla12_and293_f_u_cla12_and291_y0 = f_u_cla12_and291_y0;
  assign f_u_cla12_and293_y0 = f_u_cla12_and293_f_u_cla12_and292_y0 & f_u_cla12_and293_f_u_cla12_and291_y0;
  assign f_u_cla12_and294_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and294_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and294_y0 = f_u_cla12_and294_f_u_cla12_pg_logic5_y0 & f_u_cla12_and294_constant_wire_0;
  assign f_u_cla12_and295_f_u_cla12_and294_y0 = f_u_cla12_and294_y0;
  assign f_u_cla12_and295_f_u_cla12_and293_y0 = f_u_cla12_and293_y0;
  assign f_u_cla12_and295_y0 = f_u_cla12_and295_f_u_cla12_and294_y0 & f_u_cla12_and295_f_u_cla12_and293_y0;
  assign f_u_cla12_and296_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and296_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and296_y0 = f_u_cla12_and296_f_u_cla12_pg_logic6_y0 & f_u_cla12_and296_constant_wire_0;
  assign f_u_cla12_and297_f_u_cla12_and296_y0 = f_u_cla12_and296_y0;
  assign f_u_cla12_and297_f_u_cla12_and295_y0 = f_u_cla12_and295_y0;
  assign f_u_cla12_and297_y0 = f_u_cla12_and297_f_u_cla12_and296_y0 & f_u_cla12_and297_f_u_cla12_and295_y0;
  assign f_u_cla12_and298_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and298_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and298_y0 = f_u_cla12_and298_f_u_cla12_pg_logic7_y0 & f_u_cla12_and298_constant_wire_0;
  assign f_u_cla12_and299_f_u_cla12_and298_y0 = f_u_cla12_and298_y0;
  assign f_u_cla12_and299_f_u_cla12_and297_y0 = f_u_cla12_and297_y0;
  assign f_u_cla12_and299_y0 = f_u_cla12_and299_f_u_cla12_and298_y0 & f_u_cla12_and299_f_u_cla12_and297_y0;
  assign f_u_cla12_and300_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and300_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and300_y0 = f_u_cla12_and300_f_u_cla12_pg_logic8_y0 & f_u_cla12_and300_constant_wire_0;
  assign f_u_cla12_and301_f_u_cla12_and300_y0 = f_u_cla12_and300_y0;
  assign f_u_cla12_and301_f_u_cla12_and299_y0 = f_u_cla12_and299_y0;
  assign f_u_cla12_and301_y0 = f_u_cla12_and301_f_u_cla12_and300_y0 & f_u_cla12_and301_f_u_cla12_and299_y0;
  assign f_u_cla12_and302_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and302_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and302_y0 = f_u_cla12_and302_f_u_cla12_pg_logic9_y0 & f_u_cla12_and302_constant_wire_0;
  assign f_u_cla12_and303_f_u_cla12_and302_y0 = f_u_cla12_and302_y0;
  assign f_u_cla12_and303_f_u_cla12_and301_y0 = f_u_cla12_and301_y0;
  assign f_u_cla12_and303_y0 = f_u_cla12_and303_f_u_cla12_and302_y0 & f_u_cla12_and303_f_u_cla12_and301_y0;
  assign f_u_cla12_and304_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and304_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and304_y0 = f_u_cla12_and304_f_u_cla12_pg_logic1_y0 & f_u_cla12_and304_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and305_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and305_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and305_y0 = f_u_cla12_and305_f_u_cla12_pg_logic2_y0 & f_u_cla12_and305_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and306_f_u_cla12_and305_y0 = f_u_cla12_and305_y0;
  assign f_u_cla12_and306_f_u_cla12_and304_y0 = f_u_cla12_and304_y0;
  assign f_u_cla12_and306_y0 = f_u_cla12_and306_f_u_cla12_and305_y0 & f_u_cla12_and306_f_u_cla12_and304_y0;
  assign f_u_cla12_and307_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and307_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and307_y0 = f_u_cla12_and307_f_u_cla12_pg_logic3_y0 & f_u_cla12_and307_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and308_f_u_cla12_and307_y0 = f_u_cla12_and307_y0;
  assign f_u_cla12_and308_f_u_cla12_and306_y0 = f_u_cla12_and306_y0;
  assign f_u_cla12_and308_y0 = f_u_cla12_and308_f_u_cla12_and307_y0 & f_u_cla12_and308_f_u_cla12_and306_y0;
  assign f_u_cla12_and309_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and309_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and309_y0 = f_u_cla12_and309_f_u_cla12_pg_logic4_y0 & f_u_cla12_and309_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and310_f_u_cla12_and309_y0 = f_u_cla12_and309_y0;
  assign f_u_cla12_and310_f_u_cla12_and308_y0 = f_u_cla12_and308_y0;
  assign f_u_cla12_and310_y0 = f_u_cla12_and310_f_u_cla12_and309_y0 & f_u_cla12_and310_f_u_cla12_and308_y0;
  assign f_u_cla12_and311_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and311_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and311_y0 = f_u_cla12_and311_f_u_cla12_pg_logic5_y0 & f_u_cla12_and311_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and312_f_u_cla12_and311_y0 = f_u_cla12_and311_y0;
  assign f_u_cla12_and312_f_u_cla12_and310_y0 = f_u_cla12_and310_y0;
  assign f_u_cla12_and312_y0 = f_u_cla12_and312_f_u_cla12_and311_y0 & f_u_cla12_and312_f_u_cla12_and310_y0;
  assign f_u_cla12_and313_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and313_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and313_y0 = f_u_cla12_and313_f_u_cla12_pg_logic6_y0 & f_u_cla12_and313_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and314_f_u_cla12_and313_y0 = f_u_cla12_and313_y0;
  assign f_u_cla12_and314_f_u_cla12_and312_y0 = f_u_cla12_and312_y0;
  assign f_u_cla12_and314_y0 = f_u_cla12_and314_f_u_cla12_and313_y0 & f_u_cla12_and314_f_u_cla12_and312_y0;
  assign f_u_cla12_and315_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and315_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and315_y0 = f_u_cla12_and315_f_u_cla12_pg_logic7_y0 & f_u_cla12_and315_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and316_f_u_cla12_and315_y0 = f_u_cla12_and315_y0;
  assign f_u_cla12_and316_f_u_cla12_and314_y0 = f_u_cla12_and314_y0;
  assign f_u_cla12_and316_y0 = f_u_cla12_and316_f_u_cla12_and315_y0 & f_u_cla12_and316_f_u_cla12_and314_y0;
  assign f_u_cla12_and317_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and317_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and317_y0 = f_u_cla12_and317_f_u_cla12_pg_logic8_y0 & f_u_cla12_and317_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and318_f_u_cla12_and317_y0 = f_u_cla12_and317_y0;
  assign f_u_cla12_and318_f_u_cla12_and316_y0 = f_u_cla12_and316_y0;
  assign f_u_cla12_and318_y0 = f_u_cla12_and318_f_u_cla12_and317_y0 & f_u_cla12_and318_f_u_cla12_and316_y0;
  assign f_u_cla12_and319_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and319_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and319_y0 = f_u_cla12_and319_f_u_cla12_pg_logic9_y0 & f_u_cla12_and319_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and320_f_u_cla12_and319_y0 = f_u_cla12_and319_y0;
  assign f_u_cla12_and320_f_u_cla12_and318_y0 = f_u_cla12_and318_y0;
  assign f_u_cla12_and320_y0 = f_u_cla12_and320_f_u_cla12_and319_y0 & f_u_cla12_and320_f_u_cla12_and318_y0;
  assign f_u_cla12_and321_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and321_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and321_y0 = f_u_cla12_and321_f_u_cla12_pg_logic2_y0 & f_u_cla12_and321_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and322_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and322_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and322_y0 = f_u_cla12_and322_f_u_cla12_pg_logic3_y0 & f_u_cla12_and322_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and323_f_u_cla12_and322_y0 = f_u_cla12_and322_y0;
  assign f_u_cla12_and323_f_u_cla12_and321_y0 = f_u_cla12_and321_y0;
  assign f_u_cla12_and323_y0 = f_u_cla12_and323_f_u_cla12_and322_y0 & f_u_cla12_and323_f_u_cla12_and321_y0;
  assign f_u_cla12_and324_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and324_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and324_y0 = f_u_cla12_and324_f_u_cla12_pg_logic4_y0 & f_u_cla12_and324_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and325_f_u_cla12_and324_y0 = f_u_cla12_and324_y0;
  assign f_u_cla12_and325_f_u_cla12_and323_y0 = f_u_cla12_and323_y0;
  assign f_u_cla12_and325_y0 = f_u_cla12_and325_f_u_cla12_and324_y0 & f_u_cla12_and325_f_u_cla12_and323_y0;
  assign f_u_cla12_and326_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and326_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and326_y0 = f_u_cla12_and326_f_u_cla12_pg_logic5_y0 & f_u_cla12_and326_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and327_f_u_cla12_and326_y0 = f_u_cla12_and326_y0;
  assign f_u_cla12_and327_f_u_cla12_and325_y0 = f_u_cla12_and325_y0;
  assign f_u_cla12_and327_y0 = f_u_cla12_and327_f_u_cla12_and326_y0 & f_u_cla12_and327_f_u_cla12_and325_y0;
  assign f_u_cla12_and328_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and328_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and328_y0 = f_u_cla12_and328_f_u_cla12_pg_logic6_y0 & f_u_cla12_and328_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and329_f_u_cla12_and328_y0 = f_u_cla12_and328_y0;
  assign f_u_cla12_and329_f_u_cla12_and327_y0 = f_u_cla12_and327_y0;
  assign f_u_cla12_and329_y0 = f_u_cla12_and329_f_u_cla12_and328_y0 & f_u_cla12_and329_f_u_cla12_and327_y0;
  assign f_u_cla12_and330_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and330_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and330_y0 = f_u_cla12_and330_f_u_cla12_pg_logic7_y0 & f_u_cla12_and330_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and331_f_u_cla12_and330_y0 = f_u_cla12_and330_y0;
  assign f_u_cla12_and331_f_u_cla12_and329_y0 = f_u_cla12_and329_y0;
  assign f_u_cla12_and331_y0 = f_u_cla12_and331_f_u_cla12_and330_y0 & f_u_cla12_and331_f_u_cla12_and329_y0;
  assign f_u_cla12_and332_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and332_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and332_y0 = f_u_cla12_and332_f_u_cla12_pg_logic8_y0 & f_u_cla12_and332_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and333_f_u_cla12_and332_y0 = f_u_cla12_and332_y0;
  assign f_u_cla12_and333_f_u_cla12_and331_y0 = f_u_cla12_and331_y0;
  assign f_u_cla12_and333_y0 = f_u_cla12_and333_f_u_cla12_and332_y0 & f_u_cla12_and333_f_u_cla12_and331_y0;
  assign f_u_cla12_and334_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and334_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and334_y0 = f_u_cla12_and334_f_u_cla12_pg_logic9_y0 & f_u_cla12_and334_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and335_f_u_cla12_and334_y0 = f_u_cla12_and334_y0;
  assign f_u_cla12_and335_f_u_cla12_and333_y0 = f_u_cla12_and333_y0;
  assign f_u_cla12_and335_y0 = f_u_cla12_and335_f_u_cla12_and334_y0 & f_u_cla12_and335_f_u_cla12_and333_y0;
  assign f_u_cla12_and336_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and336_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and336_y0 = f_u_cla12_and336_f_u_cla12_pg_logic3_y0 & f_u_cla12_and336_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and337_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and337_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and337_y0 = f_u_cla12_and337_f_u_cla12_pg_logic4_y0 & f_u_cla12_and337_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and338_f_u_cla12_and337_y0 = f_u_cla12_and337_y0;
  assign f_u_cla12_and338_f_u_cla12_and336_y0 = f_u_cla12_and336_y0;
  assign f_u_cla12_and338_y0 = f_u_cla12_and338_f_u_cla12_and337_y0 & f_u_cla12_and338_f_u_cla12_and336_y0;
  assign f_u_cla12_and339_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and339_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and339_y0 = f_u_cla12_and339_f_u_cla12_pg_logic5_y0 & f_u_cla12_and339_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and340_f_u_cla12_and339_y0 = f_u_cla12_and339_y0;
  assign f_u_cla12_and340_f_u_cla12_and338_y0 = f_u_cla12_and338_y0;
  assign f_u_cla12_and340_y0 = f_u_cla12_and340_f_u_cla12_and339_y0 & f_u_cla12_and340_f_u_cla12_and338_y0;
  assign f_u_cla12_and341_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and341_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and341_y0 = f_u_cla12_and341_f_u_cla12_pg_logic6_y0 & f_u_cla12_and341_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and342_f_u_cla12_and341_y0 = f_u_cla12_and341_y0;
  assign f_u_cla12_and342_f_u_cla12_and340_y0 = f_u_cla12_and340_y0;
  assign f_u_cla12_and342_y0 = f_u_cla12_and342_f_u_cla12_and341_y0 & f_u_cla12_and342_f_u_cla12_and340_y0;
  assign f_u_cla12_and343_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and343_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and343_y0 = f_u_cla12_and343_f_u_cla12_pg_logic7_y0 & f_u_cla12_and343_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and344_f_u_cla12_and343_y0 = f_u_cla12_and343_y0;
  assign f_u_cla12_and344_f_u_cla12_and342_y0 = f_u_cla12_and342_y0;
  assign f_u_cla12_and344_y0 = f_u_cla12_and344_f_u_cla12_and343_y0 & f_u_cla12_and344_f_u_cla12_and342_y0;
  assign f_u_cla12_and345_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and345_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and345_y0 = f_u_cla12_and345_f_u_cla12_pg_logic8_y0 & f_u_cla12_and345_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and346_f_u_cla12_and345_y0 = f_u_cla12_and345_y0;
  assign f_u_cla12_and346_f_u_cla12_and344_y0 = f_u_cla12_and344_y0;
  assign f_u_cla12_and346_y0 = f_u_cla12_and346_f_u_cla12_and345_y0 & f_u_cla12_and346_f_u_cla12_and344_y0;
  assign f_u_cla12_and347_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and347_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and347_y0 = f_u_cla12_and347_f_u_cla12_pg_logic9_y0 & f_u_cla12_and347_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and348_f_u_cla12_and347_y0 = f_u_cla12_and347_y0;
  assign f_u_cla12_and348_f_u_cla12_and346_y0 = f_u_cla12_and346_y0;
  assign f_u_cla12_and348_y0 = f_u_cla12_and348_f_u_cla12_and347_y0 & f_u_cla12_and348_f_u_cla12_and346_y0;
  assign f_u_cla12_and349_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and349_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and349_y0 = f_u_cla12_and349_f_u_cla12_pg_logic4_y0 & f_u_cla12_and349_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and350_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and350_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and350_y0 = f_u_cla12_and350_f_u_cla12_pg_logic5_y0 & f_u_cla12_and350_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and351_f_u_cla12_and350_y0 = f_u_cla12_and350_y0;
  assign f_u_cla12_and351_f_u_cla12_and349_y0 = f_u_cla12_and349_y0;
  assign f_u_cla12_and351_y0 = f_u_cla12_and351_f_u_cla12_and350_y0 & f_u_cla12_and351_f_u_cla12_and349_y0;
  assign f_u_cla12_and352_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and352_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and352_y0 = f_u_cla12_and352_f_u_cla12_pg_logic6_y0 & f_u_cla12_and352_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and353_f_u_cla12_and352_y0 = f_u_cla12_and352_y0;
  assign f_u_cla12_and353_f_u_cla12_and351_y0 = f_u_cla12_and351_y0;
  assign f_u_cla12_and353_y0 = f_u_cla12_and353_f_u_cla12_and352_y0 & f_u_cla12_and353_f_u_cla12_and351_y0;
  assign f_u_cla12_and354_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and354_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and354_y0 = f_u_cla12_and354_f_u_cla12_pg_logic7_y0 & f_u_cla12_and354_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and355_f_u_cla12_and354_y0 = f_u_cla12_and354_y0;
  assign f_u_cla12_and355_f_u_cla12_and353_y0 = f_u_cla12_and353_y0;
  assign f_u_cla12_and355_y0 = f_u_cla12_and355_f_u_cla12_and354_y0 & f_u_cla12_and355_f_u_cla12_and353_y0;
  assign f_u_cla12_and356_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and356_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and356_y0 = f_u_cla12_and356_f_u_cla12_pg_logic8_y0 & f_u_cla12_and356_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and357_f_u_cla12_and356_y0 = f_u_cla12_and356_y0;
  assign f_u_cla12_and357_f_u_cla12_and355_y0 = f_u_cla12_and355_y0;
  assign f_u_cla12_and357_y0 = f_u_cla12_and357_f_u_cla12_and356_y0 & f_u_cla12_and357_f_u_cla12_and355_y0;
  assign f_u_cla12_and358_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and358_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and358_y0 = f_u_cla12_and358_f_u_cla12_pg_logic9_y0 & f_u_cla12_and358_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and359_f_u_cla12_and358_y0 = f_u_cla12_and358_y0;
  assign f_u_cla12_and359_f_u_cla12_and357_y0 = f_u_cla12_and357_y0;
  assign f_u_cla12_and359_y0 = f_u_cla12_and359_f_u_cla12_and358_y0 & f_u_cla12_and359_f_u_cla12_and357_y0;
  assign f_u_cla12_and360_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and360_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and360_y0 = f_u_cla12_and360_f_u_cla12_pg_logic5_y0 & f_u_cla12_and360_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and361_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and361_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and361_y0 = f_u_cla12_and361_f_u_cla12_pg_logic6_y0 & f_u_cla12_and361_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and362_f_u_cla12_and361_y0 = f_u_cla12_and361_y0;
  assign f_u_cla12_and362_f_u_cla12_and360_y0 = f_u_cla12_and360_y0;
  assign f_u_cla12_and362_y0 = f_u_cla12_and362_f_u_cla12_and361_y0 & f_u_cla12_and362_f_u_cla12_and360_y0;
  assign f_u_cla12_and363_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and363_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and363_y0 = f_u_cla12_and363_f_u_cla12_pg_logic7_y0 & f_u_cla12_and363_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and364_f_u_cla12_and363_y0 = f_u_cla12_and363_y0;
  assign f_u_cla12_and364_f_u_cla12_and362_y0 = f_u_cla12_and362_y0;
  assign f_u_cla12_and364_y0 = f_u_cla12_and364_f_u_cla12_and363_y0 & f_u_cla12_and364_f_u_cla12_and362_y0;
  assign f_u_cla12_and365_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and365_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and365_y0 = f_u_cla12_and365_f_u_cla12_pg_logic8_y0 & f_u_cla12_and365_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and366_f_u_cla12_and365_y0 = f_u_cla12_and365_y0;
  assign f_u_cla12_and366_f_u_cla12_and364_y0 = f_u_cla12_and364_y0;
  assign f_u_cla12_and366_y0 = f_u_cla12_and366_f_u_cla12_and365_y0 & f_u_cla12_and366_f_u_cla12_and364_y0;
  assign f_u_cla12_and367_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and367_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and367_y0 = f_u_cla12_and367_f_u_cla12_pg_logic9_y0 & f_u_cla12_and367_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and368_f_u_cla12_and367_y0 = f_u_cla12_and367_y0;
  assign f_u_cla12_and368_f_u_cla12_and366_y0 = f_u_cla12_and366_y0;
  assign f_u_cla12_and368_y0 = f_u_cla12_and368_f_u_cla12_and367_y0 & f_u_cla12_and368_f_u_cla12_and366_y0;
  assign f_u_cla12_and369_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and369_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and369_y0 = f_u_cla12_and369_f_u_cla12_pg_logic6_y0 & f_u_cla12_and369_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and370_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and370_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and370_y0 = f_u_cla12_and370_f_u_cla12_pg_logic7_y0 & f_u_cla12_and370_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and371_f_u_cla12_and370_y0 = f_u_cla12_and370_y0;
  assign f_u_cla12_and371_f_u_cla12_and369_y0 = f_u_cla12_and369_y0;
  assign f_u_cla12_and371_y0 = f_u_cla12_and371_f_u_cla12_and370_y0 & f_u_cla12_and371_f_u_cla12_and369_y0;
  assign f_u_cla12_and372_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and372_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and372_y0 = f_u_cla12_and372_f_u_cla12_pg_logic8_y0 & f_u_cla12_and372_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and373_f_u_cla12_and372_y0 = f_u_cla12_and372_y0;
  assign f_u_cla12_and373_f_u_cla12_and371_y0 = f_u_cla12_and371_y0;
  assign f_u_cla12_and373_y0 = f_u_cla12_and373_f_u_cla12_and372_y0 & f_u_cla12_and373_f_u_cla12_and371_y0;
  assign f_u_cla12_and374_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and374_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and374_y0 = f_u_cla12_and374_f_u_cla12_pg_logic9_y0 & f_u_cla12_and374_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and375_f_u_cla12_and374_y0 = f_u_cla12_and374_y0;
  assign f_u_cla12_and375_f_u_cla12_and373_y0 = f_u_cla12_and373_y0;
  assign f_u_cla12_and375_y0 = f_u_cla12_and375_f_u_cla12_and374_y0 & f_u_cla12_and375_f_u_cla12_and373_y0;
  assign f_u_cla12_and376_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and376_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and376_y0 = f_u_cla12_and376_f_u_cla12_pg_logic7_y0 & f_u_cla12_and376_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and377_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and377_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and377_y0 = f_u_cla12_and377_f_u_cla12_pg_logic8_y0 & f_u_cla12_and377_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and378_f_u_cla12_and377_y0 = f_u_cla12_and377_y0;
  assign f_u_cla12_and378_f_u_cla12_and376_y0 = f_u_cla12_and376_y0;
  assign f_u_cla12_and378_y0 = f_u_cla12_and378_f_u_cla12_and377_y0 & f_u_cla12_and378_f_u_cla12_and376_y0;
  assign f_u_cla12_and379_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and379_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and379_y0 = f_u_cla12_and379_f_u_cla12_pg_logic9_y0 & f_u_cla12_and379_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and380_f_u_cla12_and379_y0 = f_u_cla12_and379_y0;
  assign f_u_cla12_and380_f_u_cla12_and378_y0 = f_u_cla12_and378_y0;
  assign f_u_cla12_and380_y0 = f_u_cla12_and380_f_u_cla12_and379_y0 & f_u_cla12_and380_f_u_cla12_and378_y0;
  assign f_u_cla12_and381_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and381_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and381_y0 = f_u_cla12_and381_f_u_cla12_pg_logic8_y0 & f_u_cla12_and381_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and382_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and382_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and382_y0 = f_u_cla12_and382_f_u_cla12_pg_logic9_y0 & f_u_cla12_and382_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and383_f_u_cla12_and382_y0 = f_u_cla12_and382_y0;
  assign f_u_cla12_and383_f_u_cla12_and381_y0 = f_u_cla12_and381_y0;
  assign f_u_cla12_and383_y0 = f_u_cla12_and383_f_u_cla12_and382_y0 & f_u_cla12_and383_f_u_cla12_and381_y0;
  assign f_u_cla12_and384_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and384_f_u_cla12_pg_logic8_y1 = f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and384_y0 = f_u_cla12_and384_f_u_cla12_pg_logic9_y0 & f_u_cla12_and384_f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_or45_f_u_cla12_and384_y0 = f_u_cla12_and384_y0;
  assign f_u_cla12_or45_f_u_cla12_and303_y0 = f_u_cla12_and303_y0;
  assign f_u_cla12_or45_y0 = f_u_cla12_or45_f_u_cla12_and384_y0 | f_u_cla12_or45_f_u_cla12_and303_y0;
  assign f_u_cla12_or46_f_u_cla12_or45_y0 = f_u_cla12_or45_y0;
  assign f_u_cla12_or46_f_u_cla12_and320_y0 = f_u_cla12_and320_y0;
  assign f_u_cla12_or46_y0 = f_u_cla12_or46_f_u_cla12_or45_y0 | f_u_cla12_or46_f_u_cla12_and320_y0;
  assign f_u_cla12_or47_f_u_cla12_or46_y0 = f_u_cla12_or46_y0;
  assign f_u_cla12_or47_f_u_cla12_and335_y0 = f_u_cla12_and335_y0;
  assign f_u_cla12_or47_y0 = f_u_cla12_or47_f_u_cla12_or46_y0 | f_u_cla12_or47_f_u_cla12_and335_y0;
  assign f_u_cla12_or48_f_u_cla12_or47_y0 = f_u_cla12_or47_y0;
  assign f_u_cla12_or48_f_u_cla12_and348_y0 = f_u_cla12_and348_y0;
  assign f_u_cla12_or48_y0 = f_u_cla12_or48_f_u_cla12_or47_y0 | f_u_cla12_or48_f_u_cla12_and348_y0;
  assign f_u_cla12_or49_f_u_cla12_or48_y0 = f_u_cla12_or48_y0;
  assign f_u_cla12_or49_f_u_cla12_and359_y0 = f_u_cla12_and359_y0;
  assign f_u_cla12_or49_y0 = f_u_cla12_or49_f_u_cla12_or48_y0 | f_u_cla12_or49_f_u_cla12_and359_y0;
  assign f_u_cla12_or50_f_u_cla12_or49_y0 = f_u_cla12_or49_y0;
  assign f_u_cla12_or50_f_u_cla12_and368_y0 = f_u_cla12_and368_y0;
  assign f_u_cla12_or50_y0 = f_u_cla12_or50_f_u_cla12_or49_y0 | f_u_cla12_or50_f_u_cla12_and368_y0;
  assign f_u_cla12_or51_f_u_cla12_or50_y0 = f_u_cla12_or50_y0;
  assign f_u_cla12_or51_f_u_cla12_and375_y0 = f_u_cla12_and375_y0;
  assign f_u_cla12_or51_y0 = f_u_cla12_or51_f_u_cla12_or50_y0 | f_u_cla12_or51_f_u_cla12_and375_y0;
  assign f_u_cla12_or52_f_u_cla12_or51_y0 = f_u_cla12_or51_y0;
  assign f_u_cla12_or52_f_u_cla12_and380_y0 = f_u_cla12_and380_y0;
  assign f_u_cla12_or52_y0 = f_u_cla12_or52_f_u_cla12_or51_y0 | f_u_cla12_or52_f_u_cla12_and380_y0;
  assign f_u_cla12_or53_f_u_cla12_or52_y0 = f_u_cla12_or52_y0;
  assign f_u_cla12_or53_f_u_cla12_and383_y0 = f_u_cla12_and383_y0;
  assign f_u_cla12_or53_y0 = f_u_cla12_or53_f_u_cla12_or52_y0 | f_u_cla12_or53_f_u_cla12_and383_y0;
  assign f_u_cla12_or54_f_u_cla12_pg_logic9_y1 = f_u_cla12_pg_logic9_y1;
  assign f_u_cla12_or54_f_u_cla12_or53_y0 = f_u_cla12_or53_y0;
  assign f_u_cla12_or54_y0 = f_u_cla12_or54_f_u_cla12_pg_logic9_y1 | f_u_cla12_or54_f_u_cla12_or53_y0;
  assign f_u_cla12_pg_logic10_a_10 = a_10;
  assign f_u_cla12_pg_logic10_b_10 = b_10;
  assign f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_a_10 | f_u_cla12_pg_logic10_b_10;
  assign f_u_cla12_pg_logic10_y1 = f_u_cla12_pg_logic10_a_10 & f_u_cla12_pg_logic10_b_10;
  assign f_u_cla12_pg_logic10_y2 = f_u_cla12_pg_logic10_a_10 ^ f_u_cla12_pg_logic10_b_10;
  assign f_u_cla12_xor10_f_u_cla12_pg_logic10_y2 = f_u_cla12_pg_logic10_y2;
  assign f_u_cla12_xor10_f_u_cla12_or54_y0 = f_u_cla12_or54_y0;
  assign f_u_cla12_xor10_y0 = f_u_cla12_xor10_f_u_cla12_pg_logic10_y2 ^ f_u_cla12_xor10_f_u_cla12_or54_y0;
  assign f_u_cla12_and385_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and385_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and385_y0 = f_u_cla12_and385_f_u_cla12_pg_logic0_y0 & f_u_cla12_and385_constant_wire_0;
  assign f_u_cla12_and386_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and386_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and386_y0 = f_u_cla12_and386_f_u_cla12_pg_logic1_y0 & f_u_cla12_and386_constant_wire_0;
  assign f_u_cla12_and387_f_u_cla12_and386_y0 = f_u_cla12_and386_y0;
  assign f_u_cla12_and387_f_u_cla12_and385_y0 = f_u_cla12_and385_y0;
  assign f_u_cla12_and387_y0 = f_u_cla12_and387_f_u_cla12_and386_y0 & f_u_cla12_and387_f_u_cla12_and385_y0;
  assign f_u_cla12_and388_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and388_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and388_y0 = f_u_cla12_and388_f_u_cla12_pg_logic2_y0 & f_u_cla12_and388_constant_wire_0;
  assign f_u_cla12_and389_f_u_cla12_and388_y0 = f_u_cla12_and388_y0;
  assign f_u_cla12_and389_f_u_cla12_and387_y0 = f_u_cla12_and387_y0;
  assign f_u_cla12_and389_y0 = f_u_cla12_and389_f_u_cla12_and388_y0 & f_u_cla12_and389_f_u_cla12_and387_y0;
  assign f_u_cla12_and390_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and390_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and390_y0 = f_u_cla12_and390_f_u_cla12_pg_logic3_y0 & f_u_cla12_and390_constant_wire_0;
  assign f_u_cla12_and391_f_u_cla12_and390_y0 = f_u_cla12_and390_y0;
  assign f_u_cla12_and391_f_u_cla12_and389_y0 = f_u_cla12_and389_y0;
  assign f_u_cla12_and391_y0 = f_u_cla12_and391_f_u_cla12_and390_y0 & f_u_cla12_and391_f_u_cla12_and389_y0;
  assign f_u_cla12_and392_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and392_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and392_y0 = f_u_cla12_and392_f_u_cla12_pg_logic4_y0 & f_u_cla12_and392_constant_wire_0;
  assign f_u_cla12_and393_f_u_cla12_and392_y0 = f_u_cla12_and392_y0;
  assign f_u_cla12_and393_f_u_cla12_and391_y0 = f_u_cla12_and391_y0;
  assign f_u_cla12_and393_y0 = f_u_cla12_and393_f_u_cla12_and392_y0 & f_u_cla12_and393_f_u_cla12_and391_y0;
  assign f_u_cla12_and394_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and394_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and394_y0 = f_u_cla12_and394_f_u_cla12_pg_logic5_y0 & f_u_cla12_and394_constant_wire_0;
  assign f_u_cla12_and395_f_u_cla12_and394_y0 = f_u_cla12_and394_y0;
  assign f_u_cla12_and395_f_u_cla12_and393_y0 = f_u_cla12_and393_y0;
  assign f_u_cla12_and395_y0 = f_u_cla12_and395_f_u_cla12_and394_y0 & f_u_cla12_and395_f_u_cla12_and393_y0;
  assign f_u_cla12_and396_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and396_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and396_y0 = f_u_cla12_and396_f_u_cla12_pg_logic6_y0 & f_u_cla12_and396_constant_wire_0;
  assign f_u_cla12_and397_f_u_cla12_and396_y0 = f_u_cla12_and396_y0;
  assign f_u_cla12_and397_f_u_cla12_and395_y0 = f_u_cla12_and395_y0;
  assign f_u_cla12_and397_y0 = f_u_cla12_and397_f_u_cla12_and396_y0 & f_u_cla12_and397_f_u_cla12_and395_y0;
  assign f_u_cla12_and398_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and398_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and398_y0 = f_u_cla12_and398_f_u_cla12_pg_logic7_y0 & f_u_cla12_and398_constant_wire_0;
  assign f_u_cla12_and399_f_u_cla12_and398_y0 = f_u_cla12_and398_y0;
  assign f_u_cla12_and399_f_u_cla12_and397_y0 = f_u_cla12_and397_y0;
  assign f_u_cla12_and399_y0 = f_u_cla12_and399_f_u_cla12_and398_y0 & f_u_cla12_and399_f_u_cla12_and397_y0;
  assign f_u_cla12_and400_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and400_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and400_y0 = f_u_cla12_and400_f_u_cla12_pg_logic8_y0 & f_u_cla12_and400_constant_wire_0;
  assign f_u_cla12_and401_f_u_cla12_and400_y0 = f_u_cla12_and400_y0;
  assign f_u_cla12_and401_f_u_cla12_and399_y0 = f_u_cla12_and399_y0;
  assign f_u_cla12_and401_y0 = f_u_cla12_and401_f_u_cla12_and400_y0 & f_u_cla12_and401_f_u_cla12_and399_y0;
  assign f_u_cla12_and402_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and402_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and402_y0 = f_u_cla12_and402_f_u_cla12_pg_logic9_y0 & f_u_cla12_and402_constant_wire_0;
  assign f_u_cla12_and403_f_u_cla12_and402_y0 = f_u_cla12_and402_y0;
  assign f_u_cla12_and403_f_u_cla12_and401_y0 = f_u_cla12_and401_y0;
  assign f_u_cla12_and403_y0 = f_u_cla12_and403_f_u_cla12_and402_y0 & f_u_cla12_and403_f_u_cla12_and401_y0;
  assign f_u_cla12_and404_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and404_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and404_y0 = f_u_cla12_and404_f_u_cla12_pg_logic10_y0 & f_u_cla12_and404_constant_wire_0;
  assign f_u_cla12_and405_f_u_cla12_and404_y0 = f_u_cla12_and404_y0;
  assign f_u_cla12_and405_f_u_cla12_and403_y0 = f_u_cla12_and403_y0;
  assign f_u_cla12_and405_y0 = f_u_cla12_and405_f_u_cla12_and404_y0 & f_u_cla12_and405_f_u_cla12_and403_y0;
  assign f_u_cla12_and406_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and406_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and406_y0 = f_u_cla12_and406_f_u_cla12_pg_logic1_y0 & f_u_cla12_and406_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and407_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and407_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and407_y0 = f_u_cla12_and407_f_u_cla12_pg_logic2_y0 & f_u_cla12_and407_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and408_f_u_cla12_and407_y0 = f_u_cla12_and407_y0;
  assign f_u_cla12_and408_f_u_cla12_and406_y0 = f_u_cla12_and406_y0;
  assign f_u_cla12_and408_y0 = f_u_cla12_and408_f_u_cla12_and407_y0 & f_u_cla12_and408_f_u_cla12_and406_y0;
  assign f_u_cla12_and409_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and409_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and409_y0 = f_u_cla12_and409_f_u_cla12_pg_logic3_y0 & f_u_cla12_and409_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and410_f_u_cla12_and409_y0 = f_u_cla12_and409_y0;
  assign f_u_cla12_and410_f_u_cla12_and408_y0 = f_u_cla12_and408_y0;
  assign f_u_cla12_and410_y0 = f_u_cla12_and410_f_u_cla12_and409_y0 & f_u_cla12_and410_f_u_cla12_and408_y0;
  assign f_u_cla12_and411_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and411_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and411_y0 = f_u_cla12_and411_f_u_cla12_pg_logic4_y0 & f_u_cla12_and411_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and412_f_u_cla12_and411_y0 = f_u_cla12_and411_y0;
  assign f_u_cla12_and412_f_u_cla12_and410_y0 = f_u_cla12_and410_y0;
  assign f_u_cla12_and412_y0 = f_u_cla12_and412_f_u_cla12_and411_y0 & f_u_cla12_and412_f_u_cla12_and410_y0;
  assign f_u_cla12_and413_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and413_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and413_y0 = f_u_cla12_and413_f_u_cla12_pg_logic5_y0 & f_u_cla12_and413_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and414_f_u_cla12_and413_y0 = f_u_cla12_and413_y0;
  assign f_u_cla12_and414_f_u_cla12_and412_y0 = f_u_cla12_and412_y0;
  assign f_u_cla12_and414_y0 = f_u_cla12_and414_f_u_cla12_and413_y0 & f_u_cla12_and414_f_u_cla12_and412_y0;
  assign f_u_cla12_and415_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and415_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and415_y0 = f_u_cla12_and415_f_u_cla12_pg_logic6_y0 & f_u_cla12_and415_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and416_f_u_cla12_and415_y0 = f_u_cla12_and415_y0;
  assign f_u_cla12_and416_f_u_cla12_and414_y0 = f_u_cla12_and414_y0;
  assign f_u_cla12_and416_y0 = f_u_cla12_and416_f_u_cla12_and415_y0 & f_u_cla12_and416_f_u_cla12_and414_y0;
  assign f_u_cla12_and417_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and417_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and417_y0 = f_u_cla12_and417_f_u_cla12_pg_logic7_y0 & f_u_cla12_and417_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and418_f_u_cla12_and417_y0 = f_u_cla12_and417_y0;
  assign f_u_cla12_and418_f_u_cla12_and416_y0 = f_u_cla12_and416_y0;
  assign f_u_cla12_and418_y0 = f_u_cla12_and418_f_u_cla12_and417_y0 & f_u_cla12_and418_f_u_cla12_and416_y0;
  assign f_u_cla12_and419_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and419_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and419_y0 = f_u_cla12_and419_f_u_cla12_pg_logic8_y0 & f_u_cla12_and419_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and420_f_u_cla12_and419_y0 = f_u_cla12_and419_y0;
  assign f_u_cla12_and420_f_u_cla12_and418_y0 = f_u_cla12_and418_y0;
  assign f_u_cla12_and420_y0 = f_u_cla12_and420_f_u_cla12_and419_y0 & f_u_cla12_and420_f_u_cla12_and418_y0;
  assign f_u_cla12_and421_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and421_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and421_y0 = f_u_cla12_and421_f_u_cla12_pg_logic9_y0 & f_u_cla12_and421_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and422_f_u_cla12_and421_y0 = f_u_cla12_and421_y0;
  assign f_u_cla12_and422_f_u_cla12_and420_y0 = f_u_cla12_and420_y0;
  assign f_u_cla12_and422_y0 = f_u_cla12_and422_f_u_cla12_and421_y0 & f_u_cla12_and422_f_u_cla12_and420_y0;
  assign f_u_cla12_and423_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and423_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and423_y0 = f_u_cla12_and423_f_u_cla12_pg_logic10_y0 & f_u_cla12_and423_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and424_f_u_cla12_and423_y0 = f_u_cla12_and423_y0;
  assign f_u_cla12_and424_f_u_cla12_and422_y0 = f_u_cla12_and422_y0;
  assign f_u_cla12_and424_y0 = f_u_cla12_and424_f_u_cla12_and423_y0 & f_u_cla12_and424_f_u_cla12_and422_y0;
  assign f_u_cla12_and425_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and425_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and425_y0 = f_u_cla12_and425_f_u_cla12_pg_logic2_y0 & f_u_cla12_and425_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and426_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and426_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and426_y0 = f_u_cla12_and426_f_u_cla12_pg_logic3_y0 & f_u_cla12_and426_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and427_f_u_cla12_and426_y0 = f_u_cla12_and426_y0;
  assign f_u_cla12_and427_f_u_cla12_and425_y0 = f_u_cla12_and425_y0;
  assign f_u_cla12_and427_y0 = f_u_cla12_and427_f_u_cla12_and426_y0 & f_u_cla12_and427_f_u_cla12_and425_y0;
  assign f_u_cla12_and428_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and428_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and428_y0 = f_u_cla12_and428_f_u_cla12_pg_logic4_y0 & f_u_cla12_and428_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and429_f_u_cla12_and428_y0 = f_u_cla12_and428_y0;
  assign f_u_cla12_and429_f_u_cla12_and427_y0 = f_u_cla12_and427_y0;
  assign f_u_cla12_and429_y0 = f_u_cla12_and429_f_u_cla12_and428_y0 & f_u_cla12_and429_f_u_cla12_and427_y0;
  assign f_u_cla12_and430_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and430_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and430_y0 = f_u_cla12_and430_f_u_cla12_pg_logic5_y0 & f_u_cla12_and430_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and431_f_u_cla12_and430_y0 = f_u_cla12_and430_y0;
  assign f_u_cla12_and431_f_u_cla12_and429_y0 = f_u_cla12_and429_y0;
  assign f_u_cla12_and431_y0 = f_u_cla12_and431_f_u_cla12_and430_y0 & f_u_cla12_and431_f_u_cla12_and429_y0;
  assign f_u_cla12_and432_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and432_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and432_y0 = f_u_cla12_and432_f_u_cla12_pg_logic6_y0 & f_u_cla12_and432_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and433_f_u_cla12_and432_y0 = f_u_cla12_and432_y0;
  assign f_u_cla12_and433_f_u_cla12_and431_y0 = f_u_cla12_and431_y0;
  assign f_u_cla12_and433_y0 = f_u_cla12_and433_f_u_cla12_and432_y0 & f_u_cla12_and433_f_u_cla12_and431_y0;
  assign f_u_cla12_and434_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and434_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and434_y0 = f_u_cla12_and434_f_u_cla12_pg_logic7_y0 & f_u_cla12_and434_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and435_f_u_cla12_and434_y0 = f_u_cla12_and434_y0;
  assign f_u_cla12_and435_f_u_cla12_and433_y0 = f_u_cla12_and433_y0;
  assign f_u_cla12_and435_y0 = f_u_cla12_and435_f_u_cla12_and434_y0 & f_u_cla12_and435_f_u_cla12_and433_y0;
  assign f_u_cla12_and436_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and436_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and436_y0 = f_u_cla12_and436_f_u_cla12_pg_logic8_y0 & f_u_cla12_and436_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and437_f_u_cla12_and436_y0 = f_u_cla12_and436_y0;
  assign f_u_cla12_and437_f_u_cla12_and435_y0 = f_u_cla12_and435_y0;
  assign f_u_cla12_and437_y0 = f_u_cla12_and437_f_u_cla12_and436_y0 & f_u_cla12_and437_f_u_cla12_and435_y0;
  assign f_u_cla12_and438_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and438_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and438_y0 = f_u_cla12_and438_f_u_cla12_pg_logic9_y0 & f_u_cla12_and438_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and439_f_u_cla12_and438_y0 = f_u_cla12_and438_y0;
  assign f_u_cla12_and439_f_u_cla12_and437_y0 = f_u_cla12_and437_y0;
  assign f_u_cla12_and439_y0 = f_u_cla12_and439_f_u_cla12_and438_y0 & f_u_cla12_and439_f_u_cla12_and437_y0;
  assign f_u_cla12_and440_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and440_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and440_y0 = f_u_cla12_and440_f_u_cla12_pg_logic10_y0 & f_u_cla12_and440_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and441_f_u_cla12_and440_y0 = f_u_cla12_and440_y0;
  assign f_u_cla12_and441_f_u_cla12_and439_y0 = f_u_cla12_and439_y0;
  assign f_u_cla12_and441_y0 = f_u_cla12_and441_f_u_cla12_and440_y0 & f_u_cla12_and441_f_u_cla12_and439_y0;
  assign f_u_cla12_and442_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and442_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and442_y0 = f_u_cla12_and442_f_u_cla12_pg_logic3_y0 & f_u_cla12_and442_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and443_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and443_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and443_y0 = f_u_cla12_and443_f_u_cla12_pg_logic4_y0 & f_u_cla12_and443_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and444_f_u_cla12_and443_y0 = f_u_cla12_and443_y0;
  assign f_u_cla12_and444_f_u_cla12_and442_y0 = f_u_cla12_and442_y0;
  assign f_u_cla12_and444_y0 = f_u_cla12_and444_f_u_cla12_and443_y0 & f_u_cla12_and444_f_u_cla12_and442_y0;
  assign f_u_cla12_and445_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and445_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and445_y0 = f_u_cla12_and445_f_u_cla12_pg_logic5_y0 & f_u_cla12_and445_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and446_f_u_cla12_and445_y0 = f_u_cla12_and445_y0;
  assign f_u_cla12_and446_f_u_cla12_and444_y0 = f_u_cla12_and444_y0;
  assign f_u_cla12_and446_y0 = f_u_cla12_and446_f_u_cla12_and445_y0 & f_u_cla12_and446_f_u_cla12_and444_y0;
  assign f_u_cla12_and447_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and447_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and447_y0 = f_u_cla12_and447_f_u_cla12_pg_logic6_y0 & f_u_cla12_and447_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and448_f_u_cla12_and447_y0 = f_u_cla12_and447_y0;
  assign f_u_cla12_and448_f_u_cla12_and446_y0 = f_u_cla12_and446_y0;
  assign f_u_cla12_and448_y0 = f_u_cla12_and448_f_u_cla12_and447_y0 & f_u_cla12_and448_f_u_cla12_and446_y0;
  assign f_u_cla12_and449_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and449_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and449_y0 = f_u_cla12_and449_f_u_cla12_pg_logic7_y0 & f_u_cla12_and449_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and450_f_u_cla12_and449_y0 = f_u_cla12_and449_y0;
  assign f_u_cla12_and450_f_u_cla12_and448_y0 = f_u_cla12_and448_y0;
  assign f_u_cla12_and450_y0 = f_u_cla12_and450_f_u_cla12_and449_y0 & f_u_cla12_and450_f_u_cla12_and448_y0;
  assign f_u_cla12_and451_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and451_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and451_y0 = f_u_cla12_and451_f_u_cla12_pg_logic8_y0 & f_u_cla12_and451_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and452_f_u_cla12_and451_y0 = f_u_cla12_and451_y0;
  assign f_u_cla12_and452_f_u_cla12_and450_y0 = f_u_cla12_and450_y0;
  assign f_u_cla12_and452_y0 = f_u_cla12_and452_f_u_cla12_and451_y0 & f_u_cla12_and452_f_u_cla12_and450_y0;
  assign f_u_cla12_and453_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and453_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and453_y0 = f_u_cla12_and453_f_u_cla12_pg_logic9_y0 & f_u_cla12_and453_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and454_f_u_cla12_and453_y0 = f_u_cla12_and453_y0;
  assign f_u_cla12_and454_f_u_cla12_and452_y0 = f_u_cla12_and452_y0;
  assign f_u_cla12_and454_y0 = f_u_cla12_and454_f_u_cla12_and453_y0 & f_u_cla12_and454_f_u_cla12_and452_y0;
  assign f_u_cla12_and455_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and455_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and455_y0 = f_u_cla12_and455_f_u_cla12_pg_logic10_y0 & f_u_cla12_and455_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and456_f_u_cla12_and455_y0 = f_u_cla12_and455_y0;
  assign f_u_cla12_and456_f_u_cla12_and454_y0 = f_u_cla12_and454_y0;
  assign f_u_cla12_and456_y0 = f_u_cla12_and456_f_u_cla12_and455_y0 & f_u_cla12_and456_f_u_cla12_and454_y0;
  assign f_u_cla12_and457_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and457_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and457_y0 = f_u_cla12_and457_f_u_cla12_pg_logic4_y0 & f_u_cla12_and457_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and458_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and458_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and458_y0 = f_u_cla12_and458_f_u_cla12_pg_logic5_y0 & f_u_cla12_and458_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and459_f_u_cla12_and458_y0 = f_u_cla12_and458_y0;
  assign f_u_cla12_and459_f_u_cla12_and457_y0 = f_u_cla12_and457_y0;
  assign f_u_cla12_and459_y0 = f_u_cla12_and459_f_u_cla12_and458_y0 & f_u_cla12_and459_f_u_cla12_and457_y0;
  assign f_u_cla12_and460_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and460_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and460_y0 = f_u_cla12_and460_f_u_cla12_pg_logic6_y0 & f_u_cla12_and460_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and461_f_u_cla12_and460_y0 = f_u_cla12_and460_y0;
  assign f_u_cla12_and461_f_u_cla12_and459_y0 = f_u_cla12_and459_y0;
  assign f_u_cla12_and461_y0 = f_u_cla12_and461_f_u_cla12_and460_y0 & f_u_cla12_and461_f_u_cla12_and459_y0;
  assign f_u_cla12_and462_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and462_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and462_y0 = f_u_cla12_and462_f_u_cla12_pg_logic7_y0 & f_u_cla12_and462_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and463_f_u_cla12_and462_y0 = f_u_cla12_and462_y0;
  assign f_u_cla12_and463_f_u_cla12_and461_y0 = f_u_cla12_and461_y0;
  assign f_u_cla12_and463_y0 = f_u_cla12_and463_f_u_cla12_and462_y0 & f_u_cla12_and463_f_u_cla12_and461_y0;
  assign f_u_cla12_and464_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and464_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and464_y0 = f_u_cla12_and464_f_u_cla12_pg_logic8_y0 & f_u_cla12_and464_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and465_f_u_cla12_and464_y0 = f_u_cla12_and464_y0;
  assign f_u_cla12_and465_f_u_cla12_and463_y0 = f_u_cla12_and463_y0;
  assign f_u_cla12_and465_y0 = f_u_cla12_and465_f_u_cla12_and464_y0 & f_u_cla12_and465_f_u_cla12_and463_y0;
  assign f_u_cla12_and466_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and466_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and466_y0 = f_u_cla12_and466_f_u_cla12_pg_logic9_y0 & f_u_cla12_and466_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and467_f_u_cla12_and466_y0 = f_u_cla12_and466_y0;
  assign f_u_cla12_and467_f_u_cla12_and465_y0 = f_u_cla12_and465_y0;
  assign f_u_cla12_and467_y0 = f_u_cla12_and467_f_u_cla12_and466_y0 & f_u_cla12_and467_f_u_cla12_and465_y0;
  assign f_u_cla12_and468_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and468_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and468_y0 = f_u_cla12_and468_f_u_cla12_pg_logic10_y0 & f_u_cla12_and468_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and469_f_u_cla12_and468_y0 = f_u_cla12_and468_y0;
  assign f_u_cla12_and469_f_u_cla12_and467_y0 = f_u_cla12_and467_y0;
  assign f_u_cla12_and469_y0 = f_u_cla12_and469_f_u_cla12_and468_y0 & f_u_cla12_and469_f_u_cla12_and467_y0;
  assign f_u_cla12_and470_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and470_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and470_y0 = f_u_cla12_and470_f_u_cla12_pg_logic5_y0 & f_u_cla12_and470_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and471_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and471_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and471_y0 = f_u_cla12_and471_f_u_cla12_pg_logic6_y0 & f_u_cla12_and471_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and472_f_u_cla12_and471_y0 = f_u_cla12_and471_y0;
  assign f_u_cla12_and472_f_u_cla12_and470_y0 = f_u_cla12_and470_y0;
  assign f_u_cla12_and472_y0 = f_u_cla12_and472_f_u_cla12_and471_y0 & f_u_cla12_and472_f_u_cla12_and470_y0;
  assign f_u_cla12_and473_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and473_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and473_y0 = f_u_cla12_and473_f_u_cla12_pg_logic7_y0 & f_u_cla12_and473_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and474_f_u_cla12_and473_y0 = f_u_cla12_and473_y0;
  assign f_u_cla12_and474_f_u_cla12_and472_y0 = f_u_cla12_and472_y0;
  assign f_u_cla12_and474_y0 = f_u_cla12_and474_f_u_cla12_and473_y0 & f_u_cla12_and474_f_u_cla12_and472_y0;
  assign f_u_cla12_and475_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and475_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and475_y0 = f_u_cla12_and475_f_u_cla12_pg_logic8_y0 & f_u_cla12_and475_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and476_f_u_cla12_and475_y0 = f_u_cla12_and475_y0;
  assign f_u_cla12_and476_f_u_cla12_and474_y0 = f_u_cla12_and474_y0;
  assign f_u_cla12_and476_y0 = f_u_cla12_and476_f_u_cla12_and475_y0 & f_u_cla12_and476_f_u_cla12_and474_y0;
  assign f_u_cla12_and477_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and477_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and477_y0 = f_u_cla12_and477_f_u_cla12_pg_logic9_y0 & f_u_cla12_and477_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and478_f_u_cla12_and477_y0 = f_u_cla12_and477_y0;
  assign f_u_cla12_and478_f_u_cla12_and476_y0 = f_u_cla12_and476_y0;
  assign f_u_cla12_and478_y0 = f_u_cla12_and478_f_u_cla12_and477_y0 & f_u_cla12_and478_f_u_cla12_and476_y0;
  assign f_u_cla12_and479_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and479_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and479_y0 = f_u_cla12_and479_f_u_cla12_pg_logic10_y0 & f_u_cla12_and479_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and480_f_u_cla12_and479_y0 = f_u_cla12_and479_y0;
  assign f_u_cla12_and480_f_u_cla12_and478_y0 = f_u_cla12_and478_y0;
  assign f_u_cla12_and480_y0 = f_u_cla12_and480_f_u_cla12_and479_y0 & f_u_cla12_and480_f_u_cla12_and478_y0;
  assign f_u_cla12_and481_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and481_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and481_y0 = f_u_cla12_and481_f_u_cla12_pg_logic6_y0 & f_u_cla12_and481_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and482_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and482_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and482_y0 = f_u_cla12_and482_f_u_cla12_pg_logic7_y0 & f_u_cla12_and482_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and483_f_u_cla12_and482_y0 = f_u_cla12_and482_y0;
  assign f_u_cla12_and483_f_u_cla12_and481_y0 = f_u_cla12_and481_y0;
  assign f_u_cla12_and483_y0 = f_u_cla12_and483_f_u_cla12_and482_y0 & f_u_cla12_and483_f_u_cla12_and481_y0;
  assign f_u_cla12_and484_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and484_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and484_y0 = f_u_cla12_and484_f_u_cla12_pg_logic8_y0 & f_u_cla12_and484_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and485_f_u_cla12_and484_y0 = f_u_cla12_and484_y0;
  assign f_u_cla12_and485_f_u_cla12_and483_y0 = f_u_cla12_and483_y0;
  assign f_u_cla12_and485_y0 = f_u_cla12_and485_f_u_cla12_and484_y0 & f_u_cla12_and485_f_u_cla12_and483_y0;
  assign f_u_cla12_and486_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and486_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and486_y0 = f_u_cla12_and486_f_u_cla12_pg_logic9_y0 & f_u_cla12_and486_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and487_f_u_cla12_and486_y0 = f_u_cla12_and486_y0;
  assign f_u_cla12_and487_f_u_cla12_and485_y0 = f_u_cla12_and485_y0;
  assign f_u_cla12_and487_y0 = f_u_cla12_and487_f_u_cla12_and486_y0 & f_u_cla12_and487_f_u_cla12_and485_y0;
  assign f_u_cla12_and488_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and488_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and488_y0 = f_u_cla12_and488_f_u_cla12_pg_logic10_y0 & f_u_cla12_and488_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and489_f_u_cla12_and488_y0 = f_u_cla12_and488_y0;
  assign f_u_cla12_and489_f_u_cla12_and487_y0 = f_u_cla12_and487_y0;
  assign f_u_cla12_and489_y0 = f_u_cla12_and489_f_u_cla12_and488_y0 & f_u_cla12_and489_f_u_cla12_and487_y0;
  assign f_u_cla12_and490_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and490_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and490_y0 = f_u_cla12_and490_f_u_cla12_pg_logic7_y0 & f_u_cla12_and490_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and491_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and491_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and491_y0 = f_u_cla12_and491_f_u_cla12_pg_logic8_y0 & f_u_cla12_and491_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and492_f_u_cla12_and491_y0 = f_u_cla12_and491_y0;
  assign f_u_cla12_and492_f_u_cla12_and490_y0 = f_u_cla12_and490_y0;
  assign f_u_cla12_and492_y0 = f_u_cla12_and492_f_u_cla12_and491_y0 & f_u_cla12_and492_f_u_cla12_and490_y0;
  assign f_u_cla12_and493_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and493_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and493_y0 = f_u_cla12_and493_f_u_cla12_pg_logic9_y0 & f_u_cla12_and493_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and494_f_u_cla12_and493_y0 = f_u_cla12_and493_y0;
  assign f_u_cla12_and494_f_u_cla12_and492_y0 = f_u_cla12_and492_y0;
  assign f_u_cla12_and494_y0 = f_u_cla12_and494_f_u_cla12_and493_y0 & f_u_cla12_and494_f_u_cla12_and492_y0;
  assign f_u_cla12_and495_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and495_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and495_y0 = f_u_cla12_and495_f_u_cla12_pg_logic10_y0 & f_u_cla12_and495_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and496_f_u_cla12_and495_y0 = f_u_cla12_and495_y0;
  assign f_u_cla12_and496_f_u_cla12_and494_y0 = f_u_cla12_and494_y0;
  assign f_u_cla12_and496_y0 = f_u_cla12_and496_f_u_cla12_and495_y0 & f_u_cla12_and496_f_u_cla12_and494_y0;
  assign f_u_cla12_and497_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and497_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and497_y0 = f_u_cla12_and497_f_u_cla12_pg_logic8_y0 & f_u_cla12_and497_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and498_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and498_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and498_y0 = f_u_cla12_and498_f_u_cla12_pg_logic9_y0 & f_u_cla12_and498_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and499_f_u_cla12_and498_y0 = f_u_cla12_and498_y0;
  assign f_u_cla12_and499_f_u_cla12_and497_y0 = f_u_cla12_and497_y0;
  assign f_u_cla12_and499_y0 = f_u_cla12_and499_f_u_cla12_and498_y0 & f_u_cla12_and499_f_u_cla12_and497_y0;
  assign f_u_cla12_and500_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and500_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and500_y0 = f_u_cla12_and500_f_u_cla12_pg_logic10_y0 & f_u_cla12_and500_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and501_f_u_cla12_and500_y0 = f_u_cla12_and500_y0;
  assign f_u_cla12_and501_f_u_cla12_and499_y0 = f_u_cla12_and499_y0;
  assign f_u_cla12_and501_y0 = f_u_cla12_and501_f_u_cla12_and500_y0 & f_u_cla12_and501_f_u_cla12_and499_y0;
  assign f_u_cla12_and502_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and502_f_u_cla12_pg_logic8_y1 = f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and502_y0 = f_u_cla12_and502_f_u_cla12_pg_logic9_y0 & f_u_cla12_and502_f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and503_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and503_f_u_cla12_pg_logic8_y1 = f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and503_y0 = f_u_cla12_and503_f_u_cla12_pg_logic10_y0 & f_u_cla12_and503_f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and504_f_u_cla12_and503_y0 = f_u_cla12_and503_y0;
  assign f_u_cla12_and504_f_u_cla12_and502_y0 = f_u_cla12_and502_y0;
  assign f_u_cla12_and504_y0 = f_u_cla12_and504_f_u_cla12_and503_y0 & f_u_cla12_and504_f_u_cla12_and502_y0;
  assign f_u_cla12_and505_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and505_f_u_cla12_pg_logic9_y1 = f_u_cla12_pg_logic9_y1;
  assign f_u_cla12_and505_y0 = f_u_cla12_and505_f_u_cla12_pg_logic10_y0 & f_u_cla12_and505_f_u_cla12_pg_logic9_y1;
  assign f_u_cla12_or55_f_u_cla12_and505_y0 = f_u_cla12_and505_y0;
  assign f_u_cla12_or55_f_u_cla12_and405_y0 = f_u_cla12_and405_y0;
  assign f_u_cla12_or55_y0 = f_u_cla12_or55_f_u_cla12_and505_y0 | f_u_cla12_or55_f_u_cla12_and405_y0;
  assign f_u_cla12_or56_f_u_cla12_or55_y0 = f_u_cla12_or55_y0;
  assign f_u_cla12_or56_f_u_cla12_and424_y0 = f_u_cla12_and424_y0;
  assign f_u_cla12_or56_y0 = f_u_cla12_or56_f_u_cla12_or55_y0 | f_u_cla12_or56_f_u_cla12_and424_y0;
  assign f_u_cla12_or57_f_u_cla12_or56_y0 = f_u_cla12_or56_y0;
  assign f_u_cla12_or57_f_u_cla12_and441_y0 = f_u_cla12_and441_y0;
  assign f_u_cla12_or57_y0 = f_u_cla12_or57_f_u_cla12_or56_y0 | f_u_cla12_or57_f_u_cla12_and441_y0;
  assign f_u_cla12_or58_f_u_cla12_or57_y0 = f_u_cla12_or57_y0;
  assign f_u_cla12_or58_f_u_cla12_and456_y0 = f_u_cla12_and456_y0;
  assign f_u_cla12_or58_y0 = f_u_cla12_or58_f_u_cla12_or57_y0 | f_u_cla12_or58_f_u_cla12_and456_y0;
  assign f_u_cla12_or59_f_u_cla12_or58_y0 = f_u_cla12_or58_y0;
  assign f_u_cla12_or59_f_u_cla12_and469_y0 = f_u_cla12_and469_y0;
  assign f_u_cla12_or59_y0 = f_u_cla12_or59_f_u_cla12_or58_y0 | f_u_cla12_or59_f_u_cla12_and469_y0;
  assign f_u_cla12_or60_f_u_cla12_or59_y0 = f_u_cla12_or59_y0;
  assign f_u_cla12_or60_f_u_cla12_and480_y0 = f_u_cla12_and480_y0;
  assign f_u_cla12_or60_y0 = f_u_cla12_or60_f_u_cla12_or59_y0 | f_u_cla12_or60_f_u_cla12_and480_y0;
  assign f_u_cla12_or61_f_u_cla12_or60_y0 = f_u_cla12_or60_y0;
  assign f_u_cla12_or61_f_u_cla12_and489_y0 = f_u_cla12_and489_y0;
  assign f_u_cla12_or61_y0 = f_u_cla12_or61_f_u_cla12_or60_y0 | f_u_cla12_or61_f_u_cla12_and489_y0;
  assign f_u_cla12_or62_f_u_cla12_or61_y0 = f_u_cla12_or61_y0;
  assign f_u_cla12_or62_f_u_cla12_and496_y0 = f_u_cla12_and496_y0;
  assign f_u_cla12_or62_y0 = f_u_cla12_or62_f_u_cla12_or61_y0 | f_u_cla12_or62_f_u_cla12_and496_y0;
  assign f_u_cla12_or63_f_u_cla12_or62_y0 = f_u_cla12_or62_y0;
  assign f_u_cla12_or63_f_u_cla12_and501_y0 = f_u_cla12_and501_y0;
  assign f_u_cla12_or63_y0 = f_u_cla12_or63_f_u_cla12_or62_y0 | f_u_cla12_or63_f_u_cla12_and501_y0;
  assign f_u_cla12_or64_f_u_cla12_or63_y0 = f_u_cla12_or63_y0;
  assign f_u_cla12_or64_f_u_cla12_and504_y0 = f_u_cla12_and504_y0;
  assign f_u_cla12_or64_y0 = f_u_cla12_or64_f_u_cla12_or63_y0 | f_u_cla12_or64_f_u_cla12_and504_y0;
  assign f_u_cla12_or65_f_u_cla12_pg_logic10_y1 = f_u_cla12_pg_logic10_y1;
  assign f_u_cla12_or65_f_u_cla12_or64_y0 = f_u_cla12_or64_y0;
  assign f_u_cla12_or65_y0 = f_u_cla12_or65_f_u_cla12_pg_logic10_y1 | f_u_cla12_or65_f_u_cla12_or64_y0;
  assign f_u_cla12_pg_logic11_a_11 = a_11;
  assign f_u_cla12_pg_logic11_b_11 = b_11;
  assign f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_a_11 | f_u_cla12_pg_logic11_b_11;
  assign f_u_cla12_pg_logic11_y1 = f_u_cla12_pg_logic11_a_11 & f_u_cla12_pg_logic11_b_11;
  assign f_u_cla12_pg_logic11_y2 = f_u_cla12_pg_logic11_a_11 ^ f_u_cla12_pg_logic11_b_11;
  assign f_u_cla12_xor11_f_u_cla12_pg_logic11_y2 = f_u_cla12_pg_logic11_y2;
  assign f_u_cla12_xor11_f_u_cla12_or65_y0 = f_u_cla12_or65_y0;
  assign f_u_cla12_xor11_y0 = f_u_cla12_xor11_f_u_cla12_pg_logic11_y2 ^ f_u_cla12_xor11_f_u_cla12_or65_y0;
  assign f_u_cla12_and506_f_u_cla12_pg_logic0_y0 = f_u_cla12_pg_logic0_y0;
  assign f_u_cla12_and506_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and506_y0 = f_u_cla12_and506_f_u_cla12_pg_logic0_y0 & f_u_cla12_and506_constant_wire_0;
  assign f_u_cla12_and507_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and507_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and507_y0 = f_u_cla12_and507_f_u_cla12_pg_logic1_y0 & f_u_cla12_and507_constant_wire_0;
  assign f_u_cla12_and508_f_u_cla12_and507_y0 = f_u_cla12_and507_y0;
  assign f_u_cla12_and508_f_u_cla12_and506_y0 = f_u_cla12_and506_y0;
  assign f_u_cla12_and508_y0 = f_u_cla12_and508_f_u_cla12_and507_y0 & f_u_cla12_and508_f_u_cla12_and506_y0;
  assign f_u_cla12_and509_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and509_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and509_y0 = f_u_cla12_and509_f_u_cla12_pg_logic2_y0 & f_u_cla12_and509_constant_wire_0;
  assign f_u_cla12_and510_f_u_cla12_and509_y0 = f_u_cla12_and509_y0;
  assign f_u_cla12_and510_f_u_cla12_and508_y0 = f_u_cla12_and508_y0;
  assign f_u_cla12_and510_y0 = f_u_cla12_and510_f_u_cla12_and509_y0 & f_u_cla12_and510_f_u_cla12_and508_y0;
  assign f_u_cla12_and511_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and511_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and511_y0 = f_u_cla12_and511_f_u_cla12_pg_logic3_y0 & f_u_cla12_and511_constant_wire_0;
  assign f_u_cla12_and512_f_u_cla12_and511_y0 = f_u_cla12_and511_y0;
  assign f_u_cla12_and512_f_u_cla12_and510_y0 = f_u_cla12_and510_y0;
  assign f_u_cla12_and512_y0 = f_u_cla12_and512_f_u_cla12_and511_y0 & f_u_cla12_and512_f_u_cla12_and510_y0;
  assign f_u_cla12_and513_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and513_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and513_y0 = f_u_cla12_and513_f_u_cla12_pg_logic4_y0 & f_u_cla12_and513_constant_wire_0;
  assign f_u_cla12_and514_f_u_cla12_and513_y0 = f_u_cla12_and513_y0;
  assign f_u_cla12_and514_f_u_cla12_and512_y0 = f_u_cla12_and512_y0;
  assign f_u_cla12_and514_y0 = f_u_cla12_and514_f_u_cla12_and513_y0 & f_u_cla12_and514_f_u_cla12_and512_y0;
  assign f_u_cla12_and515_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and515_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and515_y0 = f_u_cla12_and515_f_u_cla12_pg_logic5_y0 & f_u_cla12_and515_constant_wire_0;
  assign f_u_cla12_and516_f_u_cla12_and515_y0 = f_u_cla12_and515_y0;
  assign f_u_cla12_and516_f_u_cla12_and514_y0 = f_u_cla12_and514_y0;
  assign f_u_cla12_and516_y0 = f_u_cla12_and516_f_u_cla12_and515_y0 & f_u_cla12_and516_f_u_cla12_and514_y0;
  assign f_u_cla12_and517_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and517_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and517_y0 = f_u_cla12_and517_f_u_cla12_pg_logic6_y0 & f_u_cla12_and517_constant_wire_0;
  assign f_u_cla12_and518_f_u_cla12_and517_y0 = f_u_cla12_and517_y0;
  assign f_u_cla12_and518_f_u_cla12_and516_y0 = f_u_cla12_and516_y0;
  assign f_u_cla12_and518_y0 = f_u_cla12_and518_f_u_cla12_and517_y0 & f_u_cla12_and518_f_u_cla12_and516_y0;
  assign f_u_cla12_and519_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and519_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and519_y0 = f_u_cla12_and519_f_u_cla12_pg_logic7_y0 & f_u_cla12_and519_constant_wire_0;
  assign f_u_cla12_and520_f_u_cla12_and519_y0 = f_u_cla12_and519_y0;
  assign f_u_cla12_and520_f_u_cla12_and518_y0 = f_u_cla12_and518_y0;
  assign f_u_cla12_and520_y0 = f_u_cla12_and520_f_u_cla12_and519_y0 & f_u_cla12_and520_f_u_cla12_and518_y0;
  assign f_u_cla12_and521_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and521_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and521_y0 = f_u_cla12_and521_f_u_cla12_pg_logic8_y0 & f_u_cla12_and521_constant_wire_0;
  assign f_u_cla12_and522_f_u_cla12_and521_y0 = f_u_cla12_and521_y0;
  assign f_u_cla12_and522_f_u_cla12_and520_y0 = f_u_cla12_and520_y0;
  assign f_u_cla12_and522_y0 = f_u_cla12_and522_f_u_cla12_and521_y0 & f_u_cla12_and522_f_u_cla12_and520_y0;
  assign f_u_cla12_and523_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and523_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and523_y0 = f_u_cla12_and523_f_u_cla12_pg_logic9_y0 & f_u_cla12_and523_constant_wire_0;
  assign f_u_cla12_and524_f_u_cla12_and523_y0 = f_u_cla12_and523_y0;
  assign f_u_cla12_and524_f_u_cla12_and522_y0 = f_u_cla12_and522_y0;
  assign f_u_cla12_and524_y0 = f_u_cla12_and524_f_u_cla12_and523_y0 & f_u_cla12_and524_f_u_cla12_and522_y0;
  assign f_u_cla12_and525_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and525_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and525_y0 = f_u_cla12_and525_f_u_cla12_pg_logic10_y0 & f_u_cla12_and525_constant_wire_0;
  assign f_u_cla12_and526_f_u_cla12_and525_y0 = f_u_cla12_and525_y0;
  assign f_u_cla12_and526_f_u_cla12_and524_y0 = f_u_cla12_and524_y0;
  assign f_u_cla12_and526_y0 = f_u_cla12_and526_f_u_cla12_and525_y0 & f_u_cla12_and526_f_u_cla12_and524_y0;
  assign f_u_cla12_and527_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and527_constant_wire_0 = constant_wire_0;
  assign f_u_cla12_and527_y0 = f_u_cla12_and527_f_u_cla12_pg_logic11_y0 & f_u_cla12_and527_constant_wire_0;
  assign f_u_cla12_and528_f_u_cla12_and527_y0 = f_u_cla12_and527_y0;
  assign f_u_cla12_and528_f_u_cla12_and526_y0 = f_u_cla12_and526_y0;
  assign f_u_cla12_and528_y0 = f_u_cla12_and528_f_u_cla12_and527_y0 & f_u_cla12_and528_f_u_cla12_and526_y0;
  assign f_u_cla12_and529_f_u_cla12_pg_logic1_y0 = f_u_cla12_pg_logic1_y0;
  assign f_u_cla12_and529_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and529_y0 = f_u_cla12_and529_f_u_cla12_pg_logic1_y0 & f_u_cla12_and529_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and530_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and530_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and530_y0 = f_u_cla12_and530_f_u_cla12_pg_logic2_y0 & f_u_cla12_and530_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and531_f_u_cla12_and530_y0 = f_u_cla12_and530_y0;
  assign f_u_cla12_and531_f_u_cla12_and529_y0 = f_u_cla12_and529_y0;
  assign f_u_cla12_and531_y0 = f_u_cla12_and531_f_u_cla12_and530_y0 & f_u_cla12_and531_f_u_cla12_and529_y0;
  assign f_u_cla12_and532_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and532_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and532_y0 = f_u_cla12_and532_f_u_cla12_pg_logic3_y0 & f_u_cla12_and532_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and533_f_u_cla12_and532_y0 = f_u_cla12_and532_y0;
  assign f_u_cla12_and533_f_u_cla12_and531_y0 = f_u_cla12_and531_y0;
  assign f_u_cla12_and533_y0 = f_u_cla12_and533_f_u_cla12_and532_y0 & f_u_cla12_and533_f_u_cla12_and531_y0;
  assign f_u_cla12_and534_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and534_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and534_y0 = f_u_cla12_and534_f_u_cla12_pg_logic4_y0 & f_u_cla12_and534_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and535_f_u_cla12_and534_y0 = f_u_cla12_and534_y0;
  assign f_u_cla12_and535_f_u_cla12_and533_y0 = f_u_cla12_and533_y0;
  assign f_u_cla12_and535_y0 = f_u_cla12_and535_f_u_cla12_and534_y0 & f_u_cla12_and535_f_u_cla12_and533_y0;
  assign f_u_cla12_and536_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and536_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and536_y0 = f_u_cla12_and536_f_u_cla12_pg_logic5_y0 & f_u_cla12_and536_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and537_f_u_cla12_and536_y0 = f_u_cla12_and536_y0;
  assign f_u_cla12_and537_f_u_cla12_and535_y0 = f_u_cla12_and535_y0;
  assign f_u_cla12_and537_y0 = f_u_cla12_and537_f_u_cla12_and536_y0 & f_u_cla12_and537_f_u_cla12_and535_y0;
  assign f_u_cla12_and538_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and538_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and538_y0 = f_u_cla12_and538_f_u_cla12_pg_logic6_y0 & f_u_cla12_and538_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and539_f_u_cla12_and538_y0 = f_u_cla12_and538_y0;
  assign f_u_cla12_and539_f_u_cla12_and537_y0 = f_u_cla12_and537_y0;
  assign f_u_cla12_and539_y0 = f_u_cla12_and539_f_u_cla12_and538_y0 & f_u_cla12_and539_f_u_cla12_and537_y0;
  assign f_u_cla12_and540_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and540_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and540_y0 = f_u_cla12_and540_f_u_cla12_pg_logic7_y0 & f_u_cla12_and540_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and541_f_u_cla12_and540_y0 = f_u_cla12_and540_y0;
  assign f_u_cla12_and541_f_u_cla12_and539_y0 = f_u_cla12_and539_y0;
  assign f_u_cla12_and541_y0 = f_u_cla12_and541_f_u_cla12_and540_y0 & f_u_cla12_and541_f_u_cla12_and539_y0;
  assign f_u_cla12_and542_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and542_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and542_y0 = f_u_cla12_and542_f_u_cla12_pg_logic8_y0 & f_u_cla12_and542_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and543_f_u_cla12_and542_y0 = f_u_cla12_and542_y0;
  assign f_u_cla12_and543_f_u_cla12_and541_y0 = f_u_cla12_and541_y0;
  assign f_u_cla12_and543_y0 = f_u_cla12_and543_f_u_cla12_and542_y0 & f_u_cla12_and543_f_u_cla12_and541_y0;
  assign f_u_cla12_and544_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and544_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and544_y0 = f_u_cla12_and544_f_u_cla12_pg_logic9_y0 & f_u_cla12_and544_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and545_f_u_cla12_and544_y0 = f_u_cla12_and544_y0;
  assign f_u_cla12_and545_f_u_cla12_and543_y0 = f_u_cla12_and543_y0;
  assign f_u_cla12_and545_y0 = f_u_cla12_and545_f_u_cla12_and544_y0 & f_u_cla12_and545_f_u_cla12_and543_y0;
  assign f_u_cla12_and546_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and546_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and546_y0 = f_u_cla12_and546_f_u_cla12_pg_logic10_y0 & f_u_cla12_and546_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and547_f_u_cla12_and546_y0 = f_u_cla12_and546_y0;
  assign f_u_cla12_and547_f_u_cla12_and545_y0 = f_u_cla12_and545_y0;
  assign f_u_cla12_and547_y0 = f_u_cla12_and547_f_u_cla12_and546_y0 & f_u_cla12_and547_f_u_cla12_and545_y0;
  assign f_u_cla12_and548_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and548_f_u_cla12_pg_logic0_y1 = f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and548_y0 = f_u_cla12_and548_f_u_cla12_pg_logic11_y0 & f_u_cla12_and548_f_u_cla12_pg_logic0_y1;
  assign f_u_cla12_and549_f_u_cla12_and548_y0 = f_u_cla12_and548_y0;
  assign f_u_cla12_and549_f_u_cla12_and547_y0 = f_u_cla12_and547_y0;
  assign f_u_cla12_and549_y0 = f_u_cla12_and549_f_u_cla12_and548_y0 & f_u_cla12_and549_f_u_cla12_and547_y0;
  assign f_u_cla12_and550_f_u_cla12_pg_logic2_y0 = f_u_cla12_pg_logic2_y0;
  assign f_u_cla12_and550_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and550_y0 = f_u_cla12_and550_f_u_cla12_pg_logic2_y0 & f_u_cla12_and550_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and551_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and551_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and551_y0 = f_u_cla12_and551_f_u_cla12_pg_logic3_y0 & f_u_cla12_and551_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and552_f_u_cla12_and551_y0 = f_u_cla12_and551_y0;
  assign f_u_cla12_and552_f_u_cla12_and550_y0 = f_u_cla12_and550_y0;
  assign f_u_cla12_and552_y0 = f_u_cla12_and552_f_u_cla12_and551_y0 & f_u_cla12_and552_f_u_cla12_and550_y0;
  assign f_u_cla12_and553_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and553_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and553_y0 = f_u_cla12_and553_f_u_cla12_pg_logic4_y0 & f_u_cla12_and553_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and554_f_u_cla12_and553_y0 = f_u_cla12_and553_y0;
  assign f_u_cla12_and554_f_u_cla12_and552_y0 = f_u_cla12_and552_y0;
  assign f_u_cla12_and554_y0 = f_u_cla12_and554_f_u_cla12_and553_y0 & f_u_cla12_and554_f_u_cla12_and552_y0;
  assign f_u_cla12_and555_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and555_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and555_y0 = f_u_cla12_and555_f_u_cla12_pg_logic5_y0 & f_u_cla12_and555_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and556_f_u_cla12_and555_y0 = f_u_cla12_and555_y0;
  assign f_u_cla12_and556_f_u_cla12_and554_y0 = f_u_cla12_and554_y0;
  assign f_u_cla12_and556_y0 = f_u_cla12_and556_f_u_cla12_and555_y0 & f_u_cla12_and556_f_u_cla12_and554_y0;
  assign f_u_cla12_and557_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and557_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and557_y0 = f_u_cla12_and557_f_u_cla12_pg_logic6_y0 & f_u_cla12_and557_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and558_f_u_cla12_and557_y0 = f_u_cla12_and557_y0;
  assign f_u_cla12_and558_f_u_cla12_and556_y0 = f_u_cla12_and556_y0;
  assign f_u_cla12_and558_y0 = f_u_cla12_and558_f_u_cla12_and557_y0 & f_u_cla12_and558_f_u_cla12_and556_y0;
  assign f_u_cla12_and559_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and559_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and559_y0 = f_u_cla12_and559_f_u_cla12_pg_logic7_y0 & f_u_cla12_and559_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and560_f_u_cla12_and559_y0 = f_u_cla12_and559_y0;
  assign f_u_cla12_and560_f_u_cla12_and558_y0 = f_u_cla12_and558_y0;
  assign f_u_cla12_and560_y0 = f_u_cla12_and560_f_u_cla12_and559_y0 & f_u_cla12_and560_f_u_cla12_and558_y0;
  assign f_u_cla12_and561_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and561_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and561_y0 = f_u_cla12_and561_f_u_cla12_pg_logic8_y0 & f_u_cla12_and561_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and562_f_u_cla12_and561_y0 = f_u_cla12_and561_y0;
  assign f_u_cla12_and562_f_u_cla12_and560_y0 = f_u_cla12_and560_y0;
  assign f_u_cla12_and562_y0 = f_u_cla12_and562_f_u_cla12_and561_y0 & f_u_cla12_and562_f_u_cla12_and560_y0;
  assign f_u_cla12_and563_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and563_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and563_y0 = f_u_cla12_and563_f_u_cla12_pg_logic9_y0 & f_u_cla12_and563_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and564_f_u_cla12_and563_y0 = f_u_cla12_and563_y0;
  assign f_u_cla12_and564_f_u_cla12_and562_y0 = f_u_cla12_and562_y0;
  assign f_u_cla12_and564_y0 = f_u_cla12_and564_f_u_cla12_and563_y0 & f_u_cla12_and564_f_u_cla12_and562_y0;
  assign f_u_cla12_and565_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and565_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and565_y0 = f_u_cla12_and565_f_u_cla12_pg_logic10_y0 & f_u_cla12_and565_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and566_f_u_cla12_and565_y0 = f_u_cla12_and565_y0;
  assign f_u_cla12_and566_f_u_cla12_and564_y0 = f_u_cla12_and564_y0;
  assign f_u_cla12_and566_y0 = f_u_cla12_and566_f_u_cla12_and565_y0 & f_u_cla12_and566_f_u_cla12_and564_y0;
  assign f_u_cla12_and567_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and567_f_u_cla12_pg_logic1_y1 = f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and567_y0 = f_u_cla12_and567_f_u_cla12_pg_logic11_y0 & f_u_cla12_and567_f_u_cla12_pg_logic1_y1;
  assign f_u_cla12_and568_f_u_cla12_and567_y0 = f_u_cla12_and567_y0;
  assign f_u_cla12_and568_f_u_cla12_and566_y0 = f_u_cla12_and566_y0;
  assign f_u_cla12_and568_y0 = f_u_cla12_and568_f_u_cla12_and567_y0 & f_u_cla12_and568_f_u_cla12_and566_y0;
  assign f_u_cla12_and569_f_u_cla12_pg_logic3_y0 = f_u_cla12_pg_logic3_y0;
  assign f_u_cla12_and569_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and569_y0 = f_u_cla12_and569_f_u_cla12_pg_logic3_y0 & f_u_cla12_and569_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and570_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and570_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and570_y0 = f_u_cla12_and570_f_u_cla12_pg_logic4_y0 & f_u_cla12_and570_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and571_f_u_cla12_and570_y0 = f_u_cla12_and570_y0;
  assign f_u_cla12_and571_f_u_cla12_and569_y0 = f_u_cla12_and569_y0;
  assign f_u_cla12_and571_y0 = f_u_cla12_and571_f_u_cla12_and570_y0 & f_u_cla12_and571_f_u_cla12_and569_y0;
  assign f_u_cla12_and572_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and572_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and572_y0 = f_u_cla12_and572_f_u_cla12_pg_logic5_y0 & f_u_cla12_and572_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and573_f_u_cla12_and572_y0 = f_u_cla12_and572_y0;
  assign f_u_cla12_and573_f_u_cla12_and571_y0 = f_u_cla12_and571_y0;
  assign f_u_cla12_and573_y0 = f_u_cla12_and573_f_u_cla12_and572_y0 & f_u_cla12_and573_f_u_cla12_and571_y0;
  assign f_u_cla12_and574_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and574_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and574_y0 = f_u_cla12_and574_f_u_cla12_pg_logic6_y0 & f_u_cla12_and574_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and575_f_u_cla12_and574_y0 = f_u_cla12_and574_y0;
  assign f_u_cla12_and575_f_u_cla12_and573_y0 = f_u_cla12_and573_y0;
  assign f_u_cla12_and575_y0 = f_u_cla12_and575_f_u_cla12_and574_y0 & f_u_cla12_and575_f_u_cla12_and573_y0;
  assign f_u_cla12_and576_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and576_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and576_y0 = f_u_cla12_and576_f_u_cla12_pg_logic7_y0 & f_u_cla12_and576_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and577_f_u_cla12_and576_y0 = f_u_cla12_and576_y0;
  assign f_u_cla12_and577_f_u_cla12_and575_y0 = f_u_cla12_and575_y0;
  assign f_u_cla12_and577_y0 = f_u_cla12_and577_f_u_cla12_and576_y0 & f_u_cla12_and577_f_u_cla12_and575_y0;
  assign f_u_cla12_and578_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and578_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and578_y0 = f_u_cla12_and578_f_u_cla12_pg_logic8_y0 & f_u_cla12_and578_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and579_f_u_cla12_and578_y0 = f_u_cla12_and578_y0;
  assign f_u_cla12_and579_f_u_cla12_and577_y0 = f_u_cla12_and577_y0;
  assign f_u_cla12_and579_y0 = f_u_cla12_and579_f_u_cla12_and578_y0 & f_u_cla12_and579_f_u_cla12_and577_y0;
  assign f_u_cla12_and580_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and580_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and580_y0 = f_u_cla12_and580_f_u_cla12_pg_logic9_y0 & f_u_cla12_and580_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and581_f_u_cla12_and580_y0 = f_u_cla12_and580_y0;
  assign f_u_cla12_and581_f_u_cla12_and579_y0 = f_u_cla12_and579_y0;
  assign f_u_cla12_and581_y0 = f_u_cla12_and581_f_u_cla12_and580_y0 & f_u_cla12_and581_f_u_cla12_and579_y0;
  assign f_u_cla12_and582_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and582_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and582_y0 = f_u_cla12_and582_f_u_cla12_pg_logic10_y0 & f_u_cla12_and582_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and583_f_u_cla12_and582_y0 = f_u_cla12_and582_y0;
  assign f_u_cla12_and583_f_u_cla12_and581_y0 = f_u_cla12_and581_y0;
  assign f_u_cla12_and583_y0 = f_u_cla12_and583_f_u_cla12_and582_y0 & f_u_cla12_and583_f_u_cla12_and581_y0;
  assign f_u_cla12_and584_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and584_f_u_cla12_pg_logic2_y1 = f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and584_y0 = f_u_cla12_and584_f_u_cla12_pg_logic11_y0 & f_u_cla12_and584_f_u_cla12_pg_logic2_y1;
  assign f_u_cla12_and585_f_u_cla12_and584_y0 = f_u_cla12_and584_y0;
  assign f_u_cla12_and585_f_u_cla12_and583_y0 = f_u_cla12_and583_y0;
  assign f_u_cla12_and585_y0 = f_u_cla12_and585_f_u_cla12_and584_y0 & f_u_cla12_and585_f_u_cla12_and583_y0;
  assign f_u_cla12_and586_f_u_cla12_pg_logic4_y0 = f_u_cla12_pg_logic4_y0;
  assign f_u_cla12_and586_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and586_y0 = f_u_cla12_and586_f_u_cla12_pg_logic4_y0 & f_u_cla12_and586_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and587_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and587_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and587_y0 = f_u_cla12_and587_f_u_cla12_pg_logic5_y0 & f_u_cla12_and587_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and588_f_u_cla12_and587_y0 = f_u_cla12_and587_y0;
  assign f_u_cla12_and588_f_u_cla12_and586_y0 = f_u_cla12_and586_y0;
  assign f_u_cla12_and588_y0 = f_u_cla12_and588_f_u_cla12_and587_y0 & f_u_cla12_and588_f_u_cla12_and586_y0;
  assign f_u_cla12_and589_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and589_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and589_y0 = f_u_cla12_and589_f_u_cla12_pg_logic6_y0 & f_u_cla12_and589_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and590_f_u_cla12_and589_y0 = f_u_cla12_and589_y0;
  assign f_u_cla12_and590_f_u_cla12_and588_y0 = f_u_cla12_and588_y0;
  assign f_u_cla12_and590_y0 = f_u_cla12_and590_f_u_cla12_and589_y0 & f_u_cla12_and590_f_u_cla12_and588_y0;
  assign f_u_cla12_and591_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and591_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and591_y0 = f_u_cla12_and591_f_u_cla12_pg_logic7_y0 & f_u_cla12_and591_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and592_f_u_cla12_and591_y0 = f_u_cla12_and591_y0;
  assign f_u_cla12_and592_f_u_cla12_and590_y0 = f_u_cla12_and590_y0;
  assign f_u_cla12_and592_y0 = f_u_cla12_and592_f_u_cla12_and591_y0 & f_u_cla12_and592_f_u_cla12_and590_y0;
  assign f_u_cla12_and593_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and593_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and593_y0 = f_u_cla12_and593_f_u_cla12_pg_logic8_y0 & f_u_cla12_and593_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and594_f_u_cla12_and593_y0 = f_u_cla12_and593_y0;
  assign f_u_cla12_and594_f_u_cla12_and592_y0 = f_u_cla12_and592_y0;
  assign f_u_cla12_and594_y0 = f_u_cla12_and594_f_u_cla12_and593_y0 & f_u_cla12_and594_f_u_cla12_and592_y0;
  assign f_u_cla12_and595_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and595_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and595_y0 = f_u_cla12_and595_f_u_cla12_pg_logic9_y0 & f_u_cla12_and595_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and596_f_u_cla12_and595_y0 = f_u_cla12_and595_y0;
  assign f_u_cla12_and596_f_u_cla12_and594_y0 = f_u_cla12_and594_y0;
  assign f_u_cla12_and596_y0 = f_u_cla12_and596_f_u_cla12_and595_y0 & f_u_cla12_and596_f_u_cla12_and594_y0;
  assign f_u_cla12_and597_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and597_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and597_y0 = f_u_cla12_and597_f_u_cla12_pg_logic10_y0 & f_u_cla12_and597_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and598_f_u_cla12_and597_y0 = f_u_cla12_and597_y0;
  assign f_u_cla12_and598_f_u_cla12_and596_y0 = f_u_cla12_and596_y0;
  assign f_u_cla12_and598_y0 = f_u_cla12_and598_f_u_cla12_and597_y0 & f_u_cla12_and598_f_u_cla12_and596_y0;
  assign f_u_cla12_and599_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and599_f_u_cla12_pg_logic3_y1 = f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and599_y0 = f_u_cla12_and599_f_u_cla12_pg_logic11_y0 & f_u_cla12_and599_f_u_cla12_pg_logic3_y1;
  assign f_u_cla12_and600_f_u_cla12_and599_y0 = f_u_cla12_and599_y0;
  assign f_u_cla12_and600_f_u_cla12_and598_y0 = f_u_cla12_and598_y0;
  assign f_u_cla12_and600_y0 = f_u_cla12_and600_f_u_cla12_and599_y0 & f_u_cla12_and600_f_u_cla12_and598_y0;
  assign f_u_cla12_and601_f_u_cla12_pg_logic5_y0 = f_u_cla12_pg_logic5_y0;
  assign f_u_cla12_and601_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and601_y0 = f_u_cla12_and601_f_u_cla12_pg_logic5_y0 & f_u_cla12_and601_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and602_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and602_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and602_y0 = f_u_cla12_and602_f_u_cla12_pg_logic6_y0 & f_u_cla12_and602_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and603_f_u_cla12_and602_y0 = f_u_cla12_and602_y0;
  assign f_u_cla12_and603_f_u_cla12_and601_y0 = f_u_cla12_and601_y0;
  assign f_u_cla12_and603_y0 = f_u_cla12_and603_f_u_cla12_and602_y0 & f_u_cla12_and603_f_u_cla12_and601_y0;
  assign f_u_cla12_and604_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and604_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and604_y0 = f_u_cla12_and604_f_u_cla12_pg_logic7_y0 & f_u_cla12_and604_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and605_f_u_cla12_and604_y0 = f_u_cla12_and604_y0;
  assign f_u_cla12_and605_f_u_cla12_and603_y0 = f_u_cla12_and603_y0;
  assign f_u_cla12_and605_y0 = f_u_cla12_and605_f_u_cla12_and604_y0 & f_u_cla12_and605_f_u_cla12_and603_y0;
  assign f_u_cla12_and606_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and606_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and606_y0 = f_u_cla12_and606_f_u_cla12_pg_logic8_y0 & f_u_cla12_and606_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and607_f_u_cla12_and606_y0 = f_u_cla12_and606_y0;
  assign f_u_cla12_and607_f_u_cla12_and605_y0 = f_u_cla12_and605_y0;
  assign f_u_cla12_and607_y0 = f_u_cla12_and607_f_u_cla12_and606_y0 & f_u_cla12_and607_f_u_cla12_and605_y0;
  assign f_u_cla12_and608_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and608_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and608_y0 = f_u_cla12_and608_f_u_cla12_pg_logic9_y0 & f_u_cla12_and608_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and609_f_u_cla12_and608_y0 = f_u_cla12_and608_y0;
  assign f_u_cla12_and609_f_u_cla12_and607_y0 = f_u_cla12_and607_y0;
  assign f_u_cla12_and609_y0 = f_u_cla12_and609_f_u_cla12_and608_y0 & f_u_cla12_and609_f_u_cla12_and607_y0;
  assign f_u_cla12_and610_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and610_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and610_y0 = f_u_cla12_and610_f_u_cla12_pg_logic10_y0 & f_u_cla12_and610_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and611_f_u_cla12_and610_y0 = f_u_cla12_and610_y0;
  assign f_u_cla12_and611_f_u_cla12_and609_y0 = f_u_cla12_and609_y0;
  assign f_u_cla12_and611_y0 = f_u_cla12_and611_f_u_cla12_and610_y0 & f_u_cla12_and611_f_u_cla12_and609_y0;
  assign f_u_cla12_and612_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and612_f_u_cla12_pg_logic4_y1 = f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and612_y0 = f_u_cla12_and612_f_u_cla12_pg_logic11_y0 & f_u_cla12_and612_f_u_cla12_pg_logic4_y1;
  assign f_u_cla12_and613_f_u_cla12_and612_y0 = f_u_cla12_and612_y0;
  assign f_u_cla12_and613_f_u_cla12_and611_y0 = f_u_cla12_and611_y0;
  assign f_u_cla12_and613_y0 = f_u_cla12_and613_f_u_cla12_and612_y0 & f_u_cla12_and613_f_u_cla12_and611_y0;
  assign f_u_cla12_and614_f_u_cla12_pg_logic6_y0 = f_u_cla12_pg_logic6_y0;
  assign f_u_cla12_and614_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and614_y0 = f_u_cla12_and614_f_u_cla12_pg_logic6_y0 & f_u_cla12_and614_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and615_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and615_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and615_y0 = f_u_cla12_and615_f_u_cla12_pg_logic7_y0 & f_u_cla12_and615_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and616_f_u_cla12_and615_y0 = f_u_cla12_and615_y0;
  assign f_u_cla12_and616_f_u_cla12_and614_y0 = f_u_cla12_and614_y0;
  assign f_u_cla12_and616_y0 = f_u_cla12_and616_f_u_cla12_and615_y0 & f_u_cla12_and616_f_u_cla12_and614_y0;
  assign f_u_cla12_and617_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and617_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and617_y0 = f_u_cla12_and617_f_u_cla12_pg_logic8_y0 & f_u_cla12_and617_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and618_f_u_cla12_and617_y0 = f_u_cla12_and617_y0;
  assign f_u_cla12_and618_f_u_cla12_and616_y0 = f_u_cla12_and616_y0;
  assign f_u_cla12_and618_y0 = f_u_cla12_and618_f_u_cla12_and617_y0 & f_u_cla12_and618_f_u_cla12_and616_y0;
  assign f_u_cla12_and619_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and619_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and619_y0 = f_u_cla12_and619_f_u_cla12_pg_logic9_y0 & f_u_cla12_and619_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and620_f_u_cla12_and619_y0 = f_u_cla12_and619_y0;
  assign f_u_cla12_and620_f_u_cla12_and618_y0 = f_u_cla12_and618_y0;
  assign f_u_cla12_and620_y0 = f_u_cla12_and620_f_u_cla12_and619_y0 & f_u_cla12_and620_f_u_cla12_and618_y0;
  assign f_u_cla12_and621_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and621_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and621_y0 = f_u_cla12_and621_f_u_cla12_pg_logic10_y0 & f_u_cla12_and621_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and622_f_u_cla12_and621_y0 = f_u_cla12_and621_y0;
  assign f_u_cla12_and622_f_u_cla12_and620_y0 = f_u_cla12_and620_y0;
  assign f_u_cla12_and622_y0 = f_u_cla12_and622_f_u_cla12_and621_y0 & f_u_cla12_and622_f_u_cla12_and620_y0;
  assign f_u_cla12_and623_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and623_f_u_cla12_pg_logic5_y1 = f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and623_y0 = f_u_cla12_and623_f_u_cla12_pg_logic11_y0 & f_u_cla12_and623_f_u_cla12_pg_logic5_y1;
  assign f_u_cla12_and624_f_u_cla12_and623_y0 = f_u_cla12_and623_y0;
  assign f_u_cla12_and624_f_u_cla12_and622_y0 = f_u_cla12_and622_y0;
  assign f_u_cla12_and624_y0 = f_u_cla12_and624_f_u_cla12_and623_y0 & f_u_cla12_and624_f_u_cla12_and622_y0;
  assign f_u_cla12_and625_f_u_cla12_pg_logic7_y0 = f_u_cla12_pg_logic7_y0;
  assign f_u_cla12_and625_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and625_y0 = f_u_cla12_and625_f_u_cla12_pg_logic7_y0 & f_u_cla12_and625_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and626_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and626_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and626_y0 = f_u_cla12_and626_f_u_cla12_pg_logic8_y0 & f_u_cla12_and626_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and627_f_u_cla12_and626_y0 = f_u_cla12_and626_y0;
  assign f_u_cla12_and627_f_u_cla12_and625_y0 = f_u_cla12_and625_y0;
  assign f_u_cla12_and627_y0 = f_u_cla12_and627_f_u_cla12_and626_y0 & f_u_cla12_and627_f_u_cla12_and625_y0;
  assign f_u_cla12_and628_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and628_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and628_y0 = f_u_cla12_and628_f_u_cla12_pg_logic9_y0 & f_u_cla12_and628_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and629_f_u_cla12_and628_y0 = f_u_cla12_and628_y0;
  assign f_u_cla12_and629_f_u_cla12_and627_y0 = f_u_cla12_and627_y0;
  assign f_u_cla12_and629_y0 = f_u_cla12_and629_f_u_cla12_and628_y0 & f_u_cla12_and629_f_u_cla12_and627_y0;
  assign f_u_cla12_and630_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and630_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and630_y0 = f_u_cla12_and630_f_u_cla12_pg_logic10_y0 & f_u_cla12_and630_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and631_f_u_cla12_and630_y0 = f_u_cla12_and630_y0;
  assign f_u_cla12_and631_f_u_cla12_and629_y0 = f_u_cla12_and629_y0;
  assign f_u_cla12_and631_y0 = f_u_cla12_and631_f_u_cla12_and630_y0 & f_u_cla12_and631_f_u_cla12_and629_y0;
  assign f_u_cla12_and632_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and632_f_u_cla12_pg_logic6_y1 = f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and632_y0 = f_u_cla12_and632_f_u_cla12_pg_logic11_y0 & f_u_cla12_and632_f_u_cla12_pg_logic6_y1;
  assign f_u_cla12_and633_f_u_cla12_and632_y0 = f_u_cla12_and632_y0;
  assign f_u_cla12_and633_f_u_cla12_and631_y0 = f_u_cla12_and631_y0;
  assign f_u_cla12_and633_y0 = f_u_cla12_and633_f_u_cla12_and632_y0 & f_u_cla12_and633_f_u_cla12_and631_y0;
  assign f_u_cla12_and634_f_u_cla12_pg_logic8_y0 = f_u_cla12_pg_logic8_y0;
  assign f_u_cla12_and634_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and634_y0 = f_u_cla12_and634_f_u_cla12_pg_logic8_y0 & f_u_cla12_and634_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and635_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and635_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and635_y0 = f_u_cla12_and635_f_u_cla12_pg_logic9_y0 & f_u_cla12_and635_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and636_f_u_cla12_and635_y0 = f_u_cla12_and635_y0;
  assign f_u_cla12_and636_f_u_cla12_and634_y0 = f_u_cla12_and634_y0;
  assign f_u_cla12_and636_y0 = f_u_cla12_and636_f_u_cla12_and635_y0 & f_u_cla12_and636_f_u_cla12_and634_y0;
  assign f_u_cla12_and637_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and637_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and637_y0 = f_u_cla12_and637_f_u_cla12_pg_logic10_y0 & f_u_cla12_and637_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and638_f_u_cla12_and637_y0 = f_u_cla12_and637_y0;
  assign f_u_cla12_and638_f_u_cla12_and636_y0 = f_u_cla12_and636_y0;
  assign f_u_cla12_and638_y0 = f_u_cla12_and638_f_u_cla12_and637_y0 & f_u_cla12_and638_f_u_cla12_and636_y0;
  assign f_u_cla12_and639_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and639_f_u_cla12_pg_logic7_y1 = f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and639_y0 = f_u_cla12_and639_f_u_cla12_pg_logic11_y0 & f_u_cla12_and639_f_u_cla12_pg_logic7_y1;
  assign f_u_cla12_and640_f_u_cla12_and639_y0 = f_u_cla12_and639_y0;
  assign f_u_cla12_and640_f_u_cla12_and638_y0 = f_u_cla12_and638_y0;
  assign f_u_cla12_and640_y0 = f_u_cla12_and640_f_u_cla12_and639_y0 & f_u_cla12_and640_f_u_cla12_and638_y0;
  assign f_u_cla12_and641_f_u_cla12_pg_logic9_y0 = f_u_cla12_pg_logic9_y0;
  assign f_u_cla12_and641_f_u_cla12_pg_logic8_y1 = f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and641_y0 = f_u_cla12_and641_f_u_cla12_pg_logic9_y0 & f_u_cla12_and641_f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and642_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and642_f_u_cla12_pg_logic8_y1 = f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and642_y0 = f_u_cla12_and642_f_u_cla12_pg_logic10_y0 & f_u_cla12_and642_f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and643_f_u_cla12_and642_y0 = f_u_cla12_and642_y0;
  assign f_u_cla12_and643_f_u_cla12_and641_y0 = f_u_cla12_and641_y0;
  assign f_u_cla12_and643_y0 = f_u_cla12_and643_f_u_cla12_and642_y0 & f_u_cla12_and643_f_u_cla12_and641_y0;
  assign f_u_cla12_and644_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and644_f_u_cla12_pg_logic8_y1 = f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and644_y0 = f_u_cla12_and644_f_u_cla12_pg_logic11_y0 & f_u_cla12_and644_f_u_cla12_pg_logic8_y1;
  assign f_u_cla12_and645_f_u_cla12_and644_y0 = f_u_cla12_and644_y0;
  assign f_u_cla12_and645_f_u_cla12_and643_y0 = f_u_cla12_and643_y0;
  assign f_u_cla12_and645_y0 = f_u_cla12_and645_f_u_cla12_and644_y0 & f_u_cla12_and645_f_u_cla12_and643_y0;
  assign f_u_cla12_and646_f_u_cla12_pg_logic10_y0 = f_u_cla12_pg_logic10_y0;
  assign f_u_cla12_and646_f_u_cla12_pg_logic9_y1 = f_u_cla12_pg_logic9_y1;
  assign f_u_cla12_and646_y0 = f_u_cla12_and646_f_u_cla12_pg_logic10_y0 & f_u_cla12_and646_f_u_cla12_pg_logic9_y1;
  assign f_u_cla12_and647_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and647_f_u_cla12_pg_logic9_y1 = f_u_cla12_pg_logic9_y1;
  assign f_u_cla12_and647_y0 = f_u_cla12_and647_f_u_cla12_pg_logic11_y0 & f_u_cla12_and647_f_u_cla12_pg_logic9_y1;
  assign f_u_cla12_and648_f_u_cla12_and647_y0 = f_u_cla12_and647_y0;
  assign f_u_cla12_and648_f_u_cla12_and646_y0 = f_u_cla12_and646_y0;
  assign f_u_cla12_and648_y0 = f_u_cla12_and648_f_u_cla12_and647_y0 & f_u_cla12_and648_f_u_cla12_and646_y0;
  assign f_u_cla12_and649_f_u_cla12_pg_logic11_y0 = f_u_cla12_pg_logic11_y0;
  assign f_u_cla12_and649_f_u_cla12_pg_logic10_y1 = f_u_cla12_pg_logic10_y1;
  assign f_u_cla12_and649_y0 = f_u_cla12_and649_f_u_cla12_pg_logic11_y0 & f_u_cla12_and649_f_u_cla12_pg_logic10_y1;
  assign f_u_cla12_or66_f_u_cla12_and649_y0 = f_u_cla12_and649_y0;
  assign f_u_cla12_or66_f_u_cla12_and528_y0 = f_u_cla12_and528_y0;
  assign f_u_cla12_or66_y0 = f_u_cla12_or66_f_u_cla12_and649_y0 | f_u_cla12_or66_f_u_cla12_and528_y0;
  assign f_u_cla12_or67_f_u_cla12_or66_y0 = f_u_cla12_or66_y0;
  assign f_u_cla12_or67_f_u_cla12_and549_y0 = f_u_cla12_and549_y0;
  assign f_u_cla12_or67_y0 = f_u_cla12_or67_f_u_cla12_or66_y0 | f_u_cla12_or67_f_u_cla12_and549_y0;
  assign f_u_cla12_or68_f_u_cla12_or67_y0 = f_u_cla12_or67_y0;
  assign f_u_cla12_or68_f_u_cla12_and568_y0 = f_u_cla12_and568_y0;
  assign f_u_cla12_or68_y0 = f_u_cla12_or68_f_u_cla12_or67_y0 | f_u_cla12_or68_f_u_cla12_and568_y0;
  assign f_u_cla12_or69_f_u_cla12_or68_y0 = f_u_cla12_or68_y0;
  assign f_u_cla12_or69_f_u_cla12_and585_y0 = f_u_cla12_and585_y0;
  assign f_u_cla12_or69_y0 = f_u_cla12_or69_f_u_cla12_or68_y0 | f_u_cla12_or69_f_u_cla12_and585_y0;
  assign f_u_cla12_or70_f_u_cla12_or69_y0 = f_u_cla12_or69_y0;
  assign f_u_cla12_or70_f_u_cla12_and600_y0 = f_u_cla12_and600_y0;
  assign f_u_cla12_or70_y0 = f_u_cla12_or70_f_u_cla12_or69_y0 | f_u_cla12_or70_f_u_cla12_and600_y0;
  assign f_u_cla12_or71_f_u_cla12_or70_y0 = f_u_cla12_or70_y0;
  assign f_u_cla12_or71_f_u_cla12_and613_y0 = f_u_cla12_and613_y0;
  assign f_u_cla12_or71_y0 = f_u_cla12_or71_f_u_cla12_or70_y0 | f_u_cla12_or71_f_u_cla12_and613_y0;
  assign f_u_cla12_or72_f_u_cla12_or71_y0 = f_u_cla12_or71_y0;
  assign f_u_cla12_or72_f_u_cla12_and624_y0 = f_u_cla12_and624_y0;
  assign f_u_cla12_or72_y0 = f_u_cla12_or72_f_u_cla12_or71_y0 | f_u_cla12_or72_f_u_cla12_and624_y0;
  assign f_u_cla12_or73_f_u_cla12_or72_y0 = f_u_cla12_or72_y0;
  assign f_u_cla12_or73_f_u_cla12_and633_y0 = f_u_cla12_and633_y0;
  assign f_u_cla12_or73_y0 = f_u_cla12_or73_f_u_cla12_or72_y0 | f_u_cla12_or73_f_u_cla12_and633_y0;
  assign f_u_cla12_or74_f_u_cla12_or73_y0 = f_u_cla12_or73_y0;
  assign f_u_cla12_or74_f_u_cla12_and640_y0 = f_u_cla12_and640_y0;
  assign f_u_cla12_or74_y0 = f_u_cla12_or74_f_u_cla12_or73_y0 | f_u_cla12_or74_f_u_cla12_and640_y0;
  assign f_u_cla12_or75_f_u_cla12_or74_y0 = f_u_cla12_or74_y0;
  assign f_u_cla12_or75_f_u_cla12_and645_y0 = f_u_cla12_and645_y0;
  assign f_u_cla12_or75_y0 = f_u_cla12_or75_f_u_cla12_or74_y0 | f_u_cla12_or75_f_u_cla12_and645_y0;
  assign f_u_cla12_or76_f_u_cla12_or75_y0 = f_u_cla12_or75_y0;
  assign f_u_cla12_or76_f_u_cla12_and648_y0 = f_u_cla12_and648_y0;
  assign f_u_cla12_or76_y0 = f_u_cla12_or76_f_u_cla12_or75_y0 | f_u_cla12_or76_f_u_cla12_and648_y0;
  assign f_u_cla12_or77_f_u_cla12_pg_logic11_y1 = f_u_cla12_pg_logic11_y1;
  assign f_u_cla12_or77_f_u_cla12_or76_y0 = f_u_cla12_or76_y0;
  assign f_u_cla12_or77_y0 = f_u_cla12_or77_f_u_cla12_pg_logic11_y1 | f_u_cla12_or77_f_u_cla12_or76_y0;

  assign out[0] = f_u_cla12_xor0_y0;
  assign out[1] = f_u_cla12_xor1_y0;
  assign out[2] = f_u_cla12_xor2_y0;
  assign out[3] = f_u_cla12_xor3_y0;
  assign out[4] = f_u_cla12_xor4_y0;
  assign out[5] = f_u_cla12_xor5_y0;
  assign out[6] = f_u_cla12_xor6_y0;
  assign out[7] = f_u_cla12_xor7_y0;
  assign out[8] = f_u_cla12_xor8_y0;
  assign out[9] = f_u_cla12_xor9_y0;
  assign out[10] = f_u_cla12_xor10_y0;
  assign out[11] = f_u_cla12_xor11_y0;
  assign out[12] = f_u_cla12_or77_y0;
endmodule