module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] fa_xor1, output [0:0] fa_or0);
  wire [0:0] fa_xor0;
  wire [0:0] fa_and0;
  wire [0:0] fa_and1;
  xor_gate xor_gate_fa_xor0(.a(a[0]), .b(b[0]), .out(fa_xor0));
  and_gate and_gate_fa_and0(.a(a[0]), .b(b[0]), .out(fa_and0));
  xor_gate xor_gate_fa_xor1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_xor1));
  and_gate and_gate_fa_and1(.a(fa_xor0[0]), .b(cin[0]), .out(fa_and1));
  or_gate or_gate_fa_or0(.a(fa_and0[0]), .b(fa_and1[0]), .out(fa_or0));
endmodule

module pg_fa(input [0:0] a, input [0:0] b, input [0:0] cin, output [0:0] pg_fa_xor0, output [0:0] pg_fa_and0, output [0:0] pg_fa_xor1);
  xor_gate xor_gate_pg_fa_xor0(.a(a[0]), .b(b[0]), .out(pg_fa_xor0));
  and_gate and_gate_pg_fa_and0(.a(a[0]), .b(b[0]), .out(pg_fa_and0));
  xor_gate xor_gate_pg_fa_xor1(.a(pg_fa_xor0[0]), .b(cin[0]), .out(pg_fa_xor1));
endmodule

module csa_component34(input [33:0] a, input [33:0] b, input [33:0] c, output [69:0] csa_component34_out);
  wire [0:0] csa_component34_fa0_xor1;
  wire [0:0] csa_component34_fa0_or0;
  wire [0:0] csa_component34_fa1_xor1;
  wire [0:0] csa_component34_fa1_or0;
  wire [0:0] csa_component34_fa2_xor1;
  wire [0:0] csa_component34_fa2_or0;
  wire [0:0] csa_component34_fa3_xor1;
  wire [0:0] csa_component34_fa3_or0;
  wire [0:0] csa_component34_fa4_xor1;
  wire [0:0] csa_component34_fa4_or0;
  wire [0:0] csa_component34_fa5_xor1;
  wire [0:0] csa_component34_fa5_or0;
  wire [0:0] csa_component34_fa6_xor1;
  wire [0:0] csa_component34_fa6_or0;
  wire [0:0] csa_component34_fa7_xor1;
  wire [0:0] csa_component34_fa7_or0;
  wire [0:0] csa_component34_fa8_xor1;
  wire [0:0] csa_component34_fa8_or0;
  wire [0:0] csa_component34_fa9_xor1;
  wire [0:0] csa_component34_fa9_or0;
  wire [0:0] csa_component34_fa10_xor1;
  wire [0:0] csa_component34_fa10_or0;
  wire [0:0] csa_component34_fa11_xor1;
  wire [0:0] csa_component34_fa11_or0;
  wire [0:0] csa_component34_fa12_xor1;
  wire [0:0] csa_component34_fa12_or0;
  wire [0:0] csa_component34_fa13_xor1;
  wire [0:0] csa_component34_fa13_or0;
  wire [0:0] csa_component34_fa14_xor1;
  wire [0:0] csa_component34_fa14_or0;
  wire [0:0] csa_component34_fa15_xor1;
  wire [0:0] csa_component34_fa15_or0;
  wire [0:0] csa_component34_fa16_xor1;
  wire [0:0] csa_component34_fa16_or0;
  wire [0:0] csa_component34_fa17_xor1;
  wire [0:0] csa_component34_fa17_or0;
  wire [0:0] csa_component34_fa18_xor1;
  wire [0:0] csa_component34_fa18_or0;
  wire [0:0] csa_component34_fa19_xor1;
  wire [0:0] csa_component34_fa19_or0;
  wire [0:0] csa_component34_fa20_xor1;
  wire [0:0] csa_component34_fa20_or0;
  wire [0:0] csa_component34_fa21_xor1;
  wire [0:0] csa_component34_fa21_or0;
  wire [0:0] csa_component34_fa22_xor1;
  wire [0:0] csa_component34_fa22_or0;
  wire [0:0] csa_component34_fa23_xor1;
  wire [0:0] csa_component34_fa23_or0;
  wire [0:0] csa_component34_fa24_xor1;
  wire [0:0] csa_component34_fa24_or0;
  wire [0:0] csa_component34_fa25_xor1;
  wire [0:0] csa_component34_fa25_or0;
  wire [0:0] csa_component34_fa26_xor1;
  wire [0:0] csa_component34_fa26_or0;
  wire [0:0] csa_component34_fa27_xor1;
  wire [0:0] csa_component34_fa27_or0;
  wire [0:0] csa_component34_fa28_xor1;
  wire [0:0] csa_component34_fa28_or0;
  wire [0:0] csa_component34_fa29_xor1;
  wire [0:0] csa_component34_fa29_or0;
  wire [0:0] csa_component34_fa30_xor1;
  wire [0:0] csa_component34_fa30_or0;
  wire [0:0] csa_component34_fa31_xor1;
  wire [0:0] csa_component34_fa31_or0;
  wire [0:0] csa_component34_fa32_xor1;
  wire [0:0] csa_component34_fa32_or0;
  wire [0:0] csa_component34_fa33_xor1;
  wire [0:0] csa_component34_fa33_or0;

  fa fa_csa_component34_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component34_fa0_xor1), .fa_or0(csa_component34_fa0_or0));
  fa fa_csa_component34_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component34_fa1_xor1), .fa_or0(csa_component34_fa1_or0));
  fa fa_csa_component34_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component34_fa2_xor1), .fa_or0(csa_component34_fa2_or0));
  fa fa_csa_component34_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component34_fa3_xor1), .fa_or0(csa_component34_fa3_or0));
  fa fa_csa_component34_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component34_fa4_xor1), .fa_or0(csa_component34_fa4_or0));
  fa fa_csa_component34_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component34_fa5_xor1), .fa_or0(csa_component34_fa5_or0));
  fa fa_csa_component34_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component34_fa6_xor1), .fa_or0(csa_component34_fa6_or0));
  fa fa_csa_component34_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component34_fa7_xor1), .fa_or0(csa_component34_fa7_or0));
  fa fa_csa_component34_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component34_fa8_xor1), .fa_or0(csa_component34_fa8_or0));
  fa fa_csa_component34_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component34_fa9_xor1), .fa_or0(csa_component34_fa9_or0));
  fa fa_csa_component34_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component34_fa10_xor1), .fa_or0(csa_component34_fa10_or0));
  fa fa_csa_component34_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component34_fa11_xor1), .fa_or0(csa_component34_fa11_or0));
  fa fa_csa_component34_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component34_fa12_xor1), .fa_or0(csa_component34_fa12_or0));
  fa fa_csa_component34_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component34_fa13_xor1), .fa_or0(csa_component34_fa13_or0));
  fa fa_csa_component34_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component34_fa14_xor1), .fa_or0(csa_component34_fa14_or0));
  fa fa_csa_component34_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component34_fa15_xor1), .fa_or0(csa_component34_fa15_or0));
  fa fa_csa_component34_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component34_fa16_xor1), .fa_or0(csa_component34_fa16_or0));
  fa fa_csa_component34_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component34_fa17_xor1), .fa_or0(csa_component34_fa17_or0));
  fa fa_csa_component34_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component34_fa18_xor1), .fa_or0(csa_component34_fa18_or0));
  fa fa_csa_component34_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component34_fa19_xor1), .fa_or0(csa_component34_fa19_or0));
  fa fa_csa_component34_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component34_fa20_xor1), .fa_or0(csa_component34_fa20_or0));
  fa fa_csa_component34_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component34_fa21_xor1), .fa_or0(csa_component34_fa21_or0));
  fa fa_csa_component34_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component34_fa22_xor1), .fa_or0(csa_component34_fa22_or0));
  fa fa_csa_component34_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component34_fa23_xor1), .fa_or0(csa_component34_fa23_or0));
  fa fa_csa_component34_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component34_fa24_xor1), .fa_or0(csa_component34_fa24_or0));
  fa fa_csa_component34_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component34_fa25_xor1), .fa_or0(csa_component34_fa25_or0));
  fa fa_csa_component34_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component34_fa26_xor1), .fa_or0(csa_component34_fa26_or0));
  fa fa_csa_component34_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component34_fa27_xor1), .fa_or0(csa_component34_fa27_or0));
  fa fa_csa_component34_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component34_fa28_xor1), .fa_or0(csa_component34_fa28_or0));
  fa fa_csa_component34_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component34_fa29_xor1), .fa_or0(csa_component34_fa29_or0));
  fa fa_csa_component34_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component34_fa30_xor1), .fa_or0(csa_component34_fa30_or0));
  fa fa_csa_component34_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component34_fa31_xor1), .fa_or0(csa_component34_fa31_or0));
  fa fa_csa_component34_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component34_fa32_xor1), .fa_or0(csa_component34_fa32_or0));
  fa fa_csa_component34_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component34_fa33_xor1), .fa_or0(csa_component34_fa33_or0));

  assign csa_component34_out[0] = csa_component34_fa0_xor1[0];
  assign csa_component34_out[1] = csa_component34_fa1_xor1[0];
  assign csa_component34_out[2] = csa_component34_fa2_xor1[0];
  assign csa_component34_out[3] = csa_component34_fa3_xor1[0];
  assign csa_component34_out[4] = csa_component34_fa4_xor1[0];
  assign csa_component34_out[5] = csa_component34_fa5_xor1[0];
  assign csa_component34_out[6] = csa_component34_fa6_xor1[0];
  assign csa_component34_out[7] = csa_component34_fa7_xor1[0];
  assign csa_component34_out[8] = csa_component34_fa8_xor1[0];
  assign csa_component34_out[9] = csa_component34_fa9_xor1[0];
  assign csa_component34_out[10] = csa_component34_fa10_xor1[0];
  assign csa_component34_out[11] = csa_component34_fa11_xor1[0];
  assign csa_component34_out[12] = csa_component34_fa12_xor1[0];
  assign csa_component34_out[13] = csa_component34_fa13_xor1[0];
  assign csa_component34_out[14] = csa_component34_fa14_xor1[0];
  assign csa_component34_out[15] = csa_component34_fa15_xor1[0];
  assign csa_component34_out[16] = csa_component34_fa16_xor1[0];
  assign csa_component34_out[17] = csa_component34_fa17_xor1[0];
  assign csa_component34_out[18] = csa_component34_fa18_xor1[0];
  assign csa_component34_out[19] = csa_component34_fa19_xor1[0];
  assign csa_component34_out[20] = csa_component34_fa20_xor1[0];
  assign csa_component34_out[21] = csa_component34_fa21_xor1[0];
  assign csa_component34_out[22] = csa_component34_fa22_xor1[0];
  assign csa_component34_out[23] = csa_component34_fa23_xor1[0];
  assign csa_component34_out[24] = csa_component34_fa24_xor1[0];
  assign csa_component34_out[25] = csa_component34_fa25_xor1[0];
  assign csa_component34_out[26] = csa_component34_fa26_xor1[0];
  assign csa_component34_out[27] = csa_component34_fa27_xor1[0];
  assign csa_component34_out[28] = csa_component34_fa28_xor1[0];
  assign csa_component34_out[29] = csa_component34_fa29_xor1[0];
  assign csa_component34_out[30] = csa_component34_fa30_xor1[0];
  assign csa_component34_out[31] = csa_component34_fa31_xor1[0];
  assign csa_component34_out[32] = csa_component34_fa32_xor1[0];
  assign csa_component34_out[33] = csa_component34_fa33_xor1[0];
  assign csa_component34_out[34] = 1'b0;
  assign csa_component34_out[35] = 1'b0;
  assign csa_component34_out[36] = csa_component34_fa0_or0[0];
  assign csa_component34_out[37] = csa_component34_fa1_or0[0];
  assign csa_component34_out[38] = csa_component34_fa2_or0[0];
  assign csa_component34_out[39] = csa_component34_fa3_or0[0];
  assign csa_component34_out[40] = csa_component34_fa4_or0[0];
  assign csa_component34_out[41] = csa_component34_fa5_or0[0];
  assign csa_component34_out[42] = csa_component34_fa6_or0[0];
  assign csa_component34_out[43] = csa_component34_fa7_or0[0];
  assign csa_component34_out[44] = csa_component34_fa8_or0[0];
  assign csa_component34_out[45] = csa_component34_fa9_or0[0];
  assign csa_component34_out[46] = csa_component34_fa10_or0[0];
  assign csa_component34_out[47] = csa_component34_fa11_or0[0];
  assign csa_component34_out[48] = csa_component34_fa12_or0[0];
  assign csa_component34_out[49] = csa_component34_fa13_or0[0];
  assign csa_component34_out[50] = csa_component34_fa14_or0[0];
  assign csa_component34_out[51] = csa_component34_fa15_or0[0];
  assign csa_component34_out[52] = csa_component34_fa16_or0[0];
  assign csa_component34_out[53] = csa_component34_fa17_or0[0];
  assign csa_component34_out[54] = csa_component34_fa18_or0[0];
  assign csa_component34_out[55] = csa_component34_fa19_or0[0];
  assign csa_component34_out[56] = csa_component34_fa20_or0[0];
  assign csa_component34_out[57] = csa_component34_fa21_or0[0];
  assign csa_component34_out[58] = csa_component34_fa22_or0[0];
  assign csa_component34_out[59] = csa_component34_fa23_or0[0];
  assign csa_component34_out[60] = csa_component34_fa24_or0[0];
  assign csa_component34_out[61] = csa_component34_fa25_or0[0];
  assign csa_component34_out[62] = csa_component34_fa26_or0[0];
  assign csa_component34_out[63] = csa_component34_fa27_or0[0];
  assign csa_component34_out[64] = csa_component34_fa28_or0[0];
  assign csa_component34_out[65] = csa_component34_fa29_or0[0];
  assign csa_component34_out[66] = csa_component34_fa30_or0[0];
  assign csa_component34_out[67] = csa_component34_fa31_or0[0];
  assign csa_component34_out[68] = csa_component34_fa32_or0[0];
  assign csa_component34_out[69] = csa_component34_fa33_or0[0];
endmodule

module csa_component37(input [36:0] a, input [36:0] b, input [36:0] c, output [75:0] csa_component37_out);
  wire [0:0] csa_component37_fa0_xor1;
  wire [0:0] csa_component37_fa0_or0;
  wire [0:0] csa_component37_fa1_xor1;
  wire [0:0] csa_component37_fa1_or0;
  wire [0:0] csa_component37_fa2_xor1;
  wire [0:0] csa_component37_fa2_or0;
  wire [0:0] csa_component37_fa3_xor1;
  wire [0:0] csa_component37_fa3_or0;
  wire [0:0] csa_component37_fa4_xor1;
  wire [0:0] csa_component37_fa4_or0;
  wire [0:0] csa_component37_fa5_xor1;
  wire [0:0] csa_component37_fa5_or0;
  wire [0:0] csa_component37_fa6_xor1;
  wire [0:0] csa_component37_fa6_or0;
  wire [0:0] csa_component37_fa7_xor1;
  wire [0:0] csa_component37_fa7_or0;
  wire [0:0] csa_component37_fa8_xor1;
  wire [0:0] csa_component37_fa8_or0;
  wire [0:0] csa_component37_fa9_xor1;
  wire [0:0] csa_component37_fa9_or0;
  wire [0:0] csa_component37_fa10_xor1;
  wire [0:0] csa_component37_fa10_or0;
  wire [0:0] csa_component37_fa11_xor1;
  wire [0:0] csa_component37_fa11_or0;
  wire [0:0] csa_component37_fa12_xor1;
  wire [0:0] csa_component37_fa12_or0;
  wire [0:0] csa_component37_fa13_xor1;
  wire [0:0] csa_component37_fa13_or0;
  wire [0:0] csa_component37_fa14_xor1;
  wire [0:0] csa_component37_fa14_or0;
  wire [0:0] csa_component37_fa15_xor1;
  wire [0:0] csa_component37_fa15_or0;
  wire [0:0] csa_component37_fa16_xor1;
  wire [0:0] csa_component37_fa16_or0;
  wire [0:0] csa_component37_fa17_xor1;
  wire [0:0] csa_component37_fa17_or0;
  wire [0:0] csa_component37_fa18_xor1;
  wire [0:0] csa_component37_fa18_or0;
  wire [0:0] csa_component37_fa19_xor1;
  wire [0:0] csa_component37_fa19_or0;
  wire [0:0] csa_component37_fa20_xor1;
  wire [0:0] csa_component37_fa20_or0;
  wire [0:0] csa_component37_fa21_xor1;
  wire [0:0] csa_component37_fa21_or0;
  wire [0:0] csa_component37_fa22_xor1;
  wire [0:0] csa_component37_fa22_or0;
  wire [0:0] csa_component37_fa23_xor1;
  wire [0:0] csa_component37_fa23_or0;
  wire [0:0] csa_component37_fa24_xor1;
  wire [0:0] csa_component37_fa24_or0;
  wire [0:0] csa_component37_fa25_xor1;
  wire [0:0] csa_component37_fa25_or0;
  wire [0:0] csa_component37_fa26_xor1;
  wire [0:0] csa_component37_fa26_or0;
  wire [0:0] csa_component37_fa27_xor1;
  wire [0:0] csa_component37_fa27_or0;
  wire [0:0] csa_component37_fa28_xor1;
  wire [0:0] csa_component37_fa28_or0;
  wire [0:0] csa_component37_fa29_xor1;
  wire [0:0] csa_component37_fa29_or0;
  wire [0:0] csa_component37_fa30_xor1;
  wire [0:0] csa_component37_fa30_or0;
  wire [0:0] csa_component37_fa31_xor1;
  wire [0:0] csa_component37_fa31_or0;
  wire [0:0] csa_component37_fa32_xor1;
  wire [0:0] csa_component37_fa32_or0;
  wire [0:0] csa_component37_fa33_xor1;
  wire [0:0] csa_component37_fa33_or0;
  wire [0:0] csa_component37_fa34_xor1;
  wire [0:0] csa_component37_fa34_or0;
  wire [0:0] csa_component37_fa35_xor1;
  wire [0:0] csa_component37_fa35_or0;
  wire [0:0] csa_component37_fa36_xor1;
  wire [0:0] csa_component37_fa36_or0;

  fa fa_csa_component37_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component37_fa0_xor1), .fa_or0(csa_component37_fa0_or0));
  fa fa_csa_component37_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component37_fa1_xor1), .fa_or0(csa_component37_fa1_or0));
  fa fa_csa_component37_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component37_fa2_xor1), .fa_or0(csa_component37_fa2_or0));
  fa fa_csa_component37_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component37_fa3_xor1), .fa_or0(csa_component37_fa3_or0));
  fa fa_csa_component37_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component37_fa4_xor1), .fa_or0(csa_component37_fa4_or0));
  fa fa_csa_component37_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component37_fa5_xor1), .fa_or0(csa_component37_fa5_or0));
  fa fa_csa_component37_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component37_fa6_xor1), .fa_or0(csa_component37_fa6_or0));
  fa fa_csa_component37_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component37_fa7_xor1), .fa_or0(csa_component37_fa7_or0));
  fa fa_csa_component37_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component37_fa8_xor1), .fa_or0(csa_component37_fa8_or0));
  fa fa_csa_component37_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component37_fa9_xor1), .fa_or0(csa_component37_fa9_or0));
  fa fa_csa_component37_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component37_fa10_xor1), .fa_or0(csa_component37_fa10_or0));
  fa fa_csa_component37_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component37_fa11_xor1), .fa_or0(csa_component37_fa11_or0));
  fa fa_csa_component37_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component37_fa12_xor1), .fa_or0(csa_component37_fa12_or0));
  fa fa_csa_component37_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component37_fa13_xor1), .fa_or0(csa_component37_fa13_or0));
  fa fa_csa_component37_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component37_fa14_xor1), .fa_or0(csa_component37_fa14_or0));
  fa fa_csa_component37_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component37_fa15_xor1), .fa_or0(csa_component37_fa15_or0));
  fa fa_csa_component37_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component37_fa16_xor1), .fa_or0(csa_component37_fa16_or0));
  fa fa_csa_component37_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component37_fa17_xor1), .fa_or0(csa_component37_fa17_or0));
  fa fa_csa_component37_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component37_fa18_xor1), .fa_or0(csa_component37_fa18_or0));
  fa fa_csa_component37_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component37_fa19_xor1), .fa_or0(csa_component37_fa19_or0));
  fa fa_csa_component37_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component37_fa20_xor1), .fa_or0(csa_component37_fa20_or0));
  fa fa_csa_component37_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component37_fa21_xor1), .fa_or0(csa_component37_fa21_or0));
  fa fa_csa_component37_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component37_fa22_xor1), .fa_or0(csa_component37_fa22_or0));
  fa fa_csa_component37_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component37_fa23_xor1), .fa_or0(csa_component37_fa23_or0));
  fa fa_csa_component37_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component37_fa24_xor1), .fa_or0(csa_component37_fa24_or0));
  fa fa_csa_component37_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component37_fa25_xor1), .fa_or0(csa_component37_fa25_or0));
  fa fa_csa_component37_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component37_fa26_xor1), .fa_or0(csa_component37_fa26_or0));
  fa fa_csa_component37_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component37_fa27_xor1), .fa_or0(csa_component37_fa27_or0));
  fa fa_csa_component37_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component37_fa28_xor1), .fa_or0(csa_component37_fa28_or0));
  fa fa_csa_component37_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component37_fa29_xor1), .fa_or0(csa_component37_fa29_or0));
  fa fa_csa_component37_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component37_fa30_xor1), .fa_or0(csa_component37_fa30_or0));
  fa fa_csa_component37_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component37_fa31_xor1), .fa_or0(csa_component37_fa31_or0));
  fa fa_csa_component37_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component37_fa32_xor1), .fa_or0(csa_component37_fa32_or0));
  fa fa_csa_component37_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component37_fa33_xor1), .fa_or0(csa_component37_fa33_or0));
  fa fa_csa_component37_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component37_fa34_xor1), .fa_or0(csa_component37_fa34_or0));
  fa fa_csa_component37_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component37_fa35_xor1), .fa_or0(csa_component37_fa35_or0));
  fa fa_csa_component37_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component37_fa36_xor1), .fa_or0(csa_component37_fa36_or0));

  assign csa_component37_out[0] = csa_component37_fa0_xor1[0];
  assign csa_component37_out[1] = csa_component37_fa1_xor1[0];
  assign csa_component37_out[2] = csa_component37_fa2_xor1[0];
  assign csa_component37_out[3] = csa_component37_fa3_xor1[0];
  assign csa_component37_out[4] = csa_component37_fa4_xor1[0];
  assign csa_component37_out[5] = csa_component37_fa5_xor1[0];
  assign csa_component37_out[6] = csa_component37_fa6_xor1[0];
  assign csa_component37_out[7] = csa_component37_fa7_xor1[0];
  assign csa_component37_out[8] = csa_component37_fa8_xor1[0];
  assign csa_component37_out[9] = csa_component37_fa9_xor1[0];
  assign csa_component37_out[10] = csa_component37_fa10_xor1[0];
  assign csa_component37_out[11] = csa_component37_fa11_xor1[0];
  assign csa_component37_out[12] = csa_component37_fa12_xor1[0];
  assign csa_component37_out[13] = csa_component37_fa13_xor1[0];
  assign csa_component37_out[14] = csa_component37_fa14_xor1[0];
  assign csa_component37_out[15] = csa_component37_fa15_xor1[0];
  assign csa_component37_out[16] = csa_component37_fa16_xor1[0];
  assign csa_component37_out[17] = csa_component37_fa17_xor1[0];
  assign csa_component37_out[18] = csa_component37_fa18_xor1[0];
  assign csa_component37_out[19] = csa_component37_fa19_xor1[0];
  assign csa_component37_out[20] = csa_component37_fa20_xor1[0];
  assign csa_component37_out[21] = csa_component37_fa21_xor1[0];
  assign csa_component37_out[22] = csa_component37_fa22_xor1[0];
  assign csa_component37_out[23] = csa_component37_fa23_xor1[0];
  assign csa_component37_out[24] = csa_component37_fa24_xor1[0];
  assign csa_component37_out[25] = csa_component37_fa25_xor1[0];
  assign csa_component37_out[26] = csa_component37_fa26_xor1[0];
  assign csa_component37_out[27] = csa_component37_fa27_xor1[0];
  assign csa_component37_out[28] = csa_component37_fa28_xor1[0];
  assign csa_component37_out[29] = csa_component37_fa29_xor1[0];
  assign csa_component37_out[30] = csa_component37_fa30_xor1[0];
  assign csa_component37_out[31] = csa_component37_fa31_xor1[0];
  assign csa_component37_out[32] = csa_component37_fa32_xor1[0];
  assign csa_component37_out[33] = csa_component37_fa33_xor1[0];
  assign csa_component37_out[34] = csa_component37_fa34_xor1[0];
  assign csa_component37_out[35] = csa_component37_fa35_xor1[0];
  assign csa_component37_out[36] = csa_component37_fa36_xor1[0];
  assign csa_component37_out[37] = 1'b0;
  assign csa_component37_out[38] = 1'b0;
  assign csa_component37_out[39] = csa_component37_fa0_or0[0];
  assign csa_component37_out[40] = csa_component37_fa1_or0[0];
  assign csa_component37_out[41] = csa_component37_fa2_or0[0];
  assign csa_component37_out[42] = csa_component37_fa3_or0[0];
  assign csa_component37_out[43] = csa_component37_fa4_or0[0];
  assign csa_component37_out[44] = csa_component37_fa5_or0[0];
  assign csa_component37_out[45] = csa_component37_fa6_or0[0];
  assign csa_component37_out[46] = csa_component37_fa7_or0[0];
  assign csa_component37_out[47] = csa_component37_fa8_or0[0];
  assign csa_component37_out[48] = csa_component37_fa9_or0[0];
  assign csa_component37_out[49] = csa_component37_fa10_or0[0];
  assign csa_component37_out[50] = csa_component37_fa11_or0[0];
  assign csa_component37_out[51] = csa_component37_fa12_or0[0];
  assign csa_component37_out[52] = csa_component37_fa13_or0[0];
  assign csa_component37_out[53] = csa_component37_fa14_or0[0];
  assign csa_component37_out[54] = csa_component37_fa15_or0[0];
  assign csa_component37_out[55] = csa_component37_fa16_or0[0];
  assign csa_component37_out[56] = csa_component37_fa17_or0[0];
  assign csa_component37_out[57] = csa_component37_fa18_or0[0];
  assign csa_component37_out[58] = csa_component37_fa19_or0[0];
  assign csa_component37_out[59] = csa_component37_fa20_or0[0];
  assign csa_component37_out[60] = csa_component37_fa21_or0[0];
  assign csa_component37_out[61] = csa_component37_fa22_or0[0];
  assign csa_component37_out[62] = csa_component37_fa23_or0[0];
  assign csa_component37_out[63] = csa_component37_fa24_or0[0];
  assign csa_component37_out[64] = csa_component37_fa25_or0[0];
  assign csa_component37_out[65] = csa_component37_fa26_or0[0];
  assign csa_component37_out[66] = csa_component37_fa27_or0[0];
  assign csa_component37_out[67] = csa_component37_fa28_or0[0];
  assign csa_component37_out[68] = csa_component37_fa29_or0[0];
  assign csa_component37_out[69] = csa_component37_fa30_or0[0];
  assign csa_component37_out[70] = csa_component37_fa31_or0[0];
  assign csa_component37_out[71] = csa_component37_fa32_or0[0];
  assign csa_component37_out[72] = csa_component37_fa33_or0[0];
  assign csa_component37_out[73] = csa_component37_fa34_or0[0];
  assign csa_component37_out[74] = csa_component37_fa35_or0[0];
  assign csa_component37_out[75] = csa_component37_fa36_or0[0];
endmodule

module csa_component40(input [39:0] a, input [39:0] b, input [39:0] c, output [81:0] csa_component40_out);
  wire [0:0] csa_component40_fa0_xor1;
  wire [0:0] csa_component40_fa0_or0;
  wire [0:0] csa_component40_fa1_xor1;
  wire [0:0] csa_component40_fa1_or0;
  wire [0:0] csa_component40_fa2_xor1;
  wire [0:0] csa_component40_fa2_or0;
  wire [0:0] csa_component40_fa3_xor1;
  wire [0:0] csa_component40_fa3_or0;
  wire [0:0] csa_component40_fa4_xor1;
  wire [0:0] csa_component40_fa4_or0;
  wire [0:0] csa_component40_fa5_xor1;
  wire [0:0] csa_component40_fa5_or0;
  wire [0:0] csa_component40_fa6_xor1;
  wire [0:0] csa_component40_fa6_or0;
  wire [0:0] csa_component40_fa7_xor1;
  wire [0:0] csa_component40_fa7_or0;
  wire [0:0] csa_component40_fa8_xor1;
  wire [0:0] csa_component40_fa8_or0;
  wire [0:0] csa_component40_fa9_xor1;
  wire [0:0] csa_component40_fa9_or0;
  wire [0:0] csa_component40_fa10_xor1;
  wire [0:0] csa_component40_fa10_or0;
  wire [0:0] csa_component40_fa11_xor1;
  wire [0:0] csa_component40_fa11_or0;
  wire [0:0] csa_component40_fa12_xor1;
  wire [0:0] csa_component40_fa12_or0;
  wire [0:0] csa_component40_fa13_xor1;
  wire [0:0] csa_component40_fa13_or0;
  wire [0:0] csa_component40_fa14_xor1;
  wire [0:0] csa_component40_fa14_or0;
  wire [0:0] csa_component40_fa15_xor1;
  wire [0:0] csa_component40_fa15_or0;
  wire [0:0] csa_component40_fa16_xor1;
  wire [0:0] csa_component40_fa16_or0;
  wire [0:0] csa_component40_fa17_xor1;
  wire [0:0] csa_component40_fa17_or0;
  wire [0:0] csa_component40_fa18_xor1;
  wire [0:0] csa_component40_fa18_or0;
  wire [0:0] csa_component40_fa19_xor1;
  wire [0:0] csa_component40_fa19_or0;
  wire [0:0] csa_component40_fa20_xor1;
  wire [0:0] csa_component40_fa20_or0;
  wire [0:0] csa_component40_fa21_xor1;
  wire [0:0] csa_component40_fa21_or0;
  wire [0:0] csa_component40_fa22_xor1;
  wire [0:0] csa_component40_fa22_or0;
  wire [0:0] csa_component40_fa23_xor1;
  wire [0:0] csa_component40_fa23_or0;
  wire [0:0] csa_component40_fa24_xor1;
  wire [0:0] csa_component40_fa24_or0;
  wire [0:0] csa_component40_fa25_xor1;
  wire [0:0] csa_component40_fa25_or0;
  wire [0:0] csa_component40_fa26_xor1;
  wire [0:0] csa_component40_fa26_or0;
  wire [0:0] csa_component40_fa27_xor1;
  wire [0:0] csa_component40_fa27_or0;
  wire [0:0] csa_component40_fa28_xor1;
  wire [0:0] csa_component40_fa28_or0;
  wire [0:0] csa_component40_fa29_xor1;
  wire [0:0] csa_component40_fa29_or0;
  wire [0:0] csa_component40_fa30_xor1;
  wire [0:0] csa_component40_fa30_or0;
  wire [0:0] csa_component40_fa31_xor1;
  wire [0:0] csa_component40_fa31_or0;
  wire [0:0] csa_component40_fa32_xor1;
  wire [0:0] csa_component40_fa32_or0;
  wire [0:0] csa_component40_fa33_xor1;
  wire [0:0] csa_component40_fa33_or0;
  wire [0:0] csa_component40_fa34_xor1;
  wire [0:0] csa_component40_fa34_or0;
  wire [0:0] csa_component40_fa35_xor1;
  wire [0:0] csa_component40_fa35_or0;
  wire [0:0] csa_component40_fa36_xor1;
  wire [0:0] csa_component40_fa36_or0;
  wire [0:0] csa_component40_fa37_xor1;
  wire [0:0] csa_component40_fa37_or0;
  wire [0:0] csa_component40_fa38_xor1;
  wire [0:0] csa_component40_fa38_or0;
  wire [0:0] csa_component40_fa39_xor1;
  wire [0:0] csa_component40_fa39_or0;

  fa fa_csa_component40_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component40_fa0_xor1), .fa_or0(csa_component40_fa0_or0));
  fa fa_csa_component40_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component40_fa1_xor1), .fa_or0(csa_component40_fa1_or0));
  fa fa_csa_component40_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component40_fa2_xor1), .fa_or0(csa_component40_fa2_or0));
  fa fa_csa_component40_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component40_fa3_xor1), .fa_or0(csa_component40_fa3_or0));
  fa fa_csa_component40_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component40_fa4_xor1), .fa_or0(csa_component40_fa4_or0));
  fa fa_csa_component40_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component40_fa5_xor1), .fa_or0(csa_component40_fa5_or0));
  fa fa_csa_component40_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component40_fa6_xor1), .fa_or0(csa_component40_fa6_or0));
  fa fa_csa_component40_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component40_fa7_xor1), .fa_or0(csa_component40_fa7_or0));
  fa fa_csa_component40_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component40_fa8_xor1), .fa_or0(csa_component40_fa8_or0));
  fa fa_csa_component40_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component40_fa9_xor1), .fa_or0(csa_component40_fa9_or0));
  fa fa_csa_component40_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component40_fa10_xor1), .fa_or0(csa_component40_fa10_or0));
  fa fa_csa_component40_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component40_fa11_xor1), .fa_or0(csa_component40_fa11_or0));
  fa fa_csa_component40_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component40_fa12_xor1), .fa_or0(csa_component40_fa12_or0));
  fa fa_csa_component40_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component40_fa13_xor1), .fa_or0(csa_component40_fa13_or0));
  fa fa_csa_component40_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component40_fa14_xor1), .fa_or0(csa_component40_fa14_or0));
  fa fa_csa_component40_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component40_fa15_xor1), .fa_or0(csa_component40_fa15_or0));
  fa fa_csa_component40_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component40_fa16_xor1), .fa_or0(csa_component40_fa16_or0));
  fa fa_csa_component40_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component40_fa17_xor1), .fa_or0(csa_component40_fa17_or0));
  fa fa_csa_component40_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component40_fa18_xor1), .fa_or0(csa_component40_fa18_or0));
  fa fa_csa_component40_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component40_fa19_xor1), .fa_or0(csa_component40_fa19_or0));
  fa fa_csa_component40_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component40_fa20_xor1), .fa_or0(csa_component40_fa20_or0));
  fa fa_csa_component40_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component40_fa21_xor1), .fa_or0(csa_component40_fa21_or0));
  fa fa_csa_component40_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component40_fa22_xor1), .fa_or0(csa_component40_fa22_or0));
  fa fa_csa_component40_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component40_fa23_xor1), .fa_or0(csa_component40_fa23_or0));
  fa fa_csa_component40_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component40_fa24_xor1), .fa_or0(csa_component40_fa24_or0));
  fa fa_csa_component40_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component40_fa25_xor1), .fa_or0(csa_component40_fa25_or0));
  fa fa_csa_component40_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component40_fa26_xor1), .fa_or0(csa_component40_fa26_or0));
  fa fa_csa_component40_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component40_fa27_xor1), .fa_or0(csa_component40_fa27_or0));
  fa fa_csa_component40_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component40_fa28_xor1), .fa_or0(csa_component40_fa28_or0));
  fa fa_csa_component40_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component40_fa29_xor1), .fa_or0(csa_component40_fa29_or0));
  fa fa_csa_component40_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component40_fa30_xor1), .fa_or0(csa_component40_fa30_or0));
  fa fa_csa_component40_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component40_fa31_xor1), .fa_or0(csa_component40_fa31_or0));
  fa fa_csa_component40_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component40_fa32_xor1), .fa_or0(csa_component40_fa32_or0));
  fa fa_csa_component40_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component40_fa33_xor1), .fa_or0(csa_component40_fa33_or0));
  fa fa_csa_component40_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component40_fa34_xor1), .fa_or0(csa_component40_fa34_or0));
  fa fa_csa_component40_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component40_fa35_xor1), .fa_or0(csa_component40_fa35_or0));
  fa fa_csa_component40_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component40_fa36_xor1), .fa_or0(csa_component40_fa36_or0));
  fa fa_csa_component40_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component40_fa37_xor1), .fa_or0(csa_component40_fa37_or0));
  fa fa_csa_component40_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component40_fa38_xor1), .fa_or0(csa_component40_fa38_or0));
  fa fa_csa_component40_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component40_fa39_xor1), .fa_or0(csa_component40_fa39_or0));

  assign csa_component40_out[0] = csa_component40_fa0_xor1[0];
  assign csa_component40_out[1] = csa_component40_fa1_xor1[0];
  assign csa_component40_out[2] = csa_component40_fa2_xor1[0];
  assign csa_component40_out[3] = csa_component40_fa3_xor1[0];
  assign csa_component40_out[4] = csa_component40_fa4_xor1[0];
  assign csa_component40_out[5] = csa_component40_fa5_xor1[0];
  assign csa_component40_out[6] = csa_component40_fa6_xor1[0];
  assign csa_component40_out[7] = csa_component40_fa7_xor1[0];
  assign csa_component40_out[8] = csa_component40_fa8_xor1[0];
  assign csa_component40_out[9] = csa_component40_fa9_xor1[0];
  assign csa_component40_out[10] = csa_component40_fa10_xor1[0];
  assign csa_component40_out[11] = csa_component40_fa11_xor1[0];
  assign csa_component40_out[12] = csa_component40_fa12_xor1[0];
  assign csa_component40_out[13] = csa_component40_fa13_xor1[0];
  assign csa_component40_out[14] = csa_component40_fa14_xor1[0];
  assign csa_component40_out[15] = csa_component40_fa15_xor1[0];
  assign csa_component40_out[16] = csa_component40_fa16_xor1[0];
  assign csa_component40_out[17] = csa_component40_fa17_xor1[0];
  assign csa_component40_out[18] = csa_component40_fa18_xor1[0];
  assign csa_component40_out[19] = csa_component40_fa19_xor1[0];
  assign csa_component40_out[20] = csa_component40_fa20_xor1[0];
  assign csa_component40_out[21] = csa_component40_fa21_xor1[0];
  assign csa_component40_out[22] = csa_component40_fa22_xor1[0];
  assign csa_component40_out[23] = csa_component40_fa23_xor1[0];
  assign csa_component40_out[24] = csa_component40_fa24_xor1[0];
  assign csa_component40_out[25] = csa_component40_fa25_xor1[0];
  assign csa_component40_out[26] = csa_component40_fa26_xor1[0];
  assign csa_component40_out[27] = csa_component40_fa27_xor1[0];
  assign csa_component40_out[28] = csa_component40_fa28_xor1[0];
  assign csa_component40_out[29] = csa_component40_fa29_xor1[0];
  assign csa_component40_out[30] = csa_component40_fa30_xor1[0];
  assign csa_component40_out[31] = csa_component40_fa31_xor1[0];
  assign csa_component40_out[32] = csa_component40_fa32_xor1[0];
  assign csa_component40_out[33] = csa_component40_fa33_xor1[0];
  assign csa_component40_out[34] = csa_component40_fa34_xor1[0];
  assign csa_component40_out[35] = csa_component40_fa35_xor1[0];
  assign csa_component40_out[36] = csa_component40_fa36_xor1[0];
  assign csa_component40_out[37] = csa_component40_fa37_xor1[0];
  assign csa_component40_out[38] = csa_component40_fa38_xor1[0];
  assign csa_component40_out[39] = csa_component40_fa39_xor1[0];
  assign csa_component40_out[40] = 1'b0;
  assign csa_component40_out[41] = 1'b0;
  assign csa_component40_out[42] = csa_component40_fa0_or0[0];
  assign csa_component40_out[43] = csa_component40_fa1_or0[0];
  assign csa_component40_out[44] = csa_component40_fa2_or0[0];
  assign csa_component40_out[45] = csa_component40_fa3_or0[0];
  assign csa_component40_out[46] = csa_component40_fa4_or0[0];
  assign csa_component40_out[47] = csa_component40_fa5_or0[0];
  assign csa_component40_out[48] = csa_component40_fa6_or0[0];
  assign csa_component40_out[49] = csa_component40_fa7_or0[0];
  assign csa_component40_out[50] = csa_component40_fa8_or0[0];
  assign csa_component40_out[51] = csa_component40_fa9_or0[0];
  assign csa_component40_out[52] = csa_component40_fa10_or0[0];
  assign csa_component40_out[53] = csa_component40_fa11_or0[0];
  assign csa_component40_out[54] = csa_component40_fa12_or0[0];
  assign csa_component40_out[55] = csa_component40_fa13_or0[0];
  assign csa_component40_out[56] = csa_component40_fa14_or0[0];
  assign csa_component40_out[57] = csa_component40_fa15_or0[0];
  assign csa_component40_out[58] = csa_component40_fa16_or0[0];
  assign csa_component40_out[59] = csa_component40_fa17_or0[0];
  assign csa_component40_out[60] = csa_component40_fa18_or0[0];
  assign csa_component40_out[61] = csa_component40_fa19_or0[0];
  assign csa_component40_out[62] = csa_component40_fa20_or0[0];
  assign csa_component40_out[63] = csa_component40_fa21_or0[0];
  assign csa_component40_out[64] = csa_component40_fa22_or0[0];
  assign csa_component40_out[65] = csa_component40_fa23_or0[0];
  assign csa_component40_out[66] = csa_component40_fa24_or0[0];
  assign csa_component40_out[67] = csa_component40_fa25_or0[0];
  assign csa_component40_out[68] = csa_component40_fa26_or0[0];
  assign csa_component40_out[69] = csa_component40_fa27_or0[0];
  assign csa_component40_out[70] = csa_component40_fa28_or0[0];
  assign csa_component40_out[71] = csa_component40_fa29_or0[0];
  assign csa_component40_out[72] = csa_component40_fa30_or0[0];
  assign csa_component40_out[73] = csa_component40_fa31_or0[0];
  assign csa_component40_out[74] = csa_component40_fa32_or0[0];
  assign csa_component40_out[75] = csa_component40_fa33_or0[0];
  assign csa_component40_out[76] = csa_component40_fa34_or0[0];
  assign csa_component40_out[77] = csa_component40_fa35_or0[0];
  assign csa_component40_out[78] = csa_component40_fa36_or0[0];
  assign csa_component40_out[79] = csa_component40_fa37_or0[0];
  assign csa_component40_out[80] = csa_component40_fa38_or0[0];
  assign csa_component40_out[81] = csa_component40_fa39_or0[0];
endmodule

module csa_component43(input [42:0] a, input [42:0] b, input [42:0] c, output [87:0] csa_component43_out);
  wire [0:0] csa_component43_fa0_xor1;
  wire [0:0] csa_component43_fa0_or0;
  wire [0:0] csa_component43_fa1_xor1;
  wire [0:0] csa_component43_fa1_or0;
  wire [0:0] csa_component43_fa2_xor1;
  wire [0:0] csa_component43_fa2_or0;
  wire [0:0] csa_component43_fa3_xor1;
  wire [0:0] csa_component43_fa3_or0;
  wire [0:0] csa_component43_fa4_xor1;
  wire [0:0] csa_component43_fa4_or0;
  wire [0:0] csa_component43_fa5_xor1;
  wire [0:0] csa_component43_fa5_or0;
  wire [0:0] csa_component43_fa6_xor1;
  wire [0:0] csa_component43_fa6_or0;
  wire [0:0] csa_component43_fa7_xor1;
  wire [0:0] csa_component43_fa7_or0;
  wire [0:0] csa_component43_fa8_xor1;
  wire [0:0] csa_component43_fa8_or0;
  wire [0:0] csa_component43_fa9_xor1;
  wire [0:0] csa_component43_fa9_or0;
  wire [0:0] csa_component43_fa10_xor1;
  wire [0:0] csa_component43_fa10_or0;
  wire [0:0] csa_component43_fa11_xor1;
  wire [0:0] csa_component43_fa11_or0;
  wire [0:0] csa_component43_fa12_xor1;
  wire [0:0] csa_component43_fa12_or0;
  wire [0:0] csa_component43_fa13_xor1;
  wire [0:0] csa_component43_fa13_or0;
  wire [0:0] csa_component43_fa14_xor1;
  wire [0:0] csa_component43_fa14_or0;
  wire [0:0] csa_component43_fa15_xor1;
  wire [0:0] csa_component43_fa15_or0;
  wire [0:0] csa_component43_fa16_xor1;
  wire [0:0] csa_component43_fa16_or0;
  wire [0:0] csa_component43_fa17_xor1;
  wire [0:0] csa_component43_fa17_or0;
  wire [0:0] csa_component43_fa18_xor1;
  wire [0:0] csa_component43_fa18_or0;
  wire [0:0] csa_component43_fa19_xor1;
  wire [0:0] csa_component43_fa19_or0;
  wire [0:0] csa_component43_fa20_xor1;
  wire [0:0] csa_component43_fa20_or0;
  wire [0:0] csa_component43_fa21_xor1;
  wire [0:0] csa_component43_fa21_or0;
  wire [0:0] csa_component43_fa22_xor1;
  wire [0:0] csa_component43_fa22_or0;
  wire [0:0] csa_component43_fa23_xor1;
  wire [0:0] csa_component43_fa23_or0;
  wire [0:0] csa_component43_fa24_xor1;
  wire [0:0] csa_component43_fa24_or0;
  wire [0:0] csa_component43_fa25_xor1;
  wire [0:0] csa_component43_fa25_or0;
  wire [0:0] csa_component43_fa26_xor1;
  wire [0:0] csa_component43_fa26_or0;
  wire [0:0] csa_component43_fa27_xor1;
  wire [0:0] csa_component43_fa27_or0;
  wire [0:0] csa_component43_fa28_xor1;
  wire [0:0] csa_component43_fa28_or0;
  wire [0:0] csa_component43_fa29_xor1;
  wire [0:0] csa_component43_fa29_or0;
  wire [0:0] csa_component43_fa30_xor1;
  wire [0:0] csa_component43_fa30_or0;
  wire [0:0] csa_component43_fa31_xor1;
  wire [0:0] csa_component43_fa31_or0;
  wire [0:0] csa_component43_fa32_xor1;
  wire [0:0] csa_component43_fa32_or0;
  wire [0:0] csa_component43_fa33_xor1;
  wire [0:0] csa_component43_fa33_or0;
  wire [0:0] csa_component43_fa34_xor1;
  wire [0:0] csa_component43_fa34_or0;
  wire [0:0] csa_component43_fa35_xor1;
  wire [0:0] csa_component43_fa35_or0;
  wire [0:0] csa_component43_fa36_xor1;
  wire [0:0] csa_component43_fa36_or0;
  wire [0:0] csa_component43_fa37_xor1;
  wire [0:0] csa_component43_fa37_or0;
  wire [0:0] csa_component43_fa38_xor1;
  wire [0:0] csa_component43_fa38_or0;
  wire [0:0] csa_component43_fa39_xor1;
  wire [0:0] csa_component43_fa39_or0;
  wire [0:0] csa_component43_fa40_xor1;
  wire [0:0] csa_component43_fa40_or0;
  wire [0:0] csa_component43_fa41_xor1;
  wire [0:0] csa_component43_fa41_or0;
  wire [0:0] csa_component43_fa42_xor1;
  wire [0:0] csa_component43_fa42_or0;

  fa fa_csa_component43_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component43_fa0_xor1), .fa_or0(csa_component43_fa0_or0));
  fa fa_csa_component43_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component43_fa1_xor1), .fa_or0(csa_component43_fa1_or0));
  fa fa_csa_component43_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component43_fa2_xor1), .fa_or0(csa_component43_fa2_or0));
  fa fa_csa_component43_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component43_fa3_xor1), .fa_or0(csa_component43_fa3_or0));
  fa fa_csa_component43_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component43_fa4_xor1), .fa_or0(csa_component43_fa4_or0));
  fa fa_csa_component43_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component43_fa5_xor1), .fa_or0(csa_component43_fa5_or0));
  fa fa_csa_component43_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component43_fa6_xor1), .fa_or0(csa_component43_fa6_or0));
  fa fa_csa_component43_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component43_fa7_xor1), .fa_or0(csa_component43_fa7_or0));
  fa fa_csa_component43_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component43_fa8_xor1), .fa_or0(csa_component43_fa8_or0));
  fa fa_csa_component43_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component43_fa9_xor1), .fa_or0(csa_component43_fa9_or0));
  fa fa_csa_component43_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component43_fa10_xor1), .fa_or0(csa_component43_fa10_or0));
  fa fa_csa_component43_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component43_fa11_xor1), .fa_or0(csa_component43_fa11_or0));
  fa fa_csa_component43_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component43_fa12_xor1), .fa_or0(csa_component43_fa12_or0));
  fa fa_csa_component43_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component43_fa13_xor1), .fa_or0(csa_component43_fa13_or0));
  fa fa_csa_component43_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component43_fa14_xor1), .fa_or0(csa_component43_fa14_or0));
  fa fa_csa_component43_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component43_fa15_xor1), .fa_or0(csa_component43_fa15_or0));
  fa fa_csa_component43_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component43_fa16_xor1), .fa_or0(csa_component43_fa16_or0));
  fa fa_csa_component43_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component43_fa17_xor1), .fa_or0(csa_component43_fa17_or0));
  fa fa_csa_component43_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component43_fa18_xor1), .fa_or0(csa_component43_fa18_or0));
  fa fa_csa_component43_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component43_fa19_xor1), .fa_or0(csa_component43_fa19_or0));
  fa fa_csa_component43_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component43_fa20_xor1), .fa_or0(csa_component43_fa20_or0));
  fa fa_csa_component43_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component43_fa21_xor1), .fa_or0(csa_component43_fa21_or0));
  fa fa_csa_component43_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component43_fa22_xor1), .fa_or0(csa_component43_fa22_or0));
  fa fa_csa_component43_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component43_fa23_xor1), .fa_or0(csa_component43_fa23_or0));
  fa fa_csa_component43_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component43_fa24_xor1), .fa_or0(csa_component43_fa24_or0));
  fa fa_csa_component43_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component43_fa25_xor1), .fa_or0(csa_component43_fa25_or0));
  fa fa_csa_component43_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component43_fa26_xor1), .fa_or0(csa_component43_fa26_or0));
  fa fa_csa_component43_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component43_fa27_xor1), .fa_or0(csa_component43_fa27_or0));
  fa fa_csa_component43_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component43_fa28_xor1), .fa_or0(csa_component43_fa28_or0));
  fa fa_csa_component43_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component43_fa29_xor1), .fa_or0(csa_component43_fa29_or0));
  fa fa_csa_component43_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component43_fa30_xor1), .fa_or0(csa_component43_fa30_or0));
  fa fa_csa_component43_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component43_fa31_xor1), .fa_or0(csa_component43_fa31_or0));
  fa fa_csa_component43_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component43_fa32_xor1), .fa_or0(csa_component43_fa32_or0));
  fa fa_csa_component43_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component43_fa33_xor1), .fa_or0(csa_component43_fa33_or0));
  fa fa_csa_component43_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component43_fa34_xor1), .fa_or0(csa_component43_fa34_or0));
  fa fa_csa_component43_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component43_fa35_xor1), .fa_or0(csa_component43_fa35_or0));
  fa fa_csa_component43_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component43_fa36_xor1), .fa_or0(csa_component43_fa36_or0));
  fa fa_csa_component43_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component43_fa37_xor1), .fa_or0(csa_component43_fa37_or0));
  fa fa_csa_component43_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component43_fa38_xor1), .fa_or0(csa_component43_fa38_or0));
  fa fa_csa_component43_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component43_fa39_xor1), .fa_or0(csa_component43_fa39_or0));
  fa fa_csa_component43_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component43_fa40_xor1), .fa_or0(csa_component43_fa40_or0));
  fa fa_csa_component43_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component43_fa41_xor1), .fa_or0(csa_component43_fa41_or0));
  fa fa_csa_component43_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component43_fa42_xor1), .fa_or0(csa_component43_fa42_or0));

  assign csa_component43_out[0] = csa_component43_fa0_xor1[0];
  assign csa_component43_out[1] = csa_component43_fa1_xor1[0];
  assign csa_component43_out[2] = csa_component43_fa2_xor1[0];
  assign csa_component43_out[3] = csa_component43_fa3_xor1[0];
  assign csa_component43_out[4] = csa_component43_fa4_xor1[0];
  assign csa_component43_out[5] = csa_component43_fa5_xor1[0];
  assign csa_component43_out[6] = csa_component43_fa6_xor1[0];
  assign csa_component43_out[7] = csa_component43_fa7_xor1[0];
  assign csa_component43_out[8] = csa_component43_fa8_xor1[0];
  assign csa_component43_out[9] = csa_component43_fa9_xor1[0];
  assign csa_component43_out[10] = csa_component43_fa10_xor1[0];
  assign csa_component43_out[11] = csa_component43_fa11_xor1[0];
  assign csa_component43_out[12] = csa_component43_fa12_xor1[0];
  assign csa_component43_out[13] = csa_component43_fa13_xor1[0];
  assign csa_component43_out[14] = csa_component43_fa14_xor1[0];
  assign csa_component43_out[15] = csa_component43_fa15_xor1[0];
  assign csa_component43_out[16] = csa_component43_fa16_xor1[0];
  assign csa_component43_out[17] = csa_component43_fa17_xor1[0];
  assign csa_component43_out[18] = csa_component43_fa18_xor1[0];
  assign csa_component43_out[19] = csa_component43_fa19_xor1[0];
  assign csa_component43_out[20] = csa_component43_fa20_xor1[0];
  assign csa_component43_out[21] = csa_component43_fa21_xor1[0];
  assign csa_component43_out[22] = csa_component43_fa22_xor1[0];
  assign csa_component43_out[23] = csa_component43_fa23_xor1[0];
  assign csa_component43_out[24] = csa_component43_fa24_xor1[0];
  assign csa_component43_out[25] = csa_component43_fa25_xor1[0];
  assign csa_component43_out[26] = csa_component43_fa26_xor1[0];
  assign csa_component43_out[27] = csa_component43_fa27_xor1[0];
  assign csa_component43_out[28] = csa_component43_fa28_xor1[0];
  assign csa_component43_out[29] = csa_component43_fa29_xor1[0];
  assign csa_component43_out[30] = csa_component43_fa30_xor1[0];
  assign csa_component43_out[31] = csa_component43_fa31_xor1[0];
  assign csa_component43_out[32] = csa_component43_fa32_xor1[0];
  assign csa_component43_out[33] = csa_component43_fa33_xor1[0];
  assign csa_component43_out[34] = csa_component43_fa34_xor1[0];
  assign csa_component43_out[35] = csa_component43_fa35_xor1[0];
  assign csa_component43_out[36] = csa_component43_fa36_xor1[0];
  assign csa_component43_out[37] = csa_component43_fa37_xor1[0];
  assign csa_component43_out[38] = csa_component43_fa38_xor1[0];
  assign csa_component43_out[39] = csa_component43_fa39_xor1[0];
  assign csa_component43_out[40] = csa_component43_fa40_xor1[0];
  assign csa_component43_out[41] = csa_component43_fa41_xor1[0];
  assign csa_component43_out[42] = csa_component43_fa42_xor1[0];
  assign csa_component43_out[43] = 1'b0;
  assign csa_component43_out[44] = 1'b0;
  assign csa_component43_out[45] = csa_component43_fa0_or0[0];
  assign csa_component43_out[46] = csa_component43_fa1_or0[0];
  assign csa_component43_out[47] = csa_component43_fa2_or0[0];
  assign csa_component43_out[48] = csa_component43_fa3_or0[0];
  assign csa_component43_out[49] = csa_component43_fa4_or0[0];
  assign csa_component43_out[50] = csa_component43_fa5_or0[0];
  assign csa_component43_out[51] = csa_component43_fa6_or0[0];
  assign csa_component43_out[52] = csa_component43_fa7_or0[0];
  assign csa_component43_out[53] = csa_component43_fa8_or0[0];
  assign csa_component43_out[54] = csa_component43_fa9_or0[0];
  assign csa_component43_out[55] = csa_component43_fa10_or0[0];
  assign csa_component43_out[56] = csa_component43_fa11_or0[0];
  assign csa_component43_out[57] = csa_component43_fa12_or0[0];
  assign csa_component43_out[58] = csa_component43_fa13_or0[0];
  assign csa_component43_out[59] = csa_component43_fa14_or0[0];
  assign csa_component43_out[60] = csa_component43_fa15_or0[0];
  assign csa_component43_out[61] = csa_component43_fa16_or0[0];
  assign csa_component43_out[62] = csa_component43_fa17_or0[0];
  assign csa_component43_out[63] = csa_component43_fa18_or0[0];
  assign csa_component43_out[64] = csa_component43_fa19_or0[0];
  assign csa_component43_out[65] = csa_component43_fa20_or0[0];
  assign csa_component43_out[66] = csa_component43_fa21_or0[0];
  assign csa_component43_out[67] = csa_component43_fa22_or0[0];
  assign csa_component43_out[68] = csa_component43_fa23_or0[0];
  assign csa_component43_out[69] = csa_component43_fa24_or0[0];
  assign csa_component43_out[70] = csa_component43_fa25_or0[0];
  assign csa_component43_out[71] = csa_component43_fa26_or0[0];
  assign csa_component43_out[72] = csa_component43_fa27_or0[0];
  assign csa_component43_out[73] = csa_component43_fa28_or0[0];
  assign csa_component43_out[74] = csa_component43_fa29_or0[0];
  assign csa_component43_out[75] = csa_component43_fa30_or0[0];
  assign csa_component43_out[76] = csa_component43_fa31_or0[0];
  assign csa_component43_out[77] = csa_component43_fa32_or0[0];
  assign csa_component43_out[78] = csa_component43_fa33_or0[0];
  assign csa_component43_out[79] = csa_component43_fa34_or0[0];
  assign csa_component43_out[80] = csa_component43_fa35_or0[0];
  assign csa_component43_out[81] = csa_component43_fa36_or0[0];
  assign csa_component43_out[82] = csa_component43_fa37_or0[0];
  assign csa_component43_out[83] = csa_component43_fa38_or0[0];
  assign csa_component43_out[84] = csa_component43_fa39_or0[0];
  assign csa_component43_out[85] = csa_component43_fa40_or0[0];
  assign csa_component43_out[86] = csa_component43_fa41_or0[0];
  assign csa_component43_out[87] = csa_component43_fa42_or0[0];
endmodule

module csa_component46(input [45:0] a, input [45:0] b, input [45:0] c, output [93:0] csa_component46_out);
  wire [0:0] csa_component46_fa0_xor1;
  wire [0:0] csa_component46_fa0_or0;
  wire [0:0] csa_component46_fa1_xor1;
  wire [0:0] csa_component46_fa1_or0;
  wire [0:0] csa_component46_fa2_xor1;
  wire [0:0] csa_component46_fa2_or0;
  wire [0:0] csa_component46_fa3_xor1;
  wire [0:0] csa_component46_fa3_or0;
  wire [0:0] csa_component46_fa4_xor1;
  wire [0:0] csa_component46_fa4_or0;
  wire [0:0] csa_component46_fa5_xor1;
  wire [0:0] csa_component46_fa5_or0;
  wire [0:0] csa_component46_fa6_xor1;
  wire [0:0] csa_component46_fa6_or0;
  wire [0:0] csa_component46_fa7_xor1;
  wire [0:0] csa_component46_fa7_or0;
  wire [0:0] csa_component46_fa8_xor1;
  wire [0:0] csa_component46_fa8_or0;
  wire [0:0] csa_component46_fa9_xor1;
  wire [0:0] csa_component46_fa9_or0;
  wire [0:0] csa_component46_fa10_xor1;
  wire [0:0] csa_component46_fa10_or0;
  wire [0:0] csa_component46_fa11_xor1;
  wire [0:0] csa_component46_fa11_or0;
  wire [0:0] csa_component46_fa12_xor1;
  wire [0:0] csa_component46_fa12_or0;
  wire [0:0] csa_component46_fa13_xor1;
  wire [0:0] csa_component46_fa13_or0;
  wire [0:0] csa_component46_fa14_xor1;
  wire [0:0] csa_component46_fa14_or0;
  wire [0:0] csa_component46_fa15_xor1;
  wire [0:0] csa_component46_fa15_or0;
  wire [0:0] csa_component46_fa16_xor1;
  wire [0:0] csa_component46_fa16_or0;
  wire [0:0] csa_component46_fa17_xor1;
  wire [0:0] csa_component46_fa17_or0;
  wire [0:0] csa_component46_fa18_xor1;
  wire [0:0] csa_component46_fa18_or0;
  wire [0:0] csa_component46_fa19_xor1;
  wire [0:0] csa_component46_fa19_or0;
  wire [0:0] csa_component46_fa20_xor1;
  wire [0:0] csa_component46_fa20_or0;
  wire [0:0] csa_component46_fa21_xor1;
  wire [0:0] csa_component46_fa21_or0;
  wire [0:0] csa_component46_fa22_xor1;
  wire [0:0] csa_component46_fa22_or0;
  wire [0:0] csa_component46_fa23_xor1;
  wire [0:0] csa_component46_fa23_or0;
  wire [0:0] csa_component46_fa24_xor1;
  wire [0:0] csa_component46_fa24_or0;
  wire [0:0] csa_component46_fa25_xor1;
  wire [0:0] csa_component46_fa25_or0;
  wire [0:0] csa_component46_fa26_xor1;
  wire [0:0] csa_component46_fa26_or0;
  wire [0:0] csa_component46_fa27_xor1;
  wire [0:0] csa_component46_fa27_or0;
  wire [0:0] csa_component46_fa28_xor1;
  wire [0:0] csa_component46_fa28_or0;
  wire [0:0] csa_component46_fa29_xor1;
  wire [0:0] csa_component46_fa29_or0;
  wire [0:0] csa_component46_fa30_xor1;
  wire [0:0] csa_component46_fa30_or0;
  wire [0:0] csa_component46_fa31_xor1;
  wire [0:0] csa_component46_fa31_or0;
  wire [0:0] csa_component46_fa32_xor1;
  wire [0:0] csa_component46_fa32_or0;
  wire [0:0] csa_component46_fa33_xor1;
  wire [0:0] csa_component46_fa33_or0;
  wire [0:0] csa_component46_fa34_xor1;
  wire [0:0] csa_component46_fa34_or0;
  wire [0:0] csa_component46_fa35_xor1;
  wire [0:0] csa_component46_fa35_or0;
  wire [0:0] csa_component46_fa36_xor1;
  wire [0:0] csa_component46_fa36_or0;
  wire [0:0] csa_component46_fa37_xor1;
  wire [0:0] csa_component46_fa37_or0;
  wire [0:0] csa_component46_fa38_xor1;
  wire [0:0] csa_component46_fa38_or0;
  wire [0:0] csa_component46_fa39_xor1;
  wire [0:0] csa_component46_fa39_or0;
  wire [0:0] csa_component46_fa40_xor1;
  wire [0:0] csa_component46_fa40_or0;
  wire [0:0] csa_component46_fa41_xor1;
  wire [0:0] csa_component46_fa41_or0;
  wire [0:0] csa_component46_fa42_xor1;
  wire [0:0] csa_component46_fa42_or0;
  wire [0:0] csa_component46_fa43_xor1;
  wire [0:0] csa_component46_fa43_or0;
  wire [0:0] csa_component46_fa44_xor1;
  wire [0:0] csa_component46_fa44_or0;
  wire [0:0] csa_component46_fa45_xor1;
  wire [0:0] csa_component46_fa45_or0;

  fa fa_csa_component46_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component46_fa0_xor1), .fa_or0(csa_component46_fa0_or0));
  fa fa_csa_component46_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component46_fa1_xor1), .fa_or0(csa_component46_fa1_or0));
  fa fa_csa_component46_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component46_fa2_xor1), .fa_or0(csa_component46_fa2_or0));
  fa fa_csa_component46_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component46_fa3_xor1), .fa_or0(csa_component46_fa3_or0));
  fa fa_csa_component46_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component46_fa4_xor1), .fa_or0(csa_component46_fa4_or0));
  fa fa_csa_component46_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component46_fa5_xor1), .fa_or0(csa_component46_fa5_or0));
  fa fa_csa_component46_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component46_fa6_xor1), .fa_or0(csa_component46_fa6_or0));
  fa fa_csa_component46_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component46_fa7_xor1), .fa_or0(csa_component46_fa7_or0));
  fa fa_csa_component46_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component46_fa8_xor1), .fa_or0(csa_component46_fa8_or0));
  fa fa_csa_component46_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component46_fa9_xor1), .fa_or0(csa_component46_fa9_or0));
  fa fa_csa_component46_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component46_fa10_xor1), .fa_or0(csa_component46_fa10_or0));
  fa fa_csa_component46_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component46_fa11_xor1), .fa_or0(csa_component46_fa11_or0));
  fa fa_csa_component46_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component46_fa12_xor1), .fa_or0(csa_component46_fa12_or0));
  fa fa_csa_component46_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component46_fa13_xor1), .fa_or0(csa_component46_fa13_or0));
  fa fa_csa_component46_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component46_fa14_xor1), .fa_or0(csa_component46_fa14_or0));
  fa fa_csa_component46_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component46_fa15_xor1), .fa_or0(csa_component46_fa15_or0));
  fa fa_csa_component46_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component46_fa16_xor1), .fa_or0(csa_component46_fa16_or0));
  fa fa_csa_component46_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component46_fa17_xor1), .fa_or0(csa_component46_fa17_or0));
  fa fa_csa_component46_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component46_fa18_xor1), .fa_or0(csa_component46_fa18_or0));
  fa fa_csa_component46_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component46_fa19_xor1), .fa_or0(csa_component46_fa19_or0));
  fa fa_csa_component46_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component46_fa20_xor1), .fa_or0(csa_component46_fa20_or0));
  fa fa_csa_component46_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component46_fa21_xor1), .fa_or0(csa_component46_fa21_or0));
  fa fa_csa_component46_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component46_fa22_xor1), .fa_or0(csa_component46_fa22_or0));
  fa fa_csa_component46_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component46_fa23_xor1), .fa_or0(csa_component46_fa23_or0));
  fa fa_csa_component46_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component46_fa24_xor1), .fa_or0(csa_component46_fa24_or0));
  fa fa_csa_component46_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component46_fa25_xor1), .fa_or0(csa_component46_fa25_or0));
  fa fa_csa_component46_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component46_fa26_xor1), .fa_or0(csa_component46_fa26_or0));
  fa fa_csa_component46_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component46_fa27_xor1), .fa_or0(csa_component46_fa27_or0));
  fa fa_csa_component46_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component46_fa28_xor1), .fa_or0(csa_component46_fa28_or0));
  fa fa_csa_component46_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component46_fa29_xor1), .fa_or0(csa_component46_fa29_or0));
  fa fa_csa_component46_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component46_fa30_xor1), .fa_or0(csa_component46_fa30_or0));
  fa fa_csa_component46_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component46_fa31_xor1), .fa_or0(csa_component46_fa31_or0));
  fa fa_csa_component46_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component46_fa32_xor1), .fa_or0(csa_component46_fa32_or0));
  fa fa_csa_component46_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component46_fa33_xor1), .fa_or0(csa_component46_fa33_or0));
  fa fa_csa_component46_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component46_fa34_xor1), .fa_or0(csa_component46_fa34_or0));
  fa fa_csa_component46_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component46_fa35_xor1), .fa_or0(csa_component46_fa35_or0));
  fa fa_csa_component46_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component46_fa36_xor1), .fa_or0(csa_component46_fa36_or0));
  fa fa_csa_component46_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component46_fa37_xor1), .fa_or0(csa_component46_fa37_or0));
  fa fa_csa_component46_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component46_fa38_xor1), .fa_or0(csa_component46_fa38_or0));
  fa fa_csa_component46_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component46_fa39_xor1), .fa_or0(csa_component46_fa39_or0));
  fa fa_csa_component46_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component46_fa40_xor1), .fa_or0(csa_component46_fa40_or0));
  fa fa_csa_component46_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component46_fa41_xor1), .fa_or0(csa_component46_fa41_or0));
  fa fa_csa_component46_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component46_fa42_xor1), .fa_or0(csa_component46_fa42_or0));
  fa fa_csa_component46_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component46_fa43_xor1), .fa_or0(csa_component46_fa43_or0));
  fa fa_csa_component46_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component46_fa44_xor1), .fa_or0(csa_component46_fa44_or0));
  fa fa_csa_component46_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component46_fa45_xor1), .fa_or0(csa_component46_fa45_or0));

  assign csa_component46_out[0] = csa_component46_fa0_xor1[0];
  assign csa_component46_out[1] = csa_component46_fa1_xor1[0];
  assign csa_component46_out[2] = csa_component46_fa2_xor1[0];
  assign csa_component46_out[3] = csa_component46_fa3_xor1[0];
  assign csa_component46_out[4] = csa_component46_fa4_xor1[0];
  assign csa_component46_out[5] = csa_component46_fa5_xor1[0];
  assign csa_component46_out[6] = csa_component46_fa6_xor1[0];
  assign csa_component46_out[7] = csa_component46_fa7_xor1[0];
  assign csa_component46_out[8] = csa_component46_fa8_xor1[0];
  assign csa_component46_out[9] = csa_component46_fa9_xor1[0];
  assign csa_component46_out[10] = csa_component46_fa10_xor1[0];
  assign csa_component46_out[11] = csa_component46_fa11_xor1[0];
  assign csa_component46_out[12] = csa_component46_fa12_xor1[0];
  assign csa_component46_out[13] = csa_component46_fa13_xor1[0];
  assign csa_component46_out[14] = csa_component46_fa14_xor1[0];
  assign csa_component46_out[15] = csa_component46_fa15_xor1[0];
  assign csa_component46_out[16] = csa_component46_fa16_xor1[0];
  assign csa_component46_out[17] = csa_component46_fa17_xor1[0];
  assign csa_component46_out[18] = csa_component46_fa18_xor1[0];
  assign csa_component46_out[19] = csa_component46_fa19_xor1[0];
  assign csa_component46_out[20] = csa_component46_fa20_xor1[0];
  assign csa_component46_out[21] = csa_component46_fa21_xor1[0];
  assign csa_component46_out[22] = csa_component46_fa22_xor1[0];
  assign csa_component46_out[23] = csa_component46_fa23_xor1[0];
  assign csa_component46_out[24] = csa_component46_fa24_xor1[0];
  assign csa_component46_out[25] = csa_component46_fa25_xor1[0];
  assign csa_component46_out[26] = csa_component46_fa26_xor1[0];
  assign csa_component46_out[27] = csa_component46_fa27_xor1[0];
  assign csa_component46_out[28] = csa_component46_fa28_xor1[0];
  assign csa_component46_out[29] = csa_component46_fa29_xor1[0];
  assign csa_component46_out[30] = csa_component46_fa30_xor1[0];
  assign csa_component46_out[31] = csa_component46_fa31_xor1[0];
  assign csa_component46_out[32] = csa_component46_fa32_xor1[0];
  assign csa_component46_out[33] = csa_component46_fa33_xor1[0];
  assign csa_component46_out[34] = csa_component46_fa34_xor1[0];
  assign csa_component46_out[35] = csa_component46_fa35_xor1[0];
  assign csa_component46_out[36] = csa_component46_fa36_xor1[0];
  assign csa_component46_out[37] = csa_component46_fa37_xor1[0];
  assign csa_component46_out[38] = csa_component46_fa38_xor1[0];
  assign csa_component46_out[39] = csa_component46_fa39_xor1[0];
  assign csa_component46_out[40] = csa_component46_fa40_xor1[0];
  assign csa_component46_out[41] = csa_component46_fa41_xor1[0];
  assign csa_component46_out[42] = csa_component46_fa42_xor1[0];
  assign csa_component46_out[43] = csa_component46_fa43_xor1[0];
  assign csa_component46_out[44] = csa_component46_fa44_xor1[0];
  assign csa_component46_out[45] = csa_component46_fa45_xor1[0];
  assign csa_component46_out[46] = 1'b0;
  assign csa_component46_out[47] = 1'b0;
  assign csa_component46_out[48] = csa_component46_fa0_or0[0];
  assign csa_component46_out[49] = csa_component46_fa1_or0[0];
  assign csa_component46_out[50] = csa_component46_fa2_or0[0];
  assign csa_component46_out[51] = csa_component46_fa3_or0[0];
  assign csa_component46_out[52] = csa_component46_fa4_or0[0];
  assign csa_component46_out[53] = csa_component46_fa5_or0[0];
  assign csa_component46_out[54] = csa_component46_fa6_or0[0];
  assign csa_component46_out[55] = csa_component46_fa7_or0[0];
  assign csa_component46_out[56] = csa_component46_fa8_or0[0];
  assign csa_component46_out[57] = csa_component46_fa9_or0[0];
  assign csa_component46_out[58] = csa_component46_fa10_or0[0];
  assign csa_component46_out[59] = csa_component46_fa11_or0[0];
  assign csa_component46_out[60] = csa_component46_fa12_or0[0];
  assign csa_component46_out[61] = csa_component46_fa13_or0[0];
  assign csa_component46_out[62] = csa_component46_fa14_or0[0];
  assign csa_component46_out[63] = csa_component46_fa15_or0[0];
  assign csa_component46_out[64] = csa_component46_fa16_or0[0];
  assign csa_component46_out[65] = csa_component46_fa17_or0[0];
  assign csa_component46_out[66] = csa_component46_fa18_or0[0];
  assign csa_component46_out[67] = csa_component46_fa19_or0[0];
  assign csa_component46_out[68] = csa_component46_fa20_or0[0];
  assign csa_component46_out[69] = csa_component46_fa21_or0[0];
  assign csa_component46_out[70] = csa_component46_fa22_or0[0];
  assign csa_component46_out[71] = csa_component46_fa23_or0[0];
  assign csa_component46_out[72] = csa_component46_fa24_or0[0];
  assign csa_component46_out[73] = csa_component46_fa25_or0[0];
  assign csa_component46_out[74] = csa_component46_fa26_or0[0];
  assign csa_component46_out[75] = csa_component46_fa27_or0[0];
  assign csa_component46_out[76] = csa_component46_fa28_or0[0];
  assign csa_component46_out[77] = csa_component46_fa29_or0[0];
  assign csa_component46_out[78] = csa_component46_fa30_or0[0];
  assign csa_component46_out[79] = csa_component46_fa31_or0[0];
  assign csa_component46_out[80] = csa_component46_fa32_or0[0];
  assign csa_component46_out[81] = csa_component46_fa33_or0[0];
  assign csa_component46_out[82] = csa_component46_fa34_or0[0];
  assign csa_component46_out[83] = csa_component46_fa35_or0[0];
  assign csa_component46_out[84] = csa_component46_fa36_or0[0];
  assign csa_component46_out[85] = csa_component46_fa37_or0[0];
  assign csa_component46_out[86] = csa_component46_fa38_or0[0];
  assign csa_component46_out[87] = csa_component46_fa39_or0[0];
  assign csa_component46_out[88] = csa_component46_fa40_or0[0];
  assign csa_component46_out[89] = csa_component46_fa41_or0[0];
  assign csa_component46_out[90] = csa_component46_fa42_or0[0];
  assign csa_component46_out[91] = csa_component46_fa43_or0[0];
  assign csa_component46_out[92] = csa_component46_fa44_or0[0];
  assign csa_component46_out[93] = csa_component46_fa45_or0[0];
endmodule

module csa_component49(input [48:0] a, input [48:0] b, input [48:0] c, output [99:0] csa_component49_out);
  wire [0:0] csa_component49_fa0_xor1;
  wire [0:0] csa_component49_fa0_or0;
  wire [0:0] csa_component49_fa1_xor1;
  wire [0:0] csa_component49_fa1_or0;
  wire [0:0] csa_component49_fa2_xor1;
  wire [0:0] csa_component49_fa2_or0;
  wire [0:0] csa_component49_fa3_xor1;
  wire [0:0] csa_component49_fa3_or0;
  wire [0:0] csa_component49_fa4_xor1;
  wire [0:0] csa_component49_fa4_or0;
  wire [0:0] csa_component49_fa5_xor1;
  wire [0:0] csa_component49_fa5_or0;
  wire [0:0] csa_component49_fa6_xor1;
  wire [0:0] csa_component49_fa6_or0;
  wire [0:0] csa_component49_fa7_xor1;
  wire [0:0] csa_component49_fa7_or0;
  wire [0:0] csa_component49_fa8_xor1;
  wire [0:0] csa_component49_fa8_or0;
  wire [0:0] csa_component49_fa9_xor1;
  wire [0:0] csa_component49_fa9_or0;
  wire [0:0] csa_component49_fa10_xor1;
  wire [0:0] csa_component49_fa10_or0;
  wire [0:0] csa_component49_fa11_xor1;
  wire [0:0] csa_component49_fa11_or0;
  wire [0:0] csa_component49_fa12_xor1;
  wire [0:0] csa_component49_fa12_or0;
  wire [0:0] csa_component49_fa13_xor1;
  wire [0:0] csa_component49_fa13_or0;
  wire [0:0] csa_component49_fa14_xor1;
  wire [0:0] csa_component49_fa14_or0;
  wire [0:0] csa_component49_fa15_xor1;
  wire [0:0] csa_component49_fa15_or0;
  wire [0:0] csa_component49_fa16_xor1;
  wire [0:0] csa_component49_fa16_or0;
  wire [0:0] csa_component49_fa17_xor1;
  wire [0:0] csa_component49_fa17_or0;
  wire [0:0] csa_component49_fa18_xor1;
  wire [0:0] csa_component49_fa18_or0;
  wire [0:0] csa_component49_fa19_xor1;
  wire [0:0] csa_component49_fa19_or0;
  wire [0:0] csa_component49_fa20_xor1;
  wire [0:0] csa_component49_fa20_or0;
  wire [0:0] csa_component49_fa21_xor1;
  wire [0:0] csa_component49_fa21_or0;
  wire [0:0] csa_component49_fa22_xor1;
  wire [0:0] csa_component49_fa22_or0;
  wire [0:0] csa_component49_fa23_xor1;
  wire [0:0] csa_component49_fa23_or0;
  wire [0:0] csa_component49_fa24_xor1;
  wire [0:0] csa_component49_fa24_or0;
  wire [0:0] csa_component49_fa25_xor1;
  wire [0:0] csa_component49_fa25_or0;
  wire [0:0] csa_component49_fa26_xor1;
  wire [0:0] csa_component49_fa26_or0;
  wire [0:0] csa_component49_fa27_xor1;
  wire [0:0] csa_component49_fa27_or0;
  wire [0:0] csa_component49_fa28_xor1;
  wire [0:0] csa_component49_fa28_or0;
  wire [0:0] csa_component49_fa29_xor1;
  wire [0:0] csa_component49_fa29_or0;
  wire [0:0] csa_component49_fa30_xor1;
  wire [0:0] csa_component49_fa30_or0;
  wire [0:0] csa_component49_fa31_xor1;
  wire [0:0] csa_component49_fa31_or0;
  wire [0:0] csa_component49_fa32_xor1;
  wire [0:0] csa_component49_fa32_or0;
  wire [0:0] csa_component49_fa33_xor1;
  wire [0:0] csa_component49_fa33_or0;
  wire [0:0] csa_component49_fa34_xor1;
  wire [0:0] csa_component49_fa34_or0;
  wire [0:0] csa_component49_fa35_xor1;
  wire [0:0] csa_component49_fa35_or0;
  wire [0:0] csa_component49_fa36_xor1;
  wire [0:0] csa_component49_fa36_or0;
  wire [0:0] csa_component49_fa37_xor1;
  wire [0:0] csa_component49_fa37_or0;
  wire [0:0] csa_component49_fa38_xor1;
  wire [0:0] csa_component49_fa38_or0;
  wire [0:0] csa_component49_fa39_xor1;
  wire [0:0] csa_component49_fa39_or0;
  wire [0:0] csa_component49_fa40_xor1;
  wire [0:0] csa_component49_fa40_or0;
  wire [0:0] csa_component49_fa41_xor1;
  wire [0:0] csa_component49_fa41_or0;
  wire [0:0] csa_component49_fa42_xor1;
  wire [0:0] csa_component49_fa42_or0;
  wire [0:0] csa_component49_fa43_xor1;
  wire [0:0] csa_component49_fa43_or0;
  wire [0:0] csa_component49_fa44_xor1;
  wire [0:0] csa_component49_fa44_or0;
  wire [0:0] csa_component49_fa45_xor1;
  wire [0:0] csa_component49_fa45_or0;
  wire [0:0] csa_component49_fa46_xor1;
  wire [0:0] csa_component49_fa46_or0;
  wire [0:0] csa_component49_fa47_xor1;
  wire [0:0] csa_component49_fa47_or0;
  wire [0:0] csa_component49_fa48_xor1;
  wire [0:0] csa_component49_fa48_or0;

  fa fa_csa_component49_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component49_fa0_xor1), .fa_or0(csa_component49_fa0_or0));
  fa fa_csa_component49_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component49_fa1_xor1), .fa_or0(csa_component49_fa1_or0));
  fa fa_csa_component49_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component49_fa2_xor1), .fa_or0(csa_component49_fa2_or0));
  fa fa_csa_component49_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component49_fa3_xor1), .fa_or0(csa_component49_fa3_or0));
  fa fa_csa_component49_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component49_fa4_xor1), .fa_or0(csa_component49_fa4_or0));
  fa fa_csa_component49_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component49_fa5_xor1), .fa_or0(csa_component49_fa5_or0));
  fa fa_csa_component49_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component49_fa6_xor1), .fa_or0(csa_component49_fa6_or0));
  fa fa_csa_component49_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component49_fa7_xor1), .fa_or0(csa_component49_fa7_or0));
  fa fa_csa_component49_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component49_fa8_xor1), .fa_or0(csa_component49_fa8_or0));
  fa fa_csa_component49_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component49_fa9_xor1), .fa_or0(csa_component49_fa9_or0));
  fa fa_csa_component49_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component49_fa10_xor1), .fa_or0(csa_component49_fa10_or0));
  fa fa_csa_component49_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component49_fa11_xor1), .fa_or0(csa_component49_fa11_or0));
  fa fa_csa_component49_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component49_fa12_xor1), .fa_or0(csa_component49_fa12_or0));
  fa fa_csa_component49_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component49_fa13_xor1), .fa_or0(csa_component49_fa13_or0));
  fa fa_csa_component49_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component49_fa14_xor1), .fa_or0(csa_component49_fa14_or0));
  fa fa_csa_component49_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component49_fa15_xor1), .fa_or0(csa_component49_fa15_or0));
  fa fa_csa_component49_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component49_fa16_xor1), .fa_or0(csa_component49_fa16_or0));
  fa fa_csa_component49_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component49_fa17_xor1), .fa_or0(csa_component49_fa17_or0));
  fa fa_csa_component49_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component49_fa18_xor1), .fa_or0(csa_component49_fa18_or0));
  fa fa_csa_component49_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component49_fa19_xor1), .fa_or0(csa_component49_fa19_or0));
  fa fa_csa_component49_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component49_fa20_xor1), .fa_or0(csa_component49_fa20_or0));
  fa fa_csa_component49_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component49_fa21_xor1), .fa_or0(csa_component49_fa21_or0));
  fa fa_csa_component49_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component49_fa22_xor1), .fa_or0(csa_component49_fa22_or0));
  fa fa_csa_component49_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component49_fa23_xor1), .fa_or0(csa_component49_fa23_or0));
  fa fa_csa_component49_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component49_fa24_xor1), .fa_or0(csa_component49_fa24_or0));
  fa fa_csa_component49_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component49_fa25_xor1), .fa_or0(csa_component49_fa25_or0));
  fa fa_csa_component49_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component49_fa26_xor1), .fa_or0(csa_component49_fa26_or0));
  fa fa_csa_component49_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component49_fa27_xor1), .fa_or0(csa_component49_fa27_or0));
  fa fa_csa_component49_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component49_fa28_xor1), .fa_or0(csa_component49_fa28_or0));
  fa fa_csa_component49_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component49_fa29_xor1), .fa_or0(csa_component49_fa29_or0));
  fa fa_csa_component49_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component49_fa30_xor1), .fa_or0(csa_component49_fa30_or0));
  fa fa_csa_component49_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component49_fa31_xor1), .fa_or0(csa_component49_fa31_or0));
  fa fa_csa_component49_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component49_fa32_xor1), .fa_or0(csa_component49_fa32_or0));
  fa fa_csa_component49_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component49_fa33_xor1), .fa_or0(csa_component49_fa33_or0));
  fa fa_csa_component49_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component49_fa34_xor1), .fa_or0(csa_component49_fa34_or0));
  fa fa_csa_component49_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component49_fa35_xor1), .fa_or0(csa_component49_fa35_or0));
  fa fa_csa_component49_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component49_fa36_xor1), .fa_or0(csa_component49_fa36_or0));
  fa fa_csa_component49_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component49_fa37_xor1), .fa_or0(csa_component49_fa37_or0));
  fa fa_csa_component49_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component49_fa38_xor1), .fa_or0(csa_component49_fa38_or0));
  fa fa_csa_component49_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component49_fa39_xor1), .fa_or0(csa_component49_fa39_or0));
  fa fa_csa_component49_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component49_fa40_xor1), .fa_or0(csa_component49_fa40_or0));
  fa fa_csa_component49_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component49_fa41_xor1), .fa_or0(csa_component49_fa41_or0));
  fa fa_csa_component49_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component49_fa42_xor1), .fa_or0(csa_component49_fa42_or0));
  fa fa_csa_component49_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component49_fa43_xor1), .fa_or0(csa_component49_fa43_or0));
  fa fa_csa_component49_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component49_fa44_xor1), .fa_or0(csa_component49_fa44_or0));
  fa fa_csa_component49_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component49_fa45_xor1), .fa_or0(csa_component49_fa45_or0));
  fa fa_csa_component49_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component49_fa46_xor1), .fa_or0(csa_component49_fa46_or0));
  fa fa_csa_component49_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component49_fa47_xor1), .fa_or0(csa_component49_fa47_or0));
  fa fa_csa_component49_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component49_fa48_xor1), .fa_or0(csa_component49_fa48_or0));

  assign csa_component49_out[0] = csa_component49_fa0_xor1[0];
  assign csa_component49_out[1] = csa_component49_fa1_xor1[0];
  assign csa_component49_out[2] = csa_component49_fa2_xor1[0];
  assign csa_component49_out[3] = csa_component49_fa3_xor1[0];
  assign csa_component49_out[4] = csa_component49_fa4_xor1[0];
  assign csa_component49_out[5] = csa_component49_fa5_xor1[0];
  assign csa_component49_out[6] = csa_component49_fa6_xor1[0];
  assign csa_component49_out[7] = csa_component49_fa7_xor1[0];
  assign csa_component49_out[8] = csa_component49_fa8_xor1[0];
  assign csa_component49_out[9] = csa_component49_fa9_xor1[0];
  assign csa_component49_out[10] = csa_component49_fa10_xor1[0];
  assign csa_component49_out[11] = csa_component49_fa11_xor1[0];
  assign csa_component49_out[12] = csa_component49_fa12_xor1[0];
  assign csa_component49_out[13] = csa_component49_fa13_xor1[0];
  assign csa_component49_out[14] = csa_component49_fa14_xor1[0];
  assign csa_component49_out[15] = csa_component49_fa15_xor1[0];
  assign csa_component49_out[16] = csa_component49_fa16_xor1[0];
  assign csa_component49_out[17] = csa_component49_fa17_xor1[0];
  assign csa_component49_out[18] = csa_component49_fa18_xor1[0];
  assign csa_component49_out[19] = csa_component49_fa19_xor1[0];
  assign csa_component49_out[20] = csa_component49_fa20_xor1[0];
  assign csa_component49_out[21] = csa_component49_fa21_xor1[0];
  assign csa_component49_out[22] = csa_component49_fa22_xor1[0];
  assign csa_component49_out[23] = csa_component49_fa23_xor1[0];
  assign csa_component49_out[24] = csa_component49_fa24_xor1[0];
  assign csa_component49_out[25] = csa_component49_fa25_xor1[0];
  assign csa_component49_out[26] = csa_component49_fa26_xor1[0];
  assign csa_component49_out[27] = csa_component49_fa27_xor1[0];
  assign csa_component49_out[28] = csa_component49_fa28_xor1[0];
  assign csa_component49_out[29] = csa_component49_fa29_xor1[0];
  assign csa_component49_out[30] = csa_component49_fa30_xor1[0];
  assign csa_component49_out[31] = csa_component49_fa31_xor1[0];
  assign csa_component49_out[32] = csa_component49_fa32_xor1[0];
  assign csa_component49_out[33] = csa_component49_fa33_xor1[0];
  assign csa_component49_out[34] = csa_component49_fa34_xor1[0];
  assign csa_component49_out[35] = csa_component49_fa35_xor1[0];
  assign csa_component49_out[36] = csa_component49_fa36_xor1[0];
  assign csa_component49_out[37] = csa_component49_fa37_xor1[0];
  assign csa_component49_out[38] = csa_component49_fa38_xor1[0];
  assign csa_component49_out[39] = csa_component49_fa39_xor1[0];
  assign csa_component49_out[40] = csa_component49_fa40_xor1[0];
  assign csa_component49_out[41] = csa_component49_fa41_xor1[0];
  assign csa_component49_out[42] = csa_component49_fa42_xor1[0];
  assign csa_component49_out[43] = csa_component49_fa43_xor1[0];
  assign csa_component49_out[44] = csa_component49_fa44_xor1[0];
  assign csa_component49_out[45] = csa_component49_fa45_xor1[0];
  assign csa_component49_out[46] = csa_component49_fa46_xor1[0];
  assign csa_component49_out[47] = csa_component49_fa47_xor1[0];
  assign csa_component49_out[48] = csa_component49_fa48_xor1[0];
  assign csa_component49_out[49] = 1'b0;
  assign csa_component49_out[50] = 1'b0;
  assign csa_component49_out[51] = csa_component49_fa0_or0[0];
  assign csa_component49_out[52] = csa_component49_fa1_or0[0];
  assign csa_component49_out[53] = csa_component49_fa2_or0[0];
  assign csa_component49_out[54] = csa_component49_fa3_or0[0];
  assign csa_component49_out[55] = csa_component49_fa4_or0[0];
  assign csa_component49_out[56] = csa_component49_fa5_or0[0];
  assign csa_component49_out[57] = csa_component49_fa6_or0[0];
  assign csa_component49_out[58] = csa_component49_fa7_or0[0];
  assign csa_component49_out[59] = csa_component49_fa8_or0[0];
  assign csa_component49_out[60] = csa_component49_fa9_or0[0];
  assign csa_component49_out[61] = csa_component49_fa10_or0[0];
  assign csa_component49_out[62] = csa_component49_fa11_or0[0];
  assign csa_component49_out[63] = csa_component49_fa12_or0[0];
  assign csa_component49_out[64] = csa_component49_fa13_or0[0];
  assign csa_component49_out[65] = csa_component49_fa14_or0[0];
  assign csa_component49_out[66] = csa_component49_fa15_or0[0];
  assign csa_component49_out[67] = csa_component49_fa16_or0[0];
  assign csa_component49_out[68] = csa_component49_fa17_or0[0];
  assign csa_component49_out[69] = csa_component49_fa18_or0[0];
  assign csa_component49_out[70] = csa_component49_fa19_or0[0];
  assign csa_component49_out[71] = csa_component49_fa20_or0[0];
  assign csa_component49_out[72] = csa_component49_fa21_or0[0];
  assign csa_component49_out[73] = csa_component49_fa22_or0[0];
  assign csa_component49_out[74] = csa_component49_fa23_or0[0];
  assign csa_component49_out[75] = csa_component49_fa24_or0[0];
  assign csa_component49_out[76] = csa_component49_fa25_or0[0];
  assign csa_component49_out[77] = csa_component49_fa26_or0[0];
  assign csa_component49_out[78] = csa_component49_fa27_or0[0];
  assign csa_component49_out[79] = csa_component49_fa28_or0[0];
  assign csa_component49_out[80] = csa_component49_fa29_or0[0];
  assign csa_component49_out[81] = csa_component49_fa30_or0[0];
  assign csa_component49_out[82] = csa_component49_fa31_or0[0];
  assign csa_component49_out[83] = csa_component49_fa32_or0[0];
  assign csa_component49_out[84] = csa_component49_fa33_or0[0];
  assign csa_component49_out[85] = csa_component49_fa34_or0[0];
  assign csa_component49_out[86] = csa_component49_fa35_or0[0];
  assign csa_component49_out[87] = csa_component49_fa36_or0[0];
  assign csa_component49_out[88] = csa_component49_fa37_or0[0];
  assign csa_component49_out[89] = csa_component49_fa38_or0[0];
  assign csa_component49_out[90] = csa_component49_fa39_or0[0];
  assign csa_component49_out[91] = csa_component49_fa40_or0[0];
  assign csa_component49_out[92] = csa_component49_fa41_or0[0];
  assign csa_component49_out[93] = csa_component49_fa42_or0[0];
  assign csa_component49_out[94] = csa_component49_fa43_or0[0];
  assign csa_component49_out[95] = csa_component49_fa44_or0[0];
  assign csa_component49_out[96] = csa_component49_fa45_or0[0];
  assign csa_component49_out[97] = csa_component49_fa46_or0[0];
  assign csa_component49_out[98] = csa_component49_fa47_or0[0];
  assign csa_component49_out[99] = csa_component49_fa48_or0[0];
endmodule

module csa_component52(input [51:0] a, input [51:0] b, input [51:0] c, output [105:0] csa_component52_out);
  wire [0:0] csa_component52_fa0_xor1;
  wire [0:0] csa_component52_fa0_or0;
  wire [0:0] csa_component52_fa1_xor1;
  wire [0:0] csa_component52_fa1_or0;
  wire [0:0] csa_component52_fa2_xor1;
  wire [0:0] csa_component52_fa2_or0;
  wire [0:0] csa_component52_fa3_xor1;
  wire [0:0] csa_component52_fa3_or0;
  wire [0:0] csa_component52_fa4_xor1;
  wire [0:0] csa_component52_fa4_or0;
  wire [0:0] csa_component52_fa5_xor1;
  wire [0:0] csa_component52_fa5_or0;
  wire [0:0] csa_component52_fa6_xor1;
  wire [0:0] csa_component52_fa6_or0;
  wire [0:0] csa_component52_fa7_xor1;
  wire [0:0] csa_component52_fa7_or0;
  wire [0:0] csa_component52_fa8_xor1;
  wire [0:0] csa_component52_fa8_or0;
  wire [0:0] csa_component52_fa9_xor1;
  wire [0:0] csa_component52_fa9_or0;
  wire [0:0] csa_component52_fa10_xor1;
  wire [0:0] csa_component52_fa10_or0;
  wire [0:0] csa_component52_fa11_xor1;
  wire [0:0] csa_component52_fa11_or0;
  wire [0:0] csa_component52_fa12_xor1;
  wire [0:0] csa_component52_fa12_or0;
  wire [0:0] csa_component52_fa13_xor1;
  wire [0:0] csa_component52_fa13_or0;
  wire [0:0] csa_component52_fa14_xor1;
  wire [0:0] csa_component52_fa14_or0;
  wire [0:0] csa_component52_fa15_xor1;
  wire [0:0] csa_component52_fa15_or0;
  wire [0:0] csa_component52_fa16_xor1;
  wire [0:0] csa_component52_fa16_or0;
  wire [0:0] csa_component52_fa17_xor1;
  wire [0:0] csa_component52_fa17_or0;
  wire [0:0] csa_component52_fa18_xor1;
  wire [0:0] csa_component52_fa18_or0;
  wire [0:0] csa_component52_fa19_xor1;
  wire [0:0] csa_component52_fa19_or0;
  wire [0:0] csa_component52_fa20_xor1;
  wire [0:0] csa_component52_fa20_or0;
  wire [0:0] csa_component52_fa21_xor1;
  wire [0:0] csa_component52_fa21_or0;
  wire [0:0] csa_component52_fa22_xor1;
  wire [0:0] csa_component52_fa22_or0;
  wire [0:0] csa_component52_fa23_xor1;
  wire [0:0] csa_component52_fa23_or0;
  wire [0:0] csa_component52_fa24_xor1;
  wire [0:0] csa_component52_fa24_or0;
  wire [0:0] csa_component52_fa25_xor1;
  wire [0:0] csa_component52_fa25_or0;
  wire [0:0] csa_component52_fa26_xor1;
  wire [0:0] csa_component52_fa26_or0;
  wire [0:0] csa_component52_fa27_xor1;
  wire [0:0] csa_component52_fa27_or0;
  wire [0:0] csa_component52_fa28_xor1;
  wire [0:0] csa_component52_fa28_or0;
  wire [0:0] csa_component52_fa29_xor1;
  wire [0:0] csa_component52_fa29_or0;
  wire [0:0] csa_component52_fa30_xor1;
  wire [0:0] csa_component52_fa30_or0;
  wire [0:0] csa_component52_fa31_xor1;
  wire [0:0] csa_component52_fa31_or0;
  wire [0:0] csa_component52_fa32_xor1;
  wire [0:0] csa_component52_fa32_or0;
  wire [0:0] csa_component52_fa33_xor1;
  wire [0:0] csa_component52_fa33_or0;
  wire [0:0] csa_component52_fa34_xor1;
  wire [0:0] csa_component52_fa34_or0;
  wire [0:0] csa_component52_fa35_xor1;
  wire [0:0] csa_component52_fa35_or0;
  wire [0:0] csa_component52_fa36_xor1;
  wire [0:0] csa_component52_fa36_or0;
  wire [0:0] csa_component52_fa37_xor1;
  wire [0:0] csa_component52_fa37_or0;
  wire [0:0] csa_component52_fa38_xor1;
  wire [0:0] csa_component52_fa38_or0;
  wire [0:0] csa_component52_fa39_xor1;
  wire [0:0] csa_component52_fa39_or0;
  wire [0:0] csa_component52_fa40_xor1;
  wire [0:0] csa_component52_fa40_or0;
  wire [0:0] csa_component52_fa41_xor1;
  wire [0:0] csa_component52_fa41_or0;
  wire [0:0] csa_component52_fa42_xor1;
  wire [0:0] csa_component52_fa42_or0;
  wire [0:0] csa_component52_fa43_xor1;
  wire [0:0] csa_component52_fa43_or0;
  wire [0:0] csa_component52_fa44_xor1;
  wire [0:0] csa_component52_fa44_or0;
  wire [0:0] csa_component52_fa45_xor1;
  wire [0:0] csa_component52_fa45_or0;
  wire [0:0] csa_component52_fa46_xor1;
  wire [0:0] csa_component52_fa46_or0;
  wire [0:0] csa_component52_fa47_xor1;
  wire [0:0] csa_component52_fa47_or0;
  wire [0:0] csa_component52_fa48_xor1;
  wire [0:0] csa_component52_fa48_or0;
  wire [0:0] csa_component52_fa49_xor1;
  wire [0:0] csa_component52_fa49_or0;
  wire [0:0] csa_component52_fa50_xor1;
  wire [0:0] csa_component52_fa50_or0;
  wire [0:0] csa_component52_fa51_xor1;
  wire [0:0] csa_component52_fa51_or0;

  fa fa_csa_component52_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component52_fa0_xor1), .fa_or0(csa_component52_fa0_or0));
  fa fa_csa_component52_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component52_fa1_xor1), .fa_or0(csa_component52_fa1_or0));
  fa fa_csa_component52_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component52_fa2_xor1), .fa_or0(csa_component52_fa2_or0));
  fa fa_csa_component52_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component52_fa3_xor1), .fa_or0(csa_component52_fa3_or0));
  fa fa_csa_component52_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component52_fa4_xor1), .fa_or0(csa_component52_fa4_or0));
  fa fa_csa_component52_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component52_fa5_xor1), .fa_or0(csa_component52_fa5_or0));
  fa fa_csa_component52_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component52_fa6_xor1), .fa_or0(csa_component52_fa6_or0));
  fa fa_csa_component52_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component52_fa7_xor1), .fa_or0(csa_component52_fa7_or0));
  fa fa_csa_component52_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component52_fa8_xor1), .fa_or0(csa_component52_fa8_or0));
  fa fa_csa_component52_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component52_fa9_xor1), .fa_or0(csa_component52_fa9_or0));
  fa fa_csa_component52_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component52_fa10_xor1), .fa_or0(csa_component52_fa10_or0));
  fa fa_csa_component52_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component52_fa11_xor1), .fa_or0(csa_component52_fa11_or0));
  fa fa_csa_component52_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component52_fa12_xor1), .fa_or0(csa_component52_fa12_or0));
  fa fa_csa_component52_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component52_fa13_xor1), .fa_or0(csa_component52_fa13_or0));
  fa fa_csa_component52_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component52_fa14_xor1), .fa_or0(csa_component52_fa14_or0));
  fa fa_csa_component52_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component52_fa15_xor1), .fa_or0(csa_component52_fa15_or0));
  fa fa_csa_component52_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component52_fa16_xor1), .fa_or0(csa_component52_fa16_or0));
  fa fa_csa_component52_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component52_fa17_xor1), .fa_or0(csa_component52_fa17_or0));
  fa fa_csa_component52_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component52_fa18_xor1), .fa_or0(csa_component52_fa18_or0));
  fa fa_csa_component52_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component52_fa19_xor1), .fa_or0(csa_component52_fa19_or0));
  fa fa_csa_component52_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component52_fa20_xor1), .fa_or0(csa_component52_fa20_or0));
  fa fa_csa_component52_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component52_fa21_xor1), .fa_or0(csa_component52_fa21_or0));
  fa fa_csa_component52_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component52_fa22_xor1), .fa_or0(csa_component52_fa22_or0));
  fa fa_csa_component52_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component52_fa23_xor1), .fa_or0(csa_component52_fa23_or0));
  fa fa_csa_component52_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component52_fa24_xor1), .fa_or0(csa_component52_fa24_or0));
  fa fa_csa_component52_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component52_fa25_xor1), .fa_or0(csa_component52_fa25_or0));
  fa fa_csa_component52_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component52_fa26_xor1), .fa_or0(csa_component52_fa26_or0));
  fa fa_csa_component52_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component52_fa27_xor1), .fa_or0(csa_component52_fa27_or0));
  fa fa_csa_component52_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component52_fa28_xor1), .fa_or0(csa_component52_fa28_or0));
  fa fa_csa_component52_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component52_fa29_xor1), .fa_or0(csa_component52_fa29_or0));
  fa fa_csa_component52_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component52_fa30_xor1), .fa_or0(csa_component52_fa30_or0));
  fa fa_csa_component52_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component52_fa31_xor1), .fa_or0(csa_component52_fa31_or0));
  fa fa_csa_component52_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component52_fa32_xor1), .fa_or0(csa_component52_fa32_or0));
  fa fa_csa_component52_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component52_fa33_xor1), .fa_or0(csa_component52_fa33_or0));
  fa fa_csa_component52_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component52_fa34_xor1), .fa_or0(csa_component52_fa34_or0));
  fa fa_csa_component52_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component52_fa35_xor1), .fa_or0(csa_component52_fa35_or0));
  fa fa_csa_component52_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component52_fa36_xor1), .fa_or0(csa_component52_fa36_or0));
  fa fa_csa_component52_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component52_fa37_xor1), .fa_or0(csa_component52_fa37_or0));
  fa fa_csa_component52_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component52_fa38_xor1), .fa_or0(csa_component52_fa38_or0));
  fa fa_csa_component52_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component52_fa39_xor1), .fa_or0(csa_component52_fa39_or0));
  fa fa_csa_component52_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component52_fa40_xor1), .fa_or0(csa_component52_fa40_or0));
  fa fa_csa_component52_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component52_fa41_xor1), .fa_or0(csa_component52_fa41_or0));
  fa fa_csa_component52_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component52_fa42_xor1), .fa_or0(csa_component52_fa42_or0));
  fa fa_csa_component52_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component52_fa43_xor1), .fa_or0(csa_component52_fa43_or0));
  fa fa_csa_component52_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component52_fa44_xor1), .fa_or0(csa_component52_fa44_or0));
  fa fa_csa_component52_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component52_fa45_xor1), .fa_or0(csa_component52_fa45_or0));
  fa fa_csa_component52_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component52_fa46_xor1), .fa_or0(csa_component52_fa46_or0));
  fa fa_csa_component52_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component52_fa47_xor1), .fa_or0(csa_component52_fa47_or0));
  fa fa_csa_component52_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component52_fa48_xor1), .fa_or0(csa_component52_fa48_or0));
  fa fa_csa_component52_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component52_fa49_xor1), .fa_or0(csa_component52_fa49_or0));
  fa fa_csa_component52_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component52_fa50_xor1), .fa_or0(csa_component52_fa50_or0));
  fa fa_csa_component52_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component52_fa51_xor1), .fa_or0(csa_component52_fa51_or0));

  assign csa_component52_out[0] = csa_component52_fa0_xor1[0];
  assign csa_component52_out[1] = csa_component52_fa1_xor1[0];
  assign csa_component52_out[2] = csa_component52_fa2_xor1[0];
  assign csa_component52_out[3] = csa_component52_fa3_xor1[0];
  assign csa_component52_out[4] = csa_component52_fa4_xor1[0];
  assign csa_component52_out[5] = csa_component52_fa5_xor1[0];
  assign csa_component52_out[6] = csa_component52_fa6_xor1[0];
  assign csa_component52_out[7] = csa_component52_fa7_xor1[0];
  assign csa_component52_out[8] = csa_component52_fa8_xor1[0];
  assign csa_component52_out[9] = csa_component52_fa9_xor1[0];
  assign csa_component52_out[10] = csa_component52_fa10_xor1[0];
  assign csa_component52_out[11] = csa_component52_fa11_xor1[0];
  assign csa_component52_out[12] = csa_component52_fa12_xor1[0];
  assign csa_component52_out[13] = csa_component52_fa13_xor1[0];
  assign csa_component52_out[14] = csa_component52_fa14_xor1[0];
  assign csa_component52_out[15] = csa_component52_fa15_xor1[0];
  assign csa_component52_out[16] = csa_component52_fa16_xor1[0];
  assign csa_component52_out[17] = csa_component52_fa17_xor1[0];
  assign csa_component52_out[18] = csa_component52_fa18_xor1[0];
  assign csa_component52_out[19] = csa_component52_fa19_xor1[0];
  assign csa_component52_out[20] = csa_component52_fa20_xor1[0];
  assign csa_component52_out[21] = csa_component52_fa21_xor1[0];
  assign csa_component52_out[22] = csa_component52_fa22_xor1[0];
  assign csa_component52_out[23] = csa_component52_fa23_xor1[0];
  assign csa_component52_out[24] = csa_component52_fa24_xor1[0];
  assign csa_component52_out[25] = csa_component52_fa25_xor1[0];
  assign csa_component52_out[26] = csa_component52_fa26_xor1[0];
  assign csa_component52_out[27] = csa_component52_fa27_xor1[0];
  assign csa_component52_out[28] = csa_component52_fa28_xor1[0];
  assign csa_component52_out[29] = csa_component52_fa29_xor1[0];
  assign csa_component52_out[30] = csa_component52_fa30_xor1[0];
  assign csa_component52_out[31] = csa_component52_fa31_xor1[0];
  assign csa_component52_out[32] = csa_component52_fa32_xor1[0];
  assign csa_component52_out[33] = csa_component52_fa33_xor1[0];
  assign csa_component52_out[34] = csa_component52_fa34_xor1[0];
  assign csa_component52_out[35] = csa_component52_fa35_xor1[0];
  assign csa_component52_out[36] = csa_component52_fa36_xor1[0];
  assign csa_component52_out[37] = csa_component52_fa37_xor1[0];
  assign csa_component52_out[38] = csa_component52_fa38_xor1[0];
  assign csa_component52_out[39] = csa_component52_fa39_xor1[0];
  assign csa_component52_out[40] = csa_component52_fa40_xor1[0];
  assign csa_component52_out[41] = csa_component52_fa41_xor1[0];
  assign csa_component52_out[42] = csa_component52_fa42_xor1[0];
  assign csa_component52_out[43] = csa_component52_fa43_xor1[0];
  assign csa_component52_out[44] = csa_component52_fa44_xor1[0];
  assign csa_component52_out[45] = csa_component52_fa45_xor1[0];
  assign csa_component52_out[46] = csa_component52_fa46_xor1[0];
  assign csa_component52_out[47] = csa_component52_fa47_xor1[0];
  assign csa_component52_out[48] = csa_component52_fa48_xor1[0];
  assign csa_component52_out[49] = csa_component52_fa49_xor1[0];
  assign csa_component52_out[50] = csa_component52_fa50_xor1[0];
  assign csa_component52_out[51] = csa_component52_fa51_xor1[0];
  assign csa_component52_out[52] = 1'b0;
  assign csa_component52_out[53] = 1'b0;
  assign csa_component52_out[54] = csa_component52_fa0_or0[0];
  assign csa_component52_out[55] = csa_component52_fa1_or0[0];
  assign csa_component52_out[56] = csa_component52_fa2_or0[0];
  assign csa_component52_out[57] = csa_component52_fa3_or0[0];
  assign csa_component52_out[58] = csa_component52_fa4_or0[0];
  assign csa_component52_out[59] = csa_component52_fa5_or0[0];
  assign csa_component52_out[60] = csa_component52_fa6_or0[0];
  assign csa_component52_out[61] = csa_component52_fa7_or0[0];
  assign csa_component52_out[62] = csa_component52_fa8_or0[0];
  assign csa_component52_out[63] = csa_component52_fa9_or0[0];
  assign csa_component52_out[64] = csa_component52_fa10_or0[0];
  assign csa_component52_out[65] = csa_component52_fa11_or0[0];
  assign csa_component52_out[66] = csa_component52_fa12_or0[0];
  assign csa_component52_out[67] = csa_component52_fa13_or0[0];
  assign csa_component52_out[68] = csa_component52_fa14_or0[0];
  assign csa_component52_out[69] = csa_component52_fa15_or0[0];
  assign csa_component52_out[70] = csa_component52_fa16_or0[0];
  assign csa_component52_out[71] = csa_component52_fa17_or0[0];
  assign csa_component52_out[72] = csa_component52_fa18_or0[0];
  assign csa_component52_out[73] = csa_component52_fa19_or0[0];
  assign csa_component52_out[74] = csa_component52_fa20_or0[0];
  assign csa_component52_out[75] = csa_component52_fa21_or0[0];
  assign csa_component52_out[76] = csa_component52_fa22_or0[0];
  assign csa_component52_out[77] = csa_component52_fa23_or0[0];
  assign csa_component52_out[78] = csa_component52_fa24_or0[0];
  assign csa_component52_out[79] = csa_component52_fa25_or0[0];
  assign csa_component52_out[80] = csa_component52_fa26_or0[0];
  assign csa_component52_out[81] = csa_component52_fa27_or0[0];
  assign csa_component52_out[82] = csa_component52_fa28_or0[0];
  assign csa_component52_out[83] = csa_component52_fa29_or0[0];
  assign csa_component52_out[84] = csa_component52_fa30_or0[0];
  assign csa_component52_out[85] = csa_component52_fa31_or0[0];
  assign csa_component52_out[86] = csa_component52_fa32_or0[0];
  assign csa_component52_out[87] = csa_component52_fa33_or0[0];
  assign csa_component52_out[88] = csa_component52_fa34_or0[0];
  assign csa_component52_out[89] = csa_component52_fa35_or0[0];
  assign csa_component52_out[90] = csa_component52_fa36_or0[0];
  assign csa_component52_out[91] = csa_component52_fa37_or0[0];
  assign csa_component52_out[92] = csa_component52_fa38_or0[0];
  assign csa_component52_out[93] = csa_component52_fa39_or0[0];
  assign csa_component52_out[94] = csa_component52_fa40_or0[0];
  assign csa_component52_out[95] = csa_component52_fa41_or0[0];
  assign csa_component52_out[96] = csa_component52_fa42_or0[0];
  assign csa_component52_out[97] = csa_component52_fa43_or0[0];
  assign csa_component52_out[98] = csa_component52_fa44_or0[0];
  assign csa_component52_out[99] = csa_component52_fa45_or0[0];
  assign csa_component52_out[100] = csa_component52_fa46_or0[0];
  assign csa_component52_out[101] = csa_component52_fa47_or0[0];
  assign csa_component52_out[102] = csa_component52_fa48_or0[0];
  assign csa_component52_out[103] = csa_component52_fa49_or0[0];
  assign csa_component52_out[104] = csa_component52_fa50_or0[0];
  assign csa_component52_out[105] = csa_component52_fa51_or0[0];
endmodule

module csa_component55(input [54:0] a, input [54:0] b, input [54:0] c, output [111:0] csa_component55_out);
  wire [0:0] csa_component55_fa0_xor1;
  wire [0:0] csa_component55_fa0_or0;
  wire [0:0] csa_component55_fa1_xor1;
  wire [0:0] csa_component55_fa1_or0;
  wire [0:0] csa_component55_fa2_xor1;
  wire [0:0] csa_component55_fa2_or0;
  wire [0:0] csa_component55_fa3_xor1;
  wire [0:0] csa_component55_fa3_or0;
  wire [0:0] csa_component55_fa4_xor1;
  wire [0:0] csa_component55_fa4_or0;
  wire [0:0] csa_component55_fa5_xor1;
  wire [0:0] csa_component55_fa5_or0;
  wire [0:0] csa_component55_fa6_xor1;
  wire [0:0] csa_component55_fa6_or0;
  wire [0:0] csa_component55_fa7_xor1;
  wire [0:0] csa_component55_fa7_or0;
  wire [0:0] csa_component55_fa8_xor1;
  wire [0:0] csa_component55_fa8_or0;
  wire [0:0] csa_component55_fa9_xor1;
  wire [0:0] csa_component55_fa9_or0;
  wire [0:0] csa_component55_fa10_xor1;
  wire [0:0] csa_component55_fa10_or0;
  wire [0:0] csa_component55_fa11_xor1;
  wire [0:0] csa_component55_fa11_or0;
  wire [0:0] csa_component55_fa12_xor1;
  wire [0:0] csa_component55_fa12_or0;
  wire [0:0] csa_component55_fa13_xor1;
  wire [0:0] csa_component55_fa13_or0;
  wire [0:0] csa_component55_fa14_xor1;
  wire [0:0] csa_component55_fa14_or0;
  wire [0:0] csa_component55_fa15_xor1;
  wire [0:0] csa_component55_fa15_or0;
  wire [0:0] csa_component55_fa16_xor1;
  wire [0:0] csa_component55_fa16_or0;
  wire [0:0] csa_component55_fa17_xor1;
  wire [0:0] csa_component55_fa17_or0;
  wire [0:0] csa_component55_fa18_xor1;
  wire [0:0] csa_component55_fa18_or0;
  wire [0:0] csa_component55_fa19_xor1;
  wire [0:0] csa_component55_fa19_or0;
  wire [0:0] csa_component55_fa20_xor1;
  wire [0:0] csa_component55_fa20_or0;
  wire [0:0] csa_component55_fa21_xor1;
  wire [0:0] csa_component55_fa21_or0;
  wire [0:0] csa_component55_fa22_xor1;
  wire [0:0] csa_component55_fa22_or0;
  wire [0:0] csa_component55_fa23_xor1;
  wire [0:0] csa_component55_fa23_or0;
  wire [0:0] csa_component55_fa24_xor1;
  wire [0:0] csa_component55_fa24_or0;
  wire [0:0] csa_component55_fa25_xor1;
  wire [0:0] csa_component55_fa25_or0;
  wire [0:0] csa_component55_fa26_xor1;
  wire [0:0] csa_component55_fa26_or0;
  wire [0:0] csa_component55_fa27_xor1;
  wire [0:0] csa_component55_fa27_or0;
  wire [0:0] csa_component55_fa28_xor1;
  wire [0:0] csa_component55_fa28_or0;
  wire [0:0] csa_component55_fa29_xor1;
  wire [0:0] csa_component55_fa29_or0;
  wire [0:0] csa_component55_fa30_xor1;
  wire [0:0] csa_component55_fa30_or0;
  wire [0:0] csa_component55_fa31_xor1;
  wire [0:0] csa_component55_fa31_or0;
  wire [0:0] csa_component55_fa32_xor1;
  wire [0:0] csa_component55_fa32_or0;
  wire [0:0] csa_component55_fa33_xor1;
  wire [0:0] csa_component55_fa33_or0;
  wire [0:0] csa_component55_fa34_xor1;
  wire [0:0] csa_component55_fa34_or0;
  wire [0:0] csa_component55_fa35_xor1;
  wire [0:0] csa_component55_fa35_or0;
  wire [0:0] csa_component55_fa36_xor1;
  wire [0:0] csa_component55_fa36_or0;
  wire [0:0] csa_component55_fa37_xor1;
  wire [0:0] csa_component55_fa37_or0;
  wire [0:0] csa_component55_fa38_xor1;
  wire [0:0] csa_component55_fa38_or0;
  wire [0:0] csa_component55_fa39_xor1;
  wire [0:0] csa_component55_fa39_or0;
  wire [0:0] csa_component55_fa40_xor1;
  wire [0:0] csa_component55_fa40_or0;
  wire [0:0] csa_component55_fa41_xor1;
  wire [0:0] csa_component55_fa41_or0;
  wire [0:0] csa_component55_fa42_xor1;
  wire [0:0] csa_component55_fa42_or0;
  wire [0:0] csa_component55_fa43_xor1;
  wire [0:0] csa_component55_fa43_or0;
  wire [0:0] csa_component55_fa44_xor1;
  wire [0:0] csa_component55_fa44_or0;
  wire [0:0] csa_component55_fa45_xor1;
  wire [0:0] csa_component55_fa45_or0;
  wire [0:0] csa_component55_fa46_xor1;
  wire [0:0] csa_component55_fa46_or0;
  wire [0:0] csa_component55_fa47_xor1;
  wire [0:0] csa_component55_fa47_or0;
  wire [0:0] csa_component55_fa48_xor1;
  wire [0:0] csa_component55_fa48_or0;
  wire [0:0] csa_component55_fa49_xor1;
  wire [0:0] csa_component55_fa49_or0;
  wire [0:0] csa_component55_fa50_xor1;
  wire [0:0] csa_component55_fa50_or0;
  wire [0:0] csa_component55_fa51_xor1;
  wire [0:0] csa_component55_fa51_or0;
  wire [0:0] csa_component55_fa52_xor1;
  wire [0:0] csa_component55_fa52_or0;
  wire [0:0] csa_component55_fa53_xor1;
  wire [0:0] csa_component55_fa53_or0;
  wire [0:0] csa_component55_fa54_xor1;
  wire [0:0] csa_component55_fa54_or0;

  fa fa_csa_component55_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component55_fa0_xor1), .fa_or0(csa_component55_fa0_or0));
  fa fa_csa_component55_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component55_fa1_xor1), .fa_or0(csa_component55_fa1_or0));
  fa fa_csa_component55_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component55_fa2_xor1), .fa_or0(csa_component55_fa2_or0));
  fa fa_csa_component55_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component55_fa3_xor1), .fa_or0(csa_component55_fa3_or0));
  fa fa_csa_component55_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component55_fa4_xor1), .fa_or0(csa_component55_fa4_or0));
  fa fa_csa_component55_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component55_fa5_xor1), .fa_or0(csa_component55_fa5_or0));
  fa fa_csa_component55_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component55_fa6_xor1), .fa_or0(csa_component55_fa6_or0));
  fa fa_csa_component55_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component55_fa7_xor1), .fa_or0(csa_component55_fa7_or0));
  fa fa_csa_component55_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component55_fa8_xor1), .fa_or0(csa_component55_fa8_or0));
  fa fa_csa_component55_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component55_fa9_xor1), .fa_or0(csa_component55_fa9_or0));
  fa fa_csa_component55_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component55_fa10_xor1), .fa_or0(csa_component55_fa10_or0));
  fa fa_csa_component55_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component55_fa11_xor1), .fa_or0(csa_component55_fa11_or0));
  fa fa_csa_component55_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component55_fa12_xor1), .fa_or0(csa_component55_fa12_or0));
  fa fa_csa_component55_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component55_fa13_xor1), .fa_or0(csa_component55_fa13_or0));
  fa fa_csa_component55_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component55_fa14_xor1), .fa_or0(csa_component55_fa14_or0));
  fa fa_csa_component55_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component55_fa15_xor1), .fa_or0(csa_component55_fa15_or0));
  fa fa_csa_component55_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component55_fa16_xor1), .fa_or0(csa_component55_fa16_or0));
  fa fa_csa_component55_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component55_fa17_xor1), .fa_or0(csa_component55_fa17_or0));
  fa fa_csa_component55_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component55_fa18_xor1), .fa_or0(csa_component55_fa18_or0));
  fa fa_csa_component55_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component55_fa19_xor1), .fa_or0(csa_component55_fa19_or0));
  fa fa_csa_component55_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component55_fa20_xor1), .fa_or0(csa_component55_fa20_or0));
  fa fa_csa_component55_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component55_fa21_xor1), .fa_or0(csa_component55_fa21_or0));
  fa fa_csa_component55_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component55_fa22_xor1), .fa_or0(csa_component55_fa22_or0));
  fa fa_csa_component55_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component55_fa23_xor1), .fa_or0(csa_component55_fa23_or0));
  fa fa_csa_component55_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component55_fa24_xor1), .fa_or0(csa_component55_fa24_or0));
  fa fa_csa_component55_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component55_fa25_xor1), .fa_or0(csa_component55_fa25_or0));
  fa fa_csa_component55_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component55_fa26_xor1), .fa_or0(csa_component55_fa26_or0));
  fa fa_csa_component55_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component55_fa27_xor1), .fa_or0(csa_component55_fa27_or0));
  fa fa_csa_component55_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component55_fa28_xor1), .fa_or0(csa_component55_fa28_or0));
  fa fa_csa_component55_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component55_fa29_xor1), .fa_or0(csa_component55_fa29_or0));
  fa fa_csa_component55_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component55_fa30_xor1), .fa_or0(csa_component55_fa30_or0));
  fa fa_csa_component55_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component55_fa31_xor1), .fa_or0(csa_component55_fa31_or0));
  fa fa_csa_component55_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component55_fa32_xor1), .fa_or0(csa_component55_fa32_or0));
  fa fa_csa_component55_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component55_fa33_xor1), .fa_or0(csa_component55_fa33_or0));
  fa fa_csa_component55_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component55_fa34_xor1), .fa_or0(csa_component55_fa34_or0));
  fa fa_csa_component55_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component55_fa35_xor1), .fa_or0(csa_component55_fa35_or0));
  fa fa_csa_component55_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component55_fa36_xor1), .fa_or0(csa_component55_fa36_or0));
  fa fa_csa_component55_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component55_fa37_xor1), .fa_or0(csa_component55_fa37_or0));
  fa fa_csa_component55_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component55_fa38_xor1), .fa_or0(csa_component55_fa38_or0));
  fa fa_csa_component55_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component55_fa39_xor1), .fa_or0(csa_component55_fa39_or0));
  fa fa_csa_component55_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component55_fa40_xor1), .fa_or0(csa_component55_fa40_or0));
  fa fa_csa_component55_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component55_fa41_xor1), .fa_or0(csa_component55_fa41_or0));
  fa fa_csa_component55_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component55_fa42_xor1), .fa_or0(csa_component55_fa42_or0));
  fa fa_csa_component55_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component55_fa43_xor1), .fa_or0(csa_component55_fa43_or0));
  fa fa_csa_component55_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component55_fa44_xor1), .fa_or0(csa_component55_fa44_or0));
  fa fa_csa_component55_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component55_fa45_xor1), .fa_or0(csa_component55_fa45_or0));
  fa fa_csa_component55_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component55_fa46_xor1), .fa_or0(csa_component55_fa46_or0));
  fa fa_csa_component55_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component55_fa47_xor1), .fa_or0(csa_component55_fa47_or0));
  fa fa_csa_component55_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component55_fa48_xor1), .fa_or0(csa_component55_fa48_or0));
  fa fa_csa_component55_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component55_fa49_xor1), .fa_or0(csa_component55_fa49_or0));
  fa fa_csa_component55_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component55_fa50_xor1), .fa_or0(csa_component55_fa50_or0));
  fa fa_csa_component55_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component55_fa51_xor1), .fa_or0(csa_component55_fa51_or0));
  fa fa_csa_component55_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component55_fa52_xor1), .fa_or0(csa_component55_fa52_or0));
  fa fa_csa_component55_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component55_fa53_xor1), .fa_or0(csa_component55_fa53_or0));
  fa fa_csa_component55_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component55_fa54_xor1), .fa_or0(csa_component55_fa54_or0));

  assign csa_component55_out[0] = csa_component55_fa0_xor1[0];
  assign csa_component55_out[1] = csa_component55_fa1_xor1[0];
  assign csa_component55_out[2] = csa_component55_fa2_xor1[0];
  assign csa_component55_out[3] = csa_component55_fa3_xor1[0];
  assign csa_component55_out[4] = csa_component55_fa4_xor1[0];
  assign csa_component55_out[5] = csa_component55_fa5_xor1[0];
  assign csa_component55_out[6] = csa_component55_fa6_xor1[0];
  assign csa_component55_out[7] = csa_component55_fa7_xor1[0];
  assign csa_component55_out[8] = csa_component55_fa8_xor1[0];
  assign csa_component55_out[9] = csa_component55_fa9_xor1[0];
  assign csa_component55_out[10] = csa_component55_fa10_xor1[0];
  assign csa_component55_out[11] = csa_component55_fa11_xor1[0];
  assign csa_component55_out[12] = csa_component55_fa12_xor1[0];
  assign csa_component55_out[13] = csa_component55_fa13_xor1[0];
  assign csa_component55_out[14] = csa_component55_fa14_xor1[0];
  assign csa_component55_out[15] = csa_component55_fa15_xor1[0];
  assign csa_component55_out[16] = csa_component55_fa16_xor1[0];
  assign csa_component55_out[17] = csa_component55_fa17_xor1[0];
  assign csa_component55_out[18] = csa_component55_fa18_xor1[0];
  assign csa_component55_out[19] = csa_component55_fa19_xor1[0];
  assign csa_component55_out[20] = csa_component55_fa20_xor1[0];
  assign csa_component55_out[21] = csa_component55_fa21_xor1[0];
  assign csa_component55_out[22] = csa_component55_fa22_xor1[0];
  assign csa_component55_out[23] = csa_component55_fa23_xor1[0];
  assign csa_component55_out[24] = csa_component55_fa24_xor1[0];
  assign csa_component55_out[25] = csa_component55_fa25_xor1[0];
  assign csa_component55_out[26] = csa_component55_fa26_xor1[0];
  assign csa_component55_out[27] = csa_component55_fa27_xor1[0];
  assign csa_component55_out[28] = csa_component55_fa28_xor1[0];
  assign csa_component55_out[29] = csa_component55_fa29_xor1[0];
  assign csa_component55_out[30] = csa_component55_fa30_xor1[0];
  assign csa_component55_out[31] = csa_component55_fa31_xor1[0];
  assign csa_component55_out[32] = csa_component55_fa32_xor1[0];
  assign csa_component55_out[33] = csa_component55_fa33_xor1[0];
  assign csa_component55_out[34] = csa_component55_fa34_xor1[0];
  assign csa_component55_out[35] = csa_component55_fa35_xor1[0];
  assign csa_component55_out[36] = csa_component55_fa36_xor1[0];
  assign csa_component55_out[37] = csa_component55_fa37_xor1[0];
  assign csa_component55_out[38] = csa_component55_fa38_xor1[0];
  assign csa_component55_out[39] = csa_component55_fa39_xor1[0];
  assign csa_component55_out[40] = csa_component55_fa40_xor1[0];
  assign csa_component55_out[41] = csa_component55_fa41_xor1[0];
  assign csa_component55_out[42] = csa_component55_fa42_xor1[0];
  assign csa_component55_out[43] = csa_component55_fa43_xor1[0];
  assign csa_component55_out[44] = csa_component55_fa44_xor1[0];
  assign csa_component55_out[45] = csa_component55_fa45_xor1[0];
  assign csa_component55_out[46] = csa_component55_fa46_xor1[0];
  assign csa_component55_out[47] = csa_component55_fa47_xor1[0];
  assign csa_component55_out[48] = csa_component55_fa48_xor1[0];
  assign csa_component55_out[49] = csa_component55_fa49_xor1[0];
  assign csa_component55_out[50] = csa_component55_fa50_xor1[0];
  assign csa_component55_out[51] = csa_component55_fa51_xor1[0];
  assign csa_component55_out[52] = csa_component55_fa52_xor1[0];
  assign csa_component55_out[53] = csa_component55_fa53_xor1[0];
  assign csa_component55_out[54] = csa_component55_fa54_xor1[0];
  assign csa_component55_out[55] = 1'b0;
  assign csa_component55_out[56] = 1'b0;
  assign csa_component55_out[57] = csa_component55_fa0_or0[0];
  assign csa_component55_out[58] = csa_component55_fa1_or0[0];
  assign csa_component55_out[59] = csa_component55_fa2_or0[0];
  assign csa_component55_out[60] = csa_component55_fa3_or0[0];
  assign csa_component55_out[61] = csa_component55_fa4_or0[0];
  assign csa_component55_out[62] = csa_component55_fa5_or0[0];
  assign csa_component55_out[63] = csa_component55_fa6_or0[0];
  assign csa_component55_out[64] = csa_component55_fa7_or0[0];
  assign csa_component55_out[65] = csa_component55_fa8_or0[0];
  assign csa_component55_out[66] = csa_component55_fa9_or0[0];
  assign csa_component55_out[67] = csa_component55_fa10_or0[0];
  assign csa_component55_out[68] = csa_component55_fa11_or0[0];
  assign csa_component55_out[69] = csa_component55_fa12_or0[0];
  assign csa_component55_out[70] = csa_component55_fa13_or0[0];
  assign csa_component55_out[71] = csa_component55_fa14_or0[0];
  assign csa_component55_out[72] = csa_component55_fa15_or0[0];
  assign csa_component55_out[73] = csa_component55_fa16_or0[0];
  assign csa_component55_out[74] = csa_component55_fa17_or0[0];
  assign csa_component55_out[75] = csa_component55_fa18_or0[0];
  assign csa_component55_out[76] = csa_component55_fa19_or0[0];
  assign csa_component55_out[77] = csa_component55_fa20_or0[0];
  assign csa_component55_out[78] = csa_component55_fa21_or0[0];
  assign csa_component55_out[79] = csa_component55_fa22_or0[0];
  assign csa_component55_out[80] = csa_component55_fa23_or0[0];
  assign csa_component55_out[81] = csa_component55_fa24_or0[0];
  assign csa_component55_out[82] = csa_component55_fa25_or0[0];
  assign csa_component55_out[83] = csa_component55_fa26_or0[0];
  assign csa_component55_out[84] = csa_component55_fa27_or0[0];
  assign csa_component55_out[85] = csa_component55_fa28_or0[0];
  assign csa_component55_out[86] = csa_component55_fa29_or0[0];
  assign csa_component55_out[87] = csa_component55_fa30_or0[0];
  assign csa_component55_out[88] = csa_component55_fa31_or0[0];
  assign csa_component55_out[89] = csa_component55_fa32_or0[0];
  assign csa_component55_out[90] = csa_component55_fa33_or0[0];
  assign csa_component55_out[91] = csa_component55_fa34_or0[0];
  assign csa_component55_out[92] = csa_component55_fa35_or0[0];
  assign csa_component55_out[93] = csa_component55_fa36_or0[0];
  assign csa_component55_out[94] = csa_component55_fa37_or0[0];
  assign csa_component55_out[95] = csa_component55_fa38_or0[0];
  assign csa_component55_out[96] = csa_component55_fa39_or0[0];
  assign csa_component55_out[97] = csa_component55_fa40_or0[0];
  assign csa_component55_out[98] = csa_component55_fa41_or0[0];
  assign csa_component55_out[99] = csa_component55_fa42_or0[0];
  assign csa_component55_out[100] = csa_component55_fa43_or0[0];
  assign csa_component55_out[101] = csa_component55_fa44_or0[0];
  assign csa_component55_out[102] = csa_component55_fa45_or0[0];
  assign csa_component55_out[103] = csa_component55_fa46_or0[0];
  assign csa_component55_out[104] = csa_component55_fa47_or0[0];
  assign csa_component55_out[105] = csa_component55_fa48_or0[0];
  assign csa_component55_out[106] = csa_component55_fa49_or0[0];
  assign csa_component55_out[107] = csa_component55_fa50_or0[0];
  assign csa_component55_out[108] = csa_component55_fa51_or0[0];
  assign csa_component55_out[109] = csa_component55_fa52_or0[0];
  assign csa_component55_out[110] = csa_component55_fa53_or0[0];
  assign csa_component55_out[111] = csa_component55_fa54_or0[0];
endmodule

module csa_component58(input [57:0] a, input [57:0] b, input [57:0] c, output [117:0] csa_component58_out);
  wire [0:0] csa_component58_fa0_xor1;
  wire [0:0] csa_component58_fa0_or0;
  wire [0:0] csa_component58_fa1_xor1;
  wire [0:0] csa_component58_fa1_or0;
  wire [0:0] csa_component58_fa2_xor1;
  wire [0:0] csa_component58_fa2_or0;
  wire [0:0] csa_component58_fa3_xor1;
  wire [0:0] csa_component58_fa3_or0;
  wire [0:0] csa_component58_fa4_xor1;
  wire [0:0] csa_component58_fa4_or0;
  wire [0:0] csa_component58_fa5_xor1;
  wire [0:0] csa_component58_fa5_or0;
  wire [0:0] csa_component58_fa6_xor1;
  wire [0:0] csa_component58_fa6_or0;
  wire [0:0] csa_component58_fa7_xor1;
  wire [0:0] csa_component58_fa7_or0;
  wire [0:0] csa_component58_fa8_xor1;
  wire [0:0] csa_component58_fa8_or0;
  wire [0:0] csa_component58_fa9_xor1;
  wire [0:0] csa_component58_fa9_or0;
  wire [0:0] csa_component58_fa10_xor1;
  wire [0:0] csa_component58_fa10_or0;
  wire [0:0] csa_component58_fa11_xor1;
  wire [0:0] csa_component58_fa11_or0;
  wire [0:0] csa_component58_fa12_xor1;
  wire [0:0] csa_component58_fa12_or0;
  wire [0:0] csa_component58_fa13_xor1;
  wire [0:0] csa_component58_fa13_or0;
  wire [0:0] csa_component58_fa14_xor1;
  wire [0:0] csa_component58_fa14_or0;
  wire [0:0] csa_component58_fa15_xor1;
  wire [0:0] csa_component58_fa15_or0;
  wire [0:0] csa_component58_fa16_xor1;
  wire [0:0] csa_component58_fa16_or0;
  wire [0:0] csa_component58_fa17_xor1;
  wire [0:0] csa_component58_fa17_or0;
  wire [0:0] csa_component58_fa18_xor1;
  wire [0:0] csa_component58_fa18_or0;
  wire [0:0] csa_component58_fa19_xor1;
  wire [0:0] csa_component58_fa19_or0;
  wire [0:0] csa_component58_fa20_xor1;
  wire [0:0] csa_component58_fa20_or0;
  wire [0:0] csa_component58_fa21_xor1;
  wire [0:0] csa_component58_fa21_or0;
  wire [0:0] csa_component58_fa22_xor1;
  wire [0:0] csa_component58_fa22_or0;
  wire [0:0] csa_component58_fa23_xor1;
  wire [0:0] csa_component58_fa23_or0;
  wire [0:0] csa_component58_fa24_xor1;
  wire [0:0] csa_component58_fa24_or0;
  wire [0:0] csa_component58_fa25_xor1;
  wire [0:0] csa_component58_fa25_or0;
  wire [0:0] csa_component58_fa26_xor1;
  wire [0:0] csa_component58_fa26_or0;
  wire [0:0] csa_component58_fa27_xor1;
  wire [0:0] csa_component58_fa27_or0;
  wire [0:0] csa_component58_fa28_xor1;
  wire [0:0] csa_component58_fa28_or0;
  wire [0:0] csa_component58_fa29_xor1;
  wire [0:0] csa_component58_fa29_or0;
  wire [0:0] csa_component58_fa30_xor1;
  wire [0:0] csa_component58_fa30_or0;
  wire [0:0] csa_component58_fa31_xor1;
  wire [0:0] csa_component58_fa31_or0;
  wire [0:0] csa_component58_fa32_xor1;
  wire [0:0] csa_component58_fa32_or0;
  wire [0:0] csa_component58_fa33_xor1;
  wire [0:0] csa_component58_fa33_or0;
  wire [0:0] csa_component58_fa34_xor1;
  wire [0:0] csa_component58_fa34_or0;
  wire [0:0] csa_component58_fa35_xor1;
  wire [0:0] csa_component58_fa35_or0;
  wire [0:0] csa_component58_fa36_xor1;
  wire [0:0] csa_component58_fa36_or0;
  wire [0:0] csa_component58_fa37_xor1;
  wire [0:0] csa_component58_fa37_or0;
  wire [0:0] csa_component58_fa38_xor1;
  wire [0:0] csa_component58_fa38_or0;
  wire [0:0] csa_component58_fa39_xor1;
  wire [0:0] csa_component58_fa39_or0;
  wire [0:0] csa_component58_fa40_xor1;
  wire [0:0] csa_component58_fa40_or0;
  wire [0:0] csa_component58_fa41_xor1;
  wire [0:0] csa_component58_fa41_or0;
  wire [0:0] csa_component58_fa42_xor1;
  wire [0:0] csa_component58_fa42_or0;
  wire [0:0] csa_component58_fa43_xor1;
  wire [0:0] csa_component58_fa43_or0;
  wire [0:0] csa_component58_fa44_xor1;
  wire [0:0] csa_component58_fa44_or0;
  wire [0:0] csa_component58_fa45_xor1;
  wire [0:0] csa_component58_fa45_or0;
  wire [0:0] csa_component58_fa46_xor1;
  wire [0:0] csa_component58_fa46_or0;
  wire [0:0] csa_component58_fa47_xor1;
  wire [0:0] csa_component58_fa47_or0;
  wire [0:0] csa_component58_fa48_xor1;
  wire [0:0] csa_component58_fa48_or0;
  wire [0:0] csa_component58_fa49_xor1;
  wire [0:0] csa_component58_fa49_or0;
  wire [0:0] csa_component58_fa50_xor1;
  wire [0:0] csa_component58_fa50_or0;
  wire [0:0] csa_component58_fa51_xor1;
  wire [0:0] csa_component58_fa51_or0;
  wire [0:0] csa_component58_fa52_xor1;
  wire [0:0] csa_component58_fa52_or0;
  wire [0:0] csa_component58_fa53_xor1;
  wire [0:0] csa_component58_fa53_or0;
  wire [0:0] csa_component58_fa54_xor1;
  wire [0:0] csa_component58_fa54_or0;
  wire [0:0] csa_component58_fa55_xor1;
  wire [0:0] csa_component58_fa55_or0;
  wire [0:0] csa_component58_fa56_xor1;
  wire [0:0] csa_component58_fa56_or0;
  wire [0:0] csa_component58_fa57_xor1;
  wire [0:0] csa_component58_fa57_or0;

  fa fa_csa_component58_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component58_fa0_xor1), .fa_or0(csa_component58_fa0_or0));
  fa fa_csa_component58_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component58_fa1_xor1), .fa_or0(csa_component58_fa1_or0));
  fa fa_csa_component58_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component58_fa2_xor1), .fa_or0(csa_component58_fa2_or0));
  fa fa_csa_component58_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component58_fa3_xor1), .fa_or0(csa_component58_fa3_or0));
  fa fa_csa_component58_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component58_fa4_xor1), .fa_or0(csa_component58_fa4_or0));
  fa fa_csa_component58_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component58_fa5_xor1), .fa_or0(csa_component58_fa5_or0));
  fa fa_csa_component58_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component58_fa6_xor1), .fa_or0(csa_component58_fa6_or0));
  fa fa_csa_component58_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component58_fa7_xor1), .fa_or0(csa_component58_fa7_or0));
  fa fa_csa_component58_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component58_fa8_xor1), .fa_or0(csa_component58_fa8_or0));
  fa fa_csa_component58_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component58_fa9_xor1), .fa_or0(csa_component58_fa9_or0));
  fa fa_csa_component58_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component58_fa10_xor1), .fa_or0(csa_component58_fa10_or0));
  fa fa_csa_component58_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component58_fa11_xor1), .fa_or0(csa_component58_fa11_or0));
  fa fa_csa_component58_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component58_fa12_xor1), .fa_or0(csa_component58_fa12_or0));
  fa fa_csa_component58_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component58_fa13_xor1), .fa_or0(csa_component58_fa13_or0));
  fa fa_csa_component58_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component58_fa14_xor1), .fa_or0(csa_component58_fa14_or0));
  fa fa_csa_component58_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component58_fa15_xor1), .fa_or0(csa_component58_fa15_or0));
  fa fa_csa_component58_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component58_fa16_xor1), .fa_or0(csa_component58_fa16_or0));
  fa fa_csa_component58_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component58_fa17_xor1), .fa_or0(csa_component58_fa17_or0));
  fa fa_csa_component58_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component58_fa18_xor1), .fa_or0(csa_component58_fa18_or0));
  fa fa_csa_component58_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component58_fa19_xor1), .fa_or0(csa_component58_fa19_or0));
  fa fa_csa_component58_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component58_fa20_xor1), .fa_or0(csa_component58_fa20_or0));
  fa fa_csa_component58_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component58_fa21_xor1), .fa_or0(csa_component58_fa21_or0));
  fa fa_csa_component58_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component58_fa22_xor1), .fa_or0(csa_component58_fa22_or0));
  fa fa_csa_component58_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component58_fa23_xor1), .fa_or0(csa_component58_fa23_or0));
  fa fa_csa_component58_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component58_fa24_xor1), .fa_or0(csa_component58_fa24_or0));
  fa fa_csa_component58_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component58_fa25_xor1), .fa_or0(csa_component58_fa25_or0));
  fa fa_csa_component58_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component58_fa26_xor1), .fa_or0(csa_component58_fa26_or0));
  fa fa_csa_component58_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component58_fa27_xor1), .fa_or0(csa_component58_fa27_or0));
  fa fa_csa_component58_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component58_fa28_xor1), .fa_or0(csa_component58_fa28_or0));
  fa fa_csa_component58_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component58_fa29_xor1), .fa_or0(csa_component58_fa29_or0));
  fa fa_csa_component58_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component58_fa30_xor1), .fa_or0(csa_component58_fa30_or0));
  fa fa_csa_component58_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component58_fa31_xor1), .fa_or0(csa_component58_fa31_or0));
  fa fa_csa_component58_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component58_fa32_xor1), .fa_or0(csa_component58_fa32_or0));
  fa fa_csa_component58_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component58_fa33_xor1), .fa_or0(csa_component58_fa33_or0));
  fa fa_csa_component58_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component58_fa34_xor1), .fa_or0(csa_component58_fa34_or0));
  fa fa_csa_component58_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component58_fa35_xor1), .fa_or0(csa_component58_fa35_or0));
  fa fa_csa_component58_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component58_fa36_xor1), .fa_or0(csa_component58_fa36_or0));
  fa fa_csa_component58_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component58_fa37_xor1), .fa_or0(csa_component58_fa37_or0));
  fa fa_csa_component58_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component58_fa38_xor1), .fa_or0(csa_component58_fa38_or0));
  fa fa_csa_component58_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component58_fa39_xor1), .fa_or0(csa_component58_fa39_or0));
  fa fa_csa_component58_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component58_fa40_xor1), .fa_or0(csa_component58_fa40_or0));
  fa fa_csa_component58_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component58_fa41_xor1), .fa_or0(csa_component58_fa41_or0));
  fa fa_csa_component58_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component58_fa42_xor1), .fa_or0(csa_component58_fa42_or0));
  fa fa_csa_component58_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component58_fa43_xor1), .fa_or0(csa_component58_fa43_or0));
  fa fa_csa_component58_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component58_fa44_xor1), .fa_or0(csa_component58_fa44_or0));
  fa fa_csa_component58_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component58_fa45_xor1), .fa_or0(csa_component58_fa45_or0));
  fa fa_csa_component58_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component58_fa46_xor1), .fa_or0(csa_component58_fa46_or0));
  fa fa_csa_component58_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component58_fa47_xor1), .fa_or0(csa_component58_fa47_or0));
  fa fa_csa_component58_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component58_fa48_xor1), .fa_or0(csa_component58_fa48_or0));
  fa fa_csa_component58_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component58_fa49_xor1), .fa_or0(csa_component58_fa49_or0));
  fa fa_csa_component58_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component58_fa50_xor1), .fa_or0(csa_component58_fa50_or0));
  fa fa_csa_component58_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component58_fa51_xor1), .fa_or0(csa_component58_fa51_or0));
  fa fa_csa_component58_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component58_fa52_xor1), .fa_or0(csa_component58_fa52_or0));
  fa fa_csa_component58_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component58_fa53_xor1), .fa_or0(csa_component58_fa53_or0));
  fa fa_csa_component58_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component58_fa54_xor1), .fa_or0(csa_component58_fa54_or0));
  fa fa_csa_component58_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component58_fa55_xor1), .fa_or0(csa_component58_fa55_or0));
  fa fa_csa_component58_fa56_out(.a(a[56]), .b(b[56]), .cin(c[56]), .fa_xor1(csa_component58_fa56_xor1), .fa_or0(csa_component58_fa56_or0));
  fa fa_csa_component58_fa57_out(.a(a[57]), .b(b[57]), .cin(c[57]), .fa_xor1(csa_component58_fa57_xor1), .fa_or0(csa_component58_fa57_or0));

  assign csa_component58_out[0] = csa_component58_fa0_xor1[0];
  assign csa_component58_out[1] = csa_component58_fa1_xor1[0];
  assign csa_component58_out[2] = csa_component58_fa2_xor1[0];
  assign csa_component58_out[3] = csa_component58_fa3_xor1[0];
  assign csa_component58_out[4] = csa_component58_fa4_xor1[0];
  assign csa_component58_out[5] = csa_component58_fa5_xor1[0];
  assign csa_component58_out[6] = csa_component58_fa6_xor1[0];
  assign csa_component58_out[7] = csa_component58_fa7_xor1[0];
  assign csa_component58_out[8] = csa_component58_fa8_xor1[0];
  assign csa_component58_out[9] = csa_component58_fa9_xor1[0];
  assign csa_component58_out[10] = csa_component58_fa10_xor1[0];
  assign csa_component58_out[11] = csa_component58_fa11_xor1[0];
  assign csa_component58_out[12] = csa_component58_fa12_xor1[0];
  assign csa_component58_out[13] = csa_component58_fa13_xor1[0];
  assign csa_component58_out[14] = csa_component58_fa14_xor1[0];
  assign csa_component58_out[15] = csa_component58_fa15_xor1[0];
  assign csa_component58_out[16] = csa_component58_fa16_xor1[0];
  assign csa_component58_out[17] = csa_component58_fa17_xor1[0];
  assign csa_component58_out[18] = csa_component58_fa18_xor1[0];
  assign csa_component58_out[19] = csa_component58_fa19_xor1[0];
  assign csa_component58_out[20] = csa_component58_fa20_xor1[0];
  assign csa_component58_out[21] = csa_component58_fa21_xor1[0];
  assign csa_component58_out[22] = csa_component58_fa22_xor1[0];
  assign csa_component58_out[23] = csa_component58_fa23_xor1[0];
  assign csa_component58_out[24] = csa_component58_fa24_xor1[0];
  assign csa_component58_out[25] = csa_component58_fa25_xor1[0];
  assign csa_component58_out[26] = csa_component58_fa26_xor1[0];
  assign csa_component58_out[27] = csa_component58_fa27_xor1[0];
  assign csa_component58_out[28] = csa_component58_fa28_xor1[0];
  assign csa_component58_out[29] = csa_component58_fa29_xor1[0];
  assign csa_component58_out[30] = csa_component58_fa30_xor1[0];
  assign csa_component58_out[31] = csa_component58_fa31_xor1[0];
  assign csa_component58_out[32] = csa_component58_fa32_xor1[0];
  assign csa_component58_out[33] = csa_component58_fa33_xor1[0];
  assign csa_component58_out[34] = csa_component58_fa34_xor1[0];
  assign csa_component58_out[35] = csa_component58_fa35_xor1[0];
  assign csa_component58_out[36] = csa_component58_fa36_xor1[0];
  assign csa_component58_out[37] = csa_component58_fa37_xor1[0];
  assign csa_component58_out[38] = csa_component58_fa38_xor1[0];
  assign csa_component58_out[39] = csa_component58_fa39_xor1[0];
  assign csa_component58_out[40] = csa_component58_fa40_xor1[0];
  assign csa_component58_out[41] = csa_component58_fa41_xor1[0];
  assign csa_component58_out[42] = csa_component58_fa42_xor1[0];
  assign csa_component58_out[43] = csa_component58_fa43_xor1[0];
  assign csa_component58_out[44] = csa_component58_fa44_xor1[0];
  assign csa_component58_out[45] = csa_component58_fa45_xor1[0];
  assign csa_component58_out[46] = csa_component58_fa46_xor1[0];
  assign csa_component58_out[47] = csa_component58_fa47_xor1[0];
  assign csa_component58_out[48] = csa_component58_fa48_xor1[0];
  assign csa_component58_out[49] = csa_component58_fa49_xor1[0];
  assign csa_component58_out[50] = csa_component58_fa50_xor1[0];
  assign csa_component58_out[51] = csa_component58_fa51_xor1[0];
  assign csa_component58_out[52] = csa_component58_fa52_xor1[0];
  assign csa_component58_out[53] = csa_component58_fa53_xor1[0];
  assign csa_component58_out[54] = csa_component58_fa54_xor1[0];
  assign csa_component58_out[55] = csa_component58_fa55_xor1[0];
  assign csa_component58_out[56] = csa_component58_fa56_xor1[0];
  assign csa_component58_out[57] = csa_component58_fa57_xor1[0];
  assign csa_component58_out[58] = 1'b0;
  assign csa_component58_out[59] = 1'b0;
  assign csa_component58_out[60] = csa_component58_fa0_or0[0];
  assign csa_component58_out[61] = csa_component58_fa1_or0[0];
  assign csa_component58_out[62] = csa_component58_fa2_or0[0];
  assign csa_component58_out[63] = csa_component58_fa3_or0[0];
  assign csa_component58_out[64] = csa_component58_fa4_or0[0];
  assign csa_component58_out[65] = csa_component58_fa5_or0[0];
  assign csa_component58_out[66] = csa_component58_fa6_or0[0];
  assign csa_component58_out[67] = csa_component58_fa7_or0[0];
  assign csa_component58_out[68] = csa_component58_fa8_or0[0];
  assign csa_component58_out[69] = csa_component58_fa9_or0[0];
  assign csa_component58_out[70] = csa_component58_fa10_or0[0];
  assign csa_component58_out[71] = csa_component58_fa11_or0[0];
  assign csa_component58_out[72] = csa_component58_fa12_or0[0];
  assign csa_component58_out[73] = csa_component58_fa13_or0[0];
  assign csa_component58_out[74] = csa_component58_fa14_or0[0];
  assign csa_component58_out[75] = csa_component58_fa15_or0[0];
  assign csa_component58_out[76] = csa_component58_fa16_or0[0];
  assign csa_component58_out[77] = csa_component58_fa17_or0[0];
  assign csa_component58_out[78] = csa_component58_fa18_or0[0];
  assign csa_component58_out[79] = csa_component58_fa19_or0[0];
  assign csa_component58_out[80] = csa_component58_fa20_or0[0];
  assign csa_component58_out[81] = csa_component58_fa21_or0[0];
  assign csa_component58_out[82] = csa_component58_fa22_or0[0];
  assign csa_component58_out[83] = csa_component58_fa23_or0[0];
  assign csa_component58_out[84] = csa_component58_fa24_or0[0];
  assign csa_component58_out[85] = csa_component58_fa25_or0[0];
  assign csa_component58_out[86] = csa_component58_fa26_or0[0];
  assign csa_component58_out[87] = csa_component58_fa27_or0[0];
  assign csa_component58_out[88] = csa_component58_fa28_or0[0];
  assign csa_component58_out[89] = csa_component58_fa29_or0[0];
  assign csa_component58_out[90] = csa_component58_fa30_or0[0];
  assign csa_component58_out[91] = csa_component58_fa31_or0[0];
  assign csa_component58_out[92] = csa_component58_fa32_or0[0];
  assign csa_component58_out[93] = csa_component58_fa33_or0[0];
  assign csa_component58_out[94] = csa_component58_fa34_or0[0];
  assign csa_component58_out[95] = csa_component58_fa35_or0[0];
  assign csa_component58_out[96] = csa_component58_fa36_or0[0];
  assign csa_component58_out[97] = csa_component58_fa37_or0[0];
  assign csa_component58_out[98] = csa_component58_fa38_or0[0];
  assign csa_component58_out[99] = csa_component58_fa39_or0[0];
  assign csa_component58_out[100] = csa_component58_fa40_or0[0];
  assign csa_component58_out[101] = csa_component58_fa41_or0[0];
  assign csa_component58_out[102] = csa_component58_fa42_or0[0];
  assign csa_component58_out[103] = csa_component58_fa43_or0[0];
  assign csa_component58_out[104] = csa_component58_fa44_or0[0];
  assign csa_component58_out[105] = csa_component58_fa45_or0[0];
  assign csa_component58_out[106] = csa_component58_fa46_or0[0];
  assign csa_component58_out[107] = csa_component58_fa47_or0[0];
  assign csa_component58_out[108] = csa_component58_fa48_or0[0];
  assign csa_component58_out[109] = csa_component58_fa49_or0[0];
  assign csa_component58_out[110] = csa_component58_fa50_or0[0];
  assign csa_component58_out[111] = csa_component58_fa51_or0[0];
  assign csa_component58_out[112] = csa_component58_fa52_or0[0];
  assign csa_component58_out[113] = csa_component58_fa53_or0[0];
  assign csa_component58_out[114] = csa_component58_fa54_or0[0];
  assign csa_component58_out[115] = csa_component58_fa55_or0[0];
  assign csa_component58_out[116] = csa_component58_fa56_or0[0];
  assign csa_component58_out[117] = csa_component58_fa57_or0[0];
endmodule

module csa_component61(input [60:0] a, input [60:0] b, input [60:0] c, output [123:0] csa_component61_out);
  wire [0:0] csa_component61_fa0_xor1;
  wire [0:0] csa_component61_fa0_or0;
  wire [0:0] csa_component61_fa1_xor1;
  wire [0:0] csa_component61_fa1_or0;
  wire [0:0] csa_component61_fa2_xor1;
  wire [0:0] csa_component61_fa2_or0;
  wire [0:0] csa_component61_fa3_xor1;
  wire [0:0] csa_component61_fa3_or0;
  wire [0:0] csa_component61_fa4_xor1;
  wire [0:0] csa_component61_fa4_or0;
  wire [0:0] csa_component61_fa5_xor1;
  wire [0:0] csa_component61_fa5_or0;
  wire [0:0] csa_component61_fa6_xor1;
  wire [0:0] csa_component61_fa6_or0;
  wire [0:0] csa_component61_fa7_xor1;
  wire [0:0] csa_component61_fa7_or0;
  wire [0:0] csa_component61_fa8_xor1;
  wire [0:0] csa_component61_fa8_or0;
  wire [0:0] csa_component61_fa9_xor1;
  wire [0:0] csa_component61_fa9_or0;
  wire [0:0] csa_component61_fa10_xor1;
  wire [0:0] csa_component61_fa10_or0;
  wire [0:0] csa_component61_fa11_xor1;
  wire [0:0] csa_component61_fa11_or0;
  wire [0:0] csa_component61_fa12_xor1;
  wire [0:0] csa_component61_fa12_or0;
  wire [0:0] csa_component61_fa13_xor1;
  wire [0:0] csa_component61_fa13_or0;
  wire [0:0] csa_component61_fa14_xor1;
  wire [0:0] csa_component61_fa14_or0;
  wire [0:0] csa_component61_fa15_xor1;
  wire [0:0] csa_component61_fa15_or0;
  wire [0:0] csa_component61_fa16_xor1;
  wire [0:0] csa_component61_fa16_or0;
  wire [0:0] csa_component61_fa17_xor1;
  wire [0:0] csa_component61_fa17_or0;
  wire [0:0] csa_component61_fa18_xor1;
  wire [0:0] csa_component61_fa18_or0;
  wire [0:0] csa_component61_fa19_xor1;
  wire [0:0] csa_component61_fa19_or0;
  wire [0:0] csa_component61_fa20_xor1;
  wire [0:0] csa_component61_fa20_or0;
  wire [0:0] csa_component61_fa21_xor1;
  wire [0:0] csa_component61_fa21_or0;
  wire [0:0] csa_component61_fa22_xor1;
  wire [0:0] csa_component61_fa22_or0;
  wire [0:0] csa_component61_fa23_xor1;
  wire [0:0] csa_component61_fa23_or0;
  wire [0:0] csa_component61_fa24_xor1;
  wire [0:0] csa_component61_fa24_or0;
  wire [0:0] csa_component61_fa25_xor1;
  wire [0:0] csa_component61_fa25_or0;
  wire [0:0] csa_component61_fa26_xor1;
  wire [0:0] csa_component61_fa26_or0;
  wire [0:0] csa_component61_fa27_xor1;
  wire [0:0] csa_component61_fa27_or0;
  wire [0:0] csa_component61_fa28_xor1;
  wire [0:0] csa_component61_fa28_or0;
  wire [0:0] csa_component61_fa29_xor1;
  wire [0:0] csa_component61_fa29_or0;
  wire [0:0] csa_component61_fa30_xor1;
  wire [0:0] csa_component61_fa30_or0;
  wire [0:0] csa_component61_fa31_xor1;
  wire [0:0] csa_component61_fa31_or0;
  wire [0:0] csa_component61_fa32_xor1;
  wire [0:0] csa_component61_fa32_or0;
  wire [0:0] csa_component61_fa33_xor1;
  wire [0:0] csa_component61_fa33_or0;
  wire [0:0] csa_component61_fa34_xor1;
  wire [0:0] csa_component61_fa34_or0;
  wire [0:0] csa_component61_fa35_xor1;
  wire [0:0] csa_component61_fa35_or0;
  wire [0:0] csa_component61_fa36_xor1;
  wire [0:0] csa_component61_fa36_or0;
  wire [0:0] csa_component61_fa37_xor1;
  wire [0:0] csa_component61_fa37_or0;
  wire [0:0] csa_component61_fa38_xor1;
  wire [0:0] csa_component61_fa38_or0;
  wire [0:0] csa_component61_fa39_xor1;
  wire [0:0] csa_component61_fa39_or0;
  wire [0:0] csa_component61_fa40_xor1;
  wire [0:0] csa_component61_fa40_or0;
  wire [0:0] csa_component61_fa41_xor1;
  wire [0:0] csa_component61_fa41_or0;
  wire [0:0] csa_component61_fa42_xor1;
  wire [0:0] csa_component61_fa42_or0;
  wire [0:0] csa_component61_fa43_xor1;
  wire [0:0] csa_component61_fa43_or0;
  wire [0:0] csa_component61_fa44_xor1;
  wire [0:0] csa_component61_fa44_or0;
  wire [0:0] csa_component61_fa45_xor1;
  wire [0:0] csa_component61_fa45_or0;
  wire [0:0] csa_component61_fa46_xor1;
  wire [0:0] csa_component61_fa46_or0;
  wire [0:0] csa_component61_fa47_xor1;
  wire [0:0] csa_component61_fa47_or0;
  wire [0:0] csa_component61_fa48_xor1;
  wire [0:0] csa_component61_fa48_or0;
  wire [0:0] csa_component61_fa49_xor1;
  wire [0:0] csa_component61_fa49_or0;
  wire [0:0] csa_component61_fa50_xor1;
  wire [0:0] csa_component61_fa50_or0;
  wire [0:0] csa_component61_fa51_xor1;
  wire [0:0] csa_component61_fa51_or0;
  wire [0:0] csa_component61_fa52_xor1;
  wire [0:0] csa_component61_fa52_or0;
  wire [0:0] csa_component61_fa53_xor1;
  wire [0:0] csa_component61_fa53_or0;
  wire [0:0] csa_component61_fa54_xor1;
  wire [0:0] csa_component61_fa54_or0;
  wire [0:0] csa_component61_fa55_xor1;
  wire [0:0] csa_component61_fa55_or0;
  wire [0:0] csa_component61_fa56_xor1;
  wire [0:0] csa_component61_fa56_or0;
  wire [0:0] csa_component61_fa57_xor1;
  wire [0:0] csa_component61_fa57_or0;
  wire [0:0] csa_component61_fa58_xor1;
  wire [0:0] csa_component61_fa58_or0;
  wire [0:0] csa_component61_fa59_xor1;
  wire [0:0] csa_component61_fa59_or0;
  wire [0:0] csa_component61_fa60_xor1;
  wire [0:0] csa_component61_fa60_or0;

  fa fa_csa_component61_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component61_fa0_xor1), .fa_or0(csa_component61_fa0_or0));
  fa fa_csa_component61_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component61_fa1_xor1), .fa_or0(csa_component61_fa1_or0));
  fa fa_csa_component61_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component61_fa2_xor1), .fa_or0(csa_component61_fa2_or0));
  fa fa_csa_component61_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component61_fa3_xor1), .fa_or0(csa_component61_fa3_or0));
  fa fa_csa_component61_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component61_fa4_xor1), .fa_or0(csa_component61_fa4_or0));
  fa fa_csa_component61_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component61_fa5_xor1), .fa_or0(csa_component61_fa5_or0));
  fa fa_csa_component61_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component61_fa6_xor1), .fa_or0(csa_component61_fa6_or0));
  fa fa_csa_component61_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component61_fa7_xor1), .fa_or0(csa_component61_fa7_or0));
  fa fa_csa_component61_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component61_fa8_xor1), .fa_or0(csa_component61_fa8_or0));
  fa fa_csa_component61_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component61_fa9_xor1), .fa_or0(csa_component61_fa9_or0));
  fa fa_csa_component61_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component61_fa10_xor1), .fa_or0(csa_component61_fa10_or0));
  fa fa_csa_component61_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component61_fa11_xor1), .fa_or0(csa_component61_fa11_or0));
  fa fa_csa_component61_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component61_fa12_xor1), .fa_or0(csa_component61_fa12_or0));
  fa fa_csa_component61_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component61_fa13_xor1), .fa_or0(csa_component61_fa13_or0));
  fa fa_csa_component61_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component61_fa14_xor1), .fa_or0(csa_component61_fa14_or0));
  fa fa_csa_component61_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component61_fa15_xor1), .fa_or0(csa_component61_fa15_or0));
  fa fa_csa_component61_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component61_fa16_xor1), .fa_or0(csa_component61_fa16_or0));
  fa fa_csa_component61_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component61_fa17_xor1), .fa_or0(csa_component61_fa17_or0));
  fa fa_csa_component61_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component61_fa18_xor1), .fa_or0(csa_component61_fa18_or0));
  fa fa_csa_component61_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component61_fa19_xor1), .fa_or0(csa_component61_fa19_or0));
  fa fa_csa_component61_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component61_fa20_xor1), .fa_or0(csa_component61_fa20_or0));
  fa fa_csa_component61_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component61_fa21_xor1), .fa_or0(csa_component61_fa21_or0));
  fa fa_csa_component61_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component61_fa22_xor1), .fa_or0(csa_component61_fa22_or0));
  fa fa_csa_component61_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component61_fa23_xor1), .fa_or0(csa_component61_fa23_or0));
  fa fa_csa_component61_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component61_fa24_xor1), .fa_or0(csa_component61_fa24_or0));
  fa fa_csa_component61_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component61_fa25_xor1), .fa_or0(csa_component61_fa25_or0));
  fa fa_csa_component61_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component61_fa26_xor1), .fa_or0(csa_component61_fa26_or0));
  fa fa_csa_component61_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component61_fa27_xor1), .fa_or0(csa_component61_fa27_or0));
  fa fa_csa_component61_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component61_fa28_xor1), .fa_or0(csa_component61_fa28_or0));
  fa fa_csa_component61_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component61_fa29_xor1), .fa_or0(csa_component61_fa29_or0));
  fa fa_csa_component61_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component61_fa30_xor1), .fa_or0(csa_component61_fa30_or0));
  fa fa_csa_component61_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component61_fa31_xor1), .fa_or0(csa_component61_fa31_or0));
  fa fa_csa_component61_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component61_fa32_xor1), .fa_or0(csa_component61_fa32_or0));
  fa fa_csa_component61_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component61_fa33_xor1), .fa_or0(csa_component61_fa33_or0));
  fa fa_csa_component61_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component61_fa34_xor1), .fa_or0(csa_component61_fa34_or0));
  fa fa_csa_component61_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component61_fa35_xor1), .fa_or0(csa_component61_fa35_or0));
  fa fa_csa_component61_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component61_fa36_xor1), .fa_or0(csa_component61_fa36_or0));
  fa fa_csa_component61_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component61_fa37_xor1), .fa_or0(csa_component61_fa37_or0));
  fa fa_csa_component61_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component61_fa38_xor1), .fa_or0(csa_component61_fa38_or0));
  fa fa_csa_component61_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component61_fa39_xor1), .fa_or0(csa_component61_fa39_or0));
  fa fa_csa_component61_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component61_fa40_xor1), .fa_or0(csa_component61_fa40_or0));
  fa fa_csa_component61_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component61_fa41_xor1), .fa_or0(csa_component61_fa41_or0));
  fa fa_csa_component61_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component61_fa42_xor1), .fa_or0(csa_component61_fa42_or0));
  fa fa_csa_component61_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component61_fa43_xor1), .fa_or0(csa_component61_fa43_or0));
  fa fa_csa_component61_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component61_fa44_xor1), .fa_or0(csa_component61_fa44_or0));
  fa fa_csa_component61_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component61_fa45_xor1), .fa_or0(csa_component61_fa45_or0));
  fa fa_csa_component61_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component61_fa46_xor1), .fa_or0(csa_component61_fa46_or0));
  fa fa_csa_component61_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component61_fa47_xor1), .fa_or0(csa_component61_fa47_or0));
  fa fa_csa_component61_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component61_fa48_xor1), .fa_or0(csa_component61_fa48_or0));
  fa fa_csa_component61_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component61_fa49_xor1), .fa_or0(csa_component61_fa49_or0));
  fa fa_csa_component61_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component61_fa50_xor1), .fa_or0(csa_component61_fa50_or0));
  fa fa_csa_component61_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component61_fa51_xor1), .fa_or0(csa_component61_fa51_or0));
  fa fa_csa_component61_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component61_fa52_xor1), .fa_or0(csa_component61_fa52_or0));
  fa fa_csa_component61_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component61_fa53_xor1), .fa_or0(csa_component61_fa53_or0));
  fa fa_csa_component61_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component61_fa54_xor1), .fa_or0(csa_component61_fa54_or0));
  fa fa_csa_component61_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component61_fa55_xor1), .fa_or0(csa_component61_fa55_or0));
  fa fa_csa_component61_fa56_out(.a(a[56]), .b(b[56]), .cin(c[56]), .fa_xor1(csa_component61_fa56_xor1), .fa_or0(csa_component61_fa56_or0));
  fa fa_csa_component61_fa57_out(.a(a[57]), .b(b[57]), .cin(c[57]), .fa_xor1(csa_component61_fa57_xor1), .fa_or0(csa_component61_fa57_or0));
  fa fa_csa_component61_fa58_out(.a(a[58]), .b(b[58]), .cin(c[58]), .fa_xor1(csa_component61_fa58_xor1), .fa_or0(csa_component61_fa58_or0));
  fa fa_csa_component61_fa59_out(.a(a[59]), .b(b[59]), .cin(c[59]), .fa_xor1(csa_component61_fa59_xor1), .fa_or0(csa_component61_fa59_or0));
  fa fa_csa_component61_fa60_out(.a(a[60]), .b(b[60]), .cin(c[60]), .fa_xor1(csa_component61_fa60_xor1), .fa_or0(csa_component61_fa60_or0));

  assign csa_component61_out[0] = csa_component61_fa0_xor1[0];
  assign csa_component61_out[1] = csa_component61_fa1_xor1[0];
  assign csa_component61_out[2] = csa_component61_fa2_xor1[0];
  assign csa_component61_out[3] = csa_component61_fa3_xor1[0];
  assign csa_component61_out[4] = csa_component61_fa4_xor1[0];
  assign csa_component61_out[5] = csa_component61_fa5_xor1[0];
  assign csa_component61_out[6] = csa_component61_fa6_xor1[0];
  assign csa_component61_out[7] = csa_component61_fa7_xor1[0];
  assign csa_component61_out[8] = csa_component61_fa8_xor1[0];
  assign csa_component61_out[9] = csa_component61_fa9_xor1[0];
  assign csa_component61_out[10] = csa_component61_fa10_xor1[0];
  assign csa_component61_out[11] = csa_component61_fa11_xor1[0];
  assign csa_component61_out[12] = csa_component61_fa12_xor1[0];
  assign csa_component61_out[13] = csa_component61_fa13_xor1[0];
  assign csa_component61_out[14] = csa_component61_fa14_xor1[0];
  assign csa_component61_out[15] = csa_component61_fa15_xor1[0];
  assign csa_component61_out[16] = csa_component61_fa16_xor1[0];
  assign csa_component61_out[17] = csa_component61_fa17_xor1[0];
  assign csa_component61_out[18] = csa_component61_fa18_xor1[0];
  assign csa_component61_out[19] = csa_component61_fa19_xor1[0];
  assign csa_component61_out[20] = csa_component61_fa20_xor1[0];
  assign csa_component61_out[21] = csa_component61_fa21_xor1[0];
  assign csa_component61_out[22] = csa_component61_fa22_xor1[0];
  assign csa_component61_out[23] = csa_component61_fa23_xor1[0];
  assign csa_component61_out[24] = csa_component61_fa24_xor1[0];
  assign csa_component61_out[25] = csa_component61_fa25_xor1[0];
  assign csa_component61_out[26] = csa_component61_fa26_xor1[0];
  assign csa_component61_out[27] = csa_component61_fa27_xor1[0];
  assign csa_component61_out[28] = csa_component61_fa28_xor1[0];
  assign csa_component61_out[29] = csa_component61_fa29_xor1[0];
  assign csa_component61_out[30] = csa_component61_fa30_xor1[0];
  assign csa_component61_out[31] = csa_component61_fa31_xor1[0];
  assign csa_component61_out[32] = csa_component61_fa32_xor1[0];
  assign csa_component61_out[33] = csa_component61_fa33_xor1[0];
  assign csa_component61_out[34] = csa_component61_fa34_xor1[0];
  assign csa_component61_out[35] = csa_component61_fa35_xor1[0];
  assign csa_component61_out[36] = csa_component61_fa36_xor1[0];
  assign csa_component61_out[37] = csa_component61_fa37_xor1[0];
  assign csa_component61_out[38] = csa_component61_fa38_xor1[0];
  assign csa_component61_out[39] = csa_component61_fa39_xor1[0];
  assign csa_component61_out[40] = csa_component61_fa40_xor1[0];
  assign csa_component61_out[41] = csa_component61_fa41_xor1[0];
  assign csa_component61_out[42] = csa_component61_fa42_xor1[0];
  assign csa_component61_out[43] = csa_component61_fa43_xor1[0];
  assign csa_component61_out[44] = csa_component61_fa44_xor1[0];
  assign csa_component61_out[45] = csa_component61_fa45_xor1[0];
  assign csa_component61_out[46] = csa_component61_fa46_xor1[0];
  assign csa_component61_out[47] = csa_component61_fa47_xor1[0];
  assign csa_component61_out[48] = csa_component61_fa48_xor1[0];
  assign csa_component61_out[49] = csa_component61_fa49_xor1[0];
  assign csa_component61_out[50] = csa_component61_fa50_xor1[0];
  assign csa_component61_out[51] = csa_component61_fa51_xor1[0];
  assign csa_component61_out[52] = csa_component61_fa52_xor1[0];
  assign csa_component61_out[53] = csa_component61_fa53_xor1[0];
  assign csa_component61_out[54] = csa_component61_fa54_xor1[0];
  assign csa_component61_out[55] = csa_component61_fa55_xor1[0];
  assign csa_component61_out[56] = csa_component61_fa56_xor1[0];
  assign csa_component61_out[57] = csa_component61_fa57_xor1[0];
  assign csa_component61_out[58] = csa_component61_fa58_xor1[0];
  assign csa_component61_out[59] = csa_component61_fa59_xor1[0];
  assign csa_component61_out[60] = csa_component61_fa60_xor1[0];
  assign csa_component61_out[61] = 1'b0;
  assign csa_component61_out[62] = 1'b0;
  assign csa_component61_out[63] = csa_component61_fa0_or0[0];
  assign csa_component61_out[64] = csa_component61_fa1_or0[0];
  assign csa_component61_out[65] = csa_component61_fa2_or0[0];
  assign csa_component61_out[66] = csa_component61_fa3_or0[0];
  assign csa_component61_out[67] = csa_component61_fa4_or0[0];
  assign csa_component61_out[68] = csa_component61_fa5_or0[0];
  assign csa_component61_out[69] = csa_component61_fa6_or0[0];
  assign csa_component61_out[70] = csa_component61_fa7_or0[0];
  assign csa_component61_out[71] = csa_component61_fa8_or0[0];
  assign csa_component61_out[72] = csa_component61_fa9_or0[0];
  assign csa_component61_out[73] = csa_component61_fa10_or0[0];
  assign csa_component61_out[74] = csa_component61_fa11_or0[0];
  assign csa_component61_out[75] = csa_component61_fa12_or0[0];
  assign csa_component61_out[76] = csa_component61_fa13_or0[0];
  assign csa_component61_out[77] = csa_component61_fa14_or0[0];
  assign csa_component61_out[78] = csa_component61_fa15_or0[0];
  assign csa_component61_out[79] = csa_component61_fa16_or0[0];
  assign csa_component61_out[80] = csa_component61_fa17_or0[0];
  assign csa_component61_out[81] = csa_component61_fa18_or0[0];
  assign csa_component61_out[82] = csa_component61_fa19_or0[0];
  assign csa_component61_out[83] = csa_component61_fa20_or0[0];
  assign csa_component61_out[84] = csa_component61_fa21_or0[0];
  assign csa_component61_out[85] = csa_component61_fa22_or0[0];
  assign csa_component61_out[86] = csa_component61_fa23_or0[0];
  assign csa_component61_out[87] = csa_component61_fa24_or0[0];
  assign csa_component61_out[88] = csa_component61_fa25_or0[0];
  assign csa_component61_out[89] = csa_component61_fa26_or0[0];
  assign csa_component61_out[90] = csa_component61_fa27_or0[0];
  assign csa_component61_out[91] = csa_component61_fa28_or0[0];
  assign csa_component61_out[92] = csa_component61_fa29_or0[0];
  assign csa_component61_out[93] = csa_component61_fa30_or0[0];
  assign csa_component61_out[94] = csa_component61_fa31_or0[0];
  assign csa_component61_out[95] = csa_component61_fa32_or0[0];
  assign csa_component61_out[96] = csa_component61_fa33_or0[0];
  assign csa_component61_out[97] = csa_component61_fa34_or0[0];
  assign csa_component61_out[98] = csa_component61_fa35_or0[0];
  assign csa_component61_out[99] = csa_component61_fa36_or0[0];
  assign csa_component61_out[100] = csa_component61_fa37_or0[0];
  assign csa_component61_out[101] = csa_component61_fa38_or0[0];
  assign csa_component61_out[102] = csa_component61_fa39_or0[0];
  assign csa_component61_out[103] = csa_component61_fa40_or0[0];
  assign csa_component61_out[104] = csa_component61_fa41_or0[0];
  assign csa_component61_out[105] = csa_component61_fa42_or0[0];
  assign csa_component61_out[106] = csa_component61_fa43_or0[0];
  assign csa_component61_out[107] = csa_component61_fa44_or0[0];
  assign csa_component61_out[108] = csa_component61_fa45_or0[0];
  assign csa_component61_out[109] = csa_component61_fa46_or0[0];
  assign csa_component61_out[110] = csa_component61_fa47_or0[0];
  assign csa_component61_out[111] = csa_component61_fa48_or0[0];
  assign csa_component61_out[112] = csa_component61_fa49_or0[0];
  assign csa_component61_out[113] = csa_component61_fa50_or0[0];
  assign csa_component61_out[114] = csa_component61_fa51_or0[0];
  assign csa_component61_out[115] = csa_component61_fa52_or0[0];
  assign csa_component61_out[116] = csa_component61_fa53_or0[0];
  assign csa_component61_out[117] = csa_component61_fa54_or0[0];
  assign csa_component61_out[118] = csa_component61_fa55_or0[0];
  assign csa_component61_out[119] = csa_component61_fa56_or0[0];
  assign csa_component61_out[120] = csa_component61_fa57_or0[0];
  assign csa_component61_out[121] = csa_component61_fa58_or0[0];
  assign csa_component61_out[122] = csa_component61_fa59_or0[0];
  assign csa_component61_out[123] = csa_component61_fa60_or0[0];
endmodule

module csa_component38(input [37:0] a, input [37:0] b, input [37:0] c, output [77:0] csa_component38_out);
  wire [0:0] csa_component38_fa0_xor1;
  wire [0:0] csa_component38_fa0_or0;
  wire [0:0] csa_component38_fa1_xor1;
  wire [0:0] csa_component38_fa1_or0;
  wire [0:0] csa_component38_fa2_xor1;
  wire [0:0] csa_component38_fa2_or0;
  wire [0:0] csa_component38_fa3_xor1;
  wire [0:0] csa_component38_fa3_or0;
  wire [0:0] csa_component38_fa4_xor1;
  wire [0:0] csa_component38_fa4_or0;
  wire [0:0] csa_component38_fa5_xor1;
  wire [0:0] csa_component38_fa5_or0;
  wire [0:0] csa_component38_fa6_xor1;
  wire [0:0] csa_component38_fa6_or0;
  wire [0:0] csa_component38_fa7_xor1;
  wire [0:0] csa_component38_fa7_or0;
  wire [0:0] csa_component38_fa8_xor1;
  wire [0:0] csa_component38_fa8_or0;
  wire [0:0] csa_component38_fa9_xor1;
  wire [0:0] csa_component38_fa9_or0;
  wire [0:0] csa_component38_fa10_xor1;
  wire [0:0] csa_component38_fa10_or0;
  wire [0:0] csa_component38_fa11_xor1;
  wire [0:0] csa_component38_fa11_or0;
  wire [0:0] csa_component38_fa12_xor1;
  wire [0:0] csa_component38_fa12_or0;
  wire [0:0] csa_component38_fa13_xor1;
  wire [0:0] csa_component38_fa13_or0;
  wire [0:0] csa_component38_fa14_xor1;
  wire [0:0] csa_component38_fa14_or0;
  wire [0:0] csa_component38_fa15_xor1;
  wire [0:0] csa_component38_fa15_or0;
  wire [0:0] csa_component38_fa16_xor1;
  wire [0:0] csa_component38_fa16_or0;
  wire [0:0] csa_component38_fa17_xor1;
  wire [0:0] csa_component38_fa17_or0;
  wire [0:0] csa_component38_fa18_xor1;
  wire [0:0] csa_component38_fa18_or0;
  wire [0:0] csa_component38_fa19_xor1;
  wire [0:0] csa_component38_fa19_or0;
  wire [0:0] csa_component38_fa20_xor1;
  wire [0:0] csa_component38_fa20_or0;
  wire [0:0] csa_component38_fa21_xor1;
  wire [0:0] csa_component38_fa21_or0;
  wire [0:0] csa_component38_fa22_xor1;
  wire [0:0] csa_component38_fa22_or0;
  wire [0:0] csa_component38_fa23_xor1;
  wire [0:0] csa_component38_fa23_or0;
  wire [0:0] csa_component38_fa24_xor1;
  wire [0:0] csa_component38_fa24_or0;
  wire [0:0] csa_component38_fa25_xor1;
  wire [0:0] csa_component38_fa25_or0;
  wire [0:0] csa_component38_fa26_xor1;
  wire [0:0] csa_component38_fa26_or0;
  wire [0:0] csa_component38_fa27_xor1;
  wire [0:0] csa_component38_fa27_or0;
  wire [0:0] csa_component38_fa28_xor1;
  wire [0:0] csa_component38_fa28_or0;
  wire [0:0] csa_component38_fa29_xor1;
  wire [0:0] csa_component38_fa29_or0;
  wire [0:0] csa_component38_fa30_xor1;
  wire [0:0] csa_component38_fa30_or0;
  wire [0:0] csa_component38_fa31_xor1;
  wire [0:0] csa_component38_fa31_or0;
  wire [0:0] csa_component38_fa32_xor1;
  wire [0:0] csa_component38_fa32_or0;
  wire [0:0] csa_component38_fa33_xor1;
  wire [0:0] csa_component38_fa33_or0;
  wire [0:0] csa_component38_fa34_xor1;
  wire [0:0] csa_component38_fa34_or0;
  wire [0:0] csa_component38_fa35_xor1;
  wire [0:0] csa_component38_fa35_or0;
  wire [0:0] csa_component38_fa36_xor1;
  wire [0:0] csa_component38_fa36_or0;
  wire [0:0] csa_component38_fa37_xor1;
  wire [0:0] csa_component38_fa37_or0;

  fa fa_csa_component38_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component38_fa0_xor1), .fa_or0(csa_component38_fa0_or0));
  fa fa_csa_component38_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component38_fa1_xor1), .fa_or0(csa_component38_fa1_or0));
  fa fa_csa_component38_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component38_fa2_xor1), .fa_or0(csa_component38_fa2_or0));
  fa fa_csa_component38_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component38_fa3_xor1), .fa_or0(csa_component38_fa3_or0));
  fa fa_csa_component38_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component38_fa4_xor1), .fa_or0(csa_component38_fa4_or0));
  fa fa_csa_component38_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component38_fa5_xor1), .fa_or0(csa_component38_fa5_or0));
  fa fa_csa_component38_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component38_fa6_xor1), .fa_or0(csa_component38_fa6_or0));
  fa fa_csa_component38_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component38_fa7_xor1), .fa_or0(csa_component38_fa7_or0));
  fa fa_csa_component38_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component38_fa8_xor1), .fa_or0(csa_component38_fa8_or0));
  fa fa_csa_component38_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component38_fa9_xor1), .fa_or0(csa_component38_fa9_or0));
  fa fa_csa_component38_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component38_fa10_xor1), .fa_or0(csa_component38_fa10_or0));
  fa fa_csa_component38_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component38_fa11_xor1), .fa_or0(csa_component38_fa11_or0));
  fa fa_csa_component38_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component38_fa12_xor1), .fa_or0(csa_component38_fa12_or0));
  fa fa_csa_component38_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component38_fa13_xor1), .fa_or0(csa_component38_fa13_or0));
  fa fa_csa_component38_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component38_fa14_xor1), .fa_or0(csa_component38_fa14_or0));
  fa fa_csa_component38_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component38_fa15_xor1), .fa_or0(csa_component38_fa15_or0));
  fa fa_csa_component38_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component38_fa16_xor1), .fa_or0(csa_component38_fa16_or0));
  fa fa_csa_component38_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component38_fa17_xor1), .fa_or0(csa_component38_fa17_or0));
  fa fa_csa_component38_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component38_fa18_xor1), .fa_or0(csa_component38_fa18_or0));
  fa fa_csa_component38_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component38_fa19_xor1), .fa_or0(csa_component38_fa19_or0));
  fa fa_csa_component38_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component38_fa20_xor1), .fa_or0(csa_component38_fa20_or0));
  fa fa_csa_component38_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component38_fa21_xor1), .fa_or0(csa_component38_fa21_or0));
  fa fa_csa_component38_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component38_fa22_xor1), .fa_or0(csa_component38_fa22_or0));
  fa fa_csa_component38_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component38_fa23_xor1), .fa_or0(csa_component38_fa23_or0));
  fa fa_csa_component38_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component38_fa24_xor1), .fa_or0(csa_component38_fa24_or0));
  fa fa_csa_component38_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component38_fa25_xor1), .fa_or0(csa_component38_fa25_or0));
  fa fa_csa_component38_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component38_fa26_xor1), .fa_or0(csa_component38_fa26_or0));
  fa fa_csa_component38_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component38_fa27_xor1), .fa_or0(csa_component38_fa27_or0));
  fa fa_csa_component38_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component38_fa28_xor1), .fa_or0(csa_component38_fa28_or0));
  fa fa_csa_component38_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component38_fa29_xor1), .fa_or0(csa_component38_fa29_or0));
  fa fa_csa_component38_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component38_fa30_xor1), .fa_or0(csa_component38_fa30_or0));
  fa fa_csa_component38_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component38_fa31_xor1), .fa_or0(csa_component38_fa31_or0));
  fa fa_csa_component38_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component38_fa32_xor1), .fa_or0(csa_component38_fa32_or0));
  fa fa_csa_component38_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component38_fa33_xor1), .fa_or0(csa_component38_fa33_or0));
  fa fa_csa_component38_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component38_fa34_xor1), .fa_or0(csa_component38_fa34_or0));
  fa fa_csa_component38_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component38_fa35_xor1), .fa_or0(csa_component38_fa35_or0));
  fa fa_csa_component38_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component38_fa36_xor1), .fa_or0(csa_component38_fa36_or0));
  fa fa_csa_component38_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component38_fa37_xor1), .fa_or0(csa_component38_fa37_or0));

  assign csa_component38_out[0] = csa_component38_fa0_xor1[0];
  assign csa_component38_out[1] = csa_component38_fa1_xor1[0];
  assign csa_component38_out[2] = csa_component38_fa2_xor1[0];
  assign csa_component38_out[3] = csa_component38_fa3_xor1[0];
  assign csa_component38_out[4] = csa_component38_fa4_xor1[0];
  assign csa_component38_out[5] = csa_component38_fa5_xor1[0];
  assign csa_component38_out[6] = csa_component38_fa6_xor1[0];
  assign csa_component38_out[7] = csa_component38_fa7_xor1[0];
  assign csa_component38_out[8] = csa_component38_fa8_xor1[0];
  assign csa_component38_out[9] = csa_component38_fa9_xor1[0];
  assign csa_component38_out[10] = csa_component38_fa10_xor1[0];
  assign csa_component38_out[11] = csa_component38_fa11_xor1[0];
  assign csa_component38_out[12] = csa_component38_fa12_xor1[0];
  assign csa_component38_out[13] = csa_component38_fa13_xor1[0];
  assign csa_component38_out[14] = csa_component38_fa14_xor1[0];
  assign csa_component38_out[15] = csa_component38_fa15_xor1[0];
  assign csa_component38_out[16] = csa_component38_fa16_xor1[0];
  assign csa_component38_out[17] = csa_component38_fa17_xor1[0];
  assign csa_component38_out[18] = csa_component38_fa18_xor1[0];
  assign csa_component38_out[19] = csa_component38_fa19_xor1[0];
  assign csa_component38_out[20] = csa_component38_fa20_xor1[0];
  assign csa_component38_out[21] = csa_component38_fa21_xor1[0];
  assign csa_component38_out[22] = csa_component38_fa22_xor1[0];
  assign csa_component38_out[23] = csa_component38_fa23_xor1[0];
  assign csa_component38_out[24] = csa_component38_fa24_xor1[0];
  assign csa_component38_out[25] = csa_component38_fa25_xor1[0];
  assign csa_component38_out[26] = csa_component38_fa26_xor1[0];
  assign csa_component38_out[27] = csa_component38_fa27_xor1[0];
  assign csa_component38_out[28] = csa_component38_fa28_xor1[0];
  assign csa_component38_out[29] = csa_component38_fa29_xor1[0];
  assign csa_component38_out[30] = csa_component38_fa30_xor1[0];
  assign csa_component38_out[31] = csa_component38_fa31_xor1[0];
  assign csa_component38_out[32] = csa_component38_fa32_xor1[0];
  assign csa_component38_out[33] = csa_component38_fa33_xor1[0];
  assign csa_component38_out[34] = csa_component38_fa34_xor1[0];
  assign csa_component38_out[35] = csa_component38_fa35_xor1[0];
  assign csa_component38_out[36] = csa_component38_fa36_xor1[0];
  assign csa_component38_out[37] = csa_component38_fa37_xor1[0];
  assign csa_component38_out[38] = 1'b0;
  assign csa_component38_out[39] = 1'b0;
  assign csa_component38_out[40] = csa_component38_fa0_or0[0];
  assign csa_component38_out[41] = csa_component38_fa1_or0[0];
  assign csa_component38_out[42] = csa_component38_fa2_or0[0];
  assign csa_component38_out[43] = csa_component38_fa3_or0[0];
  assign csa_component38_out[44] = csa_component38_fa4_or0[0];
  assign csa_component38_out[45] = csa_component38_fa5_or0[0];
  assign csa_component38_out[46] = csa_component38_fa6_or0[0];
  assign csa_component38_out[47] = csa_component38_fa7_or0[0];
  assign csa_component38_out[48] = csa_component38_fa8_or0[0];
  assign csa_component38_out[49] = csa_component38_fa9_or0[0];
  assign csa_component38_out[50] = csa_component38_fa10_or0[0];
  assign csa_component38_out[51] = csa_component38_fa11_or0[0];
  assign csa_component38_out[52] = csa_component38_fa12_or0[0];
  assign csa_component38_out[53] = csa_component38_fa13_or0[0];
  assign csa_component38_out[54] = csa_component38_fa14_or0[0];
  assign csa_component38_out[55] = csa_component38_fa15_or0[0];
  assign csa_component38_out[56] = csa_component38_fa16_or0[0];
  assign csa_component38_out[57] = csa_component38_fa17_or0[0];
  assign csa_component38_out[58] = csa_component38_fa18_or0[0];
  assign csa_component38_out[59] = csa_component38_fa19_or0[0];
  assign csa_component38_out[60] = csa_component38_fa20_or0[0];
  assign csa_component38_out[61] = csa_component38_fa21_or0[0];
  assign csa_component38_out[62] = csa_component38_fa22_or0[0];
  assign csa_component38_out[63] = csa_component38_fa23_or0[0];
  assign csa_component38_out[64] = csa_component38_fa24_or0[0];
  assign csa_component38_out[65] = csa_component38_fa25_or0[0];
  assign csa_component38_out[66] = csa_component38_fa26_or0[0];
  assign csa_component38_out[67] = csa_component38_fa27_or0[0];
  assign csa_component38_out[68] = csa_component38_fa28_or0[0];
  assign csa_component38_out[69] = csa_component38_fa29_or0[0];
  assign csa_component38_out[70] = csa_component38_fa30_or0[0];
  assign csa_component38_out[71] = csa_component38_fa31_or0[0];
  assign csa_component38_out[72] = csa_component38_fa32_or0[0];
  assign csa_component38_out[73] = csa_component38_fa33_or0[0];
  assign csa_component38_out[74] = csa_component38_fa34_or0[0];
  assign csa_component38_out[75] = csa_component38_fa35_or0[0];
  assign csa_component38_out[76] = csa_component38_fa36_or0[0];
  assign csa_component38_out[77] = csa_component38_fa37_or0[0];
endmodule

module csa_component41(input [40:0] a, input [40:0] b, input [40:0] c, output [83:0] csa_component41_out);
  wire [0:0] csa_component41_fa0_xor1;
  wire [0:0] csa_component41_fa0_or0;
  wire [0:0] csa_component41_fa1_xor1;
  wire [0:0] csa_component41_fa1_or0;
  wire [0:0] csa_component41_fa2_xor1;
  wire [0:0] csa_component41_fa2_or0;
  wire [0:0] csa_component41_fa3_xor1;
  wire [0:0] csa_component41_fa3_or0;
  wire [0:0] csa_component41_fa4_xor1;
  wire [0:0] csa_component41_fa4_or0;
  wire [0:0] csa_component41_fa5_xor1;
  wire [0:0] csa_component41_fa5_or0;
  wire [0:0] csa_component41_fa6_xor1;
  wire [0:0] csa_component41_fa6_or0;
  wire [0:0] csa_component41_fa7_xor1;
  wire [0:0] csa_component41_fa7_or0;
  wire [0:0] csa_component41_fa8_xor1;
  wire [0:0] csa_component41_fa8_or0;
  wire [0:0] csa_component41_fa9_xor1;
  wire [0:0] csa_component41_fa9_or0;
  wire [0:0] csa_component41_fa10_xor1;
  wire [0:0] csa_component41_fa10_or0;
  wire [0:0] csa_component41_fa11_xor1;
  wire [0:0] csa_component41_fa11_or0;
  wire [0:0] csa_component41_fa12_xor1;
  wire [0:0] csa_component41_fa12_or0;
  wire [0:0] csa_component41_fa13_xor1;
  wire [0:0] csa_component41_fa13_or0;
  wire [0:0] csa_component41_fa14_xor1;
  wire [0:0] csa_component41_fa14_or0;
  wire [0:0] csa_component41_fa15_xor1;
  wire [0:0] csa_component41_fa15_or0;
  wire [0:0] csa_component41_fa16_xor1;
  wire [0:0] csa_component41_fa16_or0;
  wire [0:0] csa_component41_fa17_xor1;
  wire [0:0] csa_component41_fa17_or0;
  wire [0:0] csa_component41_fa18_xor1;
  wire [0:0] csa_component41_fa18_or0;
  wire [0:0] csa_component41_fa19_xor1;
  wire [0:0] csa_component41_fa19_or0;
  wire [0:0] csa_component41_fa20_xor1;
  wire [0:0] csa_component41_fa20_or0;
  wire [0:0] csa_component41_fa21_xor1;
  wire [0:0] csa_component41_fa21_or0;
  wire [0:0] csa_component41_fa22_xor1;
  wire [0:0] csa_component41_fa22_or0;
  wire [0:0] csa_component41_fa23_xor1;
  wire [0:0] csa_component41_fa23_or0;
  wire [0:0] csa_component41_fa24_xor1;
  wire [0:0] csa_component41_fa24_or0;
  wire [0:0] csa_component41_fa25_xor1;
  wire [0:0] csa_component41_fa25_or0;
  wire [0:0] csa_component41_fa26_xor1;
  wire [0:0] csa_component41_fa26_or0;
  wire [0:0] csa_component41_fa27_xor1;
  wire [0:0] csa_component41_fa27_or0;
  wire [0:0] csa_component41_fa28_xor1;
  wire [0:0] csa_component41_fa28_or0;
  wire [0:0] csa_component41_fa29_xor1;
  wire [0:0] csa_component41_fa29_or0;
  wire [0:0] csa_component41_fa30_xor1;
  wire [0:0] csa_component41_fa30_or0;
  wire [0:0] csa_component41_fa31_xor1;
  wire [0:0] csa_component41_fa31_or0;
  wire [0:0] csa_component41_fa32_xor1;
  wire [0:0] csa_component41_fa32_or0;
  wire [0:0] csa_component41_fa33_xor1;
  wire [0:0] csa_component41_fa33_or0;
  wire [0:0] csa_component41_fa34_xor1;
  wire [0:0] csa_component41_fa34_or0;
  wire [0:0] csa_component41_fa35_xor1;
  wire [0:0] csa_component41_fa35_or0;
  wire [0:0] csa_component41_fa36_xor1;
  wire [0:0] csa_component41_fa36_or0;
  wire [0:0] csa_component41_fa37_xor1;
  wire [0:0] csa_component41_fa37_or0;
  wire [0:0] csa_component41_fa38_xor1;
  wire [0:0] csa_component41_fa38_or0;
  wire [0:0] csa_component41_fa39_xor1;
  wire [0:0] csa_component41_fa39_or0;
  wire [0:0] csa_component41_fa40_xor1;
  wire [0:0] csa_component41_fa40_or0;

  fa fa_csa_component41_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component41_fa0_xor1), .fa_or0(csa_component41_fa0_or0));
  fa fa_csa_component41_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component41_fa1_xor1), .fa_or0(csa_component41_fa1_or0));
  fa fa_csa_component41_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component41_fa2_xor1), .fa_or0(csa_component41_fa2_or0));
  fa fa_csa_component41_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component41_fa3_xor1), .fa_or0(csa_component41_fa3_or0));
  fa fa_csa_component41_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component41_fa4_xor1), .fa_or0(csa_component41_fa4_or0));
  fa fa_csa_component41_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component41_fa5_xor1), .fa_or0(csa_component41_fa5_or0));
  fa fa_csa_component41_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component41_fa6_xor1), .fa_or0(csa_component41_fa6_or0));
  fa fa_csa_component41_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component41_fa7_xor1), .fa_or0(csa_component41_fa7_or0));
  fa fa_csa_component41_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component41_fa8_xor1), .fa_or0(csa_component41_fa8_or0));
  fa fa_csa_component41_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component41_fa9_xor1), .fa_or0(csa_component41_fa9_or0));
  fa fa_csa_component41_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component41_fa10_xor1), .fa_or0(csa_component41_fa10_or0));
  fa fa_csa_component41_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component41_fa11_xor1), .fa_or0(csa_component41_fa11_or0));
  fa fa_csa_component41_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component41_fa12_xor1), .fa_or0(csa_component41_fa12_or0));
  fa fa_csa_component41_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component41_fa13_xor1), .fa_or0(csa_component41_fa13_or0));
  fa fa_csa_component41_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component41_fa14_xor1), .fa_or0(csa_component41_fa14_or0));
  fa fa_csa_component41_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component41_fa15_xor1), .fa_or0(csa_component41_fa15_or0));
  fa fa_csa_component41_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component41_fa16_xor1), .fa_or0(csa_component41_fa16_or0));
  fa fa_csa_component41_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component41_fa17_xor1), .fa_or0(csa_component41_fa17_or0));
  fa fa_csa_component41_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component41_fa18_xor1), .fa_or0(csa_component41_fa18_or0));
  fa fa_csa_component41_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component41_fa19_xor1), .fa_or0(csa_component41_fa19_or0));
  fa fa_csa_component41_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component41_fa20_xor1), .fa_or0(csa_component41_fa20_or0));
  fa fa_csa_component41_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component41_fa21_xor1), .fa_or0(csa_component41_fa21_or0));
  fa fa_csa_component41_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component41_fa22_xor1), .fa_or0(csa_component41_fa22_or0));
  fa fa_csa_component41_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component41_fa23_xor1), .fa_or0(csa_component41_fa23_or0));
  fa fa_csa_component41_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component41_fa24_xor1), .fa_or0(csa_component41_fa24_or0));
  fa fa_csa_component41_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component41_fa25_xor1), .fa_or0(csa_component41_fa25_or0));
  fa fa_csa_component41_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component41_fa26_xor1), .fa_or0(csa_component41_fa26_or0));
  fa fa_csa_component41_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component41_fa27_xor1), .fa_or0(csa_component41_fa27_or0));
  fa fa_csa_component41_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component41_fa28_xor1), .fa_or0(csa_component41_fa28_or0));
  fa fa_csa_component41_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component41_fa29_xor1), .fa_or0(csa_component41_fa29_or0));
  fa fa_csa_component41_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component41_fa30_xor1), .fa_or0(csa_component41_fa30_or0));
  fa fa_csa_component41_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component41_fa31_xor1), .fa_or0(csa_component41_fa31_or0));
  fa fa_csa_component41_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component41_fa32_xor1), .fa_or0(csa_component41_fa32_or0));
  fa fa_csa_component41_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component41_fa33_xor1), .fa_or0(csa_component41_fa33_or0));
  fa fa_csa_component41_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component41_fa34_xor1), .fa_or0(csa_component41_fa34_or0));
  fa fa_csa_component41_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component41_fa35_xor1), .fa_or0(csa_component41_fa35_or0));
  fa fa_csa_component41_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component41_fa36_xor1), .fa_or0(csa_component41_fa36_or0));
  fa fa_csa_component41_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component41_fa37_xor1), .fa_or0(csa_component41_fa37_or0));
  fa fa_csa_component41_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component41_fa38_xor1), .fa_or0(csa_component41_fa38_or0));
  fa fa_csa_component41_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component41_fa39_xor1), .fa_or0(csa_component41_fa39_or0));
  fa fa_csa_component41_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component41_fa40_xor1), .fa_or0(csa_component41_fa40_or0));

  assign csa_component41_out[0] = csa_component41_fa0_xor1[0];
  assign csa_component41_out[1] = csa_component41_fa1_xor1[0];
  assign csa_component41_out[2] = csa_component41_fa2_xor1[0];
  assign csa_component41_out[3] = csa_component41_fa3_xor1[0];
  assign csa_component41_out[4] = csa_component41_fa4_xor1[0];
  assign csa_component41_out[5] = csa_component41_fa5_xor1[0];
  assign csa_component41_out[6] = csa_component41_fa6_xor1[0];
  assign csa_component41_out[7] = csa_component41_fa7_xor1[0];
  assign csa_component41_out[8] = csa_component41_fa8_xor1[0];
  assign csa_component41_out[9] = csa_component41_fa9_xor1[0];
  assign csa_component41_out[10] = csa_component41_fa10_xor1[0];
  assign csa_component41_out[11] = csa_component41_fa11_xor1[0];
  assign csa_component41_out[12] = csa_component41_fa12_xor1[0];
  assign csa_component41_out[13] = csa_component41_fa13_xor1[0];
  assign csa_component41_out[14] = csa_component41_fa14_xor1[0];
  assign csa_component41_out[15] = csa_component41_fa15_xor1[0];
  assign csa_component41_out[16] = csa_component41_fa16_xor1[0];
  assign csa_component41_out[17] = csa_component41_fa17_xor1[0];
  assign csa_component41_out[18] = csa_component41_fa18_xor1[0];
  assign csa_component41_out[19] = csa_component41_fa19_xor1[0];
  assign csa_component41_out[20] = csa_component41_fa20_xor1[0];
  assign csa_component41_out[21] = csa_component41_fa21_xor1[0];
  assign csa_component41_out[22] = csa_component41_fa22_xor1[0];
  assign csa_component41_out[23] = csa_component41_fa23_xor1[0];
  assign csa_component41_out[24] = csa_component41_fa24_xor1[0];
  assign csa_component41_out[25] = csa_component41_fa25_xor1[0];
  assign csa_component41_out[26] = csa_component41_fa26_xor1[0];
  assign csa_component41_out[27] = csa_component41_fa27_xor1[0];
  assign csa_component41_out[28] = csa_component41_fa28_xor1[0];
  assign csa_component41_out[29] = csa_component41_fa29_xor1[0];
  assign csa_component41_out[30] = csa_component41_fa30_xor1[0];
  assign csa_component41_out[31] = csa_component41_fa31_xor1[0];
  assign csa_component41_out[32] = csa_component41_fa32_xor1[0];
  assign csa_component41_out[33] = csa_component41_fa33_xor1[0];
  assign csa_component41_out[34] = csa_component41_fa34_xor1[0];
  assign csa_component41_out[35] = csa_component41_fa35_xor1[0];
  assign csa_component41_out[36] = csa_component41_fa36_xor1[0];
  assign csa_component41_out[37] = csa_component41_fa37_xor1[0];
  assign csa_component41_out[38] = csa_component41_fa38_xor1[0];
  assign csa_component41_out[39] = csa_component41_fa39_xor1[0];
  assign csa_component41_out[40] = csa_component41_fa40_xor1[0];
  assign csa_component41_out[41] = 1'b0;
  assign csa_component41_out[42] = 1'b0;
  assign csa_component41_out[43] = csa_component41_fa0_or0[0];
  assign csa_component41_out[44] = csa_component41_fa1_or0[0];
  assign csa_component41_out[45] = csa_component41_fa2_or0[0];
  assign csa_component41_out[46] = csa_component41_fa3_or0[0];
  assign csa_component41_out[47] = csa_component41_fa4_or0[0];
  assign csa_component41_out[48] = csa_component41_fa5_or0[0];
  assign csa_component41_out[49] = csa_component41_fa6_or0[0];
  assign csa_component41_out[50] = csa_component41_fa7_or0[0];
  assign csa_component41_out[51] = csa_component41_fa8_or0[0];
  assign csa_component41_out[52] = csa_component41_fa9_or0[0];
  assign csa_component41_out[53] = csa_component41_fa10_or0[0];
  assign csa_component41_out[54] = csa_component41_fa11_or0[0];
  assign csa_component41_out[55] = csa_component41_fa12_or0[0];
  assign csa_component41_out[56] = csa_component41_fa13_or0[0];
  assign csa_component41_out[57] = csa_component41_fa14_or0[0];
  assign csa_component41_out[58] = csa_component41_fa15_or0[0];
  assign csa_component41_out[59] = csa_component41_fa16_or0[0];
  assign csa_component41_out[60] = csa_component41_fa17_or0[0];
  assign csa_component41_out[61] = csa_component41_fa18_or0[0];
  assign csa_component41_out[62] = csa_component41_fa19_or0[0];
  assign csa_component41_out[63] = csa_component41_fa20_or0[0];
  assign csa_component41_out[64] = csa_component41_fa21_or0[0];
  assign csa_component41_out[65] = csa_component41_fa22_or0[0];
  assign csa_component41_out[66] = csa_component41_fa23_or0[0];
  assign csa_component41_out[67] = csa_component41_fa24_or0[0];
  assign csa_component41_out[68] = csa_component41_fa25_or0[0];
  assign csa_component41_out[69] = csa_component41_fa26_or0[0];
  assign csa_component41_out[70] = csa_component41_fa27_or0[0];
  assign csa_component41_out[71] = csa_component41_fa28_or0[0];
  assign csa_component41_out[72] = csa_component41_fa29_or0[0];
  assign csa_component41_out[73] = csa_component41_fa30_or0[0];
  assign csa_component41_out[74] = csa_component41_fa31_or0[0];
  assign csa_component41_out[75] = csa_component41_fa32_or0[0];
  assign csa_component41_out[76] = csa_component41_fa33_or0[0];
  assign csa_component41_out[77] = csa_component41_fa34_or0[0];
  assign csa_component41_out[78] = csa_component41_fa35_or0[0];
  assign csa_component41_out[79] = csa_component41_fa36_or0[0];
  assign csa_component41_out[80] = csa_component41_fa37_or0[0];
  assign csa_component41_out[81] = csa_component41_fa38_or0[0];
  assign csa_component41_out[82] = csa_component41_fa39_or0[0];
  assign csa_component41_out[83] = csa_component41_fa40_or0[0];
endmodule

module csa_component47(input [46:0] a, input [46:0] b, input [46:0] c, output [95:0] csa_component47_out);
  wire [0:0] csa_component47_fa0_xor1;
  wire [0:0] csa_component47_fa0_or0;
  wire [0:0] csa_component47_fa1_xor1;
  wire [0:0] csa_component47_fa1_or0;
  wire [0:0] csa_component47_fa2_xor1;
  wire [0:0] csa_component47_fa2_or0;
  wire [0:0] csa_component47_fa3_xor1;
  wire [0:0] csa_component47_fa3_or0;
  wire [0:0] csa_component47_fa4_xor1;
  wire [0:0] csa_component47_fa4_or0;
  wire [0:0] csa_component47_fa5_xor1;
  wire [0:0] csa_component47_fa5_or0;
  wire [0:0] csa_component47_fa6_xor1;
  wire [0:0] csa_component47_fa6_or0;
  wire [0:0] csa_component47_fa7_xor1;
  wire [0:0] csa_component47_fa7_or0;
  wire [0:0] csa_component47_fa8_xor1;
  wire [0:0] csa_component47_fa8_or0;
  wire [0:0] csa_component47_fa9_xor1;
  wire [0:0] csa_component47_fa9_or0;
  wire [0:0] csa_component47_fa10_xor1;
  wire [0:0] csa_component47_fa10_or0;
  wire [0:0] csa_component47_fa11_xor1;
  wire [0:0] csa_component47_fa11_or0;
  wire [0:0] csa_component47_fa12_xor1;
  wire [0:0] csa_component47_fa12_or0;
  wire [0:0] csa_component47_fa13_xor1;
  wire [0:0] csa_component47_fa13_or0;
  wire [0:0] csa_component47_fa14_xor1;
  wire [0:0] csa_component47_fa14_or0;
  wire [0:0] csa_component47_fa15_xor1;
  wire [0:0] csa_component47_fa15_or0;
  wire [0:0] csa_component47_fa16_xor1;
  wire [0:0] csa_component47_fa16_or0;
  wire [0:0] csa_component47_fa17_xor1;
  wire [0:0] csa_component47_fa17_or0;
  wire [0:0] csa_component47_fa18_xor1;
  wire [0:0] csa_component47_fa18_or0;
  wire [0:0] csa_component47_fa19_xor1;
  wire [0:0] csa_component47_fa19_or0;
  wire [0:0] csa_component47_fa20_xor1;
  wire [0:0] csa_component47_fa20_or0;
  wire [0:0] csa_component47_fa21_xor1;
  wire [0:0] csa_component47_fa21_or0;
  wire [0:0] csa_component47_fa22_xor1;
  wire [0:0] csa_component47_fa22_or0;
  wire [0:0] csa_component47_fa23_xor1;
  wire [0:0] csa_component47_fa23_or0;
  wire [0:0] csa_component47_fa24_xor1;
  wire [0:0] csa_component47_fa24_or0;
  wire [0:0] csa_component47_fa25_xor1;
  wire [0:0] csa_component47_fa25_or0;
  wire [0:0] csa_component47_fa26_xor1;
  wire [0:0] csa_component47_fa26_or0;
  wire [0:0] csa_component47_fa27_xor1;
  wire [0:0] csa_component47_fa27_or0;
  wire [0:0] csa_component47_fa28_xor1;
  wire [0:0] csa_component47_fa28_or0;
  wire [0:0] csa_component47_fa29_xor1;
  wire [0:0] csa_component47_fa29_or0;
  wire [0:0] csa_component47_fa30_xor1;
  wire [0:0] csa_component47_fa30_or0;
  wire [0:0] csa_component47_fa31_xor1;
  wire [0:0] csa_component47_fa31_or0;
  wire [0:0] csa_component47_fa32_xor1;
  wire [0:0] csa_component47_fa32_or0;
  wire [0:0] csa_component47_fa33_xor1;
  wire [0:0] csa_component47_fa33_or0;
  wire [0:0] csa_component47_fa34_xor1;
  wire [0:0] csa_component47_fa34_or0;
  wire [0:0] csa_component47_fa35_xor1;
  wire [0:0] csa_component47_fa35_or0;
  wire [0:0] csa_component47_fa36_xor1;
  wire [0:0] csa_component47_fa36_or0;
  wire [0:0] csa_component47_fa37_xor1;
  wire [0:0] csa_component47_fa37_or0;
  wire [0:0] csa_component47_fa38_xor1;
  wire [0:0] csa_component47_fa38_or0;
  wire [0:0] csa_component47_fa39_xor1;
  wire [0:0] csa_component47_fa39_or0;
  wire [0:0] csa_component47_fa40_xor1;
  wire [0:0] csa_component47_fa40_or0;
  wire [0:0] csa_component47_fa41_xor1;
  wire [0:0] csa_component47_fa41_or0;
  wire [0:0] csa_component47_fa42_xor1;
  wire [0:0] csa_component47_fa42_or0;
  wire [0:0] csa_component47_fa43_xor1;
  wire [0:0] csa_component47_fa43_or0;
  wire [0:0] csa_component47_fa44_xor1;
  wire [0:0] csa_component47_fa44_or0;
  wire [0:0] csa_component47_fa45_xor1;
  wire [0:0] csa_component47_fa45_or0;
  wire [0:0] csa_component47_fa46_xor1;
  wire [0:0] csa_component47_fa46_or0;

  fa fa_csa_component47_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component47_fa0_xor1), .fa_or0(csa_component47_fa0_or0));
  fa fa_csa_component47_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component47_fa1_xor1), .fa_or0(csa_component47_fa1_or0));
  fa fa_csa_component47_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component47_fa2_xor1), .fa_or0(csa_component47_fa2_or0));
  fa fa_csa_component47_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component47_fa3_xor1), .fa_or0(csa_component47_fa3_or0));
  fa fa_csa_component47_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component47_fa4_xor1), .fa_or0(csa_component47_fa4_or0));
  fa fa_csa_component47_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component47_fa5_xor1), .fa_or0(csa_component47_fa5_or0));
  fa fa_csa_component47_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component47_fa6_xor1), .fa_or0(csa_component47_fa6_or0));
  fa fa_csa_component47_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component47_fa7_xor1), .fa_or0(csa_component47_fa7_or0));
  fa fa_csa_component47_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component47_fa8_xor1), .fa_or0(csa_component47_fa8_or0));
  fa fa_csa_component47_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component47_fa9_xor1), .fa_or0(csa_component47_fa9_or0));
  fa fa_csa_component47_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component47_fa10_xor1), .fa_or0(csa_component47_fa10_or0));
  fa fa_csa_component47_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component47_fa11_xor1), .fa_or0(csa_component47_fa11_or0));
  fa fa_csa_component47_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component47_fa12_xor1), .fa_or0(csa_component47_fa12_or0));
  fa fa_csa_component47_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component47_fa13_xor1), .fa_or0(csa_component47_fa13_or0));
  fa fa_csa_component47_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component47_fa14_xor1), .fa_or0(csa_component47_fa14_or0));
  fa fa_csa_component47_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component47_fa15_xor1), .fa_or0(csa_component47_fa15_or0));
  fa fa_csa_component47_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component47_fa16_xor1), .fa_or0(csa_component47_fa16_or0));
  fa fa_csa_component47_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component47_fa17_xor1), .fa_or0(csa_component47_fa17_or0));
  fa fa_csa_component47_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component47_fa18_xor1), .fa_or0(csa_component47_fa18_or0));
  fa fa_csa_component47_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component47_fa19_xor1), .fa_or0(csa_component47_fa19_or0));
  fa fa_csa_component47_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component47_fa20_xor1), .fa_or0(csa_component47_fa20_or0));
  fa fa_csa_component47_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component47_fa21_xor1), .fa_or0(csa_component47_fa21_or0));
  fa fa_csa_component47_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component47_fa22_xor1), .fa_or0(csa_component47_fa22_or0));
  fa fa_csa_component47_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component47_fa23_xor1), .fa_or0(csa_component47_fa23_or0));
  fa fa_csa_component47_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component47_fa24_xor1), .fa_or0(csa_component47_fa24_or0));
  fa fa_csa_component47_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component47_fa25_xor1), .fa_or0(csa_component47_fa25_or0));
  fa fa_csa_component47_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component47_fa26_xor1), .fa_or0(csa_component47_fa26_or0));
  fa fa_csa_component47_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component47_fa27_xor1), .fa_or0(csa_component47_fa27_or0));
  fa fa_csa_component47_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component47_fa28_xor1), .fa_or0(csa_component47_fa28_or0));
  fa fa_csa_component47_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component47_fa29_xor1), .fa_or0(csa_component47_fa29_or0));
  fa fa_csa_component47_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component47_fa30_xor1), .fa_or0(csa_component47_fa30_or0));
  fa fa_csa_component47_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component47_fa31_xor1), .fa_or0(csa_component47_fa31_or0));
  fa fa_csa_component47_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component47_fa32_xor1), .fa_or0(csa_component47_fa32_or0));
  fa fa_csa_component47_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component47_fa33_xor1), .fa_or0(csa_component47_fa33_or0));
  fa fa_csa_component47_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component47_fa34_xor1), .fa_or0(csa_component47_fa34_or0));
  fa fa_csa_component47_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component47_fa35_xor1), .fa_or0(csa_component47_fa35_or0));
  fa fa_csa_component47_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component47_fa36_xor1), .fa_or0(csa_component47_fa36_or0));
  fa fa_csa_component47_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component47_fa37_xor1), .fa_or0(csa_component47_fa37_or0));
  fa fa_csa_component47_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component47_fa38_xor1), .fa_or0(csa_component47_fa38_or0));
  fa fa_csa_component47_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component47_fa39_xor1), .fa_or0(csa_component47_fa39_or0));
  fa fa_csa_component47_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component47_fa40_xor1), .fa_or0(csa_component47_fa40_or0));
  fa fa_csa_component47_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component47_fa41_xor1), .fa_or0(csa_component47_fa41_or0));
  fa fa_csa_component47_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component47_fa42_xor1), .fa_or0(csa_component47_fa42_or0));
  fa fa_csa_component47_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component47_fa43_xor1), .fa_or0(csa_component47_fa43_or0));
  fa fa_csa_component47_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component47_fa44_xor1), .fa_or0(csa_component47_fa44_or0));
  fa fa_csa_component47_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component47_fa45_xor1), .fa_or0(csa_component47_fa45_or0));
  fa fa_csa_component47_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component47_fa46_xor1), .fa_or0(csa_component47_fa46_or0));

  assign csa_component47_out[0] = csa_component47_fa0_xor1[0];
  assign csa_component47_out[1] = csa_component47_fa1_xor1[0];
  assign csa_component47_out[2] = csa_component47_fa2_xor1[0];
  assign csa_component47_out[3] = csa_component47_fa3_xor1[0];
  assign csa_component47_out[4] = csa_component47_fa4_xor1[0];
  assign csa_component47_out[5] = csa_component47_fa5_xor1[0];
  assign csa_component47_out[6] = csa_component47_fa6_xor1[0];
  assign csa_component47_out[7] = csa_component47_fa7_xor1[0];
  assign csa_component47_out[8] = csa_component47_fa8_xor1[0];
  assign csa_component47_out[9] = csa_component47_fa9_xor1[0];
  assign csa_component47_out[10] = csa_component47_fa10_xor1[0];
  assign csa_component47_out[11] = csa_component47_fa11_xor1[0];
  assign csa_component47_out[12] = csa_component47_fa12_xor1[0];
  assign csa_component47_out[13] = csa_component47_fa13_xor1[0];
  assign csa_component47_out[14] = csa_component47_fa14_xor1[0];
  assign csa_component47_out[15] = csa_component47_fa15_xor1[0];
  assign csa_component47_out[16] = csa_component47_fa16_xor1[0];
  assign csa_component47_out[17] = csa_component47_fa17_xor1[0];
  assign csa_component47_out[18] = csa_component47_fa18_xor1[0];
  assign csa_component47_out[19] = csa_component47_fa19_xor1[0];
  assign csa_component47_out[20] = csa_component47_fa20_xor1[0];
  assign csa_component47_out[21] = csa_component47_fa21_xor1[0];
  assign csa_component47_out[22] = csa_component47_fa22_xor1[0];
  assign csa_component47_out[23] = csa_component47_fa23_xor1[0];
  assign csa_component47_out[24] = csa_component47_fa24_xor1[0];
  assign csa_component47_out[25] = csa_component47_fa25_xor1[0];
  assign csa_component47_out[26] = csa_component47_fa26_xor1[0];
  assign csa_component47_out[27] = csa_component47_fa27_xor1[0];
  assign csa_component47_out[28] = csa_component47_fa28_xor1[0];
  assign csa_component47_out[29] = csa_component47_fa29_xor1[0];
  assign csa_component47_out[30] = csa_component47_fa30_xor1[0];
  assign csa_component47_out[31] = csa_component47_fa31_xor1[0];
  assign csa_component47_out[32] = csa_component47_fa32_xor1[0];
  assign csa_component47_out[33] = csa_component47_fa33_xor1[0];
  assign csa_component47_out[34] = csa_component47_fa34_xor1[0];
  assign csa_component47_out[35] = csa_component47_fa35_xor1[0];
  assign csa_component47_out[36] = csa_component47_fa36_xor1[0];
  assign csa_component47_out[37] = csa_component47_fa37_xor1[0];
  assign csa_component47_out[38] = csa_component47_fa38_xor1[0];
  assign csa_component47_out[39] = csa_component47_fa39_xor1[0];
  assign csa_component47_out[40] = csa_component47_fa40_xor1[0];
  assign csa_component47_out[41] = csa_component47_fa41_xor1[0];
  assign csa_component47_out[42] = csa_component47_fa42_xor1[0];
  assign csa_component47_out[43] = csa_component47_fa43_xor1[0];
  assign csa_component47_out[44] = csa_component47_fa44_xor1[0];
  assign csa_component47_out[45] = csa_component47_fa45_xor1[0];
  assign csa_component47_out[46] = csa_component47_fa46_xor1[0];
  assign csa_component47_out[47] = 1'b0;
  assign csa_component47_out[48] = 1'b0;
  assign csa_component47_out[49] = csa_component47_fa0_or0[0];
  assign csa_component47_out[50] = csa_component47_fa1_or0[0];
  assign csa_component47_out[51] = csa_component47_fa2_or0[0];
  assign csa_component47_out[52] = csa_component47_fa3_or0[0];
  assign csa_component47_out[53] = csa_component47_fa4_or0[0];
  assign csa_component47_out[54] = csa_component47_fa5_or0[0];
  assign csa_component47_out[55] = csa_component47_fa6_or0[0];
  assign csa_component47_out[56] = csa_component47_fa7_or0[0];
  assign csa_component47_out[57] = csa_component47_fa8_or0[0];
  assign csa_component47_out[58] = csa_component47_fa9_or0[0];
  assign csa_component47_out[59] = csa_component47_fa10_or0[0];
  assign csa_component47_out[60] = csa_component47_fa11_or0[0];
  assign csa_component47_out[61] = csa_component47_fa12_or0[0];
  assign csa_component47_out[62] = csa_component47_fa13_or0[0];
  assign csa_component47_out[63] = csa_component47_fa14_or0[0];
  assign csa_component47_out[64] = csa_component47_fa15_or0[0];
  assign csa_component47_out[65] = csa_component47_fa16_or0[0];
  assign csa_component47_out[66] = csa_component47_fa17_or0[0];
  assign csa_component47_out[67] = csa_component47_fa18_or0[0];
  assign csa_component47_out[68] = csa_component47_fa19_or0[0];
  assign csa_component47_out[69] = csa_component47_fa20_or0[0];
  assign csa_component47_out[70] = csa_component47_fa21_or0[0];
  assign csa_component47_out[71] = csa_component47_fa22_or0[0];
  assign csa_component47_out[72] = csa_component47_fa23_or0[0];
  assign csa_component47_out[73] = csa_component47_fa24_or0[0];
  assign csa_component47_out[74] = csa_component47_fa25_or0[0];
  assign csa_component47_out[75] = csa_component47_fa26_or0[0];
  assign csa_component47_out[76] = csa_component47_fa27_or0[0];
  assign csa_component47_out[77] = csa_component47_fa28_or0[0];
  assign csa_component47_out[78] = csa_component47_fa29_or0[0];
  assign csa_component47_out[79] = csa_component47_fa30_or0[0];
  assign csa_component47_out[80] = csa_component47_fa31_or0[0];
  assign csa_component47_out[81] = csa_component47_fa32_or0[0];
  assign csa_component47_out[82] = csa_component47_fa33_or0[0];
  assign csa_component47_out[83] = csa_component47_fa34_or0[0];
  assign csa_component47_out[84] = csa_component47_fa35_or0[0];
  assign csa_component47_out[85] = csa_component47_fa36_or0[0];
  assign csa_component47_out[86] = csa_component47_fa37_or0[0];
  assign csa_component47_out[87] = csa_component47_fa38_or0[0];
  assign csa_component47_out[88] = csa_component47_fa39_or0[0];
  assign csa_component47_out[89] = csa_component47_fa40_or0[0];
  assign csa_component47_out[90] = csa_component47_fa41_or0[0];
  assign csa_component47_out[91] = csa_component47_fa42_or0[0];
  assign csa_component47_out[92] = csa_component47_fa43_or0[0];
  assign csa_component47_out[93] = csa_component47_fa44_or0[0];
  assign csa_component47_out[94] = csa_component47_fa45_or0[0];
  assign csa_component47_out[95] = csa_component47_fa46_or0[0];
endmodule

module csa_component50(input [49:0] a, input [49:0] b, input [49:0] c, output [101:0] csa_component50_out);
  wire [0:0] csa_component50_fa0_xor1;
  wire [0:0] csa_component50_fa0_or0;
  wire [0:0] csa_component50_fa1_xor1;
  wire [0:0] csa_component50_fa1_or0;
  wire [0:0] csa_component50_fa2_xor1;
  wire [0:0] csa_component50_fa2_or0;
  wire [0:0] csa_component50_fa3_xor1;
  wire [0:0] csa_component50_fa3_or0;
  wire [0:0] csa_component50_fa4_xor1;
  wire [0:0] csa_component50_fa4_or0;
  wire [0:0] csa_component50_fa5_xor1;
  wire [0:0] csa_component50_fa5_or0;
  wire [0:0] csa_component50_fa6_xor1;
  wire [0:0] csa_component50_fa6_or0;
  wire [0:0] csa_component50_fa7_xor1;
  wire [0:0] csa_component50_fa7_or0;
  wire [0:0] csa_component50_fa8_xor1;
  wire [0:0] csa_component50_fa8_or0;
  wire [0:0] csa_component50_fa9_xor1;
  wire [0:0] csa_component50_fa9_or0;
  wire [0:0] csa_component50_fa10_xor1;
  wire [0:0] csa_component50_fa10_or0;
  wire [0:0] csa_component50_fa11_xor1;
  wire [0:0] csa_component50_fa11_or0;
  wire [0:0] csa_component50_fa12_xor1;
  wire [0:0] csa_component50_fa12_or0;
  wire [0:0] csa_component50_fa13_xor1;
  wire [0:0] csa_component50_fa13_or0;
  wire [0:0] csa_component50_fa14_xor1;
  wire [0:0] csa_component50_fa14_or0;
  wire [0:0] csa_component50_fa15_xor1;
  wire [0:0] csa_component50_fa15_or0;
  wire [0:0] csa_component50_fa16_xor1;
  wire [0:0] csa_component50_fa16_or0;
  wire [0:0] csa_component50_fa17_xor1;
  wire [0:0] csa_component50_fa17_or0;
  wire [0:0] csa_component50_fa18_xor1;
  wire [0:0] csa_component50_fa18_or0;
  wire [0:0] csa_component50_fa19_xor1;
  wire [0:0] csa_component50_fa19_or0;
  wire [0:0] csa_component50_fa20_xor1;
  wire [0:0] csa_component50_fa20_or0;
  wire [0:0] csa_component50_fa21_xor1;
  wire [0:0] csa_component50_fa21_or0;
  wire [0:0] csa_component50_fa22_xor1;
  wire [0:0] csa_component50_fa22_or0;
  wire [0:0] csa_component50_fa23_xor1;
  wire [0:0] csa_component50_fa23_or0;
  wire [0:0] csa_component50_fa24_xor1;
  wire [0:0] csa_component50_fa24_or0;
  wire [0:0] csa_component50_fa25_xor1;
  wire [0:0] csa_component50_fa25_or0;
  wire [0:0] csa_component50_fa26_xor1;
  wire [0:0] csa_component50_fa26_or0;
  wire [0:0] csa_component50_fa27_xor1;
  wire [0:0] csa_component50_fa27_or0;
  wire [0:0] csa_component50_fa28_xor1;
  wire [0:0] csa_component50_fa28_or0;
  wire [0:0] csa_component50_fa29_xor1;
  wire [0:0] csa_component50_fa29_or0;
  wire [0:0] csa_component50_fa30_xor1;
  wire [0:0] csa_component50_fa30_or0;
  wire [0:0] csa_component50_fa31_xor1;
  wire [0:0] csa_component50_fa31_or0;
  wire [0:0] csa_component50_fa32_xor1;
  wire [0:0] csa_component50_fa32_or0;
  wire [0:0] csa_component50_fa33_xor1;
  wire [0:0] csa_component50_fa33_or0;
  wire [0:0] csa_component50_fa34_xor1;
  wire [0:0] csa_component50_fa34_or0;
  wire [0:0] csa_component50_fa35_xor1;
  wire [0:0] csa_component50_fa35_or0;
  wire [0:0] csa_component50_fa36_xor1;
  wire [0:0] csa_component50_fa36_or0;
  wire [0:0] csa_component50_fa37_xor1;
  wire [0:0] csa_component50_fa37_or0;
  wire [0:0] csa_component50_fa38_xor1;
  wire [0:0] csa_component50_fa38_or0;
  wire [0:0] csa_component50_fa39_xor1;
  wire [0:0] csa_component50_fa39_or0;
  wire [0:0] csa_component50_fa40_xor1;
  wire [0:0] csa_component50_fa40_or0;
  wire [0:0] csa_component50_fa41_xor1;
  wire [0:0] csa_component50_fa41_or0;
  wire [0:0] csa_component50_fa42_xor1;
  wire [0:0] csa_component50_fa42_or0;
  wire [0:0] csa_component50_fa43_xor1;
  wire [0:0] csa_component50_fa43_or0;
  wire [0:0] csa_component50_fa44_xor1;
  wire [0:0] csa_component50_fa44_or0;
  wire [0:0] csa_component50_fa45_xor1;
  wire [0:0] csa_component50_fa45_or0;
  wire [0:0] csa_component50_fa46_xor1;
  wire [0:0] csa_component50_fa46_or0;
  wire [0:0] csa_component50_fa47_xor1;
  wire [0:0] csa_component50_fa47_or0;
  wire [0:0] csa_component50_fa48_xor1;
  wire [0:0] csa_component50_fa48_or0;
  wire [0:0] csa_component50_fa49_xor1;
  wire [0:0] csa_component50_fa49_or0;

  fa fa_csa_component50_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component50_fa0_xor1), .fa_or0(csa_component50_fa0_or0));
  fa fa_csa_component50_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component50_fa1_xor1), .fa_or0(csa_component50_fa1_or0));
  fa fa_csa_component50_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component50_fa2_xor1), .fa_or0(csa_component50_fa2_or0));
  fa fa_csa_component50_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component50_fa3_xor1), .fa_or0(csa_component50_fa3_or0));
  fa fa_csa_component50_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component50_fa4_xor1), .fa_or0(csa_component50_fa4_or0));
  fa fa_csa_component50_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component50_fa5_xor1), .fa_or0(csa_component50_fa5_or0));
  fa fa_csa_component50_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component50_fa6_xor1), .fa_or0(csa_component50_fa6_or0));
  fa fa_csa_component50_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component50_fa7_xor1), .fa_or0(csa_component50_fa7_or0));
  fa fa_csa_component50_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component50_fa8_xor1), .fa_or0(csa_component50_fa8_or0));
  fa fa_csa_component50_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component50_fa9_xor1), .fa_or0(csa_component50_fa9_or0));
  fa fa_csa_component50_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component50_fa10_xor1), .fa_or0(csa_component50_fa10_or0));
  fa fa_csa_component50_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component50_fa11_xor1), .fa_or0(csa_component50_fa11_or0));
  fa fa_csa_component50_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component50_fa12_xor1), .fa_or0(csa_component50_fa12_or0));
  fa fa_csa_component50_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component50_fa13_xor1), .fa_or0(csa_component50_fa13_or0));
  fa fa_csa_component50_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component50_fa14_xor1), .fa_or0(csa_component50_fa14_or0));
  fa fa_csa_component50_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component50_fa15_xor1), .fa_or0(csa_component50_fa15_or0));
  fa fa_csa_component50_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component50_fa16_xor1), .fa_or0(csa_component50_fa16_or0));
  fa fa_csa_component50_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component50_fa17_xor1), .fa_or0(csa_component50_fa17_or0));
  fa fa_csa_component50_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component50_fa18_xor1), .fa_or0(csa_component50_fa18_or0));
  fa fa_csa_component50_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component50_fa19_xor1), .fa_or0(csa_component50_fa19_or0));
  fa fa_csa_component50_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component50_fa20_xor1), .fa_or0(csa_component50_fa20_or0));
  fa fa_csa_component50_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component50_fa21_xor1), .fa_or0(csa_component50_fa21_or0));
  fa fa_csa_component50_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component50_fa22_xor1), .fa_or0(csa_component50_fa22_or0));
  fa fa_csa_component50_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component50_fa23_xor1), .fa_or0(csa_component50_fa23_or0));
  fa fa_csa_component50_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component50_fa24_xor1), .fa_or0(csa_component50_fa24_or0));
  fa fa_csa_component50_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component50_fa25_xor1), .fa_or0(csa_component50_fa25_or0));
  fa fa_csa_component50_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component50_fa26_xor1), .fa_or0(csa_component50_fa26_or0));
  fa fa_csa_component50_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component50_fa27_xor1), .fa_or0(csa_component50_fa27_or0));
  fa fa_csa_component50_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component50_fa28_xor1), .fa_or0(csa_component50_fa28_or0));
  fa fa_csa_component50_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component50_fa29_xor1), .fa_or0(csa_component50_fa29_or0));
  fa fa_csa_component50_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component50_fa30_xor1), .fa_or0(csa_component50_fa30_or0));
  fa fa_csa_component50_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component50_fa31_xor1), .fa_or0(csa_component50_fa31_or0));
  fa fa_csa_component50_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component50_fa32_xor1), .fa_or0(csa_component50_fa32_or0));
  fa fa_csa_component50_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component50_fa33_xor1), .fa_or0(csa_component50_fa33_or0));
  fa fa_csa_component50_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component50_fa34_xor1), .fa_or0(csa_component50_fa34_or0));
  fa fa_csa_component50_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component50_fa35_xor1), .fa_or0(csa_component50_fa35_or0));
  fa fa_csa_component50_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component50_fa36_xor1), .fa_or0(csa_component50_fa36_or0));
  fa fa_csa_component50_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component50_fa37_xor1), .fa_or0(csa_component50_fa37_or0));
  fa fa_csa_component50_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component50_fa38_xor1), .fa_or0(csa_component50_fa38_or0));
  fa fa_csa_component50_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component50_fa39_xor1), .fa_or0(csa_component50_fa39_or0));
  fa fa_csa_component50_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component50_fa40_xor1), .fa_or0(csa_component50_fa40_or0));
  fa fa_csa_component50_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component50_fa41_xor1), .fa_or0(csa_component50_fa41_or0));
  fa fa_csa_component50_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component50_fa42_xor1), .fa_or0(csa_component50_fa42_or0));
  fa fa_csa_component50_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component50_fa43_xor1), .fa_or0(csa_component50_fa43_or0));
  fa fa_csa_component50_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component50_fa44_xor1), .fa_or0(csa_component50_fa44_or0));
  fa fa_csa_component50_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component50_fa45_xor1), .fa_or0(csa_component50_fa45_or0));
  fa fa_csa_component50_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component50_fa46_xor1), .fa_or0(csa_component50_fa46_or0));
  fa fa_csa_component50_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component50_fa47_xor1), .fa_or0(csa_component50_fa47_or0));
  fa fa_csa_component50_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component50_fa48_xor1), .fa_or0(csa_component50_fa48_or0));
  fa fa_csa_component50_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component50_fa49_xor1), .fa_or0(csa_component50_fa49_or0));

  assign csa_component50_out[0] = csa_component50_fa0_xor1[0];
  assign csa_component50_out[1] = csa_component50_fa1_xor1[0];
  assign csa_component50_out[2] = csa_component50_fa2_xor1[0];
  assign csa_component50_out[3] = csa_component50_fa3_xor1[0];
  assign csa_component50_out[4] = csa_component50_fa4_xor1[0];
  assign csa_component50_out[5] = csa_component50_fa5_xor1[0];
  assign csa_component50_out[6] = csa_component50_fa6_xor1[0];
  assign csa_component50_out[7] = csa_component50_fa7_xor1[0];
  assign csa_component50_out[8] = csa_component50_fa8_xor1[0];
  assign csa_component50_out[9] = csa_component50_fa9_xor1[0];
  assign csa_component50_out[10] = csa_component50_fa10_xor1[0];
  assign csa_component50_out[11] = csa_component50_fa11_xor1[0];
  assign csa_component50_out[12] = csa_component50_fa12_xor1[0];
  assign csa_component50_out[13] = csa_component50_fa13_xor1[0];
  assign csa_component50_out[14] = csa_component50_fa14_xor1[0];
  assign csa_component50_out[15] = csa_component50_fa15_xor1[0];
  assign csa_component50_out[16] = csa_component50_fa16_xor1[0];
  assign csa_component50_out[17] = csa_component50_fa17_xor1[0];
  assign csa_component50_out[18] = csa_component50_fa18_xor1[0];
  assign csa_component50_out[19] = csa_component50_fa19_xor1[0];
  assign csa_component50_out[20] = csa_component50_fa20_xor1[0];
  assign csa_component50_out[21] = csa_component50_fa21_xor1[0];
  assign csa_component50_out[22] = csa_component50_fa22_xor1[0];
  assign csa_component50_out[23] = csa_component50_fa23_xor1[0];
  assign csa_component50_out[24] = csa_component50_fa24_xor1[0];
  assign csa_component50_out[25] = csa_component50_fa25_xor1[0];
  assign csa_component50_out[26] = csa_component50_fa26_xor1[0];
  assign csa_component50_out[27] = csa_component50_fa27_xor1[0];
  assign csa_component50_out[28] = csa_component50_fa28_xor1[0];
  assign csa_component50_out[29] = csa_component50_fa29_xor1[0];
  assign csa_component50_out[30] = csa_component50_fa30_xor1[0];
  assign csa_component50_out[31] = csa_component50_fa31_xor1[0];
  assign csa_component50_out[32] = csa_component50_fa32_xor1[0];
  assign csa_component50_out[33] = csa_component50_fa33_xor1[0];
  assign csa_component50_out[34] = csa_component50_fa34_xor1[0];
  assign csa_component50_out[35] = csa_component50_fa35_xor1[0];
  assign csa_component50_out[36] = csa_component50_fa36_xor1[0];
  assign csa_component50_out[37] = csa_component50_fa37_xor1[0];
  assign csa_component50_out[38] = csa_component50_fa38_xor1[0];
  assign csa_component50_out[39] = csa_component50_fa39_xor1[0];
  assign csa_component50_out[40] = csa_component50_fa40_xor1[0];
  assign csa_component50_out[41] = csa_component50_fa41_xor1[0];
  assign csa_component50_out[42] = csa_component50_fa42_xor1[0];
  assign csa_component50_out[43] = csa_component50_fa43_xor1[0];
  assign csa_component50_out[44] = csa_component50_fa44_xor1[0];
  assign csa_component50_out[45] = csa_component50_fa45_xor1[0];
  assign csa_component50_out[46] = csa_component50_fa46_xor1[0];
  assign csa_component50_out[47] = csa_component50_fa47_xor1[0];
  assign csa_component50_out[48] = csa_component50_fa48_xor1[0];
  assign csa_component50_out[49] = csa_component50_fa49_xor1[0];
  assign csa_component50_out[50] = 1'b0;
  assign csa_component50_out[51] = 1'b0;
  assign csa_component50_out[52] = csa_component50_fa0_or0[0];
  assign csa_component50_out[53] = csa_component50_fa1_or0[0];
  assign csa_component50_out[54] = csa_component50_fa2_or0[0];
  assign csa_component50_out[55] = csa_component50_fa3_or0[0];
  assign csa_component50_out[56] = csa_component50_fa4_or0[0];
  assign csa_component50_out[57] = csa_component50_fa5_or0[0];
  assign csa_component50_out[58] = csa_component50_fa6_or0[0];
  assign csa_component50_out[59] = csa_component50_fa7_or0[0];
  assign csa_component50_out[60] = csa_component50_fa8_or0[0];
  assign csa_component50_out[61] = csa_component50_fa9_or0[0];
  assign csa_component50_out[62] = csa_component50_fa10_or0[0];
  assign csa_component50_out[63] = csa_component50_fa11_or0[0];
  assign csa_component50_out[64] = csa_component50_fa12_or0[0];
  assign csa_component50_out[65] = csa_component50_fa13_or0[0];
  assign csa_component50_out[66] = csa_component50_fa14_or0[0];
  assign csa_component50_out[67] = csa_component50_fa15_or0[0];
  assign csa_component50_out[68] = csa_component50_fa16_or0[0];
  assign csa_component50_out[69] = csa_component50_fa17_or0[0];
  assign csa_component50_out[70] = csa_component50_fa18_or0[0];
  assign csa_component50_out[71] = csa_component50_fa19_or0[0];
  assign csa_component50_out[72] = csa_component50_fa20_or0[0];
  assign csa_component50_out[73] = csa_component50_fa21_or0[0];
  assign csa_component50_out[74] = csa_component50_fa22_or0[0];
  assign csa_component50_out[75] = csa_component50_fa23_or0[0];
  assign csa_component50_out[76] = csa_component50_fa24_or0[0];
  assign csa_component50_out[77] = csa_component50_fa25_or0[0];
  assign csa_component50_out[78] = csa_component50_fa26_or0[0];
  assign csa_component50_out[79] = csa_component50_fa27_or0[0];
  assign csa_component50_out[80] = csa_component50_fa28_or0[0];
  assign csa_component50_out[81] = csa_component50_fa29_or0[0];
  assign csa_component50_out[82] = csa_component50_fa30_or0[0];
  assign csa_component50_out[83] = csa_component50_fa31_or0[0];
  assign csa_component50_out[84] = csa_component50_fa32_or0[0];
  assign csa_component50_out[85] = csa_component50_fa33_or0[0];
  assign csa_component50_out[86] = csa_component50_fa34_or0[0];
  assign csa_component50_out[87] = csa_component50_fa35_or0[0];
  assign csa_component50_out[88] = csa_component50_fa36_or0[0];
  assign csa_component50_out[89] = csa_component50_fa37_or0[0];
  assign csa_component50_out[90] = csa_component50_fa38_or0[0];
  assign csa_component50_out[91] = csa_component50_fa39_or0[0];
  assign csa_component50_out[92] = csa_component50_fa40_or0[0];
  assign csa_component50_out[93] = csa_component50_fa41_or0[0];
  assign csa_component50_out[94] = csa_component50_fa42_or0[0];
  assign csa_component50_out[95] = csa_component50_fa43_or0[0];
  assign csa_component50_out[96] = csa_component50_fa44_or0[0];
  assign csa_component50_out[97] = csa_component50_fa45_or0[0];
  assign csa_component50_out[98] = csa_component50_fa46_or0[0];
  assign csa_component50_out[99] = csa_component50_fa47_or0[0];
  assign csa_component50_out[100] = csa_component50_fa48_or0[0];
  assign csa_component50_out[101] = csa_component50_fa49_or0[0];
endmodule

module csa_component56(input [55:0] a, input [55:0] b, input [55:0] c, output [113:0] csa_component56_out);
  wire [0:0] csa_component56_fa0_xor1;
  wire [0:0] csa_component56_fa0_or0;
  wire [0:0] csa_component56_fa1_xor1;
  wire [0:0] csa_component56_fa1_or0;
  wire [0:0] csa_component56_fa2_xor1;
  wire [0:0] csa_component56_fa2_or0;
  wire [0:0] csa_component56_fa3_xor1;
  wire [0:0] csa_component56_fa3_or0;
  wire [0:0] csa_component56_fa4_xor1;
  wire [0:0] csa_component56_fa4_or0;
  wire [0:0] csa_component56_fa5_xor1;
  wire [0:0] csa_component56_fa5_or0;
  wire [0:0] csa_component56_fa6_xor1;
  wire [0:0] csa_component56_fa6_or0;
  wire [0:0] csa_component56_fa7_xor1;
  wire [0:0] csa_component56_fa7_or0;
  wire [0:0] csa_component56_fa8_xor1;
  wire [0:0] csa_component56_fa8_or0;
  wire [0:0] csa_component56_fa9_xor1;
  wire [0:0] csa_component56_fa9_or0;
  wire [0:0] csa_component56_fa10_xor1;
  wire [0:0] csa_component56_fa10_or0;
  wire [0:0] csa_component56_fa11_xor1;
  wire [0:0] csa_component56_fa11_or0;
  wire [0:0] csa_component56_fa12_xor1;
  wire [0:0] csa_component56_fa12_or0;
  wire [0:0] csa_component56_fa13_xor1;
  wire [0:0] csa_component56_fa13_or0;
  wire [0:0] csa_component56_fa14_xor1;
  wire [0:0] csa_component56_fa14_or0;
  wire [0:0] csa_component56_fa15_xor1;
  wire [0:0] csa_component56_fa15_or0;
  wire [0:0] csa_component56_fa16_xor1;
  wire [0:0] csa_component56_fa16_or0;
  wire [0:0] csa_component56_fa17_xor1;
  wire [0:0] csa_component56_fa17_or0;
  wire [0:0] csa_component56_fa18_xor1;
  wire [0:0] csa_component56_fa18_or0;
  wire [0:0] csa_component56_fa19_xor1;
  wire [0:0] csa_component56_fa19_or0;
  wire [0:0] csa_component56_fa20_xor1;
  wire [0:0] csa_component56_fa20_or0;
  wire [0:0] csa_component56_fa21_xor1;
  wire [0:0] csa_component56_fa21_or0;
  wire [0:0] csa_component56_fa22_xor1;
  wire [0:0] csa_component56_fa22_or0;
  wire [0:0] csa_component56_fa23_xor1;
  wire [0:0] csa_component56_fa23_or0;
  wire [0:0] csa_component56_fa24_xor1;
  wire [0:0] csa_component56_fa24_or0;
  wire [0:0] csa_component56_fa25_xor1;
  wire [0:0] csa_component56_fa25_or0;
  wire [0:0] csa_component56_fa26_xor1;
  wire [0:0] csa_component56_fa26_or0;
  wire [0:0] csa_component56_fa27_xor1;
  wire [0:0] csa_component56_fa27_or0;
  wire [0:0] csa_component56_fa28_xor1;
  wire [0:0] csa_component56_fa28_or0;
  wire [0:0] csa_component56_fa29_xor1;
  wire [0:0] csa_component56_fa29_or0;
  wire [0:0] csa_component56_fa30_xor1;
  wire [0:0] csa_component56_fa30_or0;
  wire [0:0] csa_component56_fa31_xor1;
  wire [0:0] csa_component56_fa31_or0;
  wire [0:0] csa_component56_fa32_xor1;
  wire [0:0] csa_component56_fa32_or0;
  wire [0:0] csa_component56_fa33_xor1;
  wire [0:0] csa_component56_fa33_or0;
  wire [0:0] csa_component56_fa34_xor1;
  wire [0:0] csa_component56_fa34_or0;
  wire [0:0] csa_component56_fa35_xor1;
  wire [0:0] csa_component56_fa35_or0;
  wire [0:0] csa_component56_fa36_xor1;
  wire [0:0] csa_component56_fa36_or0;
  wire [0:0] csa_component56_fa37_xor1;
  wire [0:0] csa_component56_fa37_or0;
  wire [0:0] csa_component56_fa38_xor1;
  wire [0:0] csa_component56_fa38_or0;
  wire [0:0] csa_component56_fa39_xor1;
  wire [0:0] csa_component56_fa39_or0;
  wire [0:0] csa_component56_fa40_xor1;
  wire [0:0] csa_component56_fa40_or0;
  wire [0:0] csa_component56_fa41_xor1;
  wire [0:0] csa_component56_fa41_or0;
  wire [0:0] csa_component56_fa42_xor1;
  wire [0:0] csa_component56_fa42_or0;
  wire [0:0] csa_component56_fa43_xor1;
  wire [0:0] csa_component56_fa43_or0;
  wire [0:0] csa_component56_fa44_xor1;
  wire [0:0] csa_component56_fa44_or0;
  wire [0:0] csa_component56_fa45_xor1;
  wire [0:0] csa_component56_fa45_or0;
  wire [0:0] csa_component56_fa46_xor1;
  wire [0:0] csa_component56_fa46_or0;
  wire [0:0] csa_component56_fa47_xor1;
  wire [0:0] csa_component56_fa47_or0;
  wire [0:0] csa_component56_fa48_xor1;
  wire [0:0] csa_component56_fa48_or0;
  wire [0:0] csa_component56_fa49_xor1;
  wire [0:0] csa_component56_fa49_or0;
  wire [0:0] csa_component56_fa50_xor1;
  wire [0:0] csa_component56_fa50_or0;
  wire [0:0] csa_component56_fa51_xor1;
  wire [0:0] csa_component56_fa51_or0;
  wire [0:0] csa_component56_fa52_xor1;
  wire [0:0] csa_component56_fa52_or0;
  wire [0:0] csa_component56_fa53_xor1;
  wire [0:0] csa_component56_fa53_or0;
  wire [0:0] csa_component56_fa54_xor1;
  wire [0:0] csa_component56_fa54_or0;
  wire [0:0] csa_component56_fa55_xor1;
  wire [0:0] csa_component56_fa55_or0;

  fa fa_csa_component56_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component56_fa0_xor1), .fa_or0(csa_component56_fa0_or0));
  fa fa_csa_component56_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component56_fa1_xor1), .fa_or0(csa_component56_fa1_or0));
  fa fa_csa_component56_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component56_fa2_xor1), .fa_or0(csa_component56_fa2_or0));
  fa fa_csa_component56_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component56_fa3_xor1), .fa_or0(csa_component56_fa3_or0));
  fa fa_csa_component56_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component56_fa4_xor1), .fa_or0(csa_component56_fa4_or0));
  fa fa_csa_component56_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component56_fa5_xor1), .fa_or0(csa_component56_fa5_or0));
  fa fa_csa_component56_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component56_fa6_xor1), .fa_or0(csa_component56_fa6_or0));
  fa fa_csa_component56_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component56_fa7_xor1), .fa_or0(csa_component56_fa7_or0));
  fa fa_csa_component56_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component56_fa8_xor1), .fa_or0(csa_component56_fa8_or0));
  fa fa_csa_component56_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component56_fa9_xor1), .fa_or0(csa_component56_fa9_or0));
  fa fa_csa_component56_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component56_fa10_xor1), .fa_or0(csa_component56_fa10_or0));
  fa fa_csa_component56_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component56_fa11_xor1), .fa_or0(csa_component56_fa11_or0));
  fa fa_csa_component56_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component56_fa12_xor1), .fa_or0(csa_component56_fa12_or0));
  fa fa_csa_component56_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component56_fa13_xor1), .fa_or0(csa_component56_fa13_or0));
  fa fa_csa_component56_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component56_fa14_xor1), .fa_or0(csa_component56_fa14_or0));
  fa fa_csa_component56_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component56_fa15_xor1), .fa_or0(csa_component56_fa15_or0));
  fa fa_csa_component56_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component56_fa16_xor1), .fa_or0(csa_component56_fa16_or0));
  fa fa_csa_component56_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component56_fa17_xor1), .fa_or0(csa_component56_fa17_or0));
  fa fa_csa_component56_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component56_fa18_xor1), .fa_or0(csa_component56_fa18_or0));
  fa fa_csa_component56_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component56_fa19_xor1), .fa_or0(csa_component56_fa19_or0));
  fa fa_csa_component56_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component56_fa20_xor1), .fa_or0(csa_component56_fa20_or0));
  fa fa_csa_component56_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component56_fa21_xor1), .fa_or0(csa_component56_fa21_or0));
  fa fa_csa_component56_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component56_fa22_xor1), .fa_or0(csa_component56_fa22_or0));
  fa fa_csa_component56_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component56_fa23_xor1), .fa_or0(csa_component56_fa23_or0));
  fa fa_csa_component56_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component56_fa24_xor1), .fa_or0(csa_component56_fa24_or0));
  fa fa_csa_component56_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component56_fa25_xor1), .fa_or0(csa_component56_fa25_or0));
  fa fa_csa_component56_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component56_fa26_xor1), .fa_or0(csa_component56_fa26_or0));
  fa fa_csa_component56_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component56_fa27_xor1), .fa_or0(csa_component56_fa27_or0));
  fa fa_csa_component56_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component56_fa28_xor1), .fa_or0(csa_component56_fa28_or0));
  fa fa_csa_component56_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component56_fa29_xor1), .fa_or0(csa_component56_fa29_or0));
  fa fa_csa_component56_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component56_fa30_xor1), .fa_or0(csa_component56_fa30_or0));
  fa fa_csa_component56_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component56_fa31_xor1), .fa_or0(csa_component56_fa31_or0));
  fa fa_csa_component56_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component56_fa32_xor1), .fa_or0(csa_component56_fa32_or0));
  fa fa_csa_component56_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component56_fa33_xor1), .fa_or0(csa_component56_fa33_or0));
  fa fa_csa_component56_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component56_fa34_xor1), .fa_or0(csa_component56_fa34_or0));
  fa fa_csa_component56_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component56_fa35_xor1), .fa_or0(csa_component56_fa35_or0));
  fa fa_csa_component56_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component56_fa36_xor1), .fa_or0(csa_component56_fa36_or0));
  fa fa_csa_component56_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component56_fa37_xor1), .fa_or0(csa_component56_fa37_or0));
  fa fa_csa_component56_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component56_fa38_xor1), .fa_or0(csa_component56_fa38_or0));
  fa fa_csa_component56_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component56_fa39_xor1), .fa_or0(csa_component56_fa39_or0));
  fa fa_csa_component56_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component56_fa40_xor1), .fa_or0(csa_component56_fa40_or0));
  fa fa_csa_component56_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component56_fa41_xor1), .fa_or0(csa_component56_fa41_or0));
  fa fa_csa_component56_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component56_fa42_xor1), .fa_or0(csa_component56_fa42_or0));
  fa fa_csa_component56_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component56_fa43_xor1), .fa_or0(csa_component56_fa43_or0));
  fa fa_csa_component56_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component56_fa44_xor1), .fa_or0(csa_component56_fa44_or0));
  fa fa_csa_component56_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component56_fa45_xor1), .fa_or0(csa_component56_fa45_or0));
  fa fa_csa_component56_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component56_fa46_xor1), .fa_or0(csa_component56_fa46_or0));
  fa fa_csa_component56_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component56_fa47_xor1), .fa_or0(csa_component56_fa47_or0));
  fa fa_csa_component56_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component56_fa48_xor1), .fa_or0(csa_component56_fa48_or0));
  fa fa_csa_component56_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component56_fa49_xor1), .fa_or0(csa_component56_fa49_or0));
  fa fa_csa_component56_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component56_fa50_xor1), .fa_or0(csa_component56_fa50_or0));
  fa fa_csa_component56_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component56_fa51_xor1), .fa_or0(csa_component56_fa51_or0));
  fa fa_csa_component56_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component56_fa52_xor1), .fa_or0(csa_component56_fa52_or0));
  fa fa_csa_component56_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component56_fa53_xor1), .fa_or0(csa_component56_fa53_or0));
  fa fa_csa_component56_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component56_fa54_xor1), .fa_or0(csa_component56_fa54_or0));
  fa fa_csa_component56_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component56_fa55_xor1), .fa_or0(csa_component56_fa55_or0));

  assign csa_component56_out[0] = csa_component56_fa0_xor1[0];
  assign csa_component56_out[1] = csa_component56_fa1_xor1[0];
  assign csa_component56_out[2] = csa_component56_fa2_xor1[0];
  assign csa_component56_out[3] = csa_component56_fa3_xor1[0];
  assign csa_component56_out[4] = csa_component56_fa4_xor1[0];
  assign csa_component56_out[5] = csa_component56_fa5_xor1[0];
  assign csa_component56_out[6] = csa_component56_fa6_xor1[0];
  assign csa_component56_out[7] = csa_component56_fa7_xor1[0];
  assign csa_component56_out[8] = csa_component56_fa8_xor1[0];
  assign csa_component56_out[9] = csa_component56_fa9_xor1[0];
  assign csa_component56_out[10] = csa_component56_fa10_xor1[0];
  assign csa_component56_out[11] = csa_component56_fa11_xor1[0];
  assign csa_component56_out[12] = csa_component56_fa12_xor1[0];
  assign csa_component56_out[13] = csa_component56_fa13_xor1[0];
  assign csa_component56_out[14] = csa_component56_fa14_xor1[0];
  assign csa_component56_out[15] = csa_component56_fa15_xor1[0];
  assign csa_component56_out[16] = csa_component56_fa16_xor1[0];
  assign csa_component56_out[17] = csa_component56_fa17_xor1[0];
  assign csa_component56_out[18] = csa_component56_fa18_xor1[0];
  assign csa_component56_out[19] = csa_component56_fa19_xor1[0];
  assign csa_component56_out[20] = csa_component56_fa20_xor1[0];
  assign csa_component56_out[21] = csa_component56_fa21_xor1[0];
  assign csa_component56_out[22] = csa_component56_fa22_xor1[0];
  assign csa_component56_out[23] = csa_component56_fa23_xor1[0];
  assign csa_component56_out[24] = csa_component56_fa24_xor1[0];
  assign csa_component56_out[25] = csa_component56_fa25_xor1[0];
  assign csa_component56_out[26] = csa_component56_fa26_xor1[0];
  assign csa_component56_out[27] = csa_component56_fa27_xor1[0];
  assign csa_component56_out[28] = csa_component56_fa28_xor1[0];
  assign csa_component56_out[29] = csa_component56_fa29_xor1[0];
  assign csa_component56_out[30] = csa_component56_fa30_xor1[0];
  assign csa_component56_out[31] = csa_component56_fa31_xor1[0];
  assign csa_component56_out[32] = csa_component56_fa32_xor1[0];
  assign csa_component56_out[33] = csa_component56_fa33_xor1[0];
  assign csa_component56_out[34] = csa_component56_fa34_xor1[0];
  assign csa_component56_out[35] = csa_component56_fa35_xor1[0];
  assign csa_component56_out[36] = csa_component56_fa36_xor1[0];
  assign csa_component56_out[37] = csa_component56_fa37_xor1[0];
  assign csa_component56_out[38] = csa_component56_fa38_xor1[0];
  assign csa_component56_out[39] = csa_component56_fa39_xor1[0];
  assign csa_component56_out[40] = csa_component56_fa40_xor1[0];
  assign csa_component56_out[41] = csa_component56_fa41_xor1[0];
  assign csa_component56_out[42] = csa_component56_fa42_xor1[0];
  assign csa_component56_out[43] = csa_component56_fa43_xor1[0];
  assign csa_component56_out[44] = csa_component56_fa44_xor1[0];
  assign csa_component56_out[45] = csa_component56_fa45_xor1[0];
  assign csa_component56_out[46] = csa_component56_fa46_xor1[0];
  assign csa_component56_out[47] = csa_component56_fa47_xor1[0];
  assign csa_component56_out[48] = csa_component56_fa48_xor1[0];
  assign csa_component56_out[49] = csa_component56_fa49_xor1[0];
  assign csa_component56_out[50] = csa_component56_fa50_xor1[0];
  assign csa_component56_out[51] = csa_component56_fa51_xor1[0];
  assign csa_component56_out[52] = csa_component56_fa52_xor1[0];
  assign csa_component56_out[53] = csa_component56_fa53_xor1[0];
  assign csa_component56_out[54] = csa_component56_fa54_xor1[0];
  assign csa_component56_out[55] = csa_component56_fa55_xor1[0];
  assign csa_component56_out[56] = 1'b0;
  assign csa_component56_out[57] = 1'b0;
  assign csa_component56_out[58] = csa_component56_fa0_or0[0];
  assign csa_component56_out[59] = csa_component56_fa1_or0[0];
  assign csa_component56_out[60] = csa_component56_fa2_or0[0];
  assign csa_component56_out[61] = csa_component56_fa3_or0[0];
  assign csa_component56_out[62] = csa_component56_fa4_or0[0];
  assign csa_component56_out[63] = csa_component56_fa5_or0[0];
  assign csa_component56_out[64] = csa_component56_fa6_or0[0];
  assign csa_component56_out[65] = csa_component56_fa7_or0[0];
  assign csa_component56_out[66] = csa_component56_fa8_or0[0];
  assign csa_component56_out[67] = csa_component56_fa9_or0[0];
  assign csa_component56_out[68] = csa_component56_fa10_or0[0];
  assign csa_component56_out[69] = csa_component56_fa11_or0[0];
  assign csa_component56_out[70] = csa_component56_fa12_or0[0];
  assign csa_component56_out[71] = csa_component56_fa13_or0[0];
  assign csa_component56_out[72] = csa_component56_fa14_or0[0];
  assign csa_component56_out[73] = csa_component56_fa15_or0[0];
  assign csa_component56_out[74] = csa_component56_fa16_or0[0];
  assign csa_component56_out[75] = csa_component56_fa17_or0[0];
  assign csa_component56_out[76] = csa_component56_fa18_or0[0];
  assign csa_component56_out[77] = csa_component56_fa19_or0[0];
  assign csa_component56_out[78] = csa_component56_fa20_or0[0];
  assign csa_component56_out[79] = csa_component56_fa21_or0[0];
  assign csa_component56_out[80] = csa_component56_fa22_or0[0];
  assign csa_component56_out[81] = csa_component56_fa23_or0[0];
  assign csa_component56_out[82] = csa_component56_fa24_or0[0];
  assign csa_component56_out[83] = csa_component56_fa25_or0[0];
  assign csa_component56_out[84] = csa_component56_fa26_or0[0];
  assign csa_component56_out[85] = csa_component56_fa27_or0[0];
  assign csa_component56_out[86] = csa_component56_fa28_or0[0];
  assign csa_component56_out[87] = csa_component56_fa29_or0[0];
  assign csa_component56_out[88] = csa_component56_fa30_or0[0];
  assign csa_component56_out[89] = csa_component56_fa31_or0[0];
  assign csa_component56_out[90] = csa_component56_fa32_or0[0];
  assign csa_component56_out[91] = csa_component56_fa33_or0[0];
  assign csa_component56_out[92] = csa_component56_fa34_or0[0];
  assign csa_component56_out[93] = csa_component56_fa35_or0[0];
  assign csa_component56_out[94] = csa_component56_fa36_or0[0];
  assign csa_component56_out[95] = csa_component56_fa37_or0[0];
  assign csa_component56_out[96] = csa_component56_fa38_or0[0];
  assign csa_component56_out[97] = csa_component56_fa39_or0[0];
  assign csa_component56_out[98] = csa_component56_fa40_or0[0];
  assign csa_component56_out[99] = csa_component56_fa41_or0[0];
  assign csa_component56_out[100] = csa_component56_fa42_or0[0];
  assign csa_component56_out[101] = csa_component56_fa43_or0[0];
  assign csa_component56_out[102] = csa_component56_fa44_or0[0];
  assign csa_component56_out[103] = csa_component56_fa45_or0[0];
  assign csa_component56_out[104] = csa_component56_fa46_or0[0];
  assign csa_component56_out[105] = csa_component56_fa47_or0[0];
  assign csa_component56_out[106] = csa_component56_fa48_or0[0];
  assign csa_component56_out[107] = csa_component56_fa49_or0[0];
  assign csa_component56_out[108] = csa_component56_fa50_or0[0];
  assign csa_component56_out[109] = csa_component56_fa51_or0[0];
  assign csa_component56_out[110] = csa_component56_fa52_or0[0];
  assign csa_component56_out[111] = csa_component56_fa53_or0[0];
  assign csa_component56_out[112] = csa_component56_fa54_or0[0];
  assign csa_component56_out[113] = csa_component56_fa55_or0[0];
endmodule

module csa_component59(input [58:0] a, input [58:0] b, input [58:0] c, output [119:0] csa_component59_out);
  wire [0:0] csa_component59_fa0_xor1;
  wire [0:0] csa_component59_fa0_or0;
  wire [0:0] csa_component59_fa1_xor1;
  wire [0:0] csa_component59_fa1_or0;
  wire [0:0] csa_component59_fa2_xor1;
  wire [0:0] csa_component59_fa2_or0;
  wire [0:0] csa_component59_fa3_xor1;
  wire [0:0] csa_component59_fa3_or0;
  wire [0:0] csa_component59_fa4_xor1;
  wire [0:0] csa_component59_fa4_or0;
  wire [0:0] csa_component59_fa5_xor1;
  wire [0:0] csa_component59_fa5_or0;
  wire [0:0] csa_component59_fa6_xor1;
  wire [0:0] csa_component59_fa6_or0;
  wire [0:0] csa_component59_fa7_xor1;
  wire [0:0] csa_component59_fa7_or0;
  wire [0:0] csa_component59_fa8_xor1;
  wire [0:0] csa_component59_fa8_or0;
  wire [0:0] csa_component59_fa9_xor1;
  wire [0:0] csa_component59_fa9_or0;
  wire [0:0] csa_component59_fa10_xor1;
  wire [0:0] csa_component59_fa10_or0;
  wire [0:0] csa_component59_fa11_xor1;
  wire [0:0] csa_component59_fa11_or0;
  wire [0:0] csa_component59_fa12_xor1;
  wire [0:0] csa_component59_fa12_or0;
  wire [0:0] csa_component59_fa13_xor1;
  wire [0:0] csa_component59_fa13_or0;
  wire [0:0] csa_component59_fa14_xor1;
  wire [0:0] csa_component59_fa14_or0;
  wire [0:0] csa_component59_fa15_xor1;
  wire [0:0] csa_component59_fa15_or0;
  wire [0:0] csa_component59_fa16_xor1;
  wire [0:0] csa_component59_fa16_or0;
  wire [0:0] csa_component59_fa17_xor1;
  wire [0:0] csa_component59_fa17_or0;
  wire [0:0] csa_component59_fa18_xor1;
  wire [0:0] csa_component59_fa18_or0;
  wire [0:0] csa_component59_fa19_xor1;
  wire [0:0] csa_component59_fa19_or0;
  wire [0:0] csa_component59_fa20_xor1;
  wire [0:0] csa_component59_fa20_or0;
  wire [0:0] csa_component59_fa21_xor1;
  wire [0:0] csa_component59_fa21_or0;
  wire [0:0] csa_component59_fa22_xor1;
  wire [0:0] csa_component59_fa22_or0;
  wire [0:0] csa_component59_fa23_xor1;
  wire [0:0] csa_component59_fa23_or0;
  wire [0:0] csa_component59_fa24_xor1;
  wire [0:0] csa_component59_fa24_or0;
  wire [0:0] csa_component59_fa25_xor1;
  wire [0:0] csa_component59_fa25_or0;
  wire [0:0] csa_component59_fa26_xor1;
  wire [0:0] csa_component59_fa26_or0;
  wire [0:0] csa_component59_fa27_xor1;
  wire [0:0] csa_component59_fa27_or0;
  wire [0:0] csa_component59_fa28_xor1;
  wire [0:0] csa_component59_fa28_or0;
  wire [0:0] csa_component59_fa29_xor1;
  wire [0:0] csa_component59_fa29_or0;
  wire [0:0] csa_component59_fa30_xor1;
  wire [0:0] csa_component59_fa30_or0;
  wire [0:0] csa_component59_fa31_xor1;
  wire [0:0] csa_component59_fa31_or0;
  wire [0:0] csa_component59_fa32_xor1;
  wire [0:0] csa_component59_fa32_or0;
  wire [0:0] csa_component59_fa33_xor1;
  wire [0:0] csa_component59_fa33_or0;
  wire [0:0] csa_component59_fa34_xor1;
  wire [0:0] csa_component59_fa34_or0;
  wire [0:0] csa_component59_fa35_xor1;
  wire [0:0] csa_component59_fa35_or0;
  wire [0:0] csa_component59_fa36_xor1;
  wire [0:0] csa_component59_fa36_or0;
  wire [0:0] csa_component59_fa37_xor1;
  wire [0:0] csa_component59_fa37_or0;
  wire [0:0] csa_component59_fa38_xor1;
  wire [0:0] csa_component59_fa38_or0;
  wire [0:0] csa_component59_fa39_xor1;
  wire [0:0] csa_component59_fa39_or0;
  wire [0:0] csa_component59_fa40_xor1;
  wire [0:0] csa_component59_fa40_or0;
  wire [0:0] csa_component59_fa41_xor1;
  wire [0:0] csa_component59_fa41_or0;
  wire [0:0] csa_component59_fa42_xor1;
  wire [0:0] csa_component59_fa42_or0;
  wire [0:0] csa_component59_fa43_xor1;
  wire [0:0] csa_component59_fa43_or0;
  wire [0:0] csa_component59_fa44_xor1;
  wire [0:0] csa_component59_fa44_or0;
  wire [0:0] csa_component59_fa45_xor1;
  wire [0:0] csa_component59_fa45_or0;
  wire [0:0] csa_component59_fa46_xor1;
  wire [0:0] csa_component59_fa46_or0;
  wire [0:0] csa_component59_fa47_xor1;
  wire [0:0] csa_component59_fa47_or0;
  wire [0:0] csa_component59_fa48_xor1;
  wire [0:0] csa_component59_fa48_or0;
  wire [0:0] csa_component59_fa49_xor1;
  wire [0:0] csa_component59_fa49_or0;
  wire [0:0] csa_component59_fa50_xor1;
  wire [0:0] csa_component59_fa50_or0;
  wire [0:0] csa_component59_fa51_xor1;
  wire [0:0] csa_component59_fa51_or0;
  wire [0:0] csa_component59_fa52_xor1;
  wire [0:0] csa_component59_fa52_or0;
  wire [0:0] csa_component59_fa53_xor1;
  wire [0:0] csa_component59_fa53_or0;
  wire [0:0] csa_component59_fa54_xor1;
  wire [0:0] csa_component59_fa54_or0;
  wire [0:0] csa_component59_fa55_xor1;
  wire [0:0] csa_component59_fa55_or0;
  wire [0:0] csa_component59_fa56_xor1;
  wire [0:0] csa_component59_fa56_or0;
  wire [0:0] csa_component59_fa57_xor1;
  wire [0:0] csa_component59_fa57_or0;
  wire [0:0] csa_component59_fa58_xor1;
  wire [0:0] csa_component59_fa58_or0;

  fa fa_csa_component59_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component59_fa0_xor1), .fa_or0(csa_component59_fa0_or0));
  fa fa_csa_component59_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component59_fa1_xor1), .fa_or0(csa_component59_fa1_or0));
  fa fa_csa_component59_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component59_fa2_xor1), .fa_or0(csa_component59_fa2_or0));
  fa fa_csa_component59_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component59_fa3_xor1), .fa_or0(csa_component59_fa3_or0));
  fa fa_csa_component59_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component59_fa4_xor1), .fa_or0(csa_component59_fa4_or0));
  fa fa_csa_component59_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component59_fa5_xor1), .fa_or0(csa_component59_fa5_or0));
  fa fa_csa_component59_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component59_fa6_xor1), .fa_or0(csa_component59_fa6_or0));
  fa fa_csa_component59_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component59_fa7_xor1), .fa_or0(csa_component59_fa7_or0));
  fa fa_csa_component59_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component59_fa8_xor1), .fa_or0(csa_component59_fa8_or0));
  fa fa_csa_component59_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component59_fa9_xor1), .fa_or0(csa_component59_fa9_or0));
  fa fa_csa_component59_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component59_fa10_xor1), .fa_or0(csa_component59_fa10_or0));
  fa fa_csa_component59_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component59_fa11_xor1), .fa_or0(csa_component59_fa11_or0));
  fa fa_csa_component59_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component59_fa12_xor1), .fa_or0(csa_component59_fa12_or0));
  fa fa_csa_component59_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component59_fa13_xor1), .fa_or0(csa_component59_fa13_or0));
  fa fa_csa_component59_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component59_fa14_xor1), .fa_or0(csa_component59_fa14_or0));
  fa fa_csa_component59_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component59_fa15_xor1), .fa_or0(csa_component59_fa15_or0));
  fa fa_csa_component59_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component59_fa16_xor1), .fa_or0(csa_component59_fa16_or0));
  fa fa_csa_component59_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component59_fa17_xor1), .fa_or0(csa_component59_fa17_or0));
  fa fa_csa_component59_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component59_fa18_xor1), .fa_or0(csa_component59_fa18_or0));
  fa fa_csa_component59_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component59_fa19_xor1), .fa_or0(csa_component59_fa19_or0));
  fa fa_csa_component59_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component59_fa20_xor1), .fa_or0(csa_component59_fa20_or0));
  fa fa_csa_component59_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component59_fa21_xor1), .fa_or0(csa_component59_fa21_or0));
  fa fa_csa_component59_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component59_fa22_xor1), .fa_or0(csa_component59_fa22_or0));
  fa fa_csa_component59_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component59_fa23_xor1), .fa_or0(csa_component59_fa23_or0));
  fa fa_csa_component59_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component59_fa24_xor1), .fa_or0(csa_component59_fa24_or0));
  fa fa_csa_component59_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component59_fa25_xor1), .fa_or0(csa_component59_fa25_or0));
  fa fa_csa_component59_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component59_fa26_xor1), .fa_or0(csa_component59_fa26_or0));
  fa fa_csa_component59_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component59_fa27_xor1), .fa_or0(csa_component59_fa27_or0));
  fa fa_csa_component59_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component59_fa28_xor1), .fa_or0(csa_component59_fa28_or0));
  fa fa_csa_component59_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component59_fa29_xor1), .fa_or0(csa_component59_fa29_or0));
  fa fa_csa_component59_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component59_fa30_xor1), .fa_or0(csa_component59_fa30_or0));
  fa fa_csa_component59_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component59_fa31_xor1), .fa_or0(csa_component59_fa31_or0));
  fa fa_csa_component59_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component59_fa32_xor1), .fa_or0(csa_component59_fa32_or0));
  fa fa_csa_component59_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component59_fa33_xor1), .fa_or0(csa_component59_fa33_or0));
  fa fa_csa_component59_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component59_fa34_xor1), .fa_or0(csa_component59_fa34_or0));
  fa fa_csa_component59_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component59_fa35_xor1), .fa_or0(csa_component59_fa35_or0));
  fa fa_csa_component59_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component59_fa36_xor1), .fa_or0(csa_component59_fa36_or0));
  fa fa_csa_component59_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component59_fa37_xor1), .fa_or0(csa_component59_fa37_or0));
  fa fa_csa_component59_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component59_fa38_xor1), .fa_or0(csa_component59_fa38_or0));
  fa fa_csa_component59_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component59_fa39_xor1), .fa_or0(csa_component59_fa39_or0));
  fa fa_csa_component59_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component59_fa40_xor1), .fa_or0(csa_component59_fa40_or0));
  fa fa_csa_component59_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component59_fa41_xor1), .fa_or0(csa_component59_fa41_or0));
  fa fa_csa_component59_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component59_fa42_xor1), .fa_or0(csa_component59_fa42_or0));
  fa fa_csa_component59_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component59_fa43_xor1), .fa_or0(csa_component59_fa43_or0));
  fa fa_csa_component59_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component59_fa44_xor1), .fa_or0(csa_component59_fa44_or0));
  fa fa_csa_component59_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component59_fa45_xor1), .fa_or0(csa_component59_fa45_or0));
  fa fa_csa_component59_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component59_fa46_xor1), .fa_or0(csa_component59_fa46_or0));
  fa fa_csa_component59_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component59_fa47_xor1), .fa_or0(csa_component59_fa47_or0));
  fa fa_csa_component59_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component59_fa48_xor1), .fa_or0(csa_component59_fa48_or0));
  fa fa_csa_component59_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component59_fa49_xor1), .fa_or0(csa_component59_fa49_or0));
  fa fa_csa_component59_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component59_fa50_xor1), .fa_or0(csa_component59_fa50_or0));
  fa fa_csa_component59_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component59_fa51_xor1), .fa_or0(csa_component59_fa51_or0));
  fa fa_csa_component59_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component59_fa52_xor1), .fa_or0(csa_component59_fa52_or0));
  fa fa_csa_component59_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component59_fa53_xor1), .fa_or0(csa_component59_fa53_or0));
  fa fa_csa_component59_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component59_fa54_xor1), .fa_or0(csa_component59_fa54_or0));
  fa fa_csa_component59_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component59_fa55_xor1), .fa_or0(csa_component59_fa55_or0));
  fa fa_csa_component59_fa56_out(.a(a[56]), .b(b[56]), .cin(c[56]), .fa_xor1(csa_component59_fa56_xor1), .fa_or0(csa_component59_fa56_or0));
  fa fa_csa_component59_fa57_out(.a(a[57]), .b(b[57]), .cin(c[57]), .fa_xor1(csa_component59_fa57_xor1), .fa_or0(csa_component59_fa57_or0));
  fa fa_csa_component59_fa58_out(.a(a[58]), .b(b[58]), .cin(c[58]), .fa_xor1(csa_component59_fa58_xor1), .fa_or0(csa_component59_fa58_or0));

  assign csa_component59_out[0] = csa_component59_fa0_xor1[0];
  assign csa_component59_out[1] = csa_component59_fa1_xor1[0];
  assign csa_component59_out[2] = csa_component59_fa2_xor1[0];
  assign csa_component59_out[3] = csa_component59_fa3_xor1[0];
  assign csa_component59_out[4] = csa_component59_fa4_xor1[0];
  assign csa_component59_out[5] = csa_component59_fa5_xor1[0];
  assign csa_component59_out[6] = csa_component59_fa6_xor1[0];
  assign csa_component59_out[7] = csa_component59_fa7_xor1[0];
  assign csa_component59_out[8] = csa_component59_fa8_xor1[0];
  assign csa_component59_out[9] = csa_component59_fa9_xor1[0];
  assign csa_component59_out[10] = csa_component59_fa10_xor1[0];
  assign csa_component59_out[11] = csa_component59_fa11_xor1[0];
  assign csa_component59_out[12] = csa_component59_fa12_xor1[0];
  assign csa_component59_out[13] = csa_component59_fa13_xor1[0];
  assign csa_component59_out[14] = csa_component59_fa14_xor1[0];
  assign csa_component59_out[15] = csa_component59_fa15_xor1[0];
  assign csa_component59_out[16] = csa_component59_fa16_xor1[0];
  assign csa_component59_out[17] = csa_component59_fa17_xor1[0];
  assign csa_component59_out[18] = csa_component59_fa18_xor1[0];
  assign csa_component59_out[19] = csa_component59_fa19_xor1[0];
  assign csa_component59_out[20] = csa_component59_fa20_xor1[0];
  assign csa_component59_out[21] = csa_component59_fa21_xor1[0];
  assign csa_component59_out[22] = csa_component59_fa22_xor1[0];
  assign csa_component59_out[23] = csa_component59_fa23_xor1[0];
  assign csa_component59_out[24] = csa_component59_fa24_xor1[0];
  assign csa_component59_out[25] = csa_component59_fa25_xor1[0];
  assign csa_component59_out[26] = csa_component59_fa26_xor1[0];
  assign csa_component59_out[27] = csa_component59_fa27_xor1[0];
  assign csa_component59_out[28] = csa_component59_fa28_xor1[0];
  assign csa_component59_out[29] = csa_component59_fa29_xor1[0];
  assign csa_component59_out[30] = csa_component59_fa30_xor1[0];
  assign csa_component59_out[31] = csa_component59_fa31_xor1[0];
  assign csa_component59_out[32] = csa_component59_fa32_xor1[0];
  assign csa_component59_out[33] = csa_component59_fa33_xor1[0];
  assign csa_component59_out[34] = csa_component59_fa34_xor1[0];
  assign csa_component59_out[35] = csa_component59_fa35_xor1[0];
  assign csa_component59_out[36] = csa_component59_fa36_xor1[0];
  assign csa_component59_out[37] = csa_component59_fa37_xor1[0];
  assign csa_component59_out[38] = csa_component59_fa38_xor1[0];
  assign csa_component59_out[39] = csa_component59_fa39_xor1[0];
  assign csa_component59_out[40] = csa_component59_fa40_xor1[0];
  assign csa_component59_out[41] = csa_component59_fa41_xor1[0];
  assign csa_component59_out[42] = csa_component59_fa42_xor1[0];
  assign csa_component59_out[43] = csa_component59_fa43_xor1[0];
  assign csa_component59_out[44] = csa_component59_fa44_xor1[0];
  assign csa_component59_out[45] = csa_component59_fa45_xor1[0];
  assign csa_component59_out[46] = csa_component59_fa46_xor1[0];
  assign csa_component59_out[47] = csa_component59_fa47_xor1[0];
  assign csa_component59_out[48] = csa_component59_fa48_xor1[0];
  assign csa_component59_out[49] = csa_component59_fa49_xor1[0];
  assign csa_component59_out[50] = csa_component59_fa50_xor1[0];
  assign csa_component59_out[51] = csa_component59_fa51_xor1[0];
  assign csa_component59_out[52] = csa_component59_fa52_xor1[0];
  assign csa_component59_out[53] = csa_component59_fa53_xor1[0];
  assign csa_component59_out[54] = csa_component59_fa54_xor1[0];
  assign csa_component59_out[55] = csa_component59_fa55_xor1[0];
  assign csa_component59_out[56] = csa_component59_fa56_xor1[0];
  assign csa_component59_out[57] = csa_component59_fa57_xor1[0];
  assign csa_component59_out[58] = csa_component59_fa58_xor1[0];
  assign csa_component59_out[59] = 1'b0;
  assign csa_component59_out[60] = 1'b0;
  assign csa_component59_out[61] = csa_component59_fa0_or0[0];
  assign csa_component59_out[62] = csa_component59_fa1_or0[0];
  assign csa_component59_out[63] = csa_component59_fa2_or0[0];
  assign csa_component59_out[64] = csa_component59_fa3_or0[0];
  assign csa_component59_out[65] = csa_component59_fa4_or0[0];
  assign csa_component59_out[66] = csa_component59_fa5_or0[0];
  assign csa_component59_out[67] = csa_component59_fa6_or0[0];
  assign csa_component59_out[68] = csa_component59_fa7_or0[0];
  assign csa_component59_out[69] = csa_component59_fa8_or0[0];
  assign csa_component59_out[70] = csa_component59_fa9_or0[0];
  assign csa_component59_out[71] = csa_component59_fa10_or0[0];
  assign csa_component59_out[72] = csa_component59_fa11_or0[0];
  assign csa_component59_out[73] = csa_component59_fa12_or0[0];
  assign csa_component59_out[74] = csa_component59_fa13_or0[0];
  assign csa_component59_out[75] = csa_component59_fa14_or0[0];
  assign csa_component59_out[76] = csa_component59_fa15_or0[0];
  assign csa_component59_out[77] = csa_component59_fa16_or0[0];
  assign csa_component59_out[78] = csa_component59_fa17_or0[0];
  assign csa_component59_out[79] = csa_component59_fa18_or0[0];
  assign csa_component59_out[80] = csa_component59_fa19_or0[0];
  assign csa_component59_out[81] = csa_component59_fa20_or0[0];
  assign csa_component59_out[82] = csa_component59_fa21_or0[0];
  assign csa_component59_out[83] = csa_component59_fa22_or0[0];
  assign csa_component59_out[84] = csa_component59_fa23_or0[0];
  assign csa_component59_out[85] = csa_component59_fa24_or0[0];
  assign csa_component59_out[86] = csa_component59_fa25_or0[0];
  assign csa_component59_out[87] = csa_component59_fa26_or0[0];
  assign csa_component59_out[88] = csa_component59_fa27_or0[0];
  assign csa_component59_out[89] = csa_component59_fa28_or0[0];
  assign csa_component59_out[90] = csa_component59_fa29_or0[0];
  assign csa_component59_out[91] = csa_component59_fa30_or0[0];
  assign csa_component59_out[92] = csa_component59_fa31_or0[0];
  assign csa_component59_out[93] = csa_component59_fa32_or0[0];
  assign csa_component59_out[94] = csa_component59_fa33_or0[0];
  assign csa_component59_out[95] = csa_component59_fa34_or0[0];
  assign csa_component59_out[96] = csa_component59_fa35_or0[0];
  assign csa_component59_out[97] = csa_component59_fa36_or0[0];
  assign csa_component59_out[98] = csa_component59_fa37_or0[0];
  assign csa_component59_out[99] = csa_component59_fa38_or0[0];
  assign csa_component59_out[100] = csa_component59_fa39_or0[0];
  assign csa_component59_out[101] = csa_component59_fa40_or0[0];
  assign csa_component59_out[102] = csa_component59_fa41_or0[0];
  assign csa_component59_out[103] = csa_component59_fa42_or0[0];
  assign csa_component59_out[104] = csa_component59_fa43_or0[0];
  assign csa_component59_out[105] = csa_component59_fa44_or0[0];
  assign csa_component59_out[106] = csa_component59_fa45_or0[0];
  assign csa_component59_out[107] = csa_component59_fa46_or0[0];
  assign csa_component59_out[108] = csa_component59_fa47_or0[0];
  assign csa_component59_out[109] = csa_component59_fa48_or0[0];
  assign csa_component59_out[110] = csa_component59_fa49_or0[0];
  assign csa_component59_out[111] = csa_component59_fa50_or0[0];
  assign csa_component59_out[112] = csa_component59_fa51_or0[0];
  assign csa_component59_out[113] = csa_component59_fa52_or0[0];
  assign csa_component59_out[114] = csa_component59_fa53_or0[0];
  assign csa_component59_out[115] = csa_component59_fa54_or0[0];
  assign csa_component59_out[116] = csa_component59_fa55_or0[0];
  assign csa_component59_out[117] = csa_component59_fa56_or0[0];
  assign csa_component59_out[118] = csa_component59_fa57_or0[0];
  assign csa_component59_out[119] = csa_component59_fa58_or0[0];
endmodule

module csa_component62(input [61:0] a, input [61:0] b, input [61:0] c, output [125:0] csa_component62_out);
  wire [0:0] csa_component62_fa0_xor1;
  wire [0:0] csa_component62_fa0_or0;
  wire [0:0] csa_component62_fa1_xor1;
  wire [0:0] csa_component62_fa1_or0;
  wire [0:0] csa_component62_fa2_xor1;
  wire [0:0] csa_component62_fa2_or0;
  wire [0:0] csa_component62_fa3_xor1;
  wire [0:0] csa_component62_fa3_or0;
  wire [0:0] csa_component62_fa4_xor1;
  wire [0:0] csa_component62_fa4_or0;
  wire [0:0] csa_component62_fa5_xor1;
  wire [0:0] csa_component62_fa5_or0;
  wire [0:0] csa_component62_fa6_xor1;
  wire [0:0] csa_component62_fa6_or0;
  wire [0:0] csa_component62_fa7_xor1;
  wire [0:0] csa_component62_fa7_or0;
  wire [0:0] csa_component62_fa8_xor1;
  wire [0:0] csa_component62_fa8_or0;
  wire [0:0] csa_component62_fa9_xor1;
  wire [0:0] csa_component62_fa9_or0;
  wire [0:0] csa_component62_fa10_xor1;
  wire [0:0] csa_component62_fa10_or0;
  wire [0:0] csa_component62_fa11_xor1;
  wire [0:0] csa_component62_fa11_or0;
  wire [0:0] csa_component62_fa12_xor1;
  wire [0:0] csa_component62_fa12_or0;
  wire [0:0] csa_component62_fa13_xor1;
  wire [0:0] csa_component62_fa13_or0;
  wire [0:0] csa_component62_fa14_xor1;
  wire [0:0] csa_component62_fa14_or0;
  wire [0:0] csa_component62_fa15_xor1;
  wire [0:0] csa_component62_fa15_or0;
  wire [0:0] csa_component62_fa16_xor1;
  wire [0:0] csa_component62_fa16_or0;
  wire [0:0] csa_component62_fa17_xor1;
  wire [0:0] csa_component62_fa17_or0;
  wire [0:0] csa_component62_fa18_xor1;
  wire [0:0] csa_component62_fa18_or0;
  wire [0:0] csa_component62_fa19_xor1;
  wire [0:0] csa_component62_fa19_or0;
  wire [0:0] csa_component62_fa20_xor1;
  wire [0:0] csa_component62_fa20_or0;
  wire [0:0] csa_component62_fa21_xor1;
  wire [0:0] csa_component62_fa21_or0;
  wire [0:0] csa_component62_fa22_xor1;
  wire [0:0] csa_component62_fa22_or0;
  wire [0:0] csa_component62_fa23_xor1;
  wire [0:0] csa_component62_fa23_or0;
  wire [0:0] csa_component62_fa24_xor1;
  wire [0:0] csa_component62_fa24_or0;
  wire [0:0] csa_component62_fa25_xor1;
  wire [0:0] csa_component62_fa25_or0;
  wire [0:0] csa_component62_fa26_xor1;
  wire [0:0] csa_component62_fa26_or0;
  wire [0:0] csa_component62_fa27_xor1;
  wire [0:0] csa_component62_fa27_or0;
  wire [0:0] csa_component62_fa28_xor1;
  wire [0:0] csa_component62_fa28_or0;
  wire [0:0] csa_component62_fa29_xor1;
  wire [0:0] csa_component62_fa29_or0;
  wire [0:0] csa_component62_fa30_xor1;
  wire [0:0] csa_component62_fa30_or0;
  wire [0:0] csa_component62_fa31_xor1;
  wire [0:0] csa_component62_fa31_or0;
  wire [0:0] csa_component62_fa32_xor1;
  wire [0:0] csa_component62_fa32_or0;
  wire [0:0] csa_component62_fa33_xor1;
  wire [0:0] csa_component62_fa33_or0;
  wire [0:0] csa_component62_fa34_xor1;
  wire [0:0] csa_component62_fa34_or0;
  wire [0:0] csa_component62_fa35_xor1;
  wire [0:0] csa_component62_fa35_or0;
  wire [0:0] csa_component62_fa36_xor1;
  wire [0:0] csa_component62_fa36_or0;
  wire [0:0] csa_component62_fa37_xor1;
  wire [0:0] csa_component62_fa37_or0;
  wire [0:0] csa_component62_fa38_xor1;
  wire [0:0] csa_component62_fa38_or0;
  wire [0:0] csa_component62_fa39_xor1;
  wire [0:0] csa_component62_fa39_or0;
  wire [0:0] csa_component62_fa40_xor1;
  wire [0:0] csa_component62_fa40_or0;
  wire [0:0] csa_component62_fa41_xor1;
  wire [0:0] csa_component62_fa41_or0;
  wire [0:0] csa_component62_fa42_xor1;
  wire [0:0] csa_component62_fa42_or0;
  wire [0:0] csa_component62_fa43_xor1;
  wire [0:0] csa_component62_fa43_or0;
  wire [0:0] csa_component62_fa44_xor1;
  wire [0:0] csa_component62_fa44_or0;
  wire [0:0] csa_component62_fa45_xor1;
  wire [0:0] csa_component62_fa45_or0;
  wire [0:0] csa_component62_fa46_xor1;
  wire [0:0] csa_component62_fa46_or0;
  wire [0:0] csa_component62_fa47_xor1;
  wire [0:0] csa_component62_fa47_or0;
  wire [0:0] csa_component62_fa48_xor1;
  wire [0:0] csa_component62_fa48_or0;
  wire [0:0] csa_component62_fa49_xor1;
  wire [0:0] csa_component62_fa49_or0;
  wire [0:0] csa_component62_fa50_xor1;
  wire [0:0] csa_component62_fa50_or0;
  wire [0:0] csa_component62_fa51_xor1;
  wire [0:0] csa_component62_fa51_or0;
  wire [0:0] csa_component62_fa52_xor1;
  wire [0:0] csa_component62_fa52_or0;
  wire [0:0] csa_component62_fa53_xor1;
  wire [0:0] csa_component62_fa53_or0;
  wire [0:0] csa_component62_fa54_xor1;
  wire [0:0] csa_component62_fa54_or0;
  wire [0:0] csa_component62_fa55_xor1;
  wire [0:0] csa_component62_fa55_or0;
  wire [0:0] csa_component62_fa56_xor1;
  wire [0:0] csa_component62_fa56_or0;
  wire [0:0] csa_component62_fa57_xor1;
  wire [0:0] csa_component62_fa57_or0;
  wire [0:0] csa_component62_fa58_xor1;
  wire [0:0] csa_component62_fa58_or0;
  wire [0:0] csa_component62_fa59_xor1;
  wire [0:0] csa_component62_fa59_or0;
  wire [0:0] csa_component62_fa60_xor1;
  wire [0:0] csa_component62_fa60_or0;
  wire [0:0] csa_component62_fa61_xor1;
  wire [0:0] csa_component62_fa61_or0;

  fa fa_csa_component62_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component62_fa0_xor1), .fa_or0(csa_component62_fa0_or0));
  fa fa_csa_component62_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component62_fa1_xor1), .fa_or0(csa_component62_fa1_or0));
  fa fa_csa_component62_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component62_fa2_xor1), .fa_or0(csa_component62_fa2_or0));
  fa fa_csa_component62_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component62_fa3_xor1), .fa_or0(csa_component62_fa3_or0));
  fa fa_csa_component62_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component62_fa4_xor1), .fa_or0(csa_component62_fa4_or0));
  fa fa_csa_component62_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component62_fa5_xor1), .fa_or0(csa_component62_fa5_or0));
  fa fa_csa_component62_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component62_fa6_xor1), .fa_or0(csa_component62_fa6_or0));
  fa fa_csa_component62_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component62_fa7_xor1), .fa_or0(csa_component62_fa7_or0));
  fa fa_csa_component62_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component62_fa8_xor1), .fa_or0(csa_component62_fa8_or0));
  fa fa_csa_component62_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component62_fa9_xor1), .fa_or0(csa_component62_fa9_or0));
  fa fa_csa_component62_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component62_fa10_xor1), .fa_or0(csa_component62_fa10_or0));
  fa fa_csa_component62_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component62_fa11_xor1), .fa_or0(csa_component62_fa11_or0));
  fa fa_csa_component62_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component62_fa12_xor1), .fa_or0(csa_component62_fa12_or0));
  fa fa_csa_component62_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component62_fa13_xor1), .fa_or0(csa_component62_fa13_or0));
  fa fa_csa_component62_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component62_fa14_xor1), .fa_or0(csa_component62_fa14_or0));
  fa fa_csa_component62_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component62_fa15_xor1), .fa_or0(csa_component62_fa15_or0));
  fa fa_csa_component62_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component62_fa16_xor1), .fa_or0(csa_component62_fa16_or0));
  fa fa_csa_component62_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component62_fa17_xor1), .fa_or0(csa_component62_fa17_or0));
  fa fa_csa_component62_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component62_fa18_xor1), .fa_or0(csa_component62_fa18_or0));
  fa fa_csa_component62_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component62_fa19_xor1), .fa_or0(csa_component62_fa19_or0));
  fa fa_csa_component62_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component62_fa20_xor1), .fa_or0(csa_component62_fa20_or0));
  fa fa_csa_component62_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component62_fa21_xor1), .fa_or0(csa_component62_fa21_or0));
  fa fa_csa_component62_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component62_fa22_xor1), .fa_or0(csa_component62_fa22_or0));
  fa fa_csa_component62_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component62_fa23_xor1), .fa_or0(csa_component62_fa23_or0));
  fa fa_csa_component62_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component62_fa24_xor1), .fa_or0(csa_component62_fa24_or0));
  fa fa_csa_component62_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component62_fa25_xor1), .fa_or0(csa_component62_fa25_or0));
  fa fa_csa_component62_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component62_fa26_xor1), .fa_or0(csa_component62_fa26_or0));
  fa fa_csa_component62_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component62_fa27_xor1), .fa_or0(csa_component62_fa27_or0));
  fa fa_csa_component62_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component62_fa28_xor1), .fa_or0(csa_component62_fa28_or0));
  fa fa_csa_component62_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component62_fa29_xor1), .fa_or0(csa_component62_fa29_or0));
  fa fa_csa_component62_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component62_fa30_xor1), .fa_or0(csa_component62_fa30_or0));
  fa fa_csa_component62_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component62_fa31_xor1), .fa_or0(csa_component62_fa31_or0));
  fa fa_csa_component62_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component62_fa32_xor1), .fa_or0(csa_component62_fa32_or0));
  fa fa_csa_component62_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component62_fa33_xor1), .fa_or0(csa_component62_fa33_or0));
  fa fa_csa_component62_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component62_fa34_xor1), .fa_or0(csa_component62_fa34_or0));
  fa fa_csa_component62_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component62_fa35_xor1), .fa_or0(csa_component62_fa35_or0));
  fa fa_csa_component62_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component62_fa36_xor1), .fa_or0(csa_component62_fa36_or0));
  fa fa_csa_component62_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component62_fa37_xor1), .fa_or0(csa_component62_fa37_or0));
  fa fa_csa_component62_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component62_fa38_xor1), .fa_or0(csa_component62_fa38_or0));
  fa fa_csa_component62_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component62_fa39_xor1), .fa_or0(csa_component62_fa39_or0));
  fa fa_csa_component62_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component62_fa40_xor1), .fa_or0(csa_component62_fa40_or0));
  fa fa_csa_component62_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component62_fa41_xor1), .fa_or0(csa_component62_fa41_or0));
  fa fa_csa_component62_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component62_fa42_xor1), .fa_or0(csa_component62_fa42_or0));
  fa fa_csa_component62_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component62_fa43_xor1), .fa_or0(csa_component62_fa43_or0));
  fa fa_csa_component62_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component62_fa44_xor1), .fa_or0(csa_component62_fa44_or0));
  fa fa_csa_component62_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component62_fa45_xor1), .fa_or0(csa_component62_fa45_or0));
  fa fa_csa_component62_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component62_fa46_xor1), .fa_or0(csa_component62_fa46_or0));
  fa fa_csa_component62_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component62_fa47_xor1), .fa_or0(csa_component62_fa47_or0));
  fa fa_csa_component62_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component62_fa48_xor1), .fa_or0(csa_component62_fa48_or0));
  fa fa_csa_component62_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component62_fa49_xor1), .fa_or0(csa_component62_fa49_or0));
  fa fa_csa_component62_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component62_fa50_xor1), .fa_or0(csa_component62_fa50_or0));
  fa fa_csa_component62_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component62_fa51_xor1), .fa_or0(csa_component62_fa51_or0));
  fa fa_csa_component62_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component62_fa52_xor1), .fa_or0(csa_component62_fa52_or0));
  fa fa_csa_component62_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component62_fa53_xor1), .fa_or0(csa_component62_fa53_or0));
  fa fa_csa_component62_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component62_fa54_xor1), .fa_or0(csa_component62_fa54_or0));
  fa fa_csa_component62_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component62_fa55_xor1), .fa_or0(csa_component62_fa55_or0));
  fa fa_csa_component62_fa56_out(.a(a[56]), .b(b[56]), .cin(c[56]), .fa_xor1(csa_component62_fa56_xor1), .fa_or0(csa_component62_fa56_or0));
  fa fa_csa_component62_fa57_out(.a(a[57]), .b(b[57]), .cin(c[57]), .fa_xor1(csa_component62_fa57_xor1), .fa_or0(csa_component62_fa57_or0));
  fa fa_csa_component62_fa58_out(.a(a[58]), .b(b[58]), .cin(c[58]), .fa_xor1(csa_component62_fa58_xor1), .fa_or0(csa_component62_fa58_or0));
  fa fa_csa_component62_fa59_out(.a(a[59]), .b(b[59]), .cin(c[59]), .fa_xor1(csa_component62_fa59_xor1), .fa_or0(csa_component62_fa59_or0));
  fa fa_csa_component62_fa60_out(.a(a[60]), .b(b[60]), .cin(c[60]), .fa_xor1(csa_component62_fa60_xor1), .fa_or0(csa_component62_fa60_or0));
  fa fa_csa_component62_fa61_out(.a(a[61]), .b(b[61]), .cin(c[61]), .fa_xor1(csa_component62_fa61_xor1), .fa_or0(csa_component62_fa61_or0));

  assign csa_component62_out[0] = csa_component62_fa0_xor1[0];
  assign csa_component62_out[1] = csa_component62_fa1_xor1[0];
  assign csa_component62_out[2] = csa_component62_fa2_xor1[0];
  assign csa_component62_out[3] = csa_component62_fa3_xor1[0];
  assign csa_component62_out[4] = csa_component62_fa4_xor1[0];
  assign csa_component62_out[5] = csa_component62_fa5_xor1[0];
  assign csa_component62_out[6] = csa_component62_fa6_xor1[0];
  assign csa_component62_out[7] = csa_component62_fa7_xor1[0];
  assign csa_component62_out[8] = csa_component62_fa8_xor1[0];
  assign csa_component62_out[9] = csa_component62_fa9_xor1[0];
  assign csa_component62_out[10] = csa_component62_fa10_xor1[0];
  assign csa_component62_out[11] = csa_component62_fa11_xor1[0];
  assign csa_component62_out[12] = csa_component62_fa12_xor1[0];
  assign csa_component62_out[13] = csa_component62_fa13_xor1[0];
  assign csa_component62_out[14] = csa_component62_fa14_xor1[0];
  assign csa_component62_out[15] = csa_component62_fa15_xor1[0];
  assign csa_component62_out[16] = csa_component62_fa16_xor1[0];
  assign csa_component62_out[17] = csa_component62_fa17_xor1[0];
  assign csa_component62_out[18] = csa_component62_fa18_xor1[0];
  assign csa_component62_out[19] = csa_component62_fa19_xor1[0];
  assign csa_component62_out[20] = csa_component62_fa20_xor1[0];
  assign csa_component62_out[21] = csa_component62_fa21_xor1[0];
  assign csa_component62_out[22] = csa_component62_fa22_xor1[0];
  assign csa_component62_out[23] = csa_component62_fa23_xor1[0];
  assign csa_component62_out[24] = csa_component62_fa24_xor1[0];
  assign csa_component62_out[25] = csa_component62_fa25_xor1[0];
  assign csa_component62_out[26] = csa_component62_fa26_xor1[0];
  assign csa_component62_out[27] = csa_component62_fa27_xor1[0];
  assign csa_component62_out[28] = csa_component62_fa28_xor1[0];
  assign csa_component62_out[29] = csa_component62_fa29_xor1[0];
  assign csa_component62_out[30] = csa_component62_fa30_xor1[0];
  assign csa_component62_out[31] = csa_component62_fa31_xor1[0];
  assign csa_component62_out[32] = csa_component62_fa32_xor1[0];
  assign csa_component62_out[33] = csa_component62_fa33_xor1[0];
  assign csa_component62_out[34] = csa_component62_fa34_xor1[0];
  assign csa_component62_out[35] = csa_component62_fa35_xor1[0];
  assign csa_component62_out[36] = csa_component62_fa36_xor1[0];
  assign csa_component62_out[37] = csa_component62_fa37_xor1[0];
  assign csa_component62_out[38] = csa_component62_fa38_xor1[0];
  assign csa_component62_out[39] = csa_component62_fa39_xor1[0];
  assign csa_component62_out[40] = csa_component62_fa40_xor1[0];
  assign csa_component62_out[41] = csa_component62_fa41_xor1[0];
  assign csa_component62_out[42] = csa_component62_fa42_xor1[0];
  assign csa_component62_out[43] = csa_component62_fa43_xor1[0];
  assign csa_component62_out[44] = csa_component62_fa44_xor1[0];
  assign csa_component62_out[45] = csa_component62_fa45_xor1[0];
  assign csa_component62_out[46] = csa_component62_fa46_xor1[0];
  assign csa_component62_out[47] = csa_component62_fa47_xor1[0];
  assign csa_component62_out[48] = csa_component62_fa48_xor1[0];
  assign csa_component62_out[49] = csa_component62_fa49_xor1[0];
  assign csa_component62_out[50] = csa_component62_fa50_xor1[0];
  assign csa_component62_out[51] = csa_component62_fa51_xor1[0];
  assign csa_component62_out[52] = csa_component62_fa52_xor1[0];
  assign csa_component62_out[53] = csa_component62_fa53_xor1[0];
  assign csa_component62_out[54] = csa_component62_fa54_xor1[0];
  assign csa_component62_out[55] = csa_component62_fa55_xor1[0];
  assign csa_component62_out[56] = csa_component62_fa56_xor1[0];
  assign csa_component62_out[57] = csa_component62_fa57_xor1[0];
  assign csa_component62_out[58] = csa_component62_fa58_xor1[0];
  assign csa_component62_out[59] = csa_component62_fa59_xor1[0];
  assign csa_component62_out[60] = csa_component62_fa60_xor1[0];
  assign csa_component62_out[61] = csa_component62_fa61_xor1[0];
  assign csa_component62_out[62] = 1'b0;
  assign csa_component62_out[63] = 1'b0;
  assign csa_component62_out[64] = csa_component62_fa0_or0[0];
  assign csa_component62_out[65] = csa_component62_fa1_or0[0];
  assign csa_component62_out[66] = csa_component62_fa2_or0[0];
  assign csa_component62_out[67] = csa_component62_fa3_or0[0];
  assign csa_component62_out[68] = csa_component62_fa4_or0[0];
  assign csa_component62_out[69] = csa_component62_fa5_or0[0];
  assign csa_component62_out[70] = csa_component62_fa6_or0[0];
  assign csa_component62_out[71] = csa_component62_fa7_or0[0];
  assign csa_component62_out[72] = csa_component62_fa8_or0[0];
  assign csa_component62_out[73] = csa_component62_fa9_or0[0];
  assign csa_component62_out[74] = csa_component62_fa10_or0[0];
  assign csa_component62_out[75] = csa_component62_fa11_or0[0];
  assign csa_component62_out[76] = csa_component62_fa12_or0[0];
  assign csa_component62_out[77] = csa_component62_fa13_or0[0];
  assign csa_component62_out[78] = csa_component62_fa14_or0[0];
  assign csa_component62_out[79] = csa_component62_fa15_or0[0];
  assign csa_component62_out[80] = csa_component62_fa16_or0[0];
  assign csa_component62_out[81] = csa_component62_fa17_or0[0];
  assign csa_component62_out[82] = csa_component62_fa18_or0[0];
  assign csa_component62_out[83] = csa_component62_fa19_or0[0];
  assign csa_component62_out[84] = csa_component62_fa20_or0[0];
  assign csa_component62_out[85] = csa_component62_fa21_or0[0];
  assign csa_component62_out[86] = csa_component62_fa22_or0[0];
  assign csa_component62_out[87] = csa_component62_fa23_or0[0];
  assign csa_component62_out[88] = csa_component62_fa24_or0[0];
  assign csa_component62_out[89] = csa_component62_fa25_or0[0];
  assign csa_component62_out[90] = csa_component62_fa26_or0[0];
  assign csa_component62_out[91] = csa_component62_fa27_or0[0];
  assign csa_component62_out[92] = csa_component62_fa28_or0[0];
  assign csa_component62_out[93] = csa_component62_fa29_or0[0];
  assign csa_component62_out[94] = csa_component62_fa30_or0[0];
  assign csa_component62_out[95] = csa_component62_fa31_or0[0];
  assign csa_component62_out[96] = csa_component62_fa32_or0[0];
  assign csa_component62_out[97] = csa_component62_fa33_or0[0];
  assign csa_component62_out[98] = csa_component62_fa34_or0[0];
  assign csa_component62_out[99] = csa_component62_fa35_or0[0];
  assign csa_component62_out[100] = csa_component62_fa36_or0[0];
  assign csa_component62_out[101] = csa_component62_fa37_or0[0];
  assign csa_component62_out[102] = csa_component62_fa38_or0[0];
  assign csa_component62_out[103] = csa_component62_fa39_or0[0];
  assign csa_component62_out[104] = csa_component62_fa40_or0[0];
  assign csa_component62_out[105] = csa_component62_fa41_or0[0];
  assign csa_component62_out[106] = csa_component62_fa42_or0[0];
  assign csa_component62_out[107] = csa_component62_fa43_or0[0];
  assign csa_component62_out[108] = csa_component62_fa44_or0[0];
  assign csa_component62_out[109] = csa_component62_fa45_or0[0];
  assign csa_component62_out[110] = csa_component62_fa46_or0[0];
  assign csa_component62_out[111] = csa_component62_fa47_or0[0];
  assign csa_component62_out[112] = csa_component62_fa48_or0[0];
  assign csa_component62_out[113] = csa_component62_fa49_or0[0];
  assign csa_component62_out[114] = csa_component62_fa50_or0[0];
  assign csa_component62_out[115] = csa_component62_fa51_or0[0];
  assign csa_component62_out[116] = csa_component62_fa52_or0[0];
  assign csa_component62_out[117] = csa_component62_fa53_or0[0];
  assign csa_component62_out[118] = csa_component62_fa54_or0[0];
  assign csa_component62_out[119] = csa_component62_fa55_or0[0];
  assign csa_component62_out[120] = csa_component62_fa56_or0[0];
  assign csa_component62_out[121] = csa_component62_fa57_or0[0];
  assign csa_component62_out[122] = csa_component62_fa58_or0[0];
  assign csa_component62_out[123] = csa_component62_fa59_or0[0];
  assign csa_component62_out[124] = csa_component62_fa60_or0[0];
  assign csa_component62_out[125] = csa_component62_fa61_or0[0];
endmodule

module csa_component42(input [41:0] a, input [41:0] b, input [41:0] c, output [85:0] csa_component42_out);
  wire [0:0] csa_component42_fa0_xor1;
  wire [0:0] csa_component42_fa0_or0;
  wire [0:0] csa_component42_fa1_xor1;
  wire [0:0] csa_component42_fa1_or0;
  wire [0:0] csa_component42_fa2_xor1;
  wire [0:0] csa_component42_fa2_or0;
  wire [0:0] csa_component42_fa3_xor1;
  wire [0:0] csa_component42_fa3_or0;
  wire [0:0] csa_component42_fa4_xor1;
  wire [0:0] csa_component42_fa4_or0;
  wire [0:0] csa_component42_fa5_xor1;
  wire [0:0] csa_component42_fa5_or0;
  wire [0:0] csa_component42_fa6_xor1;
  wire [0:0] csa_component42_fa6_or0;
  wire [0:0] csa_component42_fa7_xor1;
  wire [0:0] csa_component42_fa7_or0;
  wire [0:0] csa_component42_fa8_xor1;
  wire [0:0] csa_component42_fa8_or0;
  wire [0:0] csa_component42_fa9_xor1;
  wire [0:0] csa_component42_fa9_or0;
  wire [0:0] csa_component42_fa10_xor1;
  wire [0:0] csa_component42_fa10_or0;
  wire [0:0] csa_component42_fa11_xor1;
  wire [0:0] csa_component42_fa11_or0;
  wire [0:0] csa_component42_fa12_xor1;
  wire [0:0] csa_component42_fa12_or0;
  wire [0:0] csa_component42_fa13_xor1;
  wire [0:0] csa_component42_fa13_or0;
  wire [0:0] csa_component42_fa14_xor1;
  wire [0:0] csa_component42_fa14_or0;
  wire [0:0] csa_component42_fa15_xor1;
  wire [0:0] csa_component42_fa15_or0;
  wire [0:0] csa_component42_fa16_xor1;
  wire [0:0] csa_component42_fa16_or0;
  wire [0:0] csa_component42_fa17_xor1;
  wire [0:0] csa_component42_fa17_or0;
  wire [0:0] csa_component42_fa18_xor1;
  wire [0:0] csa_component42_fa18_or0;
  wire [0:0] csa_component42_fa19_xor1;
  wire [0:0] csa_component42_fa19_or0;
  wire [0:0] csa_component42_fa20_xor1;
  wire [0:0] csa_component42_fa20_or0;
  wire [0:0] csa_component42_fa21_xor1;
  wire [0:0] csa_component42_fa21_or0;
  wire [0:0] csa_component42_fa22_xor1;
  wire [0:0] csa_component42_fa22_or0;
  wire [0:0] csa_component42_fa23_xor1;
  wire [0:0] csa_component42_fa23_or0;
  wire [0:0] csa_component42_fa24_xor1;
  wire [0:0] csa_component42_fa24_or0;
  wire [0:0] csa_component42_fa25_xor1;
  wire [0:0] csa_component42_fa25_or0;
  wire [0:0] csa_component42_fa26_xor1;
  wire [0:0] csa_component42_fa26_or0;
  wire [0:0] csa_component42_fa27_xor1;
  wire [0:0] csa_component42_fa27_or0;
  wire [0:0] csa_component42_fa28_xor1;
  wire [0:0] csa_component42_fa28_or0;
  wire [0:0] csa_component42_fa29_xor1;
  wire [0:0] csa_component42_fa29_or0;
  wire [0:0] csa_component42_fa30_xor1;
  wire [0:0] csa_component42_fa30_or0;
  wire [0:0] csa_component42_fa31_xor1;
  wire [0:0] csa_component42_fa31_or0;
  wire [0:0] csa_component42_fa32_xor1;
  wire [0:0] csa_component42_fa32_or0;
  wire [0:0] csa_component42_fa33_xor1;
  wire [0:0] csa_component42_fa33_or0;
  wire [0:0] csa_component42_fa34_xor1;
  wire [0:0] csa_component42_fa34_or0;
  wire [0:0] csa_component42_fa35_xor1;
  wire [0:0] csa_component42_fa35_or0;
  wire [0:0] csa_component42_fa36_xor1;
  wire [0:0] csa_component42_fa36_or0;
  wire [0:0] csa_component42_fa37_xor1;
  wire [0:0] csa_component42_fa37_or0;
  wire [0:0] csa_component42_fa38_xor1;
  wire [0:0] csa_component42_fa38_or0;
  wire [0:0] csa_component42_fa39_xor1;
  wire [0:0] csa_component42_fa39_or0;
  wire [0:0] csa_component42_fa40_xor1;
  wire [0:0] csa_component42_fa40_or0;
  wire [0:0] csa_component42_fa41_xor1;
  wire [0:0] csa_component42_fa41_or0;

  fa fa_csa_component42_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component42_fa0_xor1), .fa_or0(csa_component42_fa0_or0));
  fa fa_csa_component42_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component42_fa1_xor1), .fa_or0(csa_component42_fa1_or0));
  fa fa_csa_component42_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component42_fa2_xor1), .fa_or0(csa_component42_fa2_or0));
  fa fa_csa_component42_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component42_fa3_xor1), .fa_or0(csa_component42_fa3_or0));
  fa fa_csa_component42_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component42_fa4_xor1), .fa_or0(csa_component42_fa4_or0));
  fa fa_csa_component42_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component42_fa5_xor1), .fa_or0(csa_component42_fa5_or0));
  fa fa_csa_component42_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component42_fa6_xor1), .fa_or0(csa_component42_fa6_or0));
  fa fa_csa_component42_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component42_fa7_xor1), .fa_or0(csa_component42_fa7_or0));
  fa fa_csa_component42_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component42_fa8_xor1), .fa_or0(csa_component42_fa8_or0));
  fa fa_csa_component42_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component42_fa9_xor1), .fa_or0(csa_component42_fa9_or0));
  fa fa_csa_component42_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component42_fa10_xor1), .fa_or0(csa_component42_fa10_or0));
  fa fa_csa_component42_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component42_fa11_xor1), .fa_or0(csa_component42_fa11_or0));
  fa fa_csa_component42_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component42_fa12_xor1), .fa_or0(csa_component42_fa12_or0));
  fa fa_csa_component42_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component42_fa13_xor1), .fa_or0(csa_component42_fa13_or0));
  fa fa_csa_component42_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component42_fa14_xor1), .fa_or0(csa_component42_fa14_or0));
  fa fa_csa_component42_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component42_fa15_xor1), .fa_or0(csa_component42_fa15_or0));
  fa fa_csa_component42_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component42_fa16_xor1), .fa_or0(csa_component42_fa16_or0));
  fa fa_csa_component42_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component42_fa17_xor1), .fa_or0(csa_component42_fa17_or0));
  fa fa_csa_component42_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component42_fa18_xor1), .fa_or0(csa_component42_fa18_or0));
  fa fa_csa_component42_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component42_fa19_xor1), .fa_or0(csa_component42_fa19_or0));
  fa fa_csa_component42_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component42_fa20_xor1), .fa_or0(csa_component42_fa20_or0));
  fa fa_csa_component42_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component42_fa21_xor1), .fa_or0(csa_component42_fa21_or0));
  fa fa_csa_component42_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component42_fa22_xor1), .fa_or0(csa_component42_fa22_or0));
  fa fa_csa_component42_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component42_fa23_xor1), .fa_or0(csa_component42_fa23_or0));
  fa fa_csa_component42_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component42_fa24_xor1), .fa_or0(csa_component42_fa24_or0));
  fa fa_csa_component42_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component42_fa25_xor1), .fa_or0(csa_component42_fa25_or0));
  fa fa_csa_component42_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component42_fa26_xor1), .fa_or0(csa_component42_fa26_or0));
  fa fa_csa_component42_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component42_fa27_xor1), .fa_or0(csa_component42_fa27_or0));
  fa fa_csa_component42_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component42_fa28_xor1), .fa_or0(csa_component42_fa28_or0));
  fa fa_csa_component42_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component42_fa29_xor1), .fa_or0(csa_component42_fa29_or0));
  fa fa_csa_component42_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component42_fa30_xor1), .fa_or0(csa_component42_fa30_or0));
  fa fa_csa_component42_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component42_fa31_xor1), .fa_or0(csa_component42_fa31_or0));
  fa fa_csa_component42_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component42_fa32_xor1), .fa_or0(csa_component42_fa32_or0));
  fa fa_csa_component42_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component42_fa33_xor1), .fa_or0(csa_component42_fa33_or0));
  fa fa_csa_component42_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component42_fa34_xor1), .fa_or0(csa_component42_fa34_or0));
  fa fa_csa_component42_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component42_fa35_xor1), .fa_or0(csa_component42_fa35_or0));
  fa fa_csa_component42_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component42_fa36_xor1), .fa_or0(csa_component42_fa36_or0));
  fa fa_csa_component42_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component42_fa37_xor1), .fa_or0(csa_component42_fa37_or0));
  fa fa_csa_component42_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component42_fa38_xor1), .fa_or0(csa_component42_fa38_or0));
  fa fa_csa_component42_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component42_fa39_xor1), .fa_or0(csa_component42_fa39_or0));
  fa fa_csa_component42_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component42_fa40_xor1), .fa_or0(csa_component42_fa40_or0));
  fa fa_csa_component42_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component42_fa41_xor1), .fa_or0(csa_component42_fa41_or0));

  assign csa_component42_out[0] = csa_component42_fa0_xor1[0];
  assign csa_component42_out[1] = csa_component42_fa1_xor1[0];
  assign csa_component42_out[2] = csa_component42_fa2_xor1[0];
  assign csa_component42_out[3] = csa_component42_fa3_xor1[0];
  assign csa_component42_out[4] = csa_component42_fa4_xor1[0];
  assign csa_component42_out[5] = csa_component42_fa5_xor1[0];
  assign csa_component42_out[6] = csa_component42_fa6_xor1[0];
  assign csa_component42_out[7] = csa_component42_fa7_xor1[0];
  assign csa_component42_out[8] = csa_component42_fa8_xor1[0];
  assign csa_component42_out[9] = csa_component42_fa9_xor1[0];
  assign csa_component42_out[10] = csa_component42_fa10_xor1[0];
  assign csa_component42_out[11] = csa_component42_fa11_xor1[0];
  assign csa_component42_out[12] = csa_component42_fa12_xor1[0];
  assign csa_component42_out[13] = csa_component42_fa13_xor1[0];
  assign csa_component42_out[14] = csa_component42_fa14_xor1[0];
  assign csa_component42_out[15] = csa_component42_fa15_xor1[0];
  assign csa_component42_out[16] = csa_component42_fa16_xor1[0];
  assign csa_component42_out[17] = csa_component42_fa17_xor1[0];
  assign csa_component42_out[18] = csa_component42_fa18_xor1[0];
  assign csa_component42_out[19] = csa_component42_fa19_xor1[0];
  assign csa_component42_out[20] = csa_component42_fa20_xor1[0];
  assign csa_component42_out[21] = csa_component42_fa21_xor1[0];
  assign csa_component42_out[22] = csa_component42_fa22_xor1[0];
  assign csa_component42_out[23] = csa_component42_fa23_xor1[0];
  assign csa_component42_out[24] = csa_component42_fa24_xor1[0];
  assign csa_component42_out[25] = csa_component42_fa25_xor1[0];
  assign csa_component42_out[26] = csa_component42_fa26_xor1[0];
  assign csa_component42_out[27] = csa_component42_fa27_xor1[0];
  assign csa_component42_out[28] = csa_component42_fa28_xor1[0];
  assign csa_component42_out[29] = csa_component42_fa29_xor1[0];
  assign csa_component42_out[30] = csa_component42_fa30_xor1[0];
  assign csa_component42_out[31] = csa_component42_fa31_xor1[0];
  assign csa_component42_out[32] = csa_component42_fa32_xor1[0];
  assign csa_component42_out[33] = csa_component42_fa33_xor1[0];
  assign csa_component42_out[34] = csa_component42_fa34_xor1[0];
  assign csa_component42_out[35] = csa_component42_fa35_xor1[0];
  assign csa_component42_out[36] = csa_component42_fa36_xor1[0];
  assign csa_component42_out[37] = csa_component42_fa37_xor1[0];
  assign csa_component42_out[38] = csa_component42_fa38_xor1[0];
  assign csa_component42_out[39] = csa_component42_fa39_xor1[0];
  assign csa_component42_out[40] = csa_component42_fa40_xor1[0];
  assign csa_component42_out[41] = csa_component42_fa41_xor1[0];
  assign csa_component42_out[42] = 1'b0;
  assign csa_component42_out[43] = 1'b0;
  assign csa_component42_out[44] = csa_component42_fa0_or0[0];
  assign csa_component42_out[45] = csa_component42_fa1_or0[0];
  assign csa_component42_out[46] = csa_component42_fa2_or0[0];
  assign csa_component42_out[47] = csa_component42_fa3_or0[0];
  assign csa_component42_out[48] = csa_component42_fa4_or0[0];
  assign csa_component42_out[49] = csa_component42_fa5_or0[0];
  assign csa_component42_out[50] = csa_component42_fa6_or0[0];
  assign csa_component42_out[51] = csa_component42_fa7_or0[0];
  assign csa_component42_out[52] = csa_component42_fa8_or0[0];
  assign csa_component42_out[53] = csa_component42_fa9_or0[0];
  assign csa_component42_out[54] = csa_component42_fa10_or0[0];
  assign csa_component42_out[55] = csa_component42_fa11_or0[0];
  assign csa_component42_out[56] = csa_component42_fa12_or0[0];
  assign csa_component42_out[57] = csa_component42_fa13_or0[0];
  assign csa_component42_out[58] = csa_component42_fa14_or0[0];
  assign csa_component42_out[59] = csa_component42_fa15_or0[0];
  assign csa_component42_out[60] = csa_component42_fa16_or0[0];
  assign csa_component42_out[61] = csa_component42_fa17_or0[0];
  assign csa_component42_out[62] = csa_component42_fa18_or0[0];
  assign csa_component42_out[63] = csa_component42_fa19_or0[0];
  assign csa_component42_out[64] = csa_component42_fa20_or0[0];
  assign csa_component42_out[65] = csa_component42_fa21_or0[0];
  assign csa_component42_out[66] = csa_component42_fa22_or0[0];
  assign csa_component42_out[67] = csa_component42_fa23_or0[0];
  assign csa_component42_out[68] = csa_component42_fa24_or0[0];
  assign csa_component42_out[69] = csa_component42_fa25_or0[0];
  assign csa_component42_out[70] = csa_component42_fa26_or0[0];
  assign csa_component42_out[71] = csa_component42_fa27_or0[0];
  assign csa_component42_out[72] = csa_component42_fa28_or0[0];
  assign csa_component42_out[73] = csa_component42_fa29_or0[0];
  assign csa_component42_out[74] = csa_component42_fa30_or0[0];
  assign csa_component42_out[75] = csa_component42_fa31_or0[0];
  assign csa_component42_out[76] = csa_component42_fa32_or0[0];
  assign csa_component42_out[77] = csa_component42_fa33_or0[0];
  assign csa_component42_out[78] = csa_component42_fa34_or0[0];
  assign csa_component42_out[79] = csa_component42_fa35_or0[0];
  assign csa_component42_out[80] = csa_component42_fa36_or0[0];
  assign csa_component42_out[81] = csa_component42_fa37_or0[0];
  assign csa_component42_out[82] = csa_component42_fa38_or0[0];
  assign csa_component42_out[83] = csa_component42_fa39_or0[0];
  assign csa_component42_out[84] = csa_component42_fa40_or0[0];
  assign csa_component42_out[85] = csa_component42_fa41_or0[0];
endmodule

module csa_component48(input [47:0] a, input [47:0] b, input [47:0] c, output [97:0] csa_component48_out);
  wire [0:0] csa_component48_fa0_xor1;
  wire [0:0] csa_component48_fa0_or0;
  wire [0:0] csa_component48_fa1_xor1;
  wire [0:0] csa_component48_fa1_or0;
  wire [0:0] csa_component48_fa2_xor1;
  wire [0:0] csa_component48_fa2_or0;
  wire [0:0] csa_component48_fa3_xor1;
  wire [0:0] csa_component48_fa3_or0;
  wire [0:0] csa_component48_fa4_xor1;
  wire [0:0] csa_component48_fa4_or0;
  wire [0:0] csa_component48_fa5_xor1;
  wire [0:0] csa_component48_fa5_or0;
  wire [0:0] csa_component48_fa6_xor1;
  wire [0:0] csa_component48_fa6_or0;
  wire [0:0] csa_component48_fa7_xor1;
  wire [0:0] csa_component48_fa7_or0;
  wire [0:0] csa_component48_fa8_xor1;
  wire [0:0] csa_component48_fa8_or0;
  wire [0:0] csa_component48_fa9_xor1;
  wire [0:0] csa_component48_fa9_or0;
  wire [0:0] csa_component48_fa10_xor1;
  wire [0:0] csa_component48_fa10_or0;
  wire [0:0] csa_component48_fa11_xor1;
  wire [0:0] csa_component48_fa11_or0;
  wire [0:0] csa_component48_fa12_xor1;
  wire [0:0] csa_component48_fa12_or0;
  wire [0:0] csa_component48_fa13_xor1;
  wire [0:0] csa_component48_fa13_or0;
  wire [0:0] csa_component48_fa14_xor1;
  wire [0:0] csa_component48_fa14_or0;
  wire [0:0] csa_component48_fa15_xor1;
  wire [0:0] csa_component48_fa15_or0;
  wire [0:0] csa_component48_fa16_xor1;
  wire [0:0] csa_component48_fa16_or0;
  wire [0:0] csa_component48_fa17_xor1;
  wire [0:0] csa_component48_fa17_or0;
  wire [0:0] csa_component48_fa18_xor1;
  wire [0:0] csa_component48_fa18_or0;
  wire [0:0] csa_component48_fa19_xor1;
  wire [0:0] csa_component48_fa19_or0;
  wire [0:0] csa_component48_fa20_xor1;
  wire [0:0] csa_component48_fa20_or0;
  wire [0:0] csa_component48_fa21_xor1;
  wire [0:0] csa_component48_fa21_or0;
  wire [0:0] csa_component48_fa22_xor1;
  wire [0:0] csa_component48_fa22_or0;
  wire [0:0] csa_component48_fa23_xor1;
  wire [0:0] csa_component48_fa23_or0;
  wire [0:0] csa_component48_fa24_xor1;
  wire [0:0] csa_component48_fa24_or0;
  wire [0:0] csa_component48_fa25_xor1;
  wire [0:0] csa_component48_fa25_or0;
  wire [0:0] csa_component48_fa26_xor1;
  wire [0:0] csa_component48_fa26_or0;
  wire [0:0] csa_component48_fa27_xor1;
  wire [0:0] csa_component48_fa27_or0;
  wire [0:0] csa_component48_fa28_xor1;
  wire [0:0] csa_component48_fa28_or0;
  wire [0:0] csa_component48_fa29_xor1;
  wire [0:0] csa_component48_fa29_or0;
  wire [0:0] csa_component48_fa30_xor1;
  wire [0:0] csa_component48_fa30_or0;
  wire [0:0] csa_component48_fa31_xor1;
  wire [0:0] csa_component48_fa31_or0;
  wire [0:0] csa_component48_fa32_xor1;
  wire [0:0] csa_component48_fa32_or0;
  wire [0:0] csa_component48_fa33_xor1;
  wire [0:0] csa_component48_fa33_or0;
  wire [0:0] csa_component48_fa34_xor1;
  wire [0:0] csa_component48_fa34_or0;
  wire [0:0] csa_component48_fa35_xor1;
  wire [0:0] csa_component48_fa35_or0;
  wire [0:0] csa_component48_fa36_xor1;
  wire [0:0] csa_component48_fa36_or0;
  wire [0:0] csa_component48_fa37_xor1;
  wire [0:0] csa_component48_fa37_or0;
  wire [0:0] csa_component48_fa38_xor1;
  wire [0:0] csa_component48_fa38_or0;
  wire [0:0] csa_component48_fa39_xor1;
  wire [0:0] csa_component48_fa39_or0;
  wire [0:0] csa_component48_fa40_xor1;
  wire [0:0] csa_component48_fa40_or0;
  wire [0:0] csa_component48_fa41_xor1;
  wire [0:0] csa_component48_fa41_or0;
  wire [0:0] csa_component48_fa42_xor1;
  wire [0:0] csa_component48_fa42_or0;
  wire [0:0] csa_component48_fa43_xor1;
  wire [0:0] csa_component48_fa43_or0;
  wire [0:0] csa_component48_fa44_xor1;
  wire [0:0] csa_component48_fa44_or0;
  wire [0:0] csa_component48_fa45_xor1;
  wire [0:0] csa_component48_fa45_or0;
  wire [0:0] csa_component48_fa46_xor1;
  wire [0:0] csa_component48_fa46_or0;
  wire [0:0] csa_component48_fa47_xor1;
  wire [0:0] csa_component48_fa47_or0;

  fa fa_csa_component48_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component48_fa0_xor1), .fa_or0(csa_component48_fa0_or0));
  fa fa_csa_component48_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component48_fa1_xor1), .fa_or0(csa_component48_fa1_or0));
  fa fa_csa_component48_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component48_fa2_xor1), .fa_or0(csa_component48_fa2_or0));
  fa fa_csa_component48_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component48_fa3_xor1), .fa_or0(csa_component48_fa3_or0));
  fa fa_csa_component48_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component48_fa4_xor1), .fa_or0(csa_component48_fa4_or0));
  fa fa_csa_component48_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component48_fa5_xor1), .fa_or0(csa_component48_fa5_or0));
  fa fa_csa_component48_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component48_fa6_xor1), .fa_or0(csa_component48_fa6_or0));
  fa fa_csa_component48_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component48_fa7_xor1), .fa_or0(csa_component48_fa7_or0));
  fa fa_csa_component48_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component48_fa8_xor1), .fa_or0(csa_component48_fa8_or0));
  fa fa_csa_component48_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component48_fa9_xor1), .fa_or0(csa_component48_fa9_or0));
  fa fa_csa_component48_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component48_fa10_xor1), .fa_or0(csa_component48_fa10_or0));
  fa fa_csa_component48_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component48_fa11_xor1), .fa_or0(csa_component48_fa11_or0));
  fa fa_csa_component48_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component48_fa12_xor1), .fa_or0(csa_component48_fa12_or0));
  fa fa_csa_component48_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component48_fa13_xor1), .fa_or0(csa_component48_fa13_or0));
  fa fa_csa_component48_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component48_fa14_xor1), .fa_or0(csa_component48_fa14_or0));
  fa fa_csa_component48_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component48_fa15_xor1), .fa_or0(csa_component48_fa15_or0));
  fa fa_csa_component48_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component48_fa16_xor1), .fa_or0(csa_component48_fa16_or0));
  fa fa_csa_component48_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component48_fa17_xor1), .fa_or0(csa_component48_fa17_or0));
  fa fa_csa_component48_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component48_fa18_xor1), .fa_or0(csa_component48_fa18_or0));
  fa fa_csa_component48_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component48_fa19_xor1), .fa_or0(csa_component48_fa19_or0));
  fa fa_csa_component48_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component48_fa20_xor1), .fa_or0(csa_component48_fa20_or0));
  fa fa_csa_component48_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component48_fa21_xor1), .fa_or0(csa_component48_fa21_or0));
  fa fa_csa_component48_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component48_fa22_xor1), .fa_or0(csa_component48_fa22_or0));
  fa fa_csa_component48_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component48_fa23_xor1), .fa_or0(csa_component48_fa23_or0));
  fa fa_csa_component48_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component48_fa24_xor1), .fa_or0(csa_component48_fa24_or0));
  fa fa_csa_component48_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component48_fa25_xor1), .fa_or0(csa_component48_fa25_or0));
  fa fa_csa_component48_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component48_fa26_xor1), .fa_or0(csa_component48_fa26_or0));
  fa fa_csa_component48_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component48_fa27_xor1), .fa_or0(csa_component48_fa27_or0));
  fa fa_csa_component48_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component48_fa28_xor1), .fa_or0(csa_component48_fa28_or0));
  fa fa_csa_component48_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component48_fa29_xor1), .fa_or0(csa_component48_fa29_or0));
  fa fa_csa_component48_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component48_fa30_xor1), .fa_or0(csa_component48_fa30_or0));
  fa fa_csa_component48_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component48_fa31_xor1), .fa_or0(csa_component48_fa31_or0));
  fa fa_csa_component48_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component48_fa32_xor1), .fa_or0(csa_component48_fa32_or0));
  fa fa_csa_component48_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component48_fa33_xor1), .fa_or0(csa_component48_fa33_or0));
  fa fa_csa_component48_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component48_fa34_xor1), .fa_or0(csa_component48_fa34_or0));
  fa fa_csa_component48_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component48_fa35_xor1), .fa_or0(csa_component48_fa35_or0));
  fa fa_csa_component48_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component48_fa36_xor1), .fa_or0(csa_component48_fa36_or0));
  fa fa_csa_component48_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component48_fa37_xor1), .fa_or0(csa_component48_fa37_or0));
  fa fa_csa_component48_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component48_fa38_xor1), .fa_or0(csa_component48_fa38_or0));
  fa fa_csa_component48_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component48_fa39_xor1), .fa_or0(csa_component48_fa39_or0));
  fa fa_csa_component48_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component48_fa40_xor1), .fa_or0(csa_component48_fa40_or0));
  fa fa_csa_component48_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component48_fa41_xor1), .fa_or0(csa_component48_fa41_or0));
  fa fa_csa_component48_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component48_fa42_xor1), .fa_or0(csa_component48_fa42_or0));
  fa fa_csa_component48_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component48_fa43_xor1), .fa_or0(csa_component48_fa43_or0));
  fa fa_csa_component48_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component48_fa44_xor1), .fa_or0(csa_component48_fa44_or0));
  fa fa_csa_component48_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component48_fa45_xor1), .fa_or0(csa_component48_fa45_or0));
  fa fa_csa_component48_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component48_fa46_xor1), .fa_or0(csa_component48_fa46_or0));
  fa fa_csa_component48_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component48_fa47_xor1), .fa_or0(csa_component48_fa47_or0));

  assign csa_component48_out[0] = csa_component48_fa0_xor1[0];
  assign csa_component48_out[1] = csa_component48_fa1_xor1[0];
  assign csa_component48_out[2] = csa_component48_fa2_xor1[0];
  assign csa_component48_out[3] = csa_component48_fa3_xor1[0];
  assign csa_component48_out[4] = csa_component48_fa4_xor1[0];
  assign csa_component48_out[5] = csa_component48_fa5_xor1[0];
  assign csa_component48_out[6] = csa_component48_fa6_xor1[0];
  assign csa_component48_out[7] = csa_component48_fa7_xor1[0];
  assign csa_component48_out[8] = csa_component48_fa8_xor1[0];
  assign csa_component48_out[9] = csa_component48_fa9_xor1[0];
  assign csa_component48_out[10] = csa_component48_fa10_xor1[0];
  assign csa_component48_out[11] = csa_component48_fa11_xor1[0];
  assign csa_component48_out[12] = csa_component48_fa12_xor1[0];
  assign csa_component48_out[13] = csa_component48_fa13_xor1[0];
  assign csa_component48_out[14] = csa_component48_fa14_xor1[0];
  assign csa_component48_out[15] = csa_component48_fa15_xor1[0];
  assign csa_component48_out[16] = csa_component48_fa16_xor1[0];
  assign csa_component48_out[17] = csa_component48_fa17_xor1[0];
  assign csa_component48_out[18] = csa_component48_fa18_xor1[0];
  assign csa_component48_out[19] = csa_component48_fa19_xor1[0];
  assign csa_component48_out[20] = csa_component48_fa20_xor1[0];
  assign csa_component48_out[21] = csa_component48_fa21_xor1[0];
  assign csa_component48_out[22] = csa_component48_fa22_xor1[0];
  assign csa_component48_out[23] = csa_component48_fa23_xor1[0];
  assign csa_component48_out[24] = csa_component48_fa24_xor1[0];
  assign csa_component48_out[25] = csa_component48_fa25_xor1[0];
  assign csa_component48_out[26] = csa_component48_fa26_xor1[0];
  assign csa_component48_out[27] = csa_component48_fa27_xor1[0];
  assign csa_component48_out[28] = csa_component48_fa28_xor1[0];
  assign csa_component48_out[29] = csa_component48_fa29_xor1[0];
  assign csa_component48_out[30] = csa_component48_fa30_xor1[0];
  assign csa_component48_out[31] = csa_component48_fa31_xor1[0];
  assign csa_component48_out[32] = csa_component48_fa32_xor1[0];
  assign csa_component48_out[33] = csa_component48_fa33_xor1[0];
  assign csa_component48_out[34] = csa_component48_fa34_xor1[0];
  assign csa_component48_out[35] = csa_component48_fa35_xor1[0];
  assign csa_component48_out[36] = csa_component48_fa36_xor1[0];
  assign csa_component48_out[37] = csa_component48_fa37_xor1[0];
  assign csa_component48_out[38] = csa_component48_fa38_xor1[0];
  assign csa_component48_out[39] = csa_component48_fa39_xor1[0];
  assign csa_component48_out[40] = csa_component48_fa40_xor1[0];
  assign csa_component48_out[41] = csa_component48_fa41_xor1[0];
  assign csa_component48_out[42] = csa_component48_fa42_xor1[0];
  assign csa_component48_out[43] = csa_component48_fa43_xor1[0];
  assign csa_component48_out[44] = csa_component48_fa44_xor1[0];
  assign csa_component48_out[45] = csa_component48_fa45_xor1[0];
  assign csa_component48_out[46] = csa_component48_fa46_xor1[0];
  assign csa_component48_out[47] = csa_component48_fa47_xor1[0];
  assign csa_component48_out[48] = 1'b0;
  assign csa_component48_out[49] = 1'b0;
  assign csa_component48_out[50] = csa_component48_fa0_or0[0];
  assign csa_component48_out[51] = csa_component48_fa1_or0[0];
  assign csa_component48_out[52] = csa_component48_fa2_or0[0];
  assign csa_component48_out[53] = csa_component48_fa3_or0[0];
  assign csa_component48_out[54] = csa_component48_fa4_or0[0];
  assign csa_component48_out[55] = csa_component48_fa5_or0[0];
  assign csa_component48_out[56] = csa_component48_fa6_or0[0];
  assign csa_component48_out[57] = csa_component48_fa7_or0[0];
  assign csa_component48_out[58] = csa_component48_fa8_or0[0];
  assign csa_component48_out[59] = csa_component48_fa9_or0[0];
  assign csa_component48_out[60] = csa_component48_fa10_or0[0];
  assign csa_component48_out[61] = csa_component48_fa11_or0[0];
  assign csa_component48_out[62] = csa_component48_fa12_or0[0];
  assign csa_component48_out[63] = csa_component48_fa13_or0[0];
  assign csa_component48_out[64] = csa_component48_fa14_or0[0];
  assign csa_component48_out[65] = csa_component48_fa15_or0[0];
  assign csa_component48_out[66] = csa_component48_fa16_or0[0];
  assign csa_component48_out[67] = csa_component48_fa17_or0[0];
  assign csa_component48_out[68] = csa_component48_fa18_or0[0];
  assign csa_component48_out[69] = csa_component48_fa19_or0[0];
  assign csa_component48_out[70] = csa_component48_fa20_or0[0];
  assign csa_component48_out[71] = csa_component48_fa21_or0[0];
  assign csa_component48_out[72] = csa_component48_fa22_or0[0];
  assign csa_component48_out[73] = csa_component48_fa23_or0[0];
  assign csa_component48_out[74] = csa_component48_fa24_or0[0];
  assign csa_component48_out[75] = csa_component48_fa25_or0[0];
  assign csa_component48_out[76] = csa_component48_fa26_or0[0];
  assign csa_component48_out[77] = csa_component48_fa27_or0[0];
  assign csa_component48_out[78] = csa_component48_fa28_or0[0];
  assign csa_component48_out[79] = csa_component48_fa29_or0[0];
  assign csa_component48_out[80] = csa_component48_fa30_or0[0];
  assign csa_component48_out[81] = csa_component48_fa31_or0[0];
  assign csa_component48_out[82] = csa_component48_fa32_or0[0];
  assign csa_component48_out[83] = csa_component48_fa33_or0[0];
  assign csa_component48_out[84] = csa_component48_fa34_or0[0];
  assign csa_component48_out[85] = csa_component48_fa35_or0[0];
  assign csa_component48_out[86] = csa_component48_fa36_or0[0];
  assign csa_component48_out[87] = csa_component48_fa37_or0[0];
  assign csa_component48_out[88] = csa_component48_fa38_or0[0];
  assign csa_component48_out[89] = csa_component48_fa39_or0[0];
  assign csa_component48_out[90] = csa_component48_fa40_or0[0];
  assign csa_component48_out[91] = csa_component48_fa41_or0[0];
  assign csa_component48_out[92] = csa_component48_fa42_or0[0];
  assign csa_component48_out[93] = csa_component48_fa43_or0[0];
  assign csa_component48_out[94] = csa_component48_fa44_or0[0];
  assign csa_component48_out[95] = csa_component48_fa45_or0[0];
  assign csa_component48_out[96] = csa_component48_fa46_or0[0];
  assign csa_component48_out[97] = csa_component48_fa47_or0[0];
endmodule

module csa_component57(input [56:0] a, input [56:0] b, input [56:0] c, output [115:0] csa_component57_out);
  wire [0:0] csa_component57_fa0_xor1;
  wire [0:0] csa_component57_fa0_or0;
  wire [0:0] csa_component57_fa1_xor1;
  wire [0:0] csa_component57_fa1_or0;
  wire [0:0] csa_component57_fa2_xor1;
  wire [0:0] csa_component57_fa2_or0;
  wire [0:0] csa_component57_fa3_xor1;
  wire [0:0] csa_component57_fa3_or0;
  wire [0:0] csa_component57_fa4_xor1;
  wire [0:0] csa_component57_fa4_or0;
  wire [0:0] csa_component57_fa5_xor1;
  wire [0:0] csa_component57_fa5_or0;
  wire [0:0] csa_component57_fa6_xor1;
  wire [0:0] csa_component57_fa6_or0;
  wire [0:0] csa_component57_fa7_xor1;
  wire [0:0] csa_component57_fa7_or0;
  wire [0:0] csa_component57_fa8_xor1;
  wire [0:0] csa_component57_fa8_or0;
  wire [0:0] csa_component57_fa9_xor1;
  wire [0:0] csa_component57_fa9_or0;
  wire [0:0] csa_component57_fa10_xor1;
  wire [0:0] csa_component57_fa10_or0;
  wire [0:0] csa_component57_fa11_xor1;
  wire [0:0] csa_component57_fa11_or0;
  wire [0:0] csa_component57_fa12_xor1;
  wire [0:0] csa_component57_fa12_or0;
  wire [0:0] csa_component57_fa13_xor1;
  wire [0:0] csa_component57_fa13_or0;
  wire [0:0] csa_component57_fa14_xor1;
  wire [0:0] csa_component57_fa14_or0;
  wire [0:0] csa_component57_fa15_xor1;
  wire [0:0] csa_component57_fa15_or0;
  wire [0:0] csa_component57_fa16_xor1;
  wire [0:0] csa_component57_fa16_or0;
  wire [0:0] csa_component57_fa17_xor1;
  wire [0:0] csa_component57_fa17_or0;
  wire [0:0] csa_component57_fa18_xor1;
  wire [0:0] csa_component57_fa18_or0;
  wire [0:0] csa_component57_fa19_xor1;
  wire [0:0] csa_component57_fa19_or0;
  wire [0:0] csa_component57_fa20_xor1;
  wire [0:0] csa_component57_fa20_or0;
  wire [0:0] csa_component57_fa21_xor1;
  wire [0:0] csa_component57_fa21_or0;
  wire [0:0] csa_component57_fa22_xor1;
  wire [0:0] csa_component57_fa22_or0;
  wire [0:0] csa_component57_fa23_xor1;
  wire [0:0] csa_component57_fa23_or0;
  wire [0:0] csa_component57_fa24_xor1;
  wire [0:0] csa_component57_fa24_or0;
  wire [0:0] csa_component57_fa25_xor1;
  wire [0:0] csa_component57_fa25_or0;
  wire [0:0] csa_component57_fa26_xor1;
  wire [0:0] csa_component57_fa26_or0;
  wire [0:0] csa_component57_fa27_xor1;
  wire [0:0] csa_component57_fa27_or0;
  wire [0:0] csa_component57_fa28_xor1;
  wire [0:0] csa_component57_fa28_or0;
  wire [0:0] csa_component57_fa29_xor1;
  wire [0:0] csa_component57_fa29_or0;
  wire [0:0] csa_component57_fa30_xor1;
  wire [0:0] csa_component57_fa30_or0;
  wire [0:0] csa_component57_fa31_xor1;
  wire [0:0] csa_component57_fa31_or0;
  wire [0:0] csa_component57_fa32_xor1;
  wire [0:0] csa_component57_fa32_or0;
  wire [0:0] csa_component57_fa33_xor1;
  wire [0:0] csa_component57_fa33_or0;
  wire [0:0] csa_component57_fa34_xor1;
  wire [0:0] csa_component57_fa34_or0;
  wire [0:0] csa_component57_fa35_xor1;
  wire [0:0] csa_component57_fa35_or0;
  wire [0:0] csa_component57_fa36_xor1;
  wire [0:0] csa_component57_fa36_or0;
  wire [0:0] csa_component57_fa37_xor1;
  wire [0:0] csa_component57_fa37_or0;
  wire [0:0] csa_component57_fa38_xor1;
  wire [0:0] csa_component57_fa38_or0;
  wire [0:0] csa_component57_fa39_xor1;
  wire [0:0] csa_component57_fa39_or0;
  wire [0:0] csa_component57_fa40_xor1;
  wire [0:0] csa_component57_fa40_or0;
  wire [0:0] csa_component57_fa41_xor1;
  wire [0:0] csa_component57_fa41_or0;
  wire [0:0] csa_component57_fa42_xor1;
  wire [0:0] csa_component57_fa42_or0;
  wire [0:0] csa_component57_fa43_xor1;
  wire [0:0] csa_component57_fa43_or0;
  wire [0:0] csa_component57_fa44_xor1;
  wire [0:0] csa_component57_fa44_or0;
  wire [0:0] csa_component57_fa45_xor1;
  wire [0:0] csa_component57_fa45_or0;
  wire [0:0] csa_component57_fa46_xor1;
  wire [0:0] csa_component57_fa46_or0;
  wire [0:0] csa_component57_fa47_xor1;
  wire [0:0] csa_component57_fa47_or0;
  wire [0:0] csa_component57_fa48_xor1;
  wire [0:0] csa_component57_fa48_or0;
  wire [0:0] csa_component57_fa49_xor1;
  wire [0:0] csa_component57_fa49_or0;
  wire [0:0] csa_component57_fa50_xor1;
  wire [0:0] csa_component57_fa50_or0;
  wire [0:0] csa_component57_fa51_xor1;
  wire [0:0] csa_component57_fa51_or0;
  wire [0:0] csa_component57_fa52_xor1;
  wire [0:0] csa_component57_fa52_or0;
  wire [0:0] csa_component57_fa53_xor1;
  wire [0:0] csa_component57_fa53_or0;
  wire [0:0] csa_component57_fa54_xor1;
  wire [0:0] csa_component57_fa54_or0;
  wire [0:0] csa_component57_fa55_xor1;
  wire [0:0] csa_component57_fa55_or0;
  wire [0:0] csa_component57_fa56_xor1;
  wire [0:0] csa_component57_fa56_or0;

  fa fa_csa_component57_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component57_fa0_xor1), .fa_or0(csa_component57_fa0_or0));
  fa fa_csa_component57_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component57_fa1_xor1), .fa_or0(csa_component57_fa1_or0));
  fa fa_csa_component57_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component57_fa2_xor1), .fa_or0(csa_component57_fa2_or0));
  fa fa_csa_component57_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component57_fa3_xor1), .fa_or0(csa_component57_fa3_or0));
  fa fa_csa_component57_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component57_fa4_xor1), .fa_or0(csa_component57_fa4_or0));
  fa fa_csa_component57_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component57_fa5_xor1), .fa_or0(csa_component57_fa5_or0));
  fa fa_csa_component57_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component57_fa6_xor1), .fa_or0(csa_component57_fa6_or0));
  fa fa_csa_component57_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component57_fa7_xor1), .fa_or0(csa_component57_fa7_or0));
  fa fa_csa_component57_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component57_fa8_xor1), .fa_or0(csa_component57_fa8_or0));
  fa fa_csa_component57_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component57_fa9_xor1), .fa_or0(csa_component57_fa9_or0));
  fa fa_csa_component57_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component57_fa10_xor1), .fa_or0(csa_component57_fa10_or0));
  fa fa_csa_component57_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component57_fa11_xor1), .fa_or0(csa_component57_fa11_or0));
  fa fa_csa_component57_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component57_fa12_xor1), .fa_or0(csa_component57_fa12_or0));
  fa fa_csa_component57_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component57_fa13_xor1), .fa_or0(csa_component57_fa13_or0));
  fa fa_csa_component57_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component57_fa14_xor1), .fa_or0(csa_component57_fa14_or0));
  fa fa_csa_component57_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component57_fa15_xor1), .fa_or0(csa_component57_fa15_or0));
  fa fa_csa_component57_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component57_fa16_xor1), .fa_or0(csa_component57_fa16_or0));
  fa fa_csa_component57_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component57_fa17_xor1), .fa_or0(csa_component57_fa17_or0));
  fa fa_csa_component57_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component57_fa18_xor1), .fa_or0(csa_component57_fa18_or0));
  fa fa_csa_component57_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component57_fa19_xor1), .fa_or0(csa_component57_fa19_or0));
  fa fa_csa_component57_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component57_fa20_xor1), .fa_or0(csa_component57_fa20_or0));
  fa fa_csa_component57_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component57_fa21_xor1), .fa_or0(csa_component57_fa21_or0));
  fa fa_csa_component57_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component57_fa22_xor1), .fa_or0(csa_component57_fa22_or0));
  fa fa_csa_component57_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component57_fa23_xor1), .fa_or0(csa_component57_fa23_or0));
  fa fa_csa_component57_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component57_fa24_xor1), .fa_or0(csa_component57_fa24_or0));
  fa fa_csa_component57_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component57_fa25_xor1), .fa_or0(csa_component57_fa25_or0));
  fa fa_csa_component57_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component57_fa26_xor1), .fa_or0(csa_component57_fa26_or0));
  fa fa_csa_component57_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component57_fa27_xor1), .fa_or0(csa_component57_fa27_or0));
  fa fa_csa_component57_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component57_fa28_xor1), .fa_or0(csa_component57_fa28_or0));
  fa fa_csa_component57_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component57_fa29_xor1), .fa_or0(csa_component57_fa29_or0));
  fa fa_csa_component57_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component57_fa30_xor1), .fa_or0(csa_component57_fa30_or0));
  fa fa_csa_component57_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component57_fa31_xor1), .fa_or0(csa_component57_fa31_or0));
  fa fa_csa_component57_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component57_fa32_xor1), .fa_or0(csa_component57_fa32_or0));
  fa fa_csa_component57_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component57_fa33_xor1), .fa_or0(csa_component57_fa33_or0));
  fa fa_csa_component57_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component57_fa34_xor1), .fa_or0(csa_component57_fa34_or0));
  fa fa_csa_component57_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component57_fa35_xor1), .fa_or0(csa_component57_fa35_or0));
  fa fa_csa_component57_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component57_fa36_xor1), .fa_or0(csa_component57_fa36_or0));
  fa fa_csa_component57_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component57_fa37_xor1), .fa_or0(csa_component57_fa37_or0));
  fa fa_csa_component57_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component57_fa38_xor1), .fa_or0(csa_component57_fa38_or0));
  fa fa_csa_component57_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component57_fa39_xor1), .fa_or0(csa_component57_fa39_or0));
  fa fa_csa_component57_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component57_fa40_xor1), .fa_or0(csa_component57_fa40_or0));
  fa fa_csa_component57_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component57_fa41_xor1), .fa_or0(csa_component57_fa41_or0));
  fa fa_csa_component57_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component57_fa42_xor1), .fa_or0(csa_component57_fa42_or0));
  fa fa_csa_component57_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component57_fa43_xor1), .fa_or0(csa_component57_fa43_or0));
  fa fa_csa_component57_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component57_fa44_xor1), .fa_or0(csa_component57_fa44_or0));
  fa fa_csa_component57_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component57_fa45_xor1), .fa_or0(csa_component57_fa45_or0));
  fa fa_csa_component57_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component57_fa46_xor1), .fa_or0(csa_component57_fa46_or0));
  fa fa_csa_component57_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component57_fa47_xor1), .fa_or0(csa_component57_fa47_or0));
  fa fa_csa_component57_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component57_fa48_xor1), .fa_or0(csa_component57_fa48_or0));
  fa fa_csa_component57_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component57_fa49_xor1), .fa_or0(csa_component57_fa49_or0));
  fa fa_csa_component57_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component57_fa50_xor1), .fa_or0(csa_component57_fa50_or0));
  fa fa_csa_component57_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component57_fa51_xor1), .fa_or0(csa_component57_fa51_or0));
  fa fa_csa_component57_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component57_fa52_xor1), .fa_or0(csa_component57_fa52_or0));
  fa fa_csa_component57_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component57_fa53_xor1), .fa_or0(csa_component57_fa53_or0));
  fa fa_csa_component57_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component57_fa54_xor1), .fa_or0(csa_component57_fa54_or0));
  fa fa_csa_component57_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component57_fa55_xor1), .fa_or0(csa_component57_fa55_or0));
  fa fa_csa_component57_fa56_out(.a(a[56]), .b(b[56]), .cin(c[56]), .fa_xor1(csa_component57_fa56_xor1), .fa_or0(csa_component57_fa56_or0));

  assign csa_component57_out[0] = csa_component57_fa0_xor1[0];
  assign csa_component57_out[1] = csa_component57_fa1_xor1[0];
  assign csa_component57_out[2] = csa_component57_fa2_xor1[0];
  assign csa_component57_out[3] = csa_component57_fa3_xor1[0];
  assign csa_component57_out[4] = csa_component57_fa4_xor1[0];
  assign csa_component57_out[5] = csa_component57_fa5_xor1[0];
  assign csa_component57_out[6] = csa_component57_fa6_xor1[0];
  assign csa_component57_out[7] = csa_component57_fa7_xor1[0];
  assign csa_component57_out[8] = csa_component57_fa8_xor1[0];
  assign csa_component57_out[9] = csa_component57_fa9_xor1[0];
  assign csa_component57_out[10] = csa_component57_fa10_xor1[0];
  assign csa_component57_out[11] = csa_component57_fa11_xor1[0];
  assign csa_component57_out[12] = csa_component57_fa12_xor1[0];
  assign csa_component57_out[13] = csa_component57_fa13_xor1[0];
  assign csa_component57_out[14] = csa_component57_fa14_xor1[0];
  assign csa_component57_out[15] = csa_component57_fa15_xor1[0];
  assign csa_component57_out[16] = csa_component57_fa16_xor1[0];
  assign csa_component57_out[17] = csa_component57_fa17_xor1[0];
  assign csa_component57_out[18] = csa_component57_fa18_xor1[0];
  assign csa_component57_out[19] = csa_component57_fa19_xor1[0];
  assign csa_component57_out[20] = csa_component57_fa20_xor1[0];
  assign csa_component57_out[21] = csa_component57_fa21_xor1[0];
  assign csa_component57_out[22] = csa_component57_fa22_xor1[0];
  assign csa_component57_out[23] = csa_component57_fa23_xor1[0];
  assign csa_component57_out[24] = csa_component57_fa24_xor1[0];
  assign csa_component57_out[25] = csa_component57_fa25_xor1[0];
  assign csa_component57_out[26] = csa_component57_fa26_xor1[0];
  assign csa_component57_out[27] = csa_component57_fa27_xor1[0];
  assign csa_component57_out[28] = csa_component57_fa28_xor1[0];
  assign csa_component57_out[29] = csa_component57_fa29_xor1[0];
  assign csa_component57_out[30] = csa_component57_fa30_xor1[0];
  assign csa_component57_out[31] = csa_component57_fa31_xor1[0];
  assign csa_component57_out[32] = csa_component57_fa32_xor1[0];
  assign csa_component57_out[33] = csa_component57_fa33_xor1[0];
  assign csa_component57_out[34] = csa_component57_fa34_xor1[0];
  assign csa_component57_out[35] = csa_component57_fa35_xor1[0];
  assign csa_component57_out[36] = csa_component57_fa36_xor1[0];
  assign csa_component57_out[37] = csa_component57_fa37_xor1[0];
  assign csa_component57_out[38] = csa_component57_fa38_xor1[0];
  assign csa_component57_out[39] = csa_component57_fa39_xor1[0];
  assign csa_component57_out[40] = csa_component57_fa40_xor1[0];
  assign csa_component57_out[41] = csa_component57_fa41_xor1[0];
  assign csa_component57_out[42] = csa_component57_fa42_xor1[0];
  assign csa_component57_out[43] = csa_component57_fa43_xor1[0];
  assign csa_component57_out[44] = csa_component57_fa44_xor1[0];
  assign csa_component57_out[45] = csa_component57_fa45_xor1[0];
  assign csa_component57_out[46] = csa_component57_fa46_xor1[0];
  assign csa_component57_out[47] = csa_component57_fa47_xor1[0];
  assign csa_component57_out[48] = csa_component57_fa48_xor1[0];
  assign csa_component57_out[49] = csa_component57_fa49_xor1[0];
  assign csa_component57_out[50] = csa_component57_fa50_xor1[0];
  assign csa_component57_out[51] = csa_component57_fa51_xor1[0];
  assign csa_component57_out[52] = csa_component57_fa52_xor1[0];
  assign csa_component57_out[53] = csa_component57_fa53_xor1[0];
  assign csa_component57_out[54] = csa_component57_fa54_xor1[0];
  assign csa_component57_out[55] = csa_component57_fa55_xor1[0];
  assign csa_component57_out[56] = csa_component57_fa56_xor1[0];
  assign csa_component57_out[57] = 1'b0;
  assign csa_component57_out[58] = 1'b0;
  assign csa_component57_out[59] = csa_component57_fa0_or0[0];
  assign csa_component57_out[60] = csa_component57_fa1_or0[0];
  assign csa_component57_out[61] = csa_component57_fa2_or0[0];
  assign csa_component57_out[62] = csa_component57_fa3_or0[0];
  assign csa_component57_out[63] = csa_component57_fa4_or0[0];
  assign csa_component57_out[64] = csa_component57_fa5_or0[0];
  assign csa_component57_out[65] = csa_component57_fa6_or0[0];
  assign csa_component57_out[66] = csa_component57_fa7_or0[0];
  assign csa_component57_out[67] = csa_component57_fa8_or0[0];
  assign csa_component57_out[68] = csa_component57_fa9_or0[0];
  assign csa_component57_out[69] = csa_component57_fa10_or0[0];
  assign csa_component57_out[70] = csa_component57_fa11_or0[0];
  assign csa_component57_out[71] = csa_component57_fa12_or0[0];
  assign csa_component57_out[72] = csa_component57_fa13_or0[0];
  assign csa_component57_out[73] = csa_component57_fa14_or0[0];
  assign csa_component57_out[74] = csa_component57_fa15_or0[0];
  assign csa_component57_out[75] = csa_component57_fa16_or0[0];
  assign csa_component57_out[76] = csa_component57_fa17_or0[0];
  assign csa_component57_out[77] = csa_component57_fa18_or0[0];
  assign csa_component57_out[78] = csa_component57_fa19_or0[0];
  assign csa_component57_out[79] = csa_component57_fa20_or0[0];
  assign csa_component57_out[80] = csa_component57_fa21_or0[0];
  assign csa_component57_out[81] = csa_component57_fa22_or0[0];
  assign csa_component57_out[82] = csa_component57_fa23_or0[0];
  assign csa_component57_out[83] = csa_component57_fa24_or0[0];
  assign csa_component57_out[84] = csa_component57_fa25_or0[0];
  assign csa_component57_out[85] = csa_component57_fa26_or0[0];
  assign csa_component57_out[86] = csa_component57_fa27_or0[0];
  assign csa_component57_out[87] = csa_component57_fa28_or0[0];
  assign csa_component57_out[88] = csa_component57_fa29_or0[0];
  assign csa_component57_out[89] = csa_component57_fa30_or0[0];
  assign csa_component57_out[90] = csa_component57_fa31_or0[0];
  assign csa_component57_out[91] = csa_component57_fa32_or0[0];
  assign csa_component57_out[92] = csa_component57_fa33_or0[0];
  assign csa_component57_out[93] = csa_component57_fa34_or0[0];
  assign csa_component57_out[94] = csa_component57_fa35_or0[0];
  assign csa_component57_out[95] = csa_component57_fa36_or0[0];
  assign csa_component57_out[96] = csa_component57_fa37_or0[0];
  assign csa_component57_out[97] = csa_component57_fa38_or0[0];
  assign csa_component57_out[98] = csa_component57_fa39_or0[0];
  assign csa_component57_out[99] = csa_component57_fa40_or0[0];
  assign csa_component57_out[100] = csa_component57_fa41_or0[0];
  assign csa_component57_out[101] = csa_component57_fa42_or0[0];
  assign csa_component57_out[102] = csa_component57_fa43_or0[0];
  assign csa_component57_out[103] = csa_component57_fa44_or0[0];
  assign csa_component57_out[104] = csa_component57_fa45_or0[0];
  assign csa_component57_out[105] = csa_component57_fa46_or0[0];
  assign csa_component57_out[106] = csa_component57_fa47_or0[0];
  assign csa_component57_out[107] = csa_component57_fa48_or0[0];
  assign csa_component57_out[108] = csa_component57_fa49_or0[0];
  assign csa_component57_out[109] = csa_component57_fa50_or0[0];
  assign csa_component57_out[110] = csa_component57_fa51_or0[0];
  assign csa_component57_out[111] = csa_component57_fa52_or0[0];
  assign csa_component57_out[112] = csa_component57_fa53_or0[0];
  assign csa_component57_out[113] = csa_component57_fa54_or0[0];
  assign csa_component57_out[114] = csa_component57_fa55_or0[0];
  assign csa_component57_out[115] = csa_component57_fa56_or0[0];
endmodule

module csa_component60(input [59:0] a, input [59:0] b, input [59:0] c, output [121:0] csa_component60_out);
  wire [0:0] csa_component60_fa0_xor1;
  wire [0:0] csa_component60_fa0_or0;
  wire [0:0] csa_component60_fa1_xor1;
  wire [0:0] csa_component60_fa1_or0;
  wire [0:0] csa_component60_fa2_xor1;
  wire [0:0] csa_component60_fa2_or0;
  wire [0:0] csa_component60_fa3_xor1;
  wire [0:0] csa_component60_fa3_or0;
  wire [0:0] csa_component60_fa4_xor1;
  wire [0:0] csa_component60_fa4_or0;
  wire [0:0] csa_component60_fa5_xor1;
  wire [0:0] csa_component60_fa5_or0;
  wire [0:0] csa_component60_fa6_xor1;
  wire [0:0] csa_component60_fa6_or0;
  wire [0:0] csa_component60_fa7_xor1;
  wire [0:0] csa_component60_fa7_or0;
  wire [0:0] csa_component60_fa8_xor1;
  wire [0:0] csa_component60_fa8_or0;
  wire [0:0] csa_component60_fa9_xor1;
  wire [0:0] csa_component60_fa9_or0;
  wire [0:0] csa_component60_fa10_xor1;
  wire [0:0] csa_component60_fa10_or0;
  wire [0:0] csa_component60_fa11_xor1;
  wire [0:0] csa_component60_fa11_or0;
  wire [0:0] csa_component60_fa12_xor1;
  wire [0:0] csa_component60_fa12_or0;
  wire [0:0] csa_component60_fa13_xor1;
  wire [0:0] csa_component60_fa13_or0;
  wire [0:0] csa_component60_fa14_xor1;
  wire [0:0] csa_component60_fa14_or0;
  wire [0:0] csa_component60_fa15_xor1;
  wire [0:0] csa_component60_fa15_or0;
  wire [0:0] csa_component60_fa16_xor1;
  wire [0:0] csa_component60_fa16_or0;
  wire [0:0] csa_component60_fa17_xor1;
  wire [0:0] csa_component60_fa17_or0;
  wire [0:0] csa_component60_fa18_xor1;
  wire [0:0] csa_component60_fa18_or0;
  wire [0:0] csa_component60_fa19_xor1;
  wire [0:0] csa_component60_fa19_or0;
  wire [0:0] csa_component60_fa20_xor1;
  wire [0:0] csa_component60_fa20_or0;
  wire [0:0] csa_component60_fa21_xor1;
  wire [0:0] csa_component60_fa21_or0;
  wire [0:0] csa_component60_fa22_xor1;
  wire [0:0] csa_component60_fa22_or0;
  wire [0:0] csa_component60_fa23_xor1;
  wire [0:0] csa_component60_fa23_or0;
  wire [0:0] csa_component60_fa24_xor1;
  wire [0:0] csa_component60_fa24_or0;
  wire [0:0] csa_component60_fa25_xor1;
  wire [0:0] csa_component60_fa25_or0;
  wire [0:0] csa_component60_fa26_xor1;
  wire [0:0] csa_component60_fa26_or0;
  wire [0:0] csa_component60_fa27_xor1;
  wire [0:0] csa_component60_fa27_or0;
  wire [0:0] csa_component60_fa28_xor1;
  wire [0:0] csa_component60_fa28_or0;
  wire [0:0] csa_component60_fa29_xor1;
  wire [0:0] csa_component60_fa29_or0;
  wire [0:0] csa_component60_fa30_xor1;
  wire [0:0] csa_component60_fa30_or0;
  wire [0:0] csa_component60_fa31_xor1;
  wire [0:0] csa_component60_fa31_or0;
  wire [0:0] csa_component60_fa32_xor1;
  wire [0:0] csa_component60_fa32_or0;
  wire [0:0] csa_component60_fa33_xor1;
  wire [0:0] csa_component60_fa33_or0;
  wire [0:0] csa_component60_fa34_xor1;
  wire [0:0] csa_component60_fa34_or0;
  wire [0:0] csa_component60_fa35_xor1;
  wire [0:0] csa_component60_fa35_or0;
  wire [0:0] csa_component60_fa36_xor1;
  wire [0:0] csa_component60_fa36_or0;
  wire [0:0] csa_component60_fa37_xor1;
  wire [0:0] csa_component60_fa37_or0;
  wire [0:0] csa_component60_fa38_xor1;
  wire [0:0] csa_component60_fa38_or0;
  wire [0:0] csa_component60_fa39_xor1;
  wire [0:0] csa_component60_fa39_or0;
  wire [0:0] csa_component60_fa40_xor1;
  wire [0:0] csa_component60_fa40_or0;
  wire [0:0] csa_component60_fa41_xor1;
  wire [0:0] csa_component60_fa41_or0;
  wire [0:0] csa_component60_fa42_xor1;
  wire [0:0] csa_component60_fa42_or0;
  wire [0:0] csa_component60_fa43_xor1;
  wire [0:0] csa_component60_fa43_or0;
  wire [0:0] csa_component60_fa44_xor1;
  wire [0:0] csa_component60_fa44_or0;
  wire [0:0] csa_component60_fa45_xor1;
  wire [0:0] csa_component60_fa45_or0;
  wire [0:0] csa_component60_fa46_xor1;
  wire [0:0] csa_component60_fa46_or0;
  wire [0:0] csa_component60_fa47_xor1;
  wire [0:0] csa_component60_fa47_or0;
  wire [0:0] csa_component60_fa48_xor1;
  wire [0:0] csa_component60_fa48_or0;
  wire [0:0] csa_component60_fa49_xor1;
  wire [0:0] csa_component60_fa49_or0;
  wire [0:0] csa_component60_fa50_xor1;
  wire [0:0] csa_component60_fa50_or0;
  wire [0:0] csa_component60_fa51_xor1;
  wire [0:0] csa_component60_fa51_or0;
  wire [0:0] csa_component60_fa52_xor1;
  wire [0:0] csa_component60_fa52_or0;
  wire [0:0] csa_component60_fa53_xor1;
  wire [0:0] csa_component60_fa53_or0;
  wire [0:0] csa_component60_fa54_xor1;
  wire [0:0] csa_component60_fa54_or0;
  wire [0:0] csa_component60_fa55_xor1;
  wire [0:0] csa_component60_fa55_or0;
  wire [0:0] csa_component60_fa56_xor1;
  wire [0:0] csa_component60_fa56_or0;
  wire [0:0] csa_component60_fa57_xor1;
  wire [0:0] csa_component60_fa57_or0;
  wire [0:0] csa_component60_fa58_xor1;
  wire [0:0] csa_component60_fa58_or0;
  wire [0:0] csa_component60_fa59_xor1;
  wire [0:0] csa_component60_fa59_or0;

  fa fa_csa_component60_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component60_fa0_xor1), .fa_or0(csa_component60_fa0_or0));
  fa fa_csa_component60_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component60_fa1_xor1), .fa_or0(csa_component60_fa1_or0));
  fa fa_csa_component60_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component60_fa2_xor1), .fa_or0(csa_component60_fa2_or0));
  fa fa_csa_component60_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component60_fa3_xor1), .fa_or0(csa_component60_fa3_or0));
  fa fa_csa_component60_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component60_fa4_xor1), .fa_or0(csa_component60_fa4_or0));
  fa fa_csa_component60_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component60_fa5_xor1), .fa_or0(csa_component60_fa5_or0));
  fa fa_csa_component60_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component60_fa6_xor1), .fa_or0(csa_component60_fa6_or0));
  fa fa_csa_component60_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component60_fa7_xor1), .fa_or0(csa_component60_fa7_or0));
  fa fa_csa_component60_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component60_fa8_xor1), .fa_or0(csa_component60_fa8_or0));
  fa fa_csa_component60_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component60_fa9_xor1), .fa_or0(csa_component60_fa9_or0));
  fa fa_csa_component60_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component60_fa10_xor1), .fa_or0(csa_component60_fa10_or0));
  fa fa_csa_component60_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component60_fa11_xor1), .fa_or0(csa_component60_fa11_or0));
  fa fa_csa_component60_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component60_fa12_xor1), .fa_or0(csa_component60_fa12_or0));
  fa fa_csa_component60_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component60_fa13_xor1), .fa_or0(csa_component60_fa13_or0));
  fa fa_csa_component60_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component60_fa14_xor1), .fa_or0(csa_component60_fa14_or0));
  fa fa_csa_component60_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component60_fa15_xor1), .fa_or0(csa_component60_fa15_or0));
  fa fa_csa_component60_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component60_fa16_xor1), .fa_or0(csa_component60_fa16_or0));
  fa fa_csa_component60_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component60_fa17_xor1), .fa_or0(csa_component60_fa17_or0));
  fa fa_csa_component60_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component60_fa18_xor1), .fa_or0(csa_component60_fa18_or0));
  fa fa_csa_component60_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component60_fa19_xor1), .fa_or0(csa_component60_fa19_or0));
  fa fa_csa_component60_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component60_fa20_xor1), .fa_or0(csa_component60_fa20_or0));
  fa fa_csa_component60_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component60_fa21_xor1), .fa_or0(csa_component60_fa21_or0));
  fa fa_csa_component60_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component60_fa22_xor1), .fa_or0(csa_component60_fa22_or0));
  fa fa_csa_component60_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component60_fa23_xor1), .fa_or0(csa_component60_fa23_or0));
  fa fa_csa_component60_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component60_fa24_xor1), .fa_or0(csa_component60_fa24_or0));
  fa fa_csa_component60_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component60_fa25_xor1), .fa_or0(csa_component60_fa25_or0));
  fa fa_csa_component60_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component60_fa26_xor1), .fa_or0(csa_component60_fa26_or0));
  fa fa_csa_component60_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component60_fa27_xor1), .fa_or0(csa_component60_fa27_or0));
  fa fa_csa_component60_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component60_fa28_xor1), .fa_or0(csa_component60_fa28_or0));
  fa fa_csa_component60_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component60_fa29_xor1), .fa_or0(csa_component60_fa29_or0));
  fa fa_csa_component60_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component60_fa30_xor1), .fa_or0(csa_component60_fa30_or0));
  fa fa_csa_component60_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component60_fa31_xor1), .fa_or0(csa_component60_fa31_or0));
  fa fa_csa_component60_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component60_fa32_xor1), .fa_or0(csa_component60_fa32_or0));
  fa fa_csa_component60_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component60_fa33_xor1), .fa_or0(csa_component60_fa33_or0));
  fa fa_csa_component60_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component60_fa34_xor1), .fa_or0(csa_component60_fa34_or0));
  fa fa_csa_component60_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component60_fa35_xor1), .fa_or0(csa_component60_fa35_or0));
  fa fa_csa_component60_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component60_fa36_xor1), .fa_or0(csa_component60_fa36_or0));
  fa fa_csa_component60_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component60_fa37_xor1), .fa_or0(csa_component60_fa37_or0));
  fa fa_csa_component60_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component60_fa38_xor1), .fa_or0(csa_component60_fa38_or0));
  fa fa_csa_component60_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component60_fa39_xor1), .fa_or0(csa_component60_fa39_or0));
  fa fa_csa_component60_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component60_fa40_xor1), .fa_or0(csa_component60_fa40_or0));
  fa fa_csa_component60_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component60_fa41_xor1), .fa_or0(csa_component60_fa41_or0));
  fa fa_csa_component60_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component60_fa42_xor1), .fa_or0(csa_component60_fa42_or0));
  fa fa_csa_component60_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component60_fa43_xor1), .fa_or0(csa_component60_fa43_or0));
  fa fa_csa_component60_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component60_fa44_xor1), .fa_or0(csa_component60_fa44_or0));
  fa fa_csa_component60_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component60_fa45_xor1), .fa_or0(csa_component60_fa45_or0));
  fa fa_csa_component60_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component60_fa46_xor1), .fa_or0(csa_component60_fa46_or0));
  fa fa_csa_component60_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component60_fa47_xor1), .fa_or0(csa_component60_fa47_or0));
  fa fa_csa_component60_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component60_fa48_xor1), .fa_or0(csa_component60_fa48_or0));
  fa fa_csa_component60_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component60_fa49_xor1), .fa_or0(csa_component60_fa49_or0));
  fa fa_csa_component60_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component60_fa50_xor1), .fa_or0(csa_component60_fa50_or0));
  fa fa_csa_component60_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component60_fa51_xor1), .fa_or0(csa_component60_fa51_or0));
  fa fa_csa_component60_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component60_fa52_xor1), .fa_or0(csa_component60_fa52_or0));
  fa fa_csa_component60_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component60_fa53_xor1), .fa_or0(csa_component60_fa53_or0));
  fa fa_csa_component60_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component60_fa54_xor1), .fa_or0(csa_component60_fa54_or0));
  fa fa_csa_component60_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component60_fa55_xor1), .fa_or0(csa_component60_fa55_or0));
  fa fa_csa_component60_fa56_out(.a(a[56]), .b(b[56]), .cin(c[56]), .fa_xor1(csa_component60_fa56_xor1), .fa_or0(csa_component60_fa56_or0));
  fa fa_csa_component60_fa57_out(.a(a[57]), .b(b[57]), .cin(c[57]), .fa_xor1(csa_component60_fa57_xor1), .fa_or0(csa_component60_fa57_or0));
  fa fa_csa_component60_fa58_out(.a(a[58]), .b(b[58]), .cin(c[58]), .fa_xor1(csa_component60_fa58_xor1), .fa_or0(csa_component60_fa58_or0));
  fa fa_csa_component60_fa59_out(.a(a[59]), .b(b[59]), .cin(c[59]), .fa_xor1(csa_component60_fa59_xor1), .fa_or0(csa_component60_fa59_or0));

  assign csa_component60_out[0] = csa_component60_fa0_xor1[0];
  assign csa_component60_out[1] = csa_component60_fa1_xor1[0];
  assign csa_component60_out[2] = csa_component60_fa2_xor1[0];
  assign csa_component60_out[3] = csa_component60_fa3_xor1[0];
  assign csa_component60_out[4] = csa_component60_fa4_xor1[0];
  assign csa_component60_out[5] = csa_component60_fa5_xor1[0];
  assign csa_component60_out[6] = csa_component60_fa6_xor1[0];
  assign csa_component60_out[7] = csa_component60_fa7_xor1[0];
  assign csa_component60_out[8] = csa_component60_fa8_xor1[0];
  assign csa_component60_out[9] = csa_component60_fa9_xor1[0];
  assign csa_component60_out[10] = csa_component60_fa10_xor1[0];
  assign csa_component60_out[11] = csa_component60_fa11_xor1[0];
  assign csa_component60_out[12] = csa_component60_fa12_xor1[0];
  assign csa_component60_out[13] = csa_component60_fa13_xor1[0];
  assign csa_component60_out[14] = csa_component60_fa14_xor1[0];
  assign csa_component60_out[15] = csa_component60_fa15_xor1[0];
  assign csa_component60_out[16] = csa_component60_fa16_xor1[0];
  assign csa_component60_out[17] = csa_component60_fa17_xor1[0];
  assign csa_component60_out[18] = csa_component60_fa18_xor1[0];
  assign csa_component60_out[19] = csa_component60_fa19_xor1[0];
  assign csa_component60_out[20] = csa_component60_fa20_xor1[0];
  assign csa_component60_out[21] = csa_component60_fa21_xor1[0];
  assign csa_component60_out[22] = csa_component60_fa22_xor1[0];
  assign csa_component60_out[23] = csa_component60_fa23_xor1[0];
  assign csa_component60_out[24] = csa_component60_fa24_xor1[0];
  assign csa_component60_out[25] = csa_component60_fa25_xor1[0];
  assign csa_component60_out[26] = csa_component60_fa26_xor1[0];
  assign csa_component60_out[27] = csa_component60_fa27_xor1[0];
  assign csa_component60_out[28] = csa_component60_fa28_xor1[0];
  assign csa_component60_out[29] = csa_component60_fa29_xor1[0];
  assign csa_component60_out[30] = csa_component60_fa30_xor1[0];
  assign csa_component60_out[31] = csa_component60_fa31_xor1[0];
  assign csa_component60_out[32] = csa_component60_fa32_xor1[0];
  assign csa_component60_out[33] = csa_component60_fa33_xor1[0];
  assign csa_component60_out[34] = csa_component60_fa34_xor1[0];
  assign csa_component60_out[35] = csa_component60_fa35_xor1[0];
  assign csa_component60_out[36] = csa_component60_fa36_xor1[0];
  assign csa_component60_out[37] = csa_component60_fa37_xor1[0];
  assign csa_component60_out[38] = csa_component60_fa38_xor1[0];
  assign csa_component60_out[39] = csa_component60_fa39_xor1[0];
  assign csa_component60_out[40] = csa_component60_fa40_xor1[0];
  assign csa_component60_out[41] = csa_component60_fa41_xor1[0];
  assign csa_component60_out[42] = csa_component60_fa42_xor1[0];
  assign csa_component60_out[43] = csa_component60_fa43_xor1[0];
  assign csa_component60_out[44] = csa_component60_fa44_xor1[0];
  assign csa_component60_out[45] = csa_component60_fa45_xor1[0];
  assign csa_component60_out[46] = csa_component60_fa46_xor1[0];
  assign csa_component60_out[47] = csa_component60_fa47_xor1[0];
  assign csa_component60_out[48] = csa_component60_fa48_xor1[0];
  assign csa_component60_out[49] = csa_component60_fa49_xor1[0];
  assign csa_component60_out[50] = csa_component60_fa50_xor1[0];
  assign csa_component60_out[51] = csa_component60_fa51_xor1[0];
  assign csa_component60_out[52] = csa_component60_fa52_xor1[0];
  assign csa_component60_out[53] = csa_component60_fa53_xor1[0];
  assign csa_component60_out[54] = csa_component60_fa54_xor1[0];
  assign csa_component60_out[55] = csa_component60_fa55_xor1[0];
  assign csa_component60_out[56] = csa_component60_fa56_xor1[0];
  assign csa_component60_out[57] = csa_component60_fa57_xor1[0];
  assign csa_component60_out[58] = csa_component60_fa58_xor1[0];
  assign csa_component60_out[59] = csa_component60_fa59_xor1[0];
  assign csa_component60_out[60] = 1'b0;
  assign csa_component60_out[61] = 1'b0;
  assign csa_component60_out[62] = csa_component60_fa0_or0[0];
  assign csa_component60_out[63] = csa_component60_fa1_or0[0];
  assign csa_component60_out[64] = csa_component60_fa2_or0[0];
  assign csa_component60_out[65] = csa_component60_fa3_or0[0];
  assign csa_component60_out[66] = csa_component60_fa4_or0[0];
  assign csa_component60_out[67] = csa_component60_fa5_or0[0];
  assign csa_component60_out[68] = csa_component60_fa6_or0[0];
  assign csa_component60_out[69] = csa_component60_fa7_or0[0];
  assign csa_component60_out[70] = csa_component60_fa8_or0[0];
  assign csa_component60_out[71] = csa_component60_fa9_or0[0];
  assign csa_component60_out[72] = csa_component60_fa10_or0[0];
  assign csa_component60_out[73] = csa_component60_fa11_or0[0];
  assign csa_component60_out[74] = csa_component60_fa12_or0[0];
  assign csa_component60_out[75] = csa_component60_fa13_or0[0];
  assign csa_component60_out[76] = csa_component60_fa14_or0[0];
  assign csa_component60_out[77] = csa_component60_fa15_or0[0];
  assign csa_component60_out[78] = csa_component60_fa16_or0[0];
  assign csa_component60_out[79] = csa_component60_fa17_or0[0];
  assign csa_component60_out[80] = csa_component60_fa18_or0[0];
  assign csa_component60_out[81] = csa_component60_fa19_or0[0];
  assign csa_component60_out[82] = csa_component60_fa20_or0[0];
  assign csa_component60_out[83] = csa_component60_fa21_or0[0];
  assign csa_component60_out[84] = csa_component60_fa22_or0[0];
  assign csa_component60_out[85] = csa_component60_fa23_or0[0];
  assign csa_component60_out[86] = csa_component60_fa24_or0[0];
  assign csa_component60_out[87] = csa_component60_fa25_or0[0];
  assign csa_component60_out[88] = csa_component60_fa26_or0[0];
  assign csa_component60_out[89] = csa_component60_fa27_or0[0];
  assign csa_component60_out[90] = csa_component60_fa28_or0[0];
  assign csa_component60_out[91] = csa_component60_fa29_or0[0];
  assign csa_component60_out[92] = csa_component60_fa30_or0[0];
  assign csa_component60_out[93] = csa_component60_fa31_or0[0];
  assign csa_component60_out[94] = csa_component60_fa32_or0[0];
  assign csa_component60_out[95] = csa_component60_fa33_or0[0];
  assign csa_component60_out[96] = csa_component60_fa34_or0[0];
  assign csa_component60_out[97] = csa_component60_fa35_or0[0];
  assign csa_component60_out[98] = csa_component60_fa36_or0[0];
  assign csa_component60_out[99] = csa_component60_fa37_or0[0];
  assign csa_component60_out[100] = csa_component60_fa38_or0[0];
  assign csa_component60_out[101] = csa_component60_fa39_or0[0];
  assign csa_component60_out[102] = csa_component60_fa40_or0[0];
  assign csa_component60_out[103] = csa_component60_fa41_or0[0];
  assign csa_component60_out[104] = csa_component60_fa42_or0[0];
  assign csa_component60_out[105] = csa_component60_fa43_or0[0];
  assign csa_component60_out[106] = csa_component60_fa44_or0[0];
  assign csa_component60_out[107] = csa_component60_fa45_or0[0];
  assign csa_component60_out[108] = csa_component60_fa46_or0[0];
  assign csa_component60_out[109] = csa_component60_fa47_or0[0];
  assign csa_component60_out[110] = csa_component60_fa48_or0[0];
  assign csa_component60_out[111] = csa_component60_fa49_or0[0];
  assign csa_component60_out[112] = csa_component60_fa50_or0[0];
  assign csa_component60_out[113] = csa_component60_fa51_or0[0];
  assign csa_component60_out[114] = csa_component60_fa52_or0[0];
  assign csa_component60_out[115] = csa_component60_fa53_or0[0];
  assign csa_component60_out[116] = csa_component60_fa54_or0[0];
  assign csa_component60_out[117] = csa_component60_fa55_or0[0];
  assign csa_component60_out[118] = csa_component60_fa56_or0[0];
  assign csa_component60_out[119] = csa_component60_fa57_or0[0];
  assign csa_component60_out[120] = csa_component60_fa58_or0[0];
  assign csa_component60_out[121] = csa_component60_fa59_or0[0];
endmodule

module csa_component63(input [62:0] a, input [62:0] b, input [62:0] c, output [127:0] csa_component63_out);
  wire [0:0] csa_component63_fa0_xor1;
  wire [0:0] csa_component63_fa0_or0;
  wire [0:0] csa_component63_fa1_xor1;
  wire [0:0] csa_component63_fa1_or0;
  wire [0:0] csa_component63_fa2_xor1;
  wire [0:0] csa_component63_fa2_or0;
  wire [0:0] csa_component63_fa3_xor1;
  wire [0:0] csa_component63_fa3_or0;
  wire [0:0] csa_component63_fa4_xor1;
  wire [0:0] csa_component63_fa4_or0;
  wire [0:0] csa_component63_fa5_xor1;
  wire [0:0] csa_component63_fa5_or0;
  wire [0:0] csa_component63_fa6_xor1;
  wire [0:0] csa_component63_fa6_or0;
  wire [0:0] csa_component63_fa7_xor1;
  wire [0:0] csa_component63_fa7_or0;
  wire [0:0] csa_component63_fa8_xor1;
  wire [0:0] csa_component63_fa8_or0;
  wire [0:0] csa_component63_fa9_xor1;
  wire [0:0] csa_component63_fa9_or0;
  wire [0:0] csa_component63_fa10_xor1;
  wire [0:0] csa_component63_fa10_or0;
  wire [0:0] csa_component63_fa11_xor1;
  wire [0:0] csa_component63_fa11_or0;
  wire [0:0] csa_component63_fa12_xor1;
  wire [0:0] csa_component63_fa12_or0;
  wire [0:0] csa_component63_fa13_xor1;
  wire [0:0] csa_component63_fa13_or0;
  wire [0:0] csa_component63_fa14_xor1;
  wire [0:0] csa_component63_fa14_or0;
  wire [0:0] csa_component63_fa15_xor1;
  wire [0:0] csa_component63_fa15_or0;
  wire [0:0] csa_component63_fa16_xor1;
  wire [0:0] csa_component63_fa16_or0;
  wire [0:0] csa_component63_fa17_xor1;
  wire [0:0] csa_component63_fa17_or0;
  wire [0:0] csa_component63_fa18_xor1;
  wire [0:0] csa_component63_fa18_or0;
  wire [0:0] csa_component63_fa19_xor1;
  wire [0:0] csa_component63_fa19_or0;
  wire [0:0] csa_component63_fa20_xor1;
  wire [0:0] csa_component63_fa20_or0;
  wire [0:0] csa_component63_fa21_xor1;
  wire [0:0] csa_component63_fa21_or0;
  wire [0:0] csa_component63_fa22_xor1;
  wire [0:0] csa_component63_fa22_or0;
  wire [0:0] csa_component63_fa23_xor1;
  wire [0:0] csa_component63_fa23_or0;
  wire [0:0] csa_component63_fa24_xor1;
  wire [0:0] csa_component63_fa24_or0;
  wire [0:0] csa_component63_fa25_xor1;
  wire [0:0] csa_component63_fa25_or0;
  wire [0:0] csa_component63_fa26_xor1;
  wire [0:0] csa_component63_fa26_or0;
  wire [0:0] csa_component63_fa27_xor1;
  wire [0:0] csa_component63_fa27_or0;
  wire [0:0] csa_component63_fa28_xor1;
  wire [0:0] csa_component63_fa28_or0;
  wire [0:0] csa_component63_fa29_xor1;
  wire [0:0] csa_component63_fa29_or0;
  wire [0:0] csa_component63_fa30_xor1;
  wire [0:0] csa_component63_fa30_or0;
  wire [0:0] csa_component63_fa31_xor1;
  wire [0:0] csa_component63_fa31_or0;
  wire [0:0] csa_component63_fa32_xor1;
  wire [0:0] csa_component63_fa32_or0;
  wire [0:0] csa_component63_fa33_xor1;
  wire [0:0] csa_component63_fa33_or0;
  wire [0:0] csa_component63_fa34_xor1;
  wire [0:0] csa_component63_fa34_or0;
  wire [0:0] csa_component63_fa35_xor1;
  wire [0:0] csa_component63_fa35_or0;
  wire [0:0] csa_component63_fa36_xor1;
  wire [0:0] csa_component63_fa36_or0;
  wire [0:0] csa_component63_fa37_xor1;
  wire [0:0] csa_component63_fa37_or0;
  wire [0:0] csa_component63_fa38_xor1;
  wire [0:0] csa_component63_fa38_or0;
  wire [0:0] csa_component63_fa39_xor1;
  wire [0:0] csa_component63_fa39_or0;
  wire [0:0] csa_component63_fa40_xor1;
  wire [0:0] csa_component63_fa40_or0;
  wire [0:0] csa_component63_fa41_xor1;
  wire [0:0] csa_component63_fa41_or0;
  wire [0:0] csa_component63_fa42_xor1;
  wire [0:0] csa_component63_fa42_or0;
  wire [0:0] csa_component63_fa43_xor1;
  wire [0:0] csa_component63_fa43_or0;
  wire [0:0] csa_component63_fa44_xor1;
  wire [0:0] csa_component63_fa44_or0;
  wire [0:0] csa_component63_fa45_xor1;
  wire [0:0] csa_component63_fa45_or0;
  wire [0:0] csa_component63_fa46_xor1;
  wire [0:0] csa_component63_fa46_or0;
  wire [0:0] csa_component63_fa47_xor1;
  wire [0:0] csa_component63_fa47_or0;
  wire [0:0] csa_component63_fa48_xor1;
  wire [0:0] csa_component63_fa48_or0;
  wire [0:0] csa_component63_fa49_xor1;
  wire [0:0] csa_component63_fa49_or0;
  wire [0:0] csa_component63_fa50_xor1;
  wire [0:0] csa_component63_fa50_or0;
  wire [0:0] csa_component63_fa51_xor1;
  wire [0:0] csa_component63_fa51_or0;
  wire [0:0] csa_component63_fa52_xor1;
  wire [0:0] csa_component63_fa52_or0;
  wire [0:0] csa_component63_fa53_xor1;
  wire [0:0] csa_component63_fa53_or0;
  wire [0:0] csa_component63_fa54_xor1;
  wire [0:0] csa_component63_fa54_or0;
  wire [0:0] csa_component63_fa55_xor1;
  wire [0:0] csa_component63_fa55_or0;
  wire [0:0] csa_component63_fa56_xor1;
  wire [0:0] csa_component63_fa56_or0;
  wire [0:0] csa_component63_fa57_xor1;
  wire [0:0] csa_component63_fa57_or0;
  wire [0:0] csa_component63_fa58_xor1;
  wire [0:0] csa_component63_fa58_or0;
  wire [0:0] csa_component63_fa59_xor1;
  wire [0:0] csa_component63_fa59_or0;
  wire [0:0] csa_component63_fa60_xor1;
  wire [0:0] csa_component63_fa60_or0;
  wire [0:0] csa_component63_fa61_xor1;
  wire [0:0] csa_component63_fa61_or0;
  wire [0:0] csa_component63_fa62_xor1;
  wire [0:0] csa_component63_fa62_or0;

  fa fa_csa_component63_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component63_fa0_xor1), .fa_or0(csa_component63_fa0_or0));
  fa fa_csa_component63_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component63_fa1_xor1), .fa_or0(csa_component63_fa1_or0));
  fa fa_csa_component63_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component63_fa2_xor1), .fa_or0(csa_component63_fa2_or0));
  fa fa_csa_component63_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component63_fa3_xor1), .fa_or0(csa_component63_fa3_or0));
  fa fa_csa_component63_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component63_fa4_xor1), .fa_or0(csa_component63_fa4_or0));
  fa fa_csa_component63_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component63_fa5_xor1), .fa_or0(csa_component63_fa5_or0));
  fa fa_csa_component63_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component63_fa6_xor1), .fa_or0(csa_component63_fa6_or0));
  fa fa_csa_component63_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component63_fa7_xor1), .fa_or0(csa_component63_fa7_or0));
  fa fa_csa_component63_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component63_fa8_xor1), .fa_or0(csa_component63_fa8_or0));
  fa fa_csa_component63_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component63_fa9_xor1), .fa_or0(csa_component63_fa9_or0));
  fa fa_csa_component63_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component63_fa10_xor1), .fa_or0(csa_component63_fa10_or0));
  fa fa_csa_component63_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component63_fa11_xor1), .fa_or0(csa_component63_fa11_or0));
  fa fa_csa_component63_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component63_fa12_xor1), .fa_or0(csa_component63_fa12_or0));
  fa fa_csa_component63_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component63_fa13_xor1), .fa_or0(csa_component63_fa13_or0));
  fa fa_csa_component63_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component63_fa14_xor1), .fa_or0(csa_component63_fa14_or0));
  fa fa_csa_component63_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component63_fa15_xor1), .fa_or0(csa_component63_fa15_or0));
  fa fa_csa_component63_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component63_fa16_xor1), .fa_or0(csa_component63_fa16_or0));
  fa fa_csa_component63_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component63_fa17_xor1), .fa_or0(csa_component63_fa17_or0));
  fa fa_csa_component63_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component63_fa18_xor1), .fa_or0(csa_component63_fa18_or0));
  fa fa_csa_component63_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component63_fa19_xor1), .fa_or0(csa_component63_fa19_or0));
  fa fa_csa_component63_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component63_fa20_xor1), .fa_or0(csa_component63_fa20_or0));
  fa fa_csa_component63_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component63_fa21_xor1), .fa_or0(csa_component63_fa21_or0));
  fa fa_csa_component63_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component63_fa22_xor1), .fa_or0(csa_component63_fa22_or0));
  fa fa_csa_component63_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component63_fa23_xor1), .fa_or0(csa_component63_fa23_or0));
  fa fa_csa_component63_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component63_fa24_xor1), .fa_or0(csa_component63_fa24_or0));
  fa fa_csa_component63_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component63_fa25_xor1), .fa_or0(csa_component63_fa25_or0));
  fa fa_csa_component63_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component63_fa26_xor1), .fa_or0(csa_component63_fa26_or0));
  fa fa_csa_component63_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component63_fa27_xor1), .fa_or0(csa_component63_fa27_or0));
  fa fa_csa_component63_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component63_fa28_xor1), .fa_or0(csa_component63_fa28_or0));
  fa fa_csa_component63_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component63_fa29_xor1), .fa_or0(csa_component63_fa29_or0));
  fa fa_csa_component63_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component63_fa30_xor1), .fa_or0(csa_component63_fa30_or0));
  fa fa_csa_component63_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component63_fa31_xor1), .fa_or0(csa_component63_fa31_or0));
  fa fa_csa_component63_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component63_fa32_xor1), .fa_or0(csa_component63_fa32_or0));
  fa fa_csa_component63_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component63_fa33_xor1), .fa_or0(csa_component63_fa33_or0));
  fa fa_csa_component63_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component63_fa34_xor1), .fa_or0(csa_component63_fa34_or0));
  fa fa_csa_component63_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component63_fa35_xor1), .fa_or0(csa_component63_fa35_or0));
  fa fa_csa_component63_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component63_fa36_xor1), .fa_or0(csa_component63_fa36_or0));
  fa fa_csa_component63_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component63_fa37_xor1), .fa_or0(csa_component63_fa37_or0));
  fa fa_csa_component63_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component63_fa38_xor1), .fa_or0(csa_component63_fa38_or0));
  fa fa_csa_component63_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component63_fa39_xor1), .fa_or0(csa_component63_fa39_or0));
  fa fa_csa_component63_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component63_fa40_xor1), .fa_or0(csa_component63_fa40_or0));
  fa fa_csa_component63_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component63_fa41_xor1), .fa_or0(csa_component63_fa41_or0));
  fa fa_csa_component63_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component63_fa42_xor1), .fa_or0(csa_component63_fa42_or0));
  fa fa_csa_component63_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component63_fa43_xor1), .fa_or0(csa_component63_fa43_or0));
  fa fa_csa_component63_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component63_fa44_xor1), .fa_or0(csa_component63_fa44_or0));
  fa fa_csa_component63_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component63_fa45_xor1), .fa_or0(csa_component63_fa45_or0));
  fa fa_csa_component63_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component63_fa46_xor1), .fa_or0(csa_component63_fa46_or0));
  fa fa_csa_component63_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component63_fa47_xor1), .fa_or0(csa_component63_fa47_or0));
  fa fa_csa_component63_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component63_fa48_xor1), .fa_or0(csa_component63_fa48_or0));
  fa fa_csa_component63_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component63_fa49_xor1), .fa_or0(csa_component63_fa49_or0));
  fa fa_csa_component63_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component63_fa50_xor1), .fa_or0(csa_component63_fa50_or0));
  fa fa_csa_component63_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component63_fa51_xor1), .fa_or0(csa_component63_fa51_or0));
  fa fa_csa_component63_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component63_fa52_xor1), .fa_or0(csa_component63_fa52_or0));
  fa fa_csa_component63_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component63_fa53_xor1), .fa_or0(csa_component63_fa53_or0));
  fa fa_csa_component63_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component63_fa54_xor1), .fa_or0(csa_component63_fa54_or0));
  fa fa_csa_component63_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component63_fa55_xor1), .fa_or0(csa_component63_fa55_or0));
  fa fa_csa_component63_fa56_out(.a(a[56]), .b(b[56]), .cin(c[56]), .fa_xor1(csa_component63_fa56_xor1), .fa_or0(csa_component63_fa56_or0));
  fa fa_csa_component63_fa57_out(.a(a[57]), .b(b[57]), .cin(c[57]), .fa_xor1(csa_component63_fa57_xor1), .fa_or0(csa_component63_fa57_or0));
  fa fa_csa_component63_fa58_out(.a(a[58]), .b(b[58]), .cin(c[58]), .fa_xor1(csa_component63_fa58_xor1), .fa_or0(csa_component63_fa58_or0));
  fa fa_csa_component63_fa59_out(.a(a[59]), .b(b[59]), .cin(c[59]), .fa_xor1(csa_component63_fa59_xor1), .fa_or0(csa_component63_fa59_or0));
  fa fa_csa_component63_fa60_out(.a(a[60]), .b(b[60]), .cin(c[60]), .fa_xor1(csa_component63_fa60_xor1), .fa_or0(csa_component63_fa60_or0));
  fa fa_csa_component63_fa61_out(.a(a[61]), .b(b[61]), .cin(c[61]), .fa_xor1(csa_component63_fa61_xor1), .fa_or0(csa_component63_fa61_or0));
  fa fa_csa_component63_fa62_out(.a(a[62]), .b(b[62]), .cin(c[62]), .fa_xor1(csa_component63_fa62_xor1), .fa_or0(csa_component63_fa62_or0));

  assign csa_component63_out[0] = csa_component63_fa0_xor1[0];
  assign csa_component63_out[1] = csa_component63_fa1_xor1[0];
  assign csa_component63_out[2] = csa_component63_fa2_xor1[0];
  assign csa_component63_out[3] = csa_component63_fa3_xor1[0];
  assign csa_component63_out[4] = csa_component63_fa4_xor1[0];
  assign csa_component63_out[5] = csa_component63_fa5_xor1[0];
  assign csa_component63_out[6] = csa_component63_fa6_xor1[0];
  assign csa_component63_out[7] = csa_component63_fa7_xor1[0];
  assign csa_component63_out[8] = csa_component63_fa8_xor1[0];
  assign csa_component63_out[9] = csa_component63_fa9_xor1[0];
  assign csa_component63_out[10] = csa_component63_fa10_xor1[0];
  assign csa_component63_out[11] = csa_component63_fa11_xor1[0];
  assign csa_component63_out[12] = csa_component63_fa12_xor1[0];
  assign csa_component63_out[13] = csa_component63_fa13_xor1[0];
  assign csa_component63_out[14] = csa_component63_fa14_xor1[0];
  assign csa_component63_out[15] = csa_component63_fa15_xor1[0];
  assign csa_component63_out[16] = csa_component63_fa16_xor1[0];
  assign csa_component63_out[17] = csa_component63_fa17_xor1[0];
  assign csa_component63_out[18] = csa_component63_fa18_xor1[0];
  assign csa_component63_out[19] = csa_component63_fa19_xor1[0];
  assign csa_component63_out[20] = csa_component63_fa20_xor1[0];
  assign csa_component63_out[21] = csa_component63_fa21_xor1[0];
  assign csa_component63_out[22] = csa_component63_fa22_xor1[0];
  assign csa_component63_out[23] = csa_component63_fa23_xor1[0];
  assign csa_component63_out[24] = csa_component63_fa24_xor1[0];
  assign csa_component63_out[25] = csa_component63_fa25_xor1[0];
  assign csa_component63_out[26] = csa_component63_fa26_xor1[0];
  assign csa_component63_out[27] = csa_component63_fa27_xor1[0];
  assign csa_component63_out[28] = csa_component63_fa28_xor1[0];
  assign csa_component63_out[29] = csa_component63_fa29_xor1[0];
  assign csa_component63_out[30] = csa_component63_fa30_xor1[0];
  assign csa_component63_out[31] = csa_component63_fa31_xor1[0];
  assign csa_component63_out[32] = csa_component63_fa32_xor1[0];
  assign csa_component63_out[33] = csa_component63_fa33_xor1[0];
  assign csa_component63_out[34] = csa_component63_fa34_xor1[0];
  assign csa_component63_out[35] = csa_component63_fa35_xor1[0];
  assign csa_component63_out[36] = csa_component63_fa36_xor1[0];
  assign csa_component63_out[37] = csa_component63_fa37_xor1[0];
  assign csa_component63_out[38] = csa_component63_fa38_xor1[0];
  assign csa_component63_out[39] = csa_component63_fa39_xor1[0];
  assign csa_component63_out[40] = csa_component63_fa40_xor1[0];
  assign csa_component63_out[41] = csa_component63_fa41_xor1[0];
  assign csa_component63_out[42] = csa_component63_fa42_xor1[0];
  assign csa_component63_out[43] = csa_component63_fa43_xor1[0];
  assign csa_component63_out[44] = csa_component63_fa44_xor1[0];
  assign csa_component63_out[45] = csa_component63_fa45_xor1[0];
  assign csa_component63_out[46] = csa_component63_fa46_xor1[0];
  assign csa_component63_out[47] = csa_component63_fa47_xor1[0];
  assign csa_component63_out[48] = csa_component63_fa48_xor1[0];
  assign csa_component63_out[49] = csa_component63_fa49_xor1[0];
  assign csa_component63_out[50] = csa_component63_fa50_xor1[0];
  assign csa_component63_out[51] = csa_component63_fa51_xor1[0];
  assign csa_component63_out[52] = csa_component63_fa52_xor1[0];
  assign csa_component63_out[53] = csa_component63_fa53_xor1[0];
  assign csa_component63_out[54] = csa_component63_fa54_xor1[0];
  assign csa_component63_out[55] = csa_component63_fa55_xor1[0];
  assign csa_component63_out[56] = csa_component63_fa56_xor1[0];
  assign csa_component63_out[57] = csa_component63_fa57_xor1[0];
  assign csa_component63_out[58] = csa_component63_fa58_xor1[0];
  assign csa_component63_out[59] = csa_component63_fa59_xor1[0];
  assign csa_component63_out[60] = csa_component63_fa60_xor1[0];
  assign csa_component63_out[61] = csa_component63_fa61_xor1[0];
  assign csa_component63_out[62] = csa_component63_fa62_xor1[0];
  assign csa_component63_out[63] = 1'b0;
  assign csa_component63_out[64] = 1'b0;
  assign csa_component63_out[65] = csa_component63_fa0_or0[0];
  assign csa_component63_out[66] = csa_component63_fa1_or0[0];
  assign csa_component63_out[67] = csa_component63_fa2_or0[0];
  assign csa_component63_out[68] = csa_component63_fa3_or0[0];
  assign csa_component63_out[69] = csa_component63_fa4_or0[0];
  assign csa_component63_out[70] = csa_component63_fa5_or0[0];
  assign csa_component63_out[71] = csa_component63_fa6_or0[0];
  assign csa_component63_out[72] = csa_component63_fa7_or0[0];
  assign csa_component63_out[73] = csa_component63_fa8_or0[0];
  assign csa_component63_out[74] = csa_component63_fa9_or0[0];
  assign csa_component63_out[75] = csa_component63_fa10_or0[0];
  assign csa_component63_out[76] = csa_component63_fa11_or0[0];
  assign csa_component63_out[77] = csa_component63_fa12_or0[0];
  assign csa_component63_out[78] = csa_component63_fa13_or0[0];
  assign csa_component63_out[79] = csa_component63_fa14_or0[0];
  assign csa_component63_out[80] = csa_component63_fa15_or0[0];
  assign csa_component63_out[81] = csa_component63_fa16_or0[0];
  assign csa_component63_out[82] = csa_component63_fa17_or0[0];
  assign csa_component63_out[83] = csa_component63_fa18_or0[0];
  assign csa_component63_out[84] = csa_component63_fa19_or0[0];
  assign csa_component63_out[85] = csa_component63_fa20_or0[0];
  assign csa_component63_out[86] = csa_component63_fa21_or0[0];
  assign csa_component63_out[87] = csa_component63_fa22_or0[0];
  assign csa_component63_out[88] = csa_component63_fa23_or0[0];
  assign csa_component63_out[89] = csa_component63_fa24_or0[0];
  assign csa_component63_out[90] = csa_component63_fa25_or0[0];
  assign csa_component63_out[91] = csa_component63_fa26_or0[0];
  assign csa_component63_out[92] = csa_component63_fa27_or0[0];
  assign csa_component63_out[93] = csa_component63_fa28_or0[0];
  assign csa_component63_out[94] = csa_component63_fa29_or0[0];
  assign csa_component63_out[95] = csa_component63_fa30_or0[0];
  assign csa_component63_out[96] = csa_component63_fa31_or0[0];
  assign csa_component63_out[97] = csa_component63_fa32_or0[0];
  assign csa_component63_out[98] = csa_component63_fa33_or0[0];
  assign csa_component63_out[99] = csa_component63_fa34_or0[0];
  assign csa_component63_out[100] = csa_component63_fa35_or0[0];
  assign csa_component63_out[101] = csa_component63_fa36_or0[0];
  assign csa_component63_out[102] = csa_component63_fa37_or0[0];
  assign csa_component63_out[103] = csa_component63_fa38_or0[0];
  assign csa_component63_out[104] = csa_component63_fa39_or0[0];
  assign csa_component63_out[105] = csa_component63_fa40_or0[0];
  assign csa_component63_out[106] = csa_component63_fa41_or0[0];
  assign csa_component63_out[107] = csa_component63_fa42_or0[0];
  assign csa_component63_out[108] = csa_component63_fa43_or0[0];
  assign csa_component63_out[109] = csa_component63_fa44_or0[0];
  assign csa_component63_out[110] = csa_component63_fa45_or0[0];
  assign csa_component63_out[111] = csa_component63_fa46_or0[0];
  assign csa_component63_out[112] = csa_component63_fa47_or0[0];
  assign csa_component63_out[113] = csa_component63_fa48_or0[0];
  assign csa_component63_out[114] = csa_component63_fa49_or0[0];
  assign csa_component63_out[115] = csa_component63_fa50_or0[0];
  assign csa_component63_out[116] = csa_component63_fa51_or0[0];
  assign csa_component63_out[117] = csa_component63_fa52_or0[0];
  assign csa_component63_out[118] = csa_component63_fa53_or0[0];
  assign csa_component63_out[119] = csa_component63_fa54_or0[0];
  assign csa_component63_out[120] = csa_component63_fa55_or0[0];
  assign csa_component63_out[121] = csa_component63_fa56_or0[0];
  assign csa_component63_out[122] = csa_component63_fa57_or0[0];
  assign csa_component63_out[123] = csa_component63_fa58_or0[0];
  assign csa_component63_out[124] = csa_component63_fa59_or0[0];
  assign csa_component63_out[125] = csa_component63_fa60_or0[0];
  assign csa_component63_out[126] = csa_component63_fa61_or0[0];
  assign csa_component63_out[127] = csa_component63_fa62_or0[0];
endmodule

module csa_component64(input [63:0] a, input [63:0] b, input [63:0] c, output [129:0] csa_component64_out);
  wire [0:0] csa_component64_fa0_xor1;
  wire [0:0] csa_component64_fa0_or0;
  wire [0:0] csa_component64_fa1_xor1;
  wire [0:0] csa_component64_fa1_or0;
  wire [0:0] csa_component64_fa2_xor1;
  wire [0:0] csa_component64_fa2_or0;
  wire [0:0] csa_component64_fa3_xor1;
  wire [0:0] csa_component64_fa3_or0;
  wire [0:0] csa_component64_fa4_xor1;
  wire [0:0] csa_component64_fa4_or0;
  wire [0:0] csa_component64_fa5_xor1;
  wire [0:0] csa_component64_fa5_or0;
  wire [0:0] csa_component64_fa6_xor1;
  wire [0:0] csa_component64_fa6_or0;
  wire [0:0] csa_component64_fa7_xor1;
  wire [0:0] csa_component64_fa7_or0;
  wire [0:0] csa_component64_fa8_xor1;
  wire [0:0] csa_component64_fa8_or0;
  wire [0:0] csa_component64_fa9_xor1;
  wire [0:0] csa_component64_fa9_or0;
  wire [0:0] csa_component64_fa10_xor1;
  wire [0:0] csa_component64_fa10_or0;
  wire [0:0] csa_component64_fa11_xor1;
  wire [0:0] csa_component64_fa11_or0;
  wire [0:0] csa_component64_fa12_xor1;
  wire [0:0] csa_component64_fa12_or0;
  wire [0:0] csa_component64_fa13_xor1;
  wire [0:0] csa_component64_fa13_or0;
  wire [0:0] csa_component64_fa14_xor1;
  wire [0:0] csa_component64_fa14_or0;
  wire [0:0] csa_component64_fa15_xor1;
  wire [0:0] csa_component64_fa15_or0;
  wire [0:0] csa_component64_fa16_xor1;
  wire [0:0] csa_component64_fa16_or0;
  wire [0:0] csa_component64_fa17_xor1;
  wire [0:0] csa_component64_fa17_or0;
  wire [0:0] csa_component64_fa18_xor1;
  wire [0:0] csa_component64_fa18_or0;
  wire [0:0] csa_component64_fa19_xor1;
  wire [0:0] csa_component64_fa19_or0;
  wire [0:0] csa_component64_fa20_xor1;
  wire [0:0] csa_component64_fa20_or0;
  wire [0:0] csa_component64_fa21_xor1;
  wire [0:0] csa_component64_fa21_or0;
  wire [0:0] csa_component64_fa22_xor1;
  wire [0:0] csa_component64_fa22_or0;
  wire [0:0] csa_component64_fa23_xor1;
  wire [0:0] csa_component64_fa23_or0;
  wire [0:0] csa_component64_fa24_xor1;
  wire [0:0] csa_component64_fa24_or0;
  wire [0:0] csa_component64_fa25_xor1;
  wire [0:0] csa_component64_fa25_or0;
  wire [0:0] csa_component64_fa26_xor1;
  wire [0:0] csa_component64_fa26_or0;
  wire [0:0] csa_component64_fa27_xor1;
  wire [0:0] csa_component64_fa27_or0;
  wire [0:0] csa_component64_fa28_xor1;
  wire [0:0] csa_component64_fa28_or0;
  wire [0:0] csa_component64_fa29_xor1;
  wire [0:0] csa_component64_fa29_or0;
  wire [0:0] csa_component64_fa30_xor1;
  wire [0:0] csa_component64_fa30_or0;
  wire [0:0] csa_component64_fa31_xor1;
  wire [0:0] csa_component64_fa31_or0;
  wire [0:0] csa_component64_fa32_xor1;
  wire [0:0] csa_component64_fa32_or0;
  wire [0:0] csa_component64_fa33_xor1;
  wire [0:0] csa_component64_fa33_or0;
  wire [0:0] csa_component64_fa34_xor1;
  wire [0:0] csa_component64_fa34_or0;
  wire [0:0] csa_component64_fa35_xor1;
  wire [0:0] csa_component64_fa35_or0;
  wire [0:0] csa_component64_fa36_xor1;
  wire [0:0] csa_component64_fa36_or0;
  wire [0:0] csa_component64_fa37_xor1;
  wire [0:0] csa_component64_fa37_or0;
  wire [0:0] csa_component64_fa38_xor1;
  wire [0:0] csa_component64_fa38_or0;
  wire [0:0] csa_component64_fa39_xor1;
  wire [0:0] csa_component64_fa39_or0;
  wire [0:0] csa_component64_fa40_xor1;
  wire [0:0] csa_component64_fa40_or0;
  wire [0:0] csa_component64_fa41_xor1;
  wire [0:0] csa_component64_fa41_or0;
  wire [0:0] csa_component64_fa42_xor1;
  wire [0:0] csa_component64_fa42_or0;
  wire [0:0] csa_component64_fa43_xor1;
  wire [0:0] csa_component64_fa43_or0;
  wire [0:0] csa_component64_fa44_xor1;
  wire [0:0] csa_component64_fa44_or0;
  wire [0:0] csa_component64_fa45_xor1;
  wire [0:0] csa_component64_fa45_or0;
  wire [0:0] csa_component64_fa46_xor1;
  wire [0:0] csa_component64_fa46_or0;
  wire [0:0] csa_component64_fa47_xor1;
  wire [0:0] csa_component64_fa47_or0;
  wire [0:0] csa_component64_fa48_xor1;
  wire [0:0] csa_component64_fa48_or0;
  wire [0:0] csa_component64_fa49_xor1;
  wire [0:0] csa_component64_fa49_or0;
  wire [0:0] csa_component64_fa50_xor1;
  wire [0:0] csa_component64_fa50_or0;
  wire [0:0] csa_component64_fa51_xor1;
  wire [0:0] csa_component64_fa51_or0;
  wire [0:0] csa_component64_fa52_xor1;
  wire [0:0] csa_component64_fa52_or0;
  wire [0:0] csa_component64_fa53_xor1;
  wire [0:0] csa_component64_fa53_or0;
  wire [0:0] csa_component64_fa54_xor1;
  wire [0:0] csa_component64_fa54_or0;
  wire [0:0] csa_component64_fa55_xor1;
  wire [0:0] csa_component64_fa55_or0;
  wire [0:0] csa_component64_fa56_xor1;
  wire [0:0] csa_component64_fa56_or0;
  wire [0:0] csa_component64_fa57_xor1;
  wire [0:0] csa_component64_fa57_or0;
  wire [0:0] csa_component64_fa58_xor1;
  wire [0:0] csa_component64_fa58_or0;
  wire [0:0] csa_component64_fa59_xor1;
  wire [0:0] csa_component64_fa59_or0;
  wire [0:0] csa_component64_fa60_xor1;
  wire [0:0] csa_component64_fa60_or0;
  wire [0:0] csa_component64_fa61_xor1;
  wire [0:0] csa_component64_fa61_or0;
  wire [0:0] csa_component64_fa62_xor1;
  wire [0:0] csa_component64_fa62_or0;
  wire [0:0] csa_component64_fa63_xor1;
  wire [0:0] csa_component64_fa63_or0;

  fa fa_csa_component64_fa0_out(.a(a[0]), .b(b[0]), .cin(c[0]), .fa_xor1(csa_component64_fa0_xor1), .fa_or0(csa_component64_fa0_or0));
  fa fa_csa_component64_fa1_out(.a(a[1]), .b(b[1]), .cin(c[1]), .fa_xor1(csa_component64_fa1_xor1), .fa_or0(csa_component64_fa1_or0));
  fa fa_csa_component64_fa2_out(.a(a[2]), .b(b[2]), .cin(c[2]), .fa_xor1(csa_component64_fa2_xor1), .fa_or0(csa_component64_fa2_or0));
  fa fa_csa_component64_fa3_out(.a(a[3]), .b(b[3]), .cin(c[3]), .fa_xor1(csa_component64_fa3_xor1), .fa_or0(csa_component64_fa3_or0));
  fa fa_csa_component64_fa4_out(.a(a[4]), .b(b[4]), .cin(c[4]), .fa_xor1(csa_component64_fa4_xor1), .fa_or0(csa_component64_fa4_or0));
  fa fa_csa_component64_fa5_out(.a(a[5]), .b(b[5]), .cin(c[5]), .fa_xor1(csa_component64_fa5_xor1), .fa_or0(csa_component64_fa5_or0));
  fa fa_csa_component64_fa6_out(.a(a[6]), .b(b[6]), .cin(c[6]), .fa_xor1(csa_component64_fa6_xor1), .fa_or0(csa_component64_fa6_or0));
  fa fa_csa_component64_fa7_out(.a(a[7]), .b(b[7]), .cin(c[7]), .fa_xor1(csa_component64_fa7_xor1), .fa_or0(csa_component64_fa7_or0));
  fa fa_csa_component64_fa8_out(.a(a[8]), .b(b[8]), .cin(c[8]), .fa_xor1(csa_component64_fa8_xor1), .fa_or0(csa_component64_fa8_or0));
  fa fa_csa_component64_fa9_out(.a(a[9]), .b(b[9]), .cin(c[9]), .fa_xor1(csa_component64_fa9_xor1), .fa_or0(csa_component64_fa9_or0));
  fa fa_csa_component64_fa10_out(.a(a[10]), .b(b[10]), .cin(c[10]), .fa_xor1(csa_component64_fa10_xor1), .fa_or0(csa_component64_fa10_or0));
  fa fa_csa_component64_fa11_out(.a(a[11]), .b(b[11]), .cin(c[11]), .fa_xor1(csa_component64_fa11_xor1), .fa_or0(csa_component64_fa11_or0));
  fa fa_csa_component64_fa12_out(.a(a[12]), .b(b[12]), .cin(c[12]), .fa_xor1(csa_component64_fa12_xor1), .fa_or0(csa_component64_fa12_or0));
  fa fa_csa_component64_fa13_out(.a(a[13]), .b(b[13]), .cin(c[13]), .fa_xor1(csa_component64_fa13_xor1), .fa_or0(csa_component64_fa13_or0));
  fa fa_csa_component64_fa14_out(.a(a[14]), .b(b[14]), .cin(c[14]), .fa_xor1(csa_component64_fa14_xor1), .fa_or0(csa_component64_fa14_or0));
  fa fa_csa_component64_fa15_out(.a(a[15]), .b(b[15]), .cin(c[15]), .fa_xor1(csa_component64_fa15_xor1), .fa_or0(csa_component64_fa15_or0));
  fa fa_csa_component64_fa16_out(.a(a[16]), .b(b[16]), .cin(c[16]), .fa_xor1(csa_component64_fa16_xor1), .fa_or0(csa_component64_fa16_or0));
  fa fa_csa_component64_fa17_out(.a(a[17]), .b(b[17]), .cin(c[17]), .fa_xor1(csa_component64_fa17_xor1), .fa_or0(csa_component64_fa17_or0));
  fa fa_csa_component64_fa18_out(.a(a[18]), .b(b[18]), .cin(c[18]), .fa_xor1(csa_component64_fa18_xor1), .fa_or0(csa_component64_fa18_or0));
  fa fa_csa_component64_fa19_out(.a(a[19]), .b(b[19]), .cin(c[19]), .fa_xor1(csa_component64_fa19_xor1), .fa_or0(csa_component64_fa19_or0));
  fa fa_csa_component64_fa20_out(.a(a[20]), .b(b[20]), .cin(c[20]), .fa_xor1(csa_component64_fa20_xor1), .fa_or0(csa_component64_fa20_or0));
  fa fa_csa_component64_fa21_out(.a(a[21]), .b(b[21]), .cin(c[21]), .fa_xor1(csa_component64_fa21_xor1), .fa_or0(csa_component64_fa21_or0));
  fa fa_csa_component64_fa22_out(.a(a[22]), .b(b[22]), .cin(c[22]), .fa_xor1(csa_component64_fa22_xor1), .fa_or0(csa_component64_fa22_or0));
  fa fa_csa_component64_fa23_out(.a(a[23]), .b(b[23]), .cin(c[23]), .fa_xor1(csa_component64_fa23_xor1), .fa_or0(csa_component64_fa23_or0));
  fa fa_csa_component64_fa24_out(.a(a[24]), .b(b[24]), .cin(c[24]), .fa_xor1(csa_component64_fa24_xor1), .fa_or0(csa_component64_fa24_or0));
  fa fa_csa_component64_fa25_out(.a(a[25]), .b(b[25]), .cin(c[25]), .fa_xor1(csa_component64_fa25_xor1), .fa_or0(csa_component64_fa25_or0));
  fa fa_csa_component64_fa26_out(.a(a[26]), .b(b[26]), .cin(c[26]), .fa_xor1(csa_component64_fa26_xor1), .fa_or0(csa_component64_fa26_or0));
  fa fa_csa_component64_fa27_out(.a(a[27]), .b(b[27]), .cin(c[27]), .fa_xor1(csa_component64_fa27_xor1), .fa_or0(csa_component64_fa27_or0));
  fa fa_csa_component64_fa28_out(.a(a[28]), .b(b[28]), .cin(c[28]), .fa_xor1(csa_component64_fa28_xor1), .fa_or0(csa_component64_fa28_or0));
  fa fa_csa_component64_fa29_out(.a(a[29]), .b(b[29]), .cin(c[29]), .fa_xor1(csa_component64_fa29_xor1), .fa_or0(csa_component64_fa29_or0));
  fa fa_csa_component64_fa30_out(.a(a[30]), .b(b[30]), .cin(c[30]), .fa_xor1(csa_component64_fa30_xor1), .fa_or0(csa_component64_fa30_or0));
  fa fa_csa_component64_fa31_out(.a(a[31]), .b(b[31]), .cin(c[31]), .fa_xor1(csa_component64_fa31_xor1), .fa_or0(csa_component64_fa31_or0));
  fa fa_csa_component64_fa32_out(.a(a[32]), .b(b[32]), .cin(c[32]), .fa_xor1(csa_component64_fa32_xor1), .fa_or0(csa_component64_fa32_or0));
  fa fa_csa_component64_fa33_out(.a(a[33]), .b(b[33]), .cin(c[33]), .fa_xor1(csa_component64_fa33_xor1), .fa_or0(csa_component64_fa33_or0));
  fa fa_csa_component64_fa34_out(.a(a[34]), .b(b[34]), .cin(c[34]), .fa_xor1(csa_component64_fa34_xor1), .fa_or0(csa_component64_fa34_or0));
  fa fa_csa_component64_fa35_out(.a(a[35]), .b(b[35]), .cin(c[35]), .fa_xor1(csa_component64_fa35_xor1), .fa_or0(csa_component64_fa35_or0));
  fa fa_csa_component64_fa36_out(.a(a[36]), .b(b[36]), .cin(c[36]), .fa_xor1(csa_component64_fa36_xor1), .fa_or0(csa_component64_fa36_or0));
  fa fa_csa_component64_fa37_out(.a(a[37]), .b(b[37]), .cin(c[37]), .fa_xor1(csa_component64_fa37_xor1), .fa_or0(csa_component64_fa37_or0));
  fa fa_csa_component64_fa38_out(.a(a[38]), .b(b[38]), .cin(c[38]), .fa_xor1(csa_component64_fa38_xor1), .fa_or0(csa_component64_fa38_or0));
  fa fa_csa_component64_fa39_out(.a(a[39]), .b(b[39]), .cin(c[39]), .fa_xor1(csa_component64_fa39_xor1), .fa_or0(csa_component64_fa39_or0));
  fa fa_csa_component64_fa40_out(.a(a[40]), .b(b[40]), .cin(c[40]), .fa_xor1(csa_component64_fa40_xor1), .fa_or0(csa_component64_fa40_or0));
  fa fa_csa_component64_fa41_out(.a(a[41]), .b(b[41]), .cin(c[41]), .fa_xor1(csa_component64_fa41_xor1), .fa_or0(csa_component64_fa41_or0));
  fa fa_csa_component64_fa42_out(.a(a[42]), .b(b[42]), .cin(c[42]), .fa_xor1(csa_component64_fa42_xor1), .fa_or0(csa_component64_fa42_or0));
  fa fa_csa_component64_fa43_out(.a(a[43]), .b(b[43]), .cin(c[43]), .fa_xor1(csa_component64_fa43_xor1), .fa_or0(csa_component64_fa43_or0));
  fa fa_csa_component64_fa44_out(.a(a[44]), .b(b[44]), .cin(c[44]), .fa_xor1(csa_component64_fa44_xor1), .fa_or0(csa_component64_fa44_or0));
  fa fa_csa_component64_fa45_out(.a(a[45]), .b(b[45]), .cin(c[45]), .fa_xor1(csa_component64_fa45_xor1), .fa_or0(csa_component64_fa45_or0));
  fa fa_csa_component64_fa46_out(.a(a[46]), .b(b[46]), .cin(c[46]), .fa_xor1(csa_component64_fa46_xor1), .fa_or0(csa_component64_fa46_or0));
  fa fa_csa_component64_fa47_out(.a(a[47]), .b(b[47]), .cin(c[47]), .fa_xor1(csa_component64_fa47_xor1), .fa_or0(csa_component64_fa47_or0));
  fa fa_csa_component64_fa48_out(.a(a[48]), .b(b[48]), .cin(c[48]), .fa_xor1(csa_component64_fa48_xor1), .fa_or0(csa_component64_fa48_or0));
  fa fa_csa_component64_fa49_out(.a(a[49]), .b(b[49]), .cin(c[49]), .fa_xor1(csa_component64_fa49_xor1), .fa_or0(csa_component64_fa49_or0));
  fa fa_csa_component64_fa50_out(.a(a[50]), .b(b[50]), .cin(c[50]), .fa_xor1(csa_component64_fa50_xor1), .fa_or0(csa_component64_fa50_or0));
  fa fa_csa_component64_fa51_out(.a(a[51]), .b(b[51]), .cin(c[51]), .fa_xor1(csa_component64_fa51_xor1), .fa_or0(csa_component64_fa51_or0));
  fa fa_csa_component64_fa52_out(.a(a[52]), .b(b[52]), .cin(c[52]), .fa_xor1(csa_component64_fa52_xor1), .fa_or0(csa_component64_fa52_or0));
  fa fa_csa_component64_fa53_out(.a(a[53]), .b(b[53]), .cin(c[53]), .fa_xor1(csa_component64_fa53_xor1), .fa_or0(csa_component64_fa53_or0));
  fa fa_csa_component64_fa54_out(.a(a[54]), .b(b[54]), .cin(c[54]), .fa_xor1(csa_component64_fa54_xor1), .fa_or0(csa_component64_fa54_or0));
  fa fa_csa_component64_fa55_out(.a(a[55]), .b(b[55]), .cin(c[55]), .fa_xor1(csa_component64_fa55_xor1), .fa_or0(csa_component64_fa55_or0));
  fa fa_csa_component64_fa56_out(.a(a[56]), .b(b[56]), .cin(c[56]), .fa_xor1(csa_component64_fa56_xor1), .fa_or0(csa_component64_fa56_or0));
  fa fa_csa_component64_fa57_out(.a(a[57]), .b(b[57]), .cin(c[57]), .fa_xor1(csa_component64_fa57_xor1), .fa_or0(csa_component64_fa57_or0));
  fa fa_csa_component64_fa58_out(.a(a[58]), .b(b[58]), .cin(c[58]), .fa_xor1(csa_component64_fa58_xor1), .fa_or0(csa_component64_fa58_or0));
  fa fa_csa_component64_fa59_out(.a(a[59]), .b(b[59]), .cin(c[59]), .fa_xor1(csa_component64_fa59_xor1), .fa_or0(csa_component64_fa59_or0));
  fa fa_csa_component64_fa60_out(.a(a[60]), .b(b[60]), .cin(c[60]), .fa_xor1(csa_component64_fa60_xor1), .fa_or0(csa_component64_fa60_or0));
  fa fa_csa_component64_fa61_out(.a(a[61]), .b(b[61]), .cin(c[61]), .fa_xor1(csa_component64_fa61_xor1), .fa_or0(csa_component64_fa61_or0));
  fa fa_csa_component64_fa62_out(.a(a[62]), .b(b[62]), .cin(c[62]), .fa_xor1(csa_component64_fa62_xor1), .fa_or0(csa_component64_fa62_or0));
  fa fa_csa_component64_fa63_out(.a(a[63]), .b(b[63]), .cin(c[63]), .fa_xor1(csa_component64_fa63_xor1), .fa_or0(csa_component64_fa63_or0));

  assign csa_component64_out[0] = csa_component64_fa0_xor1[0];
  assign csa_component64_out[1] = csa_component64_fa1_xor1[0];
  assign csa_component64_out[2] = csa_component64_fa2_xor1[0];
  assign csa_component64_out[3] = csa_component64_fa3_xor1[0];
  assign csa_component64_out[4] = csa_component64_fa4_xor1[0];
  assign csa_component64_out[5] = csa_component64_fa5_xor1[0];
  assign csa_component64_out[6] = csa_component64_fa6_xor1[0];
  assign csa_component64_out[7] = csa_component64_fa7_xor1[0];
  assign csa_component64_out[8] = csa_component64_fa8_xor1[0];
  assign csa_component64_out[9] = csa_component64_fa9_xor1[0];
  assign csa_component64_out[10] = csa_component64_fa10_xor1[0];
  assign csa_component64_out[11] = csa_component64_fa11_xor1[0];
  assign csa_component64_out[12] = csa_component64_fa12_xor1[0];
  assign csa_component64_out[13] = csa_component64_fa13_xor1[0];
  assign csa_component64_out[14] = csa_component64_fa14_xor1[0];
  assign csa_component64_out[15] = csa_component64_fa15_xor1[0];
  assign csa_component64_out[16] = csa_component64_fa16_xor1[0];
  assign csa_component64_out[17] = csa_component64_fa17_xor1[0];
  assign csa_component64_out[18] = csa_component64_fa18_xor1[0];
  assign csa_component64_out[19] = csa_component64_fa19_xor1[0];
  assign csa_component64_out[20] = csa_component64_fa20_xor1[0];
  assign csa_component64_out[21] = csa_component64_fa21_xor1[0];
  assign csa_component64_out[22] = csa_component64_fa22_xor1[0];
  assign csa_component64_out[23] = csa_component64_fa23_xor1[0];
  assign csa_component64_out[24] = csa_component64_fa24_xor1[0];
  assign csa_component64_out[25] = csa_component64_fa25_xor1[0];
  assign csa_component64_out[26] = csa_component64_fa26_xor1[0];
  assign csa_component64_out[27] = csa_component64_fa27_xor1[0];
  assign csa_component64_out[28] = csa_component64_fa28_xor1[0];
  assign csa_component64_out[29] = csa_component64_fa29_xor1[0];
  assign csa_component64_out[30] = csa_component64_fa30_xor1[0];
  assign csa_component64_out[31] = csa_component64_fa31_xor1[0];
  assign csa_component64_out[32] = csa_component64_fa32_xor1[0];
  assign csa_component64_out[33] = csa_component64_fa33_xor1[0];
  assign csa_component64_out[34] = csa_component64_fa34_xor1[0];
  assign csa_component64_out[35] = csa_component64_fa35_xor1[0];
  assign csa_component64_out[36] = csa_component64_fa36_xor1[0];
  assign csa_component64_out[37] = csa_component64_fa37_xor1[0];
  assign csa_component64_out[38] = csa_component64_fa38_xor1[0];
  assign csa_component64_out[39] = csa_component64_fa39_xor1[0];
  assign csa_component64_out[40] = csa_component64_fa40_xor1[0];
  assign csa_component64_out[41] = csa_component64_fa41_xor1[0];
  assign csa_component64_out[42] = csa_component64_fa42_xor1[0];
  assign csa_component64_out[43] = csa_component64_fa43_xor1[0];
  assign csa_component64_out[44] = csa_component64_fa44_xor1[0];
  assign csa_component64_out[45] = csa_component64_fa45_xor1[0];
  assign csa_component64_out[46] = csa_component64_fa46_xor1[0];
  assign csa_component64_out[47] = csa_component64_fa47_xor1[0];
  assign csa_component64_out[48] = csa_component64_fa48_xor1[0];
  assign csa_component64_out[49] = csa_component64_fa49_xor1[0];
  assign csa_component64_out[50] = csa_component64_fa50_xor1[0];
  assign csa_component64_out[51] = csa_component64_fa51_xor1[0];
  assign csa_component64_out[52] = csa_component64_fa52_xor1[0];
  assign csa_component64_out[53] = csa_component64_fa53_xor1[0];
  assign csa_component64_out[54] = csa_component64_fa54_xor1[0];
  assign csa_component64_out[55] = csa_component64_fa55_xor1[0];
  assign csa_component64_out[56] = csa_component64_fa56_xor1[0];
  assign csa_component64_out[57] = csa_component64_fa57_xor1[0];
  assign csa_component64_out[58] = csa_component64_fa58_xor1[0];
  assign csa_component64_out[59] = csa_component64_fa59_xor1[0];
  assign csa_component64_out[60] = csa_component64_fa60_xor1[0];
  assign csa_component64_out[61] = csa_component64_fa61_xor1[0];
  assign csa_component64_out[62] = csa_component64_fa62_xor1[0];
  assign csa_component64_out[63] = csa_component64_fa63_xor1[0];
  assign csa_component64_out[64] = 1'b0;
  assign csa_component64_out[65] = 1'b0;
  assign csa_component64_out[66] = csa_component64_fa0_or0[0];
  assign csa_component64_out[67] = csa_component64_fa1_or0[0];
  assign csa_component64_out[68] = csa_component64_fa2_or0[0];
  assign csa_component64_out[69] = csa_component64_fa3_or0[0];
  assign csa_component64_out[70] = csa_component64_fa4_or0[0];
  assign csa_component64_out[71] = csa_component64_fa5_or0[0];
  assign csa_component64_out[72] = csa_component64_fa6_or0[0];
  assign csa_component64_out[73] = csa_component64_fa7_or0[0];
  assign csa_component64_out[74] = csa_component64_fa8_or0[0];
  assign csa_component64_out[75] = csa_component64_fa9_or0[0];
  assign csa_component64_out[76] = csa_component64_fa10_or0[0];
  assign csa_component64_out[77] = csa_component64_fa11_or0[0];
  assign csa_component64_out[78] = csa_component64_fa12_or0[0];
  assign csa_component64_out[79] = csa_component64_fa13_or0[0];
  assign csa_component64_out[80] = csa_component64_fa14_or0[0];
  assign csa_component64_out[81] = csa_component64_fa15_or0[0];
  assign csa_component64_out[82] = csa_component64_fa16_or0[0];
  assign csa_component64_out[83] = csa_component64_fa17_or0[0];
  assign csa_component64_out[84] = csa_component64_fa18_or0[0];
  assign csa_component64_out[85] = csa_component64_fa19_or0[0];
  assign csa_component64_out[86] = csa_component64_fa20_or0[0];
  assign csa_component64_out[87] = csa_component64_fa21_or0[0];
  assign csa_component64_out[88] = csa_component64_fa22_or0[0];
  assign csa_component64_out[89] = csa_component64_fa23_or0[0];
  assign csa_component64_out[90] = csa_component64_fa24_or0[0];
  assign csa_component64_out[91] = csa_component64_fa25_or0[0];
  assign csa_component64_out[92] = csa_component64_fa26_or0[0];
  assign csa_component64_out[93] = csa_component64_fa27_or0[0];
  assign csa_component64_out[94] = csa_component64_fa28_or0[0];
  assign csa_component64_out[95] = csa_component64_fa29_or0[0];
  assign csa_component64_out[96] = csa_component64_fa30_or0[0];
  assign csa_component64_out[97] = csa_component64_fa31_or0[0];
  assign csa_component64_out[98] = csa_component64_fa32_or0[0];
  assign csa_component64_out[99] = csa_component64_fa33_or0[0];
  assign csa_component64_out[100] = csa_component64_fa34_or0[0];
  assign csa_component64_out[101] = csa_component64_fa35_or0[0];
  assign csa_component64_out[102] = csa_component64_fa36_or0[0];
  assign csa_component64_out[103] = csa_component64_fa37_or0[0];
  assign csa_component64_out[104] = csa_component64_fa38_or0[0];
  assign csa_component64_out[105] = csa_component64_fa39_or0[0];
  assign csa_component64_out[106] = csa_component64_fa40_or0[0];
  assign csa_component64_out[107] = csa_component64_fa41_or0[0];
  assign csa_component64_out[108] = csa_component64_fa42_or0[0];
  assign csa_component64_out[109] = csa_component64_fa43_or0[0];
  assign csa_component64_out[110] = csa_component64_fa44_or0[0];
  assign csa_component64_out[111] = csa_component64_fa45_or0[0];
  assign csa_component64_out[112] = csa_component64_fa46_or0[0];
  assign csa_component64_out[113] = csa_component64_fa47_or0[0];
  assign csa_component64_out[114] = csa_component64_fa48_or0[0];
  assign csa_component64_out[115] = csa_component64_fa49_or0[0];
  assign csa_component64_out[116] = csa_component64_fa50_or0[0];
  assign csa_component64_out[117] = csa_component64_fa51_or0[0];
  assign csa_component64_out[118] = csa_component64_fa52_or0[0];
  assign csa_component64_out[119] = csa_component64_fa53_or0[0];
  assign csa_component64_out[120] = csa_component64_fa54_or0[0];
  assign csa_component64_out[121] = csa_component64_fa55_or0[0];
  assign csa_component64_out[122] = csa_component64_fa56_or0[0];
  assign csa_component64_out[123] = csa_component64_fa57_or0[0];
  assign csa_component64_out[124] = csa_component64_fa58_or0[0];
  assign csa_component64_out[125] = csa_component64_fa59_or0[0];
  assign csa_component64_out[126] = csa_component64_fa60_or0[0];
  assign csa_component64_out[127] = csa_component64_fa61_or0[0];
  assign csa_component64_out[128] = csa_component64_fa62_or0[0];
  assign csa_component64_out[129] = csa_component64_fa63_or0[0];
endmodule

module u_pg_rca64(input [63:0] a, input [63:0] b, output [64:0] u_pg_rca64_out);
  wire [0:0] u_pg_rca64_pg_fa0_xor0;
  wire [0:0] u_pg_rca64_pg_fa0_and0;
  wire [0:0] u_pg_rca64_pg_fa1_xor0;
  wire [0:0] u_pg_rca64_pg_fa1_and0;
  wire [0:0] u_pg_rca64_pg_fa1_xor1;
  wire [0:0] u_pg_rca64_and1;
  wire [0:0] u_pg_rca64_or1;
  wire [0:0] u_pg_rca64_pg_fa2_xor0;
  wire [0:0] u_pg_rca64_pg_fa2_and0;
  wire [0:0] u_pg_rca64_pg_fa2_xor1;
  wire [0:0] u_pg_rca64_and2;
  wire [0:0] u_pg_rca64_or2;
  wire [0:0] u_pg_rca64_pg_fa3_xor0;
  wire [0:0] u_pg_rca64_pg_fa3_and0;
  wire [0:0] u_pg_rca64_pg_fa3_xor1;
  wire [0:0] u_pg_rca64_and3;
  wire [0:0] u_pg_rca64_or3;
  wire [0:0] u_pg_rca64_pg_fa4_xor0;
  wire [0:0] u_pg_rca64_pg_fa4_and0;
  wire [0:0] u_pg_rca64_pg_fa4_xor1;
  wire [0:0] u_pg_rca64_and4;
  wire [0:0] u_pg_rca64_or4;
  wire [0:0] u_pg_rca64_pg_fa5_xor0;
  wire [0:0] u_pg_rca64_pg_fa5_and0;
  wire [0:0] u_pg_rca64_pg_fa5_xor1;
  wire [0:0] u_pg_rca64_and5;
  wire [0:0] u_pg_rca64_or5;
  wire [0:0] u_pg_rca64_pg_fa6_xor0;
  wire [0:0] u_pg_rca64_pg_fa6_and0;
  wire [0:0] u_pg_rca64_pg_fa6_xor1;
  wire [0:0] u_pg_rca64_and6;
  wire [0:0] u_pg_rca64_or6;
  wire [0:0] u_pg_rca64_pg_fa7_xor0;
  wire [0:0] u_pg_rca64_pg_fa7_and0;
  wire [0:0] u_pg_rca64_pg_fa7_xor1;
  wire [0:0] u_pg_rca64_and7;
  wire [0:0] u_pg_rca64_or7;
  wire [0:0] u_pg_rca64_pg_fa8_xor0;
  wire [0:0] u_pg_rca64_pg_fa8_and0;
  wire [0:0] u_pg_rca64_pg_fa8_xor1;
  wire [0:0] u_pg_rca64_and8;
  wire [0:0] u_pg_rca64_or8;
  wire [0:0] u_pg_rca64_pg_fa9_xor0;
  wire [0:0] u_pg_rca64_pg_fa9_and0;
  wire [0:0] u_pg_rca64_pg_fa9_xor1;
  wire [0:0] u_pg_rca64_and9;
  wire [0:0] u_pg_rca64_or9;
  wire [0:0] u_pg_rca64_pg_fa10_xor0;
  wire [0:0] u_pg_rca64_pg_fa10_and0;
  wire [0:0] u_pg_rca64_pg_fa10_xor1;
  wire [0:0] u_pg_rca64_and10;
  wire [0:0] u_pg_rca64_or10;
  wire [0:0] u_pg_rca64_pg_fa11_xor0;
  wire [0:0] u_pg_rca64_pg_fa11_and0;
  wire [0:0] u_pg_rca64_pg_fa11_xor1;
  wire [0:0] u_pg_rca64_and11;
  wire [0:0] u_pg_rca64_or11;
  wire [0:0] u_pg_rca64_pg_fa12_xor0;
  wire [0:0] u_pg_rca64_pg_fa12_and0;
  wire [0:0] u_pg_rca64_pg_fa12_xor1;
  wire [0:0] u_pg_rca64_and12;
  wire [0:0] u_pg_rca64_or12;
  wire [0:0] u_pg_rca64_pg_fa13_xor0;
  wire [0:0] u_pg_rca64_pg_fa13_and0;
  wire [0:0] u_pg_rca64_pg_fa13_xor1;
  wire [0:0] u_pg_rca64_and13;
  wire [0:0] u_pg_rca64_or13;
  wire [0:0] u_pg_rca64_pg_fa14_xor0;
  wire [0:0] u_pg_rca64_pg_fa14_and0;
  wire [0:0] u_pg_rca64_pg_fa14_xor1;
  wire [0:0] u_pg_rca64_and14;
  wire [0:0] u_pg_rca64_or14;
  wire [0:0] u_pg_rca64_pg_fa15_xor0;
  wire [0:0] u_pg_rca64_pg_fa15_and0;
  wire [0:0] u_pg_rca64_pg_fa15_xor1;
  wire [0:0] u_pg_rca64_and15;
  wire [0:0] u_pg_rca64_or15;
  wire [0:0] u_pg_rca64_pg_fa16_xor0;
  wire [0:0] u_pg_rca64_pg_fa16_and0;
  wire [0:0] u_pg_rca64_pg_fa16_xor1;
  wire [0:0] u_pg_rca64_and16;
  wire [0:0] u_pg_rca64_or16;
  wire [0:0] u_pg_rca64_pg_fa17_xor0;
  wire [0:0] u_pg_rca64_pg_fa17_and0;
  wire [0:0] u_pg_rca64_pg_fa17_xor1;
  wire [0:0] u_pg_rca64_and17;
  wire [0:0] u_pg_rca64_or17;
  wire [0:0] u_pg_rca64_pg_fa18_xor0;
  wire [0:0] u_pg_rca64_pg_fa18_and0;
  wire [0:0] u_pg_rca64_pg_fa18_xor1;
  wire [0:0] u_pg_rca64_and18;
  wire [0:0] u_pg_rca64_or18;
  wire [0:0] u_pg_rca64_pg_fa19_xor0;
  wire [0:0] u_pg_rca64_pg_fa19_and0;
  wire [0:0] u_pg_rca64_pg_fa19_xor1;
  wire [0:0] u_pg_rca64_and19;
  wire [0:0] u_pg_rca64_or19;
  wire [0:0] u_pg_rca64_pg_fa20_xor0;
  wire [0:0] u_pg_rca64_pg_fa20_and0;
  wire [0:0] u_pg_rca64_pg_fa20_xor1;
  wire [0:0] u_pg_rca64_and20;
  wire [0:0] u_pg_rca64_or20;
  wire [0:0] u_pg_rca64_pg_fa21_xor0;
  wire [0:0] u_pg_rca64_pg_fa21_and0;
  wire [0:0] u_pg_rca64_pg_fa21_xor1;
  wire [0:0] u_pg_rca64_and21;
  wire [0:0] u_pg_rca64_or21;
  wire [0:0] u_pg_rca64_pg_fa22_xor0;
  wire [0:0] u_pg_rca64_pg_fa22_and0;
  wire [0:0] u_pg_rca64_pg_fa22_xor1;
  wire [0:0] u_pg_rca64_and22;
  wire [0:0] u_pg_rca64_or22;
  wire [0:0] u_pg_rca64_pg_fa23_xor0;
  wire [0:0] u_pg_rca64_pg_fa23_and0;
  wire [0:0] u_pg_rca64_pg_fa23_xor1;
  wire [0:0] u_pg_rca64_and23;
  wire [0:0] u_pg_rca64_or23;
  wire [0:0] u_pg_rca64_pg_fa24_xor0;
  wire [0:0] u_pg_rca64_pg_fa24_and0;
  wire [0:0] u_pg_rca64_pg_fa24_xor1;
  wire [0:0] u_pg_rca64_and24;
  wire [0:0] u_pg_rca64_or24;
  wire [0:0] u_pg_rca64_pg_fa25_xor0;
  wire [0:0] u_pg_rca64_pg_fa25_and0;
  wire [0:0] u_pg_rca64_pg_fa25_xor1;
  wire [0:0] u_pg_rca64_and25;
  wire [0:0] u_pg_rca64_or25;
  wire [0:0] u_pg_rca64_pg_fa26_xor0;
  wire [0:0] u_pg_rca64_pg_fa26_and0;
  wire [0:0] u_pg_rca64_pg_fa26_xor1;
  wire [0:0] u_pg_rca64_and26;
  wire [0:0] u_pg_rca64_or26;
  wire [0:0] u_pg_rca64_pg_fa27_xor0;
  wire [0:0] u_pg_rca64_pg_fa27_and0;
  wire [0:0] u_pg_rca64_pg_fa27_xor1;
  wire [0:0] u_pg_rca64_and27;
  wire [0:0] u_pg_rca64_or27;
  wire [0:0] u_pg_rca64_pg_fa28_xor0;
  wire [0:0] u_pg_rca64_pg_fa28_and0;
  wire [0:0] u_pg_rca64_pg_fa28_xor1;
  wire [0:0] u_pg_rca64_and28;
  wire [0:0] u_pg_rca64_or28;
  wire [0:0] u_pg_rca64_pg_fa29_xor0;
  wire [0:0] u_pg_rca64_pg_fa29_and0;
  wire [0:0] u_pg_rca64_pg_fa29_xor1;
  wire [0:0] u_pg_rca64_and29;
  wire [0:0] u_pg_rca64_or29;
  wire [0:0] u_pg_rca64_pg_fa30_xor0;
  wire [0:0] u_pg_rca64_pg_fa30_and0;
  wire [0:0] u_pg_rca64_pg_fa30_xor1;
  wire [0:0] u_pg_rca64_and30;
  wire [0:0] u_pg_rca64_or30;
  wire [0:0] u_pg_rca64_pg_fa31_xor0;
  wire [0:0] u_pg_rca64_pg_fa31_and0;
  wire [0:0] u_pg_rca64_pg_fa31_xor1;
  wire [0:0] u_pg_rca64_and31;
  wire [0:0] u_pg_rca64_or31;
  wire [0:0] u_pg_rca64_pg_fa32_xor0;
  wire [0:0] u_pg_rca64_pg_fa32_and0;
  wire [0:0] u_pg_rca64_pg_fa32_xor1;
  wire [0:0] u_pg_rca64_and32;
  wire [0:0] u_pg_rca64_or32;
  wire [0:0] u_pg_rca64_pg_fa33_xor0;
  wire [0:0] u_pg_rca64_pg_fa33_and0;
  wire [0:0] u_pg_rca64_pg_fa33_xor1;
  wire [0:0] u_pg_rca64_and33;
  wire [0:0] u_pg_rca64_or33;
  wire [0:0] u_pg_rca64_pg_fa34_xor0;
  wire [0:0] u_pg_rca64_pg_fa34_and0;
  wire [0:0] u_pg_rca64_pg_fa34_xor1;
  wire [0:0] u_pg_rca64_and34;
  wire [0:0] u_pg_rca64_or34;
  wire [0:0] u_pg_rca64_pg_fa35_xor0;
  wire [0:0] u_pg_rca64_pg_fa35_and0;
  wire [0:0] u_pg_rca64_pg_fa35_xor1;
  wire [0:0] u_pg_rca64_and35;
  wire [0:0] u_pg_rca64_or35;
  wire [0:0] u_pg_rca64_pg_fa36_xor0;
  wire [0:0] u_pg_rca64_pg_fa36_and0;
  wire [0:0] u_pg_rca64_pg_fa36_xor1;
  wire [0:0] u_pg_rca64_and36;
  wire [0:0] u_pg_rca64_or36;
  wire [0:0] u_pg_rca64_pg_fa37_xor0;
  wire [0:0] u_pg_rca64_pg_fa37_and0;
  wire [0:0] u_pg_rca64_pg_fa37_xor1;
  wire [0:0] u_pg_rca64_and37;
  wire [0:0] u_pg_rca64_or37;
  wire [0:0] u_pg_rca64_pg_fa38_xor0;
  wire [0:0] u_pg_rca64_pg_fa38_and0;
  wire [0:0] u_pg_rca64_pg_fa38_xor1;
  wire [0:0] u_pg_rca64_and38;
  wire [0:0] u_pg_rca64_or38;
  wire [0:0] u_pg_rca64_pg_fa39_xor0;
  wire [0:0] u_pg_rca64_pg_fa39_and0;
  wire [0:0] u_pg_rca64_pg_fa39_xor1;
  wire [0:0] u_pg_rca64_and39;
  wire [0:0] u_pg_rca64_or39;
  wire [0:0] u_pg_rca64_pg_fa40_xor0;
  wire [0:0] u_pg_rca64_pg_fa40_and0;
  wire [0:0] u_pg_rca64_pg_fa40_xor1;
  wire [0:0] u_pg_rca64_and40;
  wire [0:0] u_pg_rca64_or40;
  wire [0:0] u_pg_rca64_pg_fa41_xor0;
  wire [0:0] u_pg_rca64_pg_fa41_and0;
  wire [0:0] u_pg_rca64_pg_fa41_xor1;
  wire [0:0] u_pg_rca64_and41;
  wire [0:0] u_pg_rca64_or41;
  wire [0:0] u_pg_rca64_pg_fa42_xor0;
  wire [0:0] u_pg_rca64_pg_fa42_and0;
  wire [0:0] u_pg_rca64_pg_fa42_xor1;
  wire [0:0] u_pg_rca64_and42;
  wire [0:0] u_pg_rca64_or42;
  wire [0:0] u_pg_rca64_pg_fa43_xor0;
  wire [0:0] u_pg_rca64_pg_fa43_and0;
  wire [0:0] u_pg_rca64_pg_fa43_xor1;
  wire [0:0] u_pg_rca64_and43;
  wire [0:0] u_pg_rca64_or43;
  wire [0:0] u_pg_rca64_pg_fa44_xor0;
  wire [0:0] u_pg_rca64_pg_fa44_and0;
  wire [0:0] u_pg_rca64_pg_fa44_xor1;
  wire [0:0] u_pg_rca64_and44;
  wire [0:0] u_pg_rca64_or44;
  wire [0:0] u_pg_rca64_pg_fa45_xor0;
  wire [0:0] u_pg_rca64_pg_fa45_and0;
  wire [0:0] u_pg_rca64_pg_fa45_xor1;
  wire [0:0] u_pg_rca64_and45;
  wire [0:0] u_pg_rca64_or45;
  wire [0:0] u_pg_rca64_pg_fa46_xor0;
  wire [0:0] u_pg_rca64_pg_fa46_and0;
  wire [0:0] u_pg_rca64_pg_fa46_xor1;
  wire [0:0] u_pg_rca64_and46;
  wire [0:0] u_pg_rca64_or46;
  wire [0:0] u_pg_rca64_pg_fa47_xor0;
  wire [0:0] u_pg_rca64_pg_fa47_and0;
  wire [0:0] u_pg_rca64_pg_fa47_xor1;
  wire [0:0] u_pg_rca64_and47;
  wire [0:0] u_pg_rca64_or47;
  wire [0:0] u_pg_rca64_pg_fa48_xor0;
  wire [0:0] u_pg_rca64_pg_fa48_and0;
  wire [0:0] u_pg_rca64_pg_fa48_xor1;
  wire [0:0] u_pg_rca64_and48;
  wire [0:0] u_pg_rca64_or48;
  wire [0:0] u_pg_rca64_pg_fa49_xor0;
  wire [0:0] u_pg_rca64_pg_fa49_and0;
  wire [0:0] u_pg_rca64_pg_fa49_xor1;
  wire [0:0] u_pg_rca64_and49;
  wire [0:0] u_pg_rca64_or49;
  wire [0:0] u_pg_rca64_pg_fa50_xor0;
  wire [0:0] u_pg_rca64_pg_fa50_and0;
  wire [0:0] u_pg_rca64_pg_fa50_xor1;
  wire [0:0] u_pg_rca64_and50;
  wire [0:0] u_pg_rca64_or50;
  wire [0:0] u_pg_rca64_pg_fa51_xor0;
  wire [0:0] u_pg_rca64_pg_fa51_and0;
  wire [0:0] u_pg_rca64_pg_fa51_xor1;
  wire [0:0] u_pg_rca64_and51;
  wire [0:0] u_pg_rca64_or51;
  wire [0:0] u_pg_rca64_pg_fa52_xor0;
  wire [0:0] u_pg_rca64_pg_fa52_and0;
  wire [0:0] u_pg_rca64_pg_fa52_xor1;
  wire [0:0] u_pg_rca64_and52;
  wire [0:0] u_pg_rca64_or52;
  wire [0:0] u_pg_rca64_pg_fa53_xor0;
  wire [0:0] u_pg_rca64_pg_fa53_and0;
  wire [0:0] u_pg_rca64_pg_fa53_xor1;
  wire [0:0] u_pg_rca64_and53;
  wire [0:0] u_pg_rca64_or53;
  wire [0:0] u_pg_rca64_pg_fa54_xor0;
  wire [0:0] u_pg_rca64_pg_fa54_and0;
  wire [0:0] u_pg_rca64_pg_fa54_xor1;
  wire [0:0] u_pg_rca64_and54;
  wire [0:0] u_pg_rca64_or54;
  wire [0:0] u_pg_rca64_pg_fa55_xor0;
  wire [0:0] u_pg_rca64_pg_fa55_and0;
  wire [0:0] u_pg_rca64_pg_fa55_xor1;
  wire [0:0] u_pg_rca64_and55;
  wire [0:0] u_pg_rca64_or55;
  wire [0:0] u_pg_rca64_pg_fa56_xor0;
  wire [0:0] u_pg_rca64_pg_fa56_and0;
  wire [0:0] u_pg_rca64_pg_fa56_xor1;
  wire [0:0] u_pg_rca64_and56;
  wire [0:0] u_pg_rca64_or56;
  wire [0:0] u_pg_rca64_pg_fa57_xor0;
  wire [0:0] u_pg_rca64_pg_fa57_and0;
  wire [0:0] u_pg_rca64_pg_fa57_xor1;
  wire [0:0] u_pg_rca64_and57;
  wire [0:0] u_pg_rca64_or57;
  wire [0:0] u_pg_rca64_pg_fa58_xor0;
  wire [0:0] u_pg_rca64_pg_fa58_and0;
  wire [0:0] u_pg_rca64_pg_fa58_xor1;
  wire [0:0] u_pg_rca64_and58;
  wire [0:0] u_pg_rca64_or58;
  wire [0:0] u_pg_rca64_pg_fa59_xor0;
  wire [0:0] u_pg_rca64_pg_fa59_and0;
  wire [0:0] u_pg_rca64_pg_fa59_xor1;
  wire [0:0] u_pg_rca64_and59;
  wire [0:0] u_pg_rca64_or59;
  wire [0:0] u_pg_rca64_pg_fa60_xor0;
  wire [0:0] u_pg_rca64_pg_fa60_and0;
  wire [0:0] u_pg_rca64_pg_fa60_xor1;
  wire [0:0] u_pg_rca64_and60;
  wire [0:0] u_pg_rca64_or60;
  wire [0:0] u_pg_rca64_pg_fa61_xor0;
  wire [0:0] u_pg_rca64_pg_fa61_and0;
  wire [0:0] u_pg_rca64_pg_fa61_xor1;
  wire [0:0] u_pg_rca64_and61;
  wire [0:0] u_pg_rca64_or61;
  wire [0:0] u_pg_rca64_pg_fa62_xor0;
  wire [0:0] u_pg_rca64_pg_fa62_and0;
  wire [0:0] u_pg_rca64_pg_fa62_xor1;
  wire [0:0] u_pg_rca64_and62;
  wire [0:0] u_pg_rca64_or62;
  wire [0:0] u_pg_rca64_pg_fa63_xor0;
  wire [0:0] u_pg_rca64_pg_fa63_and0;
  wire [0:0] u_pg_rca64_pg_fa63_xor1;
  wire [0:0] u_pg_rca64_and63;
  wire [0:0] u_pg_rca64_or63;

  pg_fa pg_fa_u_pg_rca64_pg_fa0_out(.a(a[0]), .b(b[0]), .cin(1'b0), .pg_fa_xor0(u_pg_rca64_pg_fa0_xor0), .pg_fa_and0(u_pg_rca64_pg_fa0_and0), .pg_fa_xor1());
  pg_fa pg_fa_u_pg_rca64_pg_fa1_out(.a(a[1]), .b(b[1]), .cin(u_pg_rca64_pg_fa0_and0[0]), .pg_fa_xor0(u_pg_rca64_pg_fa1_xor0), .pg_fa_and0(u_pg_rca64_pg_fa1_and0), .pg_fa_xor1(u_pg_rca64_pg_fa1_xor1));
  and_gate and_gate_u_pg_rca64_and1(.a(u_pg_rca64_pg_fa0_and0[0]), .b(u_pg_rca64_pg_fa1_xor0[0]), .out(u_pg_rca64_and1));
  or_gate or_gate_u_pg_rca64_or1(.a(u_pg_rca64_and1[0]), .b(u_pg_rca64_pg_fa1_and0[0]), .out(u_pg_rca64_or1));
  pg_fa pg_fa_u_pg_rca64_pg_fa2_out(.a(a[2]), .b(b[2]), .cin(u_pg_rca64_or1[0]), .pg_fa_xor0(u_pg_rca64_pg_fa2_xor0), .pg_fa_and0(u_pg_rca64_pg_fa2_and0), .pg_fa_xor1(u_pg_rca64_pg_fa2_xor1));
  and_gate and_gate_u_pg_rca64_and2(.a(u_pg_rca64_or1[0]), .b(u_pg_rca64_pg_fa2_xor0[0]), .out(u_pg_rca64_and2));
  or_gate or_gate_u_pg_rca64_or2(.a(u_pg_rca64_and2[0]), .b(u_pg_rca64_pg_fa2_and0[0]), .out(u_pg_rca64_or2));
  pg_fa pg_fa_u_pg_rca64_pg_fa3_out(.a(a[3]), .b(b[3]), .cin(u_pg_rca64_or2[0]), .pg_fa_xor0(u_pg_rca64_pg_fa3_xor0), .pg_fa_and0(u_pg_rca64_pg_fa3_and0), .pg_fa_xor1(u_pg_rca64_pg_fa3_xor1));
  and_gate and_gate_u_pg_rca64_and3(.a(u_pg_rca64_or2[0]), .b(u_pg_rca64_pg_fa3_xor0[0]), .out(u_pg_rca64_and3));
  or_gate or_gate_u_pg_rca64_or3(.a(u_pg_rca64_and3[0]), .b(u_pg_rca64_pg_fa3_and0[0]), .out(u_pg_rca64_or3));
  pg_fa pg_fa_u_pg_rca64_pg_fa4_out(.a(a[4]), .b(b[4]), .cin(u_pg_rca64_or3[0]), .pg_fa_xor0(u_pg_rca64_pg_fa4_xor0), .pg_fa_and0(u_pg_rca64_pg_fa4_and0), .pg_fa_xor1(u_pg_rca64_pg_fa4_xor1));
  and_gate and_gate_u_pg_rca64_and4(.a(u_pg_rca64_or3[0]), .b(u_pg_rca64_pg_fa4_xor0[0]), .out(u_pg_rca64_and4));
  or_gate or_gate_u_pg_rca64_or4(.a(u_pg_rca64_and4[0]), .b(u_pg_rca64_pg_fa4_and0[0]), .out(u_pg_rca64_or4));
  pg_fa pg_fa_u_pg_rca64_pg_fa5_out(.a(a[5]), .b(b[5]), .cin(u_pg_rca64_or4[0]), .pg_fa_xor0(u_pg_rca64_pg_fa5_xor0), .pg_fa_and0(u_pg_rca64_pg_fa5_and0), .pg_fa_xor1(u_pg_rca64_pg_fa5_xor1));
  and_gate and_gate_u_pg_rca64_and5(.a(u_pg_rca64_or4[0]), .b(u_pg_rca64_pg_fa5_xor0[0]), .out(u_pg_rca64_and5));
  or_gate or_gate_u_pg_rca64_or5(.a(u_pg_rca64_and5[0]), .b(u_pg_rca64_pg_fa5_and0[0]), .out(u_pg_rca64_or5));
  pg_fa pg_fa_u_pg_rca64_pg_fa6_out(.a(a[6]), .b(b[6]), .cin(u_pg_rca64_or5[0]), .pg_fa_xor0(u_pg_rca64_pg_fa6_xor0), .pg_fa_and0(u_pg_rca64_pg_fa6_and0), .pg_fa_xor1(u_pg_rca64_pg_fa6_xor1));
  and_gate and_gate_u_pg_rca64_and6(.a(u_pg_rca64_or5[0]), .b(u_pg_rca64_pg_fa6_xor0[0]), .out(u_pg_rca64_and6));
  or_gate or_gate_u_pg_rca64_or6(.a(u_pg_rca64_and6[0]), .b(u_pg_rca64_pg_fa6_and0[0]), .out(u_pg_rca64_or6));
  pg_fa pg_fa_u_pg_rca64_pg_fa7_out(.a(a[7]), .b(b[7]), .cin(u_pg_rca64_or6[0]), .pg_fa_xor0(u_pg_rca64_pg_fa7_xor0), .pg_fa_and0(u_pg_rca64_pg_fa7_and0), .pg_fa_xor1(u_pg_rca64_pg_fa7_xor1));
  and_gate and_gate_u_pg_rca64_and7(.a(u_pg_rca64_or6[0]), .b(u_pg_rca64_pg_fa7_xor0[0]), .out(u_pg_rca64_and7));
  or_gate or_gate_u_pg_rca64_or7(.a(u_pg_rca64_and7[0]), .b(u_pg_rca64_pg_fa7_and0[0]), .out(u_pg_rca64_or7));
  pg_fa pg_fa_u_pg_rca64_pg_fa8_out(.a(a[8]), .b(b[8]), .cin(u_pg_rca64_or7[0]), .pg_fa_xor0(u_pg_rca64_pg_fa8_xor0), .pg_fa_and0(u_pg_rca64_pg_fa8_and0), .pg_fa_xor1(u_pg_rca64_pg_fa8_xor1));
  and_gate and_gate_u_pg_rca64_and8(.a(u_pg_rca64_or7[0]), .b(u_pg_rca64_pg_fa8_xor0[0]), .out(u_pg_rca64_and8));
  or_gate or_gate_u_pg_rca64_or8(.a(u_pg_rca64_and8[0]), .b(u_pg_rca64_pg_fa8_and0[0]), .out(u_pg_rca64_or8));
  pg_fa pg_fa_u_pg_rca64_pg_fa9_out(.a(a[9]), .b(b[9]), .cin(u_pg_rca64_or8[0]), .pg_fa_xor0(u_pg_rca64_pg_fa9_xor0), .pg_fa_and0(u_pg_rca64_pg_fa9_and0), .pg_fa_xor1(u_pg_rca64_pg_fa9_xor1));
  and_gate and_gate_u_pg_rca64_and9(.a(u_pg_rca64_or8[0]), .b(u_pg_rca64_pg_fa9_xor0[0]), .out(u_pg_rca64_and9));
  or_gate or_gate_u_pg_rca64_or9(.a(u_pg_rca64_and9[0]), .b(u_pg_rca64_pg_fa9_and0[0]), .out(u_pg_rca64_or9));
  pg_fa pg_fa_u_pg_rca64_pg_fa10_out(.a(a[10]), .b(b[10]), .cin(u_pg_rca64_or9[0]), .pg_fa_xor0(u_pg_rca64_pg_fa10_xor0), .pg_fa_and0(u_pg_rca64_pg_fa10_and0), .pg_fa_xor1(u_pg_rca64_pg_fa10_xor1));
  and_gate and_gate_u_pg_rca64_and10(.a(u_pg_rca64_or9[0]), .b(u_pg_rca64_pg_fa10_xor0[0]), .out(u_pg_rca64_and10));
  or_gate or_gate_u_pg_rca64_or10(.a(u_pg_rca64_and10[0]), .b(u_pg_rca64_pg_fa10_and0[0]), .out(u_pg_rca64_or10));
  pg_fa pg_fa_u_pg_rca64_pg_fa11_out(.a(a[11]), .b(b[11]), .cin(u_pg_rca64_or10[0]), .pg_fa_xor0(u_pg_rca64_pg_fa11_xor0), .pg_fa_and0(u_pg_rca64_pg_fa11_and0), .pg_fa_xor1(u_pg_rca64_pg_fa11_xor1));
  and_gate and_gate_u_pg_rca64_and11(.a(u_pg_rca64_or10[0]), .b(u_pg_rca64_pg_fa11_xor0[0]), .out(u_pg_rca64_and11));
  or_gate or_gate_u_pg_rca64_or11(.a(u_pg_rca64_and11[0]), .b(u_pg_rca64_pg_fa11_and0[0]), .out(u_pg_rca64_or11));
  pg_fa pg_fa_u_pg_rca64_pg_fa12_out(.a(a[12]), .b(b[12]), .cin(u_pg_rca64_or11[0]), .pg_fa_xor0(u_pg_rca64_pg_fa12_xor0), .pg_fa_and0(u_pg_rca64_pg_fa12_and0), .pg_fa_xor1(u_pg_rca64_pg_fa12_xor1));
  and_gate and_gate_u_pg_rca64_and12(.a(u_pg_rca64_or11[0]), .b(u_pg_rca64_pg_fa12_xor0[0]), .out(u_pg_rca64_and12));
  or_gate or_gate_u_pg_rca64_or12(.a(u_pg_rca64_and12[0]), .b(u_pg_rca64_pg_fa12_and0[0]), .out(u_pg_rca64_or12));
  pg_fa pg_fa_u_pg_rca64_pg_fa13_out(.a(a[13]), .b(b[13]), .cin(u_pg_rca64_or12[0]), .pg_fa_xor0(u_pg_rca64_pg_fa13_xor0), .pg_fa_and0(u_pg_rca64_pg_fa13_and0), .pg_fa_xor1(u_pg_rca64_pg_fa13_xor1));
  and_gate and_gate_u_pg_rca64_and13(.a(u_pg_rca64_or12[0]), .b(u_pg_rca64_pg_fa13_xor0[0]), .out(u_pg_rca64_and13));
  or_gate or_gate_u_pg_rca64_or13(.a(u_pg_rca64_and13[0]), .b(u_pg_rca64_pg_fa13_and0[0]), .out(u_pg_rca64_or13));
  pg_fa pg_fa_u_pg_rca64_pg_fa14_out(.a(a[14]), .b(b[14]), .cin(u_pg_rca64_or13[0]), .pg_fa_xor0(u_pg_rca64_pg_fa14_xor0), .pg_fa_and0(u_pg_rca64_pg_fa14_and0), .pg_fa_xor1(u_pg_rca64_pg_fa14_xor1));
  and_gate and_gate_u_pg_rca64_and14(.a(u_pg_rca64_or13[0]), .b(u_pg_rca64_pg_fa14_xor0[0]), .out(u_pg_rca64_and14));
  or_gate or_gate_u_pg_rca64_or14(.a(u_pg_rca64_and14[0]), .b(u_pg_rca64_pg_fa14_and0[0]), .out(u_pg_rca64_or14));
  pg_fa pg_fa_u_pg_rca64_pg_fa15_out(.a(a[15]), .b(b[15]), .cin(u_pg_rca64_or14[0]), .pg_fa_xor0(u_pg_rca64_pg_fa15_xor0), .pg_fa_and0(u_pg_rca64_pg_fa15_and0), .pg_fa_xor1(u_pg_rca64_pg_fa15_xor1));
  and_gate and_gate_u_pg_rca64_and15(.a(u_pg_rca64_or14[0]), .b(u_pg_rca64_pg_fa15_xor0[0]), .out(u_pg_rca64_and15));
  or_gate or_gate_u_pg_rca64_or15(.a(u_pg_rca64_and15[0]), .b(u_pg_rca64_pg_fa15_and0[0]), .out(u_pg_rca64_or15));
  pg_fa pg_fa_u_pg_rca64_pg_fa16_out(.a(a[16]), .b(b[16]), .cin(u_pg_rca64_or15[0]), .pg_fa_xor0(u_pg_rca64_pg_fa16_xor0), .pg_fa_and0(u_pg_rca64_pg_fa16_and0), .pg_fa_xor1(u_pg_rca64_pg_fa16_xor1));
  and_gate and_gate_u_pg_rca64_and16(.a(u_pg_rca64_or15[0]), .b(u_pg_rca64_pg_fa16_xor0[0]), .out(u_pg_rca64_and16));
  or_gate or_gate_u_pg_rca64_or16(.a(u_pg_rca64_and16[0]), .b(u_pg_rca64_pg_fa16_and0[0]), .out(u_pg_rca64_or16));
  pg_fa pg_fa_u_pg_rca64_pg_fa17_out(.a(a[17]), .b(b[17]), .cin(u_pg_rca64_or16[0]), .pg_fa_xor0(u_pg_rca64_pg_fa17_xor0), .pg_fa_and0(u_pg_rca64_pg_fa17_and0), .pg_fa_xor1(u_pg_rca64_pg_fa17_xor1));
  and_gate and_gate_u_pg_rca64_and17(.a(u_pg_rca64_or16[0]), .b(u_pg_rca64_pg_fa17_xor0[0]), .out(u_pg_rca64_and17));
  or_gate or_gate_u_pg_rca64_or17(.a(u_pg_rca64_and17[0]), .b(u_pg_rca64_pg_fa17_and0[0]), .out(u_pg_rca64_or17));
  pg_fa pg_fa_u_pg_rca64_pg_fa18_out(.a(a[18]), .b(b[18]), .cin(u_pg_rca64_or17[0]), .pg_fa_xor0(u_pg_rca64_pg_fa18_xor0), .pg_fa_and0(u_pg_rca64_pg_fa18_and0), .pg_fa_xor1(u_pg_rca64_pg_fa18_xor1));
  and_gate and_gate_u_pg_rca64_and18(.a(u_pg_rca64_or17[0]), .b(u_pg_rca64_pg_fa18_xor0[0]), .out(u_pg_rca64_and18));
  or_gate or_gate_u_pg_rca64_or18(.a(u_pg_rca64_and18[0]), .b(u_pg_rca64_pg_fa18_and0[0]), .out(u_pg_rca64_or18));
  pg_fa pg_fa_u_pg_rca64_pg_fa19_out(.a(a[19]), .b(b[19]), .cin(u_pg_rca64_or18[0]), .pg_fa_xor0(u_pg_rca64_pg_fa19_xor0), .pg_fa_and0(u_pg_rca64_pg_fa19_and0), .pg_fa_xor1(u_pg_rca64_pg_fa19_xor1));
  and_gate and_gate_u_pg_rca64_and19(.a(u_pg_rca64_or18[0]), .b(u_pg_rca64_pg_fa19_xor0[0]), .out(u_pg_rca64_and19));
  or_gate or_gate_u_pg_rca64_or19(.a(u_pg_rca64_and19[0]), .b(u_pg_rca64_pg_fa19_and0[0]), .out(u_pg_rca64_or19));
  pg_fa pg_fa_u_pg_rca64_pg_fa20_out(.a(a[20]), .b(b[20]), .cin(u_pg_rca64_or19[0]), .pg_fa_xor0(u_pg_rca64_pg_fa20_xor0), .pg_fa_and0(u_pg_rca64_pg_fa20_and0), .pg_fa_xor1(u_pg_rca64_pg_fa20_xor1));
  and_gate and_gate_u_pg_rca64_and20(.a(u_pg_rca64_or19[0]), .b(u_pg_rca64_pg_fa20_xor0[0]), .out(u_pg_rca64_and20));
  or_gate or_gate_u_pg_rca64_or20(.a(u_pg_rca64_and20[0]), .b(u_pg_rca64_pg_fa20_and0[0]), .out(u_pg_rca64_or20));
  pg_fa pg_fa_u_pg_rca64_pg_fa21_out(.a(a[21]), .b(b[21]), .cin(u_pg_rca64_or20[0]), .pg_fa_xor0(u_pg_rca64_pg_fa21_xor0), .pg_fa_and0(u_pg_rca64_pg_fa21_and0), .pg_fa_xor1(u_pg_rca64_pg_fa21_xor1));
  and_gate and_gate_u_pg_rca64_and21(.a(u_pg_rca64_or20[0]), .b(u_pg_rca64_pg_fa21_xor0[0]), .out(u_pg_rca64_and21));
  or_gate or_gate_u_pg_rca64_or21(.a(u_pg_rca64_and21[0]), .b(u_pg_rca64_pg_fa21_and0[0]), .out(u_pg_rca64_or21));
  pg_fa pg_fa_u_pg_rca64_pg_fa22_out(.a(a[22]), .b(b[22]), .cin(u_pg_rca64_or21[0]), .pg_fa_xor0(u_pg_rca64_pg_fa22_xor0), .pg_fa_and0(u_pg_rca64_pg_fa22_and0), .pg_fa_xor1(u_pg_rca64_pg_fa22_xor1));
  and_gate and_gate_u_pg_rca64_and22(.a(u_pg_rca64_or21[0]), .b(u_pg_rca64_pg_fa22_xor0[0]), .out(u_pg_rca64_and22));
  or_gate or_gate_u_pg_rca64_or22(.a(u_pg_rca64_and22[0]), .b(u_pg_rca64_pg_fa22_and0[0]), .out(u_pg_rca64_or22));
  pg_fa pg_fa_u_pg_rca64_pg_fa23_out(.a(a[23]), .b(b[23]), .cin(u_pg_rca64_or22[0]), .pg_fa_xor0(u_pg_rca64_pg_fa23_xor0), .pg_fa_and0(u_pg_rca64_pg_fa23_and0), .pg_fa_xor1(u_pg_rca64_pg_fa23_xor1));
  and_gate and_gate_u_pg_rca64_and23(.a(u_pg_rca64_or22[0]), .b(u_pg_rca64_pg_fa23_xor0[0]), .out(u_pg_rca64_and23));
  or_gate or_gate_u_pg_rca64_or23(.a(u_pg_rca64_and23[0]), .b(u_pg_rca64_pg_fa23_and0[0]), .out(u_pg_rca64_or23));
  pg_fa pg_fa_u_pg_rca64_pg_fa24_out(.a(a[24]), .b(b[24]), .cin(u_pg_rca64_or23[0]), .pg_fa_xor0(u_pg_rca64_pg_fa24_xor0), .pg_fa_and0(u_pg_rca64_pg_fa24_and0), .pg_fa_xor1(u_pg_rca64_pg_fa24_xor1));
  and_gate and_gate_u_pg_rca64_and24(.a(u_pg_rca64_or23[0]), .b(u_pg_rca64_pg_fa24_xor0[0]), .out(u_pg_rca64_and24));
  or_gate or_gate_u_pg_rca64_or24(.a(u_pg_rca64_and24[0]), .b(u_pg_rca64_pg_fa24_and0[0]), .out(u_pg_rca64_or24));
  pg_fa pg_fa_u_pg_rca64_pg_fa25_out(.a(a[25]), .b(b[25]), .cin(u_pg_rca64_or24[0]), .pg_fa_xor0(u_pg_rca64_pg_fa25_xor0), .pg_fa_and0(u_pg_rca64_pg_fa25_and0), .pg_fa_xor1(u_pg_rca64_pg_fa25_xor1));
  and_gate and_gate_u_pg_rca64_and25(.a(u_pg_rca64_or24[0]), .b(u_pg_rca64_pg_fa25_xor0[0]), .out(u_pg_rca64_and25));
  or_gate or_gate_u_pg_rca64_or25(.a(u_pg_rca64_and25[0]), .b(u_pg_rca64_pg_fa25_and0[0]), .out(u_pg_rca64_or25));
  pg_fa pg_fa_u_pg_rca64_pg_fa26_out(.a(a[26]), .b(b[26]), .cin(u_pg_rca64_or25[0]), .pg_fa_xor0(u_pg_rca64_pg_fa26_xor0), .pg_fa_and0(u_pg_rca64_pg_fa26_and0), .pg_fa_xor1(u_pg_rca64_pg_fa26_xor1));
  and_gate and_gate_u_pg_rca64_and26(.a(u_pg_rca64_or25[0]), .b(u_pg_rca64_pg_fa26_xor0[0]), .out(u_pg_rca64_and26));
  or_gate or_gate_u_pg_rca64_or26(.a(u_pg_rca64_and26[0]), .b(u_pg_rca64_pg_fa26_and0[0]), .out(u_pg_rca64_or26));
  pg_fa pg_fa_u_pg_rca64_pg_fa27_out(.a(a[27]), .b(b[27]), .cin(u_pg_rca64_or26[0]), .pg_fa_xor0(u_pg_rca64_pg_fa27_xor0), .pg_fa_and0(u_pg_rca64_pg_fa27_and0), .pg_fa_xor1(u_pg_rca64_pg_fa27_xor1));
  and_gate and_gate_u_pg_rca64_and27(.a(u_pg_rca64_or26[0]), .b(u_pg_rca64_pg_fa27_xor0[0]), .out(u_pg_rca64_and27));
  or_gate or_gate_u_pg_rca64_or27(.a(u_pg_rca64_and27[0]), .b(u_pg_rca64_pg_fa27_and0[0]), .out(u_pg_rca64_or27));
  pg_fa pg_fa_u_pg_rca64_pg_fa28_out(.a(a[28]), .b(b[28]), .cin(u_pg_rca64_or27[0]), .pg_fa_xor0(u_pg_rca64_pg_fa28_xor0), .pg_fa_and0(u_pg_rca64_pg_fa28_and0), .pg_fa_xor1(u_pg_rca64_pg_fa28_xor1));
  and_gate and_gate_u_pg_rca64_and28(.a(u_pg_rca64_or27[0]), .b(u_pg_rca64_pg_fa28_xor0[0]), .out(u_pg_rca64_and28));
  or_gate or_gate_u_pg_rca64_or28(.a(u_pg_rca64_and28[0]), .b(u_pg_rca64_pg_fa28_and0[0]), .out(u_pg_rca64_or28));
  pg_fa pg_fa_u_pg_rca64_pg_fa29_out(.a(a[29]), .b(b[29]), .cin(u_pg_rca64_or28[0]), .pg_fa_xor0(u_pg_rca64_pg_fa29_xor0), .pg_fa_and0(u_pg_rca64_pg_fa29_and0), .pg_fa_xor1(u_pg_rca64_pg_fa29_xor1));
  and_gate and_gate_u_pg_rca64_and29(.a(u_pg_rca64_or28[0]), .b(u_pg_rca64_pg_fa29_xor0[0]), .out(u_pg_rca64_and29));
  or_gate or_gate_u_pg_rca64_or29(.a(u_pg_rca64_and29[0]), .b(u_pg_rca64_pg_fa29_and0[0]), .out(u_pg_rca64_or29));
  pg_fa pg_fa_u_pg_rca64_pg_fa30_out(.a(a[30]), .b(b[30]), .cin(u_pg_rca64_or29[0]), .pg_fa_xor0(u_pg_rca64_pg_fa30_xor0), .pg_fa_and0(u_pg_rca64_pg_fa30_and0), .pg_fa_xor1(u_pg_rca64_pg_fa30_xor1));
  and_gate and_gate_u_pg_rca64_and30(.a(u_pg_rca64_or29[0]), .b(u_pg_rca64_pg_fa30_xor0[0]), .out(u_pg_rca64_and30));
  or_gate or_gate_u_pg_rca64_or30(.a(u_pg_rca64_and30[0]), .b(u_pg_rca64_pg_fa30_and0[0]), .out(u_pg_rca64_or30));
  pg_fa pg_fa_u_pg_rca64_pg_fa31_out(.a(a[31]), .b(b[31]), .cin(u_pg_rca64_or30[0]), .pg_fa_xor0(u_pg_rca64_pg_fa31_xor0), .pg_fa_and0(u_pg_rca64_pg_fa31_and0), .pg_fa_xor1(u_pg_rca64_pg_fa31_xor1));
  and_gate and_gate_u_pg_rca64_and31(.a(u_pg_rca64_or30[0]), .b(u_pg_rca64_pg_fa31_xor0[0]), .out(u_pg_rca64_and31));
  or_gate or_gate_u_pg_rca64_or31(.a(u_pg_rca64_and31[0]), .b(u_pg_rca64_pg_fa31_and0[0]), .out(u_pg_rca64_or31));
  pg_fa pg_fa_u_pg_rca64_pg_fa32_out(.a(a[32]), .b(b[32]), .cin(u_pg_rca64_or31[0]), .pg_fa_xor0(u_pg_rca64_pg_fa32_xor0), .pg_fa_and0(u_pg_rca64_pg_fa32_and0), .pg_fa_xor1(u_pg_rca64_pg_fa32_xor1));
  and_gate and_gate_u_pg_rca64_and32(.a(u_pg_rca64_or31[0]), .b(u_pg_rca64_pg_fa32_xor0[0]), .out(u_pg_rca64_and32));
  or_gate or_gate_u_pg_rca64_or32(.a(u_pg_rca64_and32[0]), .b(u_pg_rca64_pg_fa32_and0[0]), .out(u_pg_rca64_or32));
  pg_fa pg_fa_u_pg_rca64_pg_fa33_out(.a(a[33]), .b(b[33]), .cin(u_pg_rca64_or32[0]), .pg_fa_xor0(u_pg_rca64_pg_fa33_xor0), .pg_fa_and0(u_pg_rca64_pg_fa33_and0), .pg_fa_xor1(u_pg_rca64_pg_fa33_xor1));
  and_gate and_gate_u_pg_rca64_and33(.a(u_pg_rca64_or32[0]), .b(u_pg_rca64_pg_fa33_xor0[0]), .out(u_pg_rca64_and33));
  or_gate or_gate_u_pg_rca64_or33(.a(u_pg_rca64_and33[0]), .b(u_pg_rca64_pg_fa33_and0[0]), .out(u_pg_rca64_or33));
  pg_fa pg_fa_u_pg_rca64_pg_fa34_out(.a(a[34]), .b(b[34]), .cin(u_pg_rca64_or33[0]), .pg_fa_xor0(u_pg_rca64_pg_fa34_xor0), .pg_fa_and0(u_pg_rca64_pg_fa34_and0), .pg_fa_xor1(u_pg_rca64_pg_fa34_xor1));
  and_gate and_gate_u_pg_rca64_and34(.a(u_pg_rca64_or33[0]), .b(u_pg_rca64_pg_fa34_xor0[0]), .out(u_pg_rca64_and34));
  or_gate or_gate_u_pg_rca64_or34(.a(u_pg_rca64_and34[0]), .b(u_pg_rca64_pg_fa34_and0[0]), .out(u_pg_rca64_or34));
  pg_fa pg_fa_u_pg_rca64_pg_fa35_out(.a(a[35]), .b(b[35]), .cin(u_pg_rca64_or34[0]), .pg_fa_xor0(u_pg_rca64_pg_fa35_xor0), .pg_fa_and0(u_pg_rca64_pg_fa35_and0), .pg_fa_xor1(u_pg_rca64_pg_fa35_xor1));
  and_gate and_gate_u_pg_rca64_and35(.a(u_pg_rca64_or34[0]), .b(u_pg_rca64_pg_fa35_xor0[0]), .out(u_pg_rca64_and35));
  or_gate or_gate_u_pg_rca64_or35(.a(u_pg_rca64_and35[0]), .b(u_pg_rca64_pg_fa35_and0[0]), .out(u_pg_rca64_or35));
  pg_fa pg_fa_u_pg_rca64_pg_fa36_out(.a(a[36]), .b(b[36]), .cin(u_pg_rca64_or35[0]), .pg_fa_xor0(u_pg_rca64_pg_fa36_xor0), .pg_fa_and0(u_pg_rca64_pg_fa36_and0), .pg_fa_xor1(u_pg_rca64_pg_fa36_xor1));
  and_gate and_gate_u_pg_rca64_and36(.a(u_pg_rca64_or35[0]), .b(u_pg_rca64_pg_fa36_xor0[0]), .out(u_pg_rca64_and36));
  or_gate or_gate_u_pg_rca64_or36(.a(u_pg_rca64_and36[0]), .b(u_pg_rca64_pg_fa36_and0[0]), .out(u_pg_rca64_or36));
  pg_fa pg_fa_u_pg_rca64_pg_fa37_out(.a(a[37]), .b(b[37]), .cin(u_pg_rca64_or36[0]), .pg_fa_xor0(u_pg_rca64_pg_fa37_xor0), .pg_fa_and0(u_pg_rca64_pg_fa37_and0), .pg_fa_xor1(u_pg_rca64_pg_fa37_xor1));
  and_gate and_gate_u_pg_rca64_and37(.a(u_pg_rca64_or36[0]), .b(u_pg_rca64_pg_fa37_xor0[0]), .out(u_pg_rca64_and37));
  or_gate or_gate_u_pg_rca64_or37(.a(u_pg_rca64_and37[0]), .b(u_pg_rca64_pg_fa37_and0[0]), .out(u_pg_rca64_or37));
  pg_fa pg_fa_u_pg_rca64_pg_fa38_out(.a(a[38]), .b(b[38]), .cin(u_pg_rca64_or37[0]), .pg_fa_xor0(u_pg_rca64_pg_fa38_xor0), .pg_fa_and0(u_pg_rca64_pg_fa38_and0), .pg_fa_xor1(u_pg_rca64_pg_fa38_xor1));
  and_gate and_gate_u_pg_rca64_and38(.a(u_pg_rca64_or37[0]), .b(u_pg_rca64_pg_fa38_xor0[0]), .out(u_pg_rca64_and38));
  or_gate or_gate_u_pg_rca64_or38(.a(u_pg_rca64_and38[0]), .b(u_pg_rca64_pg_fa38_and0[0]), .out(u_pg_rca64_or38));
  pg_fa pg_fa_u_pg_rca64_pg_fa39_out(.a(a[39]), .b(b[39]), .cin(u_pg_rca64_or38[0]), .pg_fa_xor0(u_pg_rca64_pg_fa39_xor0), .pg_fa_and0(u_pg_rca64_pg_fa39_and0), .pg_fa_xor1(u_pg_rca64_pg_fa39_xor1));
  and_gate and_gate_u_pg_rca64_and39(.a(u_pg_rca64_or38[0]), .b(u_pg_rca64_pg_fa39_xor0[0]), .out(u_pg_rca64_and39));
  or_gate or_gate_u_pg_rca64_or39(.a(u_pg_rca64_and39[0]), .b(u_pg_rca64_pg_fa39_and0[0]), .out(u_pg_rca64_or39));
  pg_fa pg_fa_u_pg_rca64_pg_fa40_out(.a(a[40]), .b(b[40]), .cin(u_pg_rca64_or39[0]), .pg_fa_xor0(u_pg_rca64_pg_fa40_xor0), .pg_fa_and0(u_pg_rca64_pg_fa40_and0), .pg_fa_xor1(u_pg_rca64_pg_fa40_xor1));
  and_gate and_gate_u_pg_rca64_and40(.a(u_pg_rca64_or39[0]), .b(u_pg_rca64_pg_fa40_xor0[0]), .out(u_pg_rca64_and40));
  or_gate or_gate_u_pg_rca64_or40(.a(u_pg_rca64_and40[0]), .b(u_pg_rca64_pg_fa40_and0[0]), .out(u_pg_rca64_or40));
  pg_fa pg_fa_u_pg_rca64_pg_fa41_out(.a(a[41]), .b(b[41]), .cin(u_pg_rca64_or40[0]), .pg_fa_xor0(u_pg_rca64_pg_fa41_xor0), .pg_fa_and0(u_pg_rca64_pg_fa41_and0), .pg_fa_xor1(u_pg_rca64_pg_fa41_xor1));
  and_gate and_gate_u_pg_rca64_and41(.a(u_pg_rca64_or40[0]), .b(u_pg_rca64_pg_fa41_xor0[0]), .out(u_pg_rca64_and41));
  or_gate or_gate_u_pg_rca64_or41(.a(u_pg_rca64_and41[0]), .b(u_pg_rca64_pg_fa41_and0[0]), .out(u_pg_rca64_or41));
  pg_fa pg_fa_u_pg_rca64_pg_fa42_out(.a(a[42]), .b(b[42]), .cin(u_pg_rca64_or41[0]), .pg_fa_xor0(u_pg_rca64_pg_fa42_xor0), .pg_fa_and0(u_pg_rca64_pg_fa42_and0), .pg_fa_xor1(u_pg_rca64_pg_fa42_xor1));
  and_gate and_gate_u_pg_rca64_and42(.a(u_pg_rca64_or41[0]), .b(u_pg_rca64_pg_fa42_xor0[0]), .out(u_pg_rca64_and42));
  or_gate or_gate_u_pg_rca64_or42(.a(u_pg_rca64_and42[0]), .b(u_pg_rca64_pg_fa42_and0[0]), .out(u_pg_rca64_or42));
  pg_fa pg_fa_u_pg_rca64_pg_fa43_out(.a(a[43]), .b(b[43]), .cin(u_pg_rca64_or42[0]), .pg_fa_xor0(u_pg_rca64_pg_fa43_xor0), .pg_fa_and0(u_pg_rca64_pg_fa43_and0), .pg_fa_xor1(u_pg_rca64_pg_fa43_xor1));
  and_gate and_gate_u_pg_rca64_and43(.a(u_pg_rca64_or42[0]), .b(u_pg_rca64_pg_fa43_xor0[0]), .out(u_pg_rca64_and43));
  or_gate or_gate_u_pg_rca64_or43(.a(u_pg_rca64_and43[0]), .b(u_pg_rca64_pg_fa43_and0[0]), .out(u_pg_rca64_or43));
  pg_fa pg_fa_u_pg_rca64_pg_fa44_out(.a(a[44]), .b(b[44]), .cin(u_pg_rca64_or43[0]), .pg_fa_xor0(u_pg_rca64_pg_fa44_xor0), .pg_fa_and0(u_pg_rca64_pg_fa44_and0), .pg_fa_xor1(u_pg_rca64_pg_fa44_xor1));
  and_gate and_gate_u_pg_rca64_and44(.a(u_pg_rca64_or43[0]), .b(u_pg_rca64_pg_fa44_xor0[0]), .out(u_pg_rca64_and44));
  or_gate or_gate_u_pg_rca64_or44(.a(u_pg_rca64_and44[0]), .b(u_pg_rca64_pg_fa44_and0[0]), .out(u_pg_rca64_or44));
  pg_fa pg_fa_u_pg_rca64_pg_fa45_out(.a(a[45]), .b(b[45]), .cin(u_pg_rca64_or44[0]), .pg_fa_xor0(u_pg_rca64_pg_fa45_xor0), .pg_fa_and0(u_pg_rca64_pg_fa45_and0), .pg_fa_xor1(u_pg_rca64_pg_fa45_xor1));
  and_gate and_gate_u_pg_rca64_and45(.a(u_pg_rca64_or44[0]), .b(u_pg_rca64_pg_fa45_xor0[0]), .out(u_pg_rca64_and45));
  or_gate or_gate_u_pg_rca64_or45(.a(u_pg_rca64_and45[0]), .b(u_pg_rca64_pg_fa45_and0[0]), .out(u_pg_rca64_or45));
  pg_fa pg_fa_u_pg_rca64_pg_fa46_out(.a(a[46]), .b(b[46]), .cin(u_pg_rca64_or45[0]), .pg_fa_xor0(u_pg_rca64_pg_fa46_xor0), .pg_fa_and0(u_pg_rca64_pg_fa46_and0), .pg_fa_xor1(u_pg_rca64_pg_fa46_xor1));
  and_gate and_gate_u_pg_rca64_and46(.a(u_pg_rca64_or45[0]), .b(u_pg_rca64_pg_fa46_xor0[0]), .out(u_pg_rca64_and46));
  or_gate or_gate_u_pg_rca64_or46(.a(u_pg_rca64_and46[0]), .b(u_pg_rca64_pg_fa46_and0[0]), .out(u_pg_rca64_or46));
  pg_fa pg_fa_u_pg_rca64_pg_fa47_out(.a(a[47]), .b(b[47]), .cin(u_pg_rca64_or46[0]), .pg_fa_xor0(u_pg_rca64_pg_fa47_xor0), .pg_fa_and0(u_pg_rca64_pg_fa47_and0), .pg_fa_xor1(u_pg_rca64_pg_fa47_xor1));
  and_gate and_gate_u_pg_rca64_and47(.a(u_pg_rca64_or46[0]), .b(u_pg_rca64_pg_fa47_xor0[0]), .out(u_pg_rca64_and47));
  or_gate or_gate_u_pg_rca64_or47(.a(u_pg_rca64_and47[0]), .b(u_pg_rca64_pg_fa47_and0[0]), .out(u_pg_rca64_or47));
  pg_fa pg_fa_u_pg_rca64_pg_fa48_out(.a(a[48]), .b(b[48]), .cin(u_pg_rca64_or47[0]), .pg_fa_xor0(u_pg_rca64_pg_fa48_xor0), .pg_fa_and0(u_pg_rca64_pg_fa48_and0), .pg_fa_xor1(u_pg_rca64_pg_fa48_xor1));
  and_gate and_gate_u_pg_rca64_and48(.a(u_pg_rca64_or47[0]), .b(u_pg_rca64_pg_fa48_xor0[0]), .out(u_pg_rca64_and48));
  or_gate or_gate_u_pg_rca64_or48(.a(u_pg_rca64_and48[0]), .b(u_pg_rca64_pg_fa48_and0[0]), .out(u_pg_rca64_or48));
  pg_fa pg_fa_u_pg_rca64_pg_fa49_out(.a(a[49]), .b(b[49]), .cin(u_pg_rca64_or48[0]), .pg_fa_xor0(u_pg_rca64_pg_fa49_xor0), .pg_fa_and0(u_pg_rca64_pg_fa49_and0), .pg_fa_xor1(u_pg_rca64_pg_fa49_xor1));
  and_gate and_gate_u_pg_rca64_and49(.a(u_pg_rca64_or48[0]), .b(u_pg_rca64_pg_fa49_xor0[0]), .out(u_pg_rca64_and49));
  or_gate or_gate_u_pg_rca64_or49(.a(u_pg_rca64_and49[0]), .b(u_pg_rca64_pg_fa49_and0[0]), .out(u_pg_rca64_or49));
  pg_fa pg_fa_u_pg_rca64_pg_fa50_out(.a(a[50]), .b(b[50]), .cin(u_pg_rca64_or49[0]), .pg_fa_xor0(u_pg_rca64_pg_fa50_xor0), .pg_fa_and0(u_pg_rca64_pg_fa50_and0), .pg_fa_xor1(u_pg_rca64_pg_fa50_xor1));
  and_gate and_gate_u_pg_rca64_and50(.a(u_pg_rca64_or49[0]), .b(u_pg_rca64_pg_fa50_xor0[0]), .out(u_pg_rca64_and50));
  or_gate or_gate_u_pg_rca64_or50(.a(u_pg_rca64_and50[0]), .b(u_pg_rca64_pg_fa50_and0[0]), .out(u_pg_rca64_or50));
  pg_fa pg_fa_u_pg_rca64_pg_fa51_out(.a(a[51]), .b(b[51]), .cin(u_pg_rca64_or50[0]), .pg_fa_xor0(u_pg_rca64_pg_fa51_xor0), .pg_fa_and0(u_pg_rca64_pg_fa51_and0), .pg_fa_xor1(u_pg_rca64_pg_fa51_xor1));
  and_gate and_gate_u_pg_rca64_and51(.a(u_pg_rca64_or50[0]), .b(u_pg_rca64_pg_fa51_xor0[0]), .out(u_pg_rca64_and51));
  or_gate or_gate_u_pg_rca64_or51(.a(u_pg_rca64_and51[0]), .b(u_pg_rca64_pg_fa51_and0[0]), .out(u_pg_rca64_or51));
  pg_fa pg_fa_u_pg_rca64_pg_fa52_out(.a(a[52]), .b(b[52]), .cin(u_pg_rca64_or51[0]), .pg_fa_xor0(u_pg_rca64_pg_fa52_xor0), .pg_fa_and0(u_pg_rca64_pg_fa52_and0), .pg_fa_xor1(u_pg_rca64_pg_fa52_xor1));
  and_gate and_gate_u_pg_rca64_and52(.a(u_pg_rca64_or51[0]), .b(u_pg_rca64_pg_fa52_xor0[0]), .out(u_pg_rca64_and52));
  or_gate or_gate_u_pg_rca64_or52(.a(u_pg_rca64_and52[0]), .b(u_pg_rca64_pg_fa52_and0[0]), .out(u_pg_rca64_or52));
  pg_fa pg_fa_u_pg_rca64_pg_fa53_out(.a(a[53]), .b(b[53]), .cin(u_pg_rca64_or52[0]), .pg_fa_xor0(u_pg_rca64_pg_fa53_xor0), .pg_fa_and0(u_pg_rca64_pg_fa53_and0), .pg_fa_xor1(u_pg_rca64_pg_fa53_xor1));
  and_gate and_gate_u_pg_rca64_and53(.a(u_pg_rca64_or52[0]), .b(u_pg_rca64_pg_fa53_xor0[0]), .out(u_pg_rca64_and53));
  or_gate or_gate_u_pg_rca64_or53(.a(u_pg_rca64_and53[0]), .b(u_pg_rca64_pg_fa53_and0[0]), .out(u_pg_rca64_or53));
  pg_fa pg_fa_u_pg_rca64_pg_fa54_out(.a(a[54]), .b(b[54]), .cin(u_pg_rca64_or53[0]), .pg_fa_xor0(u_pg_rca64_pg_fa54_xor0), .pg_fa_and0(u_pg_rca64_pg_fa54_and0), .pg_fa_xor1(u_pg_rca64_pg_fa54_xor1));
  and_gate and_gate_u_pg_rca64_and54(.a(u_pg_rca64_or53[0]), .b(u_pg_rca64_pg_fa54_xor0[0]), .out(u_pg_rca64_and54));
  or_gate or_gate_u_pg_rca64_or54(.a(u_pg_rca64_and54[0]), .b(u_pg_rca64_pg_fa54_and0[0]), .out(u_pg_rca64_or54));
  pg_fa pg_fa_u_pg_rca64_pg_fa55_out(.a(a[55]), .b(b[55]), .cin(u_pg_rca64_or54[0]), .pg_fa_xor0(u_pg_rca64_pg_fa55_xor0), .pg_fa_and0(u_pg_rca64_pg_fa55_and0), .pg_fa_xor1(u_pg_rca64_pg_fa55_xor1));
  and_gate and_gate_u_pg_rca64_and55(.a(u_pg_rca64_or54[0]), .b(u_pg_rca64_pg_fa55_xor0[0]), .out(u_pg_rca64_and55));
  or_gate or_gate_u_pg_rca64_or55(.a(u_pg_rca64_and55[0]), .b(u_pg_rca64_pg_fa55_and0[0]), .out(u_pg_rca64_or55));
  pg_fa pg_fa_u_pg_rca64_pg_fa56_out(.a(a[56]), .b(b[56]), .cin(u_pg_rca64_or55[0]), .pg_fa_xor0(u_pg_rca64_pg_fa56_xor0), .pg_fa_and0(u_pg_rca64_pg_fa56_and0), .pg_fa_xor1(u_pg_rca64_pg_fa56_xor1));
  and_gate and_gate_u_pg_rca64_and56(.a(u_pg_rca64_or55[0]), .b(u_pg_rca64_pg_fa56_xor0[0]), .out(u_pg_rca64_and56));
  or_gate or_gate_u_pg_rca64_or56(.a(u_pg_rca64_and56[0]), .b(u_pg_rca64_pg_fa56_and0[0]), .out(u_pg_rca64_or56));
  pg_fa pg_fa_u_pg_rca64_pg_fa57_out(.a(a[57]), .b(b[57]), .cin(u_pg_rca64_or56[0]), .pg_fa_xor0(u_pg_rca64_pg_fa57_xor0), .pg_fa_and0(u_pg_rca64_pg_fa57_and0), .pg_fa_xor1(u_pg_rca64_pg_fa57_xor1));
  and_gate and_gate_u_pg_rca64_and57(.a(u_pg_rca64_or56[0]), .b(u_pg_rca64_pg_fa57_xor0[0]), .out(u_pg_rca64_and57));
  or_gate or_gate_u_pg_rca64_or57(.a(u_pg_rca64_and57[0]), .b(u_pg_rca64_pg_fa57_and0[0]), .out(u_pg_rca64_or57));
  pg_fa pg_fa_u_pg_rca64_pg_fa58_out(.a(a[58]), .b(b[58]), .cin(u_pg_rca64_or57[0]), .pg_fa_xor0(u_pg_rca64_pg_fa58_xor0), .pg_fa_and0(u_pg_rca64_pg_fa58_and0), .pg_fa_xor1(u_pg_rca64_pg_fa58_xor1));
  and_gate and_gate_u_pg_rca64_and58(.a(u_pg_rca64_or57[0]), .b(u_pg_rca64_pg_fa58_xor0[0]), .out(u_pg_rca64_and58));
  or_gate or_gate_u_pg_rca64_or58(.a(u_pg_rca64_and58[0]), .b(u_pg_rca64_pg_fa58_and0[0]), .out(u_pg_rca64_or58));
  pg_fa pg_fa_u_pg_rca64_pg_fa59_out(.a(a[59]), .b(b[59]), .cin(u_pg_rca64_or58[0]), .pg_fa_xor0(u_pg_rca64_pg_fa59_xor0), .pg_fa_and0(u_pg_rca64_pg_fa59_and0), .pg_fa_xor1(u_pg_rca64_pg_fa59_xor1));
  and_gate and_gate_u_pg_rca64_and59(.a(u_pg_rca64_or58[0]), .b(u_pg_rca64_pg_fa59_xor0[0]), .out(u_pg_rca64_and59));
  or_gate or_gate_u_pg_rca64_or59(.a(u_pg_rca64_and59[0]), .b(u_pg_rca64_pg_fa59_and0[0]), .out(u_pg_rca64_or59));
  pg_fa pg_fa_u_pg_rca64_pg_fa60_out(.a(a[60]), .b(b[60]), .cin(u_pg_rca64_or59[0]), .pg_fa_xor0(u_pg_rca64_pg_fa60_xor0), .pg_fa_and0(u_pg_rca64_pg_fa60_and0), .pg_fa_xor1(u_pg_rca64_pg_fa60_xor1));
  and_gate and_gate_u_pg_rca64_and60(.a(u_pg_rca64_or59[0]), .b(u_pg_rca64_pg_fa60_xor0[0]), .out(u_pg_rca64_and60));
  or_gate or_gate_u_pg_rca64_or60(.a(u_pg_rca64_and60[0]), .b(u_pg_rca64_pg_fa60_and0[0]), .out(u_pg_rca64_or60));
  pg_fa pg_fa_u_pg_rca64_pg_fa61_out(.a(a[61]), .b(b[61]), .cin(u_pg_rca64_or60[0]), .pg_fa_xor0(u_pg_rca64_pg_fa61_xor0), .pg_fa_and0(u_pg_rca64_pg_fa61_and0), .pg_fa_xor1(u_pg_rca64_pg_fa61_xor1));
  and_gate and_gate_u_pg_rca64_and61(.a(u_pg_rca64_or60[0]), .b(u_pg_rca64_pg_fa61_xor0[0]), .out(u_pg_rca64_and61));
  or_gate or_gate_u_pg_rca64_or61(.a(u_pg_rca64_and61[0]), .b(u_pg_rca64_pg_fa61_and0[0]), .out(u_pg_rca64_or61));
  pg_fa pg_fa_u_pg_rca64_pg_fa62_out(.a(a[62]), .b(b[62]), .cin(u_pg_rca64_or61[0]), .pg_fa_xor0(u_pg_rca64_pg_fa62_xor0), .pg_fa_and0(u_pg_rca64_pg_fa62_and0), .pg_fa_xor1(u_pg_rca64_pg_fa62_xor1));
  and_gate and_gate_u_pg_rca64_and62(.a(u_pg_rca64_or61[0]), .b(u_pg_rca64_pg_fa62_xor0[0]), .out(u_pg_rca64_and62));
  or_gate or_gate_u_pg_rca64_or62(.a(u_pg_rca64_and62[0]), .b(u_pg_rca64_pg_fa62_and0[0]), .out(u_pg_rca64_or62));
  pg_fa pg_fa_u_pg_rca64_pg_fa63_out(.a(a[63]), .b(b[63]), .cin(u_pg_rca64_or62[0]), .pg_fa_xor0(u_pg_rca64_pg_fa63_xor0), .pg_fa_and0(u_pg_rca64_pg_fa63_and0), .pg_fa_xor1(u_pg_rca64_pg_fa63_xor1));
  and_gate and_gate_u_pg_rca64_and63(.a(u_pg_rca64_or62[0]), .b(u_pg_rca64_pg_fa63_xor0[0]), .out(u_pg_rca64_and63));
  or_gate or_gate_u_pg_rca64_or63(.a(u_pg_rca64_and63[0]), .b(u_pg_rca64_pg_fa63_and0[0]), .out(u_pg_rca64_or63));

  assign u_pg_rca64_out[0] = u_pg_rca64_pg_fa0_xor0[0];
  assign u_pg_rca64_out[1] = u_pg_rca64_pg_fa1_xor1[0];
  assign u_pg_rca64_out[2] = u_pg_rca64_pg_fa2_xor1[0];
  assign u_pg_rca64_out[3] = u_pg_rca64_pg_fa3_xor1[0];
  assign u_pg_rca64_out[4] = u_pg_rca64_pg_fa4_xor1[0];
  assign u_pg_rca64_out[5] = u_pg_rca64_pg_fa5_xor1[0];
  assign u_pg_rca64_out[6] = u_pg_rca64_pg_fa6_xor1[0];
  assign u_pg_rca64_out[7] = u_pg_rca64_pg_fa7_xor1[0];
  assign u_pg_rca64_out[8] = u_pg_rca64_pg_fa8_xor1[0];
  assign u_pg_rca64_out[9] = u_pg_rca64_pg_fa9_xor1[0];
  assign u_pg_rca64_out[10] = u_pg_rca64_pg_fa10_xor1[0];
  assign u_pg_rca64_out[11] = u_pg_rca64_pg_fa11_xor1[0];
  assign u_pg_rca64_out[12] = u_pg_rca64_pg_fa12_xor1[0];
  assign u_pg_rca64_out[13] = u_pg_rca64_pg_fa13_xor1[0];
  assign u_pg_rca64_out[14] = u_pg_rca64_pg_fa14_xor1[0];
  assign u_pg_rca64_out[15] = u_pg_rca64_pg_fa15_xor1[0];
  assign u_pg_rca64_out[16] = u_pg_rca64_pg_fa16_xor1[0];
  assign u_pg_rca64_out[17] = u_pg_rca64_pg_fa17_xor1[0];
  assign u_pg_rca64_out[18] = u_pg_rca64_pg_fa18_xor1[0];
  assign u_pg_rca64_out[19] = u_pg_rca64_pg_fa19_xor1[0];
  assign u_pg_rca64_out[20] = u_pg_rca64_pg_fa20_xor1[0];
  assign u_pg_rca64_out[21] = u_pg_rca64_pg_fa21_xor1[0];
  assign u_pg_rca64_out[22] = u_pg_rca64_pg_fa22_xor1[0];
  assign u_pg_rca64_out[23] = u_pg_rca64_pg_fa23_xor1[0];
  assign u_pg_rca64_out[24] = u_pg_rca64_pg_fa24_xor1[0];
  assign u_pg_rca64_out[25] = u_pg_rca64_pg_fa25_xor1[0];
  assign u_pg_rca64_out[26] = u_pg_rca64_pg_fa26_xor1[0];
  assign u_pg_rca64_out[27] = u_pg_rca64_pg_fa27_xor1[0];
  assign u_pg_rca64_out[28] = u_pg_rca64_pg_fa28_xor1[0];
  assign u_pg_rca64_out[29] = u_pg_rca64_pg_fa29_xor1[0];
  assign u_pg_rca64_out[30] = u_pg_rca64_pg_fa30_xor1[0];
  assign u_pg_rca64_out[31] = u_pg_rca64_pg_fa31_xor1[0];
  assign u_pg_rca64_out[32] = u_pg_rca64_pg_fa32_xor1[0];
  assign u_pg_rca64_out[33] = u_pg_rca64_pg_fa33_xor1[0];
  assign u_pg_rca64_out[34] = u_pg_rca64_pg_fa34_xor1[0];
  assign u_pg_rca64_out[35] = u_pg_rca64_pg_fa35_xor1[0];
  assign u_pg_rca64_out[36] = u_pg_rca64_pg_fa36_xor1[0];
  assign u_pg_rca64_out[37] = u_pg_rca64_pg_fa37_xor1[0];
  assign u_pg_rca64_out[38] = u_pg_rca64_pg_fa38_xor1[0];
  assign u_pg_rca64_out[39] = u_pg_rca64_pg_fa39_xor1[0];
  assign u_pg_rca64_out[40] = u_pg_rca64_pg_fa40_xor1[0];
  assign u_pg_rca64_out[41] = u_pg_rca64_pg_fa41_xor1[0];
  assign u_pg_rca64_out[42] = u_pg_rca64_pg_fa42_xor1[0];
  assign u_pg_rca64_out[43] = u_pg_rca64_pg_fa43_xor1[0];
  assign u_pg_rca64_out[44] = u_pg_rca64_pg_fa44_xor1[0];
  assign u_pg_rca64_out[45] = u_pg_rca64_pg_fa45_xor1[0];
  assign u_pg_rca64_out[46] = u_pg_rca64_pg_fa46_xor1[0];
  assign u_pg_rca64_out[47] = u_pg_rca64_pg_fa47_xor1[0];
  assign u_pg_rca64_out[48] = u_pg_rca64_pg_fa48_xor1[0];
  assign u_pg_rca64_out[49] = u_pg_rca64_pg_fa49_xor1[0];
  assign u_pg_rca64_out[50] = u_pg_rca64_pg_fa50_xor1[0];
  assign u_pg_rca64_out[51] = u_pg_rca64_pg_fa51_xor1[0];
  assign u_pg_rca64_out[52] = u_pg_rca64_pg_fa52_xor1[0];
  assign u_pg_rca64_out[53] = u_pg_rca64_pg_fa53_xor1[0];
  assign u_pg_rca64_out[54] = u_pg_rca64_pg_fa54_xor1[0];
  assign u_pg_rca64_out[55] = u_pg_rca64_pg_fa55_xor1[0];
  assign u_pg_rca64_out[56] = u_pg_rca64_pg_fa56_xor1[0];
  assign u_pg_rca64_out[57] = u_pg_rca64_pg_fa57_xor1[0];
  assign u_pg_rca64_out[58] = u_pg_rca64_pg_fa58_xor1[0];
  assign u_pg_rca64_out[59] = u_pg_rca64_pg_fa59_xor1[0];
  assign u_pg_rca64_out[60] = u_pg_rca64_pg_fa60_xor1[0];
  assign u_pg_rca64_out[61] = u_pg_rca64_pg_fa61_xor1[0];
  assign u_pg_rca64_out[62] = u_pg_rca64_pg_fa62_xor1[0];
  assign u_pg_rca64_out[63] = u_pg_rca64_pg_fa63_xor1[0];
  assign u_pg_rca64_out[64] = u_pg_rca64_or63[0];
endmodule

module u_CSAwallace_pg_rca32(input [31:0] a, input [31:0] b, output [63:0] u_CSAwallace_pg_rca32_out);
  wire [0:0] u_CSAwallace_pg_rca32_and_0_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_0;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_1;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_2;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_3;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_4;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_5;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_6;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_7;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_8;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_9;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_10;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_11;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_12;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_13;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_14;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_15;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_16;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_17;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_18;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_19;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_20;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_21;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_22;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_23;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_24;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_25;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_26;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_27;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_28;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_29;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_30;
  wire [0:0] u_CSAwallace_pg_rca32_and_0_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_1_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_2_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_3_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_4_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_5_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_6_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_7_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_8_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_9_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_10_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_11_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_12_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_13_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_14_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_15_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_16_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_17_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_18_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_19_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_20_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_21_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_22_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_23_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_24_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_25_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_26_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_27_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_28_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_29_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_30_31;
  wire [0:0] u_CSAwallace_pg_rca32_and_31_31;
  wire [33:0] u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0;
  wire [33:0] u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1;
  wire [33:0] u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2;
  wire [69:0] u_CSAwallace_pg_rca32_csa0_csa_component_out;
  wire [36:0] u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3;
  wire [36:0] u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4;
  wire [36:0] u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5;
  wire [75:0] u_CSAwallace_pg_rca32_csa1_csa_component_out;
  wire [39:0] u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6;
  wire [39:0] u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7;
  wire [39:0] u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8;
  wire [81:0] u_CSAwallace_pg_rca32_csa2_csa_component_out;
  wire [42:0] u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9;
  wire [42:0] u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10;
  wire [42:0] u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11;
  wire [87:0] u_CSAwallace_pg_rca32_csa3_csa_component_out;
  wire [45:0] u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12;
  wire [45:0] u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13;
  wire [45:0] u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14;
  wire [93:0] u_CSAwallace_pg_rca32_csa4_csa_component_out;
  wire [48:0] u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15;
  wire [48:0] u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16;
  wire [48:0] u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17;
  wire [99:0] u_CSAwallace_pg_rca32_csa5_csa_component_out;
  wire [51:0] u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18;
  wire [51:0] u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19;
  wire [51:0] u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20;
  wire [105:0] u_CSAwallace_pg_rca32_csa6_csa_component_out;
  wire [54:0] u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21;
  wire [54:0] u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22;
  wire [54:0] u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23;
  wire [111:0] u_CSAwallace_pg_rca32_csa7_csa_component_out;
  wire [57:0] u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24;
  wire [57:0] u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25;
  wire [57:0] u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26;
  wire [117:0] u_CSAwallace_pg_rca32_csa8_csa_component_out;
  wire [60:0] u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27;
  wire [60:0] u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28;
  wire [60:0] u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29;
  wire [123:0] u_CSAwallace_pg_rca32_csa9_csa_component_out;
  wire [37:0] u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1;
  wire [37:0] u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1;
  wire [37:0] u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2;
  wire [77:0] u_CSAwallace_pg_rca32_csa10_csa_component_out;
  wire [40:0] u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2;
  wire [40:0] u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3;
  wire [40:0] u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3;
  wire [83:0] u_CSAwallace_pg_rca32_csa11_csa_component_out;
  wire [46:0] u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4;
  wire [46:0] u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4;
  wire [46:0] u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5;
  wire [95:0] u_CSAwallace_pg_rca32_csa12_csa_component_out;
  wire [49:0] u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5;
  wire [49:0] u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6;
  wire [49:0] u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6;
  wire [101:0] u_CSAwallace_pg_rca32_csa13_csa_component_out;
  wire [55:0] u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7;
  wire [55:0] u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7;
  wire [55:0] u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8;
  wire [113:0] u_CSAwallace_pg_rca32_csa14_csa_component_out;
  wire [58:0] u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8;
  wire [58:0] u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9;
  wire [58:0] u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9;
  wire [119:0] u_CSAwallace_pg_rca32_csa15_csa_component_out;
  wire [61:0] u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10;
  wire [61:0] u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10;
  wire [61:0] u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30;
  wire [125:0] u_CSAwallace_pg_rca32_csa16_csa_component_out;
  wire [41:0] u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11;
  wire [41:0] u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11;
  wire [41:0] u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12;
  wire [85:0] u_CSAwallace_pg_rca32_csa17_csa_component_out;
  wire [47:0] u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12;
  wire [47:0] u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13;
  wire [47:0] u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13;
  wire [97:0] u_CSAwallace_pg_rca32_csa18_csa_component_out;
  wire [56:0] u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14;
  wire [56:0] u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14;
  wire [56:0] u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15;
  wire [115:0] u_CSAwallace_pg_rca32_csa19_csa_component_out;
  wire [59:0] u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15;
  wire [59:0] u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16;
  wire [59:0] u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16;
  wire [121:0] u_CSAwallace_pg_rca32_csa20_csa_component_out;
  wire [62:0] u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17;
  wire [62:0] u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17;
  wire [62:0] u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31;
  wire [127:0] u_CSAwallace_pg_rca32_csa21_csa_component_out;
  wire [48:0] u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18;
  wire [48:0] u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18;
  wire [48:0] u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19;
  wire [99:0] u_CSAwallace_pg_rca32_csa22_csa_component_out;
  wire [57:0] u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19;
  wire [57:0] u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20;
  wire [57:0] u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20;
  wire [117:0] u_CSAwallace_pg_rca32_csa23_csa_component_out;
  wire [63:0] u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21;
  wire [63:0] u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21;
  wire [63:0] u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22;
  wire [129:0] u_CSAwallace_pg_rca32_csa24_csa_component_out;
  wire [58:0] u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23;
  wire [58:0] u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23;
  wire [58:0] u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24;
  wire [119:0] u_CSAwallace_pg_rca32_csa25_csa_component_out;
  wire [63:0] u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24;
  wire [63:0] u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25;
  wire [63:0] u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25;
  wire [129:0] u_CSAwallace_pg_rca32_csa26_csa_component_out;
  wire [63:0] u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26;
  wire [63:0] u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26;
  wire [63:0] u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27;
  wire [129:0] u_CSAwallace_pg_rca32_csa27_csa_component_out;
  wire [63:0] u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28;
  wire [63:0] u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28;
  wire [63:0] u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27;
  wire [129:0] u_CSAwallace_pg_rca32_csa28_csa_component_out;
  wire [63:0] u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29;
  wire [63:0] u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29;
  wire [63:0] u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22;
  wire [129:0] u_CSAwallace_pg_rca32_csa29_csa_component_out;
  wire [63:0] u_CSAwallace_pg_rca32_u_pg_rca64_a;
  wire [63:0] u_CSAwallace_pg_rca32_u_pg_rca64_b;
  wire [64:0] u_CSAwallace_pg_rca32_u_pg_rca64_out;

  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_0(.a(a[0]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_0_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_0(.a(a[1]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_1_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_0(.a(a[2]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_2_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_0(.a(a[3]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_3_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_0(.a(a[4]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_4_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_0(.a(a[5]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_5_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_0(.a(a[6]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_6_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_0(.a(a[7]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_7_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_0(.a(a[8]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_8_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_0(.a(a[9]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_9_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_0(.a(a[10]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_10_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_0(.a(a[11]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_11_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_0(.a(a[12]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_12_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_0(.a(a[13]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_13_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_0(.a(a[14]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_14_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_0(.a(a[15]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_15_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_0(.a(a[16]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_16_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_0(.a(a[17]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_17_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_0(.a(a[18]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_18_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_0(.a(a[19]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_19_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_0(.a(a[20]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_20_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_0(.a(a[21]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_21_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_0(.a(a[22]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_22_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_0(.a(a[23]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_23_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_0(.a(a[24]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_24_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_0(.a(a[25]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_25_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_0(.a(a[26]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_26_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_0(.a(a[27]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_27_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_0(.a(a[28]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_28_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_0(.a(a[29]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_29_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_0(.a(a[30]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_30_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_0(.a(a[31]), .b(b[0]), .out(u_CSAwallace_pg_rca32_and_31_0));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_1(.a(a[0]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_0_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_1(.a(a[1]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_1_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_1(.a(a[2]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_2_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_1(.a(a[3]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_3_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_1(.a(a[4]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_4_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_1(.a(a[5]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_5_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_1(.a(a[6]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_6_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_1(.a(a[7]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_7_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_1(.a(a[8]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_8_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_1(.a(a[9]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_9_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_1(.a(a[10]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_10_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_1(.a(a[11]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_11_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_1(.a(a[12]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_12_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_1(.a(a[13]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_13_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_1(.a(a[14]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_14_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_1(.a(a[15]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_15_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_1(.a(a[16]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_16_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_1(.a(a[17]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_17_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_1(.a(a[18]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_18_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_1(.a(a[19]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_19_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_1(.a(a[20]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_20_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_1(.a(a[21]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_21_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_1(.a(a[22]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_22_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_1(.a(a[23]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_23_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_1(.a(a[24]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_24_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_1(.a(a[25]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_25_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_1(.a(a[26]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_26_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_1(.a(a[27]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_27_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_1(.a(a[28]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_28_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_1(.a(a[29]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_29_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_1(.a(a[30]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_30_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_1(.a(a[31]), .b(b[1]), .out(u_CSAwallace_pg_rca32_and_31_1));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_2(.a(a[0]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_0_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_2(.a(a[1]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_1_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_2(.a(a[2]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_2_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_2(.a(a[3]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_3_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_2(.a(a[4]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_4_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_2(.a(a[5]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_5_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_2(.a(a[6]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_6_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_2(.a(a[7]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_7_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_2(.a(a[8]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_8_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_2(.a(a[9]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_9_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_2(.a(a[10]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_10_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_2(.a(a[11]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_11_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_2(.a(a[12]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_12_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_2(.a(a[13]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_13_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_2(.a(a[14]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_14_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_2(.a(a[15]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_15_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_2(.a(a[16]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_16_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_2(.a(a[17]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_17_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_2(.a(a[18]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_18_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_2(.a(a[19]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_19_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_2(.a(a[20]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_20_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_2(.a(a[21]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_21_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_2(.a(a[22]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_22_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_2(.a(a[23]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_23_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_2(.a(a[24]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_24_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_2(.a(a[25]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_25_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_2(.a(a[26]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_26_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_2(.a(a[27]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_27_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_2(.a(a[28]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_28_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_2(.a(a[29]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_29_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_2(.a(a[30]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_30_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_2(.a(a[31]), .b(b[2]), .out(u_CSAwallace_pg_rca32_and_31_2));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_3(.a(a[0]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_0_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_3(.a(a[1]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_1_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_3(.a(a[2]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_2_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_3(.a(a[3]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_3_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_3(.a(a[4]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_4_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_3(.a(a[5]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_5_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_3(.a(a[6]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_6_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_3(.a(a[7]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_7_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_3(.a(a[8]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_8_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_3(.a(a[9]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_9_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_3(.a(a[10]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_10_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_3(.a(a[11]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_11_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_3(.a(a[12]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_12_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_3(.a(a[13]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_13_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_3(.a(a[14]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_14_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_3(.a(a[15]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_15_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_3(.a(a[16]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_16_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_3(.a(a[17]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_17_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_3(.a(a[18]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_18_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_3(.a(a[19]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_19_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_3(.a(a[20]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_20_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_3(.a(a[21]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_21_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_3(.a(a[22]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_22_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_3(.a(a[23]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_23_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_3(.a(a[24]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_24_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_3(.a(a[25]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_25_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_3(.a(a[26]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_26_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_3(.a(a[27]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_27_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_3(.a(a[28]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_28_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_3(.a(a[29]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_29_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_3(.a(a[30]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_30_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_3(.a(a[31]), .b(b[3]), .out(u_CSAwallace_pg_rca32_and_31_3));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_4(.a(a[0]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_0_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_4(.a(a[1]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_1_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_4(.a(a[2]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_2_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_4(.a(a[3]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_3_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_4(.a(a[4]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_4_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_4(.a(a[5]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_5_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_4(.a(a[6]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_6_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_4(.a(a[7]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_7_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_4(.a(a[8]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_8_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_4(.a(a[9]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_9_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_4(.a(a[10]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_10_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_4(.a(a[11]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_11_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_4(.a(a[12]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_12_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_4(.a(a[13]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_13_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_4(.a(a[14]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_14_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_4(.a(a[15]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_15_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_4(.a(a[16]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_16_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_4(.a(a[17]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_17_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_4(.a(a[18]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_18_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_4(.a(a[19]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_19_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_4(.a(a[20]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_20_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_4(.a(a[21]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_21_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_4(.a(a[22]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_22_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_4(.a(a[23]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_23_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_4(.a(a[24]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_24_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_4(.a(a[25]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_25_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_4(.a(a[26]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_26_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_4(.a(a[27]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_27_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_4(.a(a[28]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_28_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_4(.a(a[29]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_29_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_4(.a(a[30]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_30_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_4(.a(a[31]), .b(b[4]), .out(u_CSAwallace_pg_rca32_and_31_4));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_5(.a(a[0]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_0_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_5(.a(a[1]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_1_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_5(.a(a[2]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_2_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_5(.a(a[3]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_3_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_5(.a(a[4]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_4_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_5(.a(a[5]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_5_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_5(.a(a[6]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_6_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_5(.a(a[7]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_7_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_5(.a(a[8]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_8_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_5(.a(a[9]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_9_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_5(.a(a[10]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_10_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_5(.a(a[11]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_11_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_5(.a(a[12]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_12_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_5(.a(a[13]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_13_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_5(.a(a[14]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_14_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_5(.a(a[15]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_15_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_5(.a(a[16]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_16_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_5(.a(a[17]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_17_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_5(.a(a[18]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_18_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_5(.a(a[19]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_19_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_5(.a(a[20]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_20_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_5(.a(a[21]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_21_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_5(.a(a[22]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_22_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_5(.a(a[23]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_23_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_5(.a(a[24]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_24_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_5(.a(a[25]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_25_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_5(.a(a[26]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_26_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_5(.a(a[27]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_27_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_5(.a(a[28]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_28_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_5(.a(a[29]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_29_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_5(.a(a[30]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_30_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_5(.a(a[31]), .b(b[5]), .out(u_CSAwallace_pg_rca32_and_31_5));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_6(.a(a[0]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_0_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_6(.a(a[1]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_1_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_6(.a(a[2]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_2_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_6(.a(a[3]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_3_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_6(.a(a[4]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_4_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_6(.a(a[5]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_5_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_6(.a(a[6]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_6_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_6(.a(a[7]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_7_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_6(.a(a[8]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_8_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_6(.a(a[9]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_9_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_6(.a(a[10]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_10_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_6(.a(a[11]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_11_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_6(.a(a[12]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_12_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_6(.a(a[13]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_13_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_6(.a(a[14]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_14_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_6(.a(a[15]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_15_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_6(.a(a[16]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_16_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_6(.a(a[17]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_17_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_6(.a(a[18]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_18_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_6(.a(a[19]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_19_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_6(.a(a[20]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_20_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_6(.a(a[21]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_21_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_6(.a(a[22]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_22_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_6(.a(a[23]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_23_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_6(.a(a[24]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_24_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_6(.a(a[25]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_25_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_6(.a(a[26]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_26_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_6(.a(a[27]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_27_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_6(.a(a[28]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_28_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_6(.a(a[29]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_29_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_6(.a(a[30]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_30_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_6(.a(a[31]), .b(b[6]), .out(u_CSAwallace_pg_rca32_and_31_6));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_7(.a(a[0]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_0_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_7(.a(a[1]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_1_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_7(.a(a[2]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_2_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_7(.a(a[3]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_3_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_7(.a(a[4]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_4_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_7(.a(a[5]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_5_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_7(.a(a[6]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_6_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_7(.a(a[7]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_7_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_7(.a(a[8]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_8_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_7(.a(a[9]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_9_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_7(.a(a[10]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_10_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_7(.a(a[11]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_11_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_7(.a(a[12]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_12_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_7(.a(a[13]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_13_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_7(.a(a[14]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_14_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_7(.a(a[15]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_15_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_7(.a(a[16]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_16_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_7(.a(a[17]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_17_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_7(.a(a[18]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_18_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_7(.a(a[19]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_19_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_7(.a(a[20]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_20_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_7(.a(a[21]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_21_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_7(.a(a[22]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_22_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_7(.a(a[23]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_23_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_7(.a(a[24]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_24_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_7(.a(a[25]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_25_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_7(.a(a[26]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_26_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_7(.a(a[27]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_27_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_7(.a(a[28]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_28_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_7(.a(a[29]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_29_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_7(.a(a[30]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_30_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_7(.a(a[31]), .b(b[7]), .out(u_CSAwallace_pg_rca32_and_31_7));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_8(.a(a[0]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_0_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_8(.a(a[1]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_1_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_8(.a(a[2]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_2_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_8(.a(a[3]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_3_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_8(.a(a[4]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_4_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_8(.a(a[5]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_5_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_8(.a(a[6]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_6_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_8(.a(a[7]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_7_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_8(.a(a[8]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_8_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_8(.a(a[9]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_9_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_8(.a(a[10]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_10_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_8(.a(a[11]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_11_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_8(.a(a[12]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_12_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_8(.a(a[13]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_13_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_8(.a(a[14]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_14_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_8(.a(a[15]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_15_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_8(.a(a[16]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_16_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_8(.a(a[17]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_17_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_8(.a(a[18]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_18_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_8(.a(a[19]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_19_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_8(.a(a[20]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_20_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_8(.a(a[21]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_21_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_8(.a(a[22]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_22_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_8(.a(a[23]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_23_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_8(.a(a[24]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_24_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_8(.a(a[25]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_25_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_8(.a(a[26]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_26_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_8(.a(a[27]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_27_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_8(.a(a[28]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_28_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_8(.a(a[29]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_29_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_8(.a(a[30]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_30_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_8(.a(a[31]), .b(b[8]), .out(u_CSAwallace_pg_rca32_and_31_8));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_9(.a(a[0]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_0_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_9(.a(a[1]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_1_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_9(.a(a[2]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_2_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_9(.a(a[3]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_3_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_9(.a(a[4]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_4_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_9(.a(a[5]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_5_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_9(.a(a[6]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_6_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_9(.a(a[7]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_7_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_9(.a(a[8]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_8_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_9(.a(a[9]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_9_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_9(.a(a[10]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_10_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_9(.a(a[11]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_11_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_9(.a(a[12]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_12_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_9(.a(a[13]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_13_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_9(.a(a[14]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_14_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_9(.a(a[15]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_15_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_9(.a(a[16]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_16_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_9(.a(a[17]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_17_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_9(.a(a[18]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_18_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_9(.a(a[19]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_19_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_9(.a(a[20]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_20_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_9(.a(a[21]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_21_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_9(.a(a[22]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_22_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_9(.a(a[23]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_23_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_9(.a(a[24]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_24_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_9(.a(a[25]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_25_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_9(.a(a[26]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_26_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_9(.a(a[27]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_27_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_9(.a(a[28]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_28_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_9(.a(a[29]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_29_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_9(.a(a[30]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_30_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_9(.a(a[31]), .b(b[9]), .out(u_CSAwallace_pg_rca32_and_31_9));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_10(.a(a[0]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_0_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_10(.a(a[1]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_1_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_10(.a(a[2]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_2_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_10(.a(a[3]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_3_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_10(.a(a[4]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_4_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_10(.a(a[5]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_5_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_10(.a(a[6]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_6_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_10(.a(a[7]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_7_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_10(.a(a[8]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_8_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_10(.a(a[9]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_9_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_10(.a(a[10]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_10_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_10(.a(a[11]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_11_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_10(.a(a[12]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_12_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_10(.a(a[13]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_13_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_10(.a(a[14]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_14_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_10(.a(a[15]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_15_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_10(.a(a[16]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_16_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_10(.a(a[17]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_17_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_10(.a(a[18]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_18_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_10(.a(a[19]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_19_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_10(.a(a[20]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_20_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_10(.a(a[21]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_21_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_10(.a(a[22]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_22_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_10(.a(a[23]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_23_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_10(.a(a[24]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_24_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_10(.a(a[25]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_25_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_10(.a(a[26]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_26_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_10(.a(a[27]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_27_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_10(.a(a[28]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_28_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_10(.a(a[29]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_29_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_10(.a(a[30]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_30_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_10(.a(a[31]), .b(b[10]), .out(u_CSAwallace_pg_rca32_and_31_10));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_11(.a(a[0]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_0_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_11(.a(a[1]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_1_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_11(.a(a[2]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_2_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_11(.a(a[3]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_3_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_11(.a(a[4]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_4_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_11(.a(a[5]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_5_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_11(.a(a[6]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_6_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_11(.a(a[7]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_7_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_11(.a(a[8]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_8_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_11(.a(a[9]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_9_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_11(.a(a[10]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_10_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_11(.a(a[11]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_11_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_11(.a(a[12]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_12_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_11(.a(a[13]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_13_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_11(.a(a[14]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_14_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_11(.a(a[15]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_15_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_11(.a(a[16]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_16_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_11(.a(a[17]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_17_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_11(.a(a[18]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_18_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_11(.a(a[19]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_19_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_11(.a(a[20]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_20_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_11(.a(a[21]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_21_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_11(.a(a[22]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_22_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_11(.a(a[23]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_23_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_11(.a(a[24]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_24_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_11(.a(a[25]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_25_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_11(.a(a[26]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_26_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_11(.a(a[27]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_27_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_11(.a(a[28]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_28_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_11(.a(a[29]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_29_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_11(.a(a[30]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_30_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_11(.a(a[31]), .b(b[11]), .out(u_CSAwallace_pg_rca32_and_31_11));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_12(.a(a[0]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_0_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_12(.a(a[1]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_1_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_12(.a(a[2]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_2_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_12(.a(a[3]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_3_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_12(.a(a[4]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_4_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_12(.a(a[5]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_5_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_12(.a(a[6]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_6_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_12(.a(a[7]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_7_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_12(.a(a[8]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_8_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_12(.a(a[9]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_9_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_12(.a(a[10]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_10_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_12(.a(a[11]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_11_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_12(.a(a[12]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_12_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_12(.a(a[13]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_13_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_12(.a(a[14]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_14_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_12(.a(a[15]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_15_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_12(.a(a[16]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_16_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_12(.a(a[17]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_17_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_12(.a(a[18]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_18_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_12(.a(a[19]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_19_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_12(.a(a[20]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_20_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_12(.a(a[21]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_21_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_12(.a(a[22]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_22_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_12(.a(a[23]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_23_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_12(.a(a[24]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_24_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_12(.a(a[25]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_25_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_12(.a(a[26]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_26_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_12(.a(a[27]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_27_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_12(.a(a[28]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_28_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_12(.a(a[29]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_29_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_12(.a(a[30]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_30_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_12(.a(a[31]), .b(b[12]), .out(u_CSAwallace_pg_rca32_and_31_12));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_13(.a(a[0]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_0_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_13(.a(a[1]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_1_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_13(.a(a[2]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_2_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_13(.a(a[3]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_3_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_13(.a(a[4]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_4_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_13(.a(a[5]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_5_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_13(.a(a[6]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_6_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_13(.a(a[7]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_7_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_13(.a(a[8]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_8_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_13(.a(a[9]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_9_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_13(.a(a[10]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_10_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_13(.a(a[11]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_11_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_13(.a(a[12]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_12_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_13(.a(a[13]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_13_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_13(.a(a[14]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_14_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_13(.a(a[15]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_15_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_13(.a(a[16]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_16_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_13(.a(a[17]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_17_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_13(.a(a[18]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_18_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_13(.a(a[19]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_19_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_13(.a(a[20]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_20_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_13(.a(a[21]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_21_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_13(.a(a[22]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_22_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_13(.a(a[23]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_23_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_13(.a(a[24]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_24_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_13(.a(a[25]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_25_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_13(.a(a[26]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_26_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_13(.a(a[27]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_27_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_13(.a(a[28]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_28_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_13(.a(a[29]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_29_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_13(.a(a[30]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_30_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_13(.a(a[31]), .b(b[13]), .out(u_CSAwallace_pg_rca32_and_31_13));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_14(.a(a[0]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_0_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_14(.a(a[1]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_1_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_14(.a(a[2]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_2_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_14(.a(a[3]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_3_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_14(.a(a[4]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_4_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_14(.a(a[5]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_5_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_14(.a(a[6]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_6_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_14(.a(a[7]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_7_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_14(.a(a[8]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_8_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_14(.a(a[9]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_9_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_14(.a(a[10]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_10_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_14(.a(a[11]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_11_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_14(.a(a[12]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_12_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_14(.a(a[13]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_13_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_14(.a(a[14]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_14_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_14(.a(a[15]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_15_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_14(.a(a[16]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_16_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_14(.a(a[17]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_17_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_14(.a(a[18]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_18_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_14(.a(a[19]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_19_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_14(.a(a[20]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_20_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_14(.a(a[21]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_21_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_14(.a(a[22]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_22_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_14(.a(a[23]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_23_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_14(.a(a[24]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_24_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_14(.a(a[25]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_25_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_14(.a(a[26]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_26_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_14(.a(a[27]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_27_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_14(.a(a[28]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_28_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_14(.a(a[29]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_29_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_14(.a(a[30]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_30_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_14(.a(a[31]), .b(b[14]), .out(u_CSAwallace_pg_rca32_and_31_14));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_15(.a(a[0]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_0_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_15(.a(a[1]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_1_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_15(.a(a[2]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_2_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_15(.a(a[3]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_3_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_15(.a(a[4]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_4_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_15(.a(a[5]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_5_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_15(.a(a[6]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_6_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_15(.a(a[7]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_7_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_15(.a(a[8]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_8_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_15(.a(a[9]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_9_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_15(.a(a[10]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_10_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_15(.a(a[11]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_11_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_15(.a(a[12]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_12_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_15(.a(a[13]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_13_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_15(.a(a[14]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_14_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_15(.a(a[15]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_15_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_15(.a(a[16]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_16_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_15(.a(a[17]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_17_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_15(.a(a[18]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_18_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_15(.a(a[19]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_19_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_15(.a(a[20]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_20_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_15(.a(a[21]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_21_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_15(.a(a[22]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_22_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_15(.a(a[23]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_23_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_15(.a(a[24]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_24_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_15(.a(a[25]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_25_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_15(.a(a[26]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_26_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_15(.a(a[27]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_27_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_15(.a(a[28]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_28_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_15(.a(a[29]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_29_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_15(.a(a[30]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_30_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_15(.a(a[31]), .b(b[15]), .out(u_CSAwallace_pg_rca32_and_31_15));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_16(.a(a[0]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_0_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_16(.a(a[1]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_1_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_16(.a(a[2]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_2_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_16(.a(a[3]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_3_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_16(.a(a[4]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_4_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_16(.a(a[5]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_5_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_16(.a(a[6]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_6_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_16(.a(a[7]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_7_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_16(.a(a[8]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_8_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_16(.a(a[9]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_9_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_16(.a(a[10]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_10_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_16(.a(a[11]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_11_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_16(.a(a[12]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_12_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_16(.a(a[13]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_13_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_16(.a(a[14]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_14_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_16(.a(a[15]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_15_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_16(.a(a[16]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_16_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_16(.a(a[17]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_17_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_16(.a(a[18]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_18_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_16(.a(a[19]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_19_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_16(.a(a[20]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_20_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_16(.a(a[21]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_21_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_16(.a(a[22]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_22_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_16(.a(a[23]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_23_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_16(.a(a[24]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_24_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_16(.a(a[25]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_25_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_16(.a(a[26]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_26_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_16(.a(a[27]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_27_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_16(.a(a[28]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_28_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_16(.a(a[29]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_29_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_16(.a(a[30]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_30_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_16(.a(a[31]), .b(b[16]), .out(u_CSAwallace_pg_rca32_and_31_16));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_17(.a(a[0]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_0_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_17(.a(a[1]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_1_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_17(.a(a[2]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_2_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_17(.a(a[3]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_3_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_17(.a(a[4]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_4_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_17(.a(a[5]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_5_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_17(.a(a[6]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_6_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_17(.a(a[7]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_7_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_17(.a(a[8]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_8_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_17(.a(a[9]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_9_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_17(.a(a[10]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_10_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_17(.a(a[11]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_11_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_17(.a(a[12]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_12_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_17(.a(a[13]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_13_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_17(.a(a[14]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_14_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_17(.a(a[15]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_15_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_17(.a(a[16]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_16_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_17(.a(a[17]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_17_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_17(.a(a[18]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_18_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_17(.a(a[19]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_19_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_17(.a(a[20]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_20_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_17(.a(a[21]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_21_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_17(.a(a[22]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_22_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_17(.a(a[23]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_23_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_17(.a(a[24]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_24_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_17(.a(a[25]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_25_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_17(.a(a[26]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_26_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_17(.a(a[27]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_27_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_17(.a(a[28]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_28_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_17(.a(a[29]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_29_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_17(.a(a[30]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_30_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_17(.a(a[31]), .b(b[17]), .out(u_CSAwallace_pg_rca32_and_31_17));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_18(.a(a[0]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_0_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_18(.a(a[1]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_1_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_18(.a(a[2]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_2_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_18(.a(a[3]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_3_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_18(.a(a[4]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_4_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_18(.a(a[5]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_5_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_18(.a(a[6]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_6_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_18(.a(a[7]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_7_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_18(.a(a[8]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_8_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_18(.a(a[9]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_9_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_18(.a(a[10]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_10_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_18(.a(a[11]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_11_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_18(.a(a[12]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_12_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_18(.a(a[13]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_13_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_18(.a(a[14]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_14_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_18(.a(a[15]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_15_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_18(.a(a[16]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_16_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_18(.a(a[17]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_17_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_18(.a(a[18]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_18_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_18(.a(a[19]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_19_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_18(.a(a[20]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_20_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_18(.a(a[21]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_21_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_18(.a(a[22]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_22_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_18(.a(a[23]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_23_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_18(.a(a[24]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_24_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_18(.a(a[25]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_25_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_18(.a(a[26]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_26_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_18(.a(a[27]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_27_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_18(.a(a[28]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_28_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_18(.a(a[29]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_29_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_18(.a(a[30]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_30_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_18(.a(a[31]), .b(b[18]), .out(u_CSAwallace_pg_rca32_and_31_18));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_19(.a(a[0]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_0_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_19(.a(a[1]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_1_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_19(.a(a[2]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_2_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_19(.a(a[3]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_3_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_19(.a(a[4]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_4_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_19(.a(a[5]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_5_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_19(.a(a[6]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_6_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_19(.a(a[7]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_7_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_19(.a(a[8]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_8_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_19(.a(a[9]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_9_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_19(.a(a[10]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_10_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_19(.a(a[11]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_11_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_19(.a(a[12]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_12_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_19(.a(a[13]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_13_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_19(.a(a[14]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_14_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_19(.a(a[15]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_15_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_19(.a(a[16]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_16_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_19(.a(a[17]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_17_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_19(.a(a[18]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_18_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_19(.a(a[19]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_19_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_19(.a(a[20]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_20_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_19(.a(a[21]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_21_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_19(.a(a[22]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_22_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_19(.a(a[23]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_23_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_19(.a(a[24]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_24_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_19(.a(a[25]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_25_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_19(.a(a[26]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_26_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_19(.a(a[27]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_27_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_19(.a(a[28]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_28_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_19(.a(a[29]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_29_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_19(.a(a[30]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_30_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_19(.a(a[31]), .b(b[19]), .out(u_CSAwallace_pg_rca32_and_31_19));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_20(.a(a[0]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_0_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_20(.a(a[1]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_1_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_20(.a(a[2]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_2_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_20(.a(a[3]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_3_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_20(.a(a[4]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_4_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_20(.a(a[5]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_5_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_20(.a(a[6]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_6_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_20(.a(a[7]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_7_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_20(.a(a[8]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_8_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_20(.a(a[9]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_9_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_20(.a(a[10]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_10_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_20(.a(a[11]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_11_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_20(.a(a[12]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_12_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_20(.a(a[13]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_13_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_20(.a(a[14]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_14_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_20(.a(a[15]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_15_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_20(.a(a[16]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_16_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_20(.a(a[17]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_17_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_20(.a(a[18]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_18_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_20(.a(a[19]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_19_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_20(.a(a[20]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_20_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_20(.a(a[21]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_21_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_20(.a(a[22]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_22_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_20(.a(a[23]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_23_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_20(.a(a[24]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_24_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_20(.a(a[25]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_25_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_20(.a(a[26]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_26_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_20(.a(a[27]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_27_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_20(.a(a[28]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_28_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_20(.a(a[29]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_29_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_20(.a(a[30]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_30_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_20(.a(a[31]), .b(b[20]), .out(u_CSAwallace_pg_rca32_and_31_20));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_21(.a(a[0]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_0_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_21(.a(a[1]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_1_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_21(.a(a[2]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_2_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_21(.a(a[3]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_3_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_21(.a(a[4]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_4_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_21(.a(a[5]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_5_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_21(.a(a[6]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_6_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_21(.a(a[7]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_7_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_21(.a(a[8]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_8_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_21(.a(a[9]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_9_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_21(.a(a[10]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_10_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_21(.a(a[11]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_11_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_21(.a(a[12]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_12_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_21(.a(a[13]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_13_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_21(.a(a[14]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_14_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_21(.a(a[15]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_15_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_21(.a(a[16]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_16_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_21(.a(a[17]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_17_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_21(.a(a[18]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_18_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_21(.a(a[19]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_19_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_21(.a(a[20]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_20_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_21(.a(a[21]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_21_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_21(.a(a[22]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_22_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_21(.a(a[23]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_23_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_21(.a(a[24]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_24_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_21(.a(a[25]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_25_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_21(.a(a[26]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_26_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_21(.a(a[27]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_27_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_21(.a(a[28]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_28_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_21(.a(a[29]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_29_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_21(.a(a[30]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_30_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_21(.a(a[31]), .b(b[21]), .out(u_CSAwallace_pg_rca32_and_31_21));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_22(.a(a[0]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_0_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_22(.a(a[1]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_1_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_22(.a(a[2]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_2_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_22(.a(a[3]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_3_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_22(.a(a[4]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_4_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_22(.a(a[5]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_5_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_22(.a(a[6]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_6_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_22(.a(a[7]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_7_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_22(.a(a[8]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_8_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_22(.a(a[9]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_9_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_22(.a(a[10]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_10_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_22(.a(a[11]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_11_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_22(.a(a[12]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_12_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_22(.a(a[13]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_13_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_22(.a(a[14]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_14_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_22(.a(a[15]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_15_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_22(.a(a[16]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_16_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_22(.a(a[17]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_17_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_22(.a(a[18]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_18_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_22(.a(a[19]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_19_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_22(.a(a[20]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_20_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_22(.a(a[21]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_21_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_22(.a(a[22]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_22_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_22(.a(a[23]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_23_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_22(.a(a[24]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_24_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_22(.a(a[25]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_25_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_22(.a(a[26]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_26_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_22(.a(a[27]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_27_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_22(.a(a[28]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_28_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_22(.a(a[29]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_29_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_22(.a(a[30]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_30_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_22(.a(a[31]), .b(b[22]), .out(u_CSAwallace_pg_rca32_and_31_22));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_23(.a(a[0]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_0_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_23(.a(a[1]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_1_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_23(.a(a[2]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_2_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_23(.a(a[3]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_3_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_23(.a(a[4]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_4_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_23(.a(a[5]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_5_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_23(.a(a[6]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_6_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_23(.a(a[7]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_7_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_23(.a(a[8]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_8_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_23(.a(a[9]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_9_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_23(.a(a[10]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_10_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_23(.a(a[11]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_11_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_23(.a(a[12]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_12_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_23(.a(a[13]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_13_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_23(.a(a[14]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_14_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_23(.a(a[15]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_15_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_23(.a(a[16]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_16_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_23(.a(a[17]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_17_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_23(.a(a[18]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_18_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_23(.a(a[19]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_19_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_23(.a(a[20]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_20_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_23(.a(a[21]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_21_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_23(.a(a[22]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_22_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_23(.a(a[23]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_23_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_23(.a(a[24]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_24_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_23(.a(a[25]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_25_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_23(.a(a[26]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_26_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_23(.a(a[27]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_27_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_23(.a(a[28]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_28_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_23(.a(a[29]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_29_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_23(.a(a[30]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_30_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_23(.a(a[31]), .b(b[23]), .out(u_CSAwallace_pg_rca32_and_31_23));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_24(.a(a[0]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_0_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_24(.a(a[1]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_1_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_24(.a(a[2]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_2_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_24(.a(a[3]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_3_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_24(.a(a[4]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_4_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_24(.a(a[5]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_5_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_24(.a(a[6]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_6_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_24(.a(a[7]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_7_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_24(.a(a[8]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_8_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_24(.a(a[9]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_9_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_24(.a(a[10]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_10_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_24(.a(a[11]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_11_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_24(.a(a[12]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_12_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_24(.a(a[13]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_13_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_24(.a(a[14]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_14_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_24(.a(a[15]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_15_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_24(.a(a[16]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_16_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_24(.a(a[17]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_17_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_24(.a(a[18]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_18_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_24(.a(a[19]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_19_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_24(.a(a[20]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_20_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_24(.a(a[21]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_21_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_24(.a(a[22]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_22_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_24(.a(a[23]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_23_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_24(.a(a[24]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_24_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_24(.a(a[25]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_25_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_24(.a(a[26]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_26_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_24(.a(a[27]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_27_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_24(.a(a[28]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_28_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_24(.a(a[29]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_29_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_24(.a(a[30]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_30_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_24(.a(a[31]), .b(b[24]), .out(u_CSAwallace_pg_rca32_and_31_24));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_25(.a(a[0]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_0_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_25(.a(a[1]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_1_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_25(.a(a[2]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_2_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_25(.a(a[3]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_3_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_25(.a(a[4]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_4_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_25(.a(a[5]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_5_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_25(.a(a[6]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_6_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_25(.a(a[7]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_7_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_25(.a(a[8]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_8_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_25(.a(a[9]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_9_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_25(.a(a[10]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_10_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_25(.a(a[11]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_11_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_25(.a(a[12]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_12_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_25(.a(a[13]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_13_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_25(.a(a[14]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_14_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_25(.a(a[15]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_15_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_25(.a(a[16]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_16_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_25(.a(a[17]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_17_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_25(.a(a[18]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_18_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_25(.a(a[19]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_19_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_25(.a(a[20]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_20_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_25(.a(a[21]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_21_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_25(.a(a[22]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_22_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_25(.a(a[23]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_23_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_25(.a(a[24]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_24_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_25(.a(a[25]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_25_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_25(.a(a[26]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_26_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_25(.a(a[27]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_27_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_25(.a(a[28]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_28_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_25(.a(a[29]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_29_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_25(.a(a[30]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_30_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_25(.a(a[31]), .b(b[25]), .out(u_CSAwallace_pg_rca32_and_31_25));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_26(.a(a[0]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_0_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_26(.a(a[1]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_1_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_26(.a(a[2]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_2_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_26(.a(a[3]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_3_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_26(.a(a[4]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_4_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_26(.a(a[5]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_5_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_26(.a(a[6]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_6_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_26(.a(a[7]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_7_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_26(.a(a[8]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_8_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_26(.a(a[9]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_9_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_26(.a(a[10]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_10_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_26(.a(a[11]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_11_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_26(.a(a[12]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_12_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_26(.a(a[13]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_13_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_26(.a(a[14]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_14_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_26(.a(a[15]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_15_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_26(.a(a[16]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_16_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_26(.a(a[17]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_17_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_26(.a(a[18]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_18_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_26(.a(a[19]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_19_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_26(.a(a[20]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_20_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_26(.a(a[21]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_21_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_26(.a(a[22]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_22_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_26(.a(a[23]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_23_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_26(.a(a[24]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_24_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_26(.a(a[25]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_25_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_26(.a(a[26]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_26_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_26(.a(a[27]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_27_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_26(.a(a[28]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_28_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_26(.a(a[29]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_29_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_26(.a(a[30]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_30_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_26(.a(a[31]), .b(b[26]), .out(u_CSAwallace_pg_rca32_and_31_26));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_27(.a(a[0]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_0_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_27(.a(a[1]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_1_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_27(.a(a[2]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_2_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_27(.a(a[3]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_3_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_27(.a(a[4]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_4_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_27(.a(a[5]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_5_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_27(.a(a[6]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_6_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_27(.a(a[7]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_7_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_27(.a(a[8]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_8_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_27(.a(a[9]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_9_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_27(.a(a[10]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_10_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_27(.a(a[11]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_11_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_27(.a(a[12]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_12_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_27(.a(a[13]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_13_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_27(.a(a[14]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_14_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_27(.a(a[15]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_15_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_27(.a(a[16]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_16_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_27(.a(a[17]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_17_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_27(.a(a[18]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_18_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_27(.a(a[19]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_19_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_27(.a(a[20]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_20_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_27(.a(a[21]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_21_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_27(.a(a[22]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_22_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_27(.a(a[23]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_23_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_27(.a(a[24]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_24_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_27(.a(a[25]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_25_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_27(.a(a[26]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_26_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_27(.a(a[27]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_27_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_27(.a(a[28]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_28_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_27(.a(a[29]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_29_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_27(.a(a[30]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_30_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_27(.a(a[31]), .b(b[27]), .out(u_CSAwallace_pg_rca32_and_31_27));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_28(.a(a[0]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_0_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_28(.a(a[1]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_1_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_28(.a(a[2]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_2_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_28(.a(a[3]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_3_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_28(.a(a[4]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_4_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_28(.a(a[5]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_5_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_28(.a(a[6]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_6_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_28(.a(a[7]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_7_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_28(.a(a[8]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_8_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_28(.a(a[9]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_9_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_28(.a(a[10]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_10_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_28(.a(a[11]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_11_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_28(.a(a[12]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_12_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_28(.a(a[13]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_13_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_28(.a(a[14]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_14_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_28(.a(a[15]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_15_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_28(.a(a[16]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_16_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_28(.a(a[17]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_17_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_28(.a(a[18]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_18_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_28(.a(a[19]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_19_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_28(.a(a[20]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_20_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_28(.a(a[21]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_21_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_28(.a(a[22]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_22_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_28(.a(a[23]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_23_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_28(.a(a[24]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_24_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_28(.a(a[25]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_25_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_28(.a(a[26]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_26_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_28(.a(a[27]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_27_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_28(.a(a[28]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_28_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_28(.a(a[29]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_29_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_28(.a(a[30]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_30_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_28(.a(a[31]), .b(b[28]), .out(u_CSAwallace_pg_rca32_and_31_28));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_29(.a(a[0]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_0_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_29(.a(a[1]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_1_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_29(.a(a[2]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_2_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_29(.a(a[3]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_3_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_29(.a(a[4]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_4_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_29(.a(a[5]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_5_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_29(.a(a[6]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_6_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_29(.a(a[7]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_7_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_29(.a(a[8]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_8_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_29(.a(a[9]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_9_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_29(.a(a[10]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_10_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_29(.a(a[11]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_11_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_29(.a(a[12]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_12_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_29(.a(a[13]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_13_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_29(.a(a[14]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_14_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_29(.a(a[15]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_15_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_29(.a(a[16]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_16_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_29(.a(a[17]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_17_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_29(.a(a[18]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_18_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_29(.a(a[19]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_19_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_29(.a(a[20]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_20_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_29(.a(a[21]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_21_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_29(.a(a[22]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_22_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_29(.a(a[23]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_23_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_29(.a(a[24]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_24_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_29(.a(a[25]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_25_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_29(.a(a[26]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_26_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_29(.a(a[27]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_27_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_29(.a(a[28]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_28_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_29(.a(a[29]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_29_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_29(.a(a[30]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_30_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_29(.a(a[31]), .b(b[29]), .out(u_CSAwallace_pg_rca32_and_31_29));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_30(.a(a[0]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_0_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_30(.a(a[1]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_1_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_30(.a(a[2]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_2_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_30(.a(a[3]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_3_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_30(.a(a[4]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_4_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_30(.a(a[5]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_5_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_30(.a(a[6]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_6_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_30(.a(a[7]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_7_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_30(.a(a[8]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_8_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_30(.a(a[9]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_9_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_30(.a(a[10]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_10_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_30(.a(a[11]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_11_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_30(.a(a[12]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_12_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_30(.a(a[13]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_13_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_30(.a(a[14]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_14_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_30(.a(a[15]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_15_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_30(.a(a[16]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_16_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_30(.a(a[17]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_17_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_30(.a(a[18]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_18_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_30(.a(a[19]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_19_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_30(.a(a[20]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_20_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_30(.a(a[21]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_21_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_30(.a(a[22]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_22_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_30(.a(a[23]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_23_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_30(.a(a[24]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_24_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_30(.a(a[25]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_25_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_30(.a(a[26]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_26_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_30(.a(a[27]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_27_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_30(.a(a[28]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_28_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_30(.a(a[29]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_29_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_30(.a(a[30]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_30_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_30(.a(a[31]), .b(b[30]), .out(u_CSAwallace_pg_rca32_and_31_30));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_0_31(.a(a[0]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_0_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_1_31(.a(a[1]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_1_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_2_31(.a(a[2]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_2_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_3_31(.a(a[3]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_3_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_4_31(.a(a[4]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_4_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_5_31(.a(a[5]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_5_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_6_31(.a(a[6]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_6_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_7_31(.a(a[7]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_7_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_8_31(.a(a[8]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_8_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_9_31(.a(a[9]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_9_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_10_31(.a(a[10]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_10_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_11_31(.a(a[11]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_11_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_12_31(.a(a[12]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_12_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_13_31(.a(a[13]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_13_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_14_31(.a(a[14]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_14_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_15_31(.a(a[15]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_15_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_16_31(.a(a[16]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_16_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_17_31(.a(a[17]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_17_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_18_31(.a(a[18]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_18_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_19_31(.a(a[19]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_19_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_20_31(.a(a[20]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_20_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_21_31(.a(a[21]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_21_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_22_31(.a(a[22]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_22_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_23_31(.a(a[23]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_23_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_24_31(.a(a[24]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_24_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_25_31(.a(a[25]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_25_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_26_31(.a(a[26]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_26_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_27_31(.a(a[27]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_27_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_28_31(.a(a[28]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_28_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_29_31(.a(a[29]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_29_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_30_31(.a(a[30]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_30_31));
  and_gate and_gate_u_CSAwallace_pg_rca32_and_31_31(.a(a[31]), .b(b[31]), .out(u_CSAwallace_pg_rca32_and_31_31));
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[0] = u_CSAwallace_pg_rca32_and_0_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[1] = u_CSAwallace_pg_rca32_and_1_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[2] = u_CSAwallace_pg_rca32_and_2_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[3] = u_CSAwallace_pg_rca32_and_3_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[4] = u_CSAwallace_pg_rca32_and_4_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[5] = u_CSAwallace_pg_rca32_and_5_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[6] = u_CSAwallace_pg_rca32_and_6_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[7] = u_CSAwallace_pg_rca32_and_7_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[8] = u_CSAwallace_pg_rca32_and_8_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[9] = u_CSAwallace_pg_rca32_and_9_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[10] = u_CSAwallace_pg_rca32_and_10_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[11] = u_CSAwallace_pg_rca32_and_11_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[12] = u_CSAwallace_pg_rca32_and_12_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[13] = u_CSAwallace_pg_rca32_and_13_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[14] = u_CSAwallace_pg_rca32_and_14_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[15] = u_CSAwallace_pg_rca32_and_15_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[16] = u_CSAwallace_pg_rca32_and_16_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[17] = u_CSAwallace_pg_rca32_and_17_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[18] = u_CSAwallace_pg_rca32_and_18_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[19] = u_CSAwallace_pg_rca32_and_19_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[20] = u_CSAwallace_pg_rca32_and_20_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[21] = u_CSAwallace_pg_rca32_and_21_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[22] = u_CSAwallace_pg_rca32_and_22_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[23] = u_CSAwallace_pg_rca32_and_23_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[24] = u_CSAwallace_pg_rca32_and_24_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[25] = u_CSAwallace_pg_rca32_and_25_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[26] = u_CSAwallace_pg_rca32_and_26_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[27] = u_CSAwallace_pg_rca32_and_27_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[28] = u_CSAwallace_pg_rca32_and_28_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[29] = u_CSAwallace_pg_rca32_and_29_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[30] = u_CSAwallace_pg_rca32_and_30_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[31] = u_CSAwallace_pg_rca32_and_31_0[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[32] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0[33] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[1] = u_CSAwallace_pg_rca32_and_0_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[2] = u_CSAwallace_pg_rca32_and_1_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[3] = u_CSAwallace_pg_rca32_and_2_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[4] = u_CSAwallace_pg_rca32_and_3_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[5] = u_CSAwallace_pg_rca32_and_4_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[6] = u_CSAwallace_pg_rca32_and_5_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[7] = u_CSAwallace_pg_rca32_and_6_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[8] = u_CSAwallace_pg_rca32_and_7_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[9] = u_CSAwallace_pg_rca32_and_8_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[10] = u_CSAwallace_pg_rca32_and_9_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[11] = u_CSAwallace_pg_rca32_and_10_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[12] = u_CSAwallace_pg_rca32_and_11_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[13] = u_CSAwallace_pg_rca32_and_12_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[14] = u_CSAwallace_pg_rca32_and_13_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[15] = u_CSAwallace_pg_rca32_and_14_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[16] = u_CSAwallace_pg_rca32_and_15_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[17] = u_CSAwallace_pg_rca32_and_16_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[18] = u_CSAwallace_pg_rca32_and_17_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[19] = u_CSAwallace_pg_rca32_and_18_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[20] = u_CSAwallace_pg_rca32_and_19_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[21] = u_CSAwallace_pg_rca32_and_20_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[22] = u_CSAwallace_pg_rca32_and_21_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[23] = u_CSAwallace_pg_rca32_and_22_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[24] = u_CSAwallace_pg_rca32_and_23_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[25] = u_CSAwallace_pg_rca32_and_24_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[26] = u_CSAwallace_pg_rca32_and_25_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[27] = u_CSAwallace_pg_rca32_and_26_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[28] = u_CSAwallace_pg_rca32_and_27_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[29] = u_CSAwallace_pg_rca32_and_28_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[30] = u_CSAwallace_pg_rca32_and_29_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[31] = u_CSAwallace_pg_rca32_and_30_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[32] = u_CSAwallace_pg_rca32_and_31_1[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1[33] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[2] = u_CSAwallace_pg_rca32_and_0_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[3] = u_CSAwallace_pg_rca32_and_1_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[4] = u_CSAwallace_pg_rca32_and_2_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[5] = u_CSAwallace_pg_rca32_and_3_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[6] = u_CSAwallace_pg_rca32_and_4_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[7] = u_CSAwallace_pg_rca32_and_5_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[8] = u_CSAwallace_pg_rca32_and_6_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[9] = u_CSAwallace_pg_rca32_and_7_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[10] = u_CSAwallace_pg_rca32_and_8_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[11] = u_CSAwallace_pg_rca32_and_9_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[12] = u_CSAwallace_pg_rca32_and_10_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[13] = u_CSAwallace_pg_rca32_and_11_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[14] = u_CSAwallace_pg_rca32_and_12_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[15] = u_CSAwallace_pg_rca32_and_13_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[16] = u_CSAwallace_pg_rca32_and_14_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[17] = u_CSAwallace_pg_rca32_and_15_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[18] = u_CSAwallace_pg_rca32_and_16_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[19] = u_CSAwallace_pg_rca32_and_17_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[20] = u_CSAwallace_pg_rca32_and_18_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[21] = u_CSAwallace_pg_rca32_and_19_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[22] = u_CSAwallace_pg_rca32_and_20_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[23] = u_CSAwallace_pg_rca32_and_21_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[24] = u_CSAwallace_pg_rca32_and_22_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[25] = u_CSAwallace_pg_rca32_and_23_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[26] = u_CSAwallace_pg_rca32_and_24_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[27] = u_CSAwallace_pg_rca32_and_25_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[28] = u_CSAwallace_pg_rca32_and_26_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[29] = u_CSAwallace_pg_rca32_and_27_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[30] = u_CSAwallace_pg_rca32_and_28_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[31] = u_CSAwallace_pg_rca32_and_29_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[32] = u_CSAwallace_pg_rca32_and_30_2[0];
  assign u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2[33] = u_CSAwallace_pg_rca32_and_31_2[0];
  csa_component34 csa_component34_u_CSAwallace_pg_rca32_csa0_csa_component_out(.a(u_CSAwallace_pg_rca32_csa0_csa_component_pp_row0), .b(u_CSAwallace_pg_rca32_csa0_csa_component_pp_row1), .c(u_CSAwallace_pg_rca32_csa0_csa_component_pp_row2), .csa_component34_out(u_CSAwallace_pg_rca32_csa0_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[3] = u_CSAwallace_pg_rca32_and_0_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[4] = u_CSAwallace_pg_rca32_and_1_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[5] = u_CSAwallace_pg_rca32_and_2_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[6] = u_CSAwallace_pg_rca32_and_3_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[7] = u_CSAwallace_pg_rca32_and_4_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[8] = u_CSAwallace_pg_rca32_and_5_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[9] = u_CSAwallace_pg_rca32_and_6_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[10] = u_CSAwallace_pg_rca32_and_7_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[11] = u_CSAwallace_pg_rca32_and_8_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[12] = u_CSAwallace_pg_rca32_and_9_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[13] = u_CSAwallace_pg_rca32_and_10_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[14] = u_CSAwallace_pg_rca32_and_11_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[15] = u_CSAwallace_pg_rca32_and_12_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[16] = u_CSAwallace_pg_rca32_and_13_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[17] = u_CSAwallace_pg_rca32_and_14_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[18] = u_CSAwallace_pg_rca32_and_15_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[19] = u_CSAwallace_pg_rca32_and_16_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[20] = u_CSAwallace_pg_rca32_and_17_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[21] = u_CSAwallace_pg_rca32_and_18_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[22] = u_CSAwallace_pg_rca32_and_19_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[23] = u_CSAwallace_pg_rca32_and_20_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[24] = u_CSAwallace_pg_rca32_and_21_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[25] = u_CSAwallace_pg_rca32_and_22_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[26] = u_CSAwallace_pg_rca32_and_23_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[27] = u_CSAwallace_pg_rca32_and_24_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[28] = u_CSAwallace_pg_rca32_and_25_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[29] = u_CSAwallace_pg_rca32_and_26_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[30] = u_CSAwallace_pg_rca32_and_27_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[31] = u_CSAwallace_pg_rca32_and_28_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[32] = u_CSAwallace_pg_rca32_and_29_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[33] = u_CSAwallace_pg_rca32_and_30_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[34] = u_CSAwallace_pg_rca32_and_31_3[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[35] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3[36] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[4] = u_CSAwallace_pg_rca32_and_0_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[5] = u_CSAwallace_pg_rca32_and_1_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[6] = u_CSAwallace_pg_rca32_and_2_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[7] = u_CSAwallace_pg_rca32_and_3_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[8] = u_CSAwallace_pg_rca32_and_4_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[9] = u_CSAwallace_pg_rca32_and_5_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[10] = u_CSAwallace_pg_rca32_and_6_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[11] = u_CSAwallace_pg_rca32_and_7_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[12] = u_CSAwallace_pg_rca32_and_8_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[13] = u_CSAwallace_pg_rca32_and_9_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[14] = u_CSAwallace_pg_rca32_and_10_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[15] = u_CSAwallace_pg_rca32_and_11_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[16] = u_CSAwallace_pg_rca32_and_12_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[17] = u_CSAwallace_pg_rca32_and_13_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[18] = u_CSAwallace_pg_rca32_and_14_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[19] = u_CSAwallace_pg_rca32_and_15_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[20] = u_CSAwallace_pg_rca32_and_16_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[21] = u_CSAwallace_pg_rca32_and_17_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[22] = u_CSAwallace_pg_rca32_and_18_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[23] = u_CSAwallace_pg_rca32_and_19_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[24] = u_CSAwallace_pg_rca32_and_20_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[25] = u_CSAwallace_pg_rca32_and_21_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[26] = u_CSAwallace_pg_rca32_and_22_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[27] = u_CSAwallace_pg_rca32_and_23_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[28] = u_CSAwallace_pg_rca32_and_24_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[29] = u_CSAwallace_pg_rca32_and_25_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[30] = u_CSAwallace_pg_rca32_and_26_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[31] = u_CSAwallace_pg_rca32_and_27_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[32] = u_CSAwallace_pg_rca32_and_28_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[33] = u_CSAwallace_pg_rca32_and_29_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[34] = u_CSAwallace_pg_rca32_and_30_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[35] = u_CSAwallace_pg_rca32_and_31_4[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4[36] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[5] = u_CSAwallace_pg_rca32_and_0_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[6] = u_CSAwallace_pg_rca32_and_1_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[7] = u_CSAwallace_pg_rca32_and_2_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[8] = u_CSAwallace_pg_rca32_and_3_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[9] = u_CSAwallace_pg_rca32_and_4_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[10] = u_CSAwallace_pg_rca32_and_5_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[11] = u_CSAwallace_pg_rca32_and_6_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[12] = u_CSAwallace_pg_rca32_and_7_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[13] = u_CSAwallace_pg_rca32_and_8_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[14] = u_CSAwallace_pg_rca32_and_9_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[15] = u_CSAwallace_pg_rca32_and_10_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[16] = u_CSAwallace_pg_rca32_and_11_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[17] = u_CSAwallace_pg_rca32_and_12_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[18] = u_CSAwallace_pg_rca32_and_13_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[19] = u_CSAwallace_pg_rca32_and_14_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[20] = u_CSAwallace_pg_rca32_and_15_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[21] = u_CSAwallace_pg_rca32_and_16_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[22] = u_CSAwallace_pg_rca32_and_17_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[23] = u_CSAwallace_pg_rca32_and_18_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[24] = u_CSAwallace_pg_rca32_and_19_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[25] = u_CSAwallace_pg_rca32_and_20_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[26] = u_CSAwallace_pg_rca32_and_21_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[27] = u_CSAwallace_pg_rca32_and_22_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[28] = u_CSAwallace_pg_rca32_and_23_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[29] = u_CSAwallace_pg_rca32_and_24_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[30] = u_CSAwallace_pg_rca32_and_25_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[31] = u_CSAwallace_pg_rca32_and_26_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[32] = u_CSAwallace_pg_rca32_and_27_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[33] = u_CSAwallace_pg_rca32_and_28_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[34] = u_CSAwallace_pg_rca32_and_29_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[35] = u_CSAwallace_pg_rca32_and_30_5[0];
  assign u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5[36] = u_CSAwallace_pg_rca32_and_31_5[0];
  csa_component37 csa_component37_u_CSAwallace_pg_rca32_csa1_csa_component_out(.a(u_CSAwallace_pg_rca32_csa1_csa_component_pp_row3), .b(u_CSAwallace_pg_rca32_csa1_csa_component_pp_row4), .c(u_CSAwallace_pg_rca32_csa1_csa_component_pp_row5), .csa_component37_out(u_CSAwallace_pg_rca32_csa1_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[6] = u_CSAwallace_pg_rca32_and_0_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[7] = u_CSAwallace_pg_rca32_and_1_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[8] = u_CSAwallace_pg_rca32_and_2_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[9] = u_CSAwallace_pg_rca32_and_3_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[10] = u_CSAwallace_pg_rca32_and_4_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[11] = u_CSAwallace_pg_rca32_and_5_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[12] = u_CSAwallace_pg_rca32_and_6_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[13] = u_CSAwallace_pg_rca32_and_7_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[14] = u_CSAwallace_pg_rca32_and_8_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[15] = u_CSAwallace_pg_rca32_and_9_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[16] = u_CSAwallace_pg_rca32_and_10_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[17] = u_CSAwallace_pg_rca32_and_11_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[18] = u_CSAwallace_pg_rca32_and_12_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[19] = u_CSAwallace_pg_rca32_and_13_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[20] = u_CSAwallace_pg_rca32_and_14_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[21] = u_CSAwallace_pg_rca32_and_15_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[22] = u_CSAwallace_pg_rca32_and_16_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[23] = u_CSAwallace_pg_rca32_and_17_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[24] = u_CSAwallace_pg_rca32_and_18_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[25] = u_CSAwallace_pg_rca32_and_19_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[26] = u_CSAwallace_pg_rca32_and_20_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[27] = u_CSAwallace_pg_rca32_and_21_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[28] = u_CSAwallace_pg_rca32_and_22_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[29] = u_CSAwallace_pg_rca32_and_23_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[30] = u_CSAwallace_pg_rca32_and_24_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[31] = u_CSAwallace_pg_rca32_and_25_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[32] = u_CSAwallace_pg_rca32_and_26_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[33] = u_CSAwallace_pg_rca32_and_27_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[34] = u_CSAwallace_pg_rca32_and_28_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[35] = u_CSAwallace_pg_rca32_and_29_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[36] = u_CSAwallace_pg_rca32_and_30_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[37] = u_CSAwallace_pg_rca32_and_31_6[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[38] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6[39] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[7] = u_CSAwallace_pg_rca32_and_0_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[8] = u_CSAwallace_pg_rca32_and_1_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[9] = u_CSAwallace_pg_rca32_and_2_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[10] = u_CSAwallace_pg_rca32_and_3_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[11] = u_CSAwallace_pg_rca32_and_4_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[12] = u_CSAwallace_pg_rca32_and_5_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[13] = u_CSAwallace_pg_rca32_and_6_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[14] = u_CSAwallace_pg_rca32_and_7_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[15] = u_CSAwallace_pg_rca32_and_8_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[16] = u_CSAwallace_pg_rca32_and_9_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[17] = u_CSAwallace_pg_rca32_and_10_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[18] = u_CSAwallace_pg_rca32_and_11_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[19] = u_CSAwallace_pg_rca32_and_12_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[20] = u_CSAwallace_pg_rca32_and_13_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[21] = u_CSAwallace_pg_rca32_and_14_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[22] = u_CSAwallace_pg_rca32_and_15_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[23] = u_CSAwallace_pg_rca32_and_16_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[24] = u_CSAwallace_pg_rca32_and_17_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[25] = u_CSAwallace_pg_rca32_and_18_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[26] = u_CSAwallace_pg_rca32_and_19_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[27] = u_CSAwallace_pg_rca32_and_20_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[28] = u_CSAwallace_pg_rca32_and_21_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[29] = u_CSAwallace_pg_rca32_and_22_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[30] = u_CSAwallace_pg_rca32_and_23_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[31] = u_CSAwallace_pg_rca32_and_24_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[32] = u_CSAwallace_pg_rca32_and_25_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[33] = u_CSAwallace_pg_rca32_and_26_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[34] = u_CSAwallace_pg_rca32_and_27_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[35] = u_CSAwallace_pg_rca32_and_28_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[36] = u_CSAwallace_pg_rca32_and_29_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[37] = u_CSAwallace_pg_rca32_and_30_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[38] = u_CSAwallace_pg_rca32_and_31_7[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7[39] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[8] = u_CSAwallace_pg_rca32_and_0_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[9] = u_CSAwallace_pg_rca32_and_1_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[10] = u_CSAwallace_pg_rca32_and_2_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[11] = u_CSAwallace_pg_rca32_and_3_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[12] = u_CSAwallace_pg_rca32_and_4_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[13] = u_CSAwallace_pg_rca32_and_5_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[14] = u_CSAwallace_pg_rca32_and_6_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[15] = u_CSAwallace_pg_rca32_and_7_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[16] = u_CSAwallace_pg_rca32_and_8_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[17] = u_CSAwallace_pg_rca32_and_9_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[18] = u_CSAwallace_pg_rca32_and_10_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[19] = u_CSAwallace_pg_rca32_and_11_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[20] = u_CSAwallace_pg_rca32_and_12_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[21] = u_CSAwallace_pg_rca32_and_13_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[22] = u_CSAwallace_pg_rca32_and_14_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[23] = u_CSAwallace_pg_rca32_and_15_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[24] = u_CSAwallace_pg_rca32_and_16_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[25] = u_CSAwallace_pg_rca32_and_17_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[26] = u_CSAwallace_pg_rca32_and_18_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[27] = u_CSAwallace_pg_rca32_and_19_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[28] = u_CSAwallace_pg_rca32_and_20_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[29] = u_CSAwallace_pg_rca32_and_21_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[30] = u_CSAwallace_pg_rca32_and_22_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[31] = u_CSAwallace_pg_rca32_and_23_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[32] = u_CSAwallace_pg_rca32_and_24_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[33] = u_CSAwallace_pg_rca32_and_25_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[34] = u_CSAwallace_pg_rca32_and_26_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[35] = u_CSAwallace_pg_rca32_and_27_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[36] = u_CSAwallace_pg_rca32_and_28_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[37] = u_CSAwallace_pg_rca32_and_29_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[38] = u_CSAwallace_pg_rca32_and_30_8[0];
  assign u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8[39] = u_CSAwallace_pg_rca32_and_31_8[0];
  csa_component40 csa_component40_u_CSAwallace_pg_rca32_csa2_csa_component_out(.a(u_CSAwallace_pg_rca32_csa2_csa_component_pp_row6), .b(u_CSAwallace_pg_rca32_csa2_csa_component_pp_row7), .c(u_CSAwallace_pg_rca32_csa2_csa_component_pp_row8), .csa_component40_out(u_CSAwallace_pg_rca32_csa2_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[9] = u_CSAwallace_pg_rca32_and_0_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[10] = u_CSAwallace_pg_rca32_and_1_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[11] = u_CSAwallace_pg_rca32_and_2_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[12] = u_CSAwallace_pg_rca32_and_3_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[13] = u_CSAwallace_pg_rca32_and_4_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[14] = u_CSAwallace_pg_rca32_and_5_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[15] = u_CSAwallace_pg_rca32_and_6_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[16] = u_CSAwallace_pg_rca32_and_7_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[17] = u_CSAwallace_pg_rca32_and_8_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[18] = u_CSAwallace_pg_rca32_and_9_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[19] = u_CSAwallace_pg_rca32_and_10_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[20] = u_CSAwallace_pg_rca32_and_11_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[21] = u_CSAwallace_pg_rca32_and_12_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[22] = u_CSAwallace_pg_rca32_and_13_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[23] = u_CSAwallace_pg_rca32_and_14_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[24] = u_CSAwallace_pg_rca32_and_15_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[25] = u_CSAwallace_pg_rca32_and_16_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[26] = u_CSAwallace_pg_rca32_and_17_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[27] = u_CSAwallace_pg_rca32_and_18_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[28] = u_CSAwallace_pg_rca32_and_19_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[29] = u_CSAwallace_pg_rca32_and_20_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[30] = u_CSAwallace_pg_rca32_and_21_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[31] = u_CSAwallace_pg_rca32_and_22_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[32] = u_CSAwallace_pg_rca32_and_23_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[33] = u_CSAwallace_pg_rca32_and_24_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[34] = u_CSAwallace_pg_rca32_and_25_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[35] = u_CSAwallace_pg_rca32_and_26_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[36] = u_CSAwallace_pg_rca32_and_27_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[37] = u_CSAwallace_pg_rca32_and_28_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[38] = u_CSAwallace_pg_rca32_and_29_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[39] = u_CSAwallace_pg_rca32_and_30_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[40] = u_CSAwallace_pg_rca32_and_31_9[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[41] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9[42] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[10] = u_CSAwallace_pg_rca32_and_0_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[11] = u_CSAwallace_pg_rca32_and_1_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[12] = u_CSAwallace_pg_rca32_and_2_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[13] = u_CSAwallace_pg_rca32_and_3_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[14] = u_CSAwallace_pg_rca32_and_4_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[15] = u_CSAwallace_pg_rca32_and_5_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[16] = u_CSAwallace_pg_rca32_and_6_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[17] = u_CSAwallace_pg_rca32_and_7_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[18] = u_CSAwallace_pg_rca32_and_8_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[19] = u_CSAwallace_pg_rca32_and_9_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[20] = u_CSAwallace_pg_rca32_and_10_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[21] = u_CSAwallace_pg_rca32_and_11_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[22] = u_CSAwallace_pg_rca32_and_12_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[23] = u_CSAwallace_pg_rca32_and_13_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[24] = u_CSAwallace_pg_rca32_and_14_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[25] = u_CSAwallace_pg_rca32_and_15_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[26] = u_CSAwallace_pg_rca32_and_16_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[27] = u_CSAwallace_pg_rca32_and_17_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[28] = u_CSAwallace_pg_rca32_and_18_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[29] = u_CSAwallace_pg_rca32_and_19_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[30] = u_CSAwallace_pg_rca32_and_20_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[31] = u_CSAwallace_pg_rca32_and_21_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[32] = u_CSAwallace_pg_rca32_and_22_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[33] = u_CSAwallace_pg_rca32_and_23_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[34] = u_CSAwallace_pg_rca32_and_24_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[35] = u_CSAwallace_pg_rca32_and_25_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[36] = u_CSAwallace_pg_rca32_and_26_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[37] = u_CSAwallace_pg_rca32_and_27_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[38] = u_CSAwallace_pg_rca32_and_28_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[39] = u_CSAwallace_pg_rca32_and_29_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[40] = u_CSAwallace_pg_rca32_and_30_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[41] = u_CSAwallace_pg_rca32_and_31_10[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10[42] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[11] = u_CSAwallace_pg_rca32_and_0_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[12] = u_CSAwallace_pg_rca32_and_1_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[13] = u_CSAwallace_pg_rca32_and_2_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[14] = u_CSAwallace_pg_rca32_and_3_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[15] = u_CSAwallace_pg_rca32_and_4_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[16] = u_CSAwallace_pg_rca32_and_5_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[17] = u_CSAwallace_pg_rca32_and_6_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[18] = u_CSAwallace_pg_rca32_and_7_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[19] = u_CSAwallace_pg_rca32_and_8_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[20] = u_CSAwallace_pg_rca32_and_9_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[21] = u_CSAwallace_pg_rca32_and_10_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[22] = u_CSAwallace_pg_rca32_and_11_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[23] = u_CSAwallace_pg_rca32_and_12_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[24] = u_CSAwallace_pg_rca32_and_13_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[25] = u_CSAwallace_pg_rca32_and_14_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[26] = u_CSAwallace_pg_rca32_and_15_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[27] = u_CSAwallace_pg_rca32_and_16_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[28] = u_CSAwallace_pg_rca32_and_17_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[29] = u_CSAwallace_pg_rca32_and_18_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[30] = u_CSAwallace_pg_rca32_and_19_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[31] = u_CSAwallace_pg_rca32_and_20_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[32] = u_CSAwallace_pg_rca32_and_21_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[33] = u_CSAwallace_pg_rca32_and_22_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[34] = u_CSAwallace_pg_rca32_and_23_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[35] = u_CSAwallace_pg_rca32_and_24_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[36] = u_CSAwallace_pg_rca32_and_25_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[37] = u_CSAwallace_pg_rca32_and_26_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[38] = u_CSAwallace_pg_rca32_and_27_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[39] = u_CSAwallace_pg_rca32_and_28_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[40] = u_CSAwallace_pg_rca32_and_29_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[41] = u_CSAwallace_pg_rca32_and_30_11[0];
  assign u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11[42] = u_CSAwallace_pg_rca32_and_31_11[0];
  csa_component43 csa_component43_u_CSAwallace_pg_rca32_csa3_csa_component_out(.a(u_CSAwallace_pg_rca32_csa3_csa_component_pp_row9), .b(u_CSAwallace_pg_rca32_csa3_csa_component_pp_row10), .c(u_CSAwallace_pg_rca32_csa3_csa_component_pp_row11), .csa_component43_out(u_CSAwallace_pg_rca32_csa3_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[12] = u_CSAwallace_pg_rca32_and_0_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[13] = u_CSAwallace_pg_rca32_and_1_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[14] = u_CSAwallace_pg_rca32_and_2_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[15] = u_CSAwallace_pg_rca32_and_3_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[16] = u_CSAwallace_pg_rca32_and_4_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[17] = u_CSAwallace_pg_rca32_and_5_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[18] = u_CSAwallace_pg_rca32_and_6_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[19] = u_CSAwallace_pg_rca32_and_7_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[20] = u_CSAwallace_pg_rca32_and_8_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[21] = u_CSAwallace_pg_rca32_and_9_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[22] = u_CSAwallace_pg_rca32_and_10_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[23] = u_CSAwallace_pg_rca32_and_11_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[24] = u_CSAwallace_pg_rca32_and_12_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[25] = u_CSAwallace_pg_rca32_and_13_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[26] = u_CSAwallace_pg_rca32_and_14_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[27] = u_CSAwallace_pg_rca32_and_15_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[28] = u_CSAwallace_pg_rca32_and_16_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[29] = u_CSAwallace_pg_rca32_and_17_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[30] = u_CSAwallace_pg_rca32_and_18_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[31] = u_CSAwallace_pg_rca32_and_19_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[32] = u_CSAwallace_pg_rca32_and_20_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[33] = u_CSAwallace_pg_rca32_and_21_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[34] = u_CSAwallace_pg_rca32_and_22_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[35] = u_CSAwallace_pg_rca32_and_23_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[36] = u_CSAwallace_pg_rca32_and_24_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[37] = u_CSAwallace_pg_rca32_and_25_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[38] = u_CSAwallace_pg_rca32_and_26_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[39] = u_CSAwallace_pg_rca32_and_27_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[40] = u_CSAwallace_pg_rca32_and_28_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[41] = u_CSAwallace_pg_rca32_and_29_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[42] = u_CSAwallace_pg_rca32_and_30_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[43] = u_CSAwallace_pg_rca32_and_31_12[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[44] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[13] = u_CSAwallace_pg_rca32_and_0_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[14] = u_CSAwallace_pg_rca32_and_1_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[15] = u_CSAwallace_pg_rca32_and_2_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[16] = u_CSAwallace_pg_rca32_and_3_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[17] = u_CSAwallace_pg_rca32_and_4_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[18] = u_CSAwallace_pg_rca32_and_5_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[19] = u_CSAwallace_pg_rca32_and_6_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[20] = u_CSAwallace_pg_rca32_and_7_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[21] = u_CSAwallace_pg_rca32_and_8_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[22] = u_CSAwallace_pg_rca32_and_9_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[23] = u_CSAwallace_pg_rca32_and_10_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[24] = u_CSAwallace_pg_rca32_and_11_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[25] = u_CSAwallace_pg_rca32_and_12_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[26] = u_CSAwallace_pg_rca32_and_13_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[27] = u_CSAwallace_pg_rca32_and_14_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[28] = u_CSAwallace_pg_rca32_and_15_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[29] = u_CSAwallace_pg_rca32_and_16_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[30] = u_CSAwallace_pg_rca32_and_17_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[31] = u_CSAwallace_pg_rca32_and_18_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[32] = u_CSAwallace_pg_rca32_and_19_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[33] = u_CSAwallace_pg_rca32_and_20_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[34] = u_CSAwallace_pg_rca32_and_21_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[35] = u_CSAwallace_pg_rca32_and_22_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[36] = u_CSAwallace_pg_rca32_and_23_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[37] = u_CSAwallace_pg_rca32_and_24_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[38] = u_CSAwallace_pg_rca32_and_25_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[39] = u_CSAwallace_pg_rca32_and_26_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[40] = u_CSAwallace_pg_rca32_and_27_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[41] = u_CSAwallace_pg_rca32_and_28_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[42] = u_CSAwallace_pg_rca32_and_29_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[43] = u_CSAwallace_pg_rca32_and_30_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[44] = u_CSAwallace_pg_rca32_and_31_13[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[14] = u_CSAwallace_pg_rca32_and_0_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[15] = u_CSAwallace_pg_rca32_and_1_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[16] = u_CSAwallace_pg_rca32_and_2_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[17] = u_CSAwallace_pg_rca32_and_3_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[18] = u_CSAwallace_pg_rca32_and_4_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[19] = u_CSAwallace_pg_rca32_and_5_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[20] = u_CSAwallace_pg_rca32_and_6_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[21] = u_CSAwallace_pg_rca32_and_7_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[22] = u_CSAwallace_pg_rca32_and_8_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[23] = u_CSAwallace_pg_rca32_and_9_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[24] = u_CSAwallace_pg_rca32_and_10_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[25] = u_CSAwallace_pg_rca32_and_11_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[26] = u_CSAwallace_pg_rca32_and_12_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[27] = u_CSAwallace_pg_rca32_and_13_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[28] = u_CSAwallace_pg_rca32_and_14_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[29] = u_CSAwallace_pg_rca32_and_15_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[30] = u_CSAwallace_pg_rca32_and_16_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[31] = u_CSAwallace_pg_rca32_and_17_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[32] = u_CSAwallace_pg_rca32_and_18_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[33] = u_CSAwallace_pg_rca32_and_19_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[34] = u_CSAwallace_pg_rca32_and_20_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[35] = u_CSAwallace_pg_rca32_and_21_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[36] = u_CSAwallace_pg_rca32_and_22_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[37] = u_CSAwallace_pg_rca32_and_23_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[38] = u_CSAwallace_pg_rca32_and_24_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[39] = u_CSAwallace_pg_rca32_and_25_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[40] = u_CSAwallace_pg_rca32_and_26_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[41] = u_CSAwallace_pg_rca32_and_27_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[42] = u_CSAwallace_pg_rca32_and_28_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[43] = u_CSAwallace_pg_rca32_and_29_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[44] = u_CSAwallace_pg_rca32_and_30_14[0];
  assign u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14[45] = u_CSAwallace_pg_rca32_and_31_14[0];
  csa_component46 csa_component46_u_CSAwallace_pg_rca32_csa4_csa_component_out(.a(u_CSAwallace_pg_rca32_csa4_csa_component_pp_row12), .b(u_CSAwallace_pg_rca32_csa4_csa_component_pp_row13), .c(u_CSAwallace_pg_rca32_csa4_csa_component_pp_row14), .csa_component46_out(u_CSAwallace_pg_rca32_csa4_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[15] = u_CSAwallace_pg_rca32_and_0_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[16] = u_CSAwallace_pg_rca32_and_1_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[17] = u_CSAwallace_pg_rca32_and_2_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[18] = u_CSAwallace_pg_rca32_and_3_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[19] = u_CSAwallace_pg_rca32_and_4_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[20] = u_CSAwallace_pg_rca32_and_5_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[21] = u_CSAwallace_pg_rca32_and_6_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[22] = u_CSAwallace_pg_rca32_and_7_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[23] = u_CSAwallace_pg_rca32_and_8_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[24] = u_CSAwallace_pg_rca32_and_9_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[25] = u_CSAwallace_pg_rca32_and_10_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[26] = u_CSAwallace_pg_rca32_and_11_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[27] = u_CSAwallace_pg_rca32_and_12_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[28] = u_CSAwallace_pg_rca32_and_13_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[29] = u_CSAwallace_pg_rca32_and_14_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[30] = u_CSAwallace_pg_rca32_and_15_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[31] = u_CSAwallace_pg_rca32_and_16_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[32] = u_CSAwallace_pg_rca32_and_17_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[33] = u_CSAwallace_pg_rca32_and_18_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[34] = u_CSAwallace_pg_rca32_and_19_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[35] = u_CSAwallace_pg_rca32_and_20_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[36] = u_CSAwallace_pg_rca32_and_21_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[37] = u_CSAwallace_pg_rca32_and_22_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[38] = u_CSAwallace_pg_rca32_and_23_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[39] = u_CSAwallace_pg_rca32_and_24_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[40] = u_CSAwallace_pg_rca32_and_25_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[41] = u_CSAwallace_pg_rca32_and_26_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[42] = u_CSAwallace_pg_rca32_and_27_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[43] = u_CSAwallace_pg_rca32_and_28_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[44] = u_CSAwallace_pg_rca32_and_29_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[45] = u_CSAwallace_pg_rca32_and_30_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[46] = u_CSAwallace_pg_rca32_and_31_15[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[16] = u_CSAwallace_pg_rca32_and_0_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[17] = u_CSAwallace_pg_rca32_and_1_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[18] = u_CSAwallace_pg_rca32_and_2_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[19] = u_CSAwallace_pg_rca32_and_3_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[20] = u_CSAwallace_pg_rca32_and_4_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[21] = u_CSAwallace_pg_rca32_and_5_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[22] = u_CSAwallace_pg_rca32_and_6_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[23] = u_CSAwallace_pg_rca32_and_7_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[24] = u_CSAwallace_pg_rca32_and_8_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[25] = u_CSAwallace_pg_rca32_and_9_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[26] = u_CSAwallace_pg_rca32_and_10_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[27] = u_CSAwallace_pg_rca32_and_11_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[28] = u_CSAwallace_pg_rca32_and_12_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[29] = u_CSAwallace_pg_rca32_and_13_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[30] = u_CSAwallace_pg_rca32_and_14_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[31] = u_CSAwallace_pg_rca32_and_15_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[32] = u_CSAwallace_pg_rca32_and_16_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[33] = u_CSAwallace_pg_rca32_and_17_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[34] = u_CSAwallace_pg_rca32_and_18_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[35] = u_CSAwallace_pg_rca32_and_19_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[36] = u_CSAwallace_pg_rca32_and_20_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[37] = u_CSAwallace_pg_rca32_and_21_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[38] = u_CSAwallace_pg_rca32_and_22_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[39] = u_CSAwallace_pg_rca32_and_23_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[40] = u_CSAwallace_pg_rca32_and_24_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[41] = u_CSAwallace_pg_rca32_and_25_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[42] = u_CSAwallace_pg_rca32_and_26_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[43] = u_CSAwallace_pg_rca32_and_27_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[44] = u_CSAwallace_pg_rca32_and_28_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[45] = u_CSAwallace_pg_rca32_and_29_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[46] = u_CSAwallace_pg_rca32_and_30_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[47] = u_CSAwallace_pg_rca32_and_31_16[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[17] = u_CSAwallace_pg_rca32_and_0_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[18] = u_CSAwallace_pg_rca32_and_1_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[19] = u_CSAwallace_pg_rca32_and_2_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[20] = u_CSAwallace_pg_rca32_and_3_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[21] = u_CSAwallace_pg_rca32_and_4_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[22] = u_CSAwallace_pg_rca32_and_5_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[23] = u_CSAwallace_pg_rca32_and_6_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[24] = u_CSAwallace_pg_rca32_and_7_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[25] = u_CSAwallace_pg_rca32_and_8_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[26] = u_CSAwallace_pg_rca32_and_9_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[27] = u_CSAwallace_pg_rca32_and_10_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[28] = u_CSAwallace_pg_rca32_and_11_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[29] = u_CSAwallace_pg_rca32_and_12_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[30] = u_CSAwallace_pg_rca32_and_13_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[31] = u_CSAwallace_pg_rca32_and_14_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[32] = u_CSAwallace_pg_rca32_and_15_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[33] = u_CSAwallace_pg_rca32_and_16_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[34] = u_CSAwallace_pg_rca32_and_17_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[35] = u_CSAwallace_pg_rca32_and_18_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[36] = u_CSAwallace_pg_rca32_and_19_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[37] = u_CSAwallace_pg_rca32_and_20_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[38] = u_CSAwallace_pg_rca32_and_21_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[39] = u_CSAwallace_pg_rca32_and_22_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[40] = u_CSAwallace_pg_rca32_and_23_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[41] = u_CSAwallace_pg_rca32_and_24_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[42] = u_CSAwallace_pg_rca32_and_25_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[43] = u_CSAwallace_pg_rca32_and_26_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[44] = u_CSAwallace_pg_rca32_and_27_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[45] = u_CSAwallace_pg_rca32_and_28_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[46] = u_CSAwallace_pg_rca32_and_29_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[47] = u_CSAwallace_pg_rca32_and_30_17[0];
  assign u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17[48] = u_CSAwallace_pg_rca32_and_31_17[0];
  csa_component49 csa_component49_u_CSAwallace_pg_rca32_csa5_csa_component_out(.a(u_CSAwallace_pg_rca32_csa5_csa_component_pp_row15), .b(u_CSAwallace_pg_rca32_csa5_csa_component_pp_row16), .c(u_CSAwallace_pg_rca32_csa5_csa_component_pp_row17), .csa_component49_out(u_CSAwallace_pg_rca32_csa5_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[18] = u_CSAwallace_pg_rca32_and_0_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[19] = u_CSAwallace_pg_rca32_and_1_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[20] = u_CSAwallace_pg_rca32_and_2_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[21] = u_CSAwallace_pg_rca32_and_3_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[22] = u_CSAwallace_pg_rca32_and_4_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[23] = u_CSAwallace_pg_rca32_and_5_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[24] = u_CSAwallace_pg_rca32_and_6_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[25] = u_CSAwallace_pg_rca32_and_7_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[26] = u_CSAwallace_pg_rca32_and_8_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[27] = u_CSAwallace_pg_rca32_and_9_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[28] = u_CSAwallace_pg_rca32_and_10_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[29] = u_CSAwallace_pg_rca32_and_11_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[30] = u_CSAwallace_pg_rca32_and_12_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[31] = u_CSAwallace_pg_rca32_and_13_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[32] = u_CSAwallace_pg_rca32_and_14_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[33] = u_CSAwallace_pg_rca32_and_15_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[34] = u_CSAwallace_pg_rca32_and_16_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[35] = u_CSAwallace_pg_rca32_and_17_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[36] = u_CSAwallace_pg_rca32_and_18_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[37] = u_CSAwallace_pg_rca32_and_19_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[38] = u_CSAwallace_pg_rca32_and_20_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[39] = u_CSAwallace_pg_rca32_and_21_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[40] = u_CSAwallace_pg_rca32_and_22_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[41] = u_CSAwallace_pg_rca32_and_23_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[42] = u_CSAwallace_pg_rca32_and_24_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[43] = u_CSAwallace_pg_rca32_and_25_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[44] = u_CSAwallace_pg_rca32_and_26_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[45] = u_CSAwallace_pg_rca32_and_27_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[46] = u_CSAwallace_pg_rca32_and_28_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[47] = u_CSAwallace_pg_rca32_and_29_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[48] = u_CSAwallace_pg_rca32_and_30_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[49] = u_CSAwallace_pg_rca32_and_31_18[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[50] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[19] = u_CSAwallace_pg_rca32_and_0_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[20] = u_CSAwallace_pg_rca32_and_1_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[21] = u_CSAwallace_pg_rca32_and_2_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[22] = u_CSAwallace_pg_rca32_and_3_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[23] = u_CSAwallace_pg_rca32_and_4_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[24] = u_CSAwallace_pg_rca32_and_5_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[25] = u_CSAwallace_pg_rca32_and_6_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[26] = u_CSAwallace_pg_rca32_and_7_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[27] = u_CSAwallace_pg_rca32_and_8_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[28] = u_CSAwallace_pg_rca32_and_9_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[29] = u_CSAwallace_pg_rca32_and_10_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[30] = u_CSAwallace_pg_rca32_and_11_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[31] = u_CSAwallace_pg_rca32_and_12_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[32] = u_CSAwallace_pg_rca32_and_13_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[33] = u_CSAwallace_pg_rca32_and_14_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[34] = u_CSAwallace_pg_rca32_and_15_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[35] = u_CSAwallace_pg_rca32_and_16_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[36] = u_CSAwallace_pg_rca32_and_17_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[37] = u_CSAwallace_pg_rca32_and_18_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[38] = u_CSAwallace_pg_rca32_and_19_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[39] = u_CSAwallace_pg_rca32_and_20_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[40] = u_CSAwallace_pg_rca32_and_21_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[41] = u_CSAwallace_pg_rca32_and_22_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[42] = u_CSAwallace_pg_rca32_and_23_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[43] = u_CSAwallace_pg_rca32_and_24_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[44] = u_CSAwallace_pg_rca32_and_25_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[45] = u_CSAwallace_pg_rca32_and_26_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[46] = u_CSAwallace_pg_rca32_and_27_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[47] = u_CSAwallace_pg_rca32_and_28_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[48] = u_CSAwallace_pg_rca32_and_29_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[49] = u_CSAwallace_pg_rca32_and_30_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[50] = u_CSAwallace_pg_rca32_and_31_19[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[20] = u_CSAwallace_pg_rca32_and_0_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[21] = u_CSAwallace_pg_rca32_and_1_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[22] = u_CSAwallace_pg_rca32_and_2_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[23] = u_CSAwallace_pg_rca32_and_3_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[24] = u_CSAwallace_pg_rca32_and_4_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[25] = u_CSAwallace_pg_rca32_and_5_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[26] = u_CSAwallace_pg_rca32_and_6_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[27] = u_CSAwallace_pg_rca32_and_7_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[28] = u_CSAwallace_pg_rca32_and_8_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[29] = u_CSAwallace_pg_rca32_and_9_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[30] = u_CSAwallace_pg_rca32_and_10_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[31] = u_CSAwallace_pg_rca32_and_11_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[32] = u_CSAwallace_pg_rca32_and_12_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[33] = u_CSAwallace_pg_rca32_and_13_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[34] = u_CSAwallace_pg_rca32_and_14_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[35] = u_CSAwallace_pg_rca32_and_15_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[36] = u_CSAwallace_pg_rca32_and_16_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[37] = u_CSAwallace_pg_rca32_and_17_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[38] = u_CSAwallace_pg_rca32_and_18_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[39] = u_CSAwallace_pg_rca32_and_19_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[40] = u_CSAwallace_pg_rca32_and_20_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[41] = u_CSAwallace_pg_rca32_and_21_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[42] = u_CSAwallace_pg_rca32_and_22_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[43] = u_CSAwallace_pg_rca32_and_23_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[44] = u_CSAwallace_pg_rca32_and_24_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[45] = u_CSAwallace_pg_rca32_and_25_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[46] = u_CSAwallace_pg_rca32_and_26_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[47] = u_CSAwallace_pg_rca32_and_27_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[48] = u_CSAwallace_pg_rca32_and_28_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[49] = u_CSAwallace_pg_rca32_and_29_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[50] = u_CSAwallace_pg_rca32_and_30_20[0];
  assign u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20[51] = u_CSAwallace_pg_rca32_and_31_20[0];
  csa_component52 csa_component52_u_CSAwallace_pg_rca32_csa6_csa_component_out(.a(u_CSAwallace_pg_rca32_csa6_csa_component_pp_row18), .b(u_CSAwallace_pg_rca32_csa6_csa_component_pp_row19), .c(u_CSAwallace_pg_rca32_csa6_csa_component_pp_row20), .csa_component52_out(u_CSAwallace_pg_rca32_csa6_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[21] = u_CSAwallace_pg_rca32_and_0_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[22] = u_CSAwallace_pg_rca32_and_1_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[23] = u_CSAwallace_pg_rca32_and_2_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[24] = u_CSAwallace_pg_rca32_and_3_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[25] = u_CSAwallace_pg_rca32_and_4_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[26] = u_CSAwallace_pg_rca32_and_5_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[27] = u_CSAwallace_pg_rca32_and_6_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[28] = u_CSAwallace_pg_rca32_and_7_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[29] = u_CSAwallace_pg_rca32_and_8_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[30] = u_CSAwallace_pg_rca32_and_9_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[31] = u_CSAwallace_pg_rca32_and_10_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[32] = u_CSAwallace_pg_rca32_and_11_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[33] = u_CSAwallace_pg_rca32_and_12_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[34] = u_CSAwallace_pg_rca32_and_13_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[35] = u_CSAwallace_pg_rca32_and_14_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[36] = u_CSAwallace_pg_rca32_and_15_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[37] = u_CSAwallace_pg_rca32_and_16_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[38] = u_CSAwallace_pg_rca32_and_17_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[39] = u_CSAwallace_pg_rca32_and_18_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[40] = u_CSAwallace_pg_rca32_and_19_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[41] = u_CSAwallace_pg_rca32_and_20_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[42] = u_CSAwallace_pg_rca32_and_21_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[43] = u_CSAwallace_pg_rca32_and_22_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[44] = u_CSAwallace_pg_rca32_and_23_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[45] = u_CSAwallace_pg_rca32_and_24_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[46] = u_CSAwallace_pg_rca32_and_25_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[47] = u_CSAwallace_pg_rca32_and_26_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[48] = u_CSAwallace_pg_rca32_and_27_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[49] = u_CSAwallace_pg_rca32_and_28_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[50] = u_CSAwallace_pg_rca32_and_29_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[51] = u_CSAwallace_pg_rca32_and_30_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[52] = u_CSAwallace_pg_rca32_and_31_21[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[22] = u_CSAwallace_pg_rca32_and_0_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[23] = u_CSAwallace_pg_rca32_and_1_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[24] = u_CSAwallace_pg_rca32_and_2_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[25] = u_CSAwallace_pg_rca32_and_3_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[26] = u_CSAwallace_pg_rca32_and_4_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[27] = u_CSAwallace_pg_rca32_and_5_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[28] = u_CSAwallace_pg_rca32_and_6_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[29] = u_CSAwallace_pg_rca32_and_7_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[30] = u_CSAwallace_pg_rca32_and_8_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[31] = u_CSAwallace_pg_rca32_and_9_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[32] = u_CSAwallace_pg_rca32_and_10_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[33] = u_CSAwallace_pg_rca32_and_11_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[34] = u_CSAwallace_pg_rca32_and_12_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[35] = u_CSAwallace_pg_rca32_and_13_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[36] = u_CSAwallace_pg_rca32_and_14_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[37] = u_CSAwallace_pg_rca32_and_15_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[38] = u_CSAwallace_pg_rca32_and_16_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[39] = u_CSAwallace_pg_rca32_and_17_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[40] = u_CSAwallace_pg_rca32_and_18_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[41] = u_CSAwallace_pg_rca32_and_19_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[42] = u_CSAwallace_pg_rca32_and_20_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[43] = u_CSAwallace_pg_rca32_and_21_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[44] = u_CSAwallace_pg_rca32_and_22_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[45] = u_CSAwallace_pg_rca32_and_23_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[46] = u_CSAwallace_pg_rca32_and_24_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[47] = u_CSAwallace_pg_rca32_and_25_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[48] = u_CSAwallace_pg_rca32_and_26_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[49] = u_CSAwallace_pg_rca32_and_27_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[50] = u_CSAwallace_pg_rca32_and_28_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[51] = u_CSAwallace_pg_rca32_and_29_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[52] = u_CSAwallace_pg_rca32_and_30_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[53] = u_CSAwallace_pg_rca32_and_31_22[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[23] = u_CSAwallace_pg_rca32_and_0_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[24] = u_CSAwallace_pg_rca32_and_1_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[25] = u_CSAwallace_pg_rca32_and_2_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[26] = u_CSAwallace_pg_rca32_and_3_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[27] = u_CSAwallace_pg_rca32_and_4_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[28] = u_CSAwallace_pg_rca32_and_5_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[29] = u_CSAwallace_pg_rca32_and_6_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[30] = u_CSAwallace_pg_rca32_and_7_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[31] = u_CSAwallace_pg_rca32_and_8_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[32] = u_CSAwallace_pg_rca32_and_9_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[33] = u_CSAwallace_pg_rca32_and_10_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[34] = u_CSAwallace_pg_rca32_and_11_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[35] = u_CSAwallace_pg_rca32_and_12_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[36] = u_CSAwallace_pg_rca32_and_13_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[37] = u_CSAwallace_pg_rca32_and_14_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[38] = u_CSAwallace_pg_rca32_and_15_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[39] = u_CSAwallace_pg_rca32_and_16_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[40] = u_CSAwallace_pg_rca32_and_17_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[41] = u_CSAwallace_pg_rca32_and_18_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[42] = u_CSAwallace_pg_rca32_and_19_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[43] = u_CSAwallace_pg_rca32_and_20_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[44] = u_CSAwallace_pg_rca32_and_21_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[45] = u_CSAwallace_pg_rca32_and_22_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[46] = u_CSAwallace_pg_rca32_and_23_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[47] = u_CSAwallace_pg_rca32_and_24_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[48] = u_CSAwallace_pg_rca32_and_25_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[49] = u_CSAwallace_pg_rca32_and_26_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[50] = u_CSAwallace_pg_rca32_and_27_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[51] = u_CSAwallace_pg_rca32_and_28_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[52] = u_CSAwallace_pg_rca32_and_29_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[53] = u_CSAwallace_pg_rca32_and_30_23[0];
  assign u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23[54] = u_CSAwallace_pg_rca32_and_31_23[0];
  csa_component55 csa_component55_u_CSAwallace_pg_rca32_csa7_csa_component_out(.a(u_CSAwallace_pg_rca32_csa7_csa_component_pp_row21), .b(u_CSAwallace_pg_rca32_csa7_csa_component_pp_row22), .c(u_CSAwallace_pg_rca32_csa7_csa_component_pp_row23), .csa_component55_out(u_CSAwallace_pg_rca32_csa7_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[24] = u_CSAwallace_pg_rca32_and_0_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[25] = u_CSAwallace_pg_rca32_and_1_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[26] = u_CSAwallace_pg_rca32_and_2_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[27] = u_CSAwallace_pg_rca32_and_3_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[28] = u_CSAwallace_pg_rca32_and_4_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[29] = u_CSAwallace_pg_rca32_and_5_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[30] = u_CSAwallace_pg_rca32_and_6_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[31] = u_CSAwallace_pg_rca32_and_7_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[32] = u_CSAwallace_pg_rca32_and_8_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[33] = u_CSAwallace_pg_rca32_and_9_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[34] = u_CSAwallace_pg_rca32_and_10_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[35] = u_CSAwallace_pg_rca32_and_11_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[36] = u_CSAwallace_pg_rca32_and_12_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[37] = u_CSAwallace_pg_rca32_and_13_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[38] = u_CSAwallace_pg_rca32_and_14_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[39] = u_CSAwallace_pg_rca32_and_15_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[40] = u_CSAwallace_pg_rca32_and_16_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[41] = u_CSAwallace_pg_rca32_and_17_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[42] = u_CSAwallace_pg_rca32_and_18_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[43] = u_CSAwallace_pg_rca32_and_19_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[44] = u_CSAwallace_pg_rca32_and_20_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[45] = u_CSAwallace_pg_rca32_and_21_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[46] = u_CSAwallace_pg_rca32_and_22_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[47] = u_CSAwallace_pg_rca32_and_23_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[48] = u_CSAwallace_pg_rca32_and_24_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[49] = u_CSAwallace_pg_rca32_and_25_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[50] = u_CSAwallace_pg_rca32_and_26_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[51] = u_CSAwallace_pg_rca32_and_27_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[52] = u_CSAwallace_pg_rca32_and_28_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[53] = u_CSAwallace_pg_rca32_and_29_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[54] = u_CSAwallace_pg_rca32_and_30_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[55] = u_CSAwallace_pg_rca32_and_31_24[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[25] = u_CSAwallace_pg_rca32_and_0_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[26] = u_CSAwallace_pg_rca32_and_1_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[27] = u_CSAwallace_pg_rca32_and_2_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[28] = u_CSAwallace_pg_rca32_and_3_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[29] = u_CSAwallace_pg_rca32_and_4_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[30] = u_CSAwallace_pg_rca32_and_5_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[31] = u_CSAwallace_pg_rca32_and_6_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[32] = u_CSAwallace_pg_rca32_and_7_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[33] = u_CSAwallace_pg_rca32_and_8_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[34] = u_CSAwallace_pg_rca32_and_9_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[35] = u_CSAwallace_pg_rca32_and_10_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[36] = u_CSAwallace_pg_rca32_and_11_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[37] = u_CSAwallace_pg_rca32_and_12_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[38] = u_CSAwallace_pg_rca32_and_13_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[39] = u_CSAwallace_pg_rca32_and_14_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[40] = u_CSAwallace_pg_rca32_and_15_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[41] = u_CSAwallace_pg_rca32_and_16_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[42] = u_CSAwallace_pg_rca32_and_17_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[43] = u_CSAwallace_pg_rca32_and_18_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[44] = u_CSAwallace_pg_rca32_and_19_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[45] = u_CSAwallace_pg_rca32_and_20_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[46] = u_CSAwallace_pg_rca32_and_21_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[47] = u_CSAwallace_pg_rca32_and_22_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[48] = u_CSAwallace_pg_rca32_and_23_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[49] = u_CSAwallace_pg_rca32_and_24_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[50] = u_CSAwallace_pg_rca32_and_25_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[51] = u_CSAwallace_pg_rca32_and_26_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[52] = u_CSAwallace_pg_rca32_and_27_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[53] = u_CSAwallace_pg_rca32_and_28_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[54] = u_CSAwallace_pg_rca32_and_29_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[55] = u_CSAwallace_pg_rca32_and_30_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[56] = u_CSAwallace_pg_rca32_and_31_25[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[26] = u_CSAwallace_pg_rca32_and_0_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[27] = u_CSAwallace_pg_rca32_and_1_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[28] = u_CSAwallace_pg_rca32_and_2_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[29] = u_CSAwallace_pg_rca32_and_3_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[30] = u_CSAwallace_pg_rca32_and_4_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[31] = u_CSAwallace_pg_rca32_and_5_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[32] = u_CSAwallace_pg_rca32_and_6_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[33] = u_CSAwallace_pg_rca32_and_7_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[34] = u_CSAwallace_pg_rca32_and_8_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[35] = u_CSAwallace_pg_rca32_and_9_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[36] = u_CSAwallace_pg_rca32_and_10_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[37] = u_CSAwallace_pg_rca32_and_11_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[38] = u_CSAwallace_pg_rca32_and_12_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[39] = u_CSAwallace_pg_rca32_and_13_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[40] = u_CSAwallace_pg_rca32_and_14_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[41] = u_CSAwallace_pg_rca32_and_15_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[42] = u_CSAwallace_pg_rca32_and_16_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[43] = u_CSAwallace_pg_rca32_and_17_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[44] = u_CSAwallace_pg_rca32_and_18_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[45] = u_CSAwallace_pg_rca32_and_19_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[46] = u_CSAwallace_pg_rca32_and_20_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[47] = u_CSAwallace_pg_rca32_and_21_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[48] = u_CSAwallace_pg_rca32_and_22_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[49] = u_CSAwallace_pg_rca32_and_23_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[50] = u_CSAwallace_pg_rca32_and_24_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[51] = u_CSAwallace_pg_rca32_and_25_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[52] = u_CSAwallace_pg_rca32_and_26_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[53] = u_CSAwallace_pg_rca32_and_27_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[54] = u_CSAwallace_pg_rca32_and_28_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[55] = u_CSAwallace_pg_rca32_and_29_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[56] = u_CSAwallace_pg_rca32_and_30_26[0];
  assign u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26[57] = u_CSAwallace_pg_rca32_and_31_26[0];
  csa_component58 csa_component58_u_CSAwallace_pg_rca32_csa8_csa_component_out(.a(u_CSAwallace_pg_rca32_csa8_csa_component_pp_row24), .b(u_CSAwallace_pg_rca32_csa8_csa_component_pp_row25), .c(u_CSAwallace_pg_rca32_csa8_csa_component_pp_row26), .csa_component58_out(u_CSAwallace_pg_rca32_csa8_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[27] = u_CSAwallace_pg_rca32_and_0_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[28] = u_CSAwallace_pg_rca32_and_1_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[29] = u_CSAwallace_pg_rca32_and_2_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[30] = u_CSAwallace_pg_rca32_and_3_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[31] = u_CSAwallace_pg_rca32_and_4_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[32] = u_CSAwallace_pg_rca32_and_5_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[33] = u_CSAwallace_pg_rca32_and_6_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[34] = u_CSAwallace_pg_rca32_and_7_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[35] = u_CSAwallace_pg_rca32_and_8_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[36] = u_CSAwallace_pg_rca32_and_9_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[37] = u_CSAwallace_pg_rca32_and_10_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[38] = u_CSAwallace_pg_rca32_and_11_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[39] = u_CSAwallace_pg_rca32_and_12_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[40] = u_CSAwallace_pg_rca32_and_13_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[41] = u_CSAwallace_pg_rca32_and_14_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[42] = u_CSAwallace_pg_rca32_and_15_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[43] = u_CSAwallace_pg_rca32_and_16_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[44] = u_CSAwallace_pg_rca32_and_17_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[45] = u_CSAwallace_pg_rca32_and_18_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[46] = u_CSAwallace_pg_rca32_and_19_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[47] = u_CSAwallace_pg_rca32_and_20_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[48] = u_CSAwallace_pg_rca32_and_21_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[49] = u_CSAwallace_pg_rca32_and_22_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[50] = u_CSAwallace_pg_rca32_and_23_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[51] = u_CSAwallace_pg_rca32_and_24_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[52] = u_CSAwallace_pg_rca32_and_25_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[53] = u_CSAwallace_pg_rca32_and_26_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[54] = u_CSAwallace_pg_rca32_and_27_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[55] = u_CSAwallace_pg_rca32_and_28_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[56] = u_CSAwallace_pg_rca32_and_29_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[57] = u_CSAwallace_pg_rca32_and_30_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[58] = u_CSAwallace_pg_rca32_and_31_27[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[27] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[28] = u_CSAwallace_pg_rca32_and_0_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[29] = u_CSAwallace_pg_rca32_and_1_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[30] = u_CSAwallace_pg_rca32_and_2_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[31] = u_CSAwallace_pg_rca32_and_3_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[32] = u_CSAwallace_pg_rca32_and_4_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[33] = u_CSAwallace_pg_rca32_and_5_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[34] = u_CSAwallace_pg_rca32_and_6_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[35] = u_CSAwallace_pg_rca32_and_7_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[36] = u_CSAwallace_pg_rca32_and_8_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[37] = u_CSAwallace_pg_rca32_and_9_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[38] = u_CSAwallace_pg_rca32_and_10_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[39] = u_CSAwallace_pg_rca32_and_11_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[40] = u_CSAwallace_pg_rca32_and_12_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[41] = u_CSAwallace_pg_rca32_and_13_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[42] = u_CSAwallace_pg_rca32_and_14_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[43] = u_CSAwallace_pg_rca32_and_15_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[44] = u_CSAwallace_pg_rca32_and_16_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[45] = u_CSAwallace_pg_rca32_and_17_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[46] = u_CSAwallace_pg_rca32_and_18_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[47] = u_CSAwallace_pg_rca32_and_19_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[48] = u_CSAwallace_pg_rca32_and_20_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[49] = u_CSAwallace_pg_rca32_and_21_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[50] = u_CSAwallace_pg_rca32_and_22_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[51] = u_CSAwallace_pg_rca32_and_23_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[52] = u_CSAwallace_pg_rca32_and_24_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[53] = u_CSAwallace_pg_rca32_and_25_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[54] = u_CSAwallace_pg_rca32_and_26_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[55] = u_CSAwallace_pg_rca32_and_27_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[56] = u_CSAwallace_pg_rca32_and_28_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[57] = u_CSAwallace_pg_rca32_and_29_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[58] = u_CSAwallace_pg_rca32_and_30_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[59] = u_CSAwallace_pg_rca32_and_31_28[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[27] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[28] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[29] = u_CSAwallace_pg_rca32_and_0_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[30] = u_CSAwallace_pg_rca32_and_1_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[31] = u_CSAwallace_pg_rca32_and_2_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[32] = u_CSAwallace_pg_rca32_and_3_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[33] = u_CSAwallace_pg_rca32_and_4_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[34] = u_CSAwallace_pg_rca32_and_5_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[35] = u_CSAwallace_pg_rca32_and_6_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[36] = u_CSAwallace_pg_rca32_and_7_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[37] = u_CSAwallace_pg_rca32_and_8_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[38] = u_CSAwallace_pg_rca32_and_9_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[39] = u_CSAwallace_pg_rca32_and_10_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[40] = u_CSAwallace_pg_rca32_and_11_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[41] = u_CSAwallace_pg_rca32_and_12_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[42] = u_CSAwallace_pg_rca32_and_13_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[43] = u_CSAwallace_pg_rca32_and_14_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[44] = u_CSAwallace_pg_rca32_and_15_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[45] = u_CSAwallace_pg_rca32_and_16_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[46] = u_CSAwallace_pg_rca32_and_17_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[47] = u_CSAwallace_pg_rca32_and_18_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[48] = u_CSAwallace_pg_rca32_and_19_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[49] = u_CSAwallace_pg_rca32_and_20_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[50] = u_CSAwallace_pg_rca32_and_21_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[51] = u_CSAwallace_pg_rca32_and_22_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[52] = u_CSAwallace_pg_rca32_and_23_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[53] = u_CSAwallace_pg_rca32_and_24_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[54] = u_CSAwallace_pg_rca32_and_25_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[55] = u_CSAwallace_pg_rca32_and_26_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[56] = u_CSAwallace_pg_rca32_and_27_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[57] = u_CSAwallace_pg_rca32_and_28_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[58] = u_CSAwallace_pg_rca32_and_29_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[59] = u_CSAwallace_pg_rca32_and_30_29[0];
  assign u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29[60] = u_CSAwallace_pg_rca32_and_31_29[0];
  csa_component61 csa_component61_u_CSAwallace_pg_rca32_csa9_csa_component_out(.a(u_CSAwallace_pg_rca32_csa9_csa_component_pp_row27), .b(u_CSAwallace_pg_rca32_csa9_csa_component_pp_row28), .c(u_CSAwallace_pg_rca32_csa9_csa_component_pp_row29), .csa_component61_out(u_CSAwallace_pg_rca32_csa9_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[0] = u_CSAwallace_pg_rca32_csa0_csa_component_out[0];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[1] = u_CSAwallace_pg_rca32_csa0_csa_component_out[1];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[2] = u_CSAwallace_pg_rca32_csa0_csa_component_out[2];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[3] = u_CSAwallace_pg_rca32_csa0_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[4] = u_CSAwallace_pg_rca32_csa0_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[5] = u_CSAwallace_pg_rca32_csa0_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[6] = u_CSAwallace_pg_rca32_csa0_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[7] = u_CSAwallace_pg_rca32_csa0_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[8] = u_CSAwallace_pg_rca32_csa0_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[9] = u_CSAwallace_pg_rca32_csa0_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[10] = u_CSAwallace_pg_rca32_csa0_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[11] = u_CSAwallace_pg_rca32_csa0_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[12] = u_CSAwallace_pg_rca32_csa0_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[13] = u_CSAwallace_pg_rca32_csa0_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[14] = u_CSAwallace_pg_rca32_csa0_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[15] = u_CSAwallace_pg_rca32_csa0_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[16] = u_CSAwallace_pg_rca32_csa0_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[17] = u_CSAwallace_pg_rca32_csa0_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[18] = u_CSAwallace_pg_rca32_csa0_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[19] = u_CSAwallace_pg_rca32_csa0_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[20] = u_CSAwallace_pg_rca32_csa0_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[21] = u_CSAwallace_pg_rca32_csa0_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[22] = u_CSAwallace_pg_rca32_csa0_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[23] = u_CSAwallace_pg_rca32_csa0_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[24] = u_CSAwallace_pg_rca32_csa0_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[25] = u_CSAwallace_pg_rca32_csa0_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[26] = u_CSAwallace_pg_rca32_csa0_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[27] = u_CSAwallace_pg_rca32_csa0_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[28] = u_CSAwallace_pg_rca32_csa0_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[29] = u_CSAwallace_pg_rca32_csa0_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[30] = u_CSAwallace_pg_rca32_csa0_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[31] = u_CSAwallace_pg_rca32_csa0_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[32] = u_CSAwallace_pg_rca32_csa0_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[33] = u_CSAwallace_pg_rca32_csa0_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[34] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[35] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[36] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1[37] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[2] = u_CSAwallace_pg_rca32_csa0_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[3] = u_CSAwallace_pg_rca32_csa0_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[4] = u_CSAwallace_pg_rca32_csa0_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[5] = u_CSAwallace_pg_rca32_csa0_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[6] = u_CSAwallace_pg_rca32_csa0_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[7] = u_CSAwallace_pg_rca32_csa0_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[8] = u_CSAwallace_pg_rca32_csa0_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[9] = u_CSAwallace_pg_rca32_csa0_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[10] = u_CSAwallace_pg_rca32_csa0_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[11] = u_CSAwallace_pg_rca32_csa0_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[12] = u_CSAwallace_pg_rca32_csa0_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[13] = u_CSAwallace_pg_rca32_csa0_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[14] = u_CSAwallace_pg_rca32_csa0_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[15] = u_CSAwallace_pg_rca32_csa0_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[16] = u_CSAwallace_pg_rca32_csa0_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[17] = u_CSAwallace_pg_rca32_csa0_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[18] = u_CSAwallace_pg_rca32_csa0_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[19] = u_CSAwallace_pg_rca32_csa0_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[20] = u_CSAwallace_pg_rca32_csa0_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[21] = u_CSAwallace_pg_rca32_csa0_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[22] = u_CSAwallace_pg_rca32_csa0_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[23] = u_CSAwallace_pg_rca32_csa0_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[24] = u_CSAwallace_pg_rca32_csa0_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[25] = u_CSAwallace_pg_rca32_csa0_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[26] = u_CSAwallace_pg_rca32_csa0_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[27] = u_CSAwallace_pg_rca32_csa0_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[28] = u_CSAwallace_pg_rca32_csa0_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[29] = u_CSAwallace_pg_rca32_csa0_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[30] = u_CSAwallace_pg_rca32_csa0_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[31] = u_CSAwallace_pg_rca32_csa0_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[32] = u_CSAwallace_pg_rca32_csa0_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[33] = u_CSAwallace_pg_rca32_csa0_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[34] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[35] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[36] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1[37] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[3] = u_CSAwallace_pg_rca32_csa1_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[4] = u_CSAwallace_pg_rca32_csa1_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[5] = u_CSAwallace_pg_rca32_csa1_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[6] = u_CSAwallace_pg_rca32_csa1_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[7] = u_CSAwallace_pg_rca32_csa1_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[8] = u_CSAwallace_pg_rca32_csa1_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[9] = u_CSAwallace_pg_rca32_csa1_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[10] = u_CSAwallace_pg_rca32_csa1_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[11] = u_CSAwallace_pg_rca32_csa1_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[12] = u_CSAwallace_pg_rca32_csa1_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[13] = u_CSAwallace_pg_rca32_csa1_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[14] = u_CSAwallace_pg_rca32_csa1_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[15] = u_CSAwallace_pg_rca32_csa1_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[16] = u_CSAwallace_pg_rca32_csa1_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[17] = u_CSAwallace_pg_rca32_csa1_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[18] = u_CSAwallace_pg_rca32_csa1_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[19] = u_CSAwallace_pg_rca32_csa1_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[20] = u_CSAwallace_pg_rca32_csa1_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[21] = u_CSAwallace_pg_rca32_csa1_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[22] = u_CSAwallace_pg_rca32_csa1_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[23] = u_CSAwallace_pg_rca32_csa1_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[24] = u_CSAwallace_pg_rca32_csa1_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[25] = u_CSAwallace_pg_rca32_csa1_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[26] = u_CSAwallace_pg_rca32_csa1_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[27] = u_CSAwallace_pg_rca32_csa1_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[28] = u_CSAwallace_pg_rca32_csa1_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[29] = u_CSAwallace_pg_rca32_csa1_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[30] = u_CSAwallace_pg_rca32_csa1_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[31] = u_CSAwallace_pg_rca32_csa1_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[32] = u_CSAwallace_pg_rca32_csa1_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[33] = u_CSAwallace_pg_rca32_csa1_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[34] = u_CSAwallace_pg_rca32_csa1_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[35] = u_CSAwallace_pg_rca32_csa1_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[36] = u_CSAwallace_pg_rca32_csa1_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2[37] = 1'b0;
  csa_component38 csa_component38_u_CSAwallace_pg_rca32_csa10_csa_component_out(.a(u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s1), .b(u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_c1), .c(u_CSAwallace_pg_rca32_csa10_csa_component_u_CSAwallace_pg_rca32_csa_s2), .csa_component38_out(u_CSAwallace_pg_rca32_csa10_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[5] = u_CSAwallace_pg_rca32_csa1_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[6] = u_CSAwallace_pg_rca32_csa1_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[7] = u_CSAwallace_pg_rca32_csa1_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[8] = u_CSAwallace_pg_rca32_csa1_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[9] = u_CSAwallace_pg_rca32_csa1_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[10] = u_CSAwallace_pg_rca32_csa1_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[11] = u_CSAwallace_pg_rca32_csa1_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[12] = u_CSAwallace_pg_rca32_csa1_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[13] = u_CSAwallace_pg_rca32_csa1_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[14] = u_CSAwallace_pg_rca32_csa1_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[15] = u_CSAwallace_pg_rca32_csa1_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[16] = u_CSAwallace_pg_rca32_csa1_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[17] = u_CSAwallace_pg_rca32_csa1_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[18] = u_CSAwallace_pg_rca32_csa1_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[19] = u_CSAwallace_pg_rca32_csa1_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[20] = u_CSAwallace_pg_rca32_csa1_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[21] = u_CSAwallace_pg_rca32_csa1_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[22] = u_CSAwallace_pg_rca32_csa1_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[23] = u_CSAwallace_pg_rca32_csa1_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[24] = u_CSAwallace_pg_rca32_csa1_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[25] = u_CSAwallace_pg_rca32_csa1_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[26] = u_CSAwallace_pg_rca32_csa1_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[27] = u_CSAwallace_pg_rca32_csa1_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[28] = u_CSAwallace_pg_rca32_csa1_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[29] = u_CSAwallace_pg_rca32_csa1_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[30] = u_CSAwallace_pg_rca32_csa1_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[31] = u_CSAwallace_pg_rca32_csa1_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[32] = u_CSAwallace_pg_rca32_csa1_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[33] = u_CSAwallace_pg_rca32_csa1_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[34] = u_CSAwallace_pg_rca32_csa1_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[35] = u_CSAwallace_pg_rca32_csa1_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[36] = u_CSAwallace_pg_rca32_csa1_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[37] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[38] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[39] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2[40] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[6] = u_CSAwallace_pg_rca32_csa2_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[7] = u_CSAwallace_pg_rca32_csa2_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[8] = u_CSAwallace_pg_rca32_csa2_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[9] = u_CSAwallace_pg_rca32_csa2_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[10] = u_CSAwallace_pg_rca32_csa2_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[11] = u_CSAwallace_pg_rca32_csa2_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[12] = u_CSAwallace_pg_rca32_csa2_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[13] = u_CSAwallace_pg_rca32_csa2_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[14] = u_CSAwallace_pg_rca32_csa2_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[15] = u_CSAwallace_pg_rca32_csa2_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[16] = u_CSAwallace_pg_rca32_csa2_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[17] = u_CSAwallace_pg_rca32_csa2_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[18] = u_CSAwallace_pg_rca32_csa2_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[19] = u_CSAwallace_pg_rca32_csa2_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[20] = u_CSAwallace_pg_rca32_csa2_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[21] = u_CSAwallace_pg_rca32_csa2_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[22] = u_CSAwallace_pg_rca32_csa2_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[23] = u_CSAwallace_pg_rca32_csa2_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[24] = u_CSAwallace_pg_rca32_csa2_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[25] = u_CSAwallace_pg_rca32_csa2_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[26] = u_CSAwallace_pg_rca32_csa2_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[27] = u_CSAwallace_pg_rca32_csa2_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[28] = u_CSAwallace_pg_rca32_csa2_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[29] = u_CSAwallace_pg_rca32_csa2_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[30] = u_CSAwallace_pg_rca32_csa2_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[31] = u_CSAwallace_pg_rca32_csa2_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[32] = u_CSAwallace_pg_rca32_csa2_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[33] = u_CSAwallace_pg_rca32_csa2_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[34] = u_CSAwallace_pg_rca32_csa2_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[35] = u_CSAwallace_pg_rca32_csa2_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[36] = u_CSAwallace_pg_rca32_csa2_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[37] = u_CSAwallace_pg_rca32_csa2_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[38] = u_CSAwallace_pg_rca32_csa2_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[39] = u_CSAwallace_pg_rca32_csa2_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3[40] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[8] = u_CSAwallace_pg_rca32_csa2_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[9] = u_CSAwallace_pg_rca32_csa2_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[10] = u_CSAwallace_pg_rca32_csa2_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[11] = u_CSAwallace_pg_rca32_csa2_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[12] = u_CSAwallace_pg_rca32_csa2_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[13] = u_CSAwallace_pg_rca32_csa2_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[14] = u_CSAwallace_pg_rca32_csa2_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[15] = u_CSAwallace_pg_rca32_csa2_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[16] = u_CSAwallace_pg_rca32_csa2_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[17] = u_CSAwallace_pg_rca32_csa2_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[18] = u_CSAwallace_pg_rca32_csa2_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[19] = u_CSAwallace_pg_rca32_csa2_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[20] = u_CSAwallace_pg_rca32_csa2_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[21] = u_CSAwallace_pg_rca32_csa2_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[22] = u_CSAwallace_pg_rca32_csa2_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[23] = u_CSAwallace_pg_rca32_csa2_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[24] = u_CSAwallace_pg_rca32_csa2_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[25] = u_CSAwallace_pg_rca32_csa2_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[26] = u_CSAwallace_pg_rca32_csa2_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[27] = u_CSAwallace_pg_rca32_csa2_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[28] = u_CSAwallace_pg_rca32_csa2_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[29] = u_CSAwallace_pg_rca32_csa2_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[30] = u_CSAwallace_pg_rca32_csa2_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[31] = u_CSAwallace_pg_rca32_csa2_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[32] = u_CSAwallace_pg_rca32_csa2_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[33] = u_CSAwallace_pg_rca32_csa2_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[34] = u_CSAwallace_pg_rca32_csa2_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[35] = u_CSAwallace_pg_rca32_csa2_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[36] = u_CSAwallace_pg_rca32_csa2_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[37] = u_CSAwallace_pg_rca32_csa2_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[38] = u_CSAwallace_pg_rca32_csa2_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[39] = u_CSAwallace_pg_rca32_csa2_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3[40] = 1'b0;
  csa_component41 csa_component41_u_CSAwallace_pg_rca32_csa11_csa_component_out(.a(u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c2), .b(u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_s3), .c(u_CSAwallace_pg_rca32_csa11_csa_component_u_CSAwallace_pg_rca32_csa_c3), .csa_component41_out(u_CSAwallace_pg_rca32_csa11_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[9] = u_CSAwallace_pg_rca32_csa3_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[10] = u_CSAwallace_pg_rca32_csa3_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[11] = u_CSAwallace_pg_rca32_csa3_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[12] = u_CSAwallace_pg_rca32_csa3_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[13] = u_CSAwallace_pg_rca32_csa3_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[14] = u_CSAwallace_pg_rca32_csa3_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[15] = u_CSAwallace_pg_rca32_csa3_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[16] = u_CSAwallace_pg_rca32_csa3_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[17] = u_CSAwallace_pg_rca32_csa3_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[18] = u_CSAwallace_pg_rca32_csa3_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[19] = u_CSAwallace_pg_rca32_csa3_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[20] = u_CSAwallace_pg_rca32_csa3_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[21] = u_CSAwallace_pg_rca32_csa3_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[22] = u_CSAwallace_pg_rca32_csa3_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[23] = u_CSAwallace_pg_rca32_csa3_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[24] = u_CSAwallace_pg_rca32_csa3_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[25] = u_CSAwallace_pg_rca32_csa3_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[26] = u_CSAwallace_pg_rca32_csa3_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[27] = u_CSAwallace_pg_rca32_csa3_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[28] = u_CSAwallace_pg_rca32_csa3_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[29] = u_CSAwallace_pg_rca32_csa3_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[30] = u_CSAwallace_pg_rca32_csa3_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[31] = u_CSAwallace_pg_rca32_csa3_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[32] = u_CSAwallace_pg_rca32_csa3_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[33] = u_CSAwallace_pg_rca32_csa3_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[34] = u_CSAwallace_pg_rca32_csa3_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[35] = u_CSAwallace_pg_rca32_csa3_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[36] = u_CSAwallace_pg_rca32_csa3_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[37] = u_CSAwallace_pg_rca32_csa3_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[38] = u_CSAwallace_pg_rca32_csa3_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[39] = u_CSAwallace_pg_rca32_csa3_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[40] = u_CSAwallace_pg_rca32_csa3_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[41] = u_CSAwallace_pg_rca32_csa3_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[42] = u_CSAwallace_pg_rca32_csa3_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[43] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[44] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[11] = u_CSAwallace_pg_rca32_csa3_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[12] = u_CSAwallace_pg_rca32_csa3_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[13] = u_CSAwallace_pg_rca32_csa3_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[14] = u_CSAwallace_pg_rca32_csa3_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[15] = u_CSAwallace_pg_rca32_csa3_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[16] = u_CSAwallace_pg_rca32_csa3_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[17] = u_CSAwallace_pg_rca32_csa3_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[18] = u_CSAwallace_pg_rca32_csa3_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[19] = u_CSAwallace_pg_rca32_csa3_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[20] = u_CSAwallace_pg_rca32_csa3_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[21] = u_CSAwallace_pg_rca32_csa3_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[22] = u_CSAwallace_pg_rca32_csa3_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[23] = u_CSAwallace_pg_rca32_csa3_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[24] = u_CSAwallace_pg_rca32_csa3_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[25] = u_CSAwallace_pg_rca32_csa3_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[26] = u_CSAwallace_pg_rca32_csa3_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[27] = u_CSAwallace_pg_rca32_csa3_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[28] = u_CSAwallace_pg_rca32_csa3_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[29] = u_CSAwallace_pg_rca32_csa3_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[30] = u_CSAwallace_pg_rca32_csa3_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[31] = u_CSAwallace_pg_rca32_csa3_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[32] = u_CSAwallace_pg_rca32_csa3_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[33] = u_CSAwallace_pg_rca32_csa3_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[34] = u_CSAwallace_pg_rca32_csa3_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[35] = u_CSAwallace_pg_rca32_csa3_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[36] = u_CSAwallace_pg_rca32_csa3_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[37] = u_CSAwallace_pg_rca32_csa3_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[38] = u_CSAwallace_pg_rca32_csa3_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[39] = u_CSAwallace_pg_rca32_csa3_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[40] = u_CSAwallace_pg_rca32_csa3_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[41] = u_CSAwallace_pg_rca32_csa3_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[42] = u_CSAwallace_pg_rca32_csa3_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[43] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[44] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[12] = u_CSAwallace_pg_rca32_csa4_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[13] = u_CSAwallace_pg_rca32_csa4_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[14] = u_CSAwallace_pg_rca32_csa4_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[15] = u_CSAwallace_pg_rca32_csa4_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[16] = u_CSAwallace_pg_rca32_csa4_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[17] = u_CSAwallace_pg_rca32_csa4_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[18] = u_CSAwallace_pg_rca32_csa4_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[19] = u_CSAwallace_pg_rca32_csa4_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[20] = u_CSAwallace_pg_rca32_csa4_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[21] = u_CSAwallace_pg_rca32_csa4_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[22] = u_CSAwallace_pg_rca32_csa4_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[23] = u_CSAwallace_pg_rca32_csa4_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[24] = u_CSAwallace_pg_rca32_csa4_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[25] = u_CSAwallace_pg_rca32_csa4_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[26] = u_CSAwallace_pg_rca32_csa4_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[27] = u_CSAwallace_pg_rca32_csa4_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[28] = u_CSAwallace_pg_rca32_csa4_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[29] = u_CSAwallace_pg_rca32_csa4_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[30] = u_CSAwallace_pg_rca32_csa4_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[31] = u_CSAwallace_pg_rca32_csa4_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[32] = u_CSAwallace_pg_rca32_csa4_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[33] = u_CSAwallace_pg_rca32_csa4_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[34] = u_CSAwallace_pg_rca32_csa4_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[35] = u_CSAwallace_pg_rca32_csa4_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[36] = u_CSAwallace_pg_rca32_csa4_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[37] = u_CSAwallace_pg_rca32_csa4_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[38] = u_CSAwallace_pg_rca32_csa4_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[39] = u_CSAwallace_pg_rca32_csa4_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[40] = u_CSAwallace_pg_rca32_csa4_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[41] = u_CSAwallace_pg_rca32_csa4_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[42] = u_CSAwallace_pg_rca32_csa4_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[43] = u_CSAwallace_pg_rca32_csa4_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[44] = u_CSAwallace_pg_rca32_csa4_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[45] = u_CSAwallace_pg_rca32_csa4_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5[46] = 1'b0;
  csa_component47 csa_component47_u_CSAwallace_pg_rca32_csa12_csa_component_out(.a(u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s4), .b(u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_c4), .c(u_CSAwallace_pg_rca32_csa12_csa_component_u_CSAwallace_pg_rca32_csa_s5), .csa_component47_out(u_CSAwallace_pg_rca32_csa12_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[14] = u_CSAwallace_pg_rca32_csa4_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[15] = u_CSAwallace_pg_rca32_csa4_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[16] = u_CSAwallace_pg_rca32_csa4_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[17] = u_CSAwallace_pg_rca32_csa4_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[18] = u_CSAwallace_pg_rca32_csa4_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[19] = u_CSAwallace_pg_rca32_csa4_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[20] = u_CSAwallace_pg_rca32_csa4_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[21] = u_CSAwallace_pg_rca32_csa4_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[22] = u_CSAwallace_pg_rca32_csa4_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[23] = u_CSAwallace_pg_rca32_csa4_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[24] = u_CSAwallace_pg_rca32_csa4_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[25] = u_CSAwallace_pg_rca32_csa4_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[26] = u_CSAwallace_pg_rca32_csa4_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[27] = u_CSAwallace_pg_rca32_csa4_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[28] = u_CSAwallace_pg_rca32_csa4_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[29] = u_CSAwallace_pg_rca32_csa4_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[30] = u_CSAwallace_pg_rca32_csa4_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[31] = u_CSAwallace_pg_rca32_csa4_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[32] = u_CSAwallace_pg_rca32_csa4_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[33] = u_CSAwallace_pg_rca32_csa4_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[34] = u_CSAwallace_pg_rca32_csa4_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[35] = u_CSAwallace_pg_rca32_csa4_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[36] = u_CSAwallace_pg_rca32_csa4_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[37] = u_CSAwallace_pg_rca32_csa4_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[38] = u_CSAwallace_pg_rca32_csa4_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[39] = u_CSAwallace_pg_rca32_csa4_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[40] = u_CSAwallace_pg_rca32_csa4_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[41] = u_CSAwallace_pg_rca32_csa4_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[42] = u_CSAwallace_pg_rca32_csa4_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[43] = u_CSAwallace_pg_rca32_csa4_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[44] = u_CSAwallace_pg_rca32_csa4_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[45] = u_CSAwallace_pg_rca32_csa4_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5[49] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[15] = u_CSAwallace_pg_rca32_csa5_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[16] = u_CSAwallace_pg_rca32_csa5_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[17] = u_CSAwallace_pg_rca32_csa5_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[18] = u_CSAwallace_pg_rca32_csa5_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[19] = u_CSAwallace_pg_rca32_csa5_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[20] = u_CSAwallace_pg_rca32_csa5_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[21] = u_CSAwallace_pg_rca32_csa5_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[22] = u_CSAwallace_pg_rca32_csa5_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[23] = u_CSAwallace_pg_rca32_csa5_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[24] = u_CSAwallace_pg_rca32_csa5_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[25] = u_CSAwallace_pg_rca32_csa5_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[26] = u_CSAwallace_pg_rca32_csa5_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[27] = u_CSAwallace_pg_rca32_csa5_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[28] = u_CSAwallace_pg_rca32_csa5_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[29] = u_CSAwallace_pg_rca32_csa5_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[30] = u_CSAwallace_pg_rca32_csa5_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[31] = u_CSAwallace_pg_rca32_csa5_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[32] = u_CSAwallace_pg_rca32_csa5_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[33] = u_CSAwallace_pg_rca32_csa5_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[34] = u_CSAwallace_pg_rca32_csa5_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[35] = u_CSAwallace_pg_rca32_csa5_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[36] = u_CSAwallace_pg_rca32_csa5_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[37] = u_CSAwallace_pg_rca32_csa5_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[38] = u_CSAwallace_pg_rca32_csa5_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[39] = u_CSAwallace_pg_rca32_csa5_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[40] = u_CSAwallace_pg_rca32_csa5_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[41] = u_CSAwallace_pg_rca32_csa5_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[42] = u_CSAwallace_pg_rca32_csa5_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[43] = u_CSAwallace_pg_rca32_csa5_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[44] = u_CSAwallace_pg_rca32_csa5_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[45] = u_CSAwallace_pg_rca32_csa5_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[46] = u_CSAwallace_pg_rca32_csa5_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[47] = u_CSAwallace_pg_rca32_csa5_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[48] = u_CSAwallace_pg_rca32_csa5_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6[49] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[17] = u_CSAwallace_pg_rca32_csa5_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[18] = u_CSAwallace_pg_rca32_csa5_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[19] = u_CSAwallace_pg_rca32_csa5_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[20] = u_CSAwallace_pg_rca32_csa5_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[21] = u_CSAwallace_pg_rca32_csa5_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[22] = u_CSAwallace_pg_rca32_csa5_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[23] = u_CSAwallace_pg_rca32_csa5_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[24] = u_CSAwallace_pg_rca32_csa5_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[25] = u_CSAwallace_pg_rca32_csa5_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[26] = u_CSAwallace_pg_rca32_csa5_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[27] = u_CSAwallace_pg_rca32_csa5_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[28] = u_CSAwallace_pg_rca32_csa5_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[29] = u_CSAwallace_pg_rca32_csa5_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[30] = u_CSAwallace_pg_rca32_csa5_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[31] = u_CSAwallace_pg_rca32_csa5_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[32] = u_CSAwallace_pg_rca32_csa5_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[33] = u_CSAwallace_pg_rca32_csa5_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[34] = u_CSAwallace_pg_rca32_csa5_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[35] = u_CSAwallace_pg_rca32_csa5_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[36] = u_CSAwallace_pg_rca32_csa5_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[37] = u_CSAwallace_pg_rca32_csa5_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[38] = u_CSAwallace_pg_rca32_csa5_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[39] = u_CSAwallace_pg_rca32_csa5_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[40] = u_CSAwallace_pg_rca32_csa5_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[41] = u_CSAwallace_pg_rca32_csa5_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[42] = u_CSAwallace_pg_rca32_csa5_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[43] = u_CSAwallace_pg_rca32_csa5_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[44] = u_CSAwallace_pg_rca32_csa5_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[45] = u_CSAwallace_pg_rca32_csa5_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[46] = u_CSAwallace_pg_rca32_csa5_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[47] = u_CSAwallace_pg_rca32_csa5_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[48] = u_CSAwallace_pg_rca32_csa5_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6[49] = 1'b0;
  csa_component50 csa_component50_u_CSAwallace_pg_rca32_csa13_csa_component_out(.a(u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c5), .b(u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_s6), .c(u_CSAwallace_pg_rca32_csa13_csa_component_u_CSAwallace_pg_rca32_csa_c6), .csa_component50_out(u_CSAwallace_pg_rca32_csa13_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[18] = u_CSAwallace_pg_rca32_csa6_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[19] = u_CSAwallace_pg_rca32_csa6_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[20] = u_CSAwallace_pg_rca32_csa6_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[21] = u_CSAwallace_pg_rca32_csa6_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[22] = u_CSAwallace_pg_rca32_csa6_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[23] = u_CSAwallace_pg_rca32_csa6_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[24] = u_CSAwallace_pg_rca32_csa6_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[25] = u_CSAwallace_pg_rca32_csa6_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[26] = u_CSAwallace_pg_rca32_csa6_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[27] = u_CSAwallace_pg_rca32_csa6_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[28] = u_CSAwallace_pg_rca32_csa6_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[29] = u_CSAwallace_pg_rca32_csa6_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[30] = u_CSAwallace_pg_rca32_csa6_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[31] = u_CSAwallace_pg_rca32_csa6_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[32] = u_CSAwallace_pg_rca32_csa6_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[33] = u_CSAwallace_pg_rca32_csa6_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[34] = u_CSAwallace_pg_rca32_csa6_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[35] = u_CSAwallace_pg_rca32_csa6_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[36] = u_CSAwallace_pg_rca32_csa6_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[37] = u_CSAwallace_pg_rca32_csa6_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[38] = u_CSAwallace_pg_rca32_csa6_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[39] = u_CSAwallace_pg_rca32_csa6_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[40] = u_CSAwallace_pg_rca32_csa6_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[41] = u_CSAwallace_pg_rca32_csa6_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[42] = u_CSAwallace_pg_rca32_csa6_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[43] = u_CSAwallace_pg_rca32_csa6_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[44] = u_CSAwallace_pg_rca32_csa6_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[45] = u_CSAwallace_pg_rca32_csa6_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[46] = u_CSAwallace_pg_rca32_csa6_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[47] = u_CSAwallace_pg_rca32_csa6_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[48] = u_CSAwallace_pg_rca32_csa6_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[49] = u_CSAwallace_pg_rca32_csa6_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[50] = u_CSAwallace_pg_rca32_csa6_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[51] = u_CSAwallace_pg_rca32_csa6_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[20] = u_CSAwallace_pg_rca32_csa6_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[21] = u_CSAwallace_pg_rca32_csa6_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[22] = u_CSAwallace_pg_rca32_csa6_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[23] = u_CSAwallace_pg_rca32_csa6_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[24] = u_CSAwallace_pg_rca32_csa6_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[25] = u_CSAwallace_pg_rca32_csa6_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[26] = u_CSAwallace_pg_rca32_csa6_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[27] = u_CSAwallace_pg_rca32_csa6_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[28] = u_CSAwallace_pg_rca32_csa6_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[29] = u_CSAwallace_pg_rca32_csa6_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[30] = u_CSAwallace_pg_rca32_csa6_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[31] = u_CSAwallace_pg_rca32_csa6_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[32] = u_CSAwallace_pg_rca32_csa6_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[33] = u_CSAwallace_pg_rca32_csa6_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[34] = u_CSAwallace_pg_rca32_csa6_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[35] = u_CSAwallace_pg_rca32_csa6_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[36] = u_CSAwallace_pg_rca32_csa6_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[37] = u_CSAwallace_pg_rca32_csa6_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[38] = u_CSAwallace_pg_rca32_csa6_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[39] = u_CSAwallace_pg_rca32_csa6_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[40] = u_CSAwallace_pg_rca32_csa6_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[41] = u_CSAwallace_pg_rca32_csa6_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[42] = u_CSAwallace_pg_rca32_csa6_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[43] = u_CSAwallace_pg_rca32_csa6_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[44] = u_CSAwallace_pg_rca32_csa6_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[45] = u_CSAwallace_pg_rca32_csa6_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[46] = u_CSAwallace_pg_rca32_csa6_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[47] = u_CSAwallace_pg_rca32_csa6_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[48] = u_CSAwallace_pg_rca32_csa6_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[49] = u_CSAwallace_pg_rca32_csa6_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[50] = u_CSAwallace_pg_rca32_csa6_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[51] = u_CSAwallace_pg_rca32_csa6_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[21] = u_CSAwallace_pg_rca32_csa7_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[22] = u_CSAwallace_pg_rca32_csa7_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[23] = u_CSAwallace_pg_rca32_csa7_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[24] = u_CSAwallace_pg_rca32_csa7_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[25] = u_CSAwallace_pg_rca32_csa7_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[26] = u_CSAwallace_pg_rca32_csa7_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[27] = u_CSAwallace_pg_rca32_csa7_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[28] = u_CSAwallace_pg_rca32_csa7_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[29] = u_CSAwallace_pg_rca32_csa7_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[30] = u_CSAwallace_pg_rca32_csa7_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[31] = u_CSAwallace_pg_rca32_csa7_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[32] = u_CSAwallace_pg_rca32_csa7_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[33] = u_CSAwallace_pg_rca32_csa7_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[34] = u_CSAwallace_pg_rca32_csa7_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[35] = u_CSAwallace_pg_rca32_csa7_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[36] = u_CSAwallace_pg_rca32_csa7_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[37] = u_CSAwallace_pg_rca32_csa7_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[38] = u_CSAwallace_pg_rca32_csa7_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[39] = u_CSAwallace_pg_rca32_csa7_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[40] = u_CSAwallace_pg_rca32_csa7_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[41] = u_CSAwallace_pg_rca32_csa7_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[42] = u_CSAwallace_pg_rca32_csa7_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[43] = u_CSAwallace_pg_rca32_csa7_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[44] = u_CSAwallace_pg_rca32_csa7_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[45] = u_CSAwallace_pg_rca32_csa7_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[46] = u_CSAwallace_pg_rca32_csa7_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[47] = u_CSAwallace_pg_rca32_csa7_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[48] = u_CSAwallace_pg_rca32_csa7_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[49] = u_CSAwallace_pg_rca32_csa7_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[50] = u_CSAwallace_pg_rca32_csa7_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[51] = u_CSAwallace_pg_rca32_csa7_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[52] = u_CSAwallace_pg_rca32_csa7_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[53] = u_CSAwallace_pg_rca32_csa7_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[54] = u_CSAwallace_pg_rca32_csa7_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8[55] = 1'b0;
  csa_component56 csa_component56_u_CSAwallace_pg_rca32_csa14_csa_component_out(.a(u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s7), .b(u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_c7), .c(u_CSAwallace_pg_rca32_csa14_csa_component_u_CSAwallace_pg_rca32_csa_s8), .csa_component56_out(u_CSAwallace_pg_rca32_csa14_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[23] = u_CSAwallace_pg_rca32_csa7_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[24] = u_CSAwallace_pg_rca32_csa7_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[25] = u_CSAwallace_pg_rca32_csa7_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[26] = u_CSAwallace_pg_rca32_csa7_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[27] = u_CSAwallace_pg_rca32_csa7_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[28] = u_CSAwallace_pg_rca32_csa7_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[29] = u_CSAwallace_pg_rca32_csa7_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[30] = u_CSAwallace_pg_rca32_csa7_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[31] = u_CSAwallace_pg_rca32_csa7_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[32] = u_CSAwallace_pg_rca32_csa7_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[33] = u_CSAwallace_pg_rca32_csa7_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[34] = u_CSAwallace_pg_rca32_csa7_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[35] = u_CSAwallace_pg_rca32_csa7_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[36] = u_CSAwallace_pg_rca32_csa7_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[37] = u_CSAwallace_pg_rca32_csa7_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[38] = u_CSAwallace_pg_rca32_csa7_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[39] = u_CSAwallace_pg_rca32_csa7_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[40] = u_CSAwallace_pg_rca32_csa7_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[41] = u_CSAwallace_pg_rca32_csa7_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[42] = u_CSAwallace_pg_rca32_csa7_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[43] = u_CSAwallace_pg_rca32_csa7_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[44] = u_CSAwallace_pg_rca32_csa7_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[45] = u_CSAwallace_pg_rca32_csa7_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[46] = u_CSAwallace_pg_rca32_csa7_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[47] = u_CSAwallace_pg_rca32_csa7_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[48] = u_CSAwallace_pg_rca32_csa7_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[49] = u_CSAwallace_pg_rca32_csa7_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[50] = u_CSAwallace_pg_rca32_csa7_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[51] = u_CSAwallace_pg_rca32_csa7_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[52] = u_CSAwallace_pg_rca32_csa7_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[53] = u_CSAwallace_pg_rca32_csa7_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[54] = u_CSAwallace_pg_rca32_csa7_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[24] = u_CSAwallace_pg_rca32_csa8_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[25] = u_CSAwallace_pg_rca32_csa8_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[26] = u_CSAwallace_pg_rca32_csa8_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[27] = u_CSAwallace_pg_rca32_csa8_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[28] = u_CSAwallace_pg_rca32_csa8_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[29] = u_CSAwallace_pg_rca32_csa8_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[30] = u_CSAwallace_pg_rca32_csa8_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[31] = u_CSAwallace_pg_rca32_csa8_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[32] = u_CSAwallace_pg_rca32_csa8_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[33] = u_CSAwallace_pg_rca32_csa8_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[34] = u_CSAwallace_pg_rca32_csa8_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[35] = u_CSAwallace_pg_rca32_csa8_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[36] = u_CSAwallace_pg_rca32_csa8_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[37] = u_CSAwallace_pg_rca32_csa8_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[38] = u_CSAwallace_pg_rca32_csa8_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[39] = u_CSAwallace_pg_rca32_csa8_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[40] = u_CSAwallace_pg_rca32_csa8_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[41] = u_CSAwallace_pg_rca32_csa8_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[42] = u_CSAwallace_pg_rca32_csa8_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[43] = u_CSAwallace_pg_rca32_csa8_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[44] = u_CSAwallace_pg_rca32_csa8_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[45] = u_CSAwallace_pg_rca32_csa8_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[46] = u_CSAwallace_pg_rca32_csa8_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[47] = u_CSAwallace_pg_rca32_csa8_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[48] = u_CSAwallace_pg_rca32_csa8_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[49] = u_CSAwallace_pg_rca32_csa8_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[50] = u_CSAwallace_pg_rca32_csa8_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[51] = u_CSAwallace_pg_rca32_csa8_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[52] = u_CSAwallace_pg_rca32_csa8_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[53] = u_CSAwallace_pg_rca32_csa8_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[54] = u_CSAwallace_pg_rca32_csa8_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[55] = u_CSAwallace_pg_rca32_csa8_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[56] = u_CSAwallace_pg_rca32_csa8_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[57] = u_CSAwallace_pg_rca32_csa8_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[26] = u_CSAwallace_pg_rca32_csa8_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[27] = u_CSAwallace_pg_rca32_csa8_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[28] = u_CSAwallace_pg_rca32_csa8_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[29] = u_CSAwallace_pg_rca32_csa8_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[30] = u_CSAwallace_pg_rca32_csa8_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[31] = u_CSAwallace_pg_rca32_csa8_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[32] = u_CSAwallace_pg_rca32_csa8_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[33] = u_CSAwallace_pg_rca32_csa8_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[34] = u_CSAwallace_pg_rca32_csa8_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[35] = u_CSAwallace_pg_rca32_csa8_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[36] = u_CSAwallace_pg_rca32_csa8_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[37] = u_CSAwallace_pg_rca32_csa8_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[38] = u_CSAwallace_pg_rca32_csa8_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[39] = u_CSAwallace_pg_rca32_csa8_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[40] = u_CSAwallace_pg_rca32_csa8_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[41] = u_CSAwallace_pg_rca32_csa8_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[42] = u_CSAwallace_pg_rca32_csa8_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[43] = u_CSAwallace_pg_rca32_csa8_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[44] = u_CSAwallace_pg_rca32_csa8_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[45] = u_CSAwallace_pg_rca32_csa8_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[46] = u_CSAwallace_pg_rca32_csa8_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[47] = u_CSAwallace_pg_rca32_csa8_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[48] = u_CSAwallace_pg_rca32_csa8_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[49] = u_CSAwallace_pg_rca32_csa8_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[50] = u_CSAwallace_pg_rca32_csa8_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[51] = u_CSAwallace_pg_rca32_csa8_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[52] = u_CSAwallace_pg_rca32_csa8_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[53] = u_CSAwallace_pg_rca32_csa8_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[54] = u_CSAwallace_pg_rca32_csa8_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[55] = u_CSAwallace_pg_rca32_csa8_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[56] = u_CSAwallace_pg_rca32_csa8_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[57] = u_CSAwallace_pg_rca32_csa8_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9[58] = 1'b0;
  csa_component59 csa_component59_u_CSAwallace_pg_rca32_csa15_csa_component_out(.a(u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c8), .b(u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_s9), .c(u_CSAwallace_pg_rca32_csa15_csa_component_u_CSAwallace_pg_rca32_csa_c9), .csa_component59_out(u_CSAwallace_pg_rca32_csa15_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[27] = u_CSAwallace_pg_rca32_csa9_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[28] = u_CSAwallace_pg_rca32_csa9_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[29] = u_CSAwallace_pg_rca32_csa9_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[30] = u_CSAwallace_pg_rca32_csa9_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[31] = u_CSAwallace_pg_rca32_csa9_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[32] = u_CSAwallace_pg_rca32_csa9_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[33] = u_CSAwallace_pg_rca32_csa9_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[34] = u_CSAwallace_pg_rca32_csa9_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[35] = u_CSAwallace_pg_rca32_csa9_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[36] = u_CSAwallace_pg_rca32_csa9_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[37] = u_CSAwallace_pg_rca32_csa9_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[38] = u_CSAwallace_pg_rca32_csa9_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[39] = u_CSAwallace_pg_rca32_csa9_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[40] = u_CSAwallace_pg_rca32_csa9_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[41] = u_CSAwallace_pg_rca32_csa9_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[42] = u_CSAwallace_pg_rca32_csa9_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[43] = u_CSAwallace_pg_rca32_csa9_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[44] = u_CSAwallace_pg_rca32_csa9_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[45] = u_CSAwallace_pg_rca32_csa9_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[46] = u_CSAwallace_pg_rca32_csa9_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[47] = u_CSAwallace_pg_rca32_csa9_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[48] = u_CSAwallace_pg_rca32_csa9_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[49] = u_CSAwallace_pg_rca32_csa9_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[50] = u_CSAwallace_pg_rca32_csa9_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[51] = u_CSAwallace_pg_rca32_csa9_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[52] = u_CSAwallace_pg_rca32_csa9_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[53] = u_CSAwallace_pg_rca32_csa9_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[54] = u_CSAwallace_pg_rca32_csa9_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[55] = u_CSAwallace_pg_rca32_csa9_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[56] = u_CSAwallace_pg_rca32_csa9_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[57] = u_CSAwallace_pg_rca32_csa9_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[58] = u_CSAwallace_pg_rca32_csa9_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[59] = u_CSAwallace_pg_rca32_csa9_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[60] = u_CSAwallace_pg_rca32_csa9_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[27] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[28] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[29] = u_CSAwallace_pg_rca32_csa9_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[30] = u_CSAwallace_pg_rca32_csa9_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[31] = u_CSAwallace_pg_rca32_csa9_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[32] = u_CSAwallace_pg_rca32_csa9_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[33] = u_CSAwallace_pg_rca32_csa9_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[34] = u_CSAwallace_pg_rca32_csa9_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[35] = u_CSAwallace_pg_rca32_csa9_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[36] = u_CSAwallace_pg_rca32_csa9_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[37] = u_CSAwallace_pg_rca32_csa9_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[38] = u_CSAwallace_pg_rca32_csa9_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[39] = u_CSAwallace_pg_rca32_csa9_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[40] = u_CSAwallace_pg_rca32_csa9_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[41] = u_CSAwallace_pg_rca32_csa9_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[42] = u_CSAwallace_pg_rca32_csa9_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[43] = u_CSAwallace_pg_rca32_csa9_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[44] = u_CSAwallace_pg_rca32_csa9_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[45] = u_CSAwallace_pg_rca32_csa9_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[46] = u_CSAwallace_pg_rca32_csa9_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[47] = u_CSAwallace_pg_rca32_csa9_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[48] = u_CSAwallace_pg_rca32_csa9_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[49] = u_CSAwallace_pg_rca32_csa9_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[50] = u_CSAwallace_pg_rca32_csa9_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[51] = u_CSAwallace_pg_rca32_csa9_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[52] = u_CSAwallace_pg_rca32_csa9_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[53] = u_CSAwallace_pg_rca32_csa9_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[54] = u_CSAwallace_pg_rca32_csa9_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[55] = u_CSAwallace_pg_rca32_csa9_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[56] = u_CSAwallace_pg_rca32_csa9_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[57] = u_CSAwallace_pg_rca32_csa9_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[58] = u_CSAwallace_pg_rca32_csa9_csa_component_out[120];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[59] = u_CSAwallace_pg_rca32_csa9_csa_component_out[121];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[60] = u_CSAwallace_pg_rca32_csa9_csa_component_out[122];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[27] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[28] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[29] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[30] = u_CSAwallace_pg_rca32_and_0_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[31] = u_CSAwallace_pg_rca32_and_1_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[32] = u_CSAwallace_pg_rca32_and_2_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[33] = u_CSAwallace_pg_rca32_and_3_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[34] = u_CSAwallace_pg_rca32_and_4_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[35] = u_CSAwallace_pg_rca32_and_5_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[36] = u_CSAwallace_pg_rca32_and_6_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[37] = u_CSAwallace_pg_rca32_and_7_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[38] = u_CSAwallace_pg_rca32_and_8_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[39] = u_CSAwallace_pg_rca32_and_9_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[40] = u_CSAwallace_pg_rca32_and_10_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[41] = u_CSAwallace_pg_rca32_and_11_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[42] = u_CSAwallace_pg_rca32_and_12_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[43] = u_CSAwallace_pg_rca32_and_13_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[44] = u_CSAwallace_pg_rca32_and_14_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[45] = u_CSAwallace_pg_rca32_and_15_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[46] = u_CSAwallace_pg_rca32_and_16_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[47] = u_CSAwallace_pg_rca32_and_17_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[48] = u_CSAwallace_pg_rca32_and_18_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[49] = u_CSAwallace_pg_rca32_and_19_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[50] = u_CSAwallace_pg_rca32_and_20_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[51] = u_CSAwallace_pg_rca32_and_21_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[52] = u_CSAwallace_pg_rca32_and_22_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[53] = u_CSAwallace_pg_rca32_and_23_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[54] = u_CSAwallace_pg_rca32_and_24_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[55] = u_CSAwallace_pg_rca32_and_25_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[56] = u_CSAwallace_pg_rca32_and_26_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[57] = u_CSAwallace_pg_rca32_and_27_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[58] = u_CSAwallace_pg_rca32_and_28_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[59] = u_CSAwallace_pg_rca32_and_29_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[60] = u_CSAwallace_pg_rca32_and_30_30[0];
  assign u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30[61] = u_CSAwallace_pg_rca32_and_31_30[0];
  csa_component62 csa_component62_u_CSAwallace_pg_rca32_csa16_csa_component_out(.a(u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_s10), .b(u_CSAwallace_pg_rca32_csa16_csa_component_u_CSAwallace_pg_rca32_csa_c10), .c(u_CSAwallace_pg_rca32_csa16_csa_component_pp_row30), .csa_component62_out(u_CSAwallace_pg_rca32_csa16_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[0] = u_CSAwallace_pg_rca32_csa10_csa_component_out[0];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[1] = u_CSAwallace_pg_rca32_csa10_csa_component_out[1];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[2] = u_CSAwallace_pg_rca32_csa10_csa_component_out[2];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[3] = u_CSAwallace_pg_rca32_csa10_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[4] = u_CSAwallace_pg_rca32_csa10_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[5] = u_CSAwallace_pg_rca32_csa10_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[6] = u_CSAwallace_pg_rca32_csa10_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[7] = u_CSAwallace_pg_rca32_csa10_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[8] = u_CSAwallace_pg_rca32_csa10_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[9] = u_CSAwallace_pg_rca32_csa10_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[10] = u_CSAwallace_pg_rca32_csa10_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[11] = u_CSAwallace_pg_rca32_csa10_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[12] = u_CSAwallace_pg_rca32_csa10_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[13] = u_CSAwallace_pg_rca32_csa10_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[14] = u_CSAwallace_pg_rca32_csa10_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[15] = u_CSAwallace_pg_rca32_csa10_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[16] = u_CSAwallace_pg_rca32_csa10_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[17] = u_CSAwallace_pg_rca32_csa10_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[18] = u_CSAwallace_pg_rca32_csa10_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[19] = u_CSAwallace_pg_rca32_csa10_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[20] = u_CSAwallace_pg_rca32_csa10_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[21] = u_CSAwallace_pg_rca32_csa10_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[22] = u_CSAwallace_pg_rca32_csa10_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[23] = u_CSAwallace_pg_rca32_csa10_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[24] = u_CSAwallace_pg_rca32_csa10_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[25] = u_CSAwallace_pg_rca32_csa10_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[26] = u_CSAwallace_pg_rca32_csa10_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[27] = u_CSAwallace_pg_rca32_csa10_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[28] = u_CSAwallace_pg_rca32_csa10_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[29] = u_CSAwallace_pg_rca32_csa10_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[30] = u_CSAwallace_pg_rca32_csa10_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[31] = u_CSAwallace_pg_rca32_csa10_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[32] = u_CSAwallace_pg_rca32_csa10_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[33] = u_CSAwallace_pg_rca32_csa10_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[34] = u_CSAwallace_pg_rca32_csa10_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[35] = u_CSAwallace_pg_rca32_csa10_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[36] = u_CSAwallace_pg_rca32_csa10_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[37] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[38] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[39] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[40] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11[41] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[3] = u_CSAwallace_pg_rca32_csa10_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[4] = u_CSAwallace_pg_rca32_csa10_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[5] = u_CSAwallace_pg_rca32_csa10_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[6] = u_CSAwallace_pg_rca32_csa10_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[7] = u_CSAwallace_pg_rca32_csa10_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[8] = u_CSAwallace_pg_rca32_csa10_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[9] = u_CSAwallace_pg_rca32_csa10_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[10] = u_CSAwallace_pg_rca32_csa10_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[11] = u_CSAwallace_pg_rca32_csa10_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[12] = u_CSAwallace_pg_rca32_csa10_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[13] = u_CSAwallace_pg_rca32_csa10_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[14] = u_CSAwallace_pg_rca32_csa10_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[15] = u_CSAwallace_pg_rca32_csa10_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[16] = u_CSAwallace_pg_rca32_csa10_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[17] = u_CSAwallace_pg_rca32_csa10_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[18] = u_CSAwallace_pg_rca32_csa10_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[19] = u_CSAwallace_pg_rca32_csa10_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[20] = u_CSAwallace_pg_rca32_csa10_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[21] = u_CSAwallace_pg_rca32_csa10_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[22] = u_CSAwallace_pg_rca32_csa10_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[23] = u_CSAwallace_pg_rca32_csa10_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[24] = u_CSAwallace_pg_rca32_csa10_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[25] = u_CSAwallace_pg_rca32_csa10_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[26] = u_CSAwallace_pg_rca32_csa10_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[27] = u_CSAwallace_pg_rca32_csa10_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[28] = u_CSAwallace_pg_rca32_csa10_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[29] = u_CSAwallace_pg_rca32_csa10_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[30] = u_CSAwallace_pg_rca32_csa10_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[31] = u_CSAwallace_pg_rca32_csa10_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[32] = u_CSAwallace_pg_rca32_csa10_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[33] = u_CSAwallace_pg_rca32_csa10_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[34] = u_CSAwallace_pg_rca32_csa10_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[35] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[36] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[37] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[38] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[39] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[40] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11[41] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[5] = u_CSAwallace_pg_rca32_csa11_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[6] = u_CSAwallace_pg_rca32_csa11_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[7] = u_CSAwallace_pg_rca32_csa11_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[8] = u_CSAwallace_pg_rca32_csa11_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[9] = u_CSAwallace_pg_rca32_csa11_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[10] = u_CSAwallace_pg_rca32_csa11_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[11] = u_CSAwallace_pg_rca32_csa11_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[12] = u_CSAwallace_pg_rca32_csa11_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[13] = u_CSAwallace_pg_rca32_csa11_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[14] = u_CSAwallace_pg_rca32_csa11_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[15] = u_CSAwallace_pg_rca32_csa11_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[16] = u_CSAwallace_pg_rca32_csa11_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[17] = u_CSAwallace_pg_rca32_csa11_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[18] = u_CSAwallace_pg_rca32_csa11_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[19] = u_CSAwallace_pg_rca32_csa11_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[20] = u_CSAwallace_pg_rca32_csa11_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[21] = u_CSAwallace_pg_rca32_csa11_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[22] = u_CSAwallace_pg_rca32_csa11_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[23] = u_CSAwallace_pg_rca32_csa11_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[24] = u_CSAwallace_pg_rca32_csa11_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[25] = u_CSAwallace_pg_rca32_csa11_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[26] = u_CSAwallace_pg_rca32_csa11_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[27] = u_CSAwallace_pg_rca32_csa11_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[28] = u_CSAwallace_pg_rca32_csa11_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[29] = u_CSAwallace_pg_rca32_csa11_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[30] = u_CSAwallace_pg_rca32_csa11_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[31] = u_CSAwallace_pg_rca32_csa11_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[32] = u_CSAwallace_pg_rca32_csa11_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[33] = u_CSAwallace_pg_rca32_csa11_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[34] = u_CSAwallace_pg_rca32_csa11_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[35] = u_CSAwallace_pg_rca32_csa11_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[36] = u_CSAwallace_pg_rca32_csa11_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[37] = u_CSAwallace_pg_rca32_csa11_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[38] = u_CSAwallace_pg_rca32_csa11_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[39] = u_CSAwallace_pg_rca32_csa11_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[40] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12[41] = 1'b0;
  csa_component42 csa_component42_u_CSAwallace_pg_rca32_csa17_csa_component_out(.a(u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s11), .b(u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_c11), .c(u_CSAwallace_pg_rca32_csa17_csa_component_u_CSAwallace_pg_rca32_csa_s12), .csa_component42_out(u_CSAwallace_pg_rca32_csa17_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[7] = u_CSAwallace_pg_rca32_csa11_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[8] = u_CSAwallace_pg_rca32_csa11_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[9] = u_CSAwallace_pg_rca32_csa11_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[10] = u_CSAwallace_pg_rca32_csa11_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[11] = u_CSAwallace_pg_rca32_csa11_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[12] = u_CSAwallace_pg_rca32_csa11_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[13] = u_CSAwallace_pg_rca32_csa11_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[14] = u_CSAwallace_pg_rca32_csa11_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[15] = u_CSAwallace_pg_rca32_csa11_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[16] = u_CSAwallace_pg_rca32_csa11_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[17] = u_CSAwallace_pg_rca32_csa11_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[18] = u_CSAwallace_pg_rca32_csa11_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[19] = u_CSAwallace_pg_rca32_csa11_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[20] = u_CSAwallace_pg_rca32_csa11_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[21] = u_CSAwallace_pg_rca32_csa11_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[22] = u_CSAwallace_pg_rca32_csa11_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[23] = u_CSAwallace_pg_rca32_csa11_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[24] = u_CSAwallace_pg_rca32_csa11_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[25] = u_CSAwallace_pg_rca32_csa11_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[26] = u_CSAwallace_pg_rca32_csa11_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[27] = u_CSAwallace_pg_rca32_csa11_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[28] = u_CSAwallace_pg_rca32_csa11_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[29] = u_CSAwallace_pg_rca32_csa11_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[30] = u_CSAwallace_pg_rca32_csa11_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[31] = u_CSAwallace_pg_rca32_csa11_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[32] = u_CSAwallace_pg_rca32_csa11_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[33] = u_CSAwallace_pg_rca32_csa11_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[34] = u_CSAwallace_pg_rca32_csa11_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[35] = u_CSAwallace_pg_rca32_csa11_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[36] = u_CSAwallace_pg_rca32_csa11_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[37] = u_CSAwallace_pg_rca32_csa11_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[38] = u_CSAwallace_pg_rca32_csa11_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[39] = u_CSAwallace_pg_rca32_csa11_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[40] = u_CSAwallace_pg_rca32_csa11_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[41] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[42] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[43] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[44] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[9] = u_CSAwallace_pg_rca32_csa12_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[10] = u_CSAwallace_pg_rca32_csa12_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[11] = u_CSAwallace_pg_rca32_csa12_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[12] = u_CSAwallace_pg_rca32_csa12_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[13] = u_CSAwallace_pg_rca32_csa12_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[14] = u_CSAwallace_pg_rca32_csa12_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[15] = u_CSAwallace_pg_rca32_csa12_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[16] = u_CSAwallace_pg_rca32_csa12_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[17] = u_CSAwallace_pg_rca32_csa12_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[18] = u_CSAwallace_pg_rca32_csa12_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[19] = u_CSAwallace_pg_rca32_csa12_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[20] = u_CSAwallace_pg_rca32_csa12_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[21] = u_CSAwallace_pg_rca32_csa12_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[22] = u_CSAwallace_pg_rca32_csa12_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[23] = u_CSAwallace_pg_rca32_csa12_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[24] = u_CSAwallace_pg_rca32_csa12_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[25] = u_CSAwallace_pg_rca32_csa12_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[26] = u_CSAwallace_pg_rca32_csa12_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[27] = u_CSAwallace_pg_rca32_csa12_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[28] = u_CSAwallace_pg_rca32_csa12_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[29] = u_CSAwallace_pg_rca32_csa12_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[30] = u_CSAwallace_pg_rca32_csa12_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[31] = u_CSAwallace_pg_rca32_csa12_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[32] = u_CSAwallace_pg_rca32_csa12_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[33] = u_CSAwallace_pg_rca32_csa12_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[34] = u_CSAwallace_pg_rca32_csa12_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[35] = u_CSAwallace_pg_rca32_csa12_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[36] = u_CSAwallace_pg_rca32_csa12_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[37] = u_CSAwallace_pg_rca32_csa12_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[38] = u_CSAwallace_pg_rca32_csa12_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[39] = u_CSAwallace_pg_rca32_csa12_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[40] = u_CSAwallace_pg_rca32_csa12_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[41] = u_CSAwallace_pg_rca32_csa12_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[42] = u_CSAwallace_pg_rca32_csa12_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[43] = u_CSAwallace_pg_rca32_csa12_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[44] = u_CSAwallace_pg_rca32_csa12_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[45] = u_CSAwallace_pg_rca32_csa12_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[12] = u_CSAwallace_pg_rca32_csa12_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[13] = u_CSAwallace_pg_rca32_csa12_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[14] = u_CSAwallace_pg_rca32_csa12_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[15] = u_CSAwallace_pg_rca32_csa12_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[16] = u_CSAwallace_pg_rca32_csa12_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[17] = u_CSAwallace_pg_rca32_csa12_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[18] = u_CSAwallace_pg_rca32_csa12_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[19] = u_CSAwallace_pg_rca32_csa12_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[20] = u_CSAwallace_pg_rca32_csa12_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[21] = u_CSAwallace_pg_rca32_csa12_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[22] = u_CSAwallace_pg_rca32_csa12_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[23] = u_CSAwallace_pg_rca32_csa12_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[24] = u_CSAwallace_pg_rca32_csa12_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[25] = u_CSAwallace_pg_rca32_csa12_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[26] = u_CSAwallace_pg_rca32_csa12_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[27] = u_CSAwallace_pg_rca32_csa12_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[28] = u_CSAwallace_pg_rca32_csa12_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[29] = u_CSAwallace_pg_rca32_csa12_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[30] = u_CSAwallace_pg_rca32_csa12_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[31] = u_CSAwallace_pg_rca32_csa12_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[32] = u_CSAwallace_pg_rca32_csa12_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[33] = u_CSAwallace_pg_rca32_csa12_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[34] = u_CSAwallace_pg_rca32_csa12_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[35] = u_CSAwallace_pg_rca32_csa12_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[36] = u_CSAwallace_pg_rca32_csa12_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[37] = u_CSAwallace_pg_rca32_csa12_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[38] = u_CSAwallace_pg_rca32_csa12_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[39] = u_CSAwallace_pg_rca32_csa12_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[40] = u_CSAwallace_pg_rca32_csa12_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[41] = u_CSAwallace_pg_rca32_csa12_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[42] = u_CSAwallace_pg_rca32_csa12_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[43] = u_CSAwallace_pg_rca32_csa12_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[44] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13[47] = 1'b0;
  csa_component48 csa_component48_u_CSAwallace_pg_rca32_csa18_csa_component_out(.a(u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c12), .b(u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_s13), .c(u_CSAwallace_pg_rca32_csa18_csa_component_u_CSAwallace_pg_rca32_csa_c13), .csa_component48_out(u_CSAwallace_pg_rca32_csa18_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[14] = u_CSAwallace_pg_rca32_csa13_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[15] = u_CSAwallace_pg_rca32_csa13_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[16] = u_CSAwallace_pg_rca32_csa13_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[17] = u_CSAwallace_pg_rca32_csa13_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[18] = u_CSAwallace_pg_rca32_csa13_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[19] = u_CSAwallace_pg_rca32_csa13_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[20] = u_CSAwallace_pg_rca32_csa13_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[21] = u_CSAwallace_pg_rca32_csa13_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[22] = u_CSAwallace_pg_rca32_csa13_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[23] = u_CSAwallace_pg_rca32_csa13_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[24] = u_CSAwallace_pg_rca32_csa13_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[25] = u_CSAwallace_pg_rca32_csa13_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[26] = u_CSAwallace_pg_rca32_csa13_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[27] = u_CSAwallace_pg_rca32_csa13_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[28] = u_CSAwallace_pg_rca32_csa13_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[29] = u_CSAwallace_pg_rca32_csa13_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[30] = u_CSAwallace_pg_rca32_csa13_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[31] = u_CSAwallace_pg_rca32_csa13_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[32] = u_CSAwallace_pg_rca32_csa13_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[33] = u_CSAwallace_pg_rca32_csa13_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[34] = u_CSAwallace_pg_rca32_csa13_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[35] = u_CSAwallace_pg_rca32_csa13_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[36] = u_CSAwallace_pg_rca32_csa13_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[37] = u_CSAwallace_pg_rca32_csa13_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[38] = u_CSAwallace_pg_rca32_csa13_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[39] = u_CSAwallace_pg_rca32_csa13_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[40] = u_CSAwallace_pg_rca32_csa13_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[41] = u_CSAwallace_pg_rca32_csa13_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[42] = u_CSAwallace_pg_rca32_csa13_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[43] = u_CSAwallace_pg_rca32_csa13_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[44] = u_CSAwallace_pg_rca32_csa13_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[45] = u_CSAwallace_pg_rca32_csa13_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[46] = u_CSAwallace_pg_rca32_csa13_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[47] = u_CSAwallace_pg_rca32_csa13_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[48] = u_CSAwallace_pg_rca32_csa13_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[49] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[50] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[16] = u_CSAwallace_pg_rca32_csa13_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[17] = u_CSAwallace_pg_rca32_csa13_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[18] = u_CSAwallace_pg_rca32_csa13_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[19] = u_CSAwallace_pg_rca32_csa13_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[20] = u_CSAwallace_pg_rca32_csa13_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[21] = u_CSAwallace_pg_rca32_csa13_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[22] = u_CSAwallace_pg_rca32_csa13_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[23] = u_CSAwallace_pg_rca32_csa13_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[24] = u_CSAwallace_pg_rca32_csa13_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[25] = u_CSAwallace_pg_rca32_csa13_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[26] = u_CSAwallace_pg_rca32_csa13_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[27] = u_CSAwallace_pg_rca32_csa13_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[28] = u_CSAwallace_pg_rca32_csa13_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[29] = u_CSAwallace_pg_rca32_csa13_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[30] = u_CSAwallace_pg_rca32_csa13_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[31] = u_CSAwallace_pg_rca32_csa13_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[32] = u_CSAwallace_pg_rca32_csa13_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[33] = u_CSAwallace_pg_rca32_csa13_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[34] = u_CSAwallace_pg_rca32_csa13_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[35] = u_CSAwallace_pg_rca32_csa13_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[36] = u_CSAwallace_pg_rca32_csa13_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[37] = u_CSAwallace_pg_rca32_csa13_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[38] = u_CSAwallace_pg_rca32_csa13_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[39] = u_CSAwallace_pg_rca32_csa13_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[40] = u_CSAwallace_pg_rca32_csa13_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[41] = u_CSAwallace_pg_rca32_csa13_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[42] = u_CSAwallace_pg_rca32_csa13_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[43] = u_CSAwallace_pg_rca32_csa13_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[44] = u_CSAwallace_pg_rca32_csa13_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[45] = u_CSAwallace_pg_rca32_csa13_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[46] = u_CSAwallace_pg_rca32_csa13_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[47] = u_CSAwallace_pg_rca32_csa13_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[48] = u_CSAwallace_pg_rca32_csa13_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[49] = u_CSAwallace_pg_rca32_csa13_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[50] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[18] = u_CSAwallace_pg_rca32_csa14_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[19] = u_CSAwallace_pg_rca32_csa14_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[20] = u_CSAwallace_pg_rca32_csa14_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[21] = u_CSAwallace_pg_rca32_csa14_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[22] = u_CSAwallace_pg_rca32_csa14_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[23] = u_CSAwallace_pg_rca32_csa14_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[24] = u_CSAwallace_pg_rca32_csa14_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[25] = u_CSAwallace_pg_rca32_csa14_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[26] = u_CSAwallace_pg_rca32_csa14_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[27] = u_CSAwallace_pg_rca32_csa14_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[28] = u_CSAwallace_pg_rca32_csa14_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[29] = u_CSAwallace_pg_rca32_csa14_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[30] = u_CSAwallace_pg_rca32_csa14_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[31] = u_CSAwallace_pg_rca32_csa14_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[32] = u_CSAwallace_pg_rca32_csa14_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[33] = u_CSAwallace_pg_rca32_csa14_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[34] = u_CSAwallace_pg_rca32_csa14_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[35] = u_CSAwallace_pg_rca32_csa14_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[36] = u_CSAwallace_pg_rca32_csa14_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[37] = u_CSAwallace_pg_rca32_csa14_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[38] = u_CSAwallace_pg_rca32_csa14_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[39] = u_CSAwallace_pg_rca32_csa14_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[40] = u_CSAwallace_pg_rca32_csa14_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[41] = u_CSAwallace_pg_rca32_csa14_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[42] = u_CSAwallace_pg_rca32_csa14_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[43] = u_CSAwallace_pg_rca32_csa14_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[44] = u_CSAwallace_pg_rca32_csa14_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[45] = u_CSAwallace_pg_rca32_csa14_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[46] = u_CSAwallace_pg_rca32_csa14_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[47] = u_CSAwallace_pg_rca32_csa14_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[48] = u_CSAwallace_pg_rca32_csa14_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[49] = u_CSAwallace_pg_rca32_csa14_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[50] = u_CSAwallace_pg_rca32_csa14_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[51] = u_CSAwallace_pg_rca32_csa14_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[52] = u_CSAwallace_pg_rca32_csa14_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[53] = u_CSAwallace_pg_rca32_csa14_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[54] = u_CSAwallace_pg_rca32_csa14_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15[56] = 1'b0;
  csa_component57 csa_component57_u_CSAwallace_pg_rca32_csa19_csa_component_out(.a(u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s14), .b(u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_c14), .c(u_CSAwallace_pg_rca32_csa19_csa_component_u_CSAwallace_pg_rca32_csa_s15), .csa_component57_out(u_CSAwallace_pg_rca32_csa19_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[21] = u_CSAwallace_pg_rca32_csa14_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[22] = u_CSAwallace_pg_rca32_csa14_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[23] = u_CSAwallace_pg_rca32_csa14_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[24] = u_CSAwallace_pg_rca32_csa14_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[25] = u_CSAwallace_pg_rca32_csa14_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[26] = u_CSAwallace_pg_rca32_csa14_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[27] = u_CSAwallace_pg_rca32_csa14_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[28] = u_CSAwallace_pg_rca32_csa14_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[29] = u_CSAwallace_pg_rca32_csa14_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[30] = u_CSAwallace_pg_rca32_csa14_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[31] = u_CSAwallace_pg_rca32_csa14_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[32] = u_CSAwallace_pg_rca32_csa14_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[33] = u_CSAwallace_pg_rca32_csa14_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[34] = u_CSAwallace_pg_rca32_csa14_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[35] = u_CSAwallace_pg_rca32_csa14_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[36] = u_CSAwallace_pg_rca32_csa14_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[37] = u_CSAwallace_pg_rca32_csa14_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[38] = u_CSAwallace_pg_rca32_csa14_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[39] = u_CSAwallace_pg_rca32_csa14_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[40] = u_CSAwallace_pg_rca32_csa14_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[41] = u_CSAwallace_pg_rca32_csa14_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[42] = u_CSAwallace_pg_rca32_csa14_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[43] = u_CSAwallace_pg_rca32_csa14_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[44] = u_CSAwallace_pg_rca32_csa14_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[45] = u_CSAwallace_pg_rca32_csa14_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[46] = u_CSAwallace_pg_rca32_csa14_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[47] = u_CSAwallace_pg_rca32_csa14_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[48] = u_CSAwallace_pg_rca32_csa14_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[49] = u_CSAwallace_pg_rca32_csa14_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[50] = u_CSAwallace_pg_rca32_csa14_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[51] = u_CSAwallace_pg_rca32_csa14_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[52] = u_CSAwallace_pg_rca32_csa14_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[23] = u_CSAwallace_pg_rca32_csa15_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[24] = u_CSAwallace_pg_rca32_csa15_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[25] = u_CSAwallace_pg_rca32_csa15_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[26] = u_CSAwallace_pg_rca32_csa15_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[27] = u_CSAwallace_pg_rca32_csa15_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[28] = u_CSAwallace_pg_rca32_csa15_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[29] = u_CSAwallace_pg_rca32_csa15_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[30] = u_CSAwallace_pg_rca32_csa15_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[31] = u_CSAwallace_pg_rca32_csa15_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[32] = u_CSAwallace_pg_rca32_csa15_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[33] = u_CSAwallace_pg_rca32_csa15_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[34] = u_CSAwallace_pg_rca32_csa15_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[35] = u_CSAwallace_pg_rca32_csa15_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[36] = u_CSAwallace_pg_rca32_csa15_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[37] = u_CSAwallace_pg_rca32_csa15_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[38] = u_CSAwallace_pg_rca32_csa15_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[39] = u_CSAwallace_pg_rca32_csa15_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[40] = u_CSAwallace_pg_rca32_csa15_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[41] = u_CSAwallace_pg_rca32_csa15_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[42] = u_CSAwallace_pg_rca32_csa15_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[43] = u_CSAwallace_pg_rca32_csa15_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[44] = u_CSAwallace_pg_rca32_csa15_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[45] = u_CSAwallace_pg_rca32_csa15_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[46] = u_CSAwallace_pg_rca32_csa15_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[47] = u_CSAwallace_pg_rca32_csa15_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[48] = u_CSAwallace_pg_rca32_csa15_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[49] = u_CSAwallace_pg_rca32_csa15_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[50] = u_CSAwallace_pg_rca32_csa15_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[51] = u_CSAwallace_pg_rca32_csa15_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[52] = u_CSAwallace_pg_rca32_csa15_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[53] = u_CSAwallace_pg_rca32_csa15_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[54] = u_CSAwallace_pg_rca32_csa15_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[55] = u_CSAwallace_pg_rca32_csa15_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[56] = u_CSAwallace_pg_rca32_csa15_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[57] = u_CSAwallace_pg_rca32_csa15_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[25] = u_CSAwallace_pg_rca32_csa15_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[26] = u_CSAwallace_pg_rca32_csa15_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[27] = u_CSAwallace_pg_rca32_csa15_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[28] = u_CSAwallace_pg_rca32_csa15_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[29] = u_CSAwallace_pg_rca32_csa15_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[30] = u_CSAwallace_pg_rca32_csa15_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[31] = u_CSAwallace_pg_rca32_csa15_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[32] = u_CSAwallace_pg_rca32_csa15_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[33] = u_CSAwallace_pg_rca32_csa15_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[34] = u_CSAwallace_pg_rca32_csa15_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[35] = u_CSAwallace_pg_rca32_csa15_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[36] = u_CSAwallace_pg_rca32_csa15_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[37] = u_CSAwallace_pg_rca32_csa15_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[38] = u_CSAwallace_pg_rca32_csa15_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[39] = u_CSAwallace_pg_rca32_csa15_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[40] = u_CSAwallace_pg_rca32_csa15_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[41] = u_CSAwallace_pg_rca32_csa15_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[42] = u_CSAwallace_pg_rca32_csa15_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[43] = u_CSAwallace_pg_rca32_csa15_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[44] = u_CSAwallace_pg_rca32_csa15_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[45] = u_CSAwallace_pg_rca32_csa15_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[46] = u_CSAwallace_pg_rca32_csa15_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[47] = u_CSAwallace_pg_rca32_csa15_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[48] = u_CSAwallace_pg_rca32_csa15_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[49] = u_CSAwallace_pg_rca32_csa15_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[50] = u_CSAwallace_pg_rca32_csa15_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[51] = u_CSAwallace_pg_rca32_csa15_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[52] = u_CSAwallace_pg_rca32_csa15_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[53] = u_CSAwallace_pg_rca32_csa15_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[54] = u_CSAwallace_pg_rca32_csa15_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[55] = u_CSAwallace_pg_rca32_csa15_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[56] = u_CSAwallace_pg_rca32_csa15_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[57] = u_CSAwallace_pg_rca32_csa15_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[58] = u_CSAwallace_pg_rca32_csa15_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16[59] = 1'b0;
  csa_component60 csa_component60_u_CSAwallace_pg_rca32_csa20_csa_component_out(.a(u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c15), .b(u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_s16), .c(u_CSAwallace_pg_rca32_csa20_csa_component_u_CSAwallace_pg_rca32_csa_c16), .csa_component60_out(u_CSAwallace_pg_rca32_csa20_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[27] = u_CSAwallace_pg_rca32_csa16_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[28] = u_CSAwallace_pg_rca32_csa16_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[29] = u_CSAwallace_pg_rca32_csa16_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[30] = u_CSAwallace_pg_rca32_csa16_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[31] = u_CSAwallace_pg_rca32_csa16_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[32] = u_CSAwallace_pg_rca32_csa16_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[33] = u_CSAwallace_pg_rca32_csa16_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[34] = u_CSAwallace_pg_rca32_csa16_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[35] = u_CSAwallace_pg_rca32_csa16_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[36] = u_CSAwallace_pg_rca32_csa16_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[37] = u_CSAwallace_pg_rca32_csa16_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[38] = u_CSAwallace_pg_rca32_csa16_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[39] = u_CSAwallace_pg_rca32_csa16_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[40] = u_CSAwallace_pg_rca32_csa16_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[41] = u_CSAwallace_pg_rca32_csa16_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[42] = u_CSAwallace_pg_rca32_csa16_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[43] = u_CSAwallace_pg_rca32_csa16_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[44] = u_CSAwallace_pg_rca32_csa16_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[45] = u_CSAwallace_pg_rca32_csa16_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[46] = u_CSAwallace_pg_rca32_csa16_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[47] = u_CSAwallace_pg_rca32_csa16_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[48] = u_CSAwallace_pg_rca32_csa16_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[49] = u_CSAwallace_pg_rca32_csa16_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[50] = u_CSAwallace_pg_rca32_csa16_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[51] = u_CSAwallace_pg_rca32_csa16_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[52] = u_CSAwallace_pg_rca32_csa16_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[53] = u_CSAwallace_pg_rca32_csa16_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[54] = u_CSAwallace_pg_rca32_csa16_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[55] = u_CSAwallace_pg_rca32_csa16_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[56] = u_CSAwallace_pg_rca32_csa16_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[57] = u_CSAwallace_pg_rca32_csa16_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[58] = u_CSAwallace_pg_rca32_csa16_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[59] = u_CSAwallace_pg_rca32_csa16_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[60] = u_CSAwallace_pg_rca32_csa16_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[61] = u_CSAwallace_pg_rca32_csa16_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[27] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[28] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[29] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[30] = u_CSAwallace_pg_rca32_csa16_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[31] = u_CSAwallace_pg_rca32_csa16_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[32] = u_CSAwallace_pg_rca32_csa16_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[33] = u_CSAwallace_pg_rca32_csa16_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[34] = u_CSAwallace_pg_rca32_csa16_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[35] = u_CSAwallace_pg_rca32_csa16_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[36] = u_CSAwallace_pg_rca32_csa16_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[37] = u_CSAwallace_pg_rca32_csa16_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[38] = u_CSAwallace_pg_rca32_csa16_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[39] = u_CSAwallace_pg_rca32_csa16_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[40] = u_CSAwallace_pg_rca32_csa16_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[41] = u_CSAwallace_pg_rca32_csa16_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[42] = u_CSAwallace_pg_rca32_csa16_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[43] = u_CSAwallace_pg_rca32_csa16_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[44] = u_CSAwallace_pg_rca32_csa16_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[45] = u_CSAwallace_pg_rca32_csa16_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[46] = u_CSAwallace_pg_rca32_csa16_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[47] = u_CSAwallace_pg_rca32_csa16_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[48] = u_CSAwallace_pg_rca32_csa16_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[49] = u_CSAwallace_pg_rca32_csa16_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[50] = u_CSAwallace_pg_rca32_csa16_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[51] = u_CSAwallace_pg_rca32_csa16_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[52] = u_CSAwallace_pg_rca32_csa16_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[53] = u_CSAwallace_pg_rca32_csa16_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[54] = u_CSAwallace_pg_rca32_csa16_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[55] = u_CSAwallace_pg_rca32_csa16_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[56] = u_CSAwallace_pg_rca32_csa16_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[57] = u_CSAwallace_pg_rca32_csa16_csa_component_out[120];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[58] = u_CSAwallace_pg_rca32_csa16_csa_component_out[121];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[59] = u_CSAwallace_pg_rca32_csa16_csa_component_out[122];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[60] = u_CSAwallace_pg_rca32_csa16_csa_component_out[123];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[61] = u_CSAwallace_pg_rca32_csa16_csa_component_out[124];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[27] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[28] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[29] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[30] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[31] = u_CSAwallace_pg_rca32_and_0_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[32] = u_CSAwallace_pg_rca32_and_1_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[33] = u_CSAwallace_pg_rca32_and_2_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[34] = u_CSAwallace_pg_rca32_and_3_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[35] = u_CSAwallace_pg_rca32_and_4_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[36] = u_CSAwallace_pg_rca32_and_5_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[37] = u_CSAwallace_pg_rca32_and_6_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[38] = u_CSAwallace_pg_rca32_and_7_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[39] = u_CSAwallace_pg_rca32_and_8_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[40] = u_CSAwallace_pg_rca32_and_9_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[41] = u_CSAwallace_pg_rca32_and_10_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[42] = u_CSAwallace_pg_rca32_and_11_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[43] = u_CSAwallace_pg_rca32_and_12_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[44] = u_CSAwallace_pg_rca32_and_13_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[45] = u_CSAwallace_pg_rca32_and_14_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[46] = u_CSAwallace_pg_rca32_and_15_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[47] = u_CSAwallace_pg_rca32_and_16_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[48] = u_CSAwallace_pg_rca32_and_17_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[49] = u_CSAwallace_pg_rca32_and_18_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[50] = u_CSAwallace_pg_rca32_and_19_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[51] = u_CSAwallace_pg_rca32_and_20_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[52] = u_CSAwallace_pg_rca32_and_21_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[53] = u_CSAwallace_pg_rca32_and_22_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[54] = u_CSAwallace_pg_rca32_and_23_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[55] = u_CSAwallace_pg_rca32_and_24_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[56] = u_CSAwallace_pg_rca32_and_25_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[57] = u_CSAwallace_pg_rca32_and_26_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[58] = u_CSAwallace_pg_rca32_and_27_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[59] = u_CSAwallace_pg_rca32_and_28_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[60] = u_CSAwallace_pg_rca32_and_29_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[61] = u_CSAwallace_pg_rca32_and_30_31[0];
  assign u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31[62] = u_CSAwallace_pg_rca32_and_31_31[0];
  csa_component63 csa_component63_u_CSAwallace_pg_rca32_csa21_csa_component_out(.a(u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_s17), .b(u_CSAwallace_pg_rca32_csa21_csa_component_u_CSAwallace_pg_rca32_csa_c17), .c(u_CSAwallace_pg_rca32_csa21_csa_component_pp_row31), .csa_component63_out(u_CSAwallace_pg_rca32_csa21_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[0] = u_CSAwallace_pg_rca32_csa17_csa_component_out[0];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[1] = u_CSAwallace_pg_rca32_csa17_csa_component_out[1];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[2] = u_CSAwallace_pg_rca32_csa17_csa_component_out[2];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[3] = u_CSAwallace_pg_rca32_csa17_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[4] = u_CSAwallace_pg_rca32_csa17_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[5] = u_CSAwallace_pg_rca32_csa17_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[6] = u_CSAwallace_pg_rca32_csa17_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[7] = u_CSAwallace_pg_rca32_csa17_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[8] = u_CSAwallace_pg_rca32_csa17_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[9] = u_CSAwallace_pg_rca32_csa17_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[10] = u_CSAwallace_pg_rca32_csa17_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[11] = u_CSAwallace_pg_rca32_csa17_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[12] = u_CSAwallace_pg_rca32_csa17_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[13] = u_CSAwallace_pg_rca32_csa17_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[14] = u_CSAwallace_pg_rca32_csa17_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[15] = u_CSAwallace_pg_rca32_csa17_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[16] = u_CSAwallace_pg_rca32_csa17_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[17] = u_CSAwallace_pg_rca32_csa17_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[18] = u_CSAwallace_pg_rca32_csa17_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[19] = u_CSAwallace_pg_rca32_csa17_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[20] = u_CSAwallace_pg_rca32_csa17_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[21] = u_CSAwallace_pg_rca32_csa17_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[22] = u_CSAwallace_pg_rca32_csa17_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[23] = u_CSAwallace_pg_rca32_csa17_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[24] = u_CSAwallace_pg_rca32_csa17_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[25] = u_CSAwallace_pg_rca32_csa17_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[26] = u_CSAwallace_pg_rca32_csa17_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[27] = u_CSAwallace_pg_rca32_csa17_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[28] = u_CSAwallace_pg_rca32_csa17_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[29] = u_CSAwallace_pg_rca32_csa17_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[30] = u_CSAwallace_pg_rca32_csa17_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[31] = u_CSAwallace_pg_rca32_csa17_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[32] = u_CSAwallace_pg_rca32_csa17_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[33] = u_CSAwallace_pg_rca32_csa17_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[34] = u_CSAwallace_pg_rca32_csa17_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[35] = u_CSAwallace_pg_rca32_csa17_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[36] = u_CSAwallace_pg_rca32_csa17_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[37] = u_CSAwallace_pg_rca32_csa17_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[38] = u_CSAwallace_pg_rca32_csa17_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[39] = u_CSAwallace_pg_rca32_csa17_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[40] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[41] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[42] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[43] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[44] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[4] = u_CSAwallace_pg_rca32_csa17_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[5] = u_CSAwallace_pg_rca32_csa17_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[6] = u_CSAwallace_pg_rca32_csa17_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[7] = u_CSAwallace_pg_rca32_csa17_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[8] = u_CSAwallace_pg_rca32_csa17_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[9] = u_CSAwallace_pg_rca32_csa17_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[10] = u_CSAwallace_pg_rca32_csa17_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[11] = u_CSAwallace_pg_rca32_csa17_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[12] = u_CSAwallace_pg_rca32_csa17_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[13] = u_CSAwallace_pg_rca32_csa17_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[14] = u_CSAwallace_pg_rca32_csa17_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[15] = u_CSAwallace_pg_rca32_csa17_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[16] = u_CSAwallace_pg_rca32_csa17_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[17] = u_CSAwallace_pg_rca32_csa17_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[18] = u_CSAwallace_pg_rca32_csa17_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[19] = u_CSAwallace_pg_rca32_csa17_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[20] = u_CSAwallace_pg_rca32_csa17_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[21] = u_CSAwallace_pg_rca32_csa17_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[22] = u_CSAwallace_pg_rca32_csa17_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[23] = u_CSAwallace_pg_rca32_csa17_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[24] = u_CSAwallace_pg_rca32_csa17_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[25] = u_CSAwallace_pg_rca32_csa17_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[26] = u_CSAwallace_pg_rca32_csa17_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[27] = u_CSAwallace_pg_rca32_csa17_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[28] = u_CSAwallace_pg_rca32_csa17_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[29] = u_CSAwallace_pg_rca32_csa17_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[30] = u_CSAwallace_pg_rca32_csa17_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[31] = u_CSAwallace_pg_rca32_csa17_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[32] = u_CSAwallace_pg_rca32_csa17_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[33] = u_CSAwallace_pg_rca32_csa17_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[34] = u_CSAwallace_pg_rca32_csa17_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[35] = u_CSAwallace_pg_rca32_csa17_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[36] = u_CSAwallace_pg_rca32_csa17_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[37] = u_CSAwallace_pg_rca32_csa17_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[38] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[39] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[40] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[41] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[42] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[43] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[44] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[7] = u_CSAwallace_pg_rca32_csa18_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[8] = u_CSAwallace_pg_rca32_csa18_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[9] = u_CSAwallace_pg_rca32_csa18_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[10] = u_CSAwallace_pg_rca32_csa18_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[11] = u_CSAwallace_pg_rca32_csa18_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[12] = u_CSAwallace_pg_rca32_csa18_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[13] = u_CSAwallace_pg_rca32_csa18_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[14] = u_CSAwallace_pg_rca32_csa18_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[15] = u_CSAwallace_pg_rca32_csa18_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[16] = u_CSAwallace_pg_rca32_csa18_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[17] = u_CSAwallace_pg_rca32_csa18_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[18] = u_CSAwallace_pg_rca32_csa18_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[19] = u_CSAwallace_pg_rca32_csa18_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[20] = u_CSAwallace_pg_rca32_csa18_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[21] = u_CSAwallace_pg_rca32_csa18_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[22] = u_CSAwallace_pg_rca32_csa18_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[23] = u_CSAwallace_pg_rca32_csa18_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[24] = u_CSAwallace_pg_rca32_csa18_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[25] = u_CSAwallace_pg_rca32_csa18_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[26] = u_CSAwallace_pg_rca32_csa18_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[27] = u_CSAwallace_pg_rca32_csa18_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[28] = u_CSAwallace_pg_rca32_csa18_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[29] = u_CSAwallace_pg_rca32_csa18_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[30] = u_CSAwallace_pg_rca32_csa18_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[31] = u_CSAwallace_pg_rca32_csa18_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[32] = u_CSAwallace_pg_rca32_csa18_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[33] = u_CSAwallace_pg_rca32_csa18_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[34] = u_CSAwallace_pg_rca32_csa18_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[35] = u_CSAwallace_pg_rca32_csa18_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[36] = u_CSAwallace_pg_rca32_csa18_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[37] = u_CSAwallace_pg_rca32_csa18_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[38] = u_CSAwallace_pg_rca32_csa18_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[39] = u_CSAwallace_pg_rca32_csa18_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[40] = u_CSAwallace_pg_rca32_csa18_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[41] = u_CSAwallace_pg_rca32_csa18_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[42] = u_CSAwallace_pg_rca32_csa18_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[43] = u_CSAwallace_pg_rca32_csa18_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[44] = u_CSAwallace_pg_rca32_csa18_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[45] = u_CSAwallace_pg_rca32_csa18_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19[48] = 1'b0;
  csa_component49 csa_component49_u_CSAwallace_pg_rca32_csa22_csa_component_out(.a(u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s18), .b(u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_c18), .c(u_CSAwallace_pg_rca32_csa22_csa_component_u_CSAwallace_pg_rca32_csa_s19), .csa_component49_out(u_CSAwallace_pg_rca32_csa22_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[10] = u_CSAwallace_pg_rca32_csa18_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[11] = u_CSAwallace_pg_rca32_csa18_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[12] = u_CSAwallace_pg_rca32_csa18_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[13] = u_CSAwallace_pg_rca32_csa18_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[14] = u_CSAwallace_pg_rca32_csa18_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[15] = u_CSAwallace_pg_rca32_csa18_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[16] = u_CSAwallace_pg_rca32_csa18_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[17] = u_CSAwallace_pg_rca32_csa18_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[18] = u_CSAwallace_pg_rca32_csa18_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[19] = u_CSAwallace_pg_rca32_csa18_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[20] = u_CSAwallace_pg_rca32_csa18_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[21] = u_CSAwallace_pg_rca32_csa18_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[22] = u_CSAwallace_pg_rca32_csa18_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[23] = u_CSAwallace_pg_rca32_csa18_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[24] = u_CSAwallace_pg_rca32_csa18_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[25] = u_CSAwallace_pg_rca32_csa18_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[26] = u_CSAwallace_pg_rca32_csa18_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[27] = u_CSAwallace_pg_rca32_csa18_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[28] = u_CSAwallace_pg_rca32_csa18_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[29] = u_CSAwallace_pg_rca32_csa18_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[30] = u_CSAwallace_pg_rca32_csa18_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[31] = u_CSAwallace_pg_rca32_csa18_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[32] = u_CSAwallace_pg_rca32_csa18_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[33] = u_CSAwallace_pg_rca32_csa18_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[34] = u_CSAwallace_pg_rca32_csa18_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[35] = u_CSAwallace_pg_rca32_csa18_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[36] = u_CSAwallace_pg_rca32_csa18_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[37] = u_CSAwallace_pg_rca32_csa18_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[38] = u_CSAwallace_pg_rca32_csa18_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[39] = u_CSAwallace_pg_rca32_csa18_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[40] = u_CSAwallace_pg_rca32_csa18_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[41] = u_CSAwallace_pg_rca32_csa18_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[42] = u_CSAwallace_pg_rca32_csa18_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[43] = u_CSAwallace_pg_rca32_csa18_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[44] = u_CSAwallace_pg_rca32_csa18_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[49] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[50] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[14] = u_CSAwallace_pg_rca32_csa19_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[15] = u_CSAwallace_pg_rca32_csa19_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[16] = u_CSAwallace_pg_rca32_csa19_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[17] = u_CSAwallace_pg_rca32_csa19_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[18] = u_CSAwallace_pg_rca32_csa19_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[19] = u_CSAwallace_pg_rca32_csa19_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[20] = u_CSAwallace_pg_rca32_csa19_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[21] = u_CSAwallace_pg_rca32_csa19_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[22] = u_CSAwallace_pg_rca32_csa19_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[23] = u_CSAwallace_pg_rca32_csa19_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[24] = u_CSAwallace_pg_rca32_csa19_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[25] = u_CSAwallace_pg_rca32_csa19_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[26] = u_CSAwallace_pg_rca32_csa19_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[27] = u_CSAwallace_pg_rca32_csa19_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[28] = u_CSAwallace_pg_rca32_csa19_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[29] = u_CSAwallace_pg_rca32_csa19_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[30] = u_CSAwallace_pg_rca32_csa19_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[31] = u_CSAwallace_pg_rca32_csa19_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[32] = u_CSAwallace_pg_rca32_csa19_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[33] = u_CSAwallace_pg_rca32_csa19_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[34] = u_CSAwallace_pg_rca32_csa19_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[35] = u_CSAwallace_pg_rca32_csa19_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[36] = u_CSAwallace_pg_rca32_csa19_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[37] = u_CSAwallace_pg_rca32_csa19_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[38] = u_CSAwallace_pg_rca32_csa19_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[39] = u_CSAwallace_pg_rca32_csa19_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[40] = u_CSAwallace_pg_rca32_csa19_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[41] = u_CSAwallace_pg_rca32_csa19_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[42] = u_CSAwallace_pg_rca32_csa19_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[43] = u_CSAwallace_pg_rca32_csa19_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[44] = u_CSAwallace_pg_rca32_csa19_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[45] = u_CSAwallace_pg_rca32_csa19_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[46] = u_CSAwallace_pg_rca32_csa19_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[47] = u_CSAwallace_pg_rca32_csa19_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[48] = u_CSAwallace_pg_rca32_csa19_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[49] = u_CSAwallace_pg_rca32_csa19_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[50] = u_CSAwallace_pg_rca32_csa19_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[51] = u_CSAwallace_pg_rca32_csa19_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[52] = u_CSAwallace_pg_rca32_csa19_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[53] = u_CSAwallace_pg_rca32_csa19_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[54] = u_CSAwallace_pg_rca32_csa19_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[17] = u_CSAwallace_pg_rca32_csa19_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[18] = u_CSAwallace_pg_rca32_csa19_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[19] = u_CSAwallace_pg_rca32_csa19_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[20] = u_CSAwallace_pg_rca32_csa19_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[21] = u_CSAwallace_pg_rca32_csa19_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[22] = u_CSAwallace_pg_rca32_csa19_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[23] = u_CSAwallace_pg_rca32_csa19_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[24] = u_CSAwallace_pg_rca32_csa19_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[25] = u_CSAwallace_pg_rca32_csa19_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[26] = u_CSAwallace_pg_rca32_csa19_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[27] = u_CSAwallace_pg_rca32_csa19_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[28] = u_CSAwallace_pg_rca32_csa19_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[29] = u_CSAwallace_pg_rca32_csa19_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[30] = u_CSAwallace_pg_rca32_csa19_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[31] = u_CSAwallace_pg_rca32_csa19_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[32] = u_CSAwallace_pg_rca32_csa19_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[33] = u_CSAwallace_pg_rca32_csa19_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[34] = u_CSAwallace_pg_rca32_csa19_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[35] = u_CSAwallace_pg_rca32_csa19_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[36] = u_CSAwallace_pg_rca32_csa19_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[37] = u_CSAwallace_pg_rca32_csa19_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[38] = u_CSAwallace_pg_rca32_csa19_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[39] = u_CSAwallace_pg_rca32_csa19_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[40] = u_CSAwallace_pg_rca32_csa19_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[41] = u_CSAwallace_pg_rca32_csa19_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[42] = u_CSAwallace_pg_rca32_csa19_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[43] = u_CSAwallace_pg_rca32_csa19_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[44] = u_CSAwallace_pg_rca32_csa19_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[45] = u_CSAwallace_pg_rca32_csa19_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[46] = u_CSAwallace_pg_rca32_csa19_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[47] = u_CSAwallace_pg_rca32_csa19_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[48] = u_CSAwallace_pg_rca32_csa19_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[49] = u_CSAwallace_pg_rca32_csa19_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[50] = u_CSAwallace_pg_rca32_csa19_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20[57] = 1'b0;
  csa_component58 csa_component58_u_CSAwallace_pg_rca32_csa23_csa_component_out(.a(u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c19), .b(u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_s20), .c(u_CSAwallace_pg_rca32_csa23_csa_component_u_CSAwallace_pg_rca32_csa_c20), .csa_component58_out(u_CSAwallace_pg_rca32_csa23_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[21] = u_CSAwallace_pg_rca32_csa20_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[22] = u_CSAwallace_pg_rca32_csa20_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[23] = u_CSAwallace_pg_rca32_csa20_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[24] = u_CSAwallace_pg_rca32_csa20_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[25] = u_CSAwallace_pg_rca32_csa20_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[26] = u_CSAwallace_pg_rca32_csa20_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[27] = u_CSAwallace_pg_rca32_csa20_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[28] = u_CSAwallace_pg_rca32_csa20_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[29] = u_CSAwallace_pg_rca32_csa20_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[30] = u_CSAwallace_pg_rca32_csa20_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[31] = u_CSAwallace_pg_rca32_csa20_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[32] = u_CSAwallace_pg_rca32_csa20_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[33] = u_CSAwallace_pg_rca32_csa20_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[34] = u_CSAwallace_pg_rca32_csa20_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[35] = u_CSAwallace_pg_rca32_csa20_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[36] = u_CSAwallace_pg_rca32_csa20_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[37] = u_CSAwallace_pg_rca32_csa20_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[38] = u_CSAwallace_pg_rca32_csa20_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[39] = u_CSAwallace_pg_rca32_csa20_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[40] = u_CSAwallace_pg_rca32_csa20_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[41] = u_CSAwallace_pg_rca32_csa20_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[42] = u_CSAwallace_pg_rca32_csa20_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[43] = u_CSAwallace_pg_rca32_csa20_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[44] = u_CSAwallace_pg_rca32_csa20_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[45] = u_CSAwallace_pg_rca32_csa20_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[46] = u_CSAwallace_pg_rca32_csa20_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[47] = u_CSAwallace_pg_rca32_csa20_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[48] = u_CSAwallace_pg_rca32_csa20_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[49] = u_CSAwallace_pg_rca32_csa20_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[50] = u_CSAwallace_pg_rca32_csa20_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[51] = u_CSAwallace_pg_rca32_csa20_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[52] = u_CSAwallace_pg_rca32_csa20_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[53] = u_CSAwallace_pg_rca32_csa20_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[54] = u_CSAwallace_pg_rca32_csa20_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[55] = u_CSAwallace_pg_rca32_csa20_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[56] = u_CSAwallace_pg_rca32_csa20_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[57] = u_CSAwallace_pg_rca32_csa20_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[58] = u_CSAwallace_pg_rca32_csa20_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[24] = u_CSAwallace_pg_rca32_csa20_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[25] = u_CSAwallace_pg_rca32_csa20_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[26] = u_CSAwallace_pg_rca32_csa20_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[27] = u_CSAwallace_pg_rca32_csa20_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[28] = u_CSAwallace_pg_rca32_csa20_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[29] = u_CSAwallace_pg_rca32_csa20_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[30] = u_CSAwallace_pg_rca32_csa20_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[31] = u_CSAwallace_pg_rca32_csa20_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[32] = u_CSAwallace_pg_rca32_csa20_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[33] = u_CSAwallace_pg_rca32_csa20_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[34] = u_CSAwallace_pg_rca32_csa20_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[35] = u_CSAwallace_pg_rca32_csa20_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[36] = u_CSAwallace_pg_rca32_csa20_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[37] = u_CSAwallace_pg_rca32_csa20_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[38] = u_CSAwallace_pg_rca32_csa20_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[39] = u_CSAwallace_pg_rca32_csa20_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[40] = u_CSAwallace_pg_rca32_csa20_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[41] = u_CSAwallace_pg_rca32_csa20_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[42] = u_CSAwallace_pg_rca32_csa20_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[43] = u_CSAwallace_pg_rca32_csa20_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[44] = u_CSAwallace_pg_rca32_csa20_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[45] = u_CSAwallace_pg_rca32_csa20_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[46] = u_CSAwallace_pg_rca32_csa20_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[47] = u_CSAwallace_pg_rca32_csa20_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[48] = u_CSAwallace_pg_rca32_csa20_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[49] = u_CSAwallace_pg_rca32_csa20_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[50] = u_CSAwallace_pg_rca32_csa20_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[51] = u_CSAwallace_pg_rca32_csa20_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[52] = u_CSAwallace_pg_rca32_csa20_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[53] = u_CSAwallace_pg_rca32_csa20_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[54] = u_CSAwallace_pg_rca32_csa20_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[55] = u_CSAwallace_pg_rca32_csa20_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[56] = u_CSAwallace_pg_rca32_csa20_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[57] = u_CSAwallace_pg_rca32_csa20_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[58] = u_CSAwallace_pg_rca32_csa20_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[27] = u_CSAwallace_pg_rca32_csa21_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[28] = u_CSAwallace_pg_rca32_csa21_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[29] = u_CSAwallace_pg_rca32_csa21_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[30] = u_CSAwallace_pg_rca32_csa21_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[31] = u_CSAwallace_pg_rca32_csa21_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[32] = u_CSAwallace_pg_rca32_csa21_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[33] = u_CSAwallace_pg_rca32_csa21_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[34] = u_CSAwallace_pg_rca32_csa21_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[35] = u_CSAwallace_pg_rca32_csa21_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[36] = u_CSAwallace_pg_rca32_csa21_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[37] = u_CSAwallace_pg_rca32_csa21_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[38] = u_CSAwallace_pg_rca32_csa21_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[39] = u_CSAwallace_pg_rca32_csa21_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[40] = u_CSAwallace_pg_rca32_csa21_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[41] = u_CSAwallace_pg_rca32_csa21_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[42] = u_CSAwallace_pg_rca32_csa21_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[43] = u_CSAwallace_pg_rca32_csa21_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[44] = u_CSAwallace_pg_rca32_csa21_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[45] = u_CSAwallace_pg_rca32_csa21_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[46] = u_CSAwallace_pg_rca32_csa21_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[47] = u_CSAwallace_pg_rca32_csa21_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[48] = u_CSAwallace_pg_rca32_csa21_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[49] = u_CSAwallace_pg_rca32_csa21_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[50] = u_CSAwallace_pg_rca32_csa21_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[51] = u_CSAwallace_pg_rca32_csa21_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[52] = u_CSAwallace_pg_rca32_csa21_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[53] = u_CSAwallace_pg_rca32_csa21_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[54] = u_CSAwallace_pg_rca32_csa21_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[55] = u_CSAwallace_pg_rca32_csa21_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[56] = u_CSAwallace_pg_rca32_csa21_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[57] = u_CSAwallace_pg_rca32_csa21_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[58] = u_CSAwallace_pg_rca32_csa21_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[59] = u_CSAwallace_pg_rca32_csa21_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[60] = u_CSAwallace_pg_rca32_csa21_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[61] = u_CSAwallace_pg_rca32_csa21_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[62] = u_CSAwallace_pg_rca32_csa21_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22[63] = 1'b0;
  csa_component64 csa_component64_u_CSAwallace_pg_rca32_csa24_csa_component_out(.a(u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s21), .b(u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_c21), .c(u_CSAwallace_pg_rca32_csa24_csa_component_u_CSAwallace_pg_rca32_csa_s22), .csa_component64_out(u_CSAwallace_pg_rca32_csa24_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[0] = u_CSAwallace_pg_rca32_csa22_csa_component_out[0];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[1] = u_CSAwallace_pg_rca32_csa22_csa_component_out[1];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[2] = u_CSAwallace_pg_rca32_csa22_csa_component_out[2];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[3] = u_CSAwallace_pg_rca32_csa22_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[4] = u_CSAwallace_pg_rca32_csa22_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[5] = u_CSAwallace_pg_rca32_csa22_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[6] = u_CSAwallace_pg_rca32_csa22_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[7] = u_CSAwallace_pg_rca32_csa22_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[8] = u_CSAwallace_pg_rca32_csa22_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[9] = u_CSAwallace_pg_rca32_csa22_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[10] = u_CSAwallace_pg_rca32_csa22_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[11] = u_CSAwallace_pg_rca32_csa22_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[12] = u_CSAwallace_pg_rca32_csa22_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[13] = u_CSAwallace_pg_rca32_csa22_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[14] = u_CSAwallace_pg_rca32_csa22_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[15] = u_CSAwallace_pg_rca32_csa22_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[16] = u_CSAwallace_pg_rca32_csa22_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[17] = u_CSAwallace_pg_rca32_csa22_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[18] = u_CSAwallace_pg_rca32_csa22_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[19] = u_CSAwallace_pg_rca32_csa22_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[20] = u_CSAwallace_pg_rca32_csa22_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[21] = u_CSAwallace_pg_rca32_csa22_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[22] = u_CSAwallace_pg_rca32_csa22_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[23] = u_CSAwallace_pg_rca32_csa22_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[24] = u_CSAwallace_pg_rca32_csa22_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[25] = u_CSAwallace_pg_rca32_csa22_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[26] = u_CSAwallace_pg_rca32_csa22_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[27] = u_CSAwallace_pg_rca32_csa22_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[28] = u_CSAwallace_pg_rca32_csa22_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[29] = u_CSAwallace_pg_rca32_csa22_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[30] = u_CSAwallace_pg_rca32_csa22_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[31] = u_CSAwallace_pg_rca32_csa22_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[32] = u_CSAwallace_pg_rca32_csa22_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[33] = u_CSAwallace_pg_rca32_csa22_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[34] = u_CSAwallace_pg_rca32_csa22_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[35] = u_CSAwallace_pg_rca32_csa22_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[36] = u_CSAwallace_pg_rca32_csa22_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[37] = u_CSAwallace_pg_rca32_csa22_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[38] = u_CSAwallace_pg_rca32_csa22_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[39] = u_CSAwallace_pg_rca32_csa22_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[40] = u_CSAwallace_pg_rca32_csa22_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[41] = u_CSAwallace_pg_rca32_csa22_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[42] = u_CSAwallace_pg_rca32_csa22_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[43] = u_CSAwallace_pg_rca32_csa22_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[44] = u_CSAwallace_pg_rca32_csa22_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[45] = u_CSAwallace_pg_rca32_csa22_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[49] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[50] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[5] = u_CSAwallace_pg_rca32_csa22_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[6] = u_CSAwallace_pg_rca32_csa22_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[7] = u_CSAwallace_pg_rca32_csa22_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[8] = u_CSAwallace_pg_rca32_csa22_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[9] = u_CSAwallace_pg_rca32_csa22_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[10] = u_CSAwallace_pg_rca32_csa22_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[11] = u_CSAwallace_pg_rca32_csa22_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[12] = u_CSAwallace_pg_rca32_csa22_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[13] = u_CSAwallace_pg_rca32_csa22_csa_component_out[63];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[14] = u_CSAwallace_pg_rca32_csa22_csa_component_out[64];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[15] = u_CSAwallace_pg_rca32_csa22_csa_component_out[65];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[16] = u_CSAwallace_pg_rca32_csa22_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[17] = u_CSAwallace_pg_rca32_csa22_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[18] = u_CSAwallace_pg_rca32_csa22_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[19] = u_CSAwallace_pg_rca32_csa22_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[20] = u_CSAwallace_pg_rca32_csa22_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[21] = u_CSAwallace_pg_rca32_csa22_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[22] = u_CSAwallace_pg_rca32_csa22_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[23] = u_CSAwallace_pg_rca32_csa22_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[24] = u_CSAwallace_pg_rca32_csa22_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[25] = u_CSAwallace_pg_rca32_csa22_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[26] = u_CSAwallace_pg_rca32_csa22_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[27] = u_CSAwallace_pg_rca32_csa22_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[28] = u_CSAwallace_pg_rca32_csa22_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[29] = u_CSAwallace_pg_rca32_csa22_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[30] = u_CSAwallace_pg_rca32_csa22_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[31] = u_CSAwallace_pg_rca32_csa22_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[32] = u_CSAwallace_pg_rca32_csa22_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[33] = u_CSAwallace_pg_rca32_csa22_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[34] = u_CSAwallace_pg_rca32_csa22_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[35] = u_CSAwallace_pg_rca32_csa22_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[36] = u_CSAwallace_pg_rca32_csa22_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[37] = u_CSAwallace_pg_rca32_csa22_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[38] = u_CSAwallace_pg_rca32_csa22_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[39] = u_CSAwallace_pg_rca32_csa22_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[40] = u_CSAwallace_pg_rca32_csa22_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[41] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[42] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[43] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[44] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[45] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[46] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[49] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[50] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[10] = u_CSAwallace_pg_rca32_csa23_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[11] = u_CSAwallace_pg_rca32_csa23_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[12] = u_CSAwallace_pg_rca32_csa23_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[13] = u_CSAwallace_pg_rca32_csa23_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[14] = u_CSAwallace_pg_rca32_csa23_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[15] = u_CSAwallace_pg_rca32_csa23_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[16] = u_CSAwallace_pg_rca32_csa23_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[17] = u_CSAwallace_pg_rca32_csa23_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[18] = u_CSAwallace_pg_rca32_csa23_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[19] = u_CSAwallace_pg_rca32_csa23_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[20] = u_CSAwallace_pg_rca32_csa23_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[21] = u_CSAwallace_pg_rca32_csa23_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[22] = u_CSAwallace_pg_rca32_csa23_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[23] = u_CSAwallace_pg_rca32_csa23_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[24] = u_CSAwallace_pg_rca32_csa23_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[25] = u_CSAwallace_pg_rca32_csa23_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[26] = u_CSAwallace_pg_rca32_csa23_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[27] = u_CSAwallace_pg_rca32_csa23_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[28] = u_CSAwallace_pg_rca32_csa23_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[29] = u_CSAwallace_pg_rca32_csa23_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[30] = u_CSAwallace_pg_rca32_csa23_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[31] = u_CSAwallace_pg_rca32_csa23_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[32] = u_CSAwallace_pg_rca32_csa23_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[33] = u_CSAwallace_pg_rca32_csa23_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[34] = u_CSAwallace_pg_rca32_csa23_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[35] = u_CSAwallace_pg_rca32_csa23_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[36] = u_CSAwallace_pg_rca32_csa23_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[37] = u_CSAwallace_pg_rca32_csa23_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[38] = u_CSAwallace_pg_rca32_csa23_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[39] = u_CSAwallace_pg_rca32_csa23_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[40] = u_CSAwallace_pg_rca32_csa23_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[41] = u_CSAwallace_pg_rca32_csa23_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[42] = u_CSAwallace_pg_rca32_csa23_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[43] = u_CSAwallace_pg_rca32_csa23_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[44] = u_CSAwallace_pg_rca32_csa23_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[45] = u_CSAwallace_pg_rca32_csa23_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[46] = u_CSAwallace_pg_rca32_csa23_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[47] = u_CSAwallace_pg_rca32_csa23_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[48] = u_CSAwallace_pg_rca32_csa23_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[49] = u_CSAwallace_pg_rca32_csa23_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[50] = u_CSAwallace_pg_rca32_csa23_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[51] = u_CSAwallace_pg_rca32_csa23_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[52] = u_CSAwallace_pg_rca32_csa23_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[53] = u_CSAwallace_pg_rca32_csa23_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[54] = u_CSAwallace_pg_rca32_csa23_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24[58] = 1'b0;
  csa_component59 csa_component59_u_CSAwallace_pg_rca32_csa25_csa_component_out(.a(u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s23), .b(u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_c23), .c(u_CSAwallace_pg_rca32_csa25_csa_component_u_CSAwallace_pg_rca32_csa_s24), .csa_component59_out(u_CSAwallace_pg_rca32_csa25_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[15] = u_CSAwallace_pg_rca32_csa23_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[16] = u_CSAwallace_pg_rca32_csa23_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[17] = u_CSAwallace_pg_rca32_csa23_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[18] = u_CSAwallace_pg_rca32_csa23_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[19] = u_CSAwallace_pg_rca32_csa23_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[20] = u_CSAwallace_pg_rca32_csa23_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[21] = u_CSAwallace_pg_rca32_csa23_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[22] = u_CSAwallace_pg_rca32_csa23_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[23] = u_CSAwallace_pg_rca32_csa23_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[24] = u_CSAwallace_pg_rca32_csa23_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[25] = u_CSAwallace_pg_rca32_csa23_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[26] = u_CSAwallace_pg_rca32_csa23_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[27] = u_CSAwallace_pg_rca32_csa23_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[28] = u_CSAwallace_pg_rca32_csa23_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[29] = u_CSAwallace_pg_rca32_csa23_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[30] = u_CSAwallace_pg_rca32_csa23_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[31] = u_CSAwallace_pg_rca32_csa23_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[32] = u_CSAwallace_pg_rca32_csa23_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[33] = u_CSAwallace_pg_rca32_csa23_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[34] = u_CSAwallace_pg_rca32_csa23_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[35] = u_CSAwallace_pg_rca32_csa23_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[36] = u_CSAwallace_pg_rca32_csa23_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[37] = u_CSAwallace_pg_rca32_csa23_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[38] = u_CSAwallace_pg_rca32_csa23_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[39] = u_CSAwallace_pg_rca32_csa23_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[40] = u_CSAwallace_pg_rca32_csa23_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[41] = u_CSAwallace_pg_rca32_csa23_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[42] = u_CSAwallace_pg_rca32_csa23_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[43] = u_CSAwallace_pg_rca32_csa23_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[44] = u_CSAwallace_pg_rca32_csa23_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[45] = u_CSAwallace_pg_rca32_csa23_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[46] = u_CSAwallace_pg_rca32_csa23_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[47] = u_CSAwallace_pg_rca32_csa23_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[48] = u_CSAwallace_pg_rca32_csa23_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[49] = u_CSAwallace_pg_rca32_csa23_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[50] = u_CSAwallace_pg_rca32_csa23_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[51] = u_CSAwallace_pg_rca32_csa23_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[21] = u_CSAwallace_pg_rca32_csa24_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[22] = u_CSAwallace_pg_rca32_csa24_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[23] = u_CSAwallace_pg_rca32_csa24_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[24] = u_CSAwallace_pg_rca32_csa24_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[25] = u_CSAwallace_pg_rca32_csa24_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[26] = u_CSAwallace_pg_rca32_csa24_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[27] = u_CSAwallace_pg_rca32_csa24_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[28] = u_CSAwallace_pg_rca32_csa24_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[29] = u_CSAwallace_pg_rca32_csa24_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[30] = u_CSAwallace_pg_rca32_csa24_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[31] = u_CSAwallace_pg_rca32_csa24_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[32] = u_CSAwallace_pg_rca32_csa24_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[33] = u_CSAwallace_pg_rca32_csa24_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[34] = u_CSAwallace_pg_rca32_csa24_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[35] = u_CSAwallace_pg_rca32_csa24_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[36] = u_CSAwallace_pg_rca32_csa24_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[37] = u_CSAwallace_pg_rca32_csa24_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[38] = u_CSAwallace_pg_rca32_csa24_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[39] = u_CSAwallace_pg_rca32_csa24_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[40] = u_CSAwallace_pg_rca32_csa24_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[41] = u_CSAwallace_pg_rca32_csa24_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[42] = u_CSAwallace_pg_rca32_csa24_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[43] = u_CSAwallace_pg_rca32_csa24_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[44] = u_CSAwallace_pg_rca32_csa24_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[45] = u_CSAwallace_pg_rca32_csa24_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[46] = u_CSAwallace_pg_rca32_csa24_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[47] = u_CSAwallace_pg_rca32_csa24_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[48] = u_CSAwallace_pg_rca32_csa24_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[49] = u_CSAwallace_pg_rca32_csa24_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[50] = u_CSAwallace_pg_rca32_csa24_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[51] = u_CSAwallace_pg_rca32_csa24_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[52] = u_CSAwallace_pg_rca32_csa24_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[53] = u_CSAwallace_pg_rca32_csa24_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[54] = u_CSAwallace_pg_rca32_csa24_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[55] = u_CSAwallace_pg_rca32_csa24_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[56] = u_CSAwallace_pg_rca32_csa24_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[57] = u_CSAwallace_pg_rca32_csa24_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[58] = u_CSAwallace_pg_rca32_csa24_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[59] = u_CSAwallace_pg_rca32_csa24_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[60] = u_CSAwallace_pg_rca32_csa24_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[61] = u_CSAwallace_pg_rca32_csa24_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[62] = u_CSAwallace_pg_rca32_csa24_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[25] = u_CSAwallace_pg_rca32_csa24_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[26] = u_CSAwallace_pg_rca32_csa24_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[27] = u_CSAwallace_pg_rca32_csa24_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[28] = u_CSAwallace_pg_rca32_csa24_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[29] = u_CSAwallace_pg_rca32_csa24_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[30] = u_CSAwallace_pg_rca32_csa24_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[31] = u_CSAwallace_pg_rca32_csa24_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[32] = u_CSAwallace_pg_rca32_csa24_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[33] = u_CSAwallace_pg_rca32_csa24_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[34] = u_CSAwallace_pg_rca32_csa24_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[35] = u_CSAwallace_pg_rca32_csa24_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[36] = u_CSAwallace_pg_rca32_csa24_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[37] = u_CSAwallace_pg_rca32_csa24_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[38] = u_CSAwallace_pg_rca32_csa24_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[39] = u_CSAwallace_pg_rca32_csa24_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[40] = u_CSAwallace_pg_rca32_csa24_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[41] = u_CSAwallace_pg_rca32_csa24_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[42] = u_CSAwallace_pg_rca32_csa24_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[43] = u_CSAwallace_pg_rca32_csa24_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[44] = u_CSAwallace_pg_rca32_csa24_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[45] = u_CSAwallace_pg_rca32_csa24_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[46] = u_CSAwallace_pg_rca32_csa24_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[47] = u_CSAwallace_pg_rca32_csa24_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[48] = u_CSAwallace_pg_rca32_csa24_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[49] = u_CSAwallace_pg_rca32_csa24_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[50] = u_CSAwallace_pg_rca32_csa24_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[51] = u_CSAwallace_pg_rca32_csa24_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[52] = u_CSAwallace_pg_rca32_csa24_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[53] = u_CSAwallace_pg_rca32_csa24_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[54] = u_CSAwallace_pg_rca32_csa24_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[55] = u_CSAwallace_pg_rca32_csa24_csa_component_out[120];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[56] = u_CSAwallace_pg_rca32_csa24_csa_component_out[121];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[57] = u_CSAwallace_pg_rca32_csa24_csa_component_out[122];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[58] = u_CSAwallace_pg_rca32_csa24_csa_component_out[123];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[59] = u_CSAwallace_pg_rca32_csa24_csa_component_out[124];
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25[63] = 1'b0;
  csa_component64 csa_component64_u_CSAwallace_pg_rca32_csa26_csa_component_out(.a(u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c24), .b(u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_s25), .c(u_CSAwallace_pg_rca32_csa26_csa_component_u_CSAwallace_pg_rca32_csa_c25), .csa_component64_out(u_CSAwallace_pg_rca32_csa26_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[0] = u_CSAwallace_pg_rca32_csa25_csa_component_out[0];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[1] = u_CSAwallace_pg_rca32_csa25_csa_component_out[1];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[2] = u_CSAwallace_pg_rca32_csa25_csa_component_out[2];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[3] = u_CSAwallace_pg_rca32_csa25_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[4] = u_CSAwallace_pg_rca32_csa25_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[5] = u_CSAwallace_pg_rca32_csa25_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[6] = u_CSAwallace_pg_rca32_csa25_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[7] = u_CSAwallace_pg_rca32_csa25_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[8] = u_CSAwallace_pg_rca32_csa25_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[9] = u_CSAwallace_pg_rca32_csa25_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[10] = u_CSAwallace_pg_rca32_csa25_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[11] = u_CSAwallace_pg_rca32_csa25_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[12] = u_CSAwallace_pg_rca32_csa25_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[13] = u_CSAwallace_pg_rca32_csa25_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[14] = u_CSAwallace_pg_rca32_csa25_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[15] = u_CSAwallace_pg_rca32_csa25_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[16] = u_CSAwallace_pg_rca32_csa25_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[17] = u_CSAwallace_pg_rca32_csa25_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[18] = u_CSAwallace_pg_rca32_csa25_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[19] = u_CSAwallace_pg_rca32_csa25_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[20] = u_CSAwallace_pg_rca32_csa25_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[21] = u_CSAwallace_pg_rca32_csa25_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[22] = u_CSAwallace_pg_rca32_csa25_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[23] = u_CSAwallace_pg_rca32_csa25_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[24] = u_CSAwallace_pg_rca32_csa25_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[25] = u_CSAwallace_pg_rca32_csa25_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[26] = u_CSAwallace_pg_rca32_csa25_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[27] = u_CSAwallace_pg_rca32_csa25_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[28] = u_CSAwallace_pg_rca32_csa25_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[29] = u_CSAwallace_pg_rca32_csa25_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[30] = u_CSAwallace_pg_rca32_csa25_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[31] = u_CSAwallace_pg_rca32_csa25_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[32] = u_CSAwallace_pg_rca32_csa25_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[33] = u_CSAwallace_pg_rca32_csa25_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[34] = u_CSAwallace_pg_rca32_csa25_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[35] = u_CSAwallace_pg_rca32_csa25_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[36] = u_CSAwallace_pg_rca32_csa25_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[37] = u_CSAwallace_pg_rca32_csa25_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[38] = u_CSAwallace_pg_rca32_csa25_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[39] = u_CSAwallace_pg_rca32_csa25_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[40] = u_CSAwallace_pg_rca32_csa25_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[41] = u_CSAwallace_pg_rca32_csa25_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[42] = u_CSAwallace_pg_rca32_csa25_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[43] = u_CSAwallace_pg_rca32_csa25_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[44] = u_CSAwallace_pg_rca32_csa25_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[45] = u_CSAwallace_pg_rca32_csa25_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[46] = u_CSAwallace_pg_rca32_csa25_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[47] = u_CSAwallace_pg_rca32_csa25_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[48] = u_CSAwallace_pg_rca32_csa25_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[49] = u_CSAwallace_pg_rca32_csa25_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[50] = u_CSAwallace_pg_rca32_csa25_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[51] = u_CSAwallace_pg_rca32_csa25_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[52] = u_CSAwallace_pg_rca32_csa25_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[53] = u_CSAwallace_pg_rca32_csa25_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[54] = u_CSAwallace_pg_rca32_csa25_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[6] = u_CSAwallace_pg_rca32_csa25_csa_component_out[66];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[7] = u_CSAwallace_pg_rca32_csa25_csa_component_out[67];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[8] = u_CSAwallace_pg_rca32_csa25_csa_component_out[68];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[9] = u_CSAwallace_pg_rca32_csa25_csa_component_out[69];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[10] = u_CSAwallace_pg_rca32_csa25_csa_component_out[70];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[11] = u_CSAwallace_pg_rca32_csa25_csa_component_out[71];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[12] = u_CSAwallace_pg_rca32_csa25_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[13] = u_CSAwallace_pg_rca32_csa25_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[14] = u_CSAwallace_pg_rca32_csa25_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[15] = u_CSAwallace_pg_rca32_csa25_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[16] = u_CSAwallace_pg_rca32_csa25_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[17] = u_CSAwallace_pg_rca32_csa25_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[18] = u_CSAwallace_pg_rca32_csa25_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[19] = u_CSAwallace_pg_rca32_csa25_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[20] = u_CSAwallace_pg_rca32_csa25_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[21] = u_CSAwallace_pg_rca32_csa25_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[22] = u_CSAwallace_pg_rca32_csa25_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[23] = u_CSAwallace_pg_rca32_csa25_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[24] = u_CSAwallace_pg_rca32_csa25_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[25] = u_CSAwallace_pg_rca32_csa25_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[26] = u_CSAwallace_pg_rca32_csa25_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[27] = u_CSAwallace_pg_rca32_csa25_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[28] = u_CSAwallace_pg_rca32_csa25_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[29] = u_CSAwallace_pg_rca32_csa25_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[30] = u_CSAwallace_pg_rca32_csa25_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[31] = u_CSAwallace_pg_rca32_csa25_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[32] = u_CSAwallace_pg_rca32_csa25_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[33] = u_CSAwallace_pg_rca32_csa25_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[34] = u_CSAwallace_pg_rca32_csa25_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[35] = u_CSAwallace_pg_rca32_csa25_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[36] = u_CSAwallace_pg_rca32_csa25_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[37] = u_CSAwallace_pg_rca32_csa25_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[38] = u_CSAwallace_pg_rca32_csa25_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[39] = u_CSAwallace_pg_rca32_csa25_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[40] = u_CSAwallace_pg_rca32_csa25_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[41] = u_CSAwallace_pg_rca32_csa25_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[42] = u_CSAwallace_pg_rca32_csa25_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[43] = u_CSAwallace_pg_rca32_csa25_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[44] = u_CSAwallace_pg_rca32_csa25_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[45] = u_CSAwallace_pg_rca32_csa25_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[46] = u_CSAwallace_pg_rca32_csa25_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[47] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[48] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[49] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[50] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[51] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[52] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[53] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[54] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[55] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[15] = u_CSAwallace_pg_rca32_csa26_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[16] = u_CSAwallace_pg_rca32_csa26_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[17] = u_CSAwallace_pg_rca32_csa26_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[18] = u_CSAwallace_pg_rca32_csa26_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[19] = u_CSAwallace_pg_rca32_csa26_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[20] = u_CSAwallace_pg_rca32_csa26_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[21] = u_CSAwallace_pg_rca32_csa26_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[22] = u_CSAwallace_pg_rca32_csa26_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[23] = u_CSAwallace_pg_rca32_csa26_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[24] = u_CSAwallace_pg_rca32_csa26_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[25] = u_CSAwallace_pg_rca32_csa26_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[26] = u_CSAwallace_pg_rca32_csa26_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[27] = u_CSAwallace_pg_rca32_csa26_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[28] = u_CSAwallace_pg_rca32_csa26_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[29] = u_CSAwallace_pg_rca32_csa26_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[30] = u_CSAwallace_pg_rca32_csa26_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[31] = u_CSAwallace_pg_rca32_csa26_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[32] = u_CSAwallace_pg_rca32_csa26_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[33] = u_CSAwallace_pg_rca32_csa26_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[34] = u_CSAwallace_pg_rca32_csa26_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[35] = u_CSAwallace_pg_rca32_csa26_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[36] = u_CSAwallace_pg_rca32_csa26_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[37] = u_CSAwallace_pg_rca32_csa26_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[38] = u_CSAwallace_pg_rca32_csa26_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[39] = u_CSAwallace_pg_rca32_csa26_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[40] = u_CSAwallace_pg_rca32_csa26_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[41] = u_CSAwallace_pg_rca32_csa26_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[42] = u_CSAwallace_pg_rca32_csa26_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[43] = u_CSAwallace_pg_rca32_csa26_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[44] = u_CSAwallace_pg_rca32_csa26_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[45] = u_CSAwallace_pg_rca32_csa26_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[46] = u_CSAwallace_pg_rca32_csa26_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[47] = u_CSAwallace_pg_rca32_csa26_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[48] = u_CSAwallace_pg_rca32_csa26_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[49] = u_CSAwallace_pg_rca32_csa26_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[50] = u_CSAwallace_pg_rca32_csa26_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[51] = u_CSAwallace_pg_rca32_csa26_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[52] = u_CSAwallace_pg_rca32_csa26_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[53] = u_CSAwallace_pg_rca32_csa26_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[54] = u_CSAwallace_pg_rca32_csa26_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[55] = u_CSAwallace_pg_rca32_csa26_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[56] = u_CSAwallace_pg_rca32_csa26_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[57] = u_CSAwallace_pg_rca32_csa26_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[58] = u_CSAwallace_pg_rca32_csa26_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[59] = u_CSAwallace_pg_rca32_csa26_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[60] = u_CSAwallace_pg_rca32_csa26_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[61] = u_CSAwallace_pg_rca32_csa26_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[62] = u_CSAwallace_pg_rca32_csa26_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27[63] = 1'b0;
  csa_component64 csa_component64_u_CSAwallace_pg_rca32_csa27_csa_component_out(.a(u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s26), .b(u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_c26), .c(u_CSAwallace_pg_rca32_csa27_csa_component_u_CSAwallace_pg_rca32_csa_s27), .csa_component64_out(u_CSAwallace_pg_rca32_csa27_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[0] = u_CSAwallace_pg_rca32_csa27_csa_component_out[0];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[1] = u_CSAwallace_pg_rca32_csa27_csa_component_out[1];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[2] = u_CSAwallace_pg_rca32_csa27_csa_component_out[2];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[3] = u_CSAwallace_pg_rca32_csa27_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[4] = u_CSAwallace_pg_rca32_csa27_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[5] = u_CSAwallace_pg_rca32_csa27_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[6] = u_CSAwallace_pg_rca32_csa27_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[7] = u_CSAwallace_pg_rca32_csa27_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[8] = u_CSAwallace_pg_rca32_csa27_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[9] = u_CSAwallace_pg_rca32_csa27_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[10] = u_CSAwallace_pg_rca32_csa27_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[11] = u_CSAwallace_pg_rca32_csa27_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[12] = u_CSAwallace_pg_rca32_csa27_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[13] = u_CSAwallace_pg_rca32_csa27_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[14] = u_CSAwallace_pg_rca32_csa27_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[15] = u_CSAwallace_pg_rca32_csa27_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[16] = u_CSAwallace_pg_rca32_csa27_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[17] = u_CSAwallace_pg_rca32_csa27_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[18] = u_CSAwallace_pg_rca32_csa27_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[19] = u_CSAwallace_pg_rca32_csa27_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[20] = u_CSAwallace_pg_rca32_csa27_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[21] = u_CSAwallace_pg_rca32_csa27_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[22] = u_CSAwallace_pg_rca32_csa27_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[23] = u_CSAwallace_pg_rca32_csa27_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[24] = u_CSAwallace_pg_rca32_csa27_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[25] = u_CSAwallace_pg_rca32_csa27_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[26] = u_CSAwallace_pg_rca32_csa27_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[27] = u_CSAwallace_pg_rca32_csa27_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[28] = u_CSAwallace_pg_rca32_csa27_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[29] = u_CSAwallace_pg_rca32_csa27_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[30] = u_CSAwallace_pg_rca32_csa27_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[31] = u_CSAwallace_pg_rca32_csa27_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[32] = u_CSAwallace_pg_rca32_csa27_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[33] = u_CSAwallace_pg_rca32_csa27_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[34] = u_CSAwallace_pg_rca32_csa27_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[35] = u_CSAwallace_pg_rca32_csa27_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[36] = u_CSAwallace_pg_rca32_csa27_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[37] = u_CSAwallace_pg_rca32_csa27_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[38] = u_CSAwallace_pg_rca32_csa27_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[39] = u_CSAwallace_pg_rca32_csa27_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[40] = u_CSAwallace_pg_rca32_csa27_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[41] = u_CSAwallace_pg_rca32_csa27_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[42] = u_CSAwallace_pg_rca32_csa27_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[43] = u_CSAwallace_pg_rca32_csa27_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[44] = u_CSAwallace_pg_rca32_csa27_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[45] = u_CSAwallace_pg_rca32_csa27_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[46] = u_CSAwallace_pg_rca32_csa27_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[47] = u_CSAwallace_pg_rca32_csa27_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[48] = u_CSAwallace_pg_rca32_csa27_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[49] = u_CSAwallace_pg_rca32_csa27_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[50] = u_CSAwallace_pg_rca32_csa27_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[51] = u_CSAwallace_pg_rca32_csa27_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[52] = u_CSAwallace_pg_rca32_csa27_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[53] = u_CSAwallace_pg_rca32_csa27_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[54] = u_CSAwallace_pg_rca32_csa27_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[55] = u_CSAwallace_pg_rca32_csa27_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[56] = u_CSAwallace_pg_rca32_csa27_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[57] = u_CSAwallace_pg_rca32_csa27_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[58] = u_CSAwallace_pg_rca32_csa27_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[59] = u_CSAwallace_pg_rca32_csa27_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[60] = u_CSAwallace_pg_rca32_csa27_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[61] = u_CSAwallace_pg_rca32_csa27_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[62] = u_CSAwallace_pg_rca32_csa27_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[7] = u_CSAwallace_pg_rca32_csa27_csa_component_out[72];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[8] = u_CSAwallace_pg_rca32_csa27_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[9] = u_CSAwallace_pg_rca32_csa27_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[10] = u_CSAwallace_pg_rca32_csa27_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[11] = u_CSAwallace_pg_rca32_csa27_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[12] = u_CSAwallace_pg_rca32_csa27_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[13] = u_CSAwallace_pg_rca32_csa27_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[14] = u_CSAwallace_pg_rca32_csa27_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[15] = u_CSAwallace_pg_rca32_csa27_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[16] = u_CSAwallace_pg_rca32_csa27_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[17] = u_CSAwallace_pg_rca32_csa27_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[18] = u_CSAwallace_pg_rca32_csa27_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[19] = u_CSAwallace_pg_rca32_csa27_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[20] = u_CSAwallace_pg_rca32_csa27_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[21] = u_CSAwallace_pg_rca32_csa27_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[22] = u_CSAwallace_pg_rca32_csa27_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[23] = u_CSAwallace_pg_rca32_csa27_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[24] = u_CSAwallace_pg_rca32_csa27_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[25] = u_CSAwallace_pg_rca32_csa27_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[26] = u_CSAwallace_pg_rca32_csa27_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[27] = u_CSAwallace_pg_rca32_csa27_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[28] = u_CSAwallace_pg_rca32_csa27_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[29] = u_CSAwallace_pg_rca32_csa27_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[30] = u_CSAwallace_pg_rca32_csa27_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[31] = u_CSAwallace_pg_rca32_csa27_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[32] = u_CSAwallace_pg_rca32_csa27_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[33] = u_CSAwallace_pg_rca32_csa27_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[34] = u_CSAwallace_pg_rca32_csa27_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[35] = u_CSAwallace_pg_rca32_csa27_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[36] = u_CSAwallace_pg_rca32_csa27_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[37] = u_CSAwallace_pg_rca32_csa27_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[38] = u_CSAwallace_pg_rca32_csa27_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[39] = u_CSAwallace_pg_rca32_csa27_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[40] = u_CSAwallace_pg_rca32_csa27_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[41] = u_CSAwallace_pg_rca32_csa27_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[42] = u_CSAwallace_pg_rca32_csa27_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[43] = u_CSAwallace_pg_rca32_csa27_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[44] = u_CSAwallace_pg_rca32_csa27_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[45] = u_CSAwallace_pg_rca32_csa27_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[46] = u_CSAwallace_pg_rca32_csa27_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[47] = u_CSAwallace_pg_rca32_csa27_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[48] = u_CSAwallace_pg_rca32_csa27_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[49] = u_CSAwallace_pg_rca32_csa27_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[50] = u_CSAwallace_pg_rca32_csa27_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[51] = u_CSAwallace_pg_rca32_csa27_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[52] = u_CSAwallace_pg_rca32_csa27_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[53] = u_CSAwallace_pg_rca32_csa27_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[54] = u_CSAwallace_pg_rca32_csa27_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[55] = u_CSAwallace_pg_rca32_csa27_csa_component_out[120];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[56] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[57] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[58] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[59] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[60] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[22] = u_CSAwallace_pg_rca32_csa26_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[23] = u_CSAwallace_pg_rca32_csa26_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[24] = u_CSAwallace_pg_rca32_csa26_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[25] = u_CSAwallace_pg_rca32_csa26_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[26] = u_CSAwallace_pg_rca32_csa26_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[27] = u_CSAwallace_pg_rca32_csa26_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[28] = u_CSAwallace_pg_rca32_csa26_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[29] = u_CSAwallace_pg_rca32_csa26_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[30] = u_CSAwallace_pg_rca32_csa26_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[31] = u_CSAwallace_pg_rca32_csa26_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[32] = u_CSAwallace_pg_rca32_csa26_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[33] = u_CSAwallace_pg_rca32_csa26_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[34] = u_CSAwallace_pg_rca32_csa26_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[35] = u_CSAwallace_pg_rca32_csa26_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[36] = u_CSAwallace_pg_rca32_csa26_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[37] = u_CSAwallace_pg_rca32_csa26_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[38] = u_CSAwallace_pg_rca32_csa26_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[39] = u_CSAwallace_pg_rca32_csa26_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[40] = u_CSAwallace_pg_rca32_csa26_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[41] = u_CSAwallace_pg_rca32_csa26_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[42] = u_CSAwallace_pg_rca32_csa26_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[43] = u_CSAwallace_pg_rca32_csa26_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[44] = u_CSAwallace_pg_rca32_csa26_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[45] = u_CSAwallace_pg_rca32_csa26_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[46] = u_CSAwallace_pg_rca32_csa26_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[47] = u_CSAwallace_pg_rca32_csa26_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[48] = u_CSAwallace_pg_rca32_csa26_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[49] = u_CSAwallace_pg_rca32_csa26_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[50] = u_CSAwallace_pg_rca32_csa26_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[51] = u_CSAwallace_pg_rca32_csa26_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[52] = u_CSAwallace_pg_rca32_csa26_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[53] = u_CSAwallace_pg_rca32_csa26_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[54] = u_CSAwallace_pg_rca32_csa26_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[55] = u_CSAwallace_pg_rca32_csa26_csa_component_out[120];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[56] = u_CSAwallace_pg_rca32_csa26_csa_component_out[121];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[57] = u_CSAwallace_pg_rca32_csa26_csa_component_out[122];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[58] = u_CSAwallace_pg_rca32_csa26_csa_component_out[123];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[59] = u_CSAwallace_pg_rca32_csa26_csa_component_out[124];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[60] = u_CSAwallace_pg_rca32_csa26_csa_component_out[125];
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[61] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27[63] = 1'b0;
  csa_component64 csa_component64_u_CSAwallace_pg_rca32_csa28_csa_component_out(.a(u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_s28), .b(u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c28), .c(u_CSAwallace_pg_rca32_csa28_csa_component_u_CSAwallace_pg_rca32_csa_c27), .csa_component64_out(u_CSAwallace_pg_rca32_csa28_csa_component_out));
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[0] = u_CSAwallace_pg_rca32_csa28_csa_component_out[0];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[1] = u_CSAwallace_pg_rca32_csa28_csa_component_out[1];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[2] = u_CSAwallace_pg_rca32_csa28_csa_component_out[2];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[3] = u_CSAwallace_pg_rca32_csa28_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[4] = u_CSAwallace_pg_rca32_csa28_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[5] = u_CSAwallace_pg_rca32_csa28_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[6] = u_CSAwallace_pg_rca32_csa28_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[7] = u_CSAwallace_pg_rca32_csa28_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[8] = u_CSAwallace_pg_rca32_csa28_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[9] = u_CSAwallace_pg_rca32_csa28_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[10] = u_CSAwallace_pg_rca32_csa28_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[11] = u_CSAwallace_pg_rca32_csa28_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[12] = u_CSAwallace_pg_rca32_csa28_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[13] = u_CSAwallace_pg_rca32_csa28_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[14] = u_CSAwallace_pg_rca32_csa28_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[15] = u_CSAwallace_pg_rca32_csa28_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[16] = u_CSAwallace_pg_rca32_csa28_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[17] = u_CSAwallace_pg_rca32_csa28_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[18] = u_CSAwallace_pg_rca32_csa28_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[19] = u_CSAwallace_pg_rca32_csa28_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[20] = u_CSAwallace_pg_rca32_csa28_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[21] = u_CSAwallace_pg_rca32_csa28_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[22] = u_CSAwallace_pg_rca32_csa28_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[23] = u_CSAwallace_pg_rca32_csa28_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[24] = u_CSAwallace_pg_rca32_csa28_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[25] = u_CSAwallace_pg_rca32_csa28_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[26] = u_CSAwallace_pg_rca32_csa28_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[27] = u_CSAwallace_pg_rca32_csa28_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[28] = u_CSAwallace_pg_rca32_csa28_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[29] = u_CSAwallace_pg_rca32_csa28_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[30] = u_CSAwallace_pg_rca32_csa28_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[31] = u_CSAwallace_pg_rca32_csa28_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[32] = u_CSAwallace_pg_rca32_csa28_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[33] = u_CSAwallace_pg_rca32_csa28_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[34] = u_CSAwallace_pg_rca32_csa28_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[35] = u_CSAwallace_pg_rca32_csa28_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[36] = u_CSAwallace_pg_rca32_csa28_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[37] = u_CSAwallace_pg_rca32_csa28_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[38] = u_CSAwallace_pg_rca32_csa28_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[39] = u_CSAwallace_pg_rca32_csa28_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[40] = u_CSAwallace_pg_rca32_csa28_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[41] = u_CSAwallace_pg_rca32_csa28_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[42] = u_CSAwallace_pg_rca32_csa28_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[43] = u_CSAwallace_pg_rca32_csa28_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[44] = u_CSAwallace_pg_rca32_csa28_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[45] = u_CSAwallace_pg_rca32_csa28_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[46] = u_CSAwallace_pg_rca32_csa28_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[47] = u_CSAwallace_pg_rca32_csa28_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[48] = u_CSAwallace_pg_rca32_csa28_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[49] = u_CSAwallace_pg_rca32_csa28_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[50] = u_CSAwallace_pg_rca32_csa28_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[51] = u_CSAwallace_pg_rca32_csa28_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[52] = u_CSAwallace_pg_rca32_csa28_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[53] = u_CSAwallace_pg_rca32_csa28_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[54] = u_CSAwallace_pg_rca32_csa28_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[55] = u_CSAwallace_pg_rca32_csa28_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[56] = u_CSAwallace_pg_rca32_csa28_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[57] = u_CSAwallace_pg_rca32_csa28_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[58] = u_CSAwallace_pg_rca32_csa28_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[59] = u_CSAwallace_pg_rca32_csa28_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[60] = u_CSAwallace_pg_rca32_csa28_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[61] = u_CSAwallace_pg_rca32_csa28_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[62] = u_CSAwallace_pg_rca32_csa28_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[8] = u_CSAwallace_pg_rca32_csa28_csa_component_out[73];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[9] = u_CSAwallace_pg_rca32_csa28_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[10] = u_CSAwallace_pg_rca32_csa28_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[11] = u_CSAwallace_pg_rca32_csa28_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[12] = u_CSAwallace_pg_rca32_csa28_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[13] = u_CSAwallace_pg_rca32_csa28_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[14] = u_CSAwallace_pg_rca32_csa28_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[15] = u_CSAwallace_pg_rca32_csa28_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[16] = u_CSAwallace_pg_rca32_csa28_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[17] = u_CSAwallace_pg_rca32_csa28_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[18] = u_CSAwallace_pg_rca32_csa28_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[19] = u_CSAwallace_pg_rca32_csa28_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[20] = u_CSAwallace_pg_rca32_csa28_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[21] = u_CSAwallace_pg_rca32_csa28_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[22] = u_CSAwallace_pg_rca32_csa28_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[23] = u_CSAwallace_pg_rca32_csa28_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[24] = u_CSAwallace_pg_rca32_csa28_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[25] = u_CSAwallace_pg_rca32_csa28_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[26] = u_CSAwallace_pg_rca32_csa28_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[27] = u_CSAwallace_pg_rca32_csa28_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[28] = u_CSAwallace_pg_rca32_csa28_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[29] = u_CSAwallace_pg_rca32_csa28_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[30] = u_CSAwallace_pg_rca32_csa28_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[31] = u_CSAwallace_pg_rca32_csa28_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[32] = u_CSAwallace_pg_rca32_csa28_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[33] = u_CSAwallace_pg_rca32_csa28_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[34] = u_CSAwallace_pg_rca32_csa28_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[35] = u_CSAwallace_pg_rca32_csa28_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[36] = u_CSAwallace_pg_rca32_csa28_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[37] = u_CSAwallace_pg_rca32_csa28_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[38] = u_CSAwallace_pg_rca32_csa28_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[39] = u_CSAwallace_pg_rca32_csa28_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[40] = u_CSAwallace_pg_rca32_csa28_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[41] = u_CSAwallace_pg_rca32_csa28_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[42] = u_CSAwallace_pg_rca32_csa28_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[43] = u_CSAwallace_pg_rca32_csa28_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[44] = u_CSAwallace_pg_rca32_csa28_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[45] = u_CSAwallace_pg_rca32_csa28_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[46] = u_CSAwallace_pg_rca32_csa28_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[47] = u_CSAwallace_pg_rca32_csa28_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[48] = u_CSAwallace_pg_rca32_csa28_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[49] = u_CSAwallace_pg_rca32_csa28_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[50] = u_CSAwallace_pg_rca32_csa28_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[51] = u_CSAwallace_pg_rca32_csa28_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[52] = u_CSAwallace_pg_rca32_csa28_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[53] = u_CSAwallace_pg_rca32_csa28_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[54] = u_CSAwallace_pg_rca32_csa28_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[55] = u_CSAwallace_pg_rca32_csa28_csa_component_out[120];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[56] = u_CSAwallace_pg_rca32_csa28_csa_component_out[121];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[57] = u_CSAwallace_pg_rca32_csa28_csa_component_out[122];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[58] = u_CSAwallace_pg_rca32_csa28_csa_component_out[123];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[59] = u_CSAwallace_pg_rca32_csa28_csa_component_out[124];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[60] = u_CSAwallace_pg_rca32_csa28_csa_component_out[125];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[61] = u_CSAwallace_pg_rca32_csa28_csa_component_out[126];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[62] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[9] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[10] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[11] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[12] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[13] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[14] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[15] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[16] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[17] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[18] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[19] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[20] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[21] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[22] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[23] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[24] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[25] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[26] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[27] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[28] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[29] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[30] = 1'b0;
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[31] = u_CSAwallace_pg_rca32_csa21_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[32] = u_CSAwallace_pg_rca32_csa21_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[33] = u_CSAwallace_pg_rca32_csa21_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[34] = u_CSAwallace_pg_rca32_csa21_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[35] = u_CSAwallace_pg_rca32_csa21_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[36] = u_CSAwallace_pg_rca32_csa21_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[37] = u_CSAwallace_pg_rca32_csa21_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[38] = u_CSAwallace_pg_rca32_csa21_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[39] = u_CSAwallace_pg_rca32_csa21_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[40] = u_CSAwallace_pg_rca32_csa21_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[41] = u_CSAwallace_pg_rca32_csa21_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[42] = u_CSAwallace_pg_rca32_csa21_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[43] = u_CSAwallace_pg_rca32_csa21_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[44] = u_CSAwallace_pg_rca32_csa21_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[45] = u_CSAwallace_pg_rca32_csa21_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[46] = u_CSAwallace_pg_rca32_csa21_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[47] = u_CSAwallace_pg_rca32_csa21_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[48] = u_CSAwallace_pg_rca32_csa21_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[49] = u_CSAwallace_pg_rca32_csa21_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[50] = u_CSAwallace_pg_rca32_csa21_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[51] = u_CSAwallace_pg_rca32_csa21_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[52] = u_CSAwallace_pg_rca32_csa21_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[53] = u_CSAwallace_pg_rca32_csa21_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[54] = u_CSAwallace_pg_rca32_csa21_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[55] = u_CSAwallace_pg_rca32_csa21_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[56] = u_CSAwallace_pg_rca32_csa21_csa_component_out[120];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[57] = u_CSAwallace_pg_rca32_csa21_csa_component_out[121];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[58] = u_CSAwallace_pg_rca32_csa21_csa_component_out[122];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[59] = u_CSAwallace_pg_rca32_csa21_csa_component_out[123];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[60] = u_CSAwallace_pg_rca32_csa21_csa_component_out[124];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[61] = u_CSAwallace_pg_rca32_csa21_csa_component_out[125];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[62] = u_CSAwallace_pg_rca32_csa21_csa_component_out[126];
  assign u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22[63] = 1'b0;
  csa_component64 csa_component64_u_CSAwallace_pg_rca32_csa29_csa_component_out(.a(u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_s29), .b(u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c29), .c(u_CSAwallace_pg_rca32_csa29_csa_component_u_CSAwallace_pg_rca32_csa_c22), .csa_component64_out(u_CSAwallace_pg_rca32_csa29_csa_component_out));
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[0] = u_CSAwallace_pg_rca32_csa29_csa_component_out[0];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[1] = u_CSAwallace_pg_rca32_csa29_csa_component_out[1];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[2] = u_CSAwallace_pg_rca32_csa29_csa_component_out[2];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[3] = u_CSAwallace_pg_rca32_csa29_csa_component_out[3];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[4] = u_CSAwallace_pg_rca32_csa29_csa_component_out[4];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[5] = u_CSAwallace_pg_rca32_csa29_csa_component_out[5];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[6] = u_CSAwallace_pg_rca32_csa29_csa_component_out[6];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[7] = u_CSAwallace_pg_rca32_csa29_csa_component_out[7];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[8] = u_CSAwallace_pg_rca32_csa29_csa_component_out[8];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[9] = u_CSAwallace_pg_rca32_csa29_csa_component_out[9];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[10] = u_CSAwallace_pg_rca32_csa29_csa_component_out[10];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[11] = u_CSAwallace_pg_rca32_csa29_csa_component_out[11];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[12] = u_CSAwallace_pg_rca32_csa29_csa_component_out[12];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[13] = u_CSAwallace_pg_rca32_csa29_csa_component_out[13];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[14] = u_CSAwallace_pg_rca32_csa29_csa_component_out[14];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[15] = u_CSAwallace_pg_rca32_csa29_csa_component_out[15];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[16] = u_CSAwallace_pg_rca32_csa29_csa_component_out[16];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[17] = u_CSAwallace_pg_rca32_csa29_csa_component_out[17];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[18] = u_CSAwallace_pg_rca32_csa29_csa_component_out[18];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[19] = u_CSAwallace_pg_rca32_csa29_csa_component_out[19];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[20] = u_CSAwallace_pg_rca32_csa29_csa_component_out[20];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[21] = u_CSAwallace_pg_rca32_csa29_csa_component_out[21];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[22] = u_CSAwallace_pg_rca32_csa29_csa_component_out[22];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[23] = u_CSAwallace_pg_rca32_csa29_csa_component_out[23];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[24] = u_CSAwallace_pg_rca32_csa29_csa_component_out[24];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[25] = u_CSAwallace_pg_rca32_csa29_csa_component_out[25];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[26] = u_CSAwallace_pg_rca32_csa29_csa_component_out[26];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[27] = u_CSAwallace_pg_rca32_csa29_csa_component_out[27];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[28] = u_CSAwallace_pg_rca32_csa29_csa_component_out[28];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[29] = u_CSAwallace_pg_rca32_csa29_csa_component_out[29];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[30] = u_CSAwallace_pg_rca32_csa29_csa_component_out[30];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[31] = u_CSAwallace_pg_rca32_csa29_csa_component_out[31];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[32] = u_CSAwallace_pg_rca32_csa29_csa_component_out[32];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[33] = u_CSAwallace_pg_rca32_csa29_csa_component_out[33];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[34] = u_CSAwallace_pg_rca32_csa29_csa_component_out[34];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[35] = u_CSAwallace_pg_rca32_csa29_csa_component_out[35];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[36] = u_CSAwallace_pg_rca32_csa29_csa_component_out[36];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[37] = u_CSAwallace_pg_rca32_csa29_csa_component_out[37];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[38] = u_CSAwallace_pg_rca32_csa29_csa_component_out[38];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[39] = u_CSAwallace_pg_rca32_csa29_csa_component_out[39];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[40] = u_CSAwallace_pg_rca32_csa29_csa_component_out[40];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[41] = u_CSAwallace_pg_rca32_csa29_csa_component_out[41];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[42] = u_CSAwallace_pg_rca32_csa29_csa_component_out[42];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[43] = u_CSAwallace_pg_rca32_csa29_csa_component_out[43];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[44] = u_CSAwallace_pg_rca32_csa29_csa_component_out[44];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[45] = u_CSAwallace_pg_rca32_csa29_csa_component_out[45];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[46] = u_CSAwallace_pg_rca32_csa29_csa_component_out[46];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[47] = u_CSAwallace_pg_rca32_csa29_csa_component_out[47];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[48] = u_CSAwallace_pg_rca32_csa29_csa_component_out[48];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[49] = u_CSAwallace_pg_rca32_csa29_csa_component_out[49];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[50] = u_CSAwallace_pg_rca32_csa29_csa_component_out[50];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[51] = u_CSAwallace_pg_rca32_csa29_csa_component_out[51];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[52] = u_CSAwallace_pg_rca32_csa29_csa_component_out[52];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[53] = u_CSAwallace_pg_rca32_csa29_csa_component_out[53];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[54] = u_CSAwallace_pg_rca32_csa29_csa_component_out[54];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[55] = u_CSAwallace_pg_rca32_csa29_csa_component_out[55];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[56] = u_CSAwallace_pg_rca32_csa29_csa_component_out[56];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[57] = u_CSAwallace_pg_rca32_csa29_csa_component_out[57];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[58] = u_CSAwallace_pg_rca32_csa29_csa_component_out[58];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[59] = u_CSAwallace_pg_rca32_csa29_csa_component_out[59];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[60] = u_CSAwallace_pg_rca32_csa29_csa_component_out[60];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[61] = u_CSAwallace_pg_rca32_csa29_csa_component_out[61];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[62] = u_CSAwallace_pg_rca32_csa29_csa_component_out[62];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_a[63] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[0] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[1] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[2] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[3] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[4] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[5] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[6] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[7] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[8] = 1'b0;
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[9] = u_CSAwallace_pg_rca32_csa29_csa_component_out[74];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[10] = u_CSAwallace_pg_rca32_csa29_csa_component_out[75];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[11] = u_CSAwallace_pg_rca32_csa29_csa_component_out[76];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[12] = u_CSAwallace_pg_rca32_csa29_csa_component_out[77];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[13] = u_CSAwallace_pg_rca32_csa29_csa_component_out[78];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[14] = u_CSAwallace_pg_rca32_csa29_csa_component_out[79];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[15] = u_CSAwallace_pg_rca32_csa29_csa_component_out[80];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[16] = u_CSAwallace_pg_rca32_csa29_csa_component_out[81];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[17] = u_CSAwallace_pg_rca32_csa29_csa_component_out[82];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[18] = u_CSAwallace_pg_rca32_csa29_csa_component_out[83];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[19] = u_CSAwallace_pg_rca32_csa29_csa_component_out[84];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[20] = u_CSAwallace_pg_rca32_csa29_csa_component_out[85];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[21] = u_CSAwallace_pg_rca32_csa29_csa_component_out[86];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[22] = u_CSAwallace_pg_rca32_csa29_csa_component_out[87];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[23] = u_CSAwallace_pg_rca32_csa29_csa_component_out[88];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[24] = u_CSAwallace_pg_rca32_csa29_csa_component_out[89];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[25] = u_CSAwallace_pg_rca32_csa29_csa_component_out[90];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[26] = u_CSAwallace_pg_rca32_csa29_csa_component_out[91];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[27] = u_CSAwallace_pg_rca32_csa29_csa_component_out[92];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[28] = u_CSAwallace_pg_rca32_csa29_csa_component_out[93];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[29] = u_CSAwallace_pg_rca32_csa29_csa_component_out[94];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[30] = u_CSAwallace_pg_rca32_csa29_csa_component_out[95];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[31] = u_CSAwallace_pg_rca32_csa29_csa_component_out[96];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[32] = u_CSAwallace_pg_rca32_csa29_csa_component_out[97];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[33] = u_CSAwallace_pg_rca32_csa29_csa_component_out[98];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[34] = u_CSAwallace_pg_rca32_csa29_csa_component_out[99];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[35] = u_CSAwallace_pg_rca32_csa29_csa_component_out[100];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[36] = u_CSAwallace_pg_rca32_csa29_csa_component_out[101];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[37] = u_CSAwallace_pg_rca32_csa29_csa_component_out[102];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[38] = u_CSAwallace_pg_rca32_csa29_csa_component_out[103];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[39] = u_CSAwallace_pg_rca32_csa29_csa_component_out[104];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[40] = u_CSAwallace_pg_rca32_csa29_csa_component_out[105];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[41] = u_CSAwallace_pg_rca32_csa29_csa_component_out[106];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[42] = u_CSAwallace_pg_rca32_csa29_csa_component_out[107];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[43] = u_CSAwallace_pg_rca32_csa29_csa_component_out[108];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[44] = u_CSAwallace_pg_rca32_csa29_csa_component_out[109];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[45] = u_CSAwallace_pg_rca32_csa29_csa_component_out[110];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[46] = u_CSAwallace_pg_rca32_csa29_csa_component_out[111];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[47] = u_CSAwallace_pg_rca32_csa29_csa_component_out[112];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[48] = u_CSAwallace_pg_rca32_csa29_csa_component_out[113];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[49] = u_CSAwallace_pg_rca32_csa29_csa_component_out[114];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[50] = u_CSAwallace_pg_rca32_csa29_csa_component_out[115];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[51] = u_CSAwallace_pg_rca32_csa29_csa_component_out[116];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[52] = u_CSAwallace_pg_rca32_csa29_csa_component_out[117];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[53] = u_CSAwallace_pg_rca32_csa29_csa_component_out[118];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[54] = u_CSAwallace_pg_rca32_csa29_csa_component_out[119];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[55] = u_CSAwallace_pg_rca32_csa29_csa_component_out[120];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[56] = u_CSAwallace_pg_rca32_csa29_csa_component_out[121];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[57] = u_CSAwallace_pg_rca32_csa29_csa_component_out[122];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[58] = u_CSAwallace_pg_rca32_csa29_csa_component_out[123];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[59] = u_CSAwallace_pg_rca32_csa29_csa_component_out[124];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[60] = u_CSAwallace_pg_rca32_csa29_csa_component_out[125];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[61] = u_CSAwallace_pg_rca32_csa29_csa_component_out[126];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[62] = u_CSAwallace_pg_rca32_csa29_csa_component_out[127];
  assign u_CSAwallace_pg_rca32_u_pg_rca64_b[63] = u_CSAwallace_pg_rca32_csa29_csa_component_out[128];
  u_pg_rca64 u_pg_rca64_u_CSAwallace_pg_rca32_u_pg_rca64_out(.a(u_CSAwallace_pg_rca32_u_pg_rca64_a), .b(u_CSAwallace_pg_rca32_u_pg_rca64_b), .u_pg_rca64_out(u_CSAwallace_pg_rca32_u_pg_rca64_out));

  assign u_CSAwallace_pg_rca32_out[0] = u_CSAwallace_pg_rca32_u_pg_rca64_out[0];
  assign u_CSAwallace_pg_rca32_out[1] = u_CSAwallace_pg_rca32_u_pg_rca64_out[1];
  assign u_CSAwallace_pg_rca32_out[2] = u_CSAwallace_pg_rca32_u_pg_rca64_out[2];
  assign u_CSAwallace_pg_rca32_out[3] = u_CSAwallace_pg_rca32_u_pg_rca64_out[3];
  assign u_CSAwallace_pg_rca32_out[4] = u_CSAwallace_pg_rca32_u_pg_rca64_out[4];
  assign u_CSAwallace_pg_rca32_out[5] = u_CSAwallace_pg_rca32_u_pg_rca64_out[5];
  assign u_CSAwallace_pg_rca32_out[6] = u_CSAwallace_pg_rca32_u_pg_rca64_out[6];
  assign u_CSAwallace_pg_rca32_out[7] = u_CSAwallace_pg_rca32_u_pg_rca64_out[7];
  assign u_CSAwallace_pg_rca32_out[8] = u_CSAwallace_pg_rca32_u_pg_rca64_out[8];
  assign u_CSAwallace_pg_rca32_out[9] = u_CSAwallace_pg_rca32_u_pg_rca64_out[9];
  assign u_CSAwallace_pg_rca32_out[10] = u_CSAwallace_pg_rca32_u_pg_rca64_out[10];
  assign u_CSAwallace_pg_rca32_out[11] = u_CSAwallace_pg_rca32_u_pg_rca64_out[11];
  assign u_CSAwallace_pg_rca32_out[12] = u_CSAwallace_pg_rca32_u_pg_rca64_out[12];
  assign u_CSAwallace_pg_rca32_out[13] = u_CSAwallace_pg_rca32_u_pg_rca64_out[13];
  assign u_CSAwallace_pg_rca32_out[14] = u_CSAwallace_pg_rca32_u_pg_rca64_out[14];
  assign u_CSAwallace_pg_rca32_out[15] = u_CSAwallace_pg_rca32_u_pg_rca64_out[15];
  assign u_CSAwallace_pg_rca32_out[16] = u_CSAwallace_pg_rca32_u_pg_rca64_out[16];
  assign u_CSAwallace_pg_rca32_out[17] = u_CSAwallace_pg_rca32_u_pg_rca64_out[17];
  assign u_CSAwallace_pg_rca32_out[18] = u_CSAwallace_pg_rca32_u_pg_rca64_out[18];
  assign u_CSAwallace_pg_rca32_out[19] = u_CSAwallace_pg_rca32_u_pg_rca64_out[19];
  assign u_CSAwallace_pg_rca32_out[20] = u_CSAwallace_pg_rca32_u_pg_rca64_out[20];
  assign u_CSAwallace_pg_rca32_out[21] = u_CSAwallace_pg_rca32_u_pg_rca64_out[21];
  assign u_CSAwallace_pg_rca32_out[22] = u_CSAwallace_pg_rca32_u_pg_rca64_out[22];
  assign u_CSAwallace_pg_rca32_out[23] = u_CSAwallace_pg_rca32_u_pg_rca64_out[23];
  assign u_CSAwallace_pg_rca32_out[24] = u_CSAwallace_pg_rca32_u_pg_rca64_out[24];
  assign u_CSAwallace_pg_rca32_out[25] = u_CSAwallace_pg_rca32_u_pg_rca64_out[25];
  assign u_CSAwallace_pg_rca32_out[26] = u_CSAwallace_pg_rca32_u_pg_rca64_out[26];
  assign u_CSAwallace_pg_rca32_out[27] = u_CSAwallace_pg_rca32_u_pg_rca64_out[27];
  assign u_CSAwallace_pg_rca32_out[28] = u_CSAwallace_pg_rca32_u_pg_rca64_out[28];
  assign u_CSAwallace_pg_rca32_out[29] = u_CSAwallace_pg_rca32_u_pg_rca64_out[29];
  assign u_CSAwallace_pg_rca32_out[30] = u_CSAwallace_pg_rca32_u_pg_rca64_out[30];
  assign u_CSAwallace_pg_rca32_out[31] = u_CSAwallace_pg_rca32_u_pg_rca64_out[31];
  assign u_CSAwallace_pg_rca32_out[32] = u_CSAwallace_pg_rca32_u_pg_rca64_out[32];
  assign u_CSAwallace_pg_rca32_out[33] = u_CSAwallace_pg_rca32_u_pg_rca64_out[33];
  assign u_CSAwallace_pg_rca32_out[34] = u_CSAwallace_pg_rca32_u_pg_rca64_out[34];
  assign u_CSAwallace_pg_rca32_out[35] = u_CSAwallace_pg_rca32_u_pg_rca64_out[35];
  assign u_CSAwallace_pg_rca32_out[36] = u_CSAwallace_pg_rca32_u_pg_rca64_out[36];
  assign u_CSAwallace_pg_rca32_out[37] = u_CSAwallace_pg_rca32_u_pg_rca64_out[37];
  assign u_CSAwallace_pg_rca32_out[38] = u_CSAwallace_pg_rca32_u_pg_rca64_out[38];
  assign u_CSAwallace_pg_rca32_out[39] = u_CSAwallace_pg_rca32_u_pg_rca64_out[39];
  assign u_CSAwallace_pg_rca32_out[40] = u_CSAwallace_pg_rca32_u_pg_rca64_out[40];
  assign u_CSAwallace_pg_rca32_out[41] = u_CSAwallace_pg_rca32_u_pg_rca64_out[41];
  assign u_CSAwallace_pg_rca32_out[42] = u_CSAwallace_pg_rca32_u_pg_rca64_out[42];
  assign u_CSAwallace_pg_rca32_out[43] = u_CSAwallace_pg_rca32_u_pg_rca64_out[43];
  assign u_CSAwallace_pg_rca32_out[44] = u_CSAwallace_pg_rca32_u_pg_rca64_out[44];
  assign u_CSAwallace_pg_rca32_out[45] = u_CSAwallace_pg_rca32_u_pg_rca64_out[45];
  assign u_CSAwallace_pg_rca32_out[46] = u_CSAwallace_pg_rca32_u_pg_rca64_out[46];
  assign u_CSAwallace_pg_rca32_out[47] = u_CSAwallace_pg_rca32_u_pg_rca64_out[47];
  assign u_CSAwallace_pg_rca32_out[48] = u_CSAwallace_pg_rca32_u_pg_rca64_out[48];
  assign u_CSAwallace_pg_rca32_out[49] = u_CSAwallace_pg_rca32_u_pg_rca64_out[49];
  assign u_CSAwallace_pg_rca32_out[50] = u_CSAwallace_pg_rca32_u_pg_rca64_out[50];
  assign u_CSAwallace_pg_rca32_out[51] = u_CSAwallace_pg_rca32_u_pg_rca64_out[51];
  assign u_CSAwallace_pg_rca32_out[52] = u_CSAwallace_pg_rca32_u_pg_rca64_out[52];
  assign u_CSAwallace_pg_rca32_out[53] = u_CSAwallace_pg_rca32_u_pg_rca64_out[53];
  assign u_CSAwallace_pg_rca32_out[54] = u_CSAwallace_pg_rca32_u_pg_rca64_out[54];
  assign u_CSAwallace_pg_rca32_out[55] = u_CSAwallace_pg_rca32_u_pg_rca64_out[55];
  assign u_CSAwallace_pg_rca32_out[56] = u_CSAwallace_pg_rca32_u_pg_rca64_out[56];
  assign u_CSAwallace_pg_rca32_out[57] = u_CSAwallace_pg_rca32_u_pg_rca64_out[57];
  assign u_CSAwallace_pg_rca32_out[58] = u_CSAwallace_pg_rca32_u_pg_rca64_out[58];
  assign u_CSAwallace_pg_rca32_out[59] = u_CSAwallace_pg_rca32_u_pg_rca64_out[59];
  assign u_CSAwallace_pg_rca32_out[60] = u_CSAwallace_pg_rca32_u_pg_rca64_out[60];
  assign u_CSAwallace_pg_rca32_out[61] = u_CSAwallace_pg_rca32_u_pg_rca64_out[61];
  assign u_CSAwallace_pg_rca32_out[62] = u_CSAwallace_pg_rca32_u_pg_rca64_out[62];
  assign u_CSAwallace_pg_rca32_out[63] = u_CSAwallace_pg_rca32_u_pg_rca64_out[63];
endmodule