module f_s_dadda_pg_rca32(input [31:0] a, input [31:0] b, output [63:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire a_24;
  wire a_25;
  wire a_26;
  wire a_27;
  wire a_28;
  wire a_29;
  wire a_30;
  wire a_31;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire b_24;
  wire b_25;
  wire b_26;
  wire b_27;
  wire b_28;
  wire b_29;
  wire b_30;
  wire b_31;
  wire constant_wire_value_1_a_0;
  wire constant_wire_value_1_b_0;
  wire constant_wire_value_1_y0;
  wire constant_wire_value_1_y1;
  wire constant_wire_1;
  wire f_s_dadda_pg_rca32_and_28_0_a_28;
  wire f_s_dadda_pg_rca32_and_28_0_b_0;
  wire f_s_dadda_pg_rca32_and_28_0_y0;
  wire f_s_dadda_pg_rca32_and_27_1_a_27;
  wire f_s_dadda_pg_rca32_and_27_1_b_1;
  wire f_s_dadda_pg_rca32_and_27_1_y0;
  wire f_s_dadda_pg_rca32_ha0_f_s_dadda_pg_rca32_and_28_0_y0;
  wire f_s_dadda_pg_rca32_ha0_f_s_dadda_pg_rca32_and_27_1_y0;
  wire f_s_dadda_pg_rca32_ha0_y0;
  wire f_s_dadda_pg_rca32_ha0_y1;
  wire f_s_dadda_pg_rca32_and_29_0_a_29;
  wire f_s_dadda_pg_rca32_and_29_0_b_0;
  wire f_s_dadda_pg_rca32_and_29_0_y0;
  wire f_s_dadda_pg_rca32_and_28_1_a_28;
  wire f_s_dadda_pg_rca32_and_28_1_b_1;
  wire f_s_dadda_pg_rca32_and_28_1_y0;
  wire f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_ha0_y1;
  wire f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_and_29_0_y0;
  wire f_s_dadda_pg_rca32_fa0_y0;
  wire f_s_dadda_pg_rca32_fa0_y1;
  wire f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_and_28_1_y0;
  wire f_s_dadda_pg_rca32_fa0_y2;
  wire f_s_dadda_pg_rca32_fa0_y3;
  wire f_s_dadda_pg_rca32_fa0_y4;
  wire f_s_dadda_pg_rca32_and_27_2_a_27;
  wire f_s_dadda_pg_rca32_and_27_2_b_2;
  wire f_s_dadda_pg_rca32_and_27_2_y0;
  wire f_s_dadda_pg_rca32_and_26_3_a_26;
  wire f_s_dadda_pg_rca32_and_26_3_b_3;
  wire f_s_dadda_pg_rca32_and_26_3_y0;
  wire f_s_dadda_pg_rca32_ha1_f_s_dadda_pg_rca32_and_27_2_y0;
  wire f_s_dadda_pg_rca32_ha1_f_s_dadda_pg_rca32_and_26_3_y0;
  wire f_s_dadda_pg_rca32_ha1_y0;
  wire f_s_dadda_pg_rca32_ha1_y1;
  wire f_s_dadda_pg_rca32_and_30_0_a_30;
  wire f_s_dadda_pg_rca32_and_30_0_b_0;
  wire f_s_dadda_pg_rca32_and_30_0_y0;
  wire f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_ha1_y1;
  wire f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_fa0_y4;
  wire f_s_dadda_pg_rca32_fa1_y0;
  wire f_s_dadda_pg_rca32_fa1_y1;
  wire f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_and_30_0_y0;
  wire f_s_dadda_pg_rca32_fa1_y2;
  wire f_s_dadda_pg_rca32_fa1_y3;
  wire f_s_dadda_pg_rca32_fa1_y4;
  wire f_s_dadda_pg_rca32_and_29_1_a_29;
  wire f_s_dadda_pg_rca32_and_29_1_b_1;
  wire f_s_dadda_pg_rca32_and_29_1_y0;
  wire f_s_dadda_pg_rca32_and_28_2_a_28;
  wire f_s_dadda_pg_rca32_and_28_2_b_2;
  wire f_s_dadda_pg_rca32_and_28_2_y0;
  wire f_s_dadda_pg_rca32_and_27_3_a_27;
  wire f_s_dadda_pg_rca32_and_27_3_b_3;
  wire f_s_dadda_pg_rca32_and_27_3_y0;
  wire f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_29_1_y0;
  wire f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_28_2_y0;
  wire f_s_dadda_pg_rca32_fa2_y0;
  wire f_s_dadda_pg_rca32_fa2_y1;
  wire f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_27_3_y0;
  wire f_s_dadda_pg_rca32_fa2_y2;
  wire f_s_dadda_pg_rca32_fa2_y3;
  wire f_s_dadda_pg_rca32_fa2_y4;
  wire f_s_dadda_pg_rca32_and_26_4_a_26;
  wire f_s_dadda_pg_rca32_and_26_4_b_4;
  wire f_s_dadda_pg_rca32_and_26_4_y0;
  wire f_s_dadda_pg_rca32_and_25_5_a_25;
  wire f_s_dadda_pg_rca32_and_25_5_b_5;
  wire f_s_dadda_pg_rca32_and_25_5_y0;
  wire f_s_dadda_pg_rca32_ha2_f_s_dadda_pg_rca32_and_26_4_y0;
  wire f_s_dadda_pg_rca32_ha2_f_s_dadda_pg_rca32_and_25_5_y0;
  wire f_s_dadda_pg_rca32_ha2_y0;
  wire f_s_dadda_pg_rca32_ha2_y1;
  wire f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_ha2_y1;
  wire f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_fa2_y4;
  wire f_s_dadda_pg_rca32_fa3_y0;
  wire f_s_dadda_pg_rca32_fa3_y1;
  wire f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_fa1_y4;
  wire f_s_dadda_pg_rca32_fa3_y2;
  wire f_s_dadda_pg_rca32_fa3_y3;
  wire f_s_dadda_pg_rca32_fa3_y4;
  wire f_s_dadda_pg_rca32_nand_31_0_a_31;
  wire f_s_dadda_pg_rca32_nand_31_0_b_0;
  wire f_s_dadda_pg_rca32_nand_31_0_y0;
  wire f_s_dadda_pg_rca32_and_30_1_a_30;
  wire f_s_dadda_pg_rca32_and_30_1_b_1;
  wire f_s_dadda_pg_rca32_and_30_1_y0;
  wire f_s_dadda_pg_rca32_and_29_2_a_29;
  wire f_s_dadda_pg_rca32_and_29_2_b_2;
  wire f_s_dadda_pg_rca32_and_29_2_y0;
  wire f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_nand_31_0_y0;
  wire f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_and_30_1_y0;
  wire f_s_dadda_pg_rca32_fa4_y0;
  wire f_s_dadda_pg_rca32_fa4_y1;
  wire f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_and_29_2_y0;
  wire f_s_dadda_pg_rca32_fa4_y2;
  wire f_s_dadda_pg_rca32_fa4_y3;
  wire f_s_dadda_pg_rca32_fa4_y4;
  wire f_s_dadda_pg_rca32_and_28_3_a_28;
  wire f_s_dadda_pg_rca32_and_28_3_b_3;
  wire f_s_dadda_pg_rca32_and_28_3_y0;
  wire f_s_dadda_pg_rca32_and_27_4_a_27;
  wire f_s_dadda_pg_rca32_and_27_4_b_4;
  wire f_s_dadda_pg_rca32_and_27_4_y0;
  wire f_s_dadda_pg_rca32_and_26_5_a_26;
  wire f_s_dadda_pg_rca32_and_26_5_b_5;
  wire f_s_dadda_pg_rca32_and_26_5_y0;
  wire f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_28_3_y0;
  wire f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_27_4_y0;
  wire f_s_dadda_pg_rca32_fa5_y0;
  wire f_s_dadda_pg_rca32_fa5_y1;
  wire f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_26_5_y0;
  wire f_s_dadda_pg_rca32_fa5_y2;
  wire f_s_dadda_pg_rca32_fa5_y3;
  wire f_s_dadda_pg_rca32_fa5_y4;
  wire f_s_dadda_pg_rca32_and_25_6_a_25;
  wire f_s_dadda_pg_rca32_and_25_6_b_6;
  wire f_s_dadda_pg_rca32_and_25_6_y0;
  wire f_s_dadda_pg_rca32_and_24_7_a_24;
  wire f_s_dadda_pg_rca32_and_24_7_b_7;
  wire f_s_dadda_pg_rca32_and_24_7_y0;
  wire f_s_dadda_pg_rca32_ha3_f_s_dadda_pg_rca32_and_25_6_y0;
  wire f_s_dadda_pg_rca32_ha3_f_s_dadda_pg_rca32_and_24_7_y0;
  wire f_s_dadda_pg_rca32_ha3_y0;
  wire f_s_dadda_pg_rca32_ha3_y1;
  wire f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_ha3_y1;
  wire f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_fa5_y4;
  wire f_s_dadda_pg_rca32_fa6_y0;
  wire f_s_dadda_pg_rca32_fa6_y1;
  wire f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_fa4_y4;
  wire f_s_dadda_pg_rca32_fa6_y2;
  wire f_s_dadda_pg_rca32_fa6_y3;
  wire f_s_dadda_pg_rca32_fa6_y4;
  wire f_s_dadda_pg_rca32_nand_31_1_a_31;
  wire f_s_dadda_pg_rca32_nand_31_1_b_1;
  wire f_s_dadda_pg_rca32_nand_31_1_y0;
  wire f_s_dadda_pg_rca32_fa7_f_s_dadda_pg_rca32_fa3_y4;
  wire f_s_dadda_pg_rca32_fa7_constant_wire_1;
  wire f_s_dadda_pg_rca32_fa7_y0;
  wire f_s_dadda_pg_rca32_fa7_y1;
  wire f_s_dadda_pg_rca32_fa7_f_s_dadda_pg_rca32_nand_31_1_y0;
  wire f_s_dadda_pg_rca32_fa7_y2;
  wire f_s_dadda_pg_rca32_fa7_y3;
  wire f_s_dadda_pg_rca32_fa7_y4;
  wire f_s_dadda_pg_rca32_and_30_2_a_30;
  wire f_s_dadda_pg_rca32_and_30_2_b_2;
  wire f_s_dadda_pg_rca32_and_30_2_y0;
  wire f_s_dadda_pg_rca32_and_29_3_a_29;
  wire f_s_dadda_pg_rca32_and_29_3_b_3;
  wire f_s_dadda_pg_rca32_and_29_3_y0;
  wire f_s_dadda_pg_rca32_and_28_4_a_28;
  wire f_s_dadda_pg_rca32_and_28_4_b_4;
  wire f_s_dadda_pg_rca32_and_28_4_y0;
  wire f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_30_2_y0;
  wire f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_29_3_y0;
  wire f_s_dadda_pg_rca32_fa8_y0;
  wire f_s_dadda_pg_rca32_fa8_y1;
  wire f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_28_4_y0;
  wire f_s_dadda_pg_rca32_fa8_y2;
  wire f_s_dadda_pg_rca32_fa8_y3;
  wire f_s_dadda_pg_rca32_fa8_y4;
  wire f_s_dadda_pg_rca32_and_27_5_a_27;
  wire f_s_dadda_pg_rca32_and_27_5_b_5;
  wire f_s_dadda_pg_rca32_and_27_5_y0;
  wire f_s_dadda_pg_rca32_and_26_6_a_26;
  wire f_s_dadda_pg_rca32_and_26_6_b_6;
  wire f_s_dadda_pg_rca32_and_26_6_y0;
  wire f_s_dadda_pg_rca32_and_25_7_a_25;
  wire f_s_dadda_pg_rca32_and_25_7_b_7;
  wire f_s_dadda_pg_rca32_and_25_7_y0;
  wire f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_27_5_y0;
  wire f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_26_6_y0;
  wire f_s_dadda_pg_rca32_fa9_y0;
  wire f_s_dadda_pg_rca32_fa9_y1;
  wire f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_25_7_y0;
  wire f_s_dadda_pg_rca32_fa9_y2;
  wire f_s_dadda_pg_rca32_fa9_y3;
  wire f_s_dadda_pg_rca32_fa9_y4;
  wire f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa9_y4;
  wire f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa8_y4;
  wire f_s_dadda_pg_rca32_fa10_y0;
  wire f_s_dadda_pg_rca32_fa10_y1;
  wire f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa7_y4;
  wire f_s_dadda_pg_rca32_fa10_y2;
  wire f_s_dadda_pg_rca32_fa10_y3;
  wire f_s_dadda_pg_rca32_fa10_y4;
  wire f_s_dadda_pg_rca32_nand_31_2_a_31;
  wire f_s_dadda_pg_rca32_nand_31_2_b_2;
  wire f_s_dadda_pg_rca32_nand_31_2_y0;
  wire f_s_dadda_pg_rca32_and_30_3_a_30;
  wire f_s_dadda_pg_rca32_and_30_3_b_3;
  wire f_s_dadda_pg_rca32_and_30_3_y0;
  wire f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_fa6_y4;
  wire f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_nand_31_2_y0;
  wire f_s_dadda_pg_rca32_fa11_y0;
  wire f_s_dadda_pg_rca32_fa11_y1;
  wire f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_and_30_3_y0;
  wire f_s_dadda_pg_rca32_fa11_y2;
  wire f_s_dadda_pg_rca32_fa11_y3;
  wire f_s_dadda_pg_rca32_fa11_y4;
  wire f_s_dadda_pg_rca32_and_29_4_a_29;
  wire f_s_dadda_pg_rca32_and_29_4_b_4;
  wire f_s_dadda_pg_rca32_and_29_4_y0;
  wire f_s_dadda_pg_rca32_and_28_5_a_28;
  wire f_s_dadda_pg_rca32_and_28_5_b_5;
  wire f_s_dadda_pg_rca32_and_28_5_y0;
  wire f_s_dadda_pg_rca32_and_27_6_a_27;
  wire f_s_dadda_pg_rca32_and_27_6_b_6;
  wire f_s_dadda_pg_rca32_and_27_6_y0;
  wire f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_29_4_y0;
  wire f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_28_5_y0;
  wire f_s_dadda_pg_rca32_fa12_y0;
  wire f_s_dadda_pg_rca32_fa12_y1;
  wire f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_27_6_y0;
  wire f_s_dadda_pg_rca32_fa12_y2;
  wire f_s_dadda_pg_rca32_fa12_y3;
  wire f_s_dadda_pg_rca32_fa12_y4;
  wire f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa12_y4;
  wire f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa11_y4;
  wire f_s_dadda_pg_rca32_fa13_y0;
  wire f_s_dadda_pg_rca32_fa13_y1;
  wire f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa10_y4;
  wire f_s_dadda_pg_rca32_fa13_y2;
  wire f_s_dadda_pg_rca32_fa13_y3;
  wire f_s_dadda_pg_rca32_fa13_y4;
  wire f_s_dadda_pg_rca32_nand_31_3_a_31;
  wire f_s_dadda_pg_rca32_nand_31_3_b_3;
  wire f_s_dadda_pg_rca32_nand_31_3_y0;
  wire f_s_dadda_pg_rca32_and_30_4_a_30;
  wire f_s_dadda_pg_rca32_and_30_4_b_4;
  wire f_s_dadda_pg_rca32_and_30_4_y0;
  wire f_s_dadda_pg_rca32_and_29_5_a_29;
  wire f_s_dadda_pg_rca32_and_29_5_b_5;
  wire f_s_dadda_pg_rca32_and_29_5_y0;
  wire f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_nand_31_3_y0;
  wire f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_and_30_4_y0;
  wire f_s_dadda_pg_rca32_fa14_y0;
  wire f_s_dadda_pg_rca32_fa14_y1;
  wire f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_and_29_5_y0;
  wire f_s_dadda_pg_rca32_fa14_y2;
  wire f_s_dadda_pg_rca32_fa14_y3;
  wire f_s_dadda_pg_rca32_fa14_y4;
  wire f_s_dadda_pg_rca32_nand_31_4_a_31;
  wire f_s_dadda_pg_rca32_nand_31_4_b_4;
  wire f_s_dadda_pg_rca32_nand_31_4_y0;
  wire f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_fa14_y4;
  wire f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_fa13_y4;
  wire f_s_dadda_pg_rca32_fa15_y0;
  wire f_s_dadda_pg_rca32_fa15_y1;
  wire f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_nand_31_4_y0;
  wire f_s_dadda_pg_rca32_fa15_y2;
  wire f_s_dadda_pg_rca32_fa15_y3;
  wire f_s_dadda_pg_rca32_fa15_y4;
  wire f_s_dadda_pg_rca32_and_6_0_a_6;
  wire f_s_dadda_pg_rca32_and_6_0_b_0;
  wire f_s_dadda_pg_rca32_and_6_0_y0;
  wire f_s_dadda_pg_rca32_and_5_1_a_5;
  wire f_s_dadda_pg_rca32_and_5_1_b_1;
  wire f_s_dadda_pg_rca32_and_5_1_y0;
  wire f_s_dadda_pg_rca32_ha4_f_s_dadda_pg_rca32_and_6_0_y0;
  wire f_s_dadda_pg_rca32_ha4_f_s_dadda_pg_rca32_and_5_1_y0;
  wire f_s_dadda_pg_rca32_ha4_y0;
  wire f_s_dadda_pg_rca32_ha4_y1;
  wire f_s_dadda_pg_rca32_and_7_0_a_7;
  wire f_s_dadda_pg_rca32_and_7_0_b_0;
  wire f_s_dadda_pg_rca32_and_7_0_y0;
  wire f_s_dadda_pg_rca32_and_6_1_a_6;
  wire f_s_dadda_pg_rca32_and_6_1_b_1;
  wire f_s_dadda_pg_rca32_and_6_1_y0;
  wire f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_ha4_y1;
  wire f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_and_7_0_y0;
  wire f_s_dadda_pg_rca32_fa16_y0;
  wire f_s_dadda_pg_rca32_fa16_y1;
  wire f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_and_6_1_y0;
  wire f_s_dadda_pg_rca32_fa16_y2;
  wire f_s_dadda_pg_rca32_fa16_y3;
  wire f_s_dadda_pg_rca32_fa16_y4;
  wire f_s_dadda_pg_rca32_and_5_2_a_5;
  wire f_s_dadda_pg_rca32_and_5_2_b_2;
  wire f_s_dadda_pg_rca32_and_5_2_y0;
  wire f_s_dadda_pg_rca32_and_4_3_a_4;
  wire f_s_dadda_pg_rca32_and_4_3_b_3;
  wire f_s_dadda_pg_rca32_and_4_3_y0;
  wire f_s_dadda_pg_rca32_ha5_f_s_dadda_pg_rca32_and_5_2_y0;
  wire f_s_dadda_pg_rca32_ha5_f_s_dadda_pg_rca32_and_4_3_y0;
  wire f_s_dadda_pg_rca32_ha5_y0;
  wire f_s_dadda_pg_rca32_ha5_y1;
  wire f_s_dadda_pg_rca32_and_8_0_a_8;
  wire f_s_dadda_pg_rca32_and_8_0_b_0;
  wire f_s_dadda_pg_rca32_and_8_0_y0;
  wire f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_ha5_y1;
  wire f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_fa16_y4;
  wire f_s_dadda_pg_rca32_fa17_y0;
  wire f_s_dadda_pg_rca32_fa17_y1;
  wire f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_and_8_0_y0;
  wire f_s_dadda_pg_rca32_fa17_y2;
  wire f_s_dadda_pg_rca32_fa17_y3;
  wire f_s_dadda_pg_rca32_fa17_y4;
  wire f_s_dadda_pg_rca32_and_7_1_a_7;
  wire f_s_dadda_pg_rca32_and_7_1_b_1;
  wire f_s_dadda_pg_rca32_and_7_1_y0;
  wire f_s_dadda_pg_rca32_and_6_2_a_6;
  wire f_s_dadda_pg_rca32_and_6_2_b_2;
  wire f_s_dadda_pg_rca32_and_6_2_y0;
  wire f_s_dadda_pg_rca32_and_5_3_a_5;
  wire f_s_dadda_pg_rca32_and_5_3_b_3;
  wire f_s_dadda_pg_rca32_and_5_3_y0;
  wire f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_7_1_y0;
  wire f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_6_2_y0;
  wire f_s_dadda_pg_rca32_fa18_y0;
  wire f_s_dadda_pg_rca32_fa18_y1;
  wire f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_5_3_y0;
  wire f_s_dadda_pg_rca32_fa18_y2;
  wire f_s_dadda_pg_rca32_fa18_y3;
  wire f_s_dadda_pg_rca32_fa18_y4;
  wire f_s_dadda_pg_rca32_and_4_4_a_4;
  wire f_s_dadda_pg_rca32_and_4_4_b_4;
  wire f_s_dadda_pg_rca32_and_4_4_y0;
  wire f_s_dadda_pg_rca32_and_3_5_a_3;
  wire f_s_dadda_pg_rca32_and_3_5_b_5;
  wire f_s_dadda_pg_rca32_and_3_5_y0;
  wire f_s_dadda_pg_rca32_ha6_f_s_dadda_pg_rca32_and_4_4_y0;
  wire f_s_dadda_pg_rca32_ha6_f_s_dadda_pg_rca32_and_3_5_y0;
  wire f_s_dadda_pg_rca32_ha6_y0;
  wire f_s_dadda_pg_rca32_ha6_y1;
  wire f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_ha6_y1;
  wire f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_fa18_y4;
  wire f_s_dadda_pg_rca32_fa19_y0;
  wire f_s_dadda_pg_rca32_fa19_y1;
  wire f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_fa17_y4;
  wire f_s_dadda_pg_rca32_fa19_y2;
  wire f_s_dadda_pg_rca32_fa19_y3;
  wire f_s_dadda_pg_rca32_fa19_y4;
  wire f_s_dadda_pg_rca32_and_9_0_a_9;
  wire f_s_dadda_pg_rca32_and_9_0_b_0;
  wire f_s_dadda_pg_rca32_and_9_0_y0;
  wire f_s_dadda_pg_rca32_and_8_1_a_8;
  wire f_s_dadda_pg_rca32_and_8_1_b_1;
  wire f_s_dadda_pg_rca32_and_8_1_y0;
  wire f_s_dadda_pg_rca32_and_7_2_a_7;
  wire f_s_dadda_pg_rca32_and_7_2_b_2;
  wire f_s_dadda_pg_rca32_and_7_2_y0;
  wire f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_9_0_y0;
  wire f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_8_1_y0;
  wire f_s_dadda_pg_rca32_fa20_y0;
  wire f_s_dadda_pg_rca32_fa20_y1;
  wire f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_7_2_y0;
  wire f_s_dadda_pg_rca32_fa20_y2;
  wire f_s_dadda_pg_rca32_fa20_y3;
  wire f_s_dadda_pg_rca32_fa20_y4;
  wire f_s_dadda_pg_rca32_and_6_3_a_6;
  wire f_s_dadda_pg_rca32_and_6_3_b_3;
  wire f_s_dadda_pg_rca32_and_6_3_y0;
  wire f_s_dadda_pg_rca32_and_5_4_a_5;
  wire f_s_dadda_pg_rca32_and_5_4_b_4;
  wire f_s_dadda_pg_rca32_and_5_4_y0;
  wire f_s_dadda_pg_rca32_and_4_5_a_4;
  wire f_s_dadda_pg_rca32_and_4_5_b_5;
  wire f_s_dadda_pg_rca32_and_4_5_y0;
  wire f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_6_3_y0;
  wire f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_5_4_y0;
  wire f_s_dadda_pg_rca32_fa21_y0;
  wire f_s_dadda_pg_rca32_fa21_y1;
  wire f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_4_5_y0;
  wire f_s_dadda_pg_rca32_fa21_y2;
  wire f_s_dadda_pg_rca32_fa21_y3;
  wire f_s_dadda_pg_rca32_fa21_y4;
  wire f_s_dadda_pg_rca32_and_3_6_a_3;
  wire f_s_dadda_pg_rca32_and_3_6_b_6;
  wire f_s_dadda_pg_rca32_and_3_6_y0;
  wire f_s_dadda_pg_rca32_and_2_7_a_2;
  wire f_s_dadda_pg_rca32_and_2_7_b_7;
  wire f_s_dadda_pg_rca32_and_2_7_y0;
  wire f_s_dadda_pg_rca32_ha7_f_s_dadda_pg_rca32_and_3_6_y0;
  wire f_s_dadda_pg_rca32_ha7_f_s_dadda_pg_rca32_and_2_7_y0;
  wire f_s_dadda_pg_rca32_ha7_y0;
  wire f_s_dadda_pg_rca32_ha7_y1;
  wire f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_ha7_y1;
  wire f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_fa21_y4;
  wire f_s_dadda_pg_rca32_fa22_y0;
  wire f_s_dadda_pg_rca32_fa22_y1;
  wire f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_fa20_y4;
  wire f_s_dadda_pg_rca32_fa22_y2;
  wire f_s_dadda_pg_rca32_fa22_y3;
  wire f_s_dadda_pg_rca32_fa22_y4;
  wire f_s_dadda_pg_rca32_and_10_0_a_10;
  wire f_s_dadda_pg_rca32_and_10_0_b_0;
  wire f_s_dadda_pg_rca32_and_10_0_y0;
  wire f_s_dadda_pg_rca32_and_9_1_a_9;
  wire f_s_dadda_pg_rca32_and_9_1_b_1;
  wire f_s_dadda_pg_rca32_and_9_1_y0;
  wire f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_fa19_y4;
  wire f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_and_10_0_y0;
  wire f_s_dadda_pg_rca32_fa23_y0;
  wire f_s_dadda_pg_rca32_fa23_y1;
  wire f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_and_9_1_y0;
  wire f_s_dadda_pg_rca32_fa23_y2;
  wire f_s_dadda_pg_rca32_fa23_y3;
  wire f_s_dadda_pg_rca32_fa23_y4;
  wire f_s_dadda_pg_rca32_and_8_2_a_8;
  wire f_s_dadda_pg_rca32_and_8_2_b_2;
  wire f_s_dadda_pg_rca32_and_8_2_y0;
  wire f_s_dadda_pg_rca32_and_7_3_a_7;
  wire f_s_dadda_pg_rca32_and_7_3_b_3;
  wire f_s_dadda_pg_rca32_and_7_3_y0;
  wire f_s_dadda_pg_rca32_and_6_4_a_6;
  wire f_s_dadda_pg_rca32_and_6_4_b_4;
  wire f_s_dadda_pg_rca32_and_6_4_y0;
  wire f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_8_2_y0;
  wire f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_7_3_y0;
  wire f_s_dadda_pg_rca32_fa24_y0;
  wire f_s_dadda_pg_rca32_fa24_y1;
  wire f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_6_4_y0;
  wire f_s_dadda_pg_rca32_fa24_y2;
  wire f_s_dadda_pg_rca32_fa24_y3;
  wire f_s_dadda_pg_rca32_fa24_y4;
  wire f_s_dadda_pg_rca32_and_5_5_a_5;
  wire f_s_dadda_pg_rca32_and_5_5_b_5;
  wire f_s_dadda_pg_rca32_and_5_5_y0;
  wire f_s_dadda_pg_rca32_and_4_6_a_4;
  wire f_s_dadda_pg_rca32_and_4_6_b_6;
  wire f_s_dadda_pg_rca32_and_4_6_y0;
  wire f_s_dadda_pg_rca32_and_3_7_a_3;
  wire f_s_dadda_pg_rca32_and_3_7_b_7;
  wire f_s_dadda_pg_rca32_and_3_7_y0;
  wire f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_5_5_y0;
  wire f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_4_6_y0;
  wire f_s_dadda_pg_rca32_fa25_y0;
  wire f_s_dadda_pg_rca32_fa25_y1;
  wire f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_3_7_y0;
  wire f_s_dadda_pg_rca32_fa25_y2;
  wire f_s_dadda_pg_rca32_fa25_y3;
  wire f_s_dadda_pg_rca32_fa25_y4;
  wire f_s_dadda_pg_rca32_and_2_8_a_2;
  wire f_s_dadda_pg_rca32_and_2_8_b_8;
  wire f_s_dadda_pg_rca32_and_2_8_y0;
  wire f_s_dadda_pg_rca32_and_1_9_a_1;
  wire f_s_dadda_pg_rca32_and_1_9_b_9;
  wire f_s_dadda_pg_rca32_and_1_9_y0;
  wire f_s_dadda_pg_rca32_ha8_f_s_dadda_pg_rca32_and_2_8_y0;
  wire f_s_dadda_pg_rca32_ha8_f_s_dadda_pg_rca32_and_1_9_y0;
  wire f_s_dadda_pg_rca32_ha8_y0;
  wire f_s_dadda_pg_rca32_ha8_y1;
  wire f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_ha8_y1;
  wire f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_fa25_y4;
  wire f_s_dadda_pg_rca32_fa26_y0;
  wire f_s_dadda_pg_rca32_fa26_y1;
  wire f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_fa24_y4;
  wire f_s_dadda_pg_rca32_fa26_y2;
  wire f_s_dadda_pg_rca32_fa26_y3;
  wire f_s_dadda_pg_rca32_fa26_y4;
  wire f_s_dadda_pg_rca32_and_11_0_a_11;
  wire f_s_dadda_pg_rca32_and_11_0_b_0;
  wire f_s_dadda_pg_rca32_and_11_0_y0;
  wire f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_fa23_y4;
  wire f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_fa22_y4;
  wire f_s_dadda_pg_rca32_fa27_y0;
  wire f_s_dadda_pg_rca32_fa27_y1;
  wire f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_and_11_0_y0;
  wire f_s_dadda_pg_rca32_fa27_y2;
  wire f_s_dadda_pg_rca32_fa27_y3;
  wire f_s_dadda_pg_rca32_fa27_y4;
  wire f_s_dadda_pg_rca32_and_10_1_a_10;
  wire f_s_dadda_pg_rca32_and_10_1_b_1;
  wire f_s_dadda_pg_rca32_and_10_1_y0;
  wire f_s_dadda_pg_rca32_and_9_2_a_9;
  wire f_s_dadda_pg_rca32_and_9_2_b_2;
  wire f_s_dadda_pg_rca32_and_9_2_y0;
  wire f_s_dadda_pg_rca32_and_8_3_a_8;
  wire f_s_dadda_pg_rca32_and_8_3_b_3;
  wire f_s_dadda_pg_rca32_and_8_3_y0;
  wire f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_10_1_y0;
  wire f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_9_2_y0;
  wire f_s_dadda_pg_rca32_fa28_y0;
  wire f_s_dadda_pg_rca32_fa28_y1;
  wire f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_8_3_y0;
  wire f_s_dadda_pg_rca32_fa28_y2;
  wire f_s_dadda_pg_rca32_fa28_y3;
  wire f_s_dadda_pg_rca32_fa28_y4;
  wire f_s_dadda_pg_rca32_and_7_4_a_7;
  wire f_s_dadda_pg_rca32_and_7_4_b_4;
  wire f_s_dadda_pg_rca32_and_7_4_y0;
  wire f_s_dadda_pg_rca32_and_6_5_a_6;
  wire f_s_dadda_pg_rca32_and_6_5_b_5;
  wire f_s_dadda_pg_rca32_and_6_5_y0;
  wire f_s_dadda_pg_rca32_and_5_6_a_5;
  wire f_s_dadda_pg_rca32_and_5_6_b_6;
  wire f_s_dadda_pg_rca32_and_5_6_y0;
  wire f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_7_4_y0;
  wire f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_6_5_y0;
  wire f_s_dadda_pg_rca32_fa29_y0;
  wire f_s_dadda_pg_rca32_fa29_y1;
  wire f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_5_6_y0;
  wire f_s_dadda_pg_rca32_fa29_y2;
  wire f_s_dadda_pg_rca32_fa29_y3;
  wire f_s_dadda_pg_rca32_fa29_y4;
  wire f_s_dadda_pg_rca32_and_4_7_a_4;
  wire f_s_dadda_pg_rca32_and_4_7_b_7;
  wire f_s_dadda_pg_rca32_and_4_7_y0;
  wire f_s_dadda_pg_rca32_and_3_8_a_3;
  wire f_s_dadda_pg_rca32_and_3_8_b_8;
  wire f_s_dadda_pg_rca32_and_3_8_y0;
  wire f_s_dadda_pg_rca32_and_2_9_a_2;
  wire f_s_dadda_pg_rca32_and_2_9_b_9;
  wire f_s_dadda_pg_rca32_and_2_9_y0;
  wire f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_4_7_y0;
  wire f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_3_8_y0;
  wire f_s_dadda_pg_rca32_fa30_y0;
  wire f_s_dadda_pg_rca32_fa30_y1;
  wire f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_2_9_y0;
  wire f_s_dadda_pg_rca32_fa30_y2;
  wire f_s_dadda_pg_rca32_fa30_y3;
  wire f_s_dadda_pg_rca32_fa30_y4;
  wire f_s_dadda_pg_rca32_and_1_10_a_1;
  wire f_s_dadda_pg_rca32_and_1_10_b_10;
  wire f_s_dadda_pg_rca32_and_1_10_y0;
  wire f_s_dadda_pg_rca32_and_0_11_a_0;
  wire f_s_dadda_pg_rca32_and_0_11_b_11;
  wire f_s_dadda_pg_rca32_and_0_11_y0;
  wire f_s_dadda_pg_rca32_ha9_f_s_dadda_pg_rca32_and_1_10_y0;
  wire f_s_dadda_pg_rca32_ha9_f_s_dadda_pg_rca32_and_0_11_y0;
  wire f_s_dadda_pg_rca32_ha9_y0;
  wire f_s_dadda_pg_rca32_ha9_y1;
  wire f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_ha9_y1;
  wire f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_fa30_y4;
  wire f_s_dadda_pg_rca32_fa31_y0;
  wire f_s_dadda_pg_rca32_fa31_y1;
  wire f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_fa29_y4;
  wire f_s_dadda_pg_rca32_fa31_y2;
  wire f_s_dadda_pg_rca32_fa31_y3;
  wire f_s_dadda_pg_rca32_fa31_y4;
  wire f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa28_y4;
  wire f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa27_y4;
  wire f_s_dadda_pg_rca32_fa32_y0;
  wire f_s_dadda_pg_rca32_fa32_y1;
  wire f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa26_y4;
  wire f_s_dadda_pg_rca32_fa32_y2;
  wire f_s_dadda_pg_rca32_fa32_y3;
  wire f_s_dadda_pg_rca32_fa32_y4;
  wire f_s_dadda_pg_rca32_and_12_0_a_12;
  wire f_s_dadda_pg_rca32_and_12_0_b_0;
  wire f_s_dadda_pg_rca32_and_12_0_y0;
  wire f_s_dadda_pg_rca32_and_11_1_a_11;
  wire f_s_dadda_pg_rca32_and_11_1_b_1;
  wire f_s_dadda_pg_rca32_and_11_1_y0;
  wire f_s_dadda_pg_rca32_and_10_2_a_10;
  wire f_s_dadda_pg_rca32_and_10_2_b_2;
  wire f_s_dadda_pg_rca32_and_10_2_y0;
  wire f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_12_0_y0;
  wire f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_11_1_y0;
  wire f_s_dadda_pg_rca32_fa33_y0;
  wire f_s_dadda_pg_rca32_fa33_y1;
  wire f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_10_2_y0;
  wire f_s_dadda_pg_rca32_fa33_y2;
  wire f_s_dadda_pg_rca32_fa33_y3;
  wire f_s_dadda_pg_rca32_fa33_y4;
  wire f_s_dadda_pg_rca32_and_9_3_a_9;
  wire f_s_dadda_pg_rca32_and_9_3_b_3;
  wire f_s_dadda_pg_rca32_and_9_3_y0;
  wire f_s_dadda_pg_rca32_and_8_4_a_8;
  wire f_s_dadda_pg_rca32_and_8_4_b_4;
  wire f_s_dadda_pg_rca32_and_8_4_y0;
  wire f_s_dadda_pg_rca32_and_7_5_a_7;
  wire f_s_dadda_pg_rca32_and_7_5_b_5;
  wire f_s_dadda_pg_rca32_and_7_5_y0;
  wire f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_9_3_y0;
  wire f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_8_4_y0;
  wire f_s_dadda_pg_rca32_fa34_y0;
  wire f_s_dadda_pg_rca32_fa34_y1;
  wire f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_7_5_y0;
  wire f_s_dadda_pg_rca32_fa34_y2;
  wire f_s_dadda_pg_rca32_fa34_y3;
  wire f_s_dadda_pg_rca32_fa34_y4;
  wire f_s_dadda_pg_rca32_and_6_6_a_6;
  wire f_s_dadda_pg_rca32_and_6_6_b_6;
  wire f_s_dadda_pg_rca32_and_6_6_y0;
  wire f_s_dadda_pg_rca32_and_5_7_a_5;
  wire f_s_dadda_pg_rca32_and_5_7_b_7;
  wire f_s_dadda_pg_rca32_and_5_7_y0;
  wire f_s_dadda_pg_rca32_and_4_8_a_4;
  wire f_s_dadda_pg_rca32_and_4_8_b_8;
  wire f_s_dadda_pg_rca32_and_4_8_y0;
  wire f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_6_6_y0;
  wire f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_5_7_y0;
  wire f_s_dadda_pg_rca32_fa35_y0;
  wire f_s_dadda_pg_rca32_fa35_y1;
  wire f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_4_8_y0;
  wire f_s_dadda_pg_rca32_fa35_y2;
  wire f_s_dadda_pg_rca32_fa35_y3;
  wire f_s_dadda_pg_rca32_fa35_y4;
  wire f_s_dadda_pg_rca32_and_3_9_a_3;
  wire f_s_dadda_pg_rca32_and_3_9_b_9;
  wire f_s_dadda_pg_rca32_and_3_9_y0;
  wire f_s_dadda_pg_rca32_and_2_10_a_2;
  wire f_s_dadda_pg_rca32_and_2_10_b_10;
  wire f_s_dadda_pg_rca32_and_2_10_y0;
  wire f_s_dadda_pg_rca32_and_1_11_a_1;
  wire f_s_dadda_pg_rca32_and_1_11_b_11;
  wire f_s_dadda_pg_rca32_and_1_11_y0;
  wire f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_3_9_y0;
  wire f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_2_10_y0;
  wire f_s_dadda_pg_rca32_fa36_y0;
  wire f_s_dadda_pg_rca32_fa36_y1;
  wire f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_1_11_y0;
  wire f_s_dadda_pg_rca32_fa36_y2;
  wire f_s_dadda_pg_rca32_fa36_y3;
  wire f_s_dadda_pg_rca32_fa36_y4;
  wire f_s_dadda_pg_rca32_and_0_12_a_0;
  wire f_s_dadda_pg_rca32_and_0_12_b_12;
  wire f_s_dadda_pg_rca32_and_0_12_y0;
  wire f_s_dadda_pg_rca32_ha10_f_s_dadda_pg_rca32_and_0_12_y0;
  wire f_s_dadda_pg_rca32_ha10_f_s_dadda_pg_rca32_fa31_y2;
  wire f_s_dadda_pg_rca32_ha10_y0;
  wire f_s_dadda_pg_rca32_ha10_y1;
  wire f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_ha10_y1;
  wire f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_fa36_y4;
  wire f_s_dadda_pg_rca32_fa37_y0;
  wire f_s_dadda_pg_rca32_fa37_y1;
  wire f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_fa35_y4;
  wire f_s_dadda_pg_rca32_fa37_y2;
  wire f_s_dadda_pg_rca32_fa37_y3;
  wire f_s_dadda_pg_rca32_fa37_y4;
  wire f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa34_y4;
  wire f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa33_y4;
  wire f_s_dadda_pg_rca32_fa38_y0;
  wire f_s_dadda_pg_rca32_fa38_y1;
  wire f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa32_y4;
  wire f_s_dadda_pg_rca32_fa38_y2;
  wire f_s_dadda_pg_rca32_fa38_y3;
  wire f_s_dadda_pg_rca32_fa38_y4;
  wire f_s_dadda_pg_rca32_and_13_0_a_13;
  wire f_s_dadda_pg_rca32_and_13_0_b_0;
  wire f_s_dadda_pg_rca32_and_13_0_y0;
  wire f_s_dadda_pg_rca32_and_12_1_a_12;
  wire f_s_dadda_pg_rca32_and_12_1_b_1;
  wire f_s_dadda_pg_rca32_and_12_1_y0;
  wire f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_fa31_y4;
  wire f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_and_13_0_y0;
  wire f_s_dadda_pg_rca32_fa39_y0;
  wire f_s_dadda_pg_rca32_fa39_y1;
  wire f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_and_12_1_y0;
  wire f_s_dadda_pg_rca32_fa39_y2;
  wire f_s_dadda_pg_rca32_fa39_y3;
  wire f_s_dadda_pg_rca32_fa39_y4;
  wire f_s_dadda_pg_rca32_and_11_2_a_11;
  wire f_s_dadda_pg_rca32_and_11_2_b_2;
  wire f_s_dadda_pg_rca32_and_11_2_y0;
  wire f_s_dadda_pg_rca32_and_10_3_a_10;
  wire f_s_dadda_pg_rca32_and_10_3_b_3;
  wire f_s_dadda_pg_rca32_and_10_3_y0;
  wire f_s_dadda_pg_rca32_and_9_4_a_9;
  wire f_s_dadda_pg_rca32_and_9_4_b_4;
  wire f_s_dadda_pg_rca32_and_9_4_y0;
  wire f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_11_2_y0;
  wire f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_10_3_y0;
  wire f_s_dadda_pg_rca32_fa40_y0;
  wire f_s_dadda_pg_rca32_fa40_y1;
  wire f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_9_4_y0;
  wire f_s_dadda_pg_rca32_fa40_y2;
  wire f_s_dadda_pg_rca32_fa40_y3;
  wire f_s_dadda_pg_rca32_fa40_y4;
  wire f_s_dadda_pg_rca32_and_8_5_a_8;
  wire f_s_dadda_pg_rca32_and_8_5_b_5;
  wire f_s_dadda_pg_rca32_and_8_5_y0;
  wire f_s_dadda_pg_rca32_and_7_6_a_7;
  wire f_s_dadda_pg_rca32_and_7_6_b_6;
  wire f_s_dadda_pg_rca32_and_7_6_y0;
  wire f_s_dadda_pg_rca32_and_6_7_a_6;
  wire f_s_dadda_pg_rca32_and_6_7_b_7;
  wire f_s_dadda_pg_rca32_and_6_7_y0;
  wire f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_8_5_y0;
  wire f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_7_6_y0;
  wire f_s_dadda_pg_rca32_fa41_y0;
  wire f_s_dadda_pg_rca32_fa41_y1;
  wire f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_6_7_y0;
  wire f_s_dadda_pg_rca32_fa41_y2;
  wire f_s_dadda_pg_rca32_fa41_y3;
  wire f_s_dadda_pg_rca32_fa41_y4;
  wire f_s_dadda_pg_rca32_and_5_8_a_5;
  wire f_s_dadda_pg_rca32_and_5_8_b_8;
  wire f_s_dadda_pg_rca32_and_5_8_y0;
  wire f_s_dadda_pg_rca32_and_4_9_a_4;
  wire f_s_dadda_pg_rca32_and_4_9_b_9;
  wire f_s_dadda_pg_rca32_and_4_9_y0;
  wire f_s_dadda_pg_rca32_and_3_10_a_3;
  wire f_s_dadda_pg_rca32_and_3_10_b_10;
  wire f_s_dadda_pg_rca32_and_3_10_y0;
  wire f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_5_8_y0;
  wire f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_4_9_y0;
  wire f_s_dadda_pg_rca32_fa42_y0;
  wire f_s_dadda_pg_rca32_fa42_y1;
  wire f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_3_10_y0;
  wire f_s_dadda_pg_rca32_fa42_y2;
  wire f_s_dadda_pg_rca32_fa42_y3;
  wire f_s_dadda_pg_rca32_fa42_y4;
  wire f_s_dadda_pg_rca32_and_2_11_a_2;
  wire f_s_dadda_pg_rca32_and_2_11_b_11;
  wire f_s_dadda_pg_rca32_and_2_11_y0;
  wire f_s_dadda_pg_rca32_and_1_12_a_1;
  wire f_s_dadda_pg_rca32_and_1_12_b_12;
  wire f_s_dadda_pg_rca32_and_1_12_y0;
  wire f_s_dadda_pg_rca32_and_0_13_a_0;
  wire f_s_dadda_pg_rca32_and_0_13_b_13;
  wire f_s_dadda_pg_rca32_and_0_13_y0;
  wire f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_2_11_y0;
  wire f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_1_12_y0;
  wire f_s_dadda_pg_rca32_fa43_y0;
  wire f_s_dadda_pg_rca32_fa43_y1;
  wire f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_0_13_y0;
  wire f_s_dadda_pg_rca32_fa43_y2;
  wire f_s_dadda_pg_rca32_fa43_y3;
  wire f_s_dadda_pg_rca32_fa43_y4;
  wire f_s_dadda_pg_rca32_ha11_f_s_dadda_pg_rca32_fa37_y2;
  wire f_s_dadda_pg_rca32_ha11_f_s_dadda_pg_rca32_fa38_y2;
  wire f_s_dadda_pg_rca32_ha11_y0;
  wire f_s_dadda_pg_rca32_ha11_y1;
  wire f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_ha11_y1;
  wire f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_fa43_y4;
  wire f_s_dadda_pg_rca32_fa44_y0;
  wire f_s_dadda_pg_rca32_fa44_y1;
  wire f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_fa42_y4;
  wire f_s_dadda_pg_rca32_fa44_y2;
  wire f_s_dadda_pg_rca32_fa44_y3;
  wire f_s_dadda_pg_rca32_fa44_y4;
  wire f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa41_y4;
  wire f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa40_y4;
  wire f_s_dadda_pg_rca32_fa45_y0;
  wire f_s_dadda_pg_rca32_fa45_y1;
  wire f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa39_y4;
  wire f_s_dadda_pg_rca32_fa45_y2;
  wire f_s_dadda_pg_rca32_fa45_y3;
  wire f_s_dadda_pg_rca32_fa45_y4;
  wire f_s_dadda_pg_rca32_and_14_0_a_14;
  wire f_s_dadda_pg_rca32_and_14_0_b_0;
  wire f_s_dadda_pg_rca32_and_14_0_y0;
  wire f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_fa38_y4;
  wire f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_fa37_y4;
  wire f_s_dadda_pg_rca32_fa46_y0;
  wire f_s_dadda_pg_rca32_fa46_y1;
  wire f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_and_14_0_y0;
  wire f_s_dadda_pg_rca32_fa46_y2;
  wire f_s_dadda_pg_rca32_fa46_y3;
  wire f_s_dadda_pg_rca32_fa46_y4;
  wire f_s_dadda_pg_rca32_and_13_1_a_13;
  wire f_s_dadda_pg_rca32_and_13_1_b_1;
  wire f_s_dadda_pg_rca32_and_13_1_y0;
  wire f_s_dadda_pg_rca32_and_12_2_a_12;
  wire f_s_dadda_pg_rca32_and_12_2_b_2;
  wire f_s_dadda_pg_rca32_and_12_2_y0;
  wire f_s_dadda_pg_rca32_and_11_3_a_11;
  wire f_s_dadda_pg_rca32_and_11_3_b_3;
  wire f_s_dadda_pg_rca32_and_11_3_y0;
  wire f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_13_1_y0;
  wire f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_12_2_y0;
  wire f_s_dadda_pg_rca32_fa47_y0;
  wire f_s_dadda_pg_rca32_fa47_y1;
  wire f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_11_3_y0;
  wire f_s_dadda_pg_rca32_fa47_y2;
  wire f_s_dadda_pg_rca32_fa47_y3;
  wire f_s_dadda_pg_rca32_fa47_y4;
  wire f_s_dadda_pg_rca32_and_10_4_a_10;
  wire f_s_dadda_pg_rca32_and_10_4_b_4;
  wire f_s_dadda_pg_rca32_and_10_4_y0;
  wire f_s_dadda_pg_rca32_and_9_5_a_9;
  wire f_s_dadda_pg_rca32_and_9_5_b_5;
  wire f_s_dadda_pg_rca32_and_9_5_y0;
  wire f_s_dadda_pg_rca32_and_8_6_a_8;
  wire f_s_dadda_pg_rca32_and_8_6_b_6;
  wire f_s_dadda_pg_rca32_and_8_6_y0;
  wire f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_10_4_y0;
  wire f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_9_5_y0;
  wire f_s_dadda_pg_rca32_fa48_y0;
  wire f_s_dadda_pg_rca32_fa48_y1;
  wire f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_8_6_y0;
  wire f_s_dadda_pg_rca32_fa48_y2;
  wire f_s_dadda_pg_rca32_fa48_y3;
  wire f_s_dadda_pg_rca32_fa48_y4;
  wire f_s_dadda_pg_rca32_and_7_7_a_7;
  wire f_s_dadda_pg_rca32_and_7_7_b_7;
  wire f_s_dadda_pg_rca32_and_7_7_y0;
  wire f_s_dadda_pg_rca32_and_6_8_a_6;
  wire f_s_dadda_pg_rca32_and_6_8_b_8;
  wire f_s_dadda_pg_rca32_and_6_8_y0;
  wire f_s_dadda_pg_rca32_and_5_9_a_5;
  wire f_s_dadda_pg_rca32_and_5_9_b_9;
  wire f_s_dadda_pg_rca32_and_5_9_y0;
  wire f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_7_7_y0;
  wire f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_6_8_y0;
  wire f_s_dadda_pg_rca32_fa49_y0;
  wire f_s_dadda_pg_rca32_fa49_y1;
  wire f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_5_9_y0;
  wire f_s_dadda_pg_rca32_fa49_y2;
  wire f_s_dadda_pg_rca32_fa49_y3;
  wire f_s_dadda_pg_rca32_fa49_y4;
  wire f_s_dadda_pg_rca32_and_4_10_a_4;
  wire f_s_dadda_pg_rca32_and_4_10_b_10;
  wire f_s_dadda_pg_rca32_and_4_10_y0;
  wire f_s_dadda_pg_rca32_and_3_11_a_3;
  wire f_s_dadda_pg_rca32_and_3_11_b_11;
  wire f_s_dadda_pg_rca32_and_3_11_y0;
  wire f_s_dadda_pg_rca32_and_2_12_a_2;
  wire f_s_dadda_pg_rca32_and_2_12_b_12;
  wire f_s_dadda_pg_rca32_and_2_12_y0;
  wire f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_4_10_y0;
  wire f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_3_11_y0;
  wire f_s_dadda_pg_rca32_fa50_y0;
  wire f_s_dadda_pg_rca32_fa50_y1;
  wire f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_2_12_y0;
  wire f_s_dadda_pg_rca32_fa50_y2;
  wire f_s_dadda_pg_rca32_fa50_y3;
  wire f_s_dadda_pg_rca32_fa50_y4;
  wire f_s_dadda_pg_rca32_and_1_13_a_1;
  wire f_s_dadda_pg_rca32_and_1_13_b_13;
  wire f_s_dadda_pg_rca32_and_1_13_y0;
  wire f_s_dadda_pg_rca32_and_0_14_a_0;
  wire f_s_dadda_pg_rca32_and_0_14_b_14;
  wire f_s_dadda_pg_rca32_and_0_14_y0;
  wire f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_and_1_13_y0;
  wire f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_and_0_14_y0;
  wire f_s_dadda_pg_rca32_fa51_y0;
  wire f_s_dadda_pg_rca32_fa51_y1;
  wire f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_fa44_y2;
  wire f_s_dadda_pg_rca32_fa51_y2;
  wire f_s_dadda_pg_rca32_fa51_y3;
  wire f_s_dadda_pg_rca32_fa51_y4;
  wire f_s_dadda_pg_rca32_ha12_f_s_dadda_pg_rca32_fa45_y2;
  wire f_s_dadda_pg_rca32_ha12_f_s_dadda_pg_rca32_fa46_y2;
  wire f_s_dadda_pg_rca32_ha12_y0;
  wire f_s_dadda_pg_rca32_ha12_y1;
  wire f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_ha12_y1;
  wire f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_fa51_y4;
  wire f_s_dadda_pg_rca32_fa52_y0;
  wire f_s_dadda_pg_rca32_fa52_y1;
  wire f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_fa50_y4;
  wire f_s_dadda_pg_rca32_fa52_y2;
  wire f_s_dadda_pg_rca32_fa52_y3;
  wire f_s_dadda_pg_rca32_fa52_y4;
  wire f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa49_y4;
  wire f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa48_y4;
  wire f_s_dadda_pg_rca32_fa53_y0;
  wire f_s_dadda_pg_rca32_fa53_y1;
  wire f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa47_y4;
  wire f_s_dadda_pg_rca32_fa53_y2;
  wire f_s_dadda_pg_rca32_fa53_y3;
  wire f_s_dadda_pg_rca32_fa53_y4;
  wire f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa46_y4;
  wire f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa45_y4;
  wire f_s_dadda_pg_rca32_fa54_y0;
  wire f_s_dadda_pg_rca32_fa54_y1;
  wire f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa44_y4;
  wire f_s_dadda_pg_rca32_fa54_y2;
  wire f_s_dadda_pg_rca32_fa54_y3;
  wire f_s_dadda_pg_rca32_fa54_y4;
  wire f_s_dadda_pg_rca32_and_15_0_a_15;
  wire f_s_dadda_pg_rca32_and_15_0_b_0;
  wire f_s_dadda_pg_rca32_and_15_0_y0;
  wire f_s_dadda_pg_rca32_and_14_1_a_14;
  wire f_s_dadda_pg_rca32_and_14_1_b_1;
  wire f_s_dadda_pg_rca32_and_14_1_y0;
  wire f_s_dadda_pg_rca32_and_13_2_a_13;
  wire f_s_dadda_pg_rca32_and_13_2_b_2;
  wire f_s_dadda_pg_rca32_and_13_2_y0;
  wire f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_15_0_y0;
  wire f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_14_1_y0;
  wire f_s_dadda_pg_rca32_fa55_y0;
  wire f_s_dadda_pg_rca32_fa55_y1;
  wire f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_13_2_y0;
  wire f_s_dadda_pg_rca32_fa55_y2;
  wire f_s_dadda_pg_rca32_fa55_y3;
  wire f_s_dadda_pg_rca32_fa55_y4;
  wire f_s_dadda_pg_rca32_and_12_3_a_12;
  wire f_s_dadda_pg_rca32_and_12_3_b_3;
  wire f_s_dadda_pg_rca32_and_12_3_y0;
  wire f_s_dadda_pg_rca32_and_11_4_a_11;
  wire f_s_dadda_pg_rca32_and_11_4_b_4;
  wire f_s_dadda_pg_rca32_and_11_4_y0;
  wire f_s_dadda_pg_rca32_and_10_5_a_10;
  wire f_s_dadda_pg_rca32_and_10_5_b_5;
  wire f_s_dadda_pg_rca32_and_10_5_y0;
  wire f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_12_3_y0;
  wire f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_11_4_y0;
  wire f_s_dadda_pg_rca32_fa56_y0;
  wire f_s_dadda_pg_rca32_fa56_y1;
  wire f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_10_5_y0;
  wire f_s_dadda_pg_rca32_fa56_y2;
  wire f_s_dadda_pg_rca32_fa56_y3;
  wire f_s_dadda_pg_rca32_fa56_y4;
  wire f_s_dadda_pg_rca32_and_9_6_a_9;
  wire f_s_dadda_pg_rca32_and_9_6_b_6;
  wire f_s_dadda_pg_rca32_and_9_6_y0;
  wire f_s_dadda_pg_rca32_and_8_7_a_8;
  wire f_s_dadda_pg_rca32_and_8_7_b_7;
  wire f_s_dadda_pg_rca32_and_8_7_y0;
  wire f_s_dadda_pg_rca32_and_7_8_a_7;
  wire f_s_dadda_pg_rca32_and_7_8_b_8;
  wire f_s_dadda_pg_rca32_and_7_8_y0;
  wire f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_9_6_y0;
  wire f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_8_7_y0;
  wire f_s_dadda_pg_rca32_fa57_y0;
  wire f_s_dadda_pg_rca32_fa57_y1;
  wire f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_7_8_y0;
  wire f_s_dadda_pg_rca32_fa57_y2;
  wire f_s_dadda_pg_rca32_fa57_y3;
  wire f_s_dadda_pg_rca32_fa57_y4;
  wire f_s_dadda_pg_rca32_and_6_9_a_6;
  wire f_s_dadda_pg_rca32_and_6_9_b_9;
  wire f_s_dadda_pg_rca32_and_6_9_y0;
  wire f_s_dadda_pg_rca32_and_5_10_a_5;
  wire f_s_dadda_pg_rca32_and_5_10_b_10;
  wire f_s_dadda_pg_rca32_and_5_10_y0;
  wire f_s_dadda_pg_rca32_and_4_11_a_4;
  wire f_s_dadda_pg_rca32_and_4_11_b_11;
  wire f_s_dadda_pg_rca32_and_4_11_y0;
  wire f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_6_9_y0;
  wire f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_5_10_y0;
  wire f_s_dadda_pg_rca32_fa58_y0;
  wire f_s_dadda_pg_rca32_fa58_y1;
  wire f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_4_11_y0;
  wire f_s_dadda_pg_rca32_fa58_y2;
  wire f_s_dadda_pg_rca32_fa58_y3;
  wire f_s_dadda_pg_rca32_fa58_y4;
  wire f_s_dadda_pg_rca32_and_3_12_a_3;
  wire f_s_dadda_pg_rca32_and_3_12_b_12;
  wire f_s_dadda_pg_rca32_and_3_12_y0;
  wire f_s_dadda_pg_rca32_and_2_13_a_2;
  wire f_s_dadda_pg_rca32_and_2_13_b_13;
  wire f_s_dadda_pg_rca32_and_2_13_y0;
  wire f_s_dadda_pg_rca32_and_1_14_a_1;
  wire f_s_dadda_pg_rca32_and_1_14_b_14;
  wire f_s_dadda_pg_rca32_and_1_14_y0;
  wire f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_3_12_y0;
  wire f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_2_13_y0;
  wire f_s_dadda_pg_rca32_fa59_y0;
  wire f_s_dadda_pg_rca32_fa59_y1;
  wire f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_1_14_y0;
  wire f_s_dadda_pg_rca32_fa59_y2;
  wire f_s_dadda_pg_rca32_fa59_y3;
  wire f_s_dadda_pg_rca32_fa59_y4;
  wire f_s_dadda_pg_rca32_and_0_15_a_0;
  wire f_s_dadda_pg_rca32_and_0_15_b_15;
  wire f_s_dadda_pg_rca32_and_0_15_y0;
  wire f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_and_0_15_y0;
  wire f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_fa52_y2;
  wire f_s_dadda_pg_rca32_fa60_y0;
  wire f_s_dadda_pg_rca32_fa60_y1;
  wire f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_fa53_y2;
  wire f_s_dadda_pg_rca32_fa60_y2;
  wire f_s_dadda_pg_rca32_fa60_y3;
  wire f_s_dadda_pg_rca32_fa60_y4;
  wire f_s_dadda_pg_rca32_ha13_f_s_dadda_pg_rca32_fa54_y2;
  wire f_s_dadda_pg_rca32_ha13_f_s_dadda_pg_rca32_fa55_y2;
  wire f_s_dadda_pg_rca32_ha13_y0;
  wire f_s_dadda_pg_rca32_ha13_y1;
  wire f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_ha13_y1;
  wire f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_fa60_y4;
  wire f_s_dadda_pg_rca32_fa61_y0;
  wire f_s_dadda_pg_rca32_fa61_y1;
  wire f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_fa59_y4;
  wire f_s_dadda_pg_rca32_fa61_y2;
  wire f_s_dadda_pg_rca32_fa61_y3;
  wire f_s_dadda_pg_rca32_fa61_y4;
  wire f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa58_y4;
  wire f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa57_y4;
  wire f_s_dadda_pg_rca32_fa62_y0;
  wire f_s_dadda_pg_rca32_fa62_y1;
  wire f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa56_y4;
  wire f_s_dadda_pg_rca32_fa62_y2;
  wire f_s_dadda_pg_rca32_fa62_y3;
  wire f_s_dadda_pg_rca32_fa62_y4;
  wire f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa55_y4;
  wire f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa54_y4;
  wire f_s_dadda_pg_rca32_fa63_y0;
  wire f_s_dadda_pg_rca32_fa63_y1;
  wire f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa53_y4;
  wire f_s_dadda_pg_rca32_fa63_y2;
  wire f_s_dadda_pg_rca32_fa63_y3;
  wire f_s_dadda_pg_rca32_fa63_y4;
  wire f_s_dadda_pg_rca32_and_16_0_a_16;
  wire f_s_dadda_pg_rca32_and_16_0_b_0;
  wire f_s_dadda_pg_rca32_and_16_0_y0;
  wire f_s_dadda_pg_rca32_and_15_1_a_15;
  wire f_s_dadda_pg_rca32_and_15_1_b_1;
  wire f_s_dadda_pg_rca32_and_15_1_y0;
  wire f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_fa52_y4;
  wire f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_and_16_0_y0;
  wire f_s_dadda_pg_rca32_fa64_y0;
  wire f_s_dadda_pg_rca32_fa64_y1;
  wire f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_and_15_1_y0;
  wire f_s_dadda_pg_rca32_fa64_y2;
  wire f_s_dadda_pg_rca32_fa64_y3;
  wire f_s_dadda_pg_rca32_fa64_y4;
  wire f_s_dadda_pg_rca32_and_14_2_a_14;
  wire f_s_dadda_pg_rca32_and_14_2_b_2;
  wire f_s_dadda_pg_rca32_and_14_2_y0;
  wire f_s_dadda_pg_rca32_and_13_3_a_13;
  wire f_s_dadda_pg_rca32_and_13_3_b_3;
  wire f_s_dadda_pg_rca32_and_13_3_y0;
  wire f_s_dadda_pg_rca32_and_12_4_a_12;
  wire f_s_dadda_pg_rca32_and_12_4_b_4;
  wire f_s_dadda_pg_rca32_and_12_4_y0;
  wire f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_14_2_y0;
  wire f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_13_3_y0;
  wire f_s_dadda_pg_rca32_fa65_y0;
  wire f_s_dadda_pg_rca32_fa65_y1;
  wire f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_12_4_y0;
  wire f_s_dadda_pg_rca32_fa65_y2;
  wire f_s_dadda_pg_rca32_fa65_y3;
  wire f_s_dadda_pg_rca32_fa65_y4;
  wire f_s_dadda_pg_rca32_and_11_5_a_11;
  wire f_s_dadda_pg_rca32_and_11_5_b_5;
  wire f_s_dadda_pg_rca32_and_11_5_y0;
  wire f_s_dadda_pg_rca32_and_10_6_a_10;
  wire f_s_dadda_pg_rca32_and_10_6_b_6;
  wire f_s_dadda_pg_rca32_and_10_6_y0;
  wire f_s_dadda_pg_rca32_and_9_7_a_9;
  wire f_s_dadda_pg_rca32_and_9_7_b_7;
  wire f_s_dadda_pg_rca32_and_9_7_y0;
  wire f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_11_5_y0;
  wire f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_10_6_y0;
  wire f_s_dadda_pg_rca32_fa66_y0;
  wire f_s_dadda_pg_rca32_fa66_y1;
  wire f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_9_7_y0;
  wire f_s_dadda_pg_rca32_fa66_y2;
  wire f_s_dadda_pg_rca32_fa66_y3;
  wire f_s_dadda_pg_rca32_fa66_y4;
  wire f_s_dadda_pg_rca32_and_8_8_a_8;
  wire f_s_dadda_pg_rca32_and_8_8_b_8;
  wire f_s_dadda_pg_rca32_and_8_8_y0;
  wire f_s_dadda_pg_rca32_and_7_9_a_7;
  wire f_s_dadda_pg_rca32_and_7_9_b_9;
  wire f_s_dadda_pg_rca32_and_7_9_y0;
  wire f_s_dadda_pg_rca32_and_6_10_a_6;
  wire f_s_dadda_pg_rca32_and_6_10_b_10;
  wire f_s_dadda_pg_rca32_and_6_10_y0;
  wire f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_8_8_y0;
  wire f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_7_9_y0;
  wire f_s_dadda_pg_rca32_fa67_y0;
  wire f_s_dadda_pg_rca32_fa67_y1;
  wire f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_6_10_y0;
  wire f_s_dadda_pg_rca32_fa67_y2;
  wire f_s_dadda_pg_rca32_fa67_y3;
  wire f_s_dadda_pg_rca32_fa67_y4;
  wire f_s_dadda_pg_rca32_and_5_11_a_5;
  wire f_s_dadda_pg_rca32_and_5_11_b_11;
  wire f_s_dadda_pg_rca32_and_5_11_y0;
  wire f_s_dadda_pg_rca32_and_4_12_a_4;
  wire f_s_dadda_pg_rca32_and_4_12_b_12;
  wire f_s_dadda_pg_rca32_and_4_12_y0;
  wire f_s_dadda_pg_rca32_and_3_13_a_3;
  wire f_s_dadda_pg_rca32_and_3_13_b_13;
  wire f_s_dadda_pg_rca32_and_3_13_y0;
  wire f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_5_11_y0;
  wire f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_4_12_y0;
  wire f_s_dadda_pg_rca32_fa68_y0;
  wire f_s_dadda_pg_rca32_fa68_y1;
  wire f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_3_13_y0;
  wire f_s_dadda_pg_rca32_fa68_y2;
  wire f_s_dadda_pg_rca32_fa68_y3;
  wire f_s_dadda_pg_rca32_fa68_y4;
  wire f_s_dadda_pg_rca32_and_2_14_a_2;
  wire f_s_dadda_pg_rca32_and_2_14_b_14;
  wire f_s_dadda_pg_rca32_and_2_14_y0;
  wire f_s_dadda_pg_rca32_and_1_15_a_1;
  wire f_s_dadda_pg_rca32_and_1_15_b_15;
  wire f_s_dadda_pg_rca32_and_1_15_y0;
  wire f_s_dadda_pg_rca32_and_0_16_a_0;
  wire f_s_dadda_pg_rca32_and_0_16_b_16;
  wire f_s_dadda_pg_rca32_and_0_16_y0;
  wire f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_2_14_y0;
  wire f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_1_15_y0;
  wire f_s_dadda_pg_rca32_fa69_y0;
  wire f_s_dadda_pg_rca32_fa69_y1;
  wire f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_0_16_y0;
  wire f_s_dadda_pg_rca32_fa69_y2;
  wire f_s_dadda_pg_rca32_fa69_y3;
  wire f_s_dadda_pg_rca32_fa69_y4;
  wire f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa61_y2;
  wire f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa62_y2;
  wire f_s_dadda_pg_rca32_fa70_y0;
  wire f_s_dadda_pg_rca32_fa70_y1;
  wire f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa63_y2;
  wire f_s_dadda_pg_rca32_fa70_y2;
  wire f_s_dadda_pg_rca32_fa70_y3;
  wire f_s_dadda_pg_rca32_fa70_y4;
  wire f_s_dadda_pg_rca32_ha14_f_s_dadda_pg_rca32_fa64_y2;
  wire f_s_dadda_pg_rca32_ha14_f_s_dadda_pg_rca32_fa65_y2;
  wire f_s_dadda_pg_rca32_ha14_y0;
  wire f_s_dadda_pg_rca32_ha14_y1;
  wire f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_ha14_y1;
  wire f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_fa70_y4;
  wire f_s_dadda_pg_rca32_fa71_y0;
  wire f_s_dadda_pg_rca32_fa71_y1;
  wire f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_fa69_y4;
  wire f_s_dadda_pg_rca32_fa71_y2;
  wire f_s_dadda_pg_rca32_fa71_y3;
  wire f_s_dadda_pg_rca32_fa71_y4;
  wire f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa68_y4;
  wire f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa67_y4;
  wire f_s_dadda_pg_rca32_fa72_y0;
  wire f_s_dadda_pg_rca32_fa72_y1;
  wire f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa66_y4;
  wire f_s_dadda_pg_rca32_fa72_y2;
  wire f_s_dadda_pg_rca32_fa72_y3;
  wire f_s_dadda_pg_rca32_fa72_y4;
  wire f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa65_y4;
  wire f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa64_y4;
  wire f_s_dadda_pg_rca32_fa73_y0;
  wire f_s_dadda_pg_rca32_fa73_y1;
  wire f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa63_y4;
  wire f_s_dadda_pg_rca32_fa73_y2;
  wire f_s_dadda_pg_rca32_fa73_y3;
  wire f_s_dadda_pg_rca32_fa73_y4;
  wire f_s_dadda_pg_rca32_and_17_0_a_17;
  wire f_s_dadda_pg_rca32_and_17_0_b_0;
  wire f_s_dadda_pg_rca32_and_17_0_y0;
  wire f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_fa62_y4;
  wire f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_fa61_y4;
  wire f_s_dadda_pg_rca32_fa74_y0;
  wire f_s_dadda_pg_rca32_fa74_y1;
  wire f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_and_17_0_y0;
  wire f_s_dadda_pg_rca32_fa74_y2;
  wire f_s_dadda_pg_rca32_fa74_y3;
  wire f_s_dadda_pg_rca32_fa74_y4;
  wire f_s_dadda_pg_rca32_and_16_1_a_16;
  wire f_s_dadda_pg_rca32_and_16_1_b_1;
  wire f_s_dadda_pg_rca32_and_16_1_y0;
  wire f_s_dadda_pg_rca32_and_15_2_a_15;
  wire f_s_dadda_pg_rca32_and_15_2_b_2;
  wire f_s_dadda_pg_rca32_and_15_2_y0;
  wire f_s_dadda_pg_rca32_and_14_3_a_14;
  wire f_s_dadda_pg_rca32_and_14_3_b_3;
  wire f_s_dadda_pg_rca32_and_14_3_y0;
  wire f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_16_1_y0;
  wire f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_15_2_y0;
  wire f_s_dadda_pg_rca32_fa75_y0;
  wire f_s_dadda_pg_rca32_fa75_y1;
  wire f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_14_3_y0;
  wire f_s_dadda_pg_rca32_fa75_y2;
  wire f_s_dadda_pg_rca32_fa75_y3;
  wire f_s_dadda_pg_rca32_fa75_y4;
  wire f_s_dadda_pg_rca32_and_13_4_a_13;
  wire f_s_dadda_pg_rca32_and_13_4_b_4;
  wire f_s_dadda_pg_rca32_and_13_4_y0;
  wire f_s_dadda_pg_rca32_and_12_5_a_12;
  wire f_s_dadda_pg_rca32_and_12_5_b_5;
  wire f_s_dadda_pg_rca32_and_12_5_y0;
  wire f_s_dadda_pg_rca32_and_11_6_a_11;
  wire f_s_dadda_pg_rca32_and_11_6_b_6;
  wire f_s_dadda_pg_rca32_and_11_6_y0;
  wire f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_13_4_y0;
  wire f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_12_5_y0;
  wire f_s_dadda_pg_rca32_fa76_y0;
  wire f_s_dadda_pg_rca32_fa76_y1;
  wire f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_11_6_y0;
  wire f_s_dadda_pg_rca32_fa76_y2;
  wire f_s_dadda_pg_rca32_fa76_y3;
  wire f_s_dadda_pg_rca32_fa76_y4;
  wire f_s_dadda_pg_rca32_and_10_7_a_10;
  wire f_s_dadda_pg_rca32_and_10_7_b_7;
  wire f_s_dadda_pg_rca32_and_10_7_y0;
  wire f_s_dadda_pg_rca32_and_9_8_a_9;
  wire f_s_dadda_pg_rca32_and_9_8_b_8;
  wire f_s_dadda_pg_rca32_and_9_8_y0;
  wire f_s_dadda_pg_rca32_and_8_9_a_8;
  wire f_s_dadda_pg_rca32_and_8_9_b_9;
  wire f_s_dadda_pg_rca32_and_8_9_y0;
  wire f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_10_7_y0;
  wire f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_9_8_y0;
  wire f_s_dadda_pg_rca32_fa77_y0;
  wire f_s_dadda_pg_rca32_fa77_y1;
  wire f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_8_9_y0;
  wire f_s_dadda_pg_rca32_fa77_y2;
  wire f_s_dadda_pg_rca32_fa77_y3;
  wire f_s_dadda_pg_rca32_fa77_y4;
  wire f_s_dadda_pg_rca32_and_7_10_a_7;
  wire f_s_dadda_pg_rca32_and_7_10_b_10;
  wire f_s_dadda_pg_rca32_and_7_10_y0;
  wire f_s_dadda_pg_rca32_and_6_11_a_6;
  wire f_s_dadda_pg_rca32_and_6_11_b_11;
  wire f_s_dadda_pg_rca32_and_6_11_y0;
  wire f_s_dadda_pg_rca32_and_5_12_a_5;
  wire f_s_dadda_pg_rca32_and_5_12_b_12;
  wire f_s_dadda_pg_rca32_and_5_12_y0;
  wire f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_7_10_y0;
  wire f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_6_11_y0;
  wire f_s_dadda_pg_rca32_fa78_y0;
  wire f_s_dadda_pg_rca32_fa78_y1;
  wire f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_5_12_y0;
  wire f_s_dadda_pg_rca32_fa78_y2;
  wire f_s_dadda_pg_rca32_fa78_y3;
  wire f_s_dadda_pg_rca32_fa78_y4;
  wire f_s_dadda_pg_rca32_and_4_13_a_4;
  wire f_s_dadda_pg_rca32_and_4_13_b_13;
  wire f_s_dadda_pg_rca32_and_4_13_y0;
  wire f_s_dadda_pg_rca32_and_3_14_a_3;
  wire f_s_dadda_pg_rca32_and_3_14_b_14;
  wire f_s_dadda_pg_rca32_and_3_14_y0;
  wire f_s_dadda_pg_rca32_and_2_15_a_2;
  wire f_s_dadda_pg_rca32_and_2_15_b_15;
  wire f_s_dadda_pg_rca32_and_2_15_y0;
  wire f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_4_13_y0;
  wire f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_3_14_y0;
  wire f_s_dadda_pg_rca32_fa79_y0;
  wire f_s_dadda_pg_rca32_fa79_y1;
  wire f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_2_15_y0;
  wire f_s_dadda_pg_rca32_fa79_y2;
  wire f_s_dadda_pg_rca32_fa79_y3;
  wire f_s_dadda_pg_rca32_fa79_y4;
  wire f_s_dadda_pg_rca32_and_1_16_a_1;
  wire f_s_dadda_pg_rca32_and_1_16_b_16;
  wire f_s_dadda_pg_rca32_and_1_16_y0;
  wire f_s_dadda_pg_rca32_and_0_17_a_0;
  wire f_s_dadda_pg_rca32_and_0_17_b_17;
  wire f_s_dadda_pg_rca32_and_0_17_y0;
  wire f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_and_1_16_y0;
  wire f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_and_0_17_y0;
  wire f_s_dadda_pg_rca32_fa80_y0;
  wire f_s_dadda_pg_rca32_fa80_y1;
  wire f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_fa71_y2;
  wire f_s_dadda_pg_rca32_fa80_y2;
  wire f_s_dadda_pg_rca32_fa80_y3;
  wire f_s_dadda_pg_rca32_fa80_y4;
  wire f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa72_y2;
  wire f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa73_y2;
  wire f_s_dadda_pg_rca32_fa81_y0;
  wire f_s_dadda_pg_rca32_fa81_y1;
  wire f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa74_y2;
  wire f_s_dadda_pg_rca32_fa81_y2;
  wire f_s_dadda_pg_rca32_fa81_y3;
  wire f_s_dadda_pg_rca32_fa81_y4;
  wire f_s_dadda_pg_rca32_ha15_f_s_dadda_pg_rca32_fa75_y2;
  wire f_s_dadda_pg_rca32_ha15_f_s_dadda_pg_rca32_fa76_y2;
  wire f_s_dadda_pg_rca32_ha15_y0;
  wire f_s_dadda_pg_rca32_ha15_y1;
  wire f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_ha15_y1;
  wire f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_fa81_y4;
  wire f_s_dadda_pg_rca32_fa82_y0;
  wire f_s_dadda_pg_rca32_fa82_y1;
  wire f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_fa80_y4;
  wire f_s_dadda_pg_rca32_fa82_y2;
  wire f_s_dadda_pg_rca32_fa82_y3;
  wire f_s_dadda_pg_rca32_fa82_y4;
  wire f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa79_y4;
  wire f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa78_y4;
  wire f_s_dadda_pg_rca32_fa83_y0;
  wire f_s_dadda_pg_rca32_fa83_y1;
  wire f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa77_y4;
  wire f_s_dadda_pg_rca32_fa83_y2;
  wire f_s_dadda_pg_rca32_fa83_y3;
  wire f_s_dadda_pg_rca32_fa83_y4;
  wire f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa76_y4;
  wire f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa75_y4;
  wire f_s_dadda_pg_rca32_fa84_y0;
  wire f_s_dadda_pg_rca32_fa84_y1;
  wire f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa74_y4;
  wire f_s_dadda_pg_rca32_fa84_y2;
  wire f_s_dadda_pg_rca32_fa84_y3;
  wire f_s_dadda_pg_rca32_fa84_y4;
  wire f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa73_y4;
  wire f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa72_y4;
  wire f_s_dadda_pg_rca32_fa85_y0;
  wire f_s_dadda_pg_rca32_fa85_y1;
  wire f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa71_y4;
  wire f_s_dadda_pg_rca32_fa85_y2;
  wire f_s_dadda_pg_rca32_fa85_y3;
  wire f_s_dadda_pg_rca32_fa85_y4;
  wire f_s_dadda_pg_rca32_and_18_0_a_18;
  wire f_s_dadda_pg_rca32_and_18_0_b_0;
  wire f_s_dadda_pg_rca32_and_18_0_y0;
  wire f_s_dadda_pg_rca32_and_17_1_a_17;
  wire f_s_dadda_pg_rca32_and_17_1_b_1;
  wire f_s_dadda_pg_rca32_and_17_1_y0;
  wire f_s_dadda_pg_rca32_and_16_2_a_16;
  wire f_s_dadda_pg_rca32_and_16_2_b_2;
  wire f_s_dadda_pg_rca32_and_16_2_y0;
  wire f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_18_0_y0;
  wire f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_17_1_y0;
  wire f_s_dadda_pg_rca32_fa86_y0;
  wire f_s_dadda_pg_rca32_fa86_y1;
  wire f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_16_2_y0;
  wire f_s_dadda_pg_rca32_fa86_y2;
  wire f_s_dadda_pg_rca32_fa86_y3;
  wire f_s_dadda_pg_rca32_fa86_y4;
  wire f_s_dadda_pg_rca32_and_15_3_a_15;
  wire f_s_dadda_pg_rca32_and_15_3_b_3;
  wire f_s_dadda_pg_rca32_and_15_3_y0;
  wire f_s_dadda_pg_rca32_and_14_4_a_14;
  wire f_s_dadda_pg_rca32_and_14_4_b_4;
  wire f_s_dadda_pg_rca32_and_14_4_y0;
  wire f_s_dadda_pg_rca32_and_13_5_a_13;
  wire f_s_dadda_pg_rca32_and_13_5_b_5;
  wire f_s_dadda_pg_rca32_and_13_5_y0;
  wire f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_15_3_y0;
  wire f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_14_4_y0;
  wire f_s_dadda_pg_rca32_fa87_y0;
  wire f_s_dadda_pg_rca32_fa87_y1;
  wire f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_13_5_y0;
  wire f_s_dadda_pg_rca32_fa87_y2;
  wire f_s_dadda_pg_rca32_fa87_y3;
  wire f_s_dadda_pg_rca32_fa87_y4;
  wire f_s_dadda_pg_rca32_and_12_6_a_12;
  wire f_s_dadda_pg_rca32_and_12_6_b_6;
  wire f_s_dadda_pg_rca32_and_12_6_y0;
  wire f_s_dadda_pg_rca32_and_11_7_a_11;
  wire f_s_dadda_pg_rca32_and_11_7_b_7;
  wire f_s_dadda_pg_rca32_and_11_7_y0;
  wire f_s_dadda_pg_rca32_and_10_8_a_10;
  wire f_s_dadda_pg_rca32_and_10_8_b_8;
  wire f_s_dadda_pg_rca32_and_10_8_y0;
  wire f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_12_6_y0;
  wire f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_11_7_y0;
  wire f_s_dadda_pg_rca32_fa88_y0;
  wire f_s_dadda_pg_rca32_fa88_y1;
  wire f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_10_8_y0;
  wire f_s_dadda_pg_rca32_fa88_y2;
  wire f_s_dadda_pg_rca32_fa88_y3;
  wire f_s_dadda_pg_rca32_fa88_y4;
  wire f_s_dadda_pg_rca32_and_9_9_a_9;
  wire f_s_dadda_pg_rca32_and_9_9_b_9;
  wire f_s_dadda_pg_rca32_and_9_9_y0;
  wire f_s_dadda_pg_rca32_and_8_10_a_8;
  wire f_s_dadda_pg_rca32_and_8_10_b_10;
  wire f_s_dadda_pg_rca32_and_8_10_y0;
  wire f_s_dadda_pg_rca32_and_7_11_a_7;
  wire f_s_dadda_pg_rca32_and_7_11_b_11;
  wire f_s_dadda_pg_rca32_and_7_11_y0;
  wire f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_9_9_y0;
  wire f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_8_10_y0;
  wire f_s_dadda_pg_rca32_fa89_y0;
  wire f_s_dadda_pg_rca32_fa89_y1;
  wire f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_7_11_y0;
  wire f_s_dadda_pg_rca32_fa89_y2;
  wire f_s_dadda_pg_rca32_fa89_y3;
  wire f_s_dadda_pg_rca32_fa89_y4;
  wire f_s_dadda_pg_rca32_and_6_12_a_6;
  wire f_s_dadda_pg_rca32_and_6_12_b_12;
  wire f_s_dadda_pg_rca32_and_6_12_y0;
  wire f_s_dadda_pg_rca32_and_5_13_a_5;
  wire f_s_dadda_pg_rca32_and_5_13_b_13;
  wire f_s_dadda_pg_rca32_and_5_13_y0;
  wire f_s_dadda_pg_rca32_and_4_14_a_4;
  wire f_s_dadda_pg_rca32_and_4_14_b_14;
  wire f_s_dadda_pg_rca32_and_4_14_y0;
  wire f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_6_12_y0;
  wire f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_5_13_y0;
  wire f_s_dadda_pg_rca32_fa90_y0;
  wire f_s_dadda_pg_rca32_fa90_y1;
  wire f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_4_14_y0;
  wire f_s_dadda_pg_rca32_fa90_y2;
  wire f_s_dadda_pg_rca32_fa90_y3;
  wire f_s_dadda_pg_rca32_fa90_y4;
  wire f_s_dadda_pg_rca32_and_3_15_a_3;
  wire f_s_dadda_pg_rca32_and_3_15_b_15;
  wire f_s_dadda_pg_rca32_and_3_15_y0;
  wire f_s_dadda_pg_rca32_and_2_16_a_2;
  wire f_s_dadda_pg_rca32_and_2_16_b_16;
  wire f_s_dadda_pg_rca32_and_2_16_y0;
  wire f_s_dadda_pg_rca32_and_1_17_a_1;
  wire f_s_dadda_pg_rca32_and_1_17_b_17;
  wire f_s_dadda_pg_rca32_and_1_17_y0;
  wire f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_3_15_y0;
  wire f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_2_16_y0;
  wire f_s_dadda_pg_rca32_fa91_y0;
  wire f_s_dadda_pg_rca32_fa91_y1;
  wire f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_1_17_y0;
  wire f_s_dadda_pg_rca32_fa91_y2;
  wire f_s_dadda_pg_rca32_fa91_y3;
  wire f_s_dadda_pg_rca32_fa91_y4;
  wire f_s_dadda_pg_rca32_and_0_18_a_0;
  wire f_s_dadda_pg_rca32_and_0_18_b_18;
  wire f_s_dadda_pg_rca32_and_0_18_y0;
  wire f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_and_0_18_y0;
  wire f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_fa82_y2;
  wire f_s_dadda_pg_rca32_fa92_y0;
  wire f_s_dadda_pg_rca32_fa92_y1;
  wire f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_fa83_y2;
  wire f_s_dadda_pg_rca32_fa92_y2;
  wire f_s_dadda_pg_rca32_fa92_y3;
  wire f_s_dadda_pg_rca32_fa92_y4;
  wire f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa84_y2;
  wire f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa85_y2;
  wire f_s_dadda_pg_rca32_fa93_y0;
  wire f_s_dadda_pg_rca32_fa93_y1;
  wire f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa86_y2;
  wire f_s_dadda_pg_rca32_fa93_y2;
  wire f_s_dadda_pg_rca32_fa93_y3;
  wire f_s_dadda_pg_rca32_fa93_y4;
  wire f_s_dadda_pg_rca32_ha16_f_s_dadda_pg_rca32_fa87_y2;
  wire f_s_dadda_pg_rca32_ha16_f_s_dadda_pg_rca32_fa88_y2;
  wire f_s_dadda_pg_rca32_ha16_y0;
  wire f_s_dadda_pg_rca32_ha16_y1;
  wire f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_ha16_y1;
  wire f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_fa93_y4;
  wire f_s_dadda_pg_rca32_fa94_y0;
  wire f_s_dadda_pg_rca32_fa94_y1;
  wire f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_fa92_y4;
  wire f_s_dadda_pg_rca32_fa94_y2;
  wire f_s_dadda_pg_rca32_fa94_y3;
  wire f_s_dadda_pg_rca32_fa94_y4;
  wire f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa91_y4;
  wire f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa90_y4;
  wire f_s_dadda_pg_rca32_fa95_y0;
  wire f_s_dadda_pg_rca32_fa95_y1;
  wire f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa89_y4;
  wire f_s_dadda_pg_rca32_fa95_y2;
  wire f_s_dadda_pg_rca32_fa95_y3;
  wire f_s_dadda_pg_rca32_fa95_y4;
  wire f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa88_y4;
  wire f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa87_y4;
  wire f_s_dadda_pg_rca32_fa96_y0;
  wire f_s_dadda_pg_rca32_fa96_y1;
  wire f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa86_y4;
  wire f_s_dadda_pg_rca32_fa96_y2;
  wire f_s_dadda_pg_rca32_fa96_y3;
  wire f_s_dadda_pg_rca32_fa96_y4;
  wire f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa85_y4;
  wire f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa84_y4;
  wire f_s_dadda_pg_rca32_fa97_y0;
  wire f_s_dadda_pg_rca32_fa97_y1;
  wire f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa83_y4;
  wire f_s_dadda_pg_rca32_fa97_y2;
  wire f_s_dadda_pg_rca32_fa97_y3;
  wire f_s_dadda_pg_rca32_fa97_y4;
  wire f_s_dadda_pg_rca32_and_19_0_a_19;
  wire f_s_dadda_pg_rca32_and_19_0_b_0;
  wire f_s_dadda_pg_rca32_and_19_0_y0;
  wire f_s_dadda_pg_rca32_and_18_1_a_18;
  wire f_s_dadda_pg_rca32_and_18_1_b_1;
  wire f_s_dadda_pg_rca32_and_18_1_y0;
  wire f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_fa82_y4;
  wire f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_and_19_0_y0;
  wire f_s_dadda_pg_rca32_fa98_y0;
  wire f_s_dadda_pg_rca32_fa98_y1;
  wire f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_and_18_1_y0;
  wire f_s_dadda_pg_rca32_fa98_y2;
  wire f_s_dadda_pg_rca32_fa98_y3;
  wire f_s_dadda_pg_rca32_fa98_y4;
  wire f_s_dadda_pg_rca32_and_17_2_a_17;
  wire f_s_dadda_pg_rca32_and_17_2_b_2;
  wire f_s_dadda_pg_rca32_and_17_2_y0;
  wire f_s_dadda_pg_rca32_and_16_3_a_16;
  wire f_s_dadda_pg_rca32_and_16_3_b_3;
  wire f_s_dadda_pg_rca32_and_16_3_y0;
  wire f_s_dadda_pg_rca32_and_15_4_a_15;
  wire f_s_dadda_pg_rca32_and_15_4_b_4;
  wire f_s_dadda_pg_rca32_and_15_4_y0;
  wire f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_17_2_y0;
  wire f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_16_3_y0;
  wire f_s_dadda_pg_rca32_fa99_y0;
  wire f_s_dadda_pg_rca32_fa99_y1;
  wire f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_15_4_y0;
  wire f_s_dadda_pg_rca32_fa99_y2;
  wire f_s_dadda_pg_rca32_fa99_y3;
  wire f_s_dadda_pg_rca32_fa99_y4;
  wire f_s_dadda_pg_rca32_and_14_5_a_14;
  wire f_s_dadda_pg_rca32_and_14_5_b_5;
  wire f_s_dadda_pg_rca32_and_14_5_y0;
  wire f_s_dadda_pg_rca32_and_13_6_a_13;
  wire f_s_dadda_pg_rca32_and_13_6_b_6;
  wire f_s_dadda_pg_rca32_and_13_6_y0;
  wire f_s_dadda_pg_rca32_and_12_7_a_12;
  wire f_s_dadda_pg_rca32_and_12_7_b_7;
  wire f_s_dadda_pg_rca32_and_12_7_y0;
  wire f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_14_5_y0;
  wire f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_13_6_y0;
  wire f_s_dadda_pg_rca32_fa100_y0;
  wire f_s_dadda_pg_rca32_fa100_y1;
  wire f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_12_7_y0;
  wire f_s_dadda_pg_rca32_fa100_y2;
  wire f_s_dadda_pg_rca32_fa100_y3;
  wire f_s_dadda_pg_rca32_fa100_y4;
  wire f_s_dadda_pg_rca32_and_11_8_a_11;
  wire f_s_dadda_pg_rca32_and_11_8_b_8;
  wire f_s_dadda_pg_rca32_and_11_8_y0;
  wire f_s_dadda_pg_rca32_and_10_9_a_10;
  wire f_s_dadda_pg_rca32_and_10_9_b_9;
  wire f_s_dadda_pg_rca32_and_10_9_y0;
  wire f_s_dadda_pg_rca32_and_9_10_a_9;
  wire f_s_dadda_pg_rca32_and_9_10_b_10;
  wire f_s_dadda_pg_rca32_and_9_10_y0;
  wire f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_11_8_y0;
  wire f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_10_9_y0;
  wire f_s_dadda_pg_rca32_fa101_y0;
  wire f_s_dadda_pg_rca32_fa101_y1;
  wire f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_9_10_y0;
  wire f_s_dadda_pg_rca32_fa101_y2;
  wire f_s_dadda_pg_rca32_fa101_y3;
  wire f_s_dadda_pg_rca32_fa101_y4;
  wire f_s_dadda_pg_rca32_and_8_11_a_8;
  wire f_s_dadda_pg_rca32_and_8_11_b_11;
  wire f_s_dadda_pg_rca32_and_8_11_y0;
  wire f_s_dadda_pg_rca32_and_7_12_a_7;
  wire f_s_dadda_pg_rca32_and_7_12_b_12;
  wire f_s_dadda_pg_rca32_and_7_12_y0;
  wire f_s_dadda_pg_rca32_and_6_13_a_6;
  wire f_s_dadda_pg_rca32_and_6_13_b_13;
  wire f_s_dadda_pg_rca32_and_6_13_y0;
  wire f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_8_11_y0;
  wire f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_7_12_y0;
  wire f_s_dadda_pg_rca32_fa102_y0;
  wire f_s_dadda_pg_rca32_fa102_y1;
  wire f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_6_13_y0;
  wire f_s_dadda_pg_rca32_fa102_y2;
  wire f_s_dadda_pg_rca32_fa102_y3;
  wire f_s_dadda_pg_rca32_fa102_y4;
  wire f_s_dadda_pg_rca32_and_5_14_a_5;
  wire f_s_dadda_pg_rca32_and_5_14_b_14;
  wire f_s_dadda_pg_rca32_and_5_14_y0;
  wire f_s_dadda_pg_rca32_and_4_15_a_4;
  wire f_s_dadda_pg_rca32_and_4_15_b_15;
  wire f_s_dadda_pg_rca32_and_4_15_y0;
  wire f_s_dadda_pg_rca32_and_3_16_a_3;
  wire f_s_dadda_pg_rca32_and_3_16_b_16;
  wire f_s_dadda_pg_rca32_and_3_16_y0;
  wire f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_5_14_y0;
  wire f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_4_15_y0;
  wire f_s_dadda_pg_rca32_fa103_y0;
  wire f_s_dadda_pg_rca32_fa103_y1;
  wire f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_3_16_y0;
  wire f_s_dadda_pg_rca32_fa103_y2;
  wire f_s_dadda_pg_rca32_fa103_y3;
  wire f_s_dadda_pg_rca32_fa103_y4;
  wire f_s_dadda_pg_rca32_and_2_17_a_2;
  wire f_s_dadda_pg_rca32_and_2_17_b_17;
  wire f_s_dadda_pg_rca32_and_2_17_y0;
  wire f_s_dadda_pg_rca32_and_1_18_a_1;
  wire f_s_dadda_pg_rca32_and_1_18_b_18;
  wire f_s_dadda_pg_rca32_and_1_18_y0;
  wire f_s_dadda_pg_rca32_and_0_19_a_0;
  wire f_s_dadda_pg_rca32_and_0_19_b_19;
  wire f_s_dadda_pg_rca32_and_0_19_y0;
  wire f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_2_17_y0;
  wire f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_1_18_y0;
  wire f_s_dadda_pg_rca32_fa104_y0;
  wire f_s_dadda_pg_rca32_fa104_y1;
  wire f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_0_19_y0;
  wire f_s_dadda_pg_rca32_fa104_y2;
  wire f_s_dadda_pg_rca32_fa104_y3;
  wire f_s_dadda_pg_rca32_fa104_y4;
  wire f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa94_y2;
  wire f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa95_y2;
  wire f_s_dadda_pg_rca32_fa105_y0;
  wire f_s_dadda_pg_rca32_fa105_y1;
  wire f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa96_y2;
  wire f_s_dadda_pg_rca32_fa105_y2;
  wire f_s_dadda_pg_rca32_fa105_y3;
  wire f_s_dadda_pg_rca32_fa105_y4;
  wire f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa97_y2;
  wire f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa98_y2;
  wire f_s_dadda_pg_rca32_fa106_y0;
  wire f_s_dadda_pg_rca32_fa106_y1;
  wire f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa99_y2;
  wire f_s_dadda_pg_rca32_fa106_y2;
  wire f_s_dadda_pg_rca32_fa106_y3;
  wire f_s_dadda_pg_rca32_fa106_y4;
  wire f_s_dadda_pg_rca32_ha17_f_s_dadda_pg_rca32_fa100_y2;
  wire f_s_dadda_pg_rca32_ha17_f_s_dadda_pg_rca32_fa101_y2;
  wire f_s_dadda_pg_rca32_ha17_y0;
  wire f_s_dadda_pg_rca32_ha17_y1;
  wire f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_ha17_y1;
  wire f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_fa106_y4;
  wire f_s_dadda_pg_rca32_fa107_y0;
  wire f_s_dadda_pg_rca32_fa107_y1;
  wire f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_fa105_y4;
  wire f_s_dadda_pg_rca32_fa107_y2;
  wire f_s_dadda_pg_rca32_fa107_y3;
  wire f_s_dadda_pg_rca32_fa107_y4;
  wire f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa104_y4;
  wire f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa103_y4;
  wire f_s_dadda_pg_rca32_fa108_y0;
  wire f_s_dadda_pg_rca32_fa108_y1;
  wire f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa102_y4;
  wire f_s_dadda_pg_rca32_fa108_y2;
  wire f_s_dadda_pg_rca32_fa108_y3;
  wire f_s_dadda_pg_rca32_fa108_y4;
  wire f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa101_y4;
  wire f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa100_y4;
  wire f_s_dadda_pg_rca32_fa109_y0;
  wire f_s_dadda_pg_rca32_fa109_y1;
  wire f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa99_y4;
  wire f_s_dadda_pg_rca32_fa109_y2;
  wire f_s_dadda_pg_rca32_fa109_y3;
  wire f_s_dadda_pg_rca32_fa109_y4;
  wire f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa98_y4;
  wire f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa97_y4;
  wire f_s_dadda_pg_rca32_fa110_y0;
  wire f_s_dadda_pg_rca32_fa110_y1;
  wire f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa96_y4;
  wire f_s_dadda_pg_rca32_fa110_y2;
  wire f_s_dadda_pg_rca32_fa110_y3;
  wire f_s_dadda_pg_rca32_fa110_y4;
  wire f_s_dadda_pg_rca32_and_20_0_a_20;
  wire f_s_dadda_pg_rca32_and_20_0_b_0;
  wire f_s_dadda_pg_rca32_and_20_0_y0;
  wire f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_fa95_y4;
  wire f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_fa94_y4;
  wire f_s_dadda_pg_rca32_fa111_y0;
  wire f_s_dadda_pg_rca32_fa111_y1;
  wire f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_and_20_0_y0;
  wire f_s_dadda_pg_rca32_fa111_y2;
  wire f_s_dadda_pg_rca32_fa111_y3;
  wire f_s_dadda_pg_rca32_fa111_y4;
  wire f_s_dadda_pg_rca32_and_19_1_a_19;
  wire f_s_dadda_pg_rca32_and_19_1_b_1;
  wire f_s_dadda_pg_rca32_and_19_1_y0;
  wire f_s_dadda_pg_rca32_and_18_2_a_18;
  wire f_s_dadda_pg_rca32_and_18_2_b_2;
  wire f_s_dadda_pg_rca32_and_18_2_y0;
  wire f_s_dadda_pg_rca32_and_17_3_a_17;
  wire f_s_dadda_pg_rca32_and_17_3_b_3;
  wire f_s_dadda_pg_rca32_and_17_3_y0;
  wire f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_19_1_y0;
  wire f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_18_2_y0;
  wire f_s_dadda_pg_rca32_fa112_y0;
  wire f_s_dadda_pg_rca32_fa112_y1;
  wire f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_17_3_y0;
  wire f_s_dadda_pg_rca32_fa112_y2;
  wire f_s_dadda_pg_rca32_fa112_y3;
  wire f_s_dadda_pg_rca32_fa112_y4;
  wire f_s_dadda_pg_rca32_and_16_4_a_16;
  wire f_s_dadda_pg_rca32_and_16_4_b_4;
  wire f_s_dadda_pg_rca32_and_16_4_y0;
  wire f_s_dadda_pg_rca32_and_15_5_a_15;
  wire f_s_dadda_pg_rca32_and_15_5_b_5;
  wire f_s_dadda_pg_rca32_and_15_5_y0;
  wire f_s_dadda_pg_rca32_and_14_6_a_14;
  wire f_s_dadda_pg_rca32_and_14_6_b_6;
  wire f_s_dadda_pg_rca32_and_14_6_y0;
  wire f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_16_4_y0;
  wire f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_15_5_y0;
  wire f_s_dadda_pg_rca32_fa113_y0;
  wire f_s_dadda_pg_rca32_fa113_y1;
  wire f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_14_6_y0;
  wire f_s_dadda_pg_rca32_fa113_y2;
  wire f_s_dadda_pg_rca32_fa113_y3;
  wire f_s_dadda_pg_rca32_fa113_y4;
  wire f_s_dadda_pg_rca32_and_13_7_a_13;
  wire f_s_dadda_pg_rca32_and_13_7_b_7;
  wire f_s_dadda_pg_rca32_and_13_7_y0;
  wire f_s_dadda_pg_rca32_and_12_8_a_12;
  wire f_s_dadda_pg_rca32_and_12_8_b_8;
  wire f_s_dadda_pg_rca32_and_12_8_y0;
  wire f_s_dadda_pg_rca32_and_11_9_a_11;
  wire f_s_dadda_pg_rca32_and_11_9_b_9;
  wire f_s_dadda_pg_rca32_and_11_9_y0;
  wire f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_13_7_y0;
  wire f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_12_8_y0;
  wire f_s_dadda_pg_rca32_fa114_y0;
  wire f_s_dadda_pg_rca32_fa114_y1;
  wire f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_11_9_y0;
  wire f_s_dadda_pg_rca32_fa114_y2;
  wire f_s_dadda_pg_rca32_fa114_y3;
  wire f_s_dadda_pg_rca32_fa114_y4;
  wire f_s_dadda_pg_rca32_and_10_10_a_10;
  wire f_s_dadda_pg_rca32_and_10_10_b_10;
  wire f_s_dadda_pg_rca32_and_10_10_y0;
  wire f_s_dadda_pg_rca32_and_9_11_a_9;
  wire f_s_dadda_pg_rca32_and_9_11_b_11;
  wire f_s_dadda_pg_rca32_and_9_11_y0;
  wire f_s_dadda_pg_rca32_and_8_12_a_8;
  wire f_s_dadda_pg_rca32_and_8_12_b_12;
  wire f_s_dadda_pg_rca32_and_8_12_y0;
  wire f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_10_10_y0;
  wire f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_9_11_y0;
  wire f_s_dadda_pg_rca32_fa115_y0;
  wire f_s_dadda_pg_rca32_fa115_y1;
  wire f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_8_12_y0;
  wire f_s_dadda_pg_rca32_fa115_y2;
  wire f_s_dadda_pg_rca32_fa115_y3;
  wire f_s_dadda_pg_rca32_fa115_y4;
  wire f_s_dadda_pg_rca32_and_7_13_a_7;
  wire f_s_dadda_pg_rca32_and_7_13_b_13;
  wire f_s_dadda_pg_rca32_and_7_13_y0;
  wire f_s_dadda_pg_rca32_and_6_14_a_6;
  wire f_s_dadda_pg_rca32_and_6_14_b_14;
  wire f_s_dadda_pg_rca32_and_6_14_y0;
  wire f_s_dadda_pg_rca32_and_5_15_a_5;
  wire f_s_dadda_pg_rca32_and_5_15_b_15;
  wire f_s_dadda_pg_rca32_and_5_15_y0;
  wire f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_7_13_y0;
  wire f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_6_14_y0;
  wire f_s_dadda_pg_rca32_fa116_y0;
  wire f_s_dadda_pg_rca32_fa116_y1;
  wire f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_5_15_y0;
  wire f_s_dadda_pg_rca32_fa116_y2;
  wire f_s_dadda_pg_rca32_fa116_y3;
  wire f_s_dadda_pg_rca32_fa116_y4;
  wire f_s_dadda_pg_rca32_and_4_16_a_4;
  wire f_s_dadda_pg_rca32_and_4_16_b_16;
  wire f_s_dadda_pg_rca32_and_4_16_y0;
  wire f_s_dadda_pg_rca32_and_3_17_a_3;
  wire f_s_dadda_pg_rca32_and_3_17_b_17;
  wire f_s_dadda_pg_rca32_and_3_17_y0;
  wire f_s_dadda_pg_rca32_and_2_18_a_2;
  wire f_s_dadda_pg_rca32_and_2_18_b_18;
  wire f_s_dadda_pg_rca32_and_2_18_y0;
  wire f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_4_16_y0;
  wire f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_3_17_y0;
  wire f_s_dadda_pg_rca32_fa117_y0;
  wire f_s_dadda_pg_rca32_fa117_y1;
  wire f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_2_18_y0;
  wire f_s_dadda_pg_rca32_fa117_y2;
  wire f_s_dadda_pg_rca32_fa117_y3;
  wire f_s_dadda_pg_rca32_fa117_y4;
  wire f_s_dadda_pg_rca32_and_1_19_a_1;
  wire f_s_dadda_pg_rca32_and_1_19_b_19;
  wire f_s_dadda_pg_rca32_and_1_19_y0;
  wire f_s_dadda_pg_rca32_and_0_20_a_0;
  wire f_s_dadda_pg_rca32_and_0_20_b_20;
  wire f_s_dadda_pg_rca32_and_0_20_y0;
  wire f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_and_1_19_y0;
  wire f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_and_0_20_y0;
  wire f_s_dadda_pg_rca32_fa118_y0;
  wire f_s_dadda_pg_rca32_fa118_y1;
  wire f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_fa107_y2;
  wire f_s_dadda_pg_rca32_fa118_y2;
  wire f_s_dadda_pg_rca32_fa118_y3;
  wire f_s_dadda_pg_rca32_fa118_y4;
  wire f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa108_y2;
  wire f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa109_y2;
  wire f_s_dadda_pg_rca32_fa119_y0;
  wire f_s_dadda_pg_rca32_fa119_y1;
  wire f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa110_y2;
  wire f_s_dadda_pg_rca32_fa119_y2;
  wire f_s_dadda_pg_rca32_fa119_y3;
  wire f_s_dadda_pg_rca32_fa119_y4;
  wire f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa111_y2;
  wire f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa112_y2;
  wire f_s_dadda_pg_rca32_fa120_y0;
  wire f_s_dadda_pg_rca32_fa120_y1;
  wire f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa113_y2;
  wire f_s_dadda_pg_rca32_fa120_y2;
  wire f_s_dadda_pg_rca32_fa120_y3;
  wire f_s_dadda_pg_rca32_fa120_y4;
  wire f_s_dadda_pg_rca32_ha18_f_s_dadda_pg_rca32_fa114_y2;
  wire f_s_dadda_pg_rca32_ha18_f_s_dadda_pg_rca32_fa115_y2;
  wire f_s_dadda_pg_rca32_ha18_y0;
  wire f_s_dadda_pg_rca32_ha18_y1;
  wire f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_ha18_y1;
  wire f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_fa120_y4;
  wire f_s_dadda_pg_rca32_fa121_y0;
  wire f_s_dadda_pg_rca32_fa121_y1;
  wire f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_fa119_y4;
  wire f_s_dadda_pg_rca32_fa121_y2;
  wire f_s_dadda_pg_rca32_fa121_y3;
  wire f_s_dadda_pg_rca32_fa121_y4;
  wire f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa118_y4;
  wire f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa117_y4;
  wire f_s_dadda_pg_rca32_fa122_y0;
  wire f_s_dadda_pg_rca32_fa122_y1;
  wire f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa116_y4;
  wire f_s_dadda_pg_rca32_fa122_y2;
  wire f_s_dadda_pg_rca32_fa122_y3;
  wire f_s_dadda_pg_rca32_fa122_y4;
  wire f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa115_y4;
  wire f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa114_y4;
  wire f_s_dadda_pg_rca32_fa123_y0;
  wire f_s_dadda_pg_rca32_fa123_y1;
  wire f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa113_y4;
  wire f_s_dadda_pg_rca32_fa123_y2;
  wire f_s_dadda_pg_rca32_fa123_y3;
  wire f_s_dadda_pg_rca32_fa123_y4;
  wire f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa112_y4;
  wire f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa111_y4;
  wire f_s_dadda_pg_rca32_fa124_y0;
  wire f_s_dadda_pg_rca32_fa124_y1;
  wire f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa110_y4;
  wire f_s_dadda_pg_rca32_fa124_y2;
  wire f_s_dadda_pg_rca32_fa124_y3;
  wire f_s_dadda_pg_rca32_fa124_y4;
  wire f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa109_y4;
  wire f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa108_y4;
  wire f_s_dadda_pg_rca32_fa125_y0;
  wire f_s_dadda_pg_rca32_fa125_y1;
  wire f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa107_y4;
  wire f_s_dadda_pg_rca32_fa125_y2;
  wire f_s_dadda_pg_rca32_fa125_y3;
  wire f_s_dadda_pg_rca32_fa125_y4;
  wire f_s_dadda_pg_rca32_and_21_0_a_21;
  wire f_s_dadda_pg_rca32_and_21_0_b_0;
  wire f_s_dadda_pg_rca32_and_21_0_y0;
  wire f_s_dadda_pg_rca32_and_20_1_a_20;
  wire f_s_dadda_pg_rca32_and_20_1_b_1;
  wire f_s_dadda_pg_rca32_and_20_1_y0;
  wire f_s_dadda_pg_rca32_and_19_2_a_19;
  wire f_s_dadda_pg_rca32_and_19_2_b_2;
  wire f_s_dadda_pg_rca32_and_19_2_y0;
  wire f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_21_0_y0;
  wire f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_20_1_y0;
  wire f_s_dadda_pg_rca32_fa126_y0;
  wire f_s_dadda_pg_rca32_fa126_y1;
  wire f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_19_2_y0;
  wire f_s_dadda_pg_rca32_fa126_y2;
  wire f_s_dadda_pg_rca32_fa126_y3;
  wire f_s_dadda_pg_rca32_fa126_y4;
  wire f_s_dadda_pg_rca32_and_18_3_a_18;
  wire f_s_dadda_pg_rca32_and_18_3_b_3;
  wire f_s_dadda_pg_rca32_and_18_3_y0;
  wire f_s_dadda_pg_rca32_and_17_4_a_17;
  wire f_s_dadda_pg_rca32_and_17_4_b_4;
  wire f_s_dadda_pg_rca32_and_17_4_y0;
  wire f_s_dadda_pg_rca32_and_16_5_a_16;
  wire f_s_dadda_pg_rca32_and_16_5_b_5;
  wire f_s_dadda_pg_rca32_and_16_5_y0;
  wire f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_18_3_y0;
  wire f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_17_4_y0;
  wire f_s_dadda_pg_rca32_fa127_y0;
  wire f_s_dadda_pg_rca32_fa127_y1;
  wire f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_16_5_y0;
  wire f_s_dadda_pg_rca32_fa127_y2;
  wire f_s_dadda_pg_rca32_fa127_y3;
  wire f_s_dadda_pg_rca32_fa127_y4;
  wire f_s_dadda_pg_rca32_and_15_6_a_15;
  wire f_s_dadda_pg_rca32_and_15_6_b_6;
  wire f_s_dadda_pg_rca32_and_15_6_y0;
  wire f_s_dadda_pg_rca32_and_14_7_a_14;
  wire f_s_dadda_pg_rca32_and_14_7_b_7;
  wire f_s_dadda_pg_rca32_and_14_7_y0;
  wire f_s_dadda_pg_rca32_and_13_8_a_13;
  wire f_s_dadda_pg_rca32_and_13_8_b_8;
  wire f_s_dadda_pg_rca32_and_13_8_y0;
  wire f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_15_6_y0;
  wire f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_14_7_y0;
  wire f_s_dadda_pg_rca32_fa128_y0;
  wire f_s_dadda_pg_rca32_fa128_y1;
  wire f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_13_8_y0;
  wire f_s_dadda_pg_rca32_fa128_y2;
  wire f_s_dadda_pg_rca32_fa128_y3;
  wire f_s_dadda_pg_rca32_fa128_y4;
  wire f_s_dadda_pg_rca32_and_12_9_a_12;
  wire f_s_dadda_pg_rca32_and_12_9_b_9;
  wire f_s_dadda_pg_rca32_and_12_9_y0;
  wire f_s_dadda_pg_rca32_and_11_10_a_11;
  wire f_s_dadda_pg_rca32_and_11_10_b_10;
  wire f_s_dadda_pg_rca32_and_11_10_y0;
  wire f_s_dadda_pg_rca32_and_10_11_a_10;
  wire f_s_dadda_pg_rca32_and_10_11_b_11;
  wire f_s_dadda_pg_rca32_and_10_11_y0;
  wire f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_12_9_y0;
  wire f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_11_10_y0;
  wire f_s_dadda_pg_rca32_fa129_y0;
  wire f_s_dadda_pg_rca32_fa129_y1;
  wire f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_10_11_y0;
  wire f_s_dadda_pg_rca32_fa129_y2;
  wire f_s_dadda_pg_rca32_fa129_y3;
  wire f_s_dadda_pg_rca32_fa129_y4;
  wire f_s_dadda_pg_rca32_and_9_12_a_9;
  wire f_s_dadda_pg_rca32_and_9_12_b_12;
  wire f_s_dadda_pg_rca32_and_9_12_y0;
  wire f_s_dadda_pg_rca32_and_8_13_a_8;
  wire f_s_dadda_pg_rca32_and_8_13_b_13;
  wire f_s_dadda_pg_rca32_and_8_13_y0;
  wire f_s_dadda_pg_rca32_and_7_14_a_7;
  wire f_s_dadda_pg_rca32_and_7_14_b_14;
  wire f_s_dadda_pg_rca32_and_7_14_y0;
  wire f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_9_12_y0;
  wire f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_8_13_y0;
  wire f_s_dadda_pg_rca32_fa130_y0;
  wire f_s_dadda_pg_rca32_fa130_y1;
  wire f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_7_14_y0;
  wire f_s_dadda_pg_rca32_fa130_y2;
  wire f_s_dadda_pg_rca32_fa130_y3;
  wire f_s_dadda_pg_rca32_fa130_y4;
  wire f_s_dadda_pg_rca32_and_6_15_a_6;
  wire f_s_dadda_pg_rca32_and_6_15_b_15;
  wire f_s_dadda_pg_rca32_and_6_15_y0;
  wire f_s_dadda_pg_rca32_and_5_16_a_5;
  wire f_s_dadda_pg_rca32_and_5_16_b_16;
  wire f_s_dadda_pg_rca32_and_5_16_y0;
  wire f_s_dadda_pg_rca32_and_4_17_a_4;
  wire f_s_dadda_pg_rca32_and_4_17_b_17;
  wire f_s_dadda_pg_rca32_and_4_17_y0;
  wire f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_6_15_y0;
  wire f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_5_16_y0;
  wire f_s_dadda_pg_rca32_fa131_y0;
  wire f_s_dadda_pg_rca32_fa131_y1;
  wire f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_4_17_y0;
  wire f_s_dadda_pg_rca32_fa131_y2;
  wire f_s_dadda_pg_rca32_fa131_y3;
  wire f_s_dadda_pg_rca32_fa131_y4;
  wire f_s_dadda_pg_rca32_and_3_18_a_3;
  wire f_s_dadda_pg_rca32_and_3_18_b_18;
  wire f_s_dadda_pg_rca32_and_3_18_y0;
  wire f_s_dadda_pg_rca32_and_2_19_a_2;
  wire f_s_dadda_pg_rca32_and_2_19_b_19;
  wire f_s_dadda_pg_rca32_and_2_19_y0;
  wire f_s_dadda_pg_rca32_and_1_20_a_1;
  wire f_s_dadda_pg_rca32_and_1_20_b_20;
  wire f_s_dadda_pg_rca32_and_1_20_y0;
  wire f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_3_18_y0;
  wire f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_2_19_y0;
  wire f_s_dadda_pg_rca32_fa132_y0;
  wire f_s_dadda_pg_rca32_fa132_y1;
  wire f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_1_20_y0;
  wire f_s_dadda_pg_rca32_fa132_y2;
  wire f_s_dadda_pg_rca32_fa132_y3;
  wire f_s_dadda_pg_rca32_fa132_y4;
  wire f_s_dadda_pg_rca32_and_0_21_a_0;
  wire f_s_dadda_pg_rca32_and_0_21_b_21;
  wire f_s_dadda_pg_rca32_and_0_21_y0;
  wire f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_and_0_21_y0;
  wire f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_fa121_y2;
  wire f_s_dadda_pg_rca32_fa133_y0;
  wire f_s_dadda_pg_rca32_fa133_y1;
  wire f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_fa122_y2;
  wire f_s_dadda_pg_rca32_fa133_y2;
  wire f_s_dadda_pg_rca32_fa133_y3;
  wire f_s_dadda_pg_rca32_fa133_y4;
  wire f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa123_y2;
  wire f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa124_y2;
  wire f_s_dadda_pg_rca32_fa134_y0;
  wire f_s_dadda_pg_rca32_fa134_y1;
  wire f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa125_y2;
  wire f_s_dadda_pg_rca32_fa134_y2;
  wire f_s_dadda_pg_rca32_fa134_y3;
  wire f_s_dadda_pg_rca32_fa134_y4;
  wire f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa126_y2;
  wire f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa127_y2;
  wire f_s_dadda_pg_rca32_fa135_y0;
  wire f_s_dadda_pg_rca32_fa135_y1;
  wire f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa128_y2;
  wire f_s_dadda_pg_rca32_fa135_y2;
  wire f_s_dadda_pg_rca32_fa135_y3;
  wire f_s_dadda_pg_rca32_fa135_y4;
  wire f_s_dadda_pg_rca32_ha19_f_s_dadda_pg_rca32_fa129_y2;
  wire f_s_dadda_pg_rca32_ha19_f_s_dadda_pg_rca32_fa130_y2;
  wire f_s_dadda_pg_rca32_ha19_y0;
  wire f_s_dadda_pg_rca32_ha19_y1;
  wire f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_ha19_y1;
  wire f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_fa135_y4;
  wire f_s_dadda_pg_rca32_fa136_y0;
  wire f_s_dadda_pg_rca32_fa136_y1;
  wire f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_fa134_y4;
  wire f_s_dadda_pg_rca32_fa136_y2;
  wire f_s_dadda_pg_rca32_fa136_y3;
  wire f_s_dadda_pg_rca32_fa136_y4;
  wire f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa133_y4;
  wire f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa132_y4;
  wire f_s_dadda_pg_rca32_fa137_y0;
  wire f_s_dadda_pg_rca32_fa137_y1;
  wire f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa131_y4;
  wire f_s_dadda_pg_rca32_fa137_y2;
  wire f_s_dadda_pg_rca32_fa137_y3;
  wire f_s_dadda_pg_rca32_fa137_y4;
  wire f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa130_y4;
  wire f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa129_y4;
  wire f_s_dadda_pg_rca32_fa138_y0;
  wire f_s_dadda_pg_rca32_fa138_y1;
  wire f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa128_y4;
  wire f_s_dadda_pg_rca32_fa138_y2;
  wire f_s_dadda_pg_rca32_fa138_y3;
  wire f_s_dadda_pg_rca32_fa138_y4;
  wire f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa127_y4;
  wire f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa126_y4;
  wire f_s_dadda_pg_rca32_fa139_y0;
  wire f_s_dadda_pg_rca32_fa139_y1;
  wire f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa125_y4;
  wire f_s_dadda_pg_rca32_fa139_y2;
  wire f_s_dadda_pg_rca32_fa139_y3;
  wire f_s_dadda_pg_rca32_fa139_y4;
  wire f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa124_y4;
  wire f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa123_y4;
  wire f_s_dadda_pg_rca32_fa140_y0;
  wire f_s_dadda_pg_rca32_fa140_y1;
  wire f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa122_y4;
  wire f_s_dadda_pg_rca32_fa140_y2;
  wire f_s_dadda_pg_rca32_fa140_y3;
  wire f_s_dadda_pg_rca32_fa140_y4;
  wire f_s_dadda_pg_rca32_and_22_0_a_22;
  wire f_s_dadda_pg_rca32_and_22_0_b_0;
  wire f_s_dadda_pg_rca32_and_22_0_y0;
  wire f_s_dadda_pg_rca32_and_21_1_a_21;
  wire f_s_dadda_pg_rca32_and_21_1_b_1;
  wire f_s_dadda_pg_rca32_and_21_1_y0;
  wire f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_fa121_y4;
  wire f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_and_22_0_y0;
  wire f_s_dadda_pg_rca32_fa141_y0;
  wire f_s_dadda_pg_rca32_fa141_y1;
  wire f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_and_21_1_y0;
  wire f_s_dadda_pg_rca32_fa141_y2;
  wire f_s_dadda_pg_rca32_fa141_y3;
  wire f_s_dadda_pg_rca32_fa141_y4;
  wire f_s_dadda_pg_rca32_and_20_2_a_20;
  wire f_s_dadda_pg_rca32_and_20_2_b_2;
  wire f_s_dadda_pg_rca32_and_20_2_y0;
  wire f_s_dadda_pg_rca32_and_19_3_a_19;
  wire f_s_dadda_pg_rca32_and_19_3_b_3;
  wire f_s_dadda_pg_rca32_and_19_3_y0;
  wire f_s_dadda_pg_rca32_and_18_4_a_18;
  wire f_s_dadda_pg_rca32_and_18_4_b_4;
  wire f_s_dadda_pg_rca32_and_18_4_y0;
  wire f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_20_2_y0;
  wire f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_19_3_y0;
  wire f_s_dadda_pg_rca32_fa142_y0;
  wire f_s_dadda_pg_rca32_fa142_y1;
  wire f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_18_4_y0;
  wire f_s_dadda_pg_rca32_fa142_y2;
  wire f_s_dadda_pg_rca32_fa142_y3;
  wire f_s_dadda_pg_rca32_fa142_y4;
  wire f_s_dadda_pg_rca32_and_17_5_a_17;
  wire f_s_dadda_pg_rca32_and_17_5_b_5;
  wire f_s_dadda_pg_rca32_and_17_5_y0;
  wire f_s_dadda_pg_rca32_and_16_6_a_16;
  wire f_s_dadda_pg_rca32_and_16_6_b_6;
  wire f_s_dadda_pg_rca32_and_16_6_y0;
  wire f_s_dadda_pg_rca32_and_15_7_a_15;
  wire f_s_dadda_pg_rca32_and_15_7_b_7;
  wire f_s_dadda_pg_rca32_and_15_7_y0;
  wire f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_17_5_y0;
  wire f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_16_6_y0;
  wire f_s_dadda_pg_rca32_fa143_y0;
  wire f_s_dadda_pg_rca32_fa143_y1;
  wire f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_15_7_y0;
  wire f_s_dadda_pg_rca32_fa143_y2;
  wire f_s_dadda_pg_rca32_fa143_y3;
  wire f_s_dadda_pg_rca32_fa143_y4;
  wire f_s_dadda_pg_rca32_and_14_8_a_14;
  wire f_s_dadda_pg_rca32_and_14_8_b_8;
  wire f_s_dadda_pg_rca32_and_14_8_y0;
  wire f_s_dadda_pg_rca32_and_13_9_a_13;
  wire f_s_dadda_pg_rca32_and_13_9_b_9;
  wire f_s_dadda_pg_rca32_and_13_9_y0;
  wire f_s_dadda_pg_rca32_and_12_10_a_12;
  wire f_s_dadda_pg_rca32_and_12_10_b_10;
  wire f_s_dadda_pg_rca32_and_12_10_y0;
  wire f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_14_8_y0;
  wire f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_13_9_y0;
  wire f_s_dadda_pg_rca32_fa144_y0;
  wire f_s_dadda_pg_rca32_fa144_y1;
  wire f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_12_10_y0;
  wire f_s_dadda_pg_rca32_fa144_y2;
  wire f_s_dadda_pg_rca32_fa144_y3;
  wire f_s_dadda_pg_rca32_fa144_y4;
  wire f_s_dadda_pg_rca32_and_11_11_a_11;
  wire f_s_dadda_pg_rca32_and_11_11_b_11;
  wire f_s_dadda_pg_rca32_and_11_11_y0;
  wire f_s_dadda_pg_rca32_and_10_12_a_10;
  wire f_s_dadda_pg_rca32_and_10_12_b_12;
  wire f_s_dadda_pg_rca32_and_10_12_y0;
  wire f_s_dadda_pg_rca32_and_9_13_a_9;
  wire f_s_dadda_pg_rca32_and_9_13_b_13;
  wire f_s_dadda_pg_rca32_and_9_13_y0;
  wire f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_11_11_y0;
  wire f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_10_12_y0;
  wire f_s_dadda_pg_rca32_fa145_y0;
  wire f_s_dadda_pg_rca32_fa145_y1;
  wire f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_9_13_y0;
  wire f_s_dadda_pg_rca32_fa145_y2;
  wire f_s_dadda_pg_rca32_fa145_y3;
  wire f_s_dadda_pg_rca32_fa145_y4;
  wire f_s_dadda_pg_rca32_and_8_14_a_8;
  wire f_s_dadda_pg_rca32_and_8_14_b_14;
  wire f_s_dadda_pg_rca32_and_8_14_y0;
  wire f_s_dadda_pg_rca32_and_7_15_a_7;
  wire f_s_dadda_pg_rca32_and_7_15_b_15;
  wire f_s_dadda_pg_rca32_and_7_15_y0;
  wire f_s_dadda_pg_rca32_and_6_16_a_6;
  wire f_s_dadda_pg_rca32_and_6_16_b_16;
  wire f_s_dadda_pg_rca32_and_6_16_y0;
  wire f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_8_14_y0;
  wire f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_7_15_y0;
  wire f_s_dadda_pg_rca32_fa146_y0;
  wire f_s_dadda_pg_rca32_fa146_y1;
  wire f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_6_16_y0;
  wire f_s_dadda_pg_rca32_fa146_y2;
  wire f_s_dadda_pg_rca32_fa146_y3;
  wire f_s_dadda_pg_rca32_fa146_y4;
  wire f_s_dadda_pg_rca32_and_5_17_a_5;
  wire f_s_dadda_pg_rca32_and_5_17_b_17;
  wire f_s_dadda_pg_rca32_and_5_17_y0;
  wire f_s_dadda_pg_rca32_and_4_18_a_4;
  wire f_s_dadda_pg_rca32_and_4_18_b_18;
  wire f_s_dadda_pg_rca32_and_4_18_y0;
  wire f_s_dadda_pg_rca32_and_3_19_a_3;
  wire f_s_dadda_pg_rca32_and_3_19_b_19;
  wire f_s_dadda_pg_rca32_and_3_19_y0;
  wire f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_5_17_y0;
  wire f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_4_18_y0;
  wire f_s_dadda_pg_rca32_fa147_y0;
  wire f_s_dadda_pg_rca32_fa147_y1;
  wire f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_3_19_y0;
  wire f_s_dadda_pg_rca32_fa147_y2;
  wire f_s_dadda_pg_rca32_fa147_y3;
  wire f_s_dadda_pg_rca32_fa147_y4;
  wire f_s_dadda_pg_rca32_and_2_20_a_2;
  wire f_s_dadda_pg_rca32_and_2_20_b_20;
  wire f_s_dadda_pg_rca32_and_2_20_y0;
  wire f_s_dadda_pg_rca32_and_1_21_a_1;
  wire f_s_dadda_pg_rca32_and_1_21_b_21;
  wire f_s_dadda_pg_rca32_and_1_21_y0;
  wire f_s_dadda_pg_rca32_and_0_22_a_0;
  wire f_s_dadda_pg_rca32_and_0_22_b_22;
  wire f_s_dadda_pg_rca32_and_0_22_y0;
  wire f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_2_20_y0;
  wire f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_1_21_y0;
  wire f_s_dadda_pg_rca32_fa148_y0;
  wire f_s_dadda_pg_rca32_fa148_y1;
  wire f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_0_22_y0;
  wire f_s_dadda_pg_rca32_fa148_y2;
  wire f_s_dadda_pg_rca32_fa148_y3;
  wire f_s_dadda_pg_rca32_fa148_y4;
  wire f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa136_y2;
  wire f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa137_y2;
  wire f_s_dadda_pg_rca32_fa149_y0;
  wire f_s_dadda_pg_rca32_fa149_y1;
  wire f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa138_y2;
  wire f_s_dadda_pg_rca32_fa149_y2;
  wire f_s_dadda_pg_rca32_fa149_y3;
  wire f_s_dadda_pg_rca32_fa149_y4;
  wire f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa139_y2;
  wire f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa140_y2;
  wire f_s_dadda_pg_rca32_fa150_y0;
  wire f_s_dadda_pg_rca32_fa150_y1;
  wire f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa141_y2;
  wire f_s_dadda_pg_rca32_fa150_y2;
  wire f_s_dadda_pg_rca32_fa150_y3;
  wire f_s_dadda_pg_rca32_fa150_y4;
  wire f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa142_y2;
  wire f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa143_y2;
  wire f_s_dadda_pg_rca32_fa151_y0;
  wire f_s_dadda_pg_rca32_fa151_y1;
  wire f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa144_y2;
  wire f_s_dadda_pg_rca32_fa151_y2;
  wire f_s_dadda_pg_rca32_fa151_y3;
  wire f_s_dadda_pg_rca32_fa151_y4;
  wire f_s_dadda_pg_rca32_ha20_f_s_dadda_pg_rca32_fa145_y2;
  wire f_s_dadda_pg_rca32_ha20_f_s_dadda_pg_rca32_fa146_y2;
  wire f_s_dadda_pg_rca32_ha20_y0;
  wire f_s_dadda_pg_rca32_ha20_y1;
  wire f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_ha20_y1;
  wire f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_fa151_y4;
  wire f_s_dadda_pg_rca32_fa152_y0;
  wire f_s_dadda_pg_rca32_fa152_y1;
  wire f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_fa150_y4;
  wire f_s_dadda_pg_rca32_fa152_y2;
  wire f_s_dadda_pg_rca32_fa152_y3;
  wire f_s_dadda_pg_rca32_fa152_y4;
  wire f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa149_y4;
  wire f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa148_y4;
  wire f_s_dadda_pg_rca32_fa153_y0;
  wire f_s_dadda_pg_rca32_fa153_y1;
  wire f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa147_y4;
  wire f_s_dadda_pg_rca32_fa153_y2;
  wire f_s_dadda_pg_rca32_fa153_y3;
  wire f_s_dadda_pg_rca32_fa153_y4;
  wire f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa146_y4;
  wire f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa145_y4;
  wire f_s_dadda_pg_rca32_fa154_y0;
  wire f_s_dadda_pg_rca32_fa154_y1;
  wire f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa144_y4;
  wire f_s_dadda_pg_rca32_fa154_y2;
  wire f_s_dadda_pg_rca32_fa154_y3;
  wire f_s_dadda_pg_rca32_fa154_y4;
  wire f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa143_y4;
  wire f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa142_y4;
  wire f_s_dadda_pg_rca32_fa155_y0;
  wire f_s_dadda_pg_rca32_fa155_y1;
  wire f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa141_y4;
  wire f_s_dadda_pg_rca32_fa155_y2;
  wire f_s_dadda_pg_rca32_fa155_y3;
  wire f_s_dadda_pg_rca32_fa155_y4;
  wire f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa140_y4;
  wire f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa139_y4;
  wire f_s_dadda_pg_rca32_fa156_y0;
  wire f_s_dadda_pg_rca32_fa156_y1;
  wire f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa138_y4;
  wire f_s_dadda_pg_rca32_fa156_y2;
  wire f_s_dadda_pg_rca32_fa156_y3;
  wire f_s_dadda_pg_rca32_fa156_y4;
  wire f_s_dadda_pg_rca32_and_23_0_a_23;
  wire f_s_dadda_pg_rca32_and_23_0_b_0;
  wire f_s_dadda_pg_rca32_and_23_0_y0;
  wire f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_fa137_y4;
  wire f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_fa136_y4;
  wire f_s_dadda_pg_rca32_fa157_y0;
  wire f_s_dadda_pg_rca32_fa157_y1;
  wire f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_and_23_0_y0;
  wire f_s_dadda_pg_rca32_fa157_y2;
  wire f_s_dadda_pg_rca32_fa157_y3;
  wire f_s_dadda_pg_rca32_fa157_y4;
  wire f_s_dadda_pg_rca32_and_22_1_a_22;
  wire f_s_dadda_pg_rca32_and_22_1_b_1;
  wire f_s_dadda_pg_rca32_and_22_1_y0;
  wire f_s_dadda_pg_rca32_and_21_2_a_21;
  wire f_s_dadda_pg_rca32_and_21_2_b_2;
  wire f_s_dadda_pg_rca32_and_21_2_y0;
  wire f_s_dadda_pg_rca32_and_20_3_a_20;
  wire f_s_dadda_pg_rca32_and_20_3_b_3;
  wire f_s_dadda_pg_rca32_and_20_3_y0;
  wire f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_22_1_y0;
  wire f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_21_2_y0;
  wire f_s_dadda_pg_rca32_fa158_y0;
  wire f_s_dadda_pg_rca32_fa158_y1;
  wire f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_20_3_y0;
  wire f_s_dadda_pg_rca32_fa158_y2;
  wire f_s_dadda_pg_rca32_fa158_y3;
  wire f_s_dadda_pg_rca32_fa158_y4;
  wire f_s_dadda_pg_rca32_and_19_4_a_19;
  wire f_s_dadda_pg_rca32_and_19_4_b_4;
  wire f_s_dadda_pg_rca32_and_19_4_y0;
  wire f_s_dadda_pg_rca32_and_18_5_a_18;
  wire f_s_dadda_pg_rca32_and_18_5_b_5;
  wire f_s_dadda_pg_rca32_and_18_5_y0;
  wire f_s_dadda_pg_rca32_and_17_6_a_17;
  wire f_s_dadda_pg_rca32_and_17_6_b_6;
  wire f_s_dadda_pg_rca32_and_17_6_y0;
  wire f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_19_4_y0;
  wire f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_18_5_y0;
  wire f_s_dadda_pg_rca32_fa159_y0;
  wire f_s_dadda_pg_rca32_fa159_y1;
  wire f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_17_6_y0;
  wire f_s_dadda_pg_rca32_fa159_y2;
  wire f_s_dadda_pg_rca32_fa159_y3;
  wire f_s_dadda_pg_rca32_fa159_y4;
  wire f_s_dadda_pg_rca32_and_16_7_a_16;
  wire f_s_dadda_pg_rca32_and_16_7_b_7;
  wire f_s_dadda_pg_rca32_and_16_7_y0;
  wire f_s_dadda_pg_rca32_and_15_8_a_15;
  wire f_s_dadda_pg_rca32_and_15_8_b_8;
  wire f_s_dadda_pg_rca32_and_15_8_y0;
  wire f_s_dadda_pg_rca32_and_14_9_a_14;
  wire f_s_dadda_pg_rca32_and_14_9_b_9;
  wire f_s_dadda_pg_rca32_and_14_9_y0;
  wire f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_16_7_y0;
  wire f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_15_8_y0;
  wire f_s_dadda_pg_rca32_fa160_y0;
  wire f_s_dadda_pg_rca32_fa160_y1;
  wire f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_14_9_y0;
  wire f_s_dadda_pg_rca32_fa160_y2;
  wire f_s_dadda_pg_rca32_fa160_y3;
  wire f_s_dadda_pg_rca32_fa160_y4;
  wire f_s_dadda_pg_rca32_and_13_10_a_13;
  wire f_s_dadda_pg_rca32_and_13_10_b_10;
  wire f_s_dadda_pg_rca32_and_13_10_y0;
  wire f_s_dadda_pg_rca32_and_12_11_a_12;
  wire f_s_dadda_pg_rca32_and_12_11_b_11;
  wire f_s_dadda_pg_rca32_and_12_11_y0;
  wire f_s_dadda_pg_rca32_and_11_12_a_11;
  wire f_s_dadda_pg_rca32_and_11_12_b_12;
  wire f_s_dadda_pg_rca32_and_11_12_y0;
  wire f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_13_10_y0;
  wire f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_12_11_y0;
  wire f_s_dadda_pg_rca32_fa161_y0;
  wire f_s_dadda_pg_rca32_fa161_y1;
  wire f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_11_12_y0;
  wire f_s_dadda_pg_rca32_fa161_y2;
  wire f_s_dadda_pg_rca32_fa161_y3;
  wire f_s_dadda_pg_rca32_fa161_y4;
  wire f_s_dadda_pg_rca32_and_10_13_a_10;
  wire f_s_dadda_pg_rca32_and_10_13_b_13;
  wire f_s_dadda_pg_rca32_and_10_13_y0;
  wire f_s_dadda_pg_rca32_and_9_14_a_9;
  wire f_s_dadda_pg_rca32_and_9_14_b_14;
  wire f_s_dadda_pg_rca32_and_9_14_y0;
  wire f_s_dadda_pg_rca32_and_8_15_a_8;
  wire f_s_dadda_pg_rca32_and_8_15_b_15;
  wire f_s_dadda_pg_rca32_and_8_15_y0;
  wire f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_10_13_y0;
  wire f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_9_14_y0;
  wire f_s_dadda_pg_rca32_fa162_y0;
  wire f_s_dadda_pg_rca32_fa162_y1;
  wire f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_8_15_y0;
  wire f_s_dadda_pg_rca32_fa162_y2;
  wire f_s_dadda_pg_rca32_fa162_y3;
  wire f_s_dadda_pg_rca32_fa162_y4;
  wire f_s_dadda_pg_rca32_and_7_16_a_7;
  wire f_s_dadda_pg_rca32_and_7_16_b_16;
  wire f_s_dadda_pg_rca32_and_7_16_y0;
  wire f_s_dadda_pg_rca32_and_6_17_a_6;
  wire f_s_dadda_pg_rca32_and_6_17_b_17;
  wire f_s_dadda_pg_rca32_and_6_17_y0;
  wire f_s_dadda_pg_rca32_and_5_18_a_5;
  wire f_s_dadda_pg_rca32_and_5_18_b_18;
  wire f_s_dadda_pg_rca32_and_5_18_y0;
  wire f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_7_16_y0;
  wire f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_6_17_y0;
  wire f_s_dadda_pg_rca32_fa163_y0;
  wire f_s_dadda_pg_rca32_fa163_y1;
  wire f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_5_18_y0;
  wire f_s_dadda_pg_rca32_fa163_y2;
  wire f_s_dadda_pg_rca32_fa163_y3;
  wire f_s_dadda_pg_rca32_fa163_y4;
  wire f_s_dadda_pg_rca32_and_4_19_a_4;
  wire f_s_dadda_pg_rca32_and_4_19_b_19;
  wire f_s_dadda_pg_rca32_and_4_19_y0;
  wire f_s_dadda_pg_rca32_and_3_20_a_3;
  wire f_s_dadda_pg_rca32_and_3_20_b_20;
  wire f_s_dadda_pg_rca32_and_3_20_y0;
  wire f_s_dadda_pg_rca32_and_2_21_a_2;
  wire f_s_dadda_pg_rca32_and_2_21_b_21;
  wire f_s_dadda_pg_rca32_and_2_21_y0;
  wire f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_4_19_y0;
  wire f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_3_20_y0;
  wire f_s_dadda_pg_rca32_fa164_y0;
  wire f_s_dadda_pg_rca32_fa164_y1;
  wire f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_2_21_y0;
  wire f_s_dadda_pg_rca32_fa164_y2;
  wire f_s_dadda_pg_rca32_fa164_y3;
  wire f_s_dadda_pg_rca32_fa164_y4;
  wire f_s_dadda_pg_rca32_and_1_22_a_1;
  wire f_s_dadda_pg_rca32_and_1_22_b_22;
  wire f_s_dadda_pg_rca32_and_1_22_y0;
  wire f_s_dadda_pg_rca32_and_0_23_a_0;
  wire f_s_dadda_pg_rca32_and_0_23_b_23;
  wire f_s_dadda_pg_rca32_and_0_23_y0;
  wire f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_and_1_22_y0;
  wire f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_and_0_23_y0;
  wire f_s_dadda_pg_rca32_fa165_y0;
  wire f_s_dadda_pg_rca32_fa165_y1;
  wire f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_fa152_y2;
  wire f_s_dadda_pg_rca32_fa165_y2;
  wire f_s_dadda_pg_rca32_fa165_y3;
  wire f_s_dadda_pg_rca32_fa165_y4;
  wire f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa153_y2;
  wire f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa154_y2;
  wire f_s_dadda_pg_rca32_fa166_y0;
  wire f_s_dadda_pg_rca32_fa166_y1;
  wire f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa155_y2;
  wire f_s_dadda_pg_rca32_fa166_y2;
  wire f_s_dadda_pg_rca32_fa166_y3;
  wire f_s_dadda_pg_rca32_fa166_y4;
  wire f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa156_y2;
  wire f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa157_y2;
  wire f_s_dadda_pg_rca32_fa167_y0;
  wire f_s_dadda_pg_rca32_fa167_y1;
  wire f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa158_y2;
  wire f_s_dadda_pg_rca32_fa167_y2;
  wire f_s_dadda_pg_rca32_fa167_y3;
  wire f_s_dadda_pg_rca32_fa167_y4;
  wire f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa159_y2;
  wire f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa160_y2;
  wire f_s_dadda_pg_rca32_fa168_y0;
  wire f_s_dadda_pg_rca32_fa168_y1;
  wire f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa161_y2;
  wire f_s_dadda_pg_rca32_fa168_y2;
  wire f_s_dadda_pg_rca32_fa168_y3;
  wire f_s_dadda_pg_rca32_fa168_y4;
  wire f_s_dadda_pg_rca32_ha21_f_s_dadda_pg_rca32_fa162_y2;
  wire f_s_dadda_pg_rca32_ha21_f_s_dadda_pg_rca32_fa163_y2;
  wire f_s_dadda_pg_rca32_ha21_y0;
  wire f_s_dadda_pg_rca32_ha21_y1;
  wire f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_ha21_y1;
  wire f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_fa168_y4;
  wire f_s_dadda_pg_rca32_fa169_y0;
  wire f_s_dadda_pg_rca32_fa169_y1;
  wire f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_fa167_y4;
  wire f_s_dadda_pg_rca32_fa169_y2;
  wire f_s_dadda_pg_rca32_fa169_y3;
  wire f_s_dadda_pg_rca32_fa169_y4;
  wire f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa166_y4;
  wire f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa165_y4;
  wire f_s_dadda_pg_rca32_fa170_y0;
  wire f_s_dadda_pg_rca32_fa170_y1;
  wire f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa164_y4;
  wire f_s_dadda_pg_rca32_fa170_y2;
  wire f_s_dadda_pg_rca32_fa170_y3;
  wire f_s_dadda_pg_rca32_fa170_y4;
  wire f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa163_y4;
  wire f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa162_y4;
  wire f_s_dadda_pg_rca32_fa171_y0;
  wire f_s_dadda_pg_rca32_fa171_y1;
  wire f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa161_y4;
  wire f_s_dadda_pg_rca32_fa171_y2;
  wire f_s_dadda_pg_rca32_fa171_y3;
  wire f_s_dadda_pg_rca32_fa171_y4;
  wire f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa160_y4;
  wire f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa159_y4;
  wire f_s_dadda_pg_rca32_fa172_y0;
  wire f_s_dadda_pg_rca32_fa172_y1;
  wire f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa158_y4;
  wire f_s_dadda_pg_rca32_fa172_y2;
  wire f_s_dadda_pg_rca32_fa172_y3;
  wire f_s_dadda_pg_rca32_fa172_y4;
  wire f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa157_y4;
  wire f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa156_y4;
  wire f_s_dadda_pg_rca32_fa173_y0;
  wire f_s_dadda_pg_rca32_fa173_y1;
  wire f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa155_y4;
  wire f_s_dadda_pg_rca32_fa173_y2;
  wire f_s_dadda_pg_rca32_fa173_y3;
  wire f_s_dadda_pg_rca32_fa173_y4;
  wire f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa154_y4;
  wire f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa153_y4;
  wire f_s_dadda_pg_rca32_fa174_y0;
  wire f_s_dadda_pg_rca32_fa174_y1;
  wire f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa152_y4;
  wire f_s_dadda_pg_rca32_fa174_y2;
  wire f_s_dadda_pg_rca32_fa174_y3;
  wire f_s_dadda_pg_rca32_fa174_y4;
  wire f_s_dadda_pg_rca32_and_24_0_a_24;
  wire f_s_dadda_pg_rca32_and_24_0_b_0;
  wire f_s_dadda_pg_rca32_and_24_0_y0;
  wire f_s_dadda_pg_rca32_and_23_1_a_23;
  wire f_s_dadda_pg_rca32_and_23_1_b_1;
  wire f_s_dadda_pg_rca32_and_23_1_y0;
  wire f_s_dadda_pg_rca32_and_22_2_a_22;
  wire f_s_dadda_pg_rca32_and_22_2_b_2;
  wire f_s_dadda_pg_rca32_and_22_2_y0;
  wire f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_24_0_y0;
  wire f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_23_1_y0;
  wire f_s_dadda_pg_rca32_fa175_y0;
  wire f_s_dadda_pg_rca32_fa175_y1;
  wire f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_22_2_y0;
  wire f_s_dadda_pg_rca32_fa175_y2;
  wire f_s_dadda_pg_rca32_fa175_y3;
  wire f_s_dadda_pg_rca32_fa175_y4;
  wire f_s_dadda_pg_rca32_and_21_3_a_21;
  wire f_s_dadda_pg_rca32_and_21_3_b_3;
  wire f_s_dadda_pg_rca32_and_21_3_y0;
  wire f_s_dadda_pg_rca32_and_20_4_a_20;
  wire f_s_dadda_pg_rca32_and_20_4_b_4;
  wire f_s_dadda_pg_rca32_and_20_4_y0;
  wire f_s_dadda_pg_rca32_and_19_5_a_19;
  wire f_s_dadda_pg_rca32_and_19_5_b_5;
  wire f_s_dadda_pg_rca32_and_19_5_y0;
  wire f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_21_3_y0;
  wire f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_20_4_y0;
  wire f_s_dadda_pg_rca32_fa176_y0;
  wire f_s_dadda_pg_rca32_fa176_y1;
  wire f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_19_5_y0;
  wire f_s_dadda_pg_rca32_fa176_y2;
  wire f_s_dadda_pg_rca32_fa176_y3;
  wire f_s_dadda_pg_rca32_fa176_y4;
  wire f_s_dadda_pg_rca32_and_18_6_a_18;
  wire f_s_dadda_pg_rca32_and_18_6_b_6;
  wire f_s_dadda_pg_rca32_and_18_6_y0;
  wire f_s_dadda_pg_rca32_and_17_7_a_17;
  wire f_s_dadda_pg_rca32_and_17_7_b_7;
  wire f_s_dadda_pg_rca32_and_17_7_y0;
  wire f_s_dadda_pg_rca32_and_16_8_a_16;
  wire f_s_dadda_pg_rca32_and_16_8_b_8;
  wire f_s_dadda_pg_rca32_and_16_8_y0;
  wire f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_18_6_y0;
  wire f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_17_7_y0;
  wire f_s_dadda_pg_rca32_fa177_y0;
  wire f_s_dadda_pg_rca32_fa177_y1;
  wire f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_16_8_y0;
  wire f_s_dadda_pg_rca32_fa177_y2;
  wire f_s_dadda_pg_rca32_fa177_y3;
  wire f_s_dadda_pg_rca32_fa177_y4;
  wire f_s_dadda_pg_rca32_and_15_9_a_15;
  wire f_s_dadda_pg_rca32_and_15_9_b_9;
  wire f_s_dadda_pg_rca32_and_15_9_y0;
  wire f_s_dadda_pg_rca32_and_14_10_a_14;
  wire f_s_dadda_pg_rca32_and_14_10_b_10;
  wire f_s_dadda_pg_rca32_and_14_10_y0;
  wire f_s_dadda_pg_rca32_and_13_11_a_13;
  wire f_s_dadda_pg_rca32_and_13_11_b_11;
  wire f_s_dadda_pg_rca32_and_13_11_y0;
  wire f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_15_9_y0;
  wire f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_14_10_y0;
  wire f_s_dadda_pg_rca32_fa178_y0;
  wire f_s_dadda_pg_rca32_fa178_y1;
  wire f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_13_11_y0;
  wire f_s_dadda_pg_rca32_fa178_y2;
  wire f_s_dadda_pg_rca32_fa178_y3;
  wire f_s_dadda_pg_rca32_fa178_y4;
  wire f_s_dadda_pg_rca32_and_12_12_a_12;
  wire f_s_dadda_pg_rca32_and_12_12_b_12;
  wire f_s_dadda_pg_rca32_and_12_12_y0;
  wire f_s_dadda_pg_rca32_and_11_13_a_11;
  wire f_s_dadda_pg_rca32_and_11_13_b_13;
  wire f_s_dadda_pg_rca32_and_11_13_y0;
  wire f_s_dadda_pg_rca32_and_10_14_a_10;
  wire f_s_dadda_pg_rca32_and_10_14_b_14;
  wire f_s_dadda_pg_rca32_and_10_14_y0;
  wire f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_12_12_y0;
  wire f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_11_13_y0;
  wire f_s_dadda_pg_rca32_fa179_y0;
  wire f_s_dadda_pg_rca32_fa179_y1;
  wire f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_10_14_y0;
  wire f_s_dadda_pg_rca32_fa179_y2;
  wire f_s_dadda_pg_rca32_fa179_y3;
  wire f_s_dadda_pg_rca32_fa179_y4;
  wire f_s_dadda_pg_rca32_and_9_15_a_9;
  wire f_s_dadda_pg_rca32_and_9_15_b_15;
  wire f_s_dadda_pg_rca32_and_9_15_y0;
  wire f_s_dadda_pg_rca32_and_8_16_a_8;
  wire f_s_dadda_pg_rca32_and_8_16_b_16;
  wire f_s_dadda_pg_rca32_and_8_16_y0;
  wire f_s_dadda_pg_rca32_and_7_17_a_7;
  wire f_s_dadda_pg_rca32_and_7_17_b_17;
  wire f_s_dadda_pg_rca32_and_7_17_y0;
  wire f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_9_15_y0;
  wire f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_8_16_y0;
  wire f_s_dadda_pg_rca32_fa180_y0;
  wire f_s_dadda_pg_rca32_fa180_y1;
  wire f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_7_17_y0;
  wire f_s_dadda_pg_rca32_fa180_y2;
  wire f_s_dadda_pg_rca32_fa180_y3;
  wire f_s_dadda_pg_rca32_fa180_y4;
  wire f_s_dadda_pg_rca32_and_6_18_a_6;
  wire f_s_dadda_pg_rca32_and_6_18_b_18;
  wire f_s_dadda_pg_rca32_and_6_18_y0;
  wire f_s_dadda_pg_rca32_and_5_19_a_5;
  wire f_s_dadda_pg_rca32_and_5_19_b_19;
  wire f_s_dadda_pg_rca32_and_5_19_y0;
  wire f_s_dadda_pg_rca32_and_4_20_a_4;
  wire f_s_dadda_pg_rca32_and_4_20_b_20;
  wire f_s_dadda_pg_rca32_and_4_20_y0;
  wire f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_6_18_y0;
  wire f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_5_19_y0;
  wire f_s_dadda_pg_rca32_fa181_y0;
  wire f_s_dadda_pg_rca32_fa181_y1;
  wire f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_4_20_y0;
  wire f_s_dadda_pg_rca32_fa181_y2;
  wire f_s_dadda_pg_rca32_fa181_y3;
  wire f_s_dadda_pg_rca32_fa181_y4;
  wire f_s_dadda_pg_rca32_and_3_21_a_3;
  wire f_s_dadda_pg_rca32_and_3_21_b_21;
  wire f_s_dadda_pg_rca32_and_3_21_y0;
  wire f_s_dadda_pg_rca32_and_2_22_a_2;
  wire f_s_dadda_pg_rca32_and_2_22_b_22;
  wire f_s_dadda_pg_rca32_and_2_22_y0;
  wire f_s_dadda_pg_rca32_and_1_23_a_1;
  wire f_s_dadda_pg_rca32_and_1_23_b_23;
  wire f_s_dadda_pg_rca32_and_1_23_y0;
  wire f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_3_21_y0;
  wire f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_2_22_y0;
  wire f_s_dadda_pg_rca32_fa182_y0;
  wire f_s_dadda_pg_rca32_fa182_y1;
  wire f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_1_23_y0;
  wire f_s_dadda_pg_rca32_fa182_y2;
  wire f_s_dadda_pg_rca32_fa182_y3;
  wire f_s_dadda_pg_rca32_fa182_y4;
  wire f_s_dadda_pg_rca32_and_0_24_a_0;
  wire f_s_dadda_pg_rca32_and_0_24_b_24;
  wire f_s_dadda_pg_rca32_and_0_24_y0;
  wire f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_and_0_24_y0;
  wire f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_fa169_y2;
  wire f_s_dadda_pg_rca32_fa183_y0;
  wire f_s_dadda_pg_rca32_fa183_y1;
  wire f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_fa170_y2;
  wire f_s_dadda_pg_rca32_fa183_y2;
  wire f_s_dadda_pg_rca32_fa183_y3;
  wire f_s_dadda_pg_rca32_fa183_y4;
  wire f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa171_y2;
  wire f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa172_y2;
  wire f_s_dadda_pg_rca32_fa184_y0;
  wire f_s_dadda_pg_rca32_fa184_y1;
  wire f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa173_y2;
  wire f_s_dadda_pg_rca32_fa184_y2;
  wire f_s_dadda_pg_rca32_fa184_y3;
  wire f_s_dadda_pg_rca32_fa184_y4;
  wire f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa174_y2;
  wire f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa175_y2;
  wire f_s_dadda_pg_rca32_fa185_y0;
  wire f_s_dadda_pg_rca32_fa185_y1;
  wire f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa176_y2;
  wire f_s_dadda_pg_rca32_fa185_y2;
  wire f_s_dadda_pg_rca32_fa185_y3;
  wire f_s_dadda_pg_rca32_fa185_y4;
  wire f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa177_y2;
  wire f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa178_y2;
  wire f_s_dadda_pg_rca32_fa186_y0;
  wire f_s_dadda_pg_rca32_fa186_y1;
  wire f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa179_y2;
  wire f_s_dadda_pg_rca32_fa186_y2;
  wire f_s_dadda_pg_rca32_fa186_y3;
  wire f_s_dadda_pg_rca32_fa186_y4;
  wire f_s_dadda_pg_rca32_ha22_f_s_dadda_pg_rca32_fa180_y2;
  wire f_s_dadda_pg_rca32_ha22_f_s_dadda_pg_rca32_fa181_y2;
  wire f_s_dadda_pg_rca32_ha22_y0;
  wire f_s_dadda_pg_rca32_ha22_y1;
  wire f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_ha22_y1;
  wire f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_fa186_y4;
  wire f_s_dadda_pg_rca32_fa187_y0;
  wire f_s_dadda_pg_rca32_fa187_y1;
  wire f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_fa185_y4;
  wire f_s_dadda_pg_rca32_fa187_y2;
  wire f_s_dadda_pg_rca32_fa187_y3;
  wire f_s_dadda_pg_rca32_fa187_y4;
  wire f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa184_y4;
  wire f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa183_y4;
  wire f_s_dadda_pg_rca32_fa188_y0;
  wire f_s_dadda_pg_rca32_fa188_y1;
  wire f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa182_y4;
  wire f_s_dadda_pg_rca32_fa188_y2;
  wire f_s_dadda_pg_rca32_fa188_y3;
  wire f_s_dadda_pg_rca32_fa188_y4;
  wire f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa181_y4;
  wire f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa180_y4;
  wire f_s_dadda_pg_rca32_fa189_y0;
  wire f_s_dadda_pg_rca32_fa189_y1;
  wire f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa179_y4;
  wire f_s_dadda_pg_rca32_fa189_y2;
  wire f_s_dadda_pg_rca32_fa189_y3;
  wire f_s_dadda_pg_rca32_fa189_y4;
  wire f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa178_y4;
  wire f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa177_y4;
  wire f_s_dadda_pg_rca32_fa190_y0;
  wire f_s_dadda_pg_rca32_fa190_y1;
  wire f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa176_y4;
  wire f_s_dadda_pg_rca32_fa190_y2;
  wire f_s_dadda_pg_rca32_fa190_y3;
  wire f_s_dadda_pg_rca32_fa190_y4;
  wire f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa175_y4;
  wire f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa174_y4;
  wire f_s_dadda_pg_rca32_fa191_y0;
  wire f_s_dadda_pg_rca32_fa191_y1;
  wire f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa173_y4;
  wire f_s_dadda_pg_rca32_fa191_y2;
  wire f_s_dadda_pg_rca32_fa191_y3;
  wire f_s_dadda_pg_rca32_fa191_y4;
  wire f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa172_y4;
  wire f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa171_y4;
  wire f_s_dadda_pg_rca32_fa192_y0;
  wire f_s_dadda_pg_rca32_fa192_y1;
  wire f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa170_y4;
  wire f_s_dadda_pg_rca32_fa192_y2;
  wire f_s_dadda_pg_rca32_fa192_y3;
  wire f_s_dadda_pg_rca32_fa192_y4;
  wire f_s_dadda_pg_rca32_and_25_0_a_25;
  wire f_s_dadda_pg_rca32_and_25_0_b_0;
  wire f_s_dadda_pg_rca32_and_25_0_y0;
  wire f_s_dadda_pg_rca32_and_24_1_a_24;
  wire f_s_dadda_pg_rca32_and_24_1_b_1;
  wire f_s_dadda_pg_rca32_and_24_1_y0;
  wire f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_fa169_y4;
  wire f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_and_25_0_y0;
  wire f_s_dadda_pg_rca32_fa193_y0;
  wire f_s_dadda_pg_rca32_fa193_y1;
  wire f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_and_24_1_y0;
  wire f_s_dadda_pg_rca32_fa193_y2;
  wire f_s_dadda_pg_rca32_fa193_y3;
  wire f_s_dadda_pg_rca32_fa193_y4;
  wire f_s_dadda_pg_rca32_and_23_2_a_23;
  wire f_s_dadda_pg_rca32_and_23_2_b_2;
  wire f_s_dadda_pg_rca32_and_23_2_y0;
  wire f_s_dadda_pg_rca32_and_22_3_a_22;
  wire f_s_dadda_pg_rca32_and_22_3_b_3;
  wire f_s_dadda_pg_rca32_and_22_3_y0;
  wire f_s_dadda_pg_rca32_and_21_4_a_21;
  wire f_s_dadda_pg_rca32_and_21_4_b_4;
  wire f_s_dadda_pg_rca32_and_21_4_y0;
  wire f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_23_2_y0;
  wire f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_22_3_y0;
  wire f_s_dadda_pg_rca32_fa194_y0;
  wire f_s_dadda_pg_rca32_fa194_y1;
  wire f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_21_4_y0;
  wire f_s_dadda_pg_rca32_fa194_y2;
  wire f_s_dadda_pg_rca32_fa194_y3;
  wire f_s_dadda_pg_rca32_fa194_y4;
  wire f_s_dadda_pg_rca32_and_20_5_a_20;
  wire f_s_dadda_pg_rca32_and_20_5_b_5;
  wire f_s_dadda_pg_rca32_and_20_5_y0;
  wire f_s_dadda_pg_rca32_and_19_6_a_19;
  wire f_s_dadda_pg_rca32_and_19_6_b_6;
  wire f_s_dadda_pg_rca32_and_19_6_y0;
  wire f_s_dadda_pg_rca32_and_18_7_a_18;
  wire f_s_dadda_pg_rca32_and_18_7_b_7;
  wire f_s_dadda_pg_rca32_and_18_7_y0;
  wire f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_20_5_y0;
  wire f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_19_6_y0;
  wire f_s_dadda_pg_rca32_fa195_y0;
  wire f_s_dadda_pg_rca32_fa195_y1;
  wire f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_18_7_y0;
  wire f_s_dadda_pg_rca32_fa195_y2;
  wire f_s_dadda_pg_rca32_fa195_y3;
  wire f_s_dadda_pg_rca32_fa195_y4;
  wire f_s_dadda_pg_rca32_and_17_8_a_17;
  wire f_s_dadda_pg_rca32_and_17_8_b_8;
  wire f_s_dadda_pg_rca32_and_17_8_y0;
  wire f_s_dadda_pg_rca32_and_16_9_a_16;
  wire f_s_dadda_pg_rca32_and_16_9_b_9;
  wire f_s_dadda_pg_rca32_and_16_9_y0;
  wire f_s_dadda_pg_rca32_and_15_10_a_15;
  wire f_s_dadda_pg_rca32_and_15_10_b_10;
  wire f_s_dadda_pg_rca32_and_15_10_y0;
  wire f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_17_8_y0;
  wire f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_16_9_y0;
  wire f_s_dadda_pg_rca32_fa196_y0;
  wire f_s_dadda_pg_rca32_fa196_y1;
  wire f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_15_10_y0;
  wire f_s_dadda_pg_rca32_fa196_y2;
  wire f_s_dadda_pg_rca32_fa196_y3;
  wire f_s_dadda_pg_rca32_fa196_y4;
  wire f_s_dadda_pg_rca32_and_14_11_a_14;
  wire f_s_dadda_pg_rca32_and_14_11_b_11;
  wire f_s_dadda_pg_rca32_and_14_11_y0;
  wire f_s_dadda_pg_rca32_and_13_12_a_13;
  wire f_s_dadda_pg_rca32_and_13_12_b_12;
  wire f_s_dadda_pg_rca32_and_13_12_y0;
  wire f_s_dadda_pg_rca32_and_12_13_a_12;
  wire f_s_dadda_pg_rca32_and_12_13_b_13;
  wire f_s_dadda_pg_rca32_and_12_13_y0;
  wire f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_14_11_y0;
  wire f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_13_12_y0;
  wire f_s_dadda_pg_rca32_fa197_y0;
  wire f_s_dadda_pg_rca32_fa197_y1;
  wire f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_12_13_y0;
  wire f_s_dadda_pg_rca32_fa197_y2;
  wire f_s_dadda_pg_rca32_fa197_y3;
  wire f_s_dadda_pg_rca32_fa197_y4;
  wire f_s_dadda_pg_rca32_and_11_14_a_11;
  wire f_s_dadda_pg_rca32_and_11_14_b_14;
  wire f_s_dadda_pg_rca32_and_11_14_y0;
  wire f_s_dadda_pg_rca32_and_10_15_a_10;
  wire f_s_dadda_pg_rca32_and_10_15_b_15;
  wire f_s_dadda_pg_rca32_and_10_15_y0;
  wire f_s_dadda_pg_rca32_and_9_16_a_9;
  wire f_s_dadda_pg_rca32_and_9_16_b_16;
  wire f_s_dadda_pg_rca32_and_9_16_y0;
  wire f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_11_14_y0;
  wire f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_10_15_y0;
  wire f_s_dadda_pg_rca32_fa198_y0;
  wire f_s_dadda_pg_rca32_fa198_y1;
  wire f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_9_16_y0;
  wire f_s_dadda_pg_rca32_fa198_y2;
  wire f_s_dadda_pg_rca32_fa198_y3;
  wire f_s_dadda_pg_rca32_fa198_y4;
  wire f_s_dadda_pg_rca32_and_8_17_a_8;
  wire f_s_dadda_pg_rca32_and_8_17_b_17;
  wire f_s_dadda_pg_rca32_and_8_17_y0;
  wire f_s_dadda_pg_rca32_and_7_18_a_7;
  wire f_s_dadda_pg_rca32_and_7_18_b_18;
  wire f_s_dadda_pg_rca32_and_7_18_y0;
  wire f_s_dadda_pg_rca32_and_6_19_a_6;
  wire f_s_dadda_pg_rca32_and_6_19_b_19;
  wire f_s_dadda_pg_rca32_and_6_19_y0;
  wire f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_8_17_y0;
  wire f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_7_18_y0;
  wire f_s_dadda_pg_rca32_fa199_y0;
  wire f_s_dadda_pg_rca32_fa199_y1;
  wire f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_6_19_y0;
  wire f_s_dadda_pg_rca32_fa199_y2;
  wire f_s_dadda_pg_rca32_fa199_y3;
  wire f_s_dadda_pg_rca32_fa199_y4;
  wire f_s_dadda_pg_rca32_and_5_20_a_5;
  wire f_s_dadda_pg_rca32_and_5_20_b_20;
  wire f_s_dadda_pg_rca32_and_5_20_y0;
  wire f_s_dadda_pg_rca32_and_4_21_a_4;
  wire f_s_dadda_pg_rca32_and_4_21_b_21;
  wire f_s_dadda_pg_rca32_and_4_21_y0;
  wire f_s_dadda_pg_rca32_and_3_22_a_3;
  wire f_s_dadda_pg_rca32_and_3_22_b_22;
  wire f_s_dadda_pg_rca32_and_3_22_y0;
  wire f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_5_20_y0;
  wire f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_4_21_y0;
  wire f_s_dadda_pg_rca32_fa200_y0;
  wire f_s_dadda_pg_rca32_fa200_y1;
  wire f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_3_22_y0;
  wire f_s_dadda_pg_rca32_fa200_y2;
  wire f_s_dadda_pg_rca32_fa200_y3;
  wire f_s_dadda_pg_rca32_fa200_y4;
  wire f_s_dadda_pg_rca32_and_2_23_a_2;
  wire f_s_dadda_pg_rca32_and_2_23_b_23;
  wire f_s_dadda_pg_rca32_and_2_23_y0;
  wire f_s_dadda_pg_rca32_and_1_24_a_1;
  wire f_s_dadda_pg_rca32_and_1_24_b_24;
  wire f_s_dadda_pg_rca32_and_1_24_y0;
  wire f_s_dadda_pg_rca32_and_0_25_a_0;
  wire f_s_dadda_pg_rca32_and_0_25_b_25;
  wire f_s_dadda_pg_rca32_and_0_25_y0;
  wire f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_2_23_y0;
  wire f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_1_24_y0;
  wire f_s_dadda_pg_rca32_fa201_y0;
  wire f_s_dadda_pg_rca32_fa201_y1;
  wire f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_0_25_y0;
  wire f_s_dadda_pg_rca32_fa201_y2;
  wire f_s_dadda_pg_rca32_fa201_y3;
  wire f_s_dadda_pg_rca32_fa201_y4;
  wire f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa187_y2;
  wire f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa188_y2;
  wire f_s_dadda_pg_rca32_fa202_y0;
  wire f_s_dadda_pg_rca32_fa202_y1;
  wire f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa189_y2;
  wire f_s_dadda_pg_rca32_fa202_y2;
  wire f_s_dadda_pg_rca32_fa202_y3;
  wire f_s_dadda_pg_rca32_fa202_y4;
  wire f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa190_y2;
  wire f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa191_y2;
  wire f_s_dadda_pg_rca32_fa203_y0;
  wire f_s_dadda_pg_rca32_fa203_y1;
  wire f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa192_y2;
  wire f_s_dadda_pg_rca32_fa203_y2;
  wire f_s_dadda_pg_rca32_fa203_y3;
  wire f_s_dadda_pg_rca32_fa203_y4;
  wire f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa193_y2;
  wire f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa194_y2;
  wire f_s_dadda_pg_rca32_fa204_y0;
  wire f_s_dadda_pg_rca32_fa204_y1;
  wire f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa195_y2;
  wire f_s_dadda_pg_rca32_fa204_y2;
  wire f_s_dadda_pg_rca32_fa204_y3;
  wire f_s_dadda_pg_rca32_fa204_y4;
  wire f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa196_y2;
  wire f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa197_y2;
  wire f_s_dadda_pg_rca32_fa205_y0;
  wire f_s_dadda_pg_rca32_fa205_y1;
  wire f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa198_y2;
  wire f_s_dadda_pg_rca32_fa205_y2;
  wire f_s_dadda_pg_rca32_fa205_y3;
  wire f_s_dadda_pg_rca32_fa205_y4;
  wire f_s_dadda_pg_rca32_ha23_f_s_dadda_pg_rca32_fa199_y2;
  wire f_s_dadda_pg_rca32_ha23_f_s_dadda_pg_rca32_fa200_y2;
  wire f_s_dadda_pg_rca32_ha23_y0;
  wire f_s_dadda_pg_rca32_ha23_y1;
  wire f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_ha23_y1;
  wire f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_fa205_y4;
  wire f_s_dadda_pg_rca32_fa206_y0;
  wire f_s_dadda_pg_rca32_fa206_y1;
  wire f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_fa204_y4;
  wire f_s_dadda_pg_rca32_fa206_y2;
  wire f_s_dadda_pg_rca32_fa206_y3;
  wire f_s_dadda_pg_rca32_fa206_y4;
  wire f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa203_y4;
  wire f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa202_y4;
  wire f_s_dadda_pg_rca32_fa207_y0;
  wire f_s_dadda_pg_rca32_fa207_y1;
  wire f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa201_y4;
  wire f_s_dadda_pg_rca32_fa207_y2;
  wire f_s_dadda_pg_rca32_fa207_y3;
  wire f_s_dadda_pg_rca32_fa207_y4;
  wire f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa200_y4;
  wire f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa199_y4;
  wire f_s_dadda_pg_rca32_fa208_y0;
  wire f_s_dadda_pg_rca32_fa208_y1;
  wire f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa198_y4;
  wire f_s_dadda_pg_rca32_fa208_y2;
  wire f_s_dadda_pg_rca32_fa208_y3;
  wire f_s_dadda_pg_rca32_fa208_y4;
  wire f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa197_y4;
  wire f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa196_y4;
  wire f_s_dadda_pg_rca32_fa209_y0;
  wire f_s_dadda_pg_rca32_fa209_y1;
  wire f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa195_y4;
  wire f_s_dadda_pg_rca32_fa209_y2;
  wire f_s_dadda_pg_rca32_fa209_y3;
  wire f_s_dadda_pg_rca32_fa209_y4;
  wire f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa194_y4;
  wire f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa193_y4;
  wire f_s_dadda_pg_rca32_fa210_y0;
  wire f_s_dadda_pg_rca32_fa210_y1;
  wire f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa192_y4;
  wire f_s_dadda_pg_rca32_fa210_y2;
  wire f_s_dadda_pg_rca32_fa210_y3;
  wire f_s_dadda_pg_rca32_fa210_y4;
  wire f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa191_y4;
  wire f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa190_y4;
  wire f_s_dadda_pg_rca32_fa211_y0;
  wire f_s_dadda_pg_rca32_fa211_y1;
  wire f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa189_y4;
  wire f_s_dadda_pg_rca32_fa211_y2;
  wire f_s_dadda_pg_rca32_fa211_y3;
  wire f_s_dadda_pg_rca32_fa211_y4;
  wire f_s_dadda_pg_rca32_and_26_0_a_26;
  wire f_s_dadda_pg_rca32_and_26_0_b_0;
  wire f_s_dadda_pg_rca32_and_26_0_y0;
  wire f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_fa188_y4;
  wire f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_fa187_y4;
  wire f_s_dadda_pg_rca32_fa212_y0;
  wire f_s_dadda_pg_rca32_fa212_y1;
  wire f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_and_26_0_y0;
  wire f_s_dadda_pg_rca32_fa212_y2;
  wire f_s_dadda_pg_rca32_fa212_y3;
  wire f_s_dadda_pg_rca32_fa212_y4;
  wire f_s_dadda_pg_rca32_and_25_1_a_25;
  wire f_s_dadda_pg_rca32_and_25_1_b_1;
  wire f_s_dadda_pg_rca32_and_25_1_y0;
  wire f_s_dadda_pg_rca32_and_24_2_a_24;
  wire f_s_dadda_pg_rca32_and_24_2_b_2;
  wire f_s_dadda_pg_rca32_and_24_2_y0;
  wire f_s_dadda_pg_rca32_and_23_3_a_23;
  wire f_s_dadda_pg_rca32_and_23_3_b_3;
  wire f_s_dadda_pg_rca32_and_23_3_y0;
  wire f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_25_1_y0;
  wire f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_24_2_y0;
  wire f_s_dadda_pg_rca32_fa213_y0;
  wire f_s_dadda_pg_rca32_fa213_y1;
  wire f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_23_3_y0;
  wire f_s_dadda_pg_rca32_fa213_y2;
  wire f_s_dadda_pg_rca32_fa213_y3;
  wire f_s_dadda_pg_rca32_fa213_y4;
  wire f_s_dadda_pg_rca32_and_22_4_a_22;
  wire f_s_dadda_pg_rca32_and_22_4_b_4;
  wire f_s_dadda_pg_rca32_and_22_4_y0;
  wire f_s_dadda_pg_rca32_and_21_5_a_21;
  wire f_s_dadda_pg_rca32_and_21_5_b_5;
  wire f_s_dadda_pg_rca32_and_21_5_y0;
  wire f_s_dadda_pg_rca32_and_20_6_a_20;
  wire f_s_dadda_pg_rca32_and_20_6_b_6;
  wire f_s_dadda_pg_rca32_and_20_6_y0;
  wire f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_22_4_y0;
  wire f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_21_5_y0;
  wire f_s_dadda_pg_rca32_fa214_y0;
  wire f_s_dadda_pg_rca32_fa214_y1;
  wire f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_20_6_y0;
  wire f_s_dadda_pg_rca32_fa214_y2;
  wire f_s_dadda_pg_rca32_fa214_y3;
  wire f_s_dadda_pg_rca32_fa214_y4;
  wire f_s_dadda_pg_rca32_and_19_7_a_19;
  wire f_s_dadda_pg_rca32_and_19_7_b_7;
  wire f_s_dadda_pg_rca32_and_19_7_y0;
  wire f_s_dadda_pg_rca32_and_18_8_a_18;
  wire f_s_dadda_pg_rca32_and_18_8_b_8;
  wire f_s_dadda_pg_rca32_and_18_8_y0;
  wire f_s_dadda_pg_rca32_and_17_9_a_17;
  wire f_s_dadda_pg_rca32_and_17_9_b_9;
  wire f_s_dadda_pg_rca32_and_17_9_y0;
  wire f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_19_7_y0;
  wire f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_18_8_y0;
  wire f_s_dadda_pg_rca32_fa215_y0;
  wire f_s_dadda_pg_rca32_fa215_y1;
  wire f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_17_9_y0;
  wire f_s_dadda_pg_rca32_fa215_y2;
  wire f_s_dadda_pg_rca32_fa215_y3;
  wire f_s_dadda_pg_rca32_fa215_y4;
  wire f_s_dadda_pg_rca32_and_16_10_a_16;
  wire f_s_dadda_pg_rca32_and_16_10_b_10;
  wire f_s_dadda_pg_rca32_and_16_10_y0;
  wire f_s_dadda_pg_rca32_and_15_11_a_15;
  wire f_s_dadda_pg_rca32_and_15_11_b_11;
  wire f_s_dadda_pg_rca32_and_15_11_y0;
  wire f_s_dadda_pg_rca32_and_14_12_a_14;
  wire f_s_dadda_pg_rca32_and_14_12_b_12;
  wire f_s_dadda_pg_rca32_and_14_12_y0;
  wire f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_16_10_y0;
  wire f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_15_11_y0;
  wire f_s_dadda_pg_rca32_fa216_y0;
  wire f_s_dadda_pg_rca32_fa216_y1;
  wire f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_14_12_y0;
  wire f_s_dadda_pg_rca32_fa216_y2;
  wire f_s_dadda_pg_rca32_fa216_y3;
  wire f_s_dadda_pg_rca32_fa216_y4;
  wire f_s_dadda_pg_rca32_and_13_13_a_13;
  wire f_s_dadda_pg_rca32_and_13_13_b_13;
  wire f_s_dadda_pg_rca32_and_13_13_y0;
  wire f_s_dadda_pg_rca32_and_12_14_a_12;
  wire f_s_dadda_pg_rca32_and_12_14_b_14;
  wire f_s_dadda_pg_rca32_and_12_14_y0;
  wire f_s_dadda_pg_rca32_and_11_15_a_11;
  wire f_s_dadda_pg_rca32_and_11_15_b_15;
  wire f_s_dadda_pg_rca32_and_11_15_y0;
  wire f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_13_13_y0;
  wire f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_12_14_y0;
  wire f_s_dadda_pg_rca32_fa217_y0;
  wire f_s_dadda_pg_rca32_fa217_y1;
  wire f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_11_15_y0;
  wire f_s_dadda_pg_rca32_fa217_y2;
  wire f_s_dadda_pg_rca32_fa217_y3;
  wire f_s_dadda_pg_rca32_fa217_y4;
  wire f_s_dadda_pg_rca32_and_10_16_a_10;
  wire f_s_dadda_pg_rca32_and_10_16_b_16;
  wire f_s_dadda_pg_rca32_and_10_16_y0;
  wire f_s_dadda_pg_rca32_and_9_17_a_9;
  wire f_s_dadda_pg_rca32_and_9_17_b_17;
  wire f_s_dadda_pg_rca32_and_9_17_y0;
  wire f_s_dadda_pg_rca32_and_8_18_a_8;
  wire f_s_dadda_pg_rca32_and_8_18_b_18;
  wire f_s_dadda_pg_rca32_and_8_18_y0;
  wire f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_10_16_y0;
  wire f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_9_17_y0;
  wire f_s_dadda_pg_rca32_fa218_y0;
  wire f_s_dadda_pg_rca32_fa218_y1;
  wire f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_8_18_y0;
  wire f_s_dadda_pg_rca32_fa218_y2;
  wire f_s_dadda_pg_rca32_fa218_y3;
  wire f_s_dadda_pg_rca32_fa218_y4;
  wire f_s_dadda_pg_rca32_and_7_19_a_7;
  wire f_s_dadda_pg_rca32_and_7_19_b_19;
  wire f_s_dadda_pg_rca32_and_7_19_y0;
  wire f_s_dadda_pg_rca32_and_6_20_a_6;
  wire f_s_dadda_pg_rca32_and_6_20_b_20;
  wire f_s_dadda_pg_rca32_and_6_20_y0;
  wire f_s_dadda_pg_rca32_and_5_21_a_5;
  wire f_s_dadda_pg_rca32_and_5_21_b_21;
  wire f_s_dadda_pg_rca32_and_5_21_y0;
  wire f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_7_19_y0;
  wire f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_6_20_y0;
  wire f_s_dadda_pg_rca32_fa219_y0;
  wire f_s_dadda_pg_rca32_fa219_y1;
  wire f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_5_21_y0;
  wire f_s_dadda_pg_rca32_fa219_y2;
  wire f_s_dadda_pg_rca32_fa219_y3;
  wire f_s_dadda_pg_rca32_fa219_y4;
  wire f_s_dadda_pg_rca32_and_4_22_a_4;
  wire f_s_dadda_pg_rca32_and_4_22_b_22;
  wire f_s_dadda_pg_rca32_and_4_22_y0;
  wire f_s_dadda_pg_rca32_and_3_23_a_3;
  wire f_s_dadda_pg_rca32_and_3_23_b_23;
  wire f_s_dadda_pg_rca32_and_3_23_y0;
  wire f_s_dadda_pg_rca32_and_2_24_a_2;
  wire f_s_dadda_pg_rca32_and_2_24_b_24;
  wire f_s_dadda_pg_rca32_and_2_24_y0;
  wire f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_4_22_y0;
  wire f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_3_23_y0;
  wire f_s_dadda_pg_rca32_fa220_y0;
  wire f_s_dadda_pg_rca32_fa220_y1;
  wire f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_2_24_y0;
  wire f_s_dadda_pg_rca32_fa220_y2;
  wire f_s_dadda_pg_rca32_fa220_y3;
  wire f_s_dadda_pg_rca32_fa220_y4;
  wire f_s_dadda_pg_rca32_and_1_25_a_1;
  wire f_s_dadda_pg_rca32_and_1_25_b_25;
  wire f_s_dadda_pg_rca32_and_1_25_y0;
  wire f_s_dadda_pg_rca32_and_0_26_a_0;
  wire f_s_dadda_pg_rca32_and_0_26_b_26;
  wire f_s_dadda_pg_rca32_and_0_26_y0;
  wire f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_and_1_25_y0;
  wire f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_and_0_26_y0;
  wire f_s_dadda_pg_rca32_fa221_y0;
  wire f_s_dadda_pg_rca32_fa221_y1;
  wire f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_fa206_y2;
  wire f_s_dadda_pg_rca32_fa221_y2;
  wire f_s_dadda_pg_rca32_fa221_y3;
  wire f_s_dadda_pg_rca32_fa221_y4;
  wire f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa207_y2;
  wire f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa208_y2;
  wire f_s_dadda_pg_rca32_fa222_y0;
  wire f_s_dadda_pg_rca32_fa222_y1;
  wire f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa209_y2;
  wire f_s_dadda_pg_rca32_fa222_y2;
  wire f_s_dadda_pg_rca32_fa222_y3;
  wire f_s_dadda_pg_rca32_fa222_y4;
  wire f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa210_y2;
  wire f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa211_y2;
  wire f_s_dadda_pg_rca32_fa223_y0;
  wire f_s_dadda_pg_rca32_fa223_y1;
  wire f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa212_y2;
  wire f_s_dadda_pg_rca32_fa223_y2;
  wire f_s_dadda_pg_rca32_fa223_y3;
  wire f_s_dadda_pg_rca32_fa223_y4;
  wire f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa213_y2;
  wire f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa214_y2;
  wire f_s_dadda_pg_rca32_fa224_y0;
  wire f_s_dadda_pg_rca32_fa224_y1;
  wire f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa215_y2;
  wire f_s_dadda_pg_rca32_fa224_y2;
  wire f_s_dadda_pg_rca32_fa224_y3;
  wire f_s_dadda_pg_rca32_fa224_y4;
  wire f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa216_y2;
  wire f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa217_y2;
  wire f_s_dadda_pg_rca32_fa225_y0;
  wire f_s_dadda_pg_rca32_fa225_y1;
  wire f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa218_y2;
  wire f_s_dadda_pg_rca32_fa225_y2;
  wire f_s_dadda_pg_rca32_fa225_y3;
  wire f_s_dadda_pg_rca32_fa225_y4;
  wire f_s_dadda_pg_rca32_ha24_f_s_dadda_pg_rca32_fa219_y2;
  wire f_s_dadda_pg_rca32_ha24_f_s_dadda_pg_rca32_fa220_y2;
  wire f_s_dadda_pg_rca32_ha24_y0;
  wire f_s_dadda_pg_rca32_ha24_y1;
  wire f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_ha24_y1;
  wire f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_fa225_y4;
  wire f_s_dadda_pg_rca32_fa226_y0;
  wire f_s_dadda_pg_rca32_fa226_y1;
  wire f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_fa224_y4;
  wire f_s_dadda_pg_rca32_fa226_y2;
  wire f_s_dadda_pg_rca32_fa226_y3;
  wire f_s_dadda_pg_rca32_fa226_y4;
  wire f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa223_y4;
  wire f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa222_y4;
  wire f_s_dadda_pg_rca32_fa227_y0;
  wire f_s_dadda_pg_rca32_fa227_y1;
  wire f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa221_y4;
  wire f_s_dadda_pg_rca32_fa227_y2;
  wire f_s_dadda_pg_rca32_fa227_y3;
  wire f_s_dadda_pg_rca32_fa227_y4;
  wire f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa220_y4;
  wire f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa219_y4;
  wire f_s_dadda_pg_rca32_fa228_y0;
  wire f_s_dadda_pg_rca32_fa228_y1;
  wire f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa218_y4;
  wire f_s_dadda_pg_rca32_fa228_y2;
  wire f_s_dadda_pg_rca32_fa228_y3;
  wire f_s_dadda_pg_rca32_fa228_y4;
  wire f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa217_y4;
  wire f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa216_y4;
  wire f_s_dadda_pg_rca32_fa229_y0;
  wire f_s_dadda_pg_rca32_fa229_y1;
  wire f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa215_y4;
  wire f_s_dadda_pg_rca32_fa229_y2;
  wire f_s_dadda_pg_rca32_fa229_y3;
  wire f_s_dadda_pg_rca32_fa229_y4;
  wire f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa214_y4;
  wire f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa213_y4;
  wire f_s_dadda_pg_rca32_fa230_y0;
  wire f_s_dadda_pg_rca32_fa230_y1;
  wire f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa212_y4;
  wire f_s_dadda_pg_rca32_fa230_y2;
  wire f_s_dadda_pg_rca32_fa230_y3;
  wire f_s_dadda_pg_rca32_fa230_y4;
  wire f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa211_y4;
  wire f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa210_y4;
  wire f_s_dadda_pg_rca32_fa231_y0;
  wire f_s_dadda_pg_rca32_fa231_y1;
  wire f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa209_y4;
  wire f_s_dadda_pg_rca32_fa231_y2;
  wire f_s_dadda_pg_rca32_fa231_y3;
  wire f_s_dadda_pg_rca32_fa231_y4;
  wire f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa208_y4;
  wire f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa207_y4;
  wire f_s_dadda_pg_rca32_fa232_y0;
  wire f_s_dadda_pg_rca32_fa232_y1;
  wire f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa206_y4;
  wire f_s_dadda_pg_rca32_fa232_y2;
  wire f_s_dadda_pg_rca32_fa232_y3;
  wire f_s_dadda_pg_rca32_fa232_y4;
  wire f_s_dadda_pg_rca32_and_27_0_a_27;
  wire f_s_dadda_pg_rca32_and_27_0_b_0;
  wire f_s_dadda_pg_rca32_and_27_0_y0;
  wire f_s_dadda_pg_rca32_and_26_1_a_26;
  wire f_s_dadda_pg_rca32_and_26_1_b_1;
  wire f_s_dadda_pg_rca32_and_26_1_y0;
  wire f_s_dadda_pg_rca32_and_25_2_a_25;
  wire f_s_dadda_pg_rca32_and_25_2_b_2;
  wire f_s_dadda_pg_rca32_and_25_2_y0;
  wire f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_27_0_y0;
  wire f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_26_1_y0;
  wire f_s_dadda_pg_rca32_fa233_y0;
  wire f_s_dadda_pg_rca32_fa233_y1;
  wire f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_25_2_y0;
  wire f_s_dadda_pg_rca32_fa233_y2;
  wire f_s_dadda_pg_rca32_fa233_y3;
  wire f_s_dadda_pg_rca32_fa233_y4;
  wire f_s_dadda_pg_rca32_and_24_3_a_24;
  wire f_s_dadda_pg_rca32_and_24_3_b_3;
  wire f_s_dadda_pg_rca32_and_24_3_y0;
  wire f_s_dadda_pg_rca32_and_23_4_a_23;
  wire f_s_dadda_pg_rca32_and_23_4_b_4;
  wire f_s_dadda_pg_rca32_and_23_4_y0;
  wire f_s_dadda_pg_rca32_and_22_5_a_22;
  wire f_s_dadda_pg_rca32_and_22_5_b_5;
  wire f_s_dadda_pg_rca32_and_22_5_y0;
  wire f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_24_3_y0;
  wire f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_23_4_y0;
  wire f_s_dadda_pg_rca32_fa234_y0;
  wire f_s_dadda_pg_rca32_fa234_y1;
  wire f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_22_5_y0;
  wire f_s_dadda_pg_rca32_fa234_y2;
  wire f_s_dadda_pg_rca32_fa234_y3;
  wire f_s_dadda_pg_rca32_fa234_y4;
  wire f_s_dadda_pg_rca32_and_21_6_a_21;
  wire f_s_dadda_pg_rca32_and_21_6_b_6;
  wire f_s_dadda_pg_rca32_and_21_6_y0;
  wire f_s_dadda_pg_rca32_and_20_7_a_20;
  wire f_s_dadda_pg_rca32_and_20_7_b_7;
  wire f_s_dadda_pg_rca32_and_20_7_y0;
  wire f_s_dadda_pg_rca32_and_19_8_a_19;
  wire f_s_dadda_pg_rca32_and_19_8_b_8;
  wire f_s_dadda_pg_rca32_and_19_8_y0;
  wire f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_21_6_y0;
  wire f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_20_7_y0;
  wire f_s_dadda_pg_rca32_fa235_y0;
  wire f_s_dadda_pg_rca32_fa235_y1;
  wire f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_19_8_y0;
  wire f_s_dadda_pg_rca32_fa235_y2;
  wire f_s_dadda_pg_rca32_fa235_y3;
  wire f_s_dadda_pg_rca32_fa235_y4;
  wire f_s_dadda_pg_rca32_and_18_9_a_18;
  wire f_s_dadda_pg_rca32_and_18_9_b_9;
  wire f_s_dadda_pg_rca32_and_18_9_y0;
  wire f_s_dadda_pg_rca32_and_17_10_a_17;
  wire f_s_dadda_pg_rca32_and_17_10_b_10;
  wire f_s_dadda_pg_rca32_and_17_10_y0;
  wire f_s_dadda_pg_rca32_and_16_11_a_16;
  wire f_s_dadda_pg_rca32_and_16_11_b_11;
  wire f_s_dadda_pg_rca32_and_16_11_y0;
  wire f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_18_9_y0;
  wire f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_17_10_y0;
  wire f_s_dadda_pg_rca32_fa236_y0;
  wire f_s_dadda_pg_rca32_fa236_y1;
  wire f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_16_11_y0;
  wire f_s_dadda_pg_rca32_fa236_y2;
  wire f_s_dadda_pg_rca32_fa236_y3;
  wire f_s_dadda_pg_rca32_fa236_y4;
  wire f_s_dadda_pg_rca32_and_15_12_a_15;
  wire f_s_dadda_pg_rca32_and_15_12_b_12;
  wire f_s_dadda_pg_rca32_and_15_12_y0;
  wire f_s_dadda_pg_rca32_and_14_13_a_14;
  wire f_s_dadda_pg_rca32_and_14_13_b_13;
  wire f_s_dadda_pg_rca32_and_14_13_y0;
  wire f_s_dadda_pg_rca32_and_13_14_a_13;
  wire f_s_dadda_pg_rca32_and_13_14_b_14;
  wire f_s_dadda_pg_rca32_and_13_14_y0;
  wire f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_15_12_y0;
  wire f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_14_13_y0;
  wire f_s_dadda_pg_rca32_fa237_y0;
  wire f_s_dadda_pg_rca32_fa237_y1;
  wire f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_13_14_y0;
  wire f_s_dadda_pg_rca32_fa237_y2;
  wire f_s_dadda_pg_rca32_fa237_y3;
  wire f_s_dadda_pg_rca32_fa237_y4;
  wire f_s_dadda_pg_rca32_and_12_15_a_12;
  wire f_s_dadda_pg_rca32_and_12_15_b_15;
  wire f_s_dadda_pg_rca32_and_12_15_y0;
  wire f_s_dadda_pg_rca32_and_11_16_a_11;
  wire f_s_dadda_pg_rca32_and_11_16_b_16;
  wire f_s_dadda_pg_rca32_and_11_16_y0;
  wire f_s_dadda_pg_rca32_and_10_17_a_10;
  wire f_s_dadda_pg_rca32_and_10_17_b_17;
  wire f_s_dadda_pg_rca32_and_10_17_y0;
  wire f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_12_15_y0;
  wire f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_11_16_y0;
  wire f_s_dadda_pg_rca32_fa238_y0;
  wire f_s_dadda_pg_rca32_fa238_y1;
  wire f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_10_17_y0;
  wire f_s_dadda_pg_rca32_fa238_y2;
  wire f_s_dadda_pg_rca32_fa238_y3;
  wire f_s_dadda_pg_rca32_fa238_y4;
  wire f_s_dadda_pg_rca32_and_9_18_a_9;
  wire f_s_dadda_pg_rca32_and_9_18_b_18;
  wire f_s_dadda_pg_rca32_and_9_18_y0;
  wire f_s_dadda_pg_rca32_and_8_19_a_8;
  wire f_s_dadda_pg_rca32_and_8_19_b_19;
  wire f_s_dadda_pg_rca32_and_8_19_y0;
  wire f_s_dadda_pg_rca32_and_7_20_a_7;
  wire f_s_dadda_pg_rca32_and_7_20_b_20;
  wire f_s_dadda_pg_rca32_and_7_20_y0;
  wire f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_9_18_y0;
  wire f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_8_19_y0;
  wire f_s_dadda_pg_rca32_fa239_y0;
  wire f_s_dadda_pg_rca32_fa239_y1;
  wire f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_7_20_y0;
  wire f_s_dadda_pg_rca32_fa239_y2;
  wire f_s_dadda_pg_rca32_fa239_y3;
  wire f_s_dadda_pg_rca32_fa239_y4;
  wire f_s_dadda_pg_rca32_and_6_21_a_6;
  wire f_s_dadda_pg_rca32_and_6_21_b_21;
  wire f_s_dadda_pg_rca32_and_6_21_y0;
  wire f_s_dadda_pg_rca32_and_5_22_a_5;
  wire f_s_dadda_pg_rca32_and_5_22_b_22;
  wire f_s_dadda_pg_rca32_and_5_22_y0;
  wire f_s_dadda_pg_rca32_and_4_23_a_4;
  wire f_s_dadda_pg_rca32_and_4_23_b_23;
  wire f_s_dadda_pg_rca32_and_4_23_y0;
  wire f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_6_21_y0;
  wire f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_5_22_y0;
  wire f_s_dadda_pg_rca32_fa240_y0;
  wire f_s_dadda_pg_rca32_fa240_y1;
  wire f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_4_23_y0;
  wire f_s_dadda_pg_rca32_fa240_y2;
  wire f_s_dadda_pg_rca32_fa240_y3;
  wire f_s_dadda_pg_rca32_fa240_y4;
  wire f_s_dadda_pg_rca32_and_3_24_a_3;
  wire f_s_dadda_pg_rca32_and_3_24_b_24;
  wire f_s_dadda_pg_rca32_and_3_24_y0;
  wire f_s_dadda_pg_rca32_and_2_25_a_2;
  wire f_s_dadda_pg_rca32_and_2_25_b_25;
  wire f_s_dadda_pg_rca32_and_2_25_y0;
  wire f_s_dadda_pg_rca32_and_1_26_a_1;
  wire f_s_dadda_pg_rca32_and_1_26_b_26;
  wire f_s_dadda_pg_rca32_and_1_26_y0;
  wire f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_3_24_y0;
  wire f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_2_25_y0;
  wire f_s_dadda_pg_rca32_fa241_y0;
  wire f_s_dadda_pg_rca32_fa241_y1;
  wire f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_1_26_y0;
  wire f_s_dadda_pg_rca32_fa241_y2;
  wire f_s_dadda_pg_rca32_fa241_y3;
  wire f_s_dadda_pg_rca32_fa241_y4;
  wire f_s_dadda_pg_rca32_and_0_27_a_0;
  wire f_s_dadda_pg_rca32_and_0_27_b_27;
  wire f_s_dadda_pg_rca32_and_0_27_y0;
  wire f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_and_0_27_y0;
  wire f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_fa226_y2;
  wire f_s_dadda_pg_rca32_fa242_y0;
  wire f_s_dadda_pg_rca32_fa242_y1;
  wire f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_fa227_y2;
  wire f_s_dadda_pg_rca32_fa242_y2;
  wire f_s_dadda_pg_rca32_fa242_y3;
  wire f_s_dadda_pg_rca32_fa242_y4;
  wire f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa228_y2;
  wire f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa229_y2;
  wire f_s_dadda_pg_rca32_fa243_y0;
  wire f_s_dadda_pg_rca32_fa243_y1;
  wire f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa230_y2;
  wire f_s_dadda_pg_rca32_fa243_y2;
  wire f_s_dadda_pg_rca32_fa243_y3;
  wire f_s_dadda_pg_rca32_fa243_y4;
  wire f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa231_y2;
  wire f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa232_y2;
  wire f_s_dadda_pg_rca32_fa244_y0;
  wire f_s_dadda_pg_rca32_fa244_y1;
  wire f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa233_y2;
  wire f_s_dadda_pg_rca32_fa244_y2;
  wire f_s_dadda_pg_rca32_fa244_y3;
  wire f_s_dadda_pg_rca32_fa244_y4;
  wire f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa234_y2;
  wire f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa235_y2;
  wire f_s_dadda_pg_rca32_fa245_y0;
  wire f_s_dadda_pg_rca32_fa245_y1;
  wire f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa236_y2;
  wire f_s_dadda_pg_rca32_fa245_y2;
  wire f_s_dadda_pg_rca32_fa245_y3;
  wire f_s_dadda_pg_rca32_fa245_y4;
  wire f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa237_y2;
  wire f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa238_y2;
  wire f_s_dadda_pg_rca32_fa246_y0;
  wire f_s_dadda_pg_rca32_fa246_y1;
  wire f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa239_y2;
  wire f_s_dadda_pg_rca32_fa246_y2;
  wire f_s_dadda_pg_rca32_fa246_y3;
  wire f_s_dadda_pg_rca32_fa246_y4;
  wire f_s_dadda_pg_rca32_ha25_f_s_dadda_pg_rca32_fa240_y2;
  wire f_s_dadda_pg_rca32_ha25_f_s_dadda_pg_rca32_fa241_y2;
  wire f_s_dadda_pg_rca32_ha25_y0;
  wire f_s_dadda_pg_rca32_ha25_y1;
  wire f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_ha25_y1;
  wire f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_fa246_y4;
  wire f_s_dadda_pg_rca32_fa247_y0;
  wire f_s_dadda_pg_rca32_fa247_y1;
  wire f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_fa245_y4;
  wire f_s_dadda_pg_rca32_fa247_y2;
  wire f_s_dadda_pg_rca32_fa247_y3;
  wire f_s_dadda_pg_rca32_fa247_y4;
  wire f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa244_y4;
  wire f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa243_y4;
  wire f_s_dadda_pg_rca32_fa248_y0;
  wire f_s_dadda_pg_rca32_fa248_y1;
  wire f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa242_y4;
  wire f_s_dadda_pg_rca32_fa248_y2;
  wire f_s_dadda_pg_rca32_fa248_y3;
  wire f_s_dadda_pg_rca32_fa248_y4;
  wire f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa241_y4;
  wire f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa240_y4;
  wire f_s_dadda_pg_rca32_fa249_y0;
  wire f_s_dadda_pg_rca32_fa249_y1;
  wire f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa239_y4;
  wire f_s_dadda_pg_rca32_fa249_y2;
  wire f_s_dadda_pg_rca32_fa249_y3;
  wire f_s_dadda_pg_rca32_fa249_y4;
  wire f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa238_y4;
  wire f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa237_y4;
  wire f_s_dadda_pg_rca32_fa250_y0;
  wire f_s_dadda_pg_rca32_fa250_y1;
  wire f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa236_y4;
  wire f_s_dadda_pg_rca32_fa250_y2;
  wire f_s_dadda_pg_rca32_fa250_y3;
  wire f_s_dadda_pg_rca32_fa250_y4;
  wire f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa235_y4;
  wire f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa234_y4;
  wire f_s_dadda_pg_rca32_fa251_y0;
  wire f_s_dadda_pg_rca32_fa251_y1;
  wire f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa233_y4;
  wire f_s_dadda_pg_rca32_fa251_y2;
  wire f_s_dadda_pg_rca32_fa251_y3;
  wire f_s_dadda_pg_rca32_fa251_y4;
  wire f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa232_y4;
  wire f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa231_y4;
  wire f_s_dadda_pg_rca32_fa252_y0;
  wire f_s_dadda_pg_rca32_fa252_y1;
  wire f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa230_y4;
  wire f_s_dadda_pg_rca32_fa252_y2;
  wire f_s_dadda_pg_rca32_fa252_y3;
  wire f_s_dadda_pg_rca32_fa252_y4;
  wire f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa229_y4;
  wire f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa228_y4;
  wire f_s_dadda_pg_rca32_fa253_y0;
  wire f_s_dadda_pg_rca32_fa253_y1;
  wire f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa227_y4;
  wire f_s_dadda_pg_rca32_fa253_y2;
  wire f_s_dadda_pg_rca32_fa253_y3;
  wire f_s_dadda_pg_rca32_fa253_y4;
  wire f_s_dadda_pg_rca32_and_26_2_a_26;
  wire f_s_dadda_pg_rca32_and_26_2_b_2;
  wire f_s_dadda_pg_rca32_and_26_2_y0;
  wire f_s_dadda_pg_rca32_and_25_3_a_25;
  wire f_s_dadda_pg_rca32_and_25_3_b_3;
  wire f_s_dadda_pg_rca32_and_25_3_y0;
  wire f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_fa226_y4;
  wire f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_and_26_2_y0;
  wire f_s_dadda_pg_rca32_fa254_y0;
  wire f_s_dadda_pg_rca32_fa254_y1;
  wire f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_and_25_3_y0;
  wire f_s_dadda_pg_rca32_fa254_y2;
  wire f_s_dadda_pg_rca32_fa254_y3;
  wire f_s_dadda_pg_rca32_fa254_y4;
  wire f_s_dadda_pg_rca32_and_24_4_a_24;
  wire f_s_dadda_pg_rca32_and_24_4_b_4;
  wire f_s_dadda_pg_rca32_and_24_4_y0;
  wire f_s_dadda_pg_rca32_and_23_5_a_23;
  wire f_s_dadda_pg_rca32_and_23_5_b_5;
  wire f_s_dadda_pg_rca32_and_23_5_y0;
  wire f_s_dadda_pg_rca32_and_22_6_a_22;
  wire f_s_dadda_pg_rca32_and_22_6_b_6;
  wire f_s_dadda_pg_rca32_and_22_6_y0;
  wire f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_24_4_y0;
  wire f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_23_5_y0;
  wire f_s_dadda_pg_rca32_fa255_y0;
  wire f_s_dadda_pg_rca32_fa255_y1;
  wire f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_22_6_y0;
  wire f_s_dadda_pg_rca32_fa255_y2;
  wire f_s_dadda_pg_rca32_fa255_y3;
  wire f_s_dadda_pg_rca32_fa255_y4;
  wire f_s_dadda_pg_rca32_and_21_7_a_21;
  wire f_s_dadda_pg_rca32_and_21_7_b_7;
  wire f_s_dadda_pg_rca32_and_21_7_y0;
  wire f_s_dadda_pg_rca32_and_20_8_a_20;
  wire f_s_dadda_pg_rca32_and_20_8_b_8;
  wire f_s_dadda_pg_rca32_and_20_8_y0;
  wire f_s_dadda_pg_rca32_and_19_9_a_19;
  wire f_s_dadda_pg_rca32_and_19_9_b_9;
  wire f_s_dadda_pg_rca32_and_19_9_y0;
  wire f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_21_7_y0;
  wire f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_20_8_y0;
  wire f_s_dadda_pg_rca32_fa256_y0;
  wire f_s_dadda_pg_rca32_fa256_y1;
  wire f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_19_9_y0;
  wire f_s_dadda_pg_rca32_fa256_y2;
  wire f_s_dadda_pg_rca32_fa256_y3;
  wire f_s_dadda_pg_rca32_fa256_y4;
  wire f_s_dadda_pg_rca32_and_18_10_a_18;
  wire f_s_dadda_pg_rca32_and_18_10_b_10;
  wire f_s_dadda_pg_rca32_and_18_10_y0;
  wire f_s_dadda_pg_rca32_and_17_11_a_17;
  wire f_s_dadda_pg_rca32_and_17_11_b_11;
  wire f_s_dadda_pg_rca32_and_17_11_y0;
  wire f_s_dadda_pg_rca32_and_16_12_a_16;
  wire f_s_dadda_pg_rca32_and_16_12_b_12;
  wire f_s_dadda_pg_rca32_and_16_12_y0;
  wire f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_18_10_y0;
  wire f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_17_11_y0;
  wire f_s_dadda_pg_rca32_fa257_y0;
  wire f_s_dadda_pg_rca32_fa257_y1;
  wire f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_16_12_y0;
  wire f_s_dadda_pg_rca32_fa257_y2;
  wire f_s_dadda_pg_rca32_fa257_y3;
  wire f_s_dadda_pg_rca32_fa257_y4;
  wire f_s_dadda_pg_rca32_and_15_13_a_15;
  wire f_s_dadda_pg_rca32_and_15_13_b_13;
  wire f_s_dadda_pg_rca32_and_15_13_y0;
  wire f_s_dadda_pg_rca32_and_14_14_a_14;
  wire f_s_dadda_pg_rca32_and_14_14_b_14;
  wire f_s_dadda_pg_rca32_and_14_14_y0;
  wire f_s_dadda_pg_rca32_and_13_15_a_13;
  wire f_s_dadda_pg_rca32_and_13_15_b_15;
  wire f_s_dadda_pg_rca32_and_13_15_y0;
  wire f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_15_13_y0;
  wire f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_14_14_y0;
  wire f_s_dadda_pg_rca32_fa258_y0;
  wire f_s_dadda_pg_rca32_fa258_y1;
  wire f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_13_15_y0;
  wire f_s_dadda_pg_rca32_fa258_y2;
  wire f_s_dadda_pg_rca32_fa258_y3;
  wire f_s_dadda_pg_rca32_fa258_y4;
  wire f_s_dadda_pg_rca32_and_12_16_a_12;
  wire f_s_dadda_pg_rca32_and_12_16_b_16;
  wire f_s_dadda_pg_rca32_and_12_16_y0;
  wire f_s_dadda_pg_rca32_and_11_17_a_11;
  wire f_s_dadda_pg_rca32_and_11_17_b_17;
  wire f_s_dadda_pg_rca32_and_11_17_y0;
  wire f_s_dadda_pg_rca32_and_10_18_a_10;
  wire f_s_dadda_pg_rca32_and_10_18_b_18;
  wire f_s_dadda_pg_rca32_and_10_18_y0;
  wire f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_12_16_y0;
  wire f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_11_17_y0;
  wire f_s_dadda_pg_rca32_fa259_y0;
  wire f_s_dadda_pg_rca32_fa259_y1;
  wire f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_10_18_y0;
  wire f_s_dadda_pg_rca32_fa259_y2;
  wire f_s_dadda_pg_rca32_fa259_y3;
  wire f_s_dadda_pg_rca32_fa259_y4;
  wire f_s_dadda_pg_rca32_and_9_19_a_9;
  wire f_s_dadda_pg_rca32_and_9_19_b_19;
  wire f_s_dadda_pg_rca32_and_9_19_y0;
  wire f_s_dadda_pg_rca32_and_8_20_a_8;
  wire f_s_dadda_pg_rca32_and_8_20_b_20;
  wire f_s_dadda_pg_rca32_and_8_20_y0;
  wire f_s_dadda_pg_rca32_and_7_21_a_7;
  wire f_s_dadda_pg_rca32_and_7_21_b_21;
  wire f_s_dadda_pg_rca32_and_7_21_y0;
  wire f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_9_19_y0;
  wire f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_8_20_y0;
  wire f_s_dadda_pg_rca32_fa260_y0;
  wire f_s_dadda_pg_rca32_fa260_y1;
  wire f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_7_21_y0;
  wire f_s_dadda_pg_rca32_fa260_y2;
  wire f_s_dadda_pg_rca32_fa260_y3;
  wire f_s_dadda_pg_rca32_fa260_y4;
  wire f_s_dadda_pg_rca32_and_6_22_a_6;
  wire f_s_dadda_pg_rca32_and_6_22_b_22;
  wire f_s_dadda_pg_rca32_and_6_22_y0;
  wire f_s_dadda_pg_rca32_and_5_23_a_5;
  wire f_s_dadda_pg_rca32_and_5_23_b_23;
  wire f_s_dadda_pg_rca32_and_5_23_y0;
  wire f_s_dadda_pg_rca32_and_4_24_a_4;
  wire f_s_dadda_pg_rca32_and_4_24_b_24;
  wire f_s_dadda_pg_rca32_and_4_24_y0;
  wire f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_6_22_y0;
  wire f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_5_23_y0;
  wire f_s_dadda_pg_rca32_fa261_y0;
  wire f_s_dadda_pg_rca32_fa261_y1;
  wire f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_4_24_y0;
  wire f_s_dadda_pg_rca32_fa261_y2;
  wire f_s_dadda_pg_rca32_fa261_y3;
  wire f_s_dadda_pg_rca32_fa261_y4;
  wire f_s_dadda_pg_rca32_and_3_25_a_3;
  wire f_s_dadda_pg_rca32_and_3_25_b_25;
  wire f_s_dadda_pg_rca32_and_3_25_y0;
  wire f_s_dadda_pg_rca32_and_2_26_a_2;
  wire f_s_dadda_pg_rca32_and_2_26_b_26;
  wire f_s_dadda_pg_rca32_and_2_26_y0;
  wire f_s_dadda_pg_rca32_and_1_27_a_1;
  wire f_s_dadda_pg_rca32_and_1_27_b_27;
  wire f_s_dadda_pg_rca32_and_1_27_y0;
  wire f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_3_25_y0;
  wire f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_2_26_y0;
  wire f_s_dadda_pg_rca32_fa262_y0;
  wire f_s_dadda_pg_rca32_fa262_y1;
  wire f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_1_27_y0;
  wire f_s_dadda_pg_rca32_fa262_y2;
  wire f_s_dadda_pg_rca32_fa262_y3;
  wire f_s_dadda_pg_rca32_fa262_y4;
  wire f_s_dadda_pg_rca32_and_0_28_a_0;
  wire f_s_dadda_pg_rca32_and_0_28_b_28;
  wire f_s_dadda_pg_rca32_and_0_28_y0;
  wire f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_and_0_28_y0;
  wire f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_ha0_y0;
  wire f_s_dadda_pg_rca32_fa263_y0;
  wire f_s_dadda_pg_rca32_fa263_y1;
  wire f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_fa247_y2;
  wire f_s_dadda_pg_rca32_fa263_y2;
  wire f_s_dadda_pg_rca32_fa263_y3;
  wire f_s_dadda_pg_rca32_fa263_y4;
  wire f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa248_y2;
  wire f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa249_y2;
  wire f_s_dadda_pg_rca32_fa264_y0;
  wire f_s_dadda_pg_rca32_fa264_y1;
  wire f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa250_y2;
  wire f_s_dadda_pg_rca32_fa264_y2;
  wire f_s_dadda_pg_rca32_fa264_y3;
  wire f_s_dadda_pg_rca32_fa264_y4;
  wire f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa251_y2;
  wire f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa252_y2;
  wire f_s_dadda_pg_rca32_fa265_y0;
  wire f_s_dadda_pg_rca32_fa265_y1;
  wire f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa253_y2;
  wire f_s_dadda_pg_rca32_fa265_y2;
  wire f_s_dadda_pg_rca32_fa265_y3;
  wire f_s_dadda_pg_rca32_fa265_y4;
  wire f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa254_y2;
  wire f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa255_y2;
  wire f_s_dadda_pg_rca32_fa266_y0;
  wire f_s_dadda_pg_rca32_fa266_y1;
  wire f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa256_y2;
  wire f_s_dadda_pg_rca32_fa266_y2;
  wire f_s_dadda_pg_rca32_fa266_y3;
  wire f_s_dadda_pg_rca32_fa266_y4;
  wire f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa257_y2;
  wire f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa258_y2;
  wire f_s_dadda_pg_rca32_fa267_y0;
  wire f_s_dadda_pg_rca32_fa267_y1;
  wire f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa259_y2;
  wire f_s_dadda_pg_rca32_fa267_y2;
  wire f_s_dadda_pg_rca32_fa267_y3;
  wire f_s_dadda_pg_rca32_fa267_y4;
  wire f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa260_y2;
  wire f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa261_y2;
  wire f_s_dadda_pg_rca32_fa268_y0;
  wire f_s_dadda_pg_rca32_fa268_y1;
  wire f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa262_y2;
  wire f_s_dadda_pg_rca32_fa268_y2;
  wire f_s_dadda_pg_rca32_fa268_y3;
  wire f_s_dadda_pg_rca32_fa268_y4;
  wire f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa268_y4;
  wire f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa267_y4;
  wire f_s_dadda_pg_rca32_fa269_y0;
  wire f_s_dadda_pg_rca32_fa269_y1;
  wire f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa266_y4;
  wire f_s_dadda_pg_rca32_fa269_y2;
  wire f_s_dadda_pg_rca32_fa269_y3;
  wire f_s_dadda_pg_rca32_fa269_y4;
  wire f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa265_y4;
  wire f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa264_y4;
  wire f_s_dadda_pg_rca32_fa270_y0;
  wire f_s_dadda_pg_rca32_fa270_y1;
  wire f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa263_y4;
  wire f_s_dadda_pg_rca32_fa270_y2;
  wire f_s_dadda_pg_rca32_fa270_y3;
  wire f_s_dadda_pg_rca32_fa270_y4;
  wire f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa262_y4;
  wire f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa261_y4;
  wire f_s_dadda_pg_rca32_fa271_y0;
  wire f_s_dadda_pg_rca32_fa271_y1;
  wire f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa260_y4;
  wire f_s_dadda_pg_rca32_fa271_y2;
  wire f_s_dadda_pg_rca32_fa271_y3;
  wire f_s_dadda_pg_rca32_fa271_y4;
  wire f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa259_y4;
  wire f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa258_y4;
  wire f_s_dadda_pg_rca32_fa272_y0;
  wire f_s_dadda_pg_rca32_fa272_y1;
  wire f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa257_y4;
  wire f_s_dadda_pg_rca32_fa272_y2;
  wire f_s_dadda_pg_rca32_fa272_y3;
  wire f_s_dadda_pg_rca32_fa272_y4;
  wire f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa256_y4;
  wire f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa255_y4;
  wire f_s_dadda_pg_rca32_fa273_y0;
  wire f_s_dadda_pg_rca32_fa273_y1;
  wire f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa254_y4;
  wire f_s_dadda_pg_rca32_fa273_y2;
  wire f_s_dadda_pg_rca32_fa273_y3;
  wire f_s_dadda_pg_rca32_fa273_y4;
  wire f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa253_y4;
  wire f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa252_y4;
  wire f_s_dadda_pg_rca32_fa274_y0;
  wire f_s_dadda_pg_rca32_fa274_y1;
  wire f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa251_y4;
  wire f_s_dadda_pg_rca32_fa274_y2;
  wire f_s_dadda_pg_rca32_fa274_y3;
  wire f_s_dadda_pg_rca32_fa274_y4;
  wire f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa250_y4;
  wire f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa249_y4;
  wire f_s_dadda_pg_rca32_fa275_y0;
  wire f_s_dadda_pg_rca32_fa275_y1;
  wire f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa248_y4;
  wire f_s_dadda_pg_rca32_fa275_y2;
  wire f_s_dadda_pg_rca32_fa275_y3;
  wire f_s_dadda_pg_rca32_fa275_y4;
  wire f_s_dadda_pg_rca32_and_25_4_a_25;
  wire f_s_dadda_pg_rca32_and_25_4_b_4;
  wire f_s_dadda_pg_rca32_and_25_4_y0;
  wire f_s_dadda_pg_rca32_and_24_5_a_24;
  wire f_s_dadda_pg_rca32_and_24_5_b_5;
  wire f_s_dadda_pg_rca32_and_24_5_y0;
  wire f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_fa247_y4;
  wire f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_and_25_4_y0;
  wire f_s_dadda_pg_rca32_fa276_y0;
  wire f_s_dadda_pg_rca32_fa276_y1;
  wire f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_and_24_5_y0;
  wire f_s_dadda_pg_rca32_fa276_y2;
  wire f_s_dadda_pg_rca32_fa276_y3;
  wire f_s_dadda_pg_rca32_fa276_y4;
  wire f_s_dadda_pg_rca32_and_23_6_a_23;
  wire f_s_dadda_pg_rca32_and_23_6_b_6;
  wire f_s_dadda_pg_rca32_and_23_6_y0;
  wire f_s_dadda_pg_rca32_and_22_7_a_22;
  wire f_s_dadda_pg_rca32_and_22_7_b_7;
  wire f_s_dadda_pg_rca32_and_22_7_y0;
  wire f_s_dadda_pg_rca32_and_21_8_a_21;
  wire f_s_dadda_pg_rca32_and_21_8_b_8;
  wire f_s_dadda_pg_rca32_and_21_8_y0;
  wire f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_23_6_y0;
  wire f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_22_7_y0;
  wire f_s_dadda_pg_rca32_fa277_y0;
  wire f_s_dadda_pg_rca32_fa277_y1;
  wire f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_21_8_y0;
  wire f_s_dadda_pg_rca32_fa277_y2;
  wire f_s_dadda_pg_rca32_fa277_y3;
  wire f_s_dadda_pg_rca32_fa277_y4;
  wire f_s_dadda_pg_rca32_and_20_9_a_20;
  wire f_s_dadda_pg_rca32_and_20_9_b_9;
  wire f_s_dadda_pg_rca32_and_20_9_y0;
  wire f_s_dadda_pg_rca32_and_19_10_a_19;
  wire f_s_dadda_pg_rca32_and_19_10_b_10;
  wire f_s_dadda_pg_rca32_and_19_10_y0;
  wire f_s_dadda_pg_rca32_and_18_11_a_18;
  wire f_s_dadda_pg_rca32_and_18_11_b_11;
  wire f_s_dadda_pg_rca32_and_18_11_y0;
  wire f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_20_9_y0;
  wire f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_19_10_y0;
  wire f_s_dadda_pg_rca32_fa278_y0;
  wire f_s_dadda_pg_rca32_fa278_y1;
  wire f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_18_11_y0;
  wire f_s_dadda_pg_rca32_fa278_y2;
  wire f_s_dadda_pg_rca32_fa278_y3;
  wire f_s_dadda_pg_rca32_fa278_y4;
  wire f_s_dadda_pg_rca32_and_17_12_a_17;
  wire f_s_dadda_pg_rca32_and_17_12_b_12;
  wire f_s_dadda_pg_rca32_and_17_12_y0;
  wire f_s_dadda_pg_rca32_and_16_13_a_16;
  wire f_s_dadda_pg_rca32_and_16_13_b_13;
  wire f_s_dadda_pg_rca32_and_16_13_y0;
  wire f_s_dadda_pg_rca32_and_15_14_a_15;
  wire f_s_dadda_pg_rca32_and_15_14_b_14;
  wire f_s_dadda_pg_rca32_and_15_14_y0;
  wire f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_17_12_y0;
  wire f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_16_13_y0;
  wire f_s_dadda_pg_rca32_fa279_y0;
  wire f_s_dadda_pg_rca32_fa279_y1;
  wire f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_15_14_y0;
  wire f_s_dadda_pg_rca32_fa279_y2;
  wire f_s_dadda_pg_rca32_fa279_y3;
  wire f_s_dadda_pg_rca32_fa279_y4;
  wire f_s_dadda_pg_rca32_and_14_15_a_14;
  wire f_s_dadda_pg_rca32_and_14_15_b_15;
  wire f_s_dadda_pg_rca32_and_14_15_y0;
  wire f_s_dadda_pg_rca32_and_13_16_a_13;
  wire f_s_dadda_pg_rca32_and_13_16_b_16;
  wire f_s_dadda_pg_rca32_and_13_16_y0;
  wire f_s_dadda_pg_rca32_and_12_17_a_12;
  wire f_s_dadda_pg_rca32_and_12_17_b_17;
  wire f_s_dadda_pg_rca32_and_12_17_y0;
  wire f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_14_15_y0;
  wire f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_13_16_y0;
  wire f_s_dadda_pg_rca32_fa280_y0;
  wire f_s_dadda_pg_rca32_fa280_y1;
  wire f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_12_17_y0;
  wire f_s_dadda_pg_rca32_fa280_y2;
  wire f_s_dadda_pg_rca32_fa280_y3;
  wire f_s_dadda_pg_rca32_fa280_y4;
  wire f_s_dadda_pg_rca32_and_11_18_a_11;
  wire f_s_dadda_pg_rca32_and_11_18_b_18;
  wire f_s_dadda_pg_rca32_and_11_18_y0;
  wire f_s_dadda_pg_rca32_and_10_19_a_10;
  wire f_s_dadda_pg_rca32_and_10_19_b_19;
  wire f_s_dadda_pg_rca32_and_10_19_y0;
  wire f_s_dadda_pg_rca32_and_9_20_a_9;
  wire f_s_dadda_pg_rca32_and_9_20_b_20;
  wire f_s_dadda_pg_rca32_and_9_20_y0;
  wire f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_11_18_y0;
  wire f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_10_19_y0;
  wire f_s_dadda_pg_rca32_fa281_y0;
  wire f_s_dadda_pg_rca32_fa281_y1;
  wire f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_9_20_y0;
  wire f_s_dadda_pg_rca32_fa281_y2;
  wire f_s_dadda_pg_rca32_fa281_y3;
  wire f_s_dadda_pg_rca32_fa281_y4;
  wire f_s_dadda_pg_rca32_and_8_21_a_8;
  wire f_s_dadda_pg_rca32_and_8_21_b_21;
  wire f_s_dadda_pg_rca32_and_8_21_y0;
  wire f_s_dadda_pg_rca32_and_7_22_a_7;
  wire f_s_dadda_pg_rca32_and_7_22_b_22;
  wire f_s_dadda_pg_rca32_and_7_22_y0;
  wire f_s_dadda_pg_rca32_and_6_23_a_6;
  wire f_s_dadda_pg_rca32_and_6_23_b_23;
  wire f_s_dadda_pg_rca32_and_6_23_y0;
  wire f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_8_21_y0;
  wire f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_7_22_y0;
  wire f_s_dadda_pg_rca32_fa282_y0;
  wire f_s_dadda_pg_rca32_fa282_y1;
  wire f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_6_23_y0;
  wire f_s_dadda_pg_rca32_fa282_y2;
  wire f_s_dadda_pg_rca32_fa282_y3;
  wire f_s_dadda_pg_rca32_fa282_y4;
  wire f_s_dadda_pg_rca32_and_5_24_a_5;
  wire f_s_dadda_pg_rca32_and_5_24_b_24;
  wire f_s_dadda_pg_rca32_and_5_24_y0;
  wire f_s_dadda_pg_rca32_and_4_25_a_4;
  wire f_s_dadda_pg_rca32_and_4_25_b_25;
  wire f_s_dadda_pg_rca32_and_4_25_y0;
  wire f_s_dadda_pg_rca32_and_3_26_a_3;
  wire f_s_dadda_pg_rca32_and_3_26_b_26;
  wire f_s_dadda_pg_rca32_and_3_26_y0;
  wire f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_5_24_y0;
  wire f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_4_25_y0;
  wire f_s_dadda_pg_rca32_fa283_y0;
  wire f_s_dadda_pg_rca32_fa283_y1;
  wire f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_3_26_y0;
  wire f_s_dadda_pg_rca32_fa283_y2;
  wire f_s_dadda_pg_rca32_fa283_y3;
  wire f_s_dadda_pg_rca32_fa283_y4;
  wire f_s_dadda_pg_rca32_and_2_27_a_2;
  wire f_s_dadda_pg_rca32_and_2_27_b_27;
  wire f_s_dadda_pg_rca32_and_2_27_y0;
  wire f_s_dadda_pg_rca32_and_1_28_a_1;
  wire f_s_dadda_pg_rca32_and_1_28_b_28;
  wire f_s_dadda_pg_rca32_and_1_28_y0;
  wire f_s_dadda_pg_rca32_and_0_29_a_0;
  wire f_s_dadda_pg_rca32_and_0_29_b_29;
  wire f_s_dadda_pg_rca32_and_0_29_y0;
  wire f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_2_27_y0;
  wire f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_1_28_y0;
  wire f_s_dadda_pg_rca32_fa284_y0;
  wire f_s_dadda_pg_rca32_fa284_y1;
  wire f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_0_29_y0;
  wire f_s_dadda_pg_rca32_fa284_y2;
  wire f_s_dadda_pg_rca32_fa284_y3;
  wire f_s_dadda_pg_rca32_fa284_y4;
  wire f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_fa0_y2;
  wire f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_ha1_y0;
  wire f_s_dadda_pg_rca32_fa285_y0;
  wire f_s_dadda_pg_rca32_fa285_y1;
  wire f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_fa269_y2;
  wire f_s_dadda_pg_rca32_fa285_y2;
  wire f_s_dadda_pg_rca32_fa285_y3;
  wire f_s_dadda_pg_rca32_fa285_y4;
  wire f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa270_y2;
  wire f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa271_y2;
  wire f_s_dadda_pg_rca32_fa286_y0;
  wire f_s_dadda_pg_rca32_fa286_y1;
  wire f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa272_y2;
  wire f_s_dadda_pg_rca32_fa286_y2;
  wire f_s_dadda_pg_rca32_fa286_y3;
  wire f_s_dadda_pg_rca32_fa286_y4;
  wire f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa273_y2;
  wire f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa274_y2;
  wire f_s_dadda_pg_rca32_fa287_y0;
  wire f_s_dadda_pg_rca32_fa287_y1;
  wire f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa275_y2;
  wire f_s_dadda_pg_rca32_fa287_y2;
  wire f_s_dadda_pg_rca32_fa287_y3;
  wire f_s_dadda_pg_rca32_fa287_y4;
  wire f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa276_y2;
  wire f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa277_y2;
  wire f_s_dadda_pg_rca32_fa288_y0;
  wire f_s_dadda_pg_rca32_fa288_y1;
  wire f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa278_y2;
  wire f_s_dadda_pg_rca32_fa288_y2;
  wire f_s_dadda_pg_rca32_fa288_y3;
  wire f_s_dadda_pg_rca32_fa288_y4;
  wire f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa279_y2;
  wire f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa280_y2;
  wire f_s_dadda_pg_rca32_fa289_y0;
  wire f_s_dadda_pg_rca32_fa289_y1;
  wire f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa281_y2;
  wire f_s_dadda_pg_rca32_fa289_y2;
  wire f_s_dadda_pg_rca32_fa289_y3;
  wire f_s_dadda_pg_rca32_fa289_y4;
  wire f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa282_y2;
  wire f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa283_y2;
  wire f_s_dadda_pg_rca32_fa290_y0;
  wire f_s_dadda_pg_rca32_fa290_y1;
  wire f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa284_y2;
  wire f_s_dadda_pg_rca32_fa290_y2;
  wire f_s_dadda_pg_rca32_fa290_y3;
  wire f_s_dadda_pg_rca32_fa290_y4;
  wire f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa290_y4;
  wire f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa289_y4;
  wire f_s_dadda_pg_rca32_fa291_y0;
  wire f_s_dadda_pg_rca32_fa291_y1;
  wire f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa288_y4;
  wire f_s_dadda_pg_rca32_fa291_y2;
  wire f_s_dadda_pg_rca32_fa291_y3;
  wire f_s_dadda_pg_rca32_fa291_y4;
  wire f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa287_y4;
  wire f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa286_y4;
  wire f_s_dadda_pg_rca32_fa292_y0;
  wire f_s_dadda_pg_rca32_fa292_y1;
  wire f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa285_y4;
  wire f_s_dadda_pg_rca32_fa292_y2;
  wire f_s_dadda_pg_rca32_fa292_y3;
  wire f_s_dadda_pg_rca32_fa292_y4;
  wire f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa284_y4;
  wire f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa283_y4;
  wire f_s_dadda_pg_rca32_fa293_y0;
  wire f_s_dadda_pg_rca32_fa293_y1;
  wire f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa282_y4;
  wire f_s_dadda_pg_rca32_fa293_y2;
  wire f_s_dadda_pg_rca32_fa293_y3;
  wire f_s_dadda_pg_rca32_fa293_y4;
  wire f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa281_y4;
  wire f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa280_y4;
  wire f_s_dadda_pg_rca32_fa294_y0;
  wire f_s_dadda_pg_rca32_fa294_y1;
  wire f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa279_y4;
  wire f_s_dadda_pg_rca32_fa294_y2;
  wire f_s_dadda_pg_rca32_fa294_y3;
  wire f_s_dadda_pg_rca32_fa294_y4;
  wire f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa278_y4;
  wire f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa277_y4;
  wire f_s_dadda_pg_rca32_fa295_y0;
  wire f_s_dadda_pg_rca32_fa295_y1;
  wire f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa276_y4;
  wire f_s_dadda_pg_rca32_fa295_y2;
  wire f_s_dadda_pg_rca32_fa295_y3;
  wire f_s_dadda_pg_rca32_fa295_y4;
  wire f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa275_y4;
  wire f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa274_y4;
  wire f_s_dadda_pg_rca32_fa296_y0;
  wire f_s_dadda_pg_rca32_fa296_y1;
  wire f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa273_y4;
  wire f_s_dadda_pg_rca32_fa296_y2;
  wire f_s_dadda_pg_rca32_fa296_y3;
  wire f_s_dadda_pg_rca32_fa296_y4;
  wire f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa272_y4;
  wire f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa271_y4;
  wire f_s_dadda_pg_rca32_fa297_y0;
  wire f_s_dadda_pg_rca32_fa297_y1;
  wire f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa270_y4;
  wire f_s_dadda_pg_rca32_fa297_y2;
  wire f_s_dadda_pg_rca32_fa297_y3;
  wire f_s_dadda_pg_rca32_fa297_y4;
  wire f_s_dadda_pg_rca32_and_24_6_a_24;
  wire f_s_dadda_pg_rca32_and_24_6_b_6;
  wire f_s_dadda_pg_rca32_and_24_6_y0;
  wire f_s_dadda_pg_rca32_and_23_7_a_23;
  wire f_s_dadda_pg_rca32_and_23_7_b_7;
  wire f_s_dadda_pg_rca32_and_23_7_y0;
  wire f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_fa269_y4;
  wire f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_and_24_6_y0;
  wire f_s_dadda_pg_rca32_fa298_y0;
  wire f_s_dadda_pg_rca32_fa298_y1;
  wire f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_and_23_7_y0;
  wire f_s_dadda_pg_rca32_fa298_y2;
  wire f_s_dadda_pg_rca32_fa298_y3;
  wire f_s_dadda_pg_rca32_fa298_y4;
  wire f_s_dadda_pg_rca32_and_22_8_a_22;
  wire f_s_dadda_pg_rca32_and_22_8_b_8;
  wire f_s_dadda_pg_rca32_and_22_8_y0;
  wire f_s_dadda_pg_rca32_and_21_9_a_21;
  wire f_s_dadda_pg_rca32_and_21_9_b_9;
  wire f_s_dadda_pg_rca32_and_21_9_y0;
  wire f_s_dadda_pg_rca32_and_20_10_a_20;
  wire f_s_dadda_pg_rca32_and_20_10_b_10;
  wire f_s_dadda_pg_rca32_and_20_10_y0;
  wire f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_22_8_y0;
  wire f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_21_9_y0;
  wire f_s_dadda_pg_rca32_fa299_y0;
  wire f_s_dadda_pg_rca32_fa299_y1;
  wire f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_20_10_y0;
  wire f_s_dadda_pg_rca32_fa299_y2;
  wire f_s_dadda_pg_rca32_fa299_y3;
  wire f_s_dadda_pg_rca32_fa299_y4;
  wire f_s_dadda_pg_rca32_and_19_11_a_19;
  wire f_s_dadda_pg_rca32_and_19_11_b_11;
  wire f_s_dadda_pg_rca32_and_19_11_y0;
  wire f_s_dadda_pg_rca32_and_18_12_a_18;
  wire f_s_dadda_pg_rca32_and_18_12_b_12;
  wire f_s_dadda_pg_rca32_and_18_12_y0;
  wire f_s_dadda_pg_rca32_and_17_13_a_17;
  wire f_s_dadda_pg_rca32_and_17_13_b_13;
  wire f_s_dadda_pg_rca32_and_17_13_y0;
  wire f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_19_11_y0;
  wire f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_18_12_y0;
  wire f_s_dadda_pg_rca32_fa300_y0;
  wire f_s_dadda_pg_rca32_fa300_y1;
  wire f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_17_13_y0;
  wire f_s_dadda_pg_rca32_fa300_y2;
  wire f_s_dadda_pg_rca32_fa300_y3;
  wire f_s_dadda_pg_rca32_fa300_y4;
  wire f_s_dadda_pg_rca32_and_16_14_a_16;
  wire f_s_dadda_pg_rca32_and_16_14_b_14;
  wire f_s_dadda_pg_rca32_and_16_14_y0;
  wire f_s_dadda_pg_rca32_and_15_15_a_15;
  wire f_s_dadda_pg_rca32_and_15_15_b_15;
  wire f_s_dadda_pg_rca32_and_15_15_y0;
  wire f_s_dadda_pg_rca32_and_14_16_a_14;
  wire f_s_dadda_pg_rca32_and_14_16_b_16;
  wire f_s_dadda_pg_rca32_and_14_16_y0;
  wire f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_16_14_y0;
  wire f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_15_15_y0;
  wire f_s_dadda_pg_rca32_fa301_y0;
  wire f_s_dadda_pg_rca32_fa301_y1;
  wire f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_14_16_y0;
  wire f_s_dadda_pg_rca32_fa301_y2;
  wire f_s_dadda_pg_rca32_fa301_y3;
  wire f_s_dadda_pg_rca32_fa301_y4;
  wire f_s_dadda_pg_rca32_and_13_17_a_13;
  wire f_s_dadda_pg_rca32_and_13_17_b_17;
  wire f_s_dadda_pg_rca32_and_13_17_y0;
  wire f_s_dadda_pg_rca32_and_12_18_a_12;
  wire f_s_dadda_pg_rca32_and_12_18_b_18;
  wire f_s_dadda_pg_rca32_and_12_18_y0;
  wire f_s_dadda_pg_rca32_and_11_19_a_11;
  wire f_s_dadda_pg_rca32_and_11_19_b_19;
  wire f_s_dadda_pg_rca32_and_11_19_y0;
  wire f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_13_17_y0;
  wire f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_12_18_y0;
  wire f_s_dadda_pg_rca32_fa302_y0;
  wire f_s_dadda_pg_rca32_fa302_y1;
  wire f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_11_19_y0;
  wire f_s_dadda_pg_rca32_fa302_y2;
  wire f_s_dadda_pg_rca32_fa302_y3;
  wire f_s_dadda_pg_rca32_fa302_y4;
  wire f_s_dadda_pg_rca32_and_10_20_a_10;
  wire f_s_dadda_pg_rca32_and_10_20_b_20;
  wire f_s_dadda_pg_rca32_and_10_20_y0;
  wire f_s_dadda_pg_rca32_and_9_21_a_9;
  wire f_s_dadda_pg_rca32_and_9_21_b_21;
  wire f_s_dadda_pg_rca32_and_9_21_y0;
  wire f_s_dadda_pg_rca32_and_8_22_a_8;
  wire f_s_dadda_pg_rca32_and_8_22_b_22;
  wire f_s_dadda_pg_rca32_and_8_22_y0;
  wire f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_10_20_y0;
  wire f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_9_21_y0;
  wire f_s_dadda_pg_rca32_fa303_y0;
  wire f_s_dadda_pg_rca32_fa303_y1;
  wire f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_8_22_y0;
  wire f_s_dadda_pg_rca32_fa303_y2;
  wire f_s_dadda_pg_rca32_fa303_y3;
  wire f_s_dadda_pg_rca32_fa303_y4;
  wire f_s_dadda_pg_rca32_and_7_23_a_7;
  wire f_s_dadda_pg_rca32_and_7_23_b_23;
  wire f_s_dadda_pg_rca32_and_7_23_y0;
  wire f_s_dadda_pg_rca32_and_6_24_a_6;
  wire f_s_dadda_pg_rca32_and_6_24_b_24;
  wire f_s_dadda_pg_rca32_and_6_24_y0;
  wire f_s_dadda_pg_rca32_and_5_25_a_5;
  wire f_s_dadda_pg_rca32_and_5_25_b_25;
  wire f_s_dadda_pg_rca32_and_5_25_y0;
  wire f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_7_23_y0;
  wire f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_6_24_y0;
  wire f_s_dadda_pg_rca32_fa304_y0;
  wire f_s_dadda_pg_rca32_fa304_y1;
  wire f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_5_25_y0;
  wire f_s_dadda_pg_rca32_fa304_y2;
  wire f_s_dadda_pg_rca32_fa304_y3;
  wire f_s_dadda_pg_rca32_fa304_y4;
  wire f_s_dadda_pg_rca32_and_4_26_a_4;
  wire f_s_dadda_pg_rca32_and_4_26_b_26;
  wire f_s_dadda_pg_rca32_and_4_26_y0;
  wire f_s_dadda_pg_rca32_and_3_27_a_3;
  wire f_s_dadda_pg_rca32_and_3_27_b_27;
  wire f_s_dadda_pg_rca32_and_3_27_y0;
  wire f_s_dadda_pg_rca32_and_2_28_a_2;
  wire f_s_dadda_pg_rca32_and_2_28_b_28;
  wire f_s_dadda_pg_rca32_and_2_28_y0;
  wire f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_4_26_y0;
  wire f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_3_27_y0;
  wire f_s_dadda_pg_rca32_fa305_y0;
  wire f_s_dadda_pg_rca32_fa305_y1;
  wire f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_2_28_y0;
  wire f_s_dadda_pg_rca32_fa305_y2;
  wire f_s_dadda_pg_rca32_fa305_y3;
  wire f_s_dadda_pg_rca32_fa305_y4;
  wire f_s_dadda_pg_rca32_and_1_29_a_1;
  wire f_s_dadda_pg_rca32_and_1_29_b_29;
  wire f_s_dadda_pg_rca32_and_1_29_y0;
  wire f_s_dadda_pg_rca32_and_0_30_a_0;
  wire f_s_dadda_pg_rca32_and_0_30_b_30;
  wire f_s_dadda_pg_rca32_and_0_30_y0;
  wire f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_and_1_29_y0;
  wire f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_and_0_30_y0;
  wire f_s_dadda_pg_rca32_fa306_y0;
  wire f_s_dadda_pg_rca32_fa306_y1;
  wire f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_fa1_y2;
  wire f_s_dadda_pg_rca32_fa306_y2;
  wire f_s_dadda_pg_rca32_fa306_y3;
  wire f_s_dadda_pg_rca32_fa306_y4;
  wire f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_fa2_y2;
  wire f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_ha2_y0;
  wire f_s_dadda_pg_rca32_fa307_y0;
  wire f_s_dadda_pg_rca32_fa307_y1;
  wire f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_fa291_y2;
  wire f_s_dadda_pg_rca32_fa307_y2;
  wire f_s_dadda_pg_rca32_fa307_y3;
  wire f_s_dadda_pg_rca32_fa307_y4;
  wire f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa292_y2;
  wire f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa293_y2;
  wire f_s_dadda_pg_rca32_fa308_y0;
  wire f_s_dadda_pg_rca32_fa308_y1;
  wire f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa294_y2;
  wire f_s_dadda_pg_rca32_fa308_y2;
  wire f_s_dadda_pg_rca32_fa308_y3;
  wire f_s_dadda_pg_rca32_fa308_y4;
  wire f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa295_y2;
  wire f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa296_y2;
  wire f_s_dadda_pg_rca32_fa309_y0;
  wire f_s_dadda_pg_rca32_fa309_y1;
  wire f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa297_y2;
  wire f_s_dadda_pg_rca32_fa309_y2;
  wire f_s_dadda_pg_rca32_fa309_y3;
  wire f_s_dadda_pg_rca32_fa309_y4;
  wire f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa298_y2;
  wire f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa299_y2;
  wire f_s_dadda_pg_rca32_fa310_y0;
  wire f_s_dadda_pg_rca32_fa310_y1;
  wire f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa300_y2;
  wire f_s_dadda_pg_rca32_fa310_y2;
  wire f_s_dadda_pg_rca32_fa310_y3;
  wire f_s_dadda_pg_rca32_fa310_y4;
  wire f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa301_y2;
  wire f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa302_y2;
  wire f_s_dadda_pg_rca32_fa311_y0;
  wire f_s_dadda_pg_rca32_fa311_y1;
  wire f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa303_y2;
  wire f_s_dadda_pg_rca32_fa311_y2;
  wire f_s_dadda_pg_rca32_fa311_y3;
  wire f_s_dadda_pg_rca32_fa311_y4;
  wire f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa304_y2;
  wire f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa305_y2;
  wire f_s_dadda_pg_rca32_fa312_y0;
  wire f_s_dadda_pg_rca32_fa312_y1;
  wire f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa306_y2;
  wire f_s_dadda_pg_rca32_fa312_y2;
  wire f_s_dadda_pg_rca32_fa312_y3;
  wire f_s_dadda_pg_rca32_fa312_y4;
  wire f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa312_y4;
  wire f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa311_y4;
  wire f_s_dadda_pg_rca32_fa313_y0;
  wire f_s_dadda_pg_rca32_fa313_y1;
  wire f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa310_y4;
  wire f_s_dadda_pg_rca32_fa313_y2;
  wire f_s_dadda_pg_rca32_fa313_y3;
  wire f_s_dadda_pg_rca32_fa313_y4;
  wire f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa309_y4;
  wire f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa308_y4;
  wire f_s_dadda_pg_rca32_fa314_y0;
  wire f_s_dadda_pg_rca32_fa314_y1;
  wire f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa307_y4;
  wire f_s_dadda_pg_rca32_fa314_y2;
  wire f_s_dadda_pg_rca32_fa314_y3;
  wire f_s_dadda_pg_rca32_fa314_y4;
  wire f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa306_y4;
  wire f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa305_y4;
  wire f_s_dadda_pg_rca32_fa315_y0;
  wire f_s_dadda_pg_rca32_fa315_y1;
  wire f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa304_y4;
  wire f_s_dadda_pg_rca32_fa315_y2;
  wire f_s_dadda_pg_rca32_fa315_y3;
  wire f_s_dadda_pg_rca32_fa315_y4;
  wire f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa303_y4;
  wire f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa302_y4;
  wire f_s_dadda_pg_rca32_fa316_y0;
  wire f_s_dadda_pg_rca32_fa316_y1;
  wire f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa301_y4;
  wire f_s_dadda_pg_rca32_fa316_y2;
  wire f_s_dadda_pg_rca32_fa316_y3;
  wire f_s_dadda_pg_rca32_fa316_y4;
  wire f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa300_y4;
  wire f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa299_y4;
  wire f_s_dadda_pg_rca32_fa317_y0;
  wire f_s_dadda_pg_rca32_fa317_y1;
  wire f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa298_y4;
  wire f_s_dadda_pg_rca32_fa317_y2;
  wire f_s_dadda_pg_rca32_fa317_y3;
  wire f_s_dadda_pg_rca32_fa317_y4;
  wire f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa297_y4;
  wire f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa296_y4;
  wire f_s_dadda_pg_rca32_fa318_y0;
  wire f_s_dadda_pg_rca32_fa318_y1;
  wire f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa295_y4;
  wire f_s_dadda_pg_rca32_fa318_y2;
  wire f_s_dadda_pg_rca32_fa318_y3;
  wire f_s_dadda_pg_rca32_fa318_y4;
  wire f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa294_y4;
  wire f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa293_y4;
  wire f_s_dadda_pg_rca32_fa319_y0;
  wire f_s_dadda_pg_rca32_fa319_y1;
  wire f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa292_y4;
  wire f_s_dadda_pg_rca32_fa319_y2;
  wire f_s_dadda_pg_rca32_fa319_y3;
  wire f_s_dadda_pg_rca32_fa319_y4;
  wire f_s_dadda_pg_rca32_and_23_8_a_23;
  wire f_s_dadda_pg_rca32_and_23_8_b_8;
  wire f_s_dadda_pg_rca32_and_23_8_y0;
  wire f_s_dadda_pg_rca32_and_22_9_a_22;
  wire f_s_dadda_pg_rca32_and_22_9_b_9;
  wire f_s_dadda_pg_rca32_and_22_9_y0;
  wire f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_fa291_y4;
  wire f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_and_23_8_y0;
  wire f_s_dadda_pg_rca32_fa320_y0;
  wire f_s_dadda_pg_rca32_fa320_y1;
  wire f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_and_22_9_y0;
  wire f_s_dadda_pg_rca32_fa320_y2;
  wire f_s_dadda_pg_rca32_fa320_y3;
  wire f_s_dadda_pg_rca32_fa320_y4;
  wire f_s_dadda_pg_rca32_and_21_10_a_21;
  wire f_s_dadda_pg_rca32_and_21_10_b_10;
  wire f_s_dadda_pg_rca32_and_21_10_y0;
  wire f_s_dadda_pg_rca32_and_20_11_a_20;
  wire f_s_dadda_pg_rca32_and_20_11_b_11;
  wire f_s_dadda_pg_rca32_and_20_11_y0;
  wire f_s_dadda_pg_rca32_and_19_12_a_19;
  wire f_s_dadda_pg_rca32_and_19_12_b_12;
  wire f_s_dadda_pg_rca32_and_19_12_y0;
  wire f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_21_10_y0;
  wire f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_20_11_y0;
  wire f_s_dadda_pg_rca32_fa321_y0;
  wire f_s_dadda_pg_rca32_fa321_y1;
  wire f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_19_12_y0;
  wire f_s_dadda_pg_rca32_fa321_y2;
  wire f_s_dadda_pg_rca32_fa321_y3;
  wire f_s_dadda_pg_rca32_fa321_y4;
  wire f_s_dadda_pg_rca32_and_18_13_a_18;
  wire f_s_dadda_pg_rca32_and_18_13_b_13;
  wire f_s_dadda_pg_rca32_and_18_13_y0;
  wire f_s_dadda_pg_rca32_and_17_14_a_17;
  wire f_s_dadda_pg_rca32_and_17_14_b_14;
  wire f_s_dadda_pg_rca32_and_17_14_y0;
  wire f_s_dadda_pg_rca32_and_16_15_a_16;
  wire f_s_dadda_pg_rca32_and_16_15_b_15;
  wire f_s_dadda_pg_rca32_and_16_15_y0;
  wire f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_18_13_y0;
  wire f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_17_14_y0;
  wire f_s_dadda_pg_rca32_fa322_y0;
  wire f_s_dadda_pg_rca32_fa322_y1;
  wire f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_16_15_y0;
  wire f_s_dadda_pg_rca32_fa322_y2;
  wire f_s_dadda_pg_rca32_fa322_y3;
  wire f_s_dadda_pg_rca32_fa322_y4;
  wire f_s_dadda_pg_rca32_and_15_16_a_15;
  wire f_s_dadda_pg_rca32_and_15_16_b_16;
  wire f_s_dadda_pg_rca32_and_15_16_y0;
  wire f_s_dadda_pg_rca32_and_14_17_a_14;
  wire f_s_dadda_pg_rca32_and_14_17_b_17;
  wire f_s_dadda_pg_rca32_and_14_17_y0;
  wire f_s_dadda_pg_rca32_and_13_18_a_13;
  wire f_s_dadda_pg_rca32_and_13_18_b_18;
  wire f_s_dadda_pg_rca32_and_13_18_y0;
  wire f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_15_16_y0;
  wire f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_14_17_y0;
  wire f_s_dadda_pg_rca32_fa323_y0;
  wire f_s_dadda_pg_rca32_fa323_y1;
  wire f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_13_18_y0;
  wire f_s_dadda_pg_rca32_fa323_y2;
  wire f_s_dadda_pg_rca32_fa323_y3;
  wire f_s_dadda_pg_rca32_fa323_y4;
  wire f_s_dadda_pg_rca32_and_12_19_a_12;
  wire f_s_dadda_pg_rca32_and_12_19_b_19;
  wire f_s_dadda_pg_rca32_and_12_19_y0;
  wire f_s_dadda_pg_rca32_and_11_20_a_11;
  wire f_s_dadda_pg_rca32_and_11_20_b_20;
  wire f_s_dadda_pg_rca32_and_11_20_y0;
  wire f_s_dadda_pg_rca32_and_10_21_a_10;
  wire f_s_dadda_pg_rca32_and_10_21_b_21;
  wire f_s_dadda_pg_rca32_and_10_21_y0;
  wire f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_12_19_y0;
  wire f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_11_20_y0;
  wire f_s_dadda_pg_rca32_fa324_y0;
  wire f_s_dadda_pg_rca32_fa324_y1;
  wire f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_10_21_y0;
  wire f_s_dadda_pg_rca32_fa324_y2;
  wire f_s_dadda_pg_rca32_fa324_y3;
  wire f_s_dadda_pg_rca32_fa324_y4;
  wire f_s_dadda_pg_rca32_and_9_22_a_9;
  wire f_s_dadda_pg_rca32_and_9_22_b_22;
  wire f_s_dadda_pg_rca32_and_9_22_y0;
  wire f_s_dadda_pg_rca32_and_8_23_a_8;
  wire f_s_dadda_pg_rca32_and_8_23_b_23;
  wire f_s_dadda_pg_rca32_and_8_23_y0;
  wire f_s_dadda_pg_rca32_and_7_24_a_7;
  wire f_s_dadda_pg_rca32_and_7_24_b_24;
  wire f_s_dadda_pg_rca32_and_7_24_y0;
  wire f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_9_22_y0;
  wire f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_8_23_y0;
  wire f_s_dadda_pg_rca32_fa325_y0;
  wire f_s_dadda_pg_rca32_fa325_y1;
  wire f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_7_24_y0;
  wire f_s_dadda_pg_rca32_fa325_y2;
  wire f_s_dadda_pg_rca32_fa325_y3;
  wire f_s_dadda_pg_rca32_fa325_y4;
  wire f_s_dadda_pg_rca32_and_6_25_a_6;
  wire f_s_dadda_pg_rca32_and_6_25_b_25;
  wire f_s_dadda_pg_rca32_and_6_25_y0;
  wire f_s_dadda_pg_rca32_and_5_26_a_5;
  wire f_s_dadda_pg_rca32_and_5_26_b_26;
  wire f_s_dadda_pg_rca32_and_5_26_y0;
  wire f_s_dadda_pg_rca32_and_4_27_a_4;
  wire f_s_dadda_pg_rca32_and_4_27_b_27;
  wire f_s_dadda_pg_rca32_and_4_27_y0;
  wire f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_6_25_y0;
  wire f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_5_26_y0;
  wire f_s_dadda_pg_rca32_fa326_y0;
  wire f_s_dadda_pg_rca32_fa326_y1;
  wire f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_4_27_y0;
  wire f_s_dadda_pg_rca32_fa326_y2;
  wire f_s_dadda_pg_rca32_fa326_y3;
  wire f_s_dadda_pg_rca32_fa326_y4;
  wire f_s_dadda_pg_rca32_and_3_28_a_3;
  wire f_s_dadda_pg_rca32_and_3_28_b_28;
  wire f_s_dadda_pg_rca32_and_3_28_y0;
  wire f_s_dadda_pg_rca32_and_2_29_a_2;
  wire f_s_dadda_pg_rca32_and_2_29_b_29;
  wire f_s_dadda_pg_rca32_and_2_29_y0;
  wire f_s_dadda_pg_rca32_and_1_30_a_1;
  wire f_s_dadda_pg_rca32_and_1_30_b_30;
  wire f_s_dadda_pg_rca32_and_1_30_y0;
  wire f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_3_28_y0;
  wire f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_2_29_y0;
  wire f_s_dadda_pg_rca32_fa327_y0;
  wire f_s_dadda_pg_rca32_fa327_y1;
  wire f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_1_30_y0;
  wire f_s_dadda_pg_rca32_fa327_y2;
  wire f_s_dadda_pg_rca32_fa327_y3;
  wire f_s_dadda_pg_rca32_fa327_y4;
  wire f_s_dadda_pg_rca32_nand_0_31_a_0;
  wire f_s_dadda_pg_rca32_nand_0_31_b_31;
  wire f_s_dadda_pg_rca32_nand_0_31_y0;
  wire f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_nand_0_31_y0;
  wire f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_fa3_y2;
  wire f_s_dadda_pg_rca32_fa328_y0;
  wire f_s_dadda_pg_rca32_fa328_y1;
  wire f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_fa4_y2;
  wire f_s_dadda_pg_rca32_fa328_y2;
  wire f_s_dadda_pg_rca32_fa328_y3;
  wire f_s_dadda_pg_rca32_fa328_y4;
  wire f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_fa5_y2;
  wire f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_ha3_y0;
  wire f_s_dadda_pg_rca32_fa329_y0;
  wire f_s_dadda_pg_rca32_fa329_y1;
  wire f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_fa313_y2;
  wire f_s_dadda_pg_rca32_fa329_y2;
  wire f_s_dadda_pg_rca32_fa329_y3;
  wire f_s_dadda_pg_rca32_fa329_y4;
  wire f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa314_y2;
  wire f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa315_y2;
  wire f_s_dadda_pg_rca32_fa330_y0;
  wire f_s_dadda_pg_rca32_fa330_y1;
  wire f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa316_y2;
  wire f_s_dadda_pg_rca32_fa330_y2;
  wire f_s_dadda_pg_rca32_fa330_y3;
  wire f_s_dadda_pg_rca32_fa330_y4;
  wire f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa317_y2;
  wire f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa318_y2;
  wire f_s_dadda_pg_rca32_fa331_y0;
  wire f_s_dadda_pg_rca32_fa331_y1;
  wire f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa319_y2;
  wire f_s_dadda_pg_rca32_fa331_y2;
  wire f_s_dadda_pg_rca32_fa331_y3;
  wire f_s_dadda_pg_rca32_fa331_y4;
  wire f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa320_y2;
  wire f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa321_y2;
  wire f_s_dadda_pg_rca32_fa332_y0;
  wire f_s_dadda_pg_rca32_fa332_y1;
  wire f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa322_y2;
  wire f_s_dadda_pg_rca32_fa332_y2;
  wire f_s_dadda_pg_rca32_fa332_y3;
  wire f_s_dadda_pg_rca32_fa332_y4;
  wire f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa323_y2;
  wire f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa324_y2;
  wire f_s_dadda_pg_rca32_fa333_y0;
  wire f_s_dadda_pg_rca32_fa333_y1;
  wire f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa325_y2;
  wire f_s_dadda_pg_rca32_fa333_y2;
  wire f_s_dadda_pg_rca32_fa333_y3;
  wire f_s_dadda_pg_rca32_fa333_y4;
  wire f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa326_y2;
  wire f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa327_y2;
  wire f_s_dadda_pg_rca32_fa334_y0;
  wire f_s_dadda_pg_rca32_fa334_y1;
  wire f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa328_y2;
  wire f_s_dadda_pg_rca32_fa334_y2;
  wire f_s_dadda_pg_rca32_fa334_y3;
  wire f_s_dadda_pg_rca32_fa334_y4;
  wire f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa334_y4;
  wire f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa333_y4;
  wire f_s_dadda_pg_rca32_fa335_y0;
  wire f_s_dadda_pg_rca32_fa335_y1;
  wire f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa332_y4;
  wire f_s_dadda_pg_rca32_fa335_y2;
  wire f_s_dadda_pg_rca32_fa335_y3;
  wire f_s_dadda_pg_rca32_fa335_y4;
  wire f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa331_y4;
  wire f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa330_y4;
  wire f_s_dadda_pg_rca32_fa336_y0;
  wire f_s_dadda_pg_rca32_fa336_y1;
  wire f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa329_y4;
  wire f_s_dadda_pg_rca32_fa336_y2;
  wire f_s_dadda_pg_rca32_fa336_y3;
  wire f_s_dadda_pg_rca32_fa336_y4;
  wire f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa328_y4;
  wire f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa327_y4;
  wire f_s_dadda_pg_rca32_fa337_y0;
  wire f_s_dadda_pg_rca32_fa337_y1;
  wire f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa326_y4;
  wire f_s_dadda_pg_rca32_fa337_y2;
  wire f_s_dadda_pg_rca32_fa337_y3;
  wire f_s_dadda_pg_rca32_fa337_y4;
  wire f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa325_y4;
  wire f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa324_y4;
  wire f_s_dadda_pg_rca32_fa338_y0;
  wire f_s_dadda_pg_rca32_fa338_y1;
  wire f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa323_y4;
  wire f_s_dadda_pg_rca32_fa338_y2;
  wire f_s_dadda_pg_rca32_fa338_y3;
  wire f_s_dadda_pg_rca32_fa338_y4;
  wire f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa322_y4;
  wire f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa321_y4;
  wire f_s_dadda_pg_rca32_fa339_y0;
  wire f_s_dadda_pg_rca32_fa339_y1;
  wire f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa320_y4;
  wire f_s_dadda_pg_rca32_fa339_y2;
  wire f_s_dadda_pg_rca32_fa339_y3;
  wire f_s_dadda_pg_rca32_fa339_y4;
  wire f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa319_y4;
  wire f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa318_y4;
  wire f_s_dadda_pg_rca32_fa340_y0;
  wire f_s_dadda_pg_rca32_fa340_y1;
  wire f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa317_y4;
  wire f_s_dadda_pg_rca32_fa340_y2;
  wire f_s_dadda_pg_rca32_fa340_y3;
  wire f_s_dadda_pg_rca32_fa340_y4;
  wire f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa316_y4;
  wire f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa315_y4;
  wire f_s_dadda_pg_rca32_fa341_y0;
  wire f_s_dadda_pg_rca32_fa341_y1;
  wire f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa314_y4;
  wire f_s_dadda_pg_rca32_fa341_y2;
  wire f_s_dadda_pg_rca32_fa341_y3;
  wire f_s_dadda_pg_rca32_fa341_y4;
  wire f_s_dadda_pg_rca32_and_24_8_a_24;
  wire f_s_dadda_pg_rca32_and_24_8_b_8;
  wire f_s_dadda_pg_rca32_and_24_8_y0;
  wire f_s_dadda_pg_rca32_and_23_9_a_23;
  wire f_s_dadda_pg_rca32_and_23_9_b_9;
  wire f_s_dadda_pg_rca32_and_23_9_y0;
  wire f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_fa313_y4;
  wire f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_and_24_8_y0;
  wire f_s_dadda_pg_rca32_fa342_y0;
  wire f_s_dadda_pg_rca32_fa342_y1;
  wire f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_and_23_9_y0;
  wire f_s_dadda_pg_rca32_fa342_y2;
  wire f_s_dadda_pg_rca32_fa342_y3;
  wire f_s_dadda_pg_rca32_fa342_y4;
  wire f_s_dadda_pg_rca32_and_22_10_a_22;
  wire f_s_dadda_pg_rca32_and_22_10_b_10;
  wire f_s_dadda_pg_rca32_and_22_10_y0;
  wire f_s_dadda_pg_rca32_and_21_11_a_21;
  wire f_s_dadda_pg_rca32_and_21_11_b_11;
  wire f_s_dadda_pg_rca32_and_21_11_y0;
  wire f_s_dadda_pg_rca32_and_20_12_a_20;
  wire f_s_dadda_pg_rca32_and_20_12_b_12;
  wire f_s_dadda_pg_rca32_and_20_12_y0;
  wire f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_22_10_y0;
  wire f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_21_11_y0;
  wire f_s_dadda_pg_rca32_fa343_y0;
  wire f_s_dadda_pg_rca32_fa343_y1;
  wire f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_20_12_y0;
  wire f_s_dadda_pg_rca32_fa343_y2;
  wire f_s_dadda_pg_rca32_fa343_y3;
  wire f_s_dadda_pg_rca32_fa343_y4;
  wire f_s_dadda_pg_rca32_and_19_13_a_19;
  wire f_s_dadda_pg_rca32_and_19_13_b_13;
  wire f_s_dadda_pg_rca32_and_19_13_y0;
  wire f_s_dadda_pg_rca32_and_18_14_a_18;
  wire f_s_dadda_pg_rca32_and_18_14_b_14;
  wire f_s_dadda_pg_rca32_and_18_14_y0;
  wire f_s_dadda_pg_rca32_and_17_15_a_17;
  wire f_s_dadda_pg_rca32_and_17_15_b_15;
  wire f_s_dadda_pg_rca32_and_17_15_y0;
  wire f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_19_13_y0;
  wire f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_18_14_y0;
  wire f_s_dadda_pg_rca32_fa344_y0;
  wire f_s_dadda_pg_rca32_fa344_y1;
  wire f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_17_15_y0;
  wire f_s_dadda_pg_rca32_fa344_y2;
  wire f_s_dadda_pg_rca32_fa344_y3;
  wire f_s_dadda_pg_rca32_fa344_y4;
  wire f_s_dadda_pg_rca32_and_16_16_a_16;
  wire f_s_dadda_pg_rca32_and_16_16_b_16;
  wire f_s_dadda_pg_rca32_and_16_16_y0;
  wire f_s_dadda_pg_rca32_and_15_17_a_15;
  wire f_s_dadda_pg_rca32_and_15_17_b_17;
  wire f_s_dadda_pg_rca32_and_15_17_y0;
  wire f_s_dadda_pg_rca32_and_14_18_a_14;
  wire f_s_dadda_pg_rca32_and_14_18_b_18;
  wire f_s_dadda_pg_rca32_and_14_18_y0;
  wire f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_16_16_y0;
  wire f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_15_17_y0;
  wire f_s_dadda_pg_rca32_fa345_y0;
  wire f_s_dadda_pg_rca32_fa345_y1;
  wire f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_14_18_y0;
  wire f_s_dadda_pg_rca32_fa345_y2;
  wire f_s_dadda_pg_rca32_fa345_y3;
  wire f_s_dadda_pg_rca32_fa345_y4;
  wire f_s_dadda_pg_rca32_and_13_19_a_13;
  wire f_s_dadda_pg_rca32_and_13_19_b_19;
  wire f_s_dadda_pg_rca32_and_13_19_y0;
  wire f_s_dadda_pg_rca32_and_12_20_a_12;
  wire f_s_dadda_pg_rca32_and_12_20_b_20;
  wire f_s_dadda_pg_rca32_and_12_20_y0;
  wire f_s_dadda_pg_rca32_and_11_21_a_11;
  wire f_s_dadda_pg_rca32_and_11_21_b_21;
  wire f_s_dadda_pg_rca32_and_11_21_y0;
  wire f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_13_19_y0;
  wire f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_12_20_y0;
  wire f_s_dadda_pg_rca32_fa346_y0;
  wire f_s_dadda_pg_rca32_fa346_y1;
  wire f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_11_21_y0;
  wire f_s_dadda_pg_rca32_fa346_y2;
  wire f_s_dadda_pg_rca32_fa346_y3;
  wire f_s_dadda_pg_rca32_fa346_y4;
  wire f_s_dadda_pg_rca32_and_10_22_a_10;
  wire f_s_dadda_pg_rca32_and_10_22_b_22;
  wire f_s_dadda_pg_rca32_and_10_22_y0;
  wire f_s_dadda_pg_rca32_and_9_23_a_9;
  wire f_s_dadda_pg_rca32_and_9_23_b_23;
  wire f_s_dadda_pg_rca32_and_9_23_y0;
  wire f_s_dadda_pg_rca32_and_8_24_a_8;
  wire f_s_dadda_pg_rca32_and_8_24_b_24;
  wire f_s_dadda_pg_rca32_and_8_24_y0;
  wire f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_10_22_y0;
  wire f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_9_23_y0;
  wire f_s_dadda_pg_rca32_fa347_y0;
  wire f_s_dadda_pg_rca32_fa347_y1;
  wire f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_8_24_y0;
  wire f_s_dadda_pg_rca32_fa347_y2;
  wire f_s_dadda_pg_rca32_fa347_y3;
  wire f_s_dadda_pg_rca32_fa347_y4;
  wire f_s_dadda_pg_rca32_and_7_25_a_7;
  wire f_s_dadda_pg_rca32_and_7_25_b_25;
  wire f_s_dadda_pg_rca32_and_7_25_y0;
  wire f_s_dadda_pg_rca32_and_6_26_a_6;
  wire f_s_dadda_pg_rca32_and_6_26_b_26;
  wire f_s_dadda_pg_rca32_and_6_26_y0;
  wire f_s_dadda_pg_rca32_and_5_27_a_5;
  wire f_s_dadda_pg_rca32_and_5_27_b_27;
  wire f_s_dadda_pg_rca32_and_5_27_y0;
  wire f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_7_25_y0;
  wire f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_6_26_y0;
  wire f_s_dadda_pg_rca32_fa348_y0;
  wire f_s_dadda_pg_rca32_fa348_y1;
  wire f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_5_27_y0;
  wire f_s_dadda_pg_rca32_fa348_y2;
  wire f_s_dadda_pg_rca32_fa348_y3;
  wire f_s_dadda_pg_rca32_fa348_y4;
  wire f_s_dadda_pg_rca32_and_4_28_a_4;
  wire f_s_dadda_pg_rca32_and_4_28_b_28;
  wire f_s_dadda_pg_rca32_and_4_28_y0;
  wire f_s_dadda_pg_rca32_and_3_29_a_3;
  wire f_s_dadda_pg_rca32_and_3_29_b_29;
  wire f_s_dadda_pg_rca32_and_3_29_y0;
  wire f_s_dadda_pg_rca32_and_2_30_a_2;
  wire f_s_dadda_pg_rca32_and_2_30_b_30;
  wire f_s_dadda_pg_rca32_and_2_30_y0;
  wire f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_4_28_y0;
  wire f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_3_29_y0;
  wire f_s_dadda_pg_rca32_fa349_y0;
  wire f_s_dadda_pg_rca32_fa349_y1;
  wire f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_2_30_y0;
  wire f_s_dadda_pg_rca32_fa349_y2;
  wire f_s_dadda_pg_rca32_fa349_y3;
  wire f_s_dadda_pg_rca32_fa349_y4;
  wire f_s_dadda_pg_rca32_nand_1_31_a_1;
  wire f_s_dadda_pg_rca32_nand_1_31_b_31;
  wire f_s_dadda_pg_rca32_nand_1_31_y0;
  wire f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_nand_1_31_y0;
  wire f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_fa6_y2;
  wire f_s_dadda_pg_rca32_fa350_y0;
  wire f_s_dadda_pg_rca32_fa350_y1;
  wire f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_fa7_y2;
  wire f_s_dadda_pg_rca32_fa350_y2;
  wire f_s_dadda_pg_rca32_fa350_y3;
  wire f_s_dadda_pg_rca32_fa350_y4;
  wire f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa8_y2;
  wire f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa9_y2;
  wire f_s_dadda_pg_rca32_fa351_y0;
  wire f_s_dadda_pg_rca32_fa351_y1;
  wire f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa335_y2;
  wire f_s_dadda_pg_rca32_fa351_y2;
  wire f_s_dadda_pg_rca32_fa351_y3;
  wire f_s_dadda_pg_rca32_fa351_y4;
  wire f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa336_y2;
  wire f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa337_y2;
  wire f_s_dadda_pg_rca32_fa352_y0;
  wire f_s_dadda_pg_rca32_fa352_y1;
  wire f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa338_y2;
  wire f_s_dadda_pg_rca32_fa352_y2;
  wire f_s_dadda_pg_rca32_fa352_y3;
  wire f_s_dadda_pg_rca32_fa352_y4;
  wire f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa339_y2;
  wire f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa340_y2;
  wire f_s_dadda_pg_rca32_fa353_y0;
  wire f_s_dadda_pg_rca32_fa353_y1;
  wire f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa341_y2;
  wire f_s_dadda_pg_rca32_fa353_y2;
  wire f_s_dadda_pg_rca32_fa353_y3;
  wire f_s_dadda_pg_rca32_fa353_y4;
  wire f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa342_y2;
  wire f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa343_y2;
  wire f_s_dadda_pg_rca32_fa354_y0;
  wire f_s_dadda_pg_rca32_fa354_y1;
  wire f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa344_y2;
  wire f_s_dadda_pg_rca32_fa354_y2;
  wire f_s_dadda_pg_rca32_fa354_y3;
  wire f_s_dadda_pg_rca32_fa354_y4;
  wire f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa345_y2;
  wire f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa346_y2;
  wire f_s_dadda_pg_rca32_fa355_y0;
  wire f_s_dadda_pg_rca32_fa355_y1;
  wire f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa347_y2;
  wire f_s_dadda_pg_rca32_fa355_y2;
  wire f_s_dadda_pg_rca32_fa355_y3;
  wire f_s_dadda_pg_rca32_fa355_y4;
  wire f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa348_y2;
  wire f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa349_y2;
  wire f_s_dadda_pg_rca32_fa356_y0;
  wire f_s_dadda_pg_rca32_fa356_y1;
  wire f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa350_y2;
  wire f_s_dadda_pg_rca32_fa356_y2;
  wire f_s_dadda_pg_rca32_fa356_y3;
  wire f_s_dadda_pg_rca32_fa356_y4;
  wire f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa356_y4;
  wire f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa355_y4;
  wire f_s_dadda_pg_rca32_fa357_y0;
  wire f_s_dadda_pg_rca32_fa357_y1;
  wire f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa354_y4;
  wire f_s_dadda_pg_rca32_fa357_y2;
  wire f_s_dadda_pg_rca32_fa357_y3;
  wire f_s_dadda_pg_rca32_fa357_y4;
  wire f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa353_y4;
  wire f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa352_y4;
  wire f_s_dadda_pg_rca32_fa358_y0;
  wire f_s_dadda_pg_rca32_fa358_y1;
  wire f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa351_y4;
  wire f_s_dadda_pg_rca32_fa358_y2;
  wire f_s_dadda_pg_rca32_fa358_y3;
  wire f_s_dadda_pg_rca32_fa358_y4;
  wire f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa350_y4;
  wire f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa349_y4;
  wire f_s_dadda_pg_rca32_fa359_y0;
  wire f_s_dadda_pg_rca32_fa359_y1;
  wire f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa348_y4;
  wire f_s_dadda_pg_rca32_fa359_y2;
  wire f_s_dadda_pg_rca32_fa359_y3;
  wire f_s_dadda_pg_rca32_fa359_y4;
  wire f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa347_y4;
  wire f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa346_y4;
  wire f_s_dadda_pg_rca32_fa360_y0;
  wire f_s_dadda_pg_rca32_fa360_y1;
  wire f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa345_y4;
  wire f_s_dadda_pg_rca32_fa360_y2;
  wire f_s_dadda_pg_rca32_fa360_y3;
  wire f_s_dadda_pg_rca32_fa360_y4;
  wire f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa344_y4;
  wire f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa343_y4;
  wire f_s_dadda_pg_rca32_fa361_y0;
  wire f_s_dadda_pg_rca32_fa361_y1;
  wire f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa342_y4;
  wire f_s_dadda_pg_rca32_fa361_y2;
  wire f_s_dadda_pg_rca32_fa361_y3;
  wire f_s_dadda_pg_rca32_fa361_y4;
  wire f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa341_y4;
  wire f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa340_y4;
  wire f_s_dadda_pg_rca32_fa362_y0;
  wire f_s_dadda_pg_rca32_fa362_y1;
  wire f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa339_y4;
  wire f_s_dadda_pg_rca32_fa362_y2;
  wire f_s_dadda_pg_rca32_fa362_y3;
  wire f_s_dadda_pg_rca32_fa362_y4;
  wire f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa338_y4;
  wire f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa337_y4;
  wire f_s_dadda_pg_rca32_fa363_y0;
  wire f_s_dadda_pg_rca32_fa363_y1;
  wire f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa336_y4;
  wire f_s_dadda_pg_rca32_fa363_y2;
  wire f_s_dadda_pg_rca32_fa363_y3;
  wire f_s_dadda_pg_rca32_fa363_y4;
  wire f_s_dadda_pg_rca32_and_26_7_a_26;
  wire f_s_dadda_pg_rca32_and_26_7_b_7;
  wire f_s_dadda_pg_rca32_and_26_7_y0;
  wire f_s_dadda_pg_rca32_and_25_8_a_25;
  wire f_s_dadda_pg_rca32_and_25_8_b_8;
  wire f_s_dadda_pg_rca32_and_25_8_y0;
  wire f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_fa335_y4;
  wire f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_and_26_7_y0;
  wire f_s_dadda_pg_rca32_fa364_y0;
  wire f_s_dadda_pg_rca32_fa364_y1;
  wire f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_and_25_8_y0;
  wire f_s_dadda_pg_rca32_fa364_y2;
  wire f_s_dadda_pg_rca32_fa364_y3;
  wire f_s_dadda_pg_rca32_fa364_y4;
  wire f_s_dadda_pg_rca32_and_24_9_a_24;
  wire f_s_dadda_pg_rca32_and_24_9_b_9;
  wire f_s_dadda_pg_rca32_and_24_9_y0;
  wire f_s_dadda_pg_rca32_and_23_10_a_23;
  wire f_s_dadda_pg_rca32_and_23_10_b_10;
  wire f_s_dadda_pg_rca32_and_23_10_y0;
  wire f_s_dadda_pg_rca32_and_22_11_a_22;
  wire f_s_dadda_pg_rca32_and_22_11_b_11;
  wire f_s_dadda_pg_rca32_and_22_11_y0;
  wire f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_24_9_y0;
  wire f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_23_10_y0;
  wire f_s_dadda_pg_rca32_fa365_y0;
  wire f_s_dadda_pg_rca32_fa365_y1;
  wire f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_22_11_y0;
  wire f_s_dadda_pg_rca32_fa365_y2;
  wire f_s_dadda_pg_rca32_fa365_y3;
  wire f_s_dadda_pg_rca32_fa365_y4;
  wire f_s_dadda_pg_rca32_and_21_12_a_21;
  wire f_s_dadda_pg_rca32_and_21_12_b_12;
  wire f_s_dadda_pg_rca32_and_21_12_y0;
  wire f_s_dadda_pg_rca32_and_20_13_a_20;
  wire f_s_dadda_pg_rca32_and_20_13_b_13;
  wire f_s_dadda_pg_rca32_and_20_13_y0;
  wire f_s_dadda_pg_rca32_and_19_14_a_19;
  wire f_s_dadda_pg_rca32_and_19_14_b_14;
  wire f_s_dadda_pg_rca32_and_19_14_y0;
  wire f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_21_12_y0;
  wire f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_20_13_y0;
  wire f_s_dadda_pg_rca32_fa366_y0;
  wire f_s_dadda_pg_rca32_fa366_y1;
  wire f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_19_14_y0;
  wire f_s_dadda_pg_rca32_fa366_y2;
  wire f_s_dadda_pg_rca32_fa366_y3;
  wire f_s_dadda_pg_rca32_fa366_y4;
  wire f_s_dadda_pg_rca32_and_18_15_a_18;
  wire f_s_dadda_pg_rca32_and_18_15_b_15;
  wire f_s_dadda_pg_rca32_and_18_15_y0;
  wire f_s_dadda_pg_rca32_and_17_16_a_17;
  wire f_s_dadda_pg_rca32_and_17_16_b_16;
  wire f_s_dadda_pg_rca32_and_17_16_y0;
  wire f_s_dadda_pg_rca32_and_16_17_a_16;
  wire f_s_dadda_pg_rca32_and_16_17_b_17;
  wire f_s_dadda_pg_rca32_and_16_17_y0;
  wire f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_18_15_y0;
  wire f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_17_16_y0;
  wire f_s_dadda_pg_rca32_fa367_y0;
  wire f_s_dadda_pg_rca32_fa367_y1;
  wire f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_16_17_y0;
  wire f_s_dadda_pg_rca32_fa367_y2;
  wire f_s_dadda_pg_rca32_fa367_y3;
  wire f_s_dadda_pg_rca32_fa367_y4;
  wire f_s_dadda_pg_rca32_and_15_18_a_15;
  wire f_s_dadda_pg_rca32_and_15_18_b_18;
  wire f_s_dadda_pg_rca32_and_15_18_y0;
  wire f_s_dadda_pg_rca32_and_14_19_a_14;
  wire f_s_dadda_pg_rca32_and_14_19_b_19;
  wire f_s_dadda_pg_rca32_and_14_19_y0;
  wire f_s_dadda_pg_rca32_and_13_20_a_13;
  wire f_s_dadda_pg_rca32_and_13_20_b_20;
  wire f_s_dadda_pg_rca32_and_13_20_y0;
  wire f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_15_18_y0;
  wire f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_14_19_y0;
  wire f_s_dadda_pg_rca32_fa368_y0;
  wire f_s_dadda_pg_rca32_fa368_y1;
  wire f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_13_20_y0;
  wire f_s_dadda_pg_rca32_fa368_y2;
  wire f_s_dadda_pg_rca32_fa368_y3;
  wire f_s_dadda_pg_rca32_fa368_y4;
  wire f_s_dadda_pg_rca32_and_12_21_a_12;
  wire f_s_dadda_pg_rca32_and_12_21_b_21;
  wire f_s_dadda_pg_rca32_and_12_21_y0;
  wire f_s_dadda_pg_rca32_and_11_22_a_11;
  wire f_s_dadda_pg_rca32_and_11_22_b_22;
  wire f_s_dadda_pg_rca32_and_11_22_y0;
  wire f_s_dadda_pg_rca32_and_10_23_a_10;
  wire f_s_dadda_pg_rca32_and_10_23_b_23;
  wire f_s_dadda_pg_rca32_and_10_23_y0;
  wire f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_12_21_y0;
  wire f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_11_22_y0;
  wire f_s_dadda_pg_rca32_fa369_y0;
  wire f_s_dadda_pg_rca32_fa369_y1;
  wire f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_10_23_y0;
  wire f_s_dadda_pg_rca32_fa369_y2;
  wire f_s_dadda_pg_rca32_fa369_y3;
  wire f_s_dadda_pg_rca32_fa369_y4;
  wire f_s_dadda_pg_rca32_and_9_24_a_9;
  wire f_s_dadda_pg_rca32_and_9_24_b_24;
  wire f_s_dadda_pg_rca32_and_9_24_y0;
  wire f_s_dadda_pg_rca32_and_8_25_a_8;
  wire f_s_dadda_pg_rca32_and_8_25_b_25;
  wire f_s_dadda_pg_rca32_and_8_25_y0;
  wire f_s_dadda_pg_rca32_and_7_26_a_7;
  wire f_s_dadda_pg_rca32_and_7_26_b_26;
  wire f_s_dadda_pg_rca32_and_7_26_y0;
  wire f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_9_24_y0;
  wire f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_8_25_y0;
  wire f_s_dadda_pg_rca32_fa370_y0;
  wire f_s_dadda_pg_rca32_fa370_y1;
  wire f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_7_26_y0;
  wire f_s_dadda_pg_rca32_fa370_y2;
  wire f_s_dadda_pg_rca32_fa370_y3;
  wire f_s_dadda_pg_rca32_fa370_y4;
  wire f_s_dadda_pg_rca32_and_6_27_a_6;
  wire f_s_dadda_pg_rca32_and_6_27_b_27;
  wire f_s_dadda_pg_rca32_and_6_27_y0;
  wire f_s_dadda_pg_rca32_and_5_28_a_5;
  wire f_s_dadda_pg_rca32_and_5_28_b_28;
  wire f_s_dadda_pg_rca32_and_5_28_y0;
  wire f_s_dadda_pg_rca32_and_4_29_a_4;
  wire f_s_dadda_pg_rca32_and_4_29_b_29;
  wire f_s_dadda_pg_rca32_and_4_29_y0;
  wire f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_6_27_y0;
  wire f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_5_28_y0;
  wire f_s_dadda_pg_rca32_fa371_y0;
  wire f_s_dadda_pg_rca32_fa371_y1;
  wire f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_4_29_y0;
  wire f_s_dadda_pg_rca32_fa371_y2;
  wire f_s_dadda_pg_rca32_fa371_y3;
  wire f_s_dadda_pg_rca32_fa371_y4;
  wire f_s_dadda_pg_rca32_and_3_30_a_3;
  wire f_s_dadda_pg_rca32_and_3_30_b_30;
  wire f_s_dadda_pg_rca32_and_3_30_y0;
  wire f_s_dadda_pg_rca32_nand_2_31_a_2;
  wire f_s_dadda_pg_rca32_nand_2_31_b_31;
  wire f_s_dadda_pg_rca32_nand_2_31_y0;
  wire f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_and_3_30_y0;
  wire f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_nand_2_31_y0;
  wire f_s_dadda_pg_rca32_fa372_y0;
  wire f_s_dadda_pg_rca32_fa372_y1;
  wire f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_fa10_y2;
  wire f_s_dadda_pg_rca32_fa372_y2;
  wire f_s_dadda_pg_rca32_fa372_y3;
  wire f_s_dadda_pg_rca32_fa372_y4;
  wire f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa11_y2;
  wire f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa12_y2;
  wire f_s_dadda_pg_rca32_fa373_y0;
  wire f_s_dadda_pg_rca32_fa373_y1;
  wire f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa357_y2;
  wire f_s_dadda_pg_rca32_fa373_y2;
  wire f_s_dadda_pg_rca32_fa373_y3;
  wire f_s_dadda_pg_rca32_fa373_y4;
  wire f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa358_y2;
  wire f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa359_y2;
  wire f_s_dadda_pg_rca32_fa374_y0;
  wire f_s_dadda_pg_rca32_fa374_y1;
  wire f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa360_y2;
  wire f_s_dadda_pg_rca32_fa374_y2;
  wire f_s_dadda_pg_rca32_fa374_y3;
  wire f_s_dadda_pg_rca32_fa374_y4;
  wire f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa361_y2;
  wire f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa362_y2;
  wire f_s_dadda_pg_rca32_fa375_y0;
  wire f_s_dadda_pg_rca32_fa375_y1;
  wire f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa363_y2;
  wire f_s_dadda_pg_rca32_fa375_y2;
  wire f_s_dadda_pg_rca32_fa375_y3;
  wire f_s_dadda_pg_rca32_fa375_y4;
  wire f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa364_y2;
  wire f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa365_y2;
  wire f_s_dadda_pg_rca32_fa376_y0;
  wire f_s_dadda_pg_rca32_fa376_y1;
  wire f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa366_y2;
  wire f_s_dadda_pg_rca32_fa376_y2;
  wire f_s_dadda_pg_rca32_fa376_y3;
  wire f_s_dadda_pg_rca32_fa376_y4;
  wire f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa367_y2;
  wire f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa368_y2;
  wire f_s_dadda_pg_rca32_fa377_y0;
  wire f_s_dadda_pg_rca32_fa377_y1;
  wire f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa369_y2;
  wire f_s_dadda_pg_rca32_fa377_y2;
  wire f_s_dadda_pg_rca32_fa377_y3;
  wire f_s_dadda_pg_rca32_fa377_y4;
  wire f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa370_y2;
  wire f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa371_y2;
  wire f_s_dadda_pg_rca32_fa378_y0;
  wire f_s_dadda_pg_rca32_fa378_y1;
  wire f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa372_y2;
  wire f_s_dadda_pg_rca32_fa378_y2;
  wire f_s_dadda_pg_rca32_fa378_y3;
  wire f_s_dadda_pg_rca32_fa378_y4;
  wire f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa378_y4;
  wire f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa377_y4;
  wire f_s_dadda_pg_rca32_fa379_y0;
  wire f_s_dadda_pg_rca32_fa379_y1;
  wire f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa376_y4;
  wire f_s_dadda_pg_rca32_fa379_y2;
  wire f_s_dadda_pg_rca32_fa379_y3;
  wire f_s_dadda_pg_rca32_fa379_y4;
  wire f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa375_y4;
  wire f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa374_y4;
  wire f_s_dadda_pg_rca32_fa380_y0;
  wire f_s_dadda_pg_rca32_fa380_y1;
  wire f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa373_y4;
  wire f_s_dadda_pg_rca32_fa380_y2;
  wire f_s_dadda_pg_rca32_fa380_y3;
  wire f_s_dadda_pg_rca32_fa380_y4;
  wire f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa372_y4;
  wire f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa371_y4;
  wire f_s_dadda_pg_rca32_fa381_y0;
  wire f_s_dadda_pg_rca32_fa381_y1;
  wire f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa370_y4;
  wire f_s_dadda_pg_rca32_fa381_y2;
  wire f_s_dadda_pg_rca32_fa381_y3;
  wire f_s_dadda_pg_rca32_fa381_y4;
  wire f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa369_y4;
  wire f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa368_y4;
  wire f_s_dadda_pg_rca32_fa382_y0;
  wire f_s_dadda_pg_rca32_fa382_y1;
  wire f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa367_y4;
  wire f_s_dadda_pg_rca32_fa382_y2;
  wire f_s_dadda_pg_rca32_fa382_y3;
  wire f_s_dadda_pg_rca32_fa382_y4;
  wire f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa366_y4;
  wire f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa365_y4;
  wire f_s_dadda_pg_rca32_fa383_y0;
  wire f_s_dadda_pg_rca32_fa383_y1;
  wire f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa364_y4;
  wire f_s_dadda_pg_rca32_fa383_y2;
  wire f_s_dadda_pg_rca32_fa383_y3;
  wire f_s_dadda_pg_rca32_fa383_y4;
  wire f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa363_y4;
  wire f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa362_y4;
  wire f_s_dadda_pg_rca32_fa384_y0;
  wire f_s_dadda_pg_rca32_fa384_y1;
  wire f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa361_y4;
  wire f_s_dadda_pg_rca32_fa384_y2;
  wire f_s_dadda_pg_rca32_fa384_y3;
  wire f_s_dadda_pg_rca32_fa384_y4;
  wire f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa360_y4;
  wire f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa359_y4;
  wire f_s_dadda_pg_rca32_fa385_y0;
  wire f_s_dadda_pg_rca32_fa385_y1;
  wire f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa358_y4;
  wire f_s_dadda_pg_rca32_fa385_y2;
  wire f_s_dadda_pg_rca32_fa385_y3;
  wire f_s_dadda_pg_rca32_fa385_y4;
  wire f_s_dadda_pg_rca32_and_28_6_a_28;
  wire f_s_dadda_pg_rca32_and_28_6_b_6;
  wire f_s_dadda_pg_rca32_and_28_6_y0;
  wire f_s_dadda_pg_rca32_and_27_7_a_27;
  wire f_s_dadda_pg_rca32_and_27_7_b_7;
  wire f_s_dadda_pg_rca32_and_27_7_y0;
  wire f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_fa357_y4;
  wire f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_and_28_6_y0;
  wire f_s_dadda_pg_rca32_fa386_y0;
  wire f_s_dadda_pg_rca32_fa386_y1;
  wire f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_and_27_7_y0;
  wire f_s_dadda_pg_rca32_fa386_y2;
  wire f_s_dadda_pg_rca32_fa386_y3;
  wire f_s_dadda_pg_rca32_fa386_y4;
  wire f_s_dadda_pg_rca32_and_26_8_a_26;
  wire f_s_dadda_pg_rca32_and_26_8_b_8;
  wire f_s_dadda_pg_rca32_and_26_8_y0;
  wire f_s_dadda_pg_rca32_and_25_9_a_25;
  wire f_s_dadda_pg_rca32_and_25_9_b_9;
  wire f_s_dadda_pg_rca32_and_25_9_y0;
  wire f_s_dadda_pg_rca32_and_24_10_a_24;
  wire f_s_dadda_pg_rca32_and_24_10_b_10;
  wire f_s_dadda_pg_rca32_and_24_10_y0;
  wire f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_26_8_y0;
  wire f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_25_9_y0;
  wire f_s_dadda_pg_rca32_fa387_y0;
  wire f_s_dadda_pg_rca32_fa387_y1;
  wire f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_24_10_y0;
  wire f_s_dadda_pg_rca32_fa387_y2;
  wire f_s_dadda_pg_rca32_fa387_y3;
  wire f_s_dadda_pg_rca32_fa387_y4;
  wire f_s_dadda_pg_rca32_and_23_11_a_23;
  wire f_s_dadda_pg_rca32_and_23_11_b_11;
  wire f_s_dadda_pg_rca32_and_23_11_y0;
  wire f_s_dadda_pg_rca32_and_22_12_a_22;
  wire f_s_dadda_pg_rca32_and_22_12_b_12;
  wire f_s_dadda_pg_rca32_and_22_12_y0;
  wire f_s_dadda_pg_rca32_and_21_13_a_21;
  wire f_s_dadda_pg_rca32_and_21_13_b_13;
  wire f_s_dadda_pg_rca32_and_21_13_y0;
  wire f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_23_11_y0;
  wire f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_22_12_y0;
  wire f_s_dadda_pg_rca32_fa388_y0;
  wire f_s_dadda_pg_rca32_fa388_y1;
  wire f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_21_13_y0;
  wire f_s_dadda_pg_rca32_fa388_y2;
  wire f_s_dadda_pg_rca32_fa388_y3;
  wire f_s_dadda_pg_rca32_fa388_y4;
  wire f_s_dadda_pg_rca32_and_20_14_a_20;
  wire f_s_dadda_pg_rca32_and_20_14_b_14;
  wire f_s_dadda_pg_rca32_and_20_14_y0;
  wire f_s_dadda_pg_rca32_and_19_15_a_19;
  wire f_s_dadda_pg_rca32_and_19_15_b_15;
  wire f_s_dadda_pg_rca32_and_19_15_y0;
  wire f_s_dadda_pg_rca32_and_18_16_a_18;
  wire f_s_dadda_pg_rca32_and_18_16_b_16;
  wire f_s_dadda_pg_rca32_and_18_16_y0;
  wire f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_20_14_y0;
  wire f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_19_15_y0;
  wire f_s_dadda_pg_rca32_fa389_y0;
  wire f_s_dadda_pg_rca32_fa389_y1;
  wire f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_18_16_y0;
  wire f_s_dadda_pg_rca32_fa389_y2;
  wire f_s_dadda_pg_rca32_fa389_y3;
  wire f_s_dadda_pg_rca32_fa389_y4;
  wire f_s_dadda_pg_rca32_and_17_17_a_17;
  wire f_s_dadda_pg_rca32_and_17_17_b_17;
  wire f_s_dadda_pg_rca32_and_17_17_y0;
  wire f_s_dadda_pg_rca32_and_16_18_a_16;
  wire f_s_dadda_pg_rca32_and_16_18_b_18;
  wire f_s_dadda_pg_rca32_and_16_18_y0;
  wire f_s_dadda_pg_rca32_and_15_19_a_15;
  wire f_s_dadda_pg_rca32_and_15_19_b_19;
  wire f_s_dadda_pg_rca32_and_15_19_y0;
  wire f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_17_17_y0;
  wire f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_16_18_y0;
  wire f_s_dadda_pg_rca32_fa390_y0;
  wire f_s_dadda_pg_rca32_fa390_y1;
  wire f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_15_19_y0;
  wire f_s_dadda_pg_rca32_fa390_y2;
  wire f_s_dadda_pg_rca32_fa390_y3;
  wire f_s_dadda_pg_rca32_fa390_y4;
  wire f_s_dadda_pg_rca32_and_14_20_a_14;
  wire f_s_dadda_pg_rca32_and_14_20_b_20;
  wire f_s_dadda_pg_rca32_and_14_20_y0;
  wire f_s_dadda_pg_rca32_and_13_21_a_13;
  wire f_s_dadda_pg_rca32_and_13_21_b_21;
  wire f_s_dadda_pg_rca32_and_13_21_y0;
  wire f_s_dadda_pg_rca32_and_12_22_a_12;
  wire f_s_dadda_pg_rca32_and_12_22_b_22;
  wire f_s_dadda_pg_rca32_and_12_22_y0;
  wire f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_14_20_y0;
  wire f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_13_21_y0;
  wire f_s_dadda_pg_rca32_fa391_y0;
  wire f_s_dadda_pg_rca32_fa391_y1;
  wire f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_12_22_y0;
  wire f_s_dadda_pg_rca32_fa391_y2;
  wire f_s_dadda_pg_rca32_fa391_y3;
  wire f_s_dadda_pg_rca32_fa391_y4;
  wire f_s_dadda_pg_rca32_and_11_23_a_11;
  wire f_s_dadda_pg_rca32_and_11_23_b_23;
  wire f_s_dadda_pg_rca32_and_11_23_y0;
  wire f_s_dadda_pg_rca32_and_10_24_a_10;
  wire f_s_dadda_pg_rca32_and_10_24_b_24;
  wire f_s_dadda_pg_rca32_and_10_24_y0;
  wire f_s_dadda_pg_rca32_and_9_25_a_9;
  wire f_s_dadda_pg_rca32_and_9_25_b_25;
  wire f_s_dadda_pg_rca32_and_9_25_y0;
  wire f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_11_23_y0;
  wire f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_10_24_y0;
  wire f_s_dadda_pg_rca32_fa392_y0;
  wire f_s_dadda_pg_rca32_fa392_y1;
  wire f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_9_25_y0;
  wire f_s_dadda_pg_rca32_fa392_y2;
  wire f_s_dadda_pg_rca32_fa392_y3;
  wire f_s_dadda_pg_rca32_fa392_y4;
  wire f_s_dadda_pg_rca32_and_8_26_a_8;
  wire f_s_dadda_pg_rca32_and_8_26_b_26;
  wire f_s_dadda_pg_rca32_and_8_26_y0;
  wire f_s_dadda_pg_rca32_and_7_27_a_7;
  wire f_s_dadda_pg_rca32_and_7_27_b_27;
  wire f_s_dadda_pg_rca32_and_7_27_y0;
  wire f_s_dadda_pg_rca32_and_6_28_a_6;
  wire f_s_dadda_pg_rca32_and_6_28_b_28;
  wire f_s_dadda_pg_rca32_and_6_28_y0;
  wire f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_8_26_y0;
  wire f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_7_27_y0;
  wire f_s_dadda_pg_rca32_fa393_y0;
  wire f_s_dadda_pg_rca32_fa393_y1;
  wire f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_6_28_y0;
  wire f_s_dadda_pg_rca32_fa393_y2;
  wire f_s_dadda_pg_rca32_fa393_y3;
  wire f_s_dadda_pg_rca32_fa393_y4;
  wire f_s_dadda_pg_rca32_and_5_29_a_5;
  wire f_s_dadda_pg_rca32_and_5_29_b_29;
  wire f_s_dadda_pg_rca32_and_5_29_y0;
  wire f_s_dadda_pg_rca32_and_4_30_a_4;
  wire f_s_dadda_pg_rca32_and_4_30_b_30;
  wire f_s_dadda_pg_rca32_and_4_30_y0;
  wire f_s_dadda_pg_rca32_nand_3_31_a_3;
  wire f_s_dadda_pg_rca32_nand_3_31_b_31;
  wire f_s_dadda_pg_rca32_nand_3_31_y0;
  wire f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_and_5_29_y0;
  wire f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_and_4_30_y0;
  wire f_s_dadda_pg_rca32_fa394_y0;
  wire f_s_dadda_pg_rca32_fa394_y1;
  wire f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_nand_3_31_y0;
  wire f_s_dadda_pg_rca32_fa394_y2;
  wire f_s_dadda_pg_rca32_fa394_y3;
  wire f_s_dadda_pg_rca32_fa394_y4;
  wire f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa13_y2;
  wire f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa14_y2;
  wire f_s_dadda_pg_rca32_fa395_y0;
  wire f_s_dadda_pg_rca32_fa395_y1;
  wire f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa379_y2;
  wire f_s_dadda_pg_rca32_fa395_y2;
  wire f_s_dadda_pg_rca32_fa395_y3;
  wire f_s_dadda_pg_rca32_fa395_y4;
  wire f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa380_y2;
  wire f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa381_y2;
  wire f_s_dadda_pg_rca32_fa396_y0;
  wire f_s_dadda_pg_rca32_fa396_y1;
  wire f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa382_y2;
  wire f_s_dadda_pg_rca32_fa396_y2;
  wire f_s_dadda_pg_rca32_fa396_y3;
  wire f_s_dadda_pg_rca32_fa396_y4;
  wire f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa383_y2;
  wire f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa384_y2;
  wire f_s_dadda_pg_rca32_fa397_y0;
  wire f_s_dadda_pg_rca32_fa397_y1;
  wire f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa385_y2;
  wire f_s_dadda_pg_rca32_fa397_y2;
  wire f_s_dadda_pg_rca32_fa397_y3;
  wire f_s_dadda_pg_rca32_fa397_y4;
  wire f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa386_y2;
  wire f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa387_y2;
  wire f_s_dadda_pg_rca32_fa398_y0;
  wire f_s_dadda_pg_rca32_fa398_y1;
  wire f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa388_y2;
  wire f_s_dadda_pg_rca32_fa398_y2;
  wire f_s_dadda_pg_rca32_fa398_y3;
  wire f_s_dadda_pg_rca32_fa398_y4;
  wire f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa389_y2;
  wire f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa390_y2;
  wire f_s_dadda_pg_rca32_fa399_y0;
  wire f_s_dadda_pg_rca32_fa399_y1;
  wire f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa391_y2;
  wire f_s_dadda_pg_rca32_fa399_y2;
  wire f_s_dadda_pg_rca32_fa399_y3;
  wire f_s_dadda_pg_rca32_fa399_y4;
  wire f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa392_y2;
  wire f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa393_y2;
  wire f_s_dadda_pg_rca32_fa400_y0;
  wire f_s_dadda_pg_rca32_fa400_y1;
  wire f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa394_y2;
  wire f_s_dadda_pg_rca32_fa400_y2;
  wire f_s_dadda_pg_rca32_fa400_y3;
  wire f_s_dadda_pg_rca32_fa400_y4;
  wire f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa400_y4;
  wire f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa399_y4;
  wire f_s_dadda_pg_rca32_fa401_y0;
  wire f_s_dadda_pg_rca32_fa401_y1;
  wire f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa398_y4;
  wire f_s_dadda_pg_rca32_fa401_y2;
  wire f_s_dadda_pg_rca32_fa401_y3;
  wire f_s_dadda_pg_rca32_fa401_y4;
  wire f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa397_y4;
  wire f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa396_y4;
  wire f_s_dadda_pg_rca32_fa402_y0;
  wire f_s_dadda_pg_rca32_fa402_y1;
  wire f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa395_y4;
  wire f_s_dadda_pg_rca32_fa402_y2;
  wire f_s_dadda_pg_rca32_fa402_y3;
  wire f_s_dadda_pg_rca32_fa402_y4;
  wire f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa394_y4;
  wire f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa393_y4;
  wire f_s_dadda_pg_rca32_fa403_y0;
  wire f_s_dadda_pg_rca32_fa403_y1;
  wire f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa392_y4;
  wire f_s_dadda_pg_rca32_fa403_y2;
  wire f_s_dadda_pg_rca32_fa403_y3;
  wire f_s_dadda_pg_rca32_fa403_y4;
  wire f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa391_y4;
  wire f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa390_y4;
  wire f_s_dadda_pg_rca32_fa404_y0;
  wire f_s_dadda_pg_rca32_fa404_y1;
  wire f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa389_y4;
  wire f_s_dadda_pg_rca32_fa404_y2;
  wire f_s_dadda_pg_rca32_fa404_y3;
  wire f_s_dadda_pg_rca32_fa404_y4;
  wire f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa388_y4;
  wire f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa387_y4;
  wire f_s_dadda_pg_rca32_fa405_y0;
  wire f_s_dadda_pg_rca32_fa405_y1;
  wire f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa386_y4;
  wire f_s_dadda_pg_rca32_fa405_y2;
  wire f_s_dadda_pg_rca32_fa405_y3;
  wire f_s_dadda_pg_rca32_fa405_y4;
  wire f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa385_y4;
  wire f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa384_y4;
  wire f_s_dadda_pg_rca32_fa406_y0;
  wire f_s_dadda_pg_rca32_fa406_y1;
  wire f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa383_y4;
  wire f_s_dadda_pg_rca32_fa406_y2;
  wire f_s_dadda_pg_rca32_fa406_y3;
  wire f_s_dadda_pg_rca32_fa406_y4;
  wire f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa382_y4;
  wire f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa381_y4;
  wire f_s_dadda_pg_rca32_fa407_y0;
  wire f_s_dadda_pg_rca32_fa407_y1;
  wire f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa380_y4;
  wire f_s_dadda_pg_rca32_fa407_y2;
  wire f_s_dadda_pg_rca32_fa407_y3;
  wire f_s_dadda_pg_rca32_fa407_y4;
  wire f_s_dadda_pg_rca32_and_30_5_a_30;
  wire f_s_dadda_pg_rca32_and_30_5_b_5;
  wire f_s_dadda_pg_rca32_and_30_5_y0;
  wire f_s_dadda_pg_rca32_and_29_6_a_29;
  wire f_s_dadda_pg_rca32_and_29_6_b_6;
  wire f_s_dadda_pg_rca32_and_29_6_y0;
  wire f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_fa379_y4;
  wire f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_and_30_5_y0;
  wire f_s_dadda_pg_rca32_fa408_y0;
  wire f_s_dadda_pg_rca32_fa408_y1;
  wire f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_and_29_6_y0;
  wire f_s_dadda_pg_rca32_fa408_y2;
  wire f_s_dadda_pg_rca32_fa408_y3;
  wire f_s_dadda_pg_rca32_fa408_y4;
  wire f_s_dadda_pg_rca32_and_28_7_a_28;
  wire f_s_dadda_pg_rca32_and_28_7_b_7;
  wire f_s_dadda_pg_rca32_and_28_7_y0;
  wire f_s_dadda_pg_rca32_and_27_8_a_27;
  wire f_s_dadda_pg_rca32_and_27_8_b_8;
  wire f_s_dadda_pg_rca32_and_27_8_y0;
  wire f_s_dadda_pg_rca32_and_26_9_a_26;
  wire f_s_dadda_pg_rca32_and_26_9_b_9;
  wire f_s_dadda_pg_rca32_and_26_9_y0;
  wire f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_28_7_y0;
  wire f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_27_8_y0;
  wire f_s_dadda_pg_rca32_fa409_y0;
  wire f_s_dadda_pg_rca32_fa409_y1;
  wire f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_26_9_y0;
  wire f_s_dadda_pg_rca32_fa409_y2;
  wire f_s_dadda_pg_rca32_fa409_y3;
  wire f_s_dadda_pg_rca32_fa409_y4;
  wire f_s_dadda_pg_rca32_and_25_10_a_25;
  wire f_s_dadda_pg_rca32_and_25_10_b_10;
  wire f_s_dadda_pg_rca32_and_25_10_y0;
  wire f_s_dadda_pg_rca32_and_24_11_a_24;
  wire f_s_dadda_pg_rca32_and_24_11_b_11;
  wire f_s_dadda_pg_rca32_and_24_11_y0;
  wire f_s_dadda_pg_rca32_and_23_12_a_23;
  wire f_s_dadda_pg_rca32_and_23_12_b_12;
  wire f_s_dadda_pg_rca32_and_23_12_y0;
  wire f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_25_10_y0;
  wire f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_24_11_y0;
  wire f_s_dadda_pg_rca32_fa410_y0;
  wire f_s_dadda_pg_rca32_fa410_y1;
  wire f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_23_12_y0;
  wire f_s_dadda_pg_rca32_fa410_y2;
  wire f_s_dadda_pg_rca32_fa410_y3;
  wire f_s_dadda_pg_rca32_fa410_y4;
  wire f_s_dadda_pg_rca32_and_22_13_a_22;
  wire f_s_dadda_pg_rca32_and_22_13_b_13;
  wire f_s_dadda_pg_rca32_and_22_13_y0;
  wire f_s_dadda_pg_rca32_and_21_14_a_21;
  wire f_s_dadda_pg_rca32_and_21_14_b_14;
  wire f_s_dadda_pg_rca32_and_21_14_y0;
  wire f_s_dadda_pg_rca32_and_20_15_a_20;
  wire f_s_dadda_pg_rca32_and_20_15_b_15;
  wire f_s_dadda_pg_rca32_and_20_15_y0;
  wire f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_22_13_y0;
  wire f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_21_14_y0;
  wire f_s_dadda_pg_rca32_fa411_y0;
  wire f_s_dadda_pg_rca32_fa411_y1;
  wire f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_20_15_y0;
  wire f_s_dadda_pg_rca32_fa411_y2;
  wire f_s_dadda_pg_rca32_fa411_y3;
  wire f_s_dadda_pg_rca32_fa411_y4;
  wire f_s_dadda_pg_rca32_and_19_16_a_19;
  wire f_s_dadda_pg_rca32_and_19_16_b_16;
  wire f_s_dadda_pg_rca32_and_19_16_y0;
  wire f_s_dadda_pg_rca32_and_18_17_a_18;
  wire f_s_dadda_pg_rca32_and_18_17_b_17;
  wire f_s_dadda_pg_rca32_and_18_17_y0;
  wire f_s_dadda_pg_rca32_and_17_18_a_17;
  wire f_s_dadda_pg_rca32_and_17_18_b_18;
  wire f_s_dadda_pg_rca32_and_17_18_y0;
  wire f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_19_16_y0;
  wire f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_18_17_y0;
  wire f_s_dadda_pg_rca32_fa412_y0;
  wire f_s_dadda_pg_rca32_fa412_y1;
  wire f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_17_18_y0;
  wire f_s_dadda_pg_rca32_fa412_y2;
  wire f_s_dadda_pg_rca32_fa412_y3;
  wire f_s_dadda_pg_rca32_fa412_y4;
  wire f_s_dadda_pg_rca32_and_16_19_a_16;
  wire f_s_dadda_pg_rca32_and_16_19_b_19;
  wire f_s_dadda_pg_rca32_and_16_19_y0;
  wire f_s_dadda_pg_rca32_and_15_20_a_15;
  wire f_s_dadda_pg_rca32_and_15_20_b_20;
  wire f_s_dadda_pg_rca32_and_15_20_y0;
  wire f_s_dadda_pg_rca32_and_14_21_a_14;
  wire f_s_dadda_pg_rca32_and_14_21_b_21;
  wire f_s_dadda_pg_rca32_and_14_21_y0;
  wire f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_16_19_y0;
  wire f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_15_20_y0;
  wire f_s_dadda_pg_rca32_fa413_y0;
  wire f_s_dadda_pg_rca32_fa413_y1;
  wire f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_14_21_y0;
  wire f_s_dadda_pg_rca32_fa413_y2;
  wire f_s_dadda_pg_rca32_fa413_y3;
  wire f_s_dadda_pg_rca32_fa413_y4;
  wire f_s_dadda_pg_rca32_and_13_22_a_13;
  wire f_s_dadda_pg_rca32_and_13_22_b_22;
  wire f_s_dadda_pg_rca32_and_13_22_y0;
  wire f_s_dadda_pg_rca32_and_12_23_a_12;
  wire f_s_dadda_pg_rca32_and_12_23_b_23;
  wire f_s_dadda_pg_rca32_and_12_23_y0;
  wire f_s_dadda_pg_rca32_and_11_24_a_11;
  wire f_s_dadda_pg_rca32_and_11_24_b_24;
  wire f_s_dadda_pg_rca32_and_11_24_y0;
  wire f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_13_22_y0;
  wire f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_12_23_y0;
  wire f_s_dadda_pg_rca32_fa414_y0;
  wire f_s_dadda_pg_rca32_fa414_y1;
  wire f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_11_24_y0;
  wire f_s_dadda_pg_rca32_fa414_y2;
  wire f_s_dadda_pg_rca32_fa414_y3;
  wire f_s_dadda_pg_rca32_fa414_y4;
  wire f_s_dadda_pg_rca32_and_10_25_a_10;
  wire f_s_dadda_pg_rca32_and_10_25_b_25;
  wire f_s_dadda_pg_rca32_and_10_25_y0;
  wire f_s_dadda_pg_rca32_and_9_26_a_9;
  wire f_s_dadda_pg_rca32_and_9_26_b_26;
  wire f_s_dadda_pg_rca32_and_9_26_y0;
  wire f_s_dadda_pg_rca32_and_8_27_a_8;
  wire f_s_dadda_pg_rca32_and_8_27_b_27;
  wire f_s_dadda_pg_rca32_and_8_27_y0;
  wire f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_10_25_y0;
  wire f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_9_26_y0;
  wire f_s_dadda_pg_rca32_fa415_y0;
  wire f_s_dadda_pg_rca32_fa415_y1;
  wire f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_8_27_y0;
  wire f_s_dadda_pg_rca32_fa415_y2;
  wire f_s_dadda_pg_rca32_fa415_y3;
  wire f_s_dadda_pg_rca32_fa415_y4;
  wire f_s_dadda_pg_rca32_and_7_28_a_7;
  wire f_s_dadda_pg_rca32_and_7_28_b_28;
  wire f_s_dadda_pg_rca32_and_7_28_y0;
  wire f_s_dadda_pg_rca32_and_6_29_a_6;
  wire f_s_dadda_pg_rca32_and_6_29_b_29;
  wire f_s_dadda_pg_rca32_and_6_29_y0;
  wire f_s_dadda_pg_rca32_and_5_30_a_5;
  wire f_s_dadda_pg_rca32_and_5_30_b_30;
  wire f_s_dadda_pg_rca32_and_5_30_y0;
  wire f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_7_28_y0;
  wire f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_6_29_y0;
  wire f_s_dadda_pg_rca32_fa416_y0;
  wire f_s_dadda_pg_rca32_fa416_y1;
  wire f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_5_30_y0;
  wire f_s_dadda_pg_rca32_fa416_y2;
  wire f_s_dadda_pg_rca32_fa416_y3;
  wire f_s_dadda_pg_rca32_fa416_y4;
  wire f_s_dadda_pg_rca32_nand_4_31_a_4;
  wire f_s_dadda_pg_rca32_nand_4_31_b_31;
  wire f_s_dadda_pg_rca32_nand_4_31_y0;
  wire f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_nand_4_31_y0;
  wire f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_fa15_y2;
  wire f_s_dadda_pg_rca32_fa417_y0;
  wire f_s_dadda_pg_rca32_fa417_y1;
  wire f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_fa401_y2;
  wire f_s_dadda_pg_rca32_fa417_y2;
  wire f_s_dadda_pg_rca32_fa417_y3;
  wire f_s_dadda_pg_rca32_fa417_y4;
  wire f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa402_y2;
  wire f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa403_y2;
  wire f_s_dadda_pg_rca32_fa418_y0;
  wire f_s_dadda_pg_rca32_fa418_y1;
  wire f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa404_y2;
  wire f_s_dadda_pg_rca32_fa418_y2;
  wire f_s_dadda_pg_rca32_fa418_y3;
  wire f_s_dadda_pg_rca32_fa418_y4;
  wire f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa405_y2;
  wire f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa406_y2;
  wire f_s_dadda_pg_rca32_fa419_y0;
  wire f_s_dadda_pg_rca32_fa419_y1;
  wire f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa407_y2;
  wire f_s_dadda_pg_rca32_fa419_y2;
  wire f_s_dadda_pg_rca32_fa419_y3;
  wire f_s_dadda_pg_rca32_fa419_y4;
  wire f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa408_y2;
  wire f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa409_y2;
  wire f_s_dadda_pg_rca32_fa420_y0;
  wire f_s_dadda_pg_rca32_fa420_y1;
  wire f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa410_y2;
  wire f_s_dadda_pg_rca32_fa420_y2;
  wire f_s_dadda_pg_rca32_fa420_y3;
  wire f_s_dadda_pg_rca32_fa420_y4;
  wire f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa411_y2;
  wire f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa412_y2;
  wire f_s_dadda_pg_rca32_fa421_y0;
  wire f_s_dadda_pg_rca32_fa421_y1;
  wire f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa413_y2;
  wire f_s_dadda_pg_rca32_fa421_y2;
  wire f_s_dadda_pg_rca32_fa421_y3;
  wire f_s_dadda_pg_rca32_fa421_y4;
  wire f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa414_y2;
  wire f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa415_y2;
  wire f_s_dadda_pg_rca32_fa422_y0;
  wire f_s_dadda_pg_rca32_fa422_y1;
  wire f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa416_y2;
  wire f_s_dadda_pg_rca32_fa422_y2;
  wire f_s_dadda_pg_rca32_fa422_y3;
  wire f_s_dadda_pg_rca32_fa422_y4;
  wire f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa422_y4;
  wire f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa421_y4;
  wire f_s_dadda_pg_rca32_fa423_y0;
  wire f_s_dadda_pg_rca32_fa423_y1;
  wire f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa420_y4;
  wire f_s_dadda_pg_rca32_fa423_y2;
  wire f_s_dadda_pg_rca32_fa423_y3;
  wire f_s_dadda_pg_rca32_fa423_y4;
  wire f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa419_y4;
  wire f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa418_y4;
  wire f_s_dadda_pg_rca32_fa424_y0;
  wire f_s_dadda_pg_rca32_fa424_y1;
  wire f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa417_y4;
  wire f_s_dadda_pg_rca32_fa424_y2;
  wire f_s_dadda_pg_rca32_fa424_y3;
  wire f_s_dadda_pg_rca32_fa424_y4;
  wire f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa416_y4;
  wire f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa415_y4;
  wire f_s_dadda_pg_rca32_fa425_y0;
  wire f_s_dadda_pg_rca32_fa425_y1;
  wire f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa414_y4;
  wire f_s_dadda_pg_rca32_fa425_y2;
  wire f_s_dadda_pg_rca32_fa425_y3;
  wire f_s_dadda_pg_rca32_fa425_y4;
  wire f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa413_y4;
  wire f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa412_y4;
  wire f_s_dadda_pg_rca32_fa426_y0;
  wire f_s_dadda_pg_rca32_fa426_y1;
  wire f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa411_y4;
  wire f_s_dadda_pg_rca32_fa426_y2;
  wire f_s_dadda_pg_rca32_fa426_y3;
  wire f_s_dadda_pg_rca32_fa426_y4;
  wire f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa410_y4;
  wire f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa409_y4;
  wire f_s_dadda_pg_rca32_fa427_y0;
  wire f_s_dadda_pg_rca32_fa427_y1;
  wire f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa408_y4;
  wire f_s_dadda_pg_rca32_fa427_y2;
  wire f_s_dadda_pg_rca32_fa427_y3;
  wire f_s_dadda_pg_rca32_fa427_y4;
  wire f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa407_y4;
  wire f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa406_y4;
  wire f_s_dadda_pg_rca32_fa428_y0;
  wire f_s_dadda_pg_rca32_fa428_y1;
  wire f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa405_y4;
  wire f_s_dadda_pg_rca32_fa428_y2;
  wire f_s_dadda_pg_rca32_fa428_y3;
  wire f_s_dadda_pg_rca32_fa428_y4;
  wire f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa404_y4;
  wire f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa403_y4;
  wire f_s_dadda_pg_rca32_fa429_y0;
  wire f_s_dadda_pg_rca32_fa429_y1;
  wire f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa402_y4;
  wire f_s_dadda_pg_rca32_fa429_y2;
  wire f_s_dadda_pg_rca32_fa429_y3;
  wire f_s_dadda_pg_rca32_fa429_y4;
  wire f_s_dadda_pg_rca32_nand_31_5_a_31;
  wire f_s_dadda_pg_rca32_nand_31_5_b_5;
  wire f_s_dadda_pg_rca32_nand_31_5_y0;
  wire f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_fa401_y4;
  wire f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_fa15_y4;
  wire f_s_dadda_pg_rca32_fa430_y0;
  wire f_s_dadda_pg_rca32_fa430_y1;
  wire f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_nand_31_5_y0;
  wire f_s_dadda_pg_rca32_fa430_y2;
  wire f_s_dadda_pg_rca32_fa430_y3;
  wire f_s_dadda_pg_rca32_fa430_y4;
  wire f_s_dadda_pg_rca32_and_30_6_a_30;
  wire f_s_dadda_pg_rca32_and_30_6_b_6;
  wire f_s_dadda_pg_rca32_and_30_6_y0;
  wire f_s_dadda_pg_rca32_and_29_7_a_29;
  wire f_s_dadda_pg_rca32_and_29_7_b_7;
  wire f_s_dadda_pg_rca32_and_29_7_y0;
  wire f_s_dadda_pg_rca32_and_28_8_a_28;
  wire f_s_dadda_pg_rca32_and_28_8_b_8;
  wire f_s_dadda_pg_rca32_and_28_8_y0;
  wire f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_30_6_y0;
  wire f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_29_7_y0;
  wire f_s_dadda_pg_rca32_fa431_y0;
  wire f_s_dadda_pg_rca32_fa431_y1;
  wire f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_28_8_y0;
  wire f_s_dadda_pg_rca32_fa431_y2;
  wire f_s_dadda_pg_rca32_fa431_y3;
  wire f_s_dadda_pg_rca32_fa431_y4;
  wire f_s_dadda_pg_rca32_and_27_9_a_27;
  wire f_s_dadda_pg_rca32_and_27_9_b_9;
  wire f_s_dadda_pg_rca32_and_27_9_y0;
  wire f_s_dadda_pg_rca32_and_26_10_a_26;
  wire f_s_dadda_pg_rca32_and_26_10_b_10;
  wire f_s_dadda_pg_rca32_and_26_10_y0;
  wire f_s_dadda_pg_rca32_and_25_11_a_25;
  wire f_s_dadda_pg_rca32_and_25_11_b_11;
  wire f_s_dadda_pg_rca32_and_25_11_y0;
  wire f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_27_9_y0;
  wire f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_26_10_y0;
  wire f_s_dadda_pg_rca32_fa432_y0;
  wire f_s_dadda_pg_rca32_fa432_y1;
  wire f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_25_11_y0;
  wire f_s_dadda_pg_rca32_fa432_y2;
  wire f_s_dadda_pg_rca32_fa432_y3;
  wire f_s_dadda_pg_rca32_fa432_y4;
  wire f_s_dadda_pg_rca32_and_24_12_a_24;
  wire f_s_dadda_pg_rca32_and_24_12_b_12;
  wire f_s_dadda_pg_rca32_and_24_12_y0;
  wire f_s_dadda_pg_rca32_and_23_13_a_23;
  wire f_s_dadda_pg_rca32_and_23_13_b_13;
  wire f_s_dadda_pg_rca32_and_23_13_y0;
  wire f_s_dadda_pg_rca32_and_22_14_a_22;
  wire f_s_dadda_pg_rca32_and_22_14_b_14;
  wire f_s_dadda_pg_rca32_and_22_14_y0;
  wire f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_24_12_y0;
  wire f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_23_13_y0;
  wire f_s_dadda_pg_rca32_fa433_y0;
  wire f_s_dadda_pg_rca32_fa433_y1;
  wire f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_22_14_y0;
  wire f_s_dadda_pg_rca32_fa433_y2;
  wire f_s_dadda_pg_rca32_fa433_y3;
  wire f_s_dadda_pg_rca32_fa433_y4;
  wire f_s_dadda_pg_rca32_and_21_15_a_21;
  wire f_s_dadda_pg_rca32_and_21_15_b_15;
  wire f_s_dadda_pg_rca32_and_21_15_y0;
  wire f_s_dadda_pg_rca32_and_20_16_a_20;
  wire f_s_dadda_pg_rca32_and_20_16_b_16;
  wire f_s_dadda_pg_rca32_and_20_16_y0;
  wire f_s_dadda_pg_rca32_and_19_17_a_19;
  wire f_s_dadda_pg_rca32_and_19_17_b_17;
  wire f_s_dadda_pg_rca32_and_19_17_y0;
  wire f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_21_15_y0;
  wire f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_20_16_y0;
  wire f_s_dadda_pg_rca32_fa434_y0;
  wire f_s_dadda_pg_rca32_fa434_y1;
  wire f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_19_17_y0;
  wire f_s_dadda_pg_rca32_fa434_y2;
  wire f_s_dadda_pg_rca32_fa434_y3;
  wire f_s_dadda_pg_rca32_fa434_y4;
  wire f_s_dadda_pg_rca32_and_18_18_a_18;
  wire f_s_dadda_pg_rca32_and_18_18_b_18;
  wire f_s_dadda_pg_rca32_and_18_18_y0;
  wire f_s_dadda_pg_rca32_and_17_19_a_17;
  wire f_s_dadda_pg_rca32_and_17_19_b_19;
  wire f_s_dadda_pg_rca32_and_17_19_y0;
  wire f_s_dadda_pg_rca32_and_16_20_a_16;
  wire f_s_dadda_pg_rca32_and_16_20_b_20;
  wire f_s_dadda_pg_rca32_and_16_20_y0;
  wire f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_18_18_y0;
  wire f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_17_19_y0;
  wire f_s_dadda_pg_rca32_fa435_y0;
  wire f_s_dadda_pg_rca32_fa435_y1;
  wire f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_16_20_y0;
  wire f_s_dadda_pg_rca32_fa435_y2;
  wire f_s_dadda_pg_rca32_fa435_y3;
  wire f_s_dadda_pg_rca32_fa435_y4;
  wire f_s_dadda_pg_rca32_and_15_21_a_15;
  wire f_s_dadda_pg_rca32_and_15_21_b_21;
  wire f_s_dadda_pg_rca32_and_15_21_y0;
  wire f_s_dadda_pg_rca32_and_14_22_a_14;
  wire f_s_dadda_pg_rca32_and_14_22_b_22;
  wire f_s_dadda_pg_rca32_and_14_22_y0;
  wire f_s_dadda_pg_rca32_and_13_23_a_13;
  wire f_s_dadda_pg_rca32_and_13_23_b_23;
  wire f_s_dadda_pg_rca32_and_13_23_y0;
  wire f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_15_21_y0;
  wire f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_14_22_y0;
  wire f_s_dadda_pg_rca32_fa436_y0;
  wire f_s_dadda_pg_rca32_fa436_y1;
  wire f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_13_23_y0;
  wire f_s_dadda_pg_rca32_fa436_y2;
  wire f_s_dadda_pg_rca32_fa436_y3;
  wire f_s_dadda_pg_rca32_fa436_y4;
  wire f_s_dadda_pg_rca32_and_12_24_a_12;
  wire f_s_dadda_pg_rca32_and_12_24_b_24;
  wire f_s_dadda_pg_rca32_and_12_24_y0;
  wire f_s_dadda_pg_rca32_and_11_25_a_11;
  wire f_s_dadda_pg_rca32_and_11_25_b_25;
  wire f_s_dadda_pg_rca32_and_11_25_y0;
  wire f_s_dadda_pg_rca32_and_10_26_a_10;
  wire f_s_dadda_pg_rca32_and_10_26_b_26;
  wire f_s_dadda_pg_rca32_and_10_26_y0;
  wire f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_12_24_y0;
  wire f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_11_25_y0;
  wire f_s_dadda_pg_rca32_fa437_y0;
  wire f_s_dadda_pg_rca32_fa437_y1;
  wire f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_10_26_y0;
  wire f_s_dadda_pg_rca32_fa437_y2;
  wire f_s_dadda_pg_rca32_fa437_y3;
  wire f_s_dadda_pg_rca32_fa437_y4;
  wire f_s_dadda_pg_rca32_and_9_27_a_9;
  wire f_s_dadda_pg_rca32_and_9_27_b_27;
  wire f_s_dadda_pg_rca32_and_9_27_y0;
  wire f_s_dadda_pg_rca32_and_8_28_a_8;
  wire f_s_dadda_pg_rca32_and_8_28_b_28;
  wire f_s_dadda_pg_rca32_and_8_28_y0;
  wire f_s_dadda_pg_rca32_and_7_29_a_7;
  wire f_s_dadda_pg_rca32_and_7_29_b_29;
  wire f_s_dadda_pg_rca32_and_7_29_y0;
  wire f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_9_27_y0;
  wire f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_8_28_y0;
  wire f_s_dadda_pg_rca32_fa438_y0;
  wire f_s_dadda_pg_rca32_fa438_y1;
  wire f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_7_29_y0;
  wire f_s_dadda_pg_rca32_fa438_y2;
  wire f_s_dadda_pg_rca32_fa438_y3;
  wire f_s_dadda_pg_rca32_fa438_y4;
  wire f_s_dadda_pg_rca32_and_6_30_a_6;
  wire f_s_dadda_pg_rca32_and_6_30_b_30;
  wire f_s_dadda_pg_rca32_and_6_30_y0;
  wire f_s_dadda_pg_rca32_nand_5_31_a_5;
  wire f_s_dadda_pg_rca32_nand_5_31_b_31;
  wire f_s_dadda_pg_rca32_nand_5_31_y0;
  wire f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_and_6_30_y0;
  wire f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_nand_5_31_y0;
  wire f_s_dadda_pg_rca32_fa439_y0;
  wire f_s_dadda_pg_rca32_fa439_y1;
  wire f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_fa423_y2;
  wire f_s_dadda_pg_rca32_fa439_y2;
  wire f_s_dadda_pg_rca32_fa439_y3;
  wire f_s_dadda_pg_rca32_fa439_y4;
  wire f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa424_y2;
  wire f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa425_y2;
  wire f_s_dadda_pg_rca32_fa440_y0;
  wire f_s_dadda_pg_rca32_fa440_y1;
  wire f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa426_y2;
  wire f_s_dadda_pg_rca32_fa440_y2;
  wire f_s_dadda_pg_rca32_fa440_y3;
  wire f_s_dadda_pg_rca32_fa440_y4;
  wire f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa427_y2;
  wire f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa428_y2;
  wire f_s_dadda_pg_rca32_fa441_y0;
  wire f_s_dadda_pg_rca32_fa441_y1;
  wire f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa429_y2;
  wire f_s_dadda_pg_rca32_fa441_y2;
  wire f_s_dadda_pg_rca32_fa441_y3;
  wire f_s_dadda_pg_rca32_fa441_y4;
  wire f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa430_y2;
  wire f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa431_y2;
  wire f_s_dadda_pg_rca32_fa442_y0;
  wire f_s_dadda_pg_rca32_fa442_y1;
  wire f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa432_y2;
  wire f_s_dadda_pg_rca32_fa442_y2;
  wire f_s_dadda_pg_rca32_fa442_y3;
  wire f_s_dadda_pg_rca32_fa442_y4;
  wire f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa433_y2;
  wire f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa434_y2;
  wire f_s_dadda_pg_rca32_fa443_y0;
  wire f_s_dadda_pg_rca32_fa443_y1;
  wire f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa435_y2;
  wire f_s_dadda_pg_rca32_fa443_y2;
  wire f_s_dadda_pg_rca32_fa443_y3;
  wire f_s_dadda_pg_rca32_fa443_y4;
  wire f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa436_y2;
  wire f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa437_y2;
  wire f_s_dadda_pg_rca32_fa444_y0;
  wire f_s_dadda_pg_rca32_fa444_y1;
  wire f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa438_y2;
  wire f_s_dadda_pg_rca32_fa444_y2;
  wire f_s_dadda_pg_rca32_fa444_y3;
  wire f_s_dadda_pg_rca32_fa444_y4;
  wire f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa444_y4;
  wire f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa443_y4;
  wire f_s_dadda_pg_rca32_fa445_y0;
  wire f_s_dadda_pg_rca32_fa445_y1;
  wire f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa442_y4;
  wire f_s_dadda_pg_rca32_fa445_y2;
  wire f_s_dadda_pg_rca32_fa445_y3;
  wire f_s_dadda_pg_rca32_fa445_y4;
  wire f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa441_y4;
  wire f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa440_y4;
  wire f_s_dadda_pg_rca32_fa446_y0;
  wire f_s_dadda_pg_rca32_fa446_y1;
  wire f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa439_y4;
  wire f_s_dadda_pg_rca32_fa446_y2;
  wire f_s_dadda_pg_rca32_fa446_y3;
  wire f_s_dadda_pg_rca32_fa446_y4;
  wire f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa438_y4;
  wire f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa437_y4;
  wire f_s_dadda_pg_rca32_fa447_y0;
  wire f_s_dadda_pg_rca32_fa447_y1;
  wire f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa436_y4;
  wire f_s_dadda_pg_rca32_fa447_y2;
  wire f_s_dadda_pg_rca32_fa447_y3;
  wire f_s_dadda_pg_rca32_fa447_y4;
  wire f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa435_y4;
  wire f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa434_y4;
  wire f_s_dadda_pg_rca32_fa448_y0;
  wire f_s_dadda_pg_rca32_fa448_y1;
  wire f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa433_y4;
  wire f_s_dadda_pg_rca32_fa448_y2;
  wire f_s_dadda_pg_rca32_fa448_y3;
  wire f_s_dadda_pg_rca32_fa448_y4;
  wire f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa432_y4;
  wire f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa431_y4;
  wire f_s_dadda_pg_rca32_fa449_y0;
  wire f_s_dadda_pg_rca32_fa449_y1;
  wire f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa430_y4;
  wire f_s_dadda_pg_rca32_fa449_y2;
  wire f_s_dadda_pg_rca32_fa449_y3;
  wire f_s_dadda_pg_rca32_fa449_y4;
  wire f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa429_y4;
  wire f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa428_y4;
  wire f_s_dadda_pg_rca32_fa450_y0;
  wire f_s_dadda_pg_rca32_fa450_y1;
  wire f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa427_y4;
  wire f_s_dadda_pg_rca32_fa450_y2;
  wire f_s_dadda_pg_rca32_fa450_y3;
  wire f_s_dadda_pg_rca32_fa450_y4;
  wire f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa426_y4;
  wire f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa425_y4;
  wire f_s_dadda_pg_rca32_fa451_y0;
  wire f_s_dadda_pg_rca32_fa451_y1;
  wire f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa424_y4;
  wire f_s_dadda_pg_rca32_fa451_y2;
  wire f_s_dadda_pg_rca32_fa451_y3;
  wire f_s_dadda_pg_rca32_fa451_y4;
  wire f_s_dadda_pg_rca32_nand_31_6_a_31;
  wire f_s_dadda_pg_rca32_nand_31_6_b_6;
  wire f_s_dadda_pg_rca32_nand_31_6_y0;
  wire f_s_dadda_pg_rca32_and_30_7_a_30;
  wire f_s_dadda_pg_rca32_and_30_7_b_7;
  wire f_s_dadda_pg_rca32_and_30_7_y0;
  wire f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_fa423_y4;
  wire f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_nand_31_6_y0;
  wire f_s_dadda_pg_rca32_fa452_y0;
  wire f_s_dadda_pg_rca32_fa452_y1;
  wire f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_and_30_7_y0;
  wire f_s_dadda_pg_rca32_fa452_y2;
  wire f_s_dadda_pg_rca32_fa452_y3;
  wire f_s_dadda_pg_rca32_fa452_y4;
  wire f_s_dadda_pg_rca32_and_29_8_a_29;
  wire f_s_dadda_pg_rca32_and_29_8_b_8;
  wire f_s_dadda_pg_rca32_and_29_8_y0;
  wire f_s_dadda_pg_rca32_and_28_9_a_28;
  wire f_s_dadda_pg_rca32_and_28_9_b_9;
  wire f_s_dadda_pg_rca32_and_28_9_y0;
  wire f_s_dadda_pg_rca32_and_27_10_a_27;
  wire f_s_dadda_pg_rca32_and_27_10_b_10;
  wire f_s_dadda_pg_rca32_and_27_10_y0;
  wire f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_29_8_y0;
  wire f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_28_9_y0;
  wire f_s_dadda_pg_rca32_fa453_y0;
  wire f_s_dadda_pg_rca32_fa453_y1;
  wire f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_27_10_y0;
  wire f_s_dadda_pg_rca32_fa453_y2;
  wire f_s_dadda_pg_rca32_fa453_y3;
  wire f_s_dadda_pg_rca32_fa453_y4;
  wire f_s_dadda_pg_rca32_and_26_11_a_26;
  wire f_s_dadda_pg_rca32_and_26_11_b_11;
  wire f_s_dadda_pg_rca32_and_26_11_y0;
  wire f_s_dadda_pg_rca32_and_25_12_a_25;
  wire f_s_dadda_pg_rca32_and_25_12_b_12;
  wire f_s_dadda_pg_rca32_and_25_12_y0;
  wire f_s_dadda_pg_rca32_and_24_13_a_24;
  wire f_s_dadda_pg_rca32_and_24_13_b_13;
  wire f_s_dadda_pg_rca32_and_24_13_y0;
  wire f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_26_11_y0;
  wire f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_25_12_y0;
  wire f_s_dadda_pg_rca32_fa454_y0;
  wire f_s_dadda_pg_rca32_fa454_y1;
  wire f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_24_13_y0;
  wire f_s_dadda_pg_rca32_fa454_y2;
  wire f_s_dadda_pg_rca32_fa454_y3;
  wire f_s_dadda_pg_rca32_fa454_y4;
  wire f_s_dadda_pg_rca32_and_23_14_a_23;
  wire f_s_dadda_pg_rca32_and_23_14_b_14;
  wire f_s_dadda_pg_rca32_and_23_14_y0;
  wire f_s_dadda_pg_rca32_and_22_15_a_22;
  wire f_s_dadda_pg_rca32_and_22_15_b_15;
  wire f_s_dadda_pg_rca32_and_22_15_y0;
  wire f_s_dadda_pg_rca32_and_21_16_a_21;
  wire f_s_dadda_pg_rca32_and_21_16_b_16;
  wire f_s_dadda_pg_rca32_and_21_16_y0;
  wire f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_23_14_y0;
  wire f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_22_15_y0;
  wire f_s_dadda_pg_rca32_fa455_y0;
  wire f_s_dadda_pg_rca32_fa455_y1;
  wire f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_21_16_y0;
  wire f_s_dadda_pg_rca32_fa455_y2;
  wire f_s_dadda_pg_rca32_fa455_y3;
  wire f_s_dadda_pg_rca32_fa455_y4;
  wire f_s_dadda_pg_rca32_and_20_17_a_20;
  wire f_s_dadda_pg_rca32_and_20_17_b_17;
  wire f_s_dadda_pg_rca32_and_20_17_y0;
  wire f_s_dadda_pg_rca32_and_19_18_a_19;
  wire f_s_dadda_pg_rca32_and_19_18_b_18;
  wire f_s_dadda_pg_rca32_and_19_18_y0;
  wire f_s_dadda_pg_rca32_and_18_19_a_18;
  wire f_s_dadda_pg_rca32_and_18_19_b_19;
  wire f_s_dadda_pg_rca32_and_18_19_y0;
  wire f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_20_17_y0;
  wire f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_19_18_y0;
  wire f_s_dadda_pg_rca32_fa456_y0;
  wire f_s_dadda_pg_rca32_fa456_y1;
  wire f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_18_19_y0;
  wire f_s_dadda_pg_rca32_fa456_y2;
  wire f_s_dadda_pg_rca32_fa456_y3;
  wire f_s_dadda_pg_rca32_fa456_y4;
  wire f_s_dadda_pg_rca32_and_17_20_a_17;
  wire f_s_dadda_pg_rca32_and_17_20_b_20;
  wire f_s_dadda_pg_rca32_and_17_20_y0;
  wire f_s_dadda_pg_rca32_and_16_21_a_16;
  wire f_s_dadda_pg_rca32_and_16_21_b_21;
  wire f_s_dadda_pg_rca32_and_16_21_y0;
  wire f_s_dadda_pg_rca32_and_15_22_a_15;
  wire f_s_dadda_pg_rca32_and_15_22_b_22;
  wire f_s_dadda_pg_rca32_and_15_22_y0;
  wire f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_17_20_y0;
  wire f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_16_21_y0;
  wire f_s_dadda_pg_rca32_fa457_y0;
  wire f_s_dadda_pg_rca32_fa457_y1;
  wire f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_15_22_y0;
  wire f_s_dadda_pg_rca32_fa457_y2;
  wire f_s_dadda_pg_rca32_fa457_y3;
  wire f_s_dadda_pg_rca32_fa457_y4;
  wire f_s_dadda_pg_rca32_and_14_23_a_14;
  wire f_s_dadda_pg_rca32_and_14_23_b_23;
  wire f_s_dadda_pg_rca32_and_14_23_y0;
  wire f_s_dadda_pg_rca32_and_13_24_a_13;
  wire f_s_dadda_pg_rca32_and_13_24_b_24;
  wire f_s_dadda_pg_rca32_and_13_24_y0;
  wire f_s_dadda_pg_rca32_and_12_25_a_12;
  wire f_s_dadda_pg_rca32_and_12_25_b_25;
  wire f_s_dadda_pg_rca32_and_12_25_y0;
  wire f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_14_23_y0;
  wire f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_13_24_y0;
  wire f_s_dadda_pg_rca32_fa458_y0;
  wire f_s_dadda_pg_rca32_fa458_y1;
  wire f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_12_25_y0;
  wire f_s_dadda_pg_rca32_fa458_y2;
  wire f_s_dadda_pg_rca32_fa458_y3;
  wire f_s_dadda_pg_rca32_fa458_y4;
  wire f_s_dadda_pg_rca32_and_11_26_a_11;
  wire f_s_dadda_pg_rca32_and_11_26_b_26;
  wire f_s_dadda_pg_rca32_and_11_26_y0;
  wire f_s_dadda_pg_rca32_and_10_27_a_10;
  wire f_s_dadda_pg_rca32_and_10_27_b_27;
  wire f_s_dadda_pg_rca32_and_10_27_y0;
  wire f_s_dadda_pg_rca32_and_9_28_a_9;
  wire f_s_dadda_pg_rca32_and_9_28_b_28;
  wire f_s_dadda_pg_rca32_and_9_28_y0;
  wire f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_11_26_y0;
  wire f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_10_27_y0;
  wire f_s_dadda_pg_rca32_fa459_y0;
  wire f_s_dadda_pg_rca32_fa459_y1;
  wire f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_9_28_y0;
  wire f_s_dadda_pg_rca32_fa459_y2;
  wire f_s_dadda_pg_rca32_fa459_y3;
  wire f_s_dadda_pg_rca32_fa459_y4;
  wire f_s_dadda_pg_rca32_and_8_29_a_8;
  wire f_s_dadda_pg_rca32_and_8_29_b_29;
  wire f_s_dadda_pg_rca32_and_8_29_y0;
  wire f_s_dadda_pg_rca32_and_7_30_a_7;
  wire f_s_dadda_pg_rca32_and_7_30_b_30;
  wire f_s_dadda_pg_rca32_and_7_30_y0;
  wire f_s_dadda_pg_rca32_nand_6_31_a_6;
  wire f_s_dadda_pg_rca32_nand_6_31_b_31;
  wire f_s_dadda_pg_rca32_nand_6_31_y0;
  wire f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_and_8_29_y0;
  wire f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_and_7_30_y0;
  wire f_s_dadda_pg_rca32_fa460_y0;
  wire f_s_dadda_pg_rca32_fa460_y1;
  wire f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_nand_6_31_y0;
  wire f_s_dadda_pg_rca32_fa460_y2;
  wire f_s_dadda_pg_rca32_fa460_y3;
  wire f_s_dadda_pg_rca32_fa460_y4;
  wire f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa445_y2;
  wire f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa446_y2;
  wire f_s_dadda_pg_rca32_fa461_y0;
  wire f_s_dadda_pg_rca32_fa461_y1;
  wire f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa447_y2;
  wire f_s_dadda_pg_rca32_fa461_y2;
  wire f_s_dadda_pg_rca32_fa461_y3;
  wire f_s_dadda_pg_rca32_fa461_y4;
  wire f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa448_y2;
  wire f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa449_y2;
  wire f_s_dadda_pg_rca32_fa462_y0;
  wire f_s_dadda_pg_rca32_fa462_y1;
  wire f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa450_y2;
  wire f_s_dadda_pg_rca32_fa462_y2;
  wire f_s_dadda_pg_rca32_fa462_y3;
  wire f_s_dadda_pg_rca32_fa462_y4;
  wire f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa451_y2;
  wire f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa452_y2;
  wire f_s_dadda_pg_rca32_fa463_y0;
  wire f_s_dadda_pg_rca32_fa463_y1;
  wire f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa453_y2;
  wire f_s_dadda_pg_rca32_fa463_y2;
  wire f_s_dadda_pg_rca32_fa463_y3;
  wire f_s_dadda_pg_rca32_fa463_y4;
  wire f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa454_y2;
  wire f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa455_y2;
  wire f_s_dadda_pg_rca32_fa464_y0;
  wire f_s_dadda_pg_rca32_fa464_y1;
  wire f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa456_y2;
  wire f_s_dadda_pg_rca32_fa464_y2;
  wire f_s_dadda_pg_rca32_fa464_y3;
  wire f_s_dadda_pg_rca32_fa464_y4;
  wire f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa457_y2;
  wire f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa458_y2;
  wire f_s_dadda_pg_rca32_fa465_y0;
  wire f_s_dadda_pg_rca32_fa465_y1;
  wire f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa459_y2;
  wire f_s_dadda_pg_rca32_fa465_y2;
  wire f_s_dadda_pg_rca32_fa465_y3;
  wire f_s_dadda_pg_rca32_fa465_y4;
  wire f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa465_y4;
  wire f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa464_y4;
  wire f_s_dadda_pg_rca32_fa466_y0;
  wire f_s_dadda_pg_rca32_fa466_y1;
  wire f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa463_y4;
  wire f_s_dadda_pg_rca32_fa466_y2;
  wire f_s_dadda_pg_rca32_fa466_y3;
  wire f_s_dadda_pg_rca32_fa466_y4;
  wire f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa462_y4;
  wire f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa461_y4;
  wire f_s_dadda_pg_rca32_fa467_y0;
  wire f_s_dadda_pg_rca32_fa467_y1;
  wire f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa460_y4;
  wire f_s_dadda_pg_rca32_fa467_y2;
  wire f_s_dadda_pg_rca32_fa467_y3;
  wire f_s_dadda_pg_rca32_fa467_y4;
  wire f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa459_y4;
  wire f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa458_y4;
  wire f_s_dadda_pg_rca32_fa468_y0;
  wire f_s_dadda_pg_rca32_fa468_y1;
  wire f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa457_y4;
  wire f_s_dadda_pg_rca32_fa468_y2;
  wire f_s_dadda_pg_rca32_fa468_y3;
  wire f_s_dadda_pg_rca32_fa468_y4;
  wire f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa456_y4;
  wire f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa455_y4;
  wire f_s_dadda_pg_rca32_fa469_y0;
  wire f_s_dadda_pg_rca32_fa469_y1;
  wire f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa454_y4;
  wire f_s_dadda_pg_rca32_fa469_y2;
  wire f_s_dadda_pg_rca32_fa469_y3;
  wire f_s_dadda_pg_rca32_fa469_y4;
  wire f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa453_y4;
  wire f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa452_y4;
  wire f_s_dadda_pg_rca32_fa470_y0;
  wire f_s_dadda_pg_rca32_fa470_y1;
  wire f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa451_y4;
  wire f_s_dadda_pg_rca32_fa470_y2;
  wire f_s_dadda_pg_rca32_fa470_y3;
  wire f_s_dadda_pg_rca32_fa470_y4;
  wire f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa450_y4;
  wire f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa449_y4;
  wire f_s_dadda_pg_rca32_fa471_y0;
  wire f_s_dadda_pg_rca32_fa471_y1;
  wire f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa448_y4;
  wire f_s_dadda_pg_rca32_fa471_y2;
  wire f_s_dadda_pg_rca32_fa471_y3;
  wire f_s_dadda_pg_rca32_fa471_y4;
  wire f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa447_y4;
  wire f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa446_y4;
  wire f_s_dadda_pg_rca32_fa472_y0;
  wire f_s_dadda_pg_rca32_fa472_y1;
  wire f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa445_y4;
  wire f_s_dadda_pg_rca32_fa472_y2;
  wire f_s_dadda_pg_rca32_fa472_y3;
  wire f_s_dadda_pg_rca32_fa472_y4;
  wire f_s_dadda_pg_rca32_nand_31_7_a_31;
  wire f_s_dadda_pg_rca32_nand_31_7_b_7;
  wire f_s_dadda_pg_rca32_nand_31_7_y0;
  wire f_s_dadda_pg_rca32_and_30_8_a_30;
  wire f_s_dadda_pg_rca32_and_30_8_b_8;
  wire f_s_dadda_pg_rca32_and_30_8_y0;
  wire f_s_dadda_pg_rca32_and_29_9_a_29;
  wire f_s_dadda_pg_rca32_and_29_9_b_9;
  wire f_s_dadda_pg_rca32_and_29_9_y0;
  wire f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_nand_31_7_y0;
  wire f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_and_30_8_y0;
  wire f_s_dadda_pg_rca32_fa473_y0;
  wire f_s_dadda_pg_rca32_fa473_y1;
  wire f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_and_29_9_y0;
  wire f_s_dadda_pg_rca32_fa473_y2;
  wire f_s_dadda_pg_rca32_fa473_y3;
  wire f_s_dadda_pg_rca32_fa473_y4;
  wire f_s_dadda_pg_rca32_and_28_10_a_28;
  wire f_s_dadda_pg_rca32_and_28_10_b_10;
  wire f_s_dadda_pg_rca32_and_28_10_y0;
  wire f_s_dadda_pg_rca32_and_27_11_a_27;
  wire f_s_dadda_pg_rca32_and_27_11_b_11;
  wire f_s_dadda_pg_rca32_and_27_11_y0;
  wire f_s_dadda_pg_rca32_and_26_12_a_26;
  wire f_s_dadda_pg_rca32_and_26_12_b_12;
  wire f_s_dadda_pg_rca32_and_26_12_y0;
  wire f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_28_10_y0;
  wire f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_27_11_y0;
  wire f_s_dadda_pg_rca32_fa474_y0;
  wire f_s_dadda_pg_rca32_fa474_y1;
  wire f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_26_12_y0;
  wire f_s_dadda_pg_rca32_fa474_y2;
  wire f_s_dadda_pg_rca32_fa474_y3;
  wire f_s_dadda_pg_rca32_fa474_y4;
  wire f_s_dadda_pg_rca32_and_25_13_a_25;
  wire f_s_dadda_pg_rca32_and_25_13_b_13;
  wire f_s_dadda_pg_rca32_and_25_13_y0;
  wire f_s_dadda_pg_rca32_and_24_14_a_24;
  wire f_s_dadda_pg_rca32_and_24_14_b_14;
  wire f_s_dadda_pg_rca32_and_24_14_y0;
  wire f_s_dadda_pg_rca32_and_23_15_a_23;
  wire f_s_dadda_pg_rca32_and_23_15_b_15;
  wire f_s_dadda_pg_rca32_and_23_15_y0;
  wire f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_25_13_y0;
  wire f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_24_14_y0;
  wire f_s_dadda_pg_rca32_fa475_y0;
  wire f_s_dadda_pg_rca32_fa475_y1;
  wire f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_23_15_y0;
  wire f_s_dadda_pg_rca32_fa475_y2;
  wire f_s_dadda_pg_rca32_fa475_y3;
  wire f_s_dadda_pg_rca32_fa475_y4;
  wire f_s_dadda_pg_rca32_and_22_16_a_22;
  wire f_s_dadda_pg_rca32_and_22_16_b_16;
  wire f_s_dadda_pg_rca32_and_22_16_y0;
  wire f_s_dadda_pg_rca32_and_21_17_a_21;
  wire f_s_dadda_pg_rca32_and_21_17_b_17;
  wire f_s_dadda_pg_rca32_and_21_17_y0;
  wire f_s_dadda_pg_rca32_and_20_18_a_20;
  wire f_s_dadda_pg_rca32_and_20_18_b_18;
  wire f_s_dadda_pg_rca32_and_20_18_y0;
  wire f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_22_16_y0;
  wire f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_21_17_y0;
  wire f_s_dadda_pg_rca32_fa476_y0;
  wire f_s_dadda_pg_rca32_fa476_y1;
  wire f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_20_18_y0;
  wire f_s_dadda_pg_rca32_fa476_y2;
  wire f_s_dadda_pg_rca32_fa476_y3;
  wire f_s_dadda_pg_rca32_fa476_y4;
  wire f_s_dadda_pg_rca32_and_19_19_a_19;
  wire f_s_dadda_pg_rca32_and_19_19_b_19;
  wire f_s_dadda_pg_rca32_and_19_19_y0;
  wire f_s_dadda_pg_rca32_and_18_20_a_18;
  wire f_s_dadda_pg_rca32_and_18_20_b_20;
  wire f_s_dadda_pg_rca32_and_18_20_y0;
  wire f_s_dadda_pg_rca32_and_17_21_a_17;
  wire f_s_dadda_pg_rca32_and_17_21_b_21;
  wire f_s_dadda_pg_rca32_and_17_21_y0;
  wire f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_19_19_y0;
  wire f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_18_20_y0;
  wire f_s_dadda_pg_rca32_fa477_y0;
  wire f_s_dadda_pg_rca32_fa477_y1;
  wire f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_17_21_y0;
  wire f_s_dadda_pg_rca32_fa477_y2;
  wire f_s_dadda_pg_rca32_fa477_y3;
  wire f_s_dadda_pg_rca32_fa477_y4;
  wire f_s_dadda_pg_rca32_and_16_22_a_16;
  wire f_s_dadda_pg_rca32_and_16_22_b_22;
  wire f_s_dadda_pg_rca32_and_16_22_y0;
  wire f_s_dadda_pg_rca32_and_15_23_a_15;
  wire f_s_dadda_pg_rca32_and_15_23_b_23;
  wire f_s_dadda_pg_rca32_and_15_23_y0;
  wire f_s_dadda_pg_rca32_and_14_24_a_14;
  wire f_s_dadda_pg_rca32_and_14_24_b_24;
  wire f_s_dadda_pg_rca32_and_14_24_y0;
  wire f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_16_22_y0;
  wire f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_15_23_y0;
  wire f_s_dadda_pg_rca32_fa478_y0;
  wire f_s_dadda_pg_rca32_fa478_y1;
  wire f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_14_24_y0;
  wire f_s_dadda_pg_rca32_fa478_y2;
  wire f_s_dadda_pg_rca32_fa478_y3;
  wire f_s_dadda_pg_rca32_fa478_y4;
  wire f_s_dadda_pg_rca32_and_13_25_a_13;
  wire f_s_dadda_pg_rca32_and_13_25_b_25;
  wire f_s_dadda_pg_rca32_and_13_25_y0;
  wire f_s_dadda_pg_rca32_and_12_26_a_12;
  wire f_s_dadda_pg_rca32_and_12_26_b_26;
  wire f_s_dadda_pg_rca32_and_12_26_y0;
  wire f_s_dadda_pg_rca32_and_11_27_a_11;
  wire f_s_dadda_pg_rca32_and_11_27_b_27;
  wire f_s_dadda_pg_rca32_and_11_27_y0;
  wire f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_13_25_y0;
  wire f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_12_26_y0;
  wire f_s_dadda_pg_rca32_fa479_y0;
  wire f_s_dadda_pg_rca32_fa479_y1;
  wire f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_11_27_y0;
  wire f_s_dadda_pg_rca32_fa479_y2;
  wire f_s_dadda_pg_rca32_fa479_y3;
  wire f_s_dadda_pg_rca32_fa479_y4;
  wire f_s_dadda_pg_rca32_and_10_28_a_10;
  wire f_s_dadda_pg_rca32_and_10_28_b_28;
  wire f_s_dadda_pg_rca32_and_10_28_y0;
  wire f_s_dadda_pg_rca32_and_9_29_a_9;
  wire f_s_dadda_pg_rca32_and_9_29_b_29;
  wire f_s_dadda_pg_rca32_and_9_29_y0;
  wire f_s_dadda_pg_rca32_and_8_30_a_8;
  wire f_s_dadda_pg_rca32_and_8_30_b_30;
  wire f_s_dadda_pg_rca32_and_8_30_y0;
  wire f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_10_28_y0;
  wire f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_9_29_y0;
  wire f_s_dadda_pg_rca32_fa480_y0;
  wire f_s_dadda_pg_rca32_fa480_y1;
  wire f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_8_30_y0;
  wire f_s_dadda_pg_rca32_fa480_y2;
  wire f_s_dadda_pg_rca32_fa480_y3;
  wire f_s_dadda_pg_rca32_fa480_y4;
  wire f_s_dadda_pg_rca32_nand_7_31_a_7;
  wire f_s_dadda_pg_rca32_nand_7_31_b_31;
  wire f_s_dadda_pg_rca32_nand_7_31_y0;
  wire f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_nand_7_31_y0;
  wire f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_fa466_y2;
  wire f_s_dadda_pg_rca32_fa481_y0;
  wire f_s_dadda_pg_rca32_fa481_y1;
  wire f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_fa467_y2;
  wire f_s_dadda_pg_rca32_fa481_y2;
  wire f_s_dadda_pg_rca32_fa481_y3;
  wire f_s_dadda_pg_rca32_fa481_y4;
  wire f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa468_y2;
  wire f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa469_y2;
  wire f_s_dadda_pg_rca32_fa482_y0;
  wire f_s_dadda_pg_rca32_fa482_y1;
  wire f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa470_y2;
  wire f_s_dadda_pg_rca32_fa482_y2;
  wire f_s_dadda_pg_rca32_fa482_y3;
  wire f_s_dadda_pg_rca32_fa482_y4;
  wire f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa471_y2;
  wire f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa472_y2;
  wire f_s_dadda_pg_rca32_fa483_y0;
  wire f_s_dadda_pg_rca32_fa483_y1;
  wire f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa473_y2;
  wire f_s_dadda_pg_rca32_fa483_y2;
  wire f_s_dadda_pg_rca32_fa483_y3;
  wire f_s_dadda_pg_rca32_fa483_y4;
  wire f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa474_y2;
  wire f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa475_y2;
  wire f_s_dadda_pg_rca32_fa484_y0;
  wire f_s_dadda_pg_rca32_fa484_y1;
  wire f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa476_y2;
  wire f_s_dadda_pg_rca32_fa484_y2;
  wire f_s_dadda_pg_rca32_fa484_y3;
  wire f_s_dadda_pg_rca32_fa484_y4;
  wire f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa477_y2;
  wire f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa478_y2;
  wire f_s_dadda_pg_rca32_fa485_y0;
  wire f_s_dadda_pg_rca32_fa485_y1;
  wire f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa479_y2;
  wire f_s_dadda_pg_rca32_fa485_y2;
  wire f_s_dadda_pg_rca32_fa485_y3;
  wire f_s_dadda_pg_rca32_fa485_y4;
  wire f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa485_y4;
  wire f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa484_y4;
  wire f_s_dadda_pg_rca32_fa486_y0;
  wire f_s_dadda_pg_rca32_fa486_y1;
  wire f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa483_y4;
  wire f_s_dadda_pg_rca32_fa486_y2;
  wire f_s_dadda_pg_rca32_fa486_y3;
  wire f_s_dadda_pg_rca32_fa486_y4;
  wire f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa482_y4;
  wire f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa481_y4;
  wire f_s_dadda_pg_rca32_fa487_y0;
  wire f_s_dadda_pg_rca32_fa487_y1;
  wire f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa480_y4;
  wire f_s_dadda_pg_rca32_fa487_y2;
  wire f_s_dadda_pg_rca32_fa487_y3;
  wire f_s_dadda_pg_rca32_fa487_y4;
  wire f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa479_y4;
  wire f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa478_y4;
  wire f_s_dadda_pg_rca32_fa488_y0;
  wire f_s_dadda_pg_rca32_fa488_y1;
  wire f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa477_y4;
  wire f_s_dadda_pg_rca32_fa488_y2;
  wire f_s_dadda_pg_rca32_fa488_y3;
  wire f_s_dadda_pg_rca32_fa488_y4;
  wire f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa476_y4;
  wire f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa475_y4;
  wire f_s_dadda_pg_rca32_fa489_y0;
  wire f_s_dadda_pg_rca32_fa489_y1;
  wire f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa474_y4;
  wire f_s_dadda_pg_rca32_fa489_y2;
  wire f_s_dadda_pg_rca32_fa489_y3;
  wire f_s_dadda_pg_rca32_fa489_y4;
  wire f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa473_y4;
  wire f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa472_y4;
  wire f_s_dadda_pg_rca32_fa490_y0;
  wire f_s_dadda_pg_rca32_fa490_y1;
  wire f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa471_y4;
  wire f_s_dadda_pg_rca32_fa490_y2;
  wire f_s_dadda_pg_rca32_fa490_y3;
  wire f_s_dadda_pg_rca32_fa490_y4;
  wire f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa470_y4;
  wire f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa469_y4;
  wire f_s_dadda_pg_rca32_fa491_y0;
  wire f_s_dadda_pg_rca32_fa491_y1;
  wire f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa468_y4;
  wire f_s_dadda_pg_rca32_fa491_y2;
  wire f_s_dadda_pg_rca32_fa491_y3;
  wire f_s_dadda_pg_rca32_fa491_y4;
  wire f_s_dadda_pg_rca32_nand_31_8_a_31;
  wire f_s_dadda_pg_rca32_nand_31_8_b_8;
  wire f_s_dadda_pg_rca32_nand_31_8_y0;
  wire f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_fa467_y4;
  wire f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_fa466_y4;
  wire f_s_dadda_pg_rca32_fa492_y0;
  wire f_s_dadda_pg_rca32_fa492_y1;
  wire f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_nand_31_8_y0;
  wire f_s_dadda_pg_rca32_fa492_y2;
  wire f_s_dadda_pg_rca32_fa492_y3;
  wire f_s_dadda_pg_rca32_fa492_y4;
  wire f_s_dadda_pg_rca32_and_30_9_a_30;
  wire f_s_dadda_pg_rca32_and_30_9_b_9;
  wire f_s_dadda_pg_rca32_and_30_9_y0;
  wire f_s_dadda_pg_rca32_and_29_10_a_29;
  wire f_s_dadda_pg_rca32_and_29_10_b_10;
  wire f_s_dadda_pg_rca32_and_29_10_y0;
  wire f_s_dadda_pg_rca32_and_28_11_a_28;
  wire f_s_dadda_pg_rca32_and_28_11_b_11;
  wire f_s_dadda_pg_rca32_and_28_11_y0;
  wire f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_30_9_y0;
  wire f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_29_10_y0;
  wire f_s_dadda_pg_rca32_fa493_y0;
  wire f_s_dadda_pg_rca32_fa493_y1;
  wire f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_28_11_y0;
  wire f_s_dadda_pg_rca32_fa493_y2;
  wire f_s_dadda_pg_rca32_fa493_y3;
  wire f_s_dadda_pg_rca32_fa493_y4;
  wire f_s_dadda_pg_rca32_and_27_12_a_27;
  wire f_s_dadda_pg_rca32_and_27_12_b_12;
  wire f_s_dadda_pg_rca32_and_27_12_y0;
  wire f_s_dadda_pg_rca32_and_26_13_a_26;
  wire f_s_dadda_pg_rca32_and_26_13_b_13;
  wire f_s_dadda_pg_rca32_and_26_13_y0;
  wire f_s_dadda_pg_rca32_and_25_14_a_25;
  wire f_s_dadda_pg_rca32_and_25_14_b_14;
  wire f_s_dadda_pg_rca32_and_25_14_y0;
  wire f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_27_12_y0;
  wire f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_26_13_y0;
  wire f_s_dadda_pg_rca32_fa494_y0;
  wire f_s_dadda_pg_rca32_fa494_y1;
  wire f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_25_14_y0;
  wire f_s_dadda_pg_rca32_fa494_y2;
  wire f_s_dadda_pg_rca32_fa494_y3;
  wire f_s_dadda_pg_rca32_fa494_y4;
  wire f_s_dadda_pg_rca32_and_24_15_a_24;
  wire f_s_dadda_pg_rca32_and_24_15_b_15;
  wire f_s_dadda_pg_rca32_and_24_15_y0;
  wire f_s_dadda_pg_rca32_and_23_16_a_23;
  wire f_s_dadda_pg_rca32_and_23_16_b_16;
  wire f_s_dadda_pg_rca32_and_23_16_y0;
  wire f_s_dadda_pg_rca32_and_22_17_a_22;
  wire f_s_dadda_pg_rca32_and_22_17_b_17;
  wire f_s_dadda_pg_rca32_and_22_17_y0;
  wire f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_24_15_y0;
  wire f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_23_16_y0;
  wire f_s_dadda_pg_rca32_fa495_y0;
  wire f_s_dadda_pg_rca32_fa495_y1;
  wire f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_22_17_y0;
  wire f_s_dadda_pg_rca32_fa495_y2;
  wire f_s_dadda_pg_rca32_fa495_y3;
  wire f_s_dadda_pg_rca32_fa495_y4;
  wire f_s_dadda_pg_rca32_and_21_18_a_21;
  wire f_s_dadda_pg_rca32_and_21_18_b_18;
  wire f_s_dadda_pg_rca32_and_21_18_y0;
  wire f_s_dadda_pg_rca32_and_20_19_a_20;
  wire f_s_dadda_pg_rca32_and_20_19_b_19;
  wire f_s_dadda_pg_rca32_and_20_19_y0;
  wire f_s_dadda_pg_rca32_and_19_20_a_19;
  wire f_s_dadda_pg_rca32_and_19_20_b_20;
  wire f_s_dadda_pg_rca32_and_19_20_y0;
  wire f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_21_18_y0;
  wire f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_20_19_y0;
  wire f_s_dadda_pg_rca32_fa496_y0;
  wire f_s_dadda_pg_rca32_fa496_y1;
  wire f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_19_20_y0;
  wire f_s_dadda_pg_rca32_fa496_y2;
  wire f_s_dadda_pg_rca32_fa496_y3;
  wire f_s_dadda_pg_rca32_fa496_y4;
  wire f_s_dadda_pg_rca32_and_18_21_a_18;
  wire f_s_dadda_pg_rca32_and_18_21_b_21;
  wire f_s_dadda_pg_rca32_and_18_21_y0;
  wire f_s_dadda_pg_rca32_and_17_22_a_17;
  wire f_s_dadda_pg_rca32_and_17_22_b_22;
  wire f_s_dadda_pg_rca32_and_17_22_y0;
  wire f_s_dadda_pg_rca32_and_16_23_a_16;
  wire f_s_dadda_pg_rca32_and_16_23_b_23;
  wire f_s_dadda_pg_rca32_and_16_23_y0;
  wire f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_18_21_y0;
  wire f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_17_22_y0;
  wire f_s_dadda_pg_rca32_fa497_y0;
  wire f_s_dadda_pg_rca32_fa497_y1;
  wire f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_16_23_y0;
  wire f_s_dadda_pg_rca32_fa497_y2;
  wire f_s_dadda_pg_rca32_fa497_y3;
  wire f_s_dadda_pg_rca32_fa497_y4;
  wire f_s_dadda_pg_rca32_and_15_24_a_15;
  wire f_s_dadda_pg_rca32_and_15_24_b_24;
  wire f_s_dadda_pg_rca32_and_15_24_y0;
  wire f_s_dadda_pg_rca32_and_14_25_a_14;
  wire f_s_dadda_pg_rca32_and_14_25_b_25;
  wire f_s_dadda_pg_rca32_and_14_25_y0;
  wire f_s_dadda_pg_rca32_and_13_26_a_13;
  wire f_s_dadda_pg_rca32_and_13_26_b_26;
  wire f_s_dadda_pg_rca32_and_13_26_y0;
  wire f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_15_24_y0;
  wire f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_14_25_y0;
  wire f_s_dadda_pg_rca32_fa498_y0;
  wire f_s_dadda_pg_rca32_fa498_y1;
  wire f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_13_26_y0;
  wire f_s_dadda_pg_rca32_fa498_y2;
  wire f_s_dadda_pg_rca32_fa498_y3;
  wire f_s_dadda_pg_rca32_fa498_y4;
  wire f_s_dadda_pg_rca32_and_12_27_a_12;
  wire f_s_dadda_pg_rca32_and_12_27_b_27;
  wire f_s_dadda_pg_rca32_and_12_27_y0;
  wire f_s_dadda_pg_rca32_and_11_28_a_11;
  wire f_s_dadda_pg_rca32_and_11_28_b_28;
  wire f_s_dadda_pg_rca32_and_11_28_y0;
  wire f_s_dadda_pg_rca32_and_10_29_a_10;
  wire f_s_dadda_pg_rca32_and_10_29_b_29;
  wire f_s_dadda_pg_rca32_and_10_29_y0;
  wire f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_12_27_y0;
  wire f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_11_28_y0;
  wire f_s_dadda_pg_rca32_fa499_y0;
  wire f_s_dadda_pg_rca32_fa499_y1;
  wire f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_10_29_y0;
  wire f_s_dadda_pg_rca32_fa499_y2;
  wire f_s_dadda_pg_rca32_fa499_y3;
  wire f_s_dadda_pg_rca32_fa499_y4;
  wire f_s_dadda_pg_rca32_and_9_30_a_9;
  wire f_s_dadda_pg_rca32_and_9_30_b_30;
  wire f_s_dadda_pg_rca32_and_9_30_y0;
  wire f_s_dadda_pg_rca32_nand_8_31_a_8;
  wire f_s_dadda_pg_rca32_nand_8_31_b_31;
  wire f_s_dadda_pg_rca32_nand_8_31_y0;
  wire f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_and_9_30_y0;
  wire f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_nand_8_31_y0;
  wire f_s_dadda_pg_rca32_fa500_y0;
  wire f_s_dadda_pg_rca32_fa500_y1;
  wire f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_fa486_y2;
  wire f_s_dadda_pg_rca32_fa500_y2;
  wire f_s_dadda_pg_rca32_fa500_y3;
  wire f_s_dadda_pg_rca32_fa500_y4;
  wire f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa487_y2;
  wire f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa488_y2;
  wire f_s_dadda_pg_rca32_fa501_y0;
  wire f_s_dadda_pg_rca32_fa501_y1;
  wire f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa489_y2;
  wire f_s_dadda_pg_rca32_fa501_y2;
  wire f_s_dadda_pg_rca32_fa501_y3;
  wire f_s_dadda_pg_rca32_fa501_y4;
  wire f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa490_y2;
  wire f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa491_y2;
  wire f_s_dadda_pg_rca32_fa502_y0;
  wire f_s_dadda_pg_rca32_fa502_y1;
  wire f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa492_y2;
  wire f_s_dadda_pg_rca32_fa502_y2;
  wire f_s_dadda_pg_rca32_fa502_y3;
  wire f_s_dadda_pg_rca32_fa502_y4;
  wire f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa493_y2;
  wire f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa494_y2;
  wire f_s_dadda_pg_rca32_fa503_y0;
  wire f_s_dadda_pg_rca32_fa503_y1;
  wire f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa495_y2;
  wire f_s_dadda_pg_rca32_fa503_y2;
  wire f_s_dadda_pg_rca32_fa503_y3;
  wire f_s_dadda_pg_rca32_fa503_y4;
  wire f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa496_y2;
  wire f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa497_y2;
  wire f_s_dadda_pg_rca32_fa504_y0;
  wire f_s_dadda_pg_rca32_fa504_y1;
  wire f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa498_y2;
  wire f_s_dadda_pg_rca32_fa504_y2;
  wire f_s_dadda_pg_rca32_fa504_y3;
  wire f_s_dadda_pg_rca32_fa504_y4;
  wire f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa504_y4;
  wire f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa503_y4;
  wire f_s_dadda_pg_rca32_fa505_y0;
  wire f_s_dadda_pg_rca32_fa505_y1;
  wire f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa502_y4;
  wire f_s_dadda_pg_rca32_fa505_y2;
  wire f_s_dadda_pg_rca32_fa505_y3;
  wire f_s_dadda_pg_rca32_fa505_y4;
  wire f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa501_y4;
  wire f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa500_y4;
  wire f_s_dadda_pg_rca32_fa506_y0;
  wire f_s_dadda_pg_rca32_fa506_y1;
  wire f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa499_y4;
  wire f_s_dadda_pg_rca32_fa506_y2;
  wire f_s_dadda_pg_rca32_fa506_y3;
  wire f_s_dadda_pg_rca32_fa506_y4;
  wire f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa498_y4;
  wire f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa497_y4;
  wire f_s_dadda_pg_rca32_fa507_y0;
  wire f_s_dadda_pg_rca32_fa507_y1;
  wire f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa496_y4;
  wire f_s_dadda_pg_rca32_fa507_y2;
  wire f_s_dadda_pg_rca32_fa507_y3;
  wire f_s_dadda_pg_rca32_fa507_y4;
  wire f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa495_y4;
  wire f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa494_y4;
  wire f_s_dadda_pg_rca32_fa508_y0;
  wire f_s_dadda_pg_rca32_fa508_y1;
  wire f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa493_y4;
  wire f_s_dadda_pg_rca32_fa508_y2;
  wire f_s_dadda_pg_rca32_fa508_y3;
  wire f_s_dadda_pg_rca32_fa508_y4;
  wire f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa492_y4;
  wire f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa491_y4;
  wire f_s_dadda_pg_rca32_fa509_y0;
  wire f_s_dadda_pg_rca32_fa509_y1;
  wire f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa490_y4;
  wire f_s_dadda_pg_rca32_fa509_y2;
  wire f_s_dadda_pg_rca32_fa509_y3;
  wire f_s_dadda_pg_rca32_fa509_y4;
  wire f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa489_y4;
  wire f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa488_y4;
  wire f_s_dadda_pg_rca32_fa510_y0;
  wire f_s_dadda_pg_rca32_fa510_y1;
  wire f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa487_y4;
  wire f_s_dadda_pg_rca32_fa510_y2;
  wire f_s_dadda_pg_rca32_fa510_y3;
  wire f_s_dadda_pg_rca32_fa510_y4;
  wire f_s_dadda_pg_rca32_nand_31_9_a_31;
  wire f_s_dadda_pg_rca32_nand_31_9_b_9;
  wire f_s_dadda_pg_rca32_nand_31_9_y0;
  wire f_s_dadda_pg_rca32_and_30_10_a_30;
  wire f_s_dadda_pg_rca32_and_30_10_b_10;
  wire f_s_dadda_pg_rca32_and_30_10_y0;
  wire f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_fa486_y4;
  wire f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_nand_31_9_y0;
  wire f_s_dadda_pg_rca32_fa511_y0;
  wire f_s_dadda_pg_rca32_fa511_y1;
  wire f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_and_30_10_y0;
  wire f_s_dadda_pg_rca32_fa511_y2;
  wire f_s_dadda_pg_rca32_fa511_y3;
  wire f_s_dadda_pg_rca32_fa511_y4;
  wire f_s_dadda_pg_rca32_and_29_11_a_29;
  wire f_s_dadda_pg_rca32_and_29_11_b_11;
  wire f_s_dadda_pg_rca32_and_29_11_y0;
  wire f_s_dadda_pg_rca32_and_28_12_a_28;
  wire f_s_dadda_pg_rca32_and_28_12_b_12;
  wire f_s_dadda_pg_rca32_and_28_12_y0;
  wire f_s_dadda_pg_rca32_and_27_13_a_27;
  wire f_s_dadda_pg_rca32_and_27_13_b_13;
  wire f_s_dadda_pg_rca32_and_27_13_y0;
  wire f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_29_11_y0;
  wire f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_28_12_y0;
  wire f_s_dadda_pg_rca32_fa512_y0;
  wire f_s_dadda_pg_rca32_fa512_y1;
  wire f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_27_13_y0;
  wire f_s_dadda_pg_rca32_fa512_y2;
  wire f_s_dadda_pg_rca32_fa512_y3;
  wire f_s_dadda_pg_rca32_fa512_y4;
  wire f_s_dadda_pg_rca32_and_26_14_a_26;
  wire f_s_dadda_pg_rca32_and_26_14_b_14;
  wire f_s_dadda_pg_rca32_and_26_14_y0;
  wire f_s_dadda_pg_rca32_and_25_15_a_25;
  wire f_s_dadda_pg_rca32_and_25_15_b_15;
  wire f_s_dadda_pg_rca32_and_25_15_y0;
  wire f_s_dadda_pg_rca32_and_24_16_a_24;
  wire f_s_dadda_pg_rca32_and_24_16_b_16;
  wire f_s_dadda_pg_rca32_and_24_16_y0;
  wire f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_26_14_y0;
  wire f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_25_15_y0;
  wire f_s_dadda_pg_rca32_fa513_y0;
  wire f_s_dadda_pg_rca32_fa513_y1;
  wire f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_24_16_y0;
  wire f_s_dadda_pg_rca32_fa513_y2;
  wire f_s_dadda_pg_rca32_fa513_y3;
  wire f_s_dadda_pg_rca32_fa513_y4;
  wire f_s_dadda_pg_rca32_and_23_17_a_23;
  wire f_s_dadda_pg_rca32_and_23_17_b_17;
  wire f_s_dadda_pg_rca32_and_23_17_y0;
  wire f_s_dadda_pg_rca32_and_22_18_a_22;
  wire f_s_dadda_pg_rca32_and_22_18_b_18;
  wire f_s_dadda_pg_rca32_and_22_18_y0;
  wire f_s_dadda_pg_rca32_and_21_19_a_21;
  wire f_s_dadda_pg_rca32_and_21_19_b_19;
  wire f_s_dadda_pg_rca32_and_21_19_y0;
  wire f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_23_17_y0;
  wire f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_22_18_y0;
  wire f_s_dadda_pg_rca32_fa514_y0;
  wire f_s_dadda_pg_rca32_fa514_y1;
  wire f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_21_19_y0;
  wire f_s_dadda_pg_rca32_fa514_y2;
  wire f_s_dadda_pg_rca32_fa514_y3;
  wire f_s_dadda_pg_rca32_fa514_y4;
  wire f_s_dadda_pg_rca32_and_20_20_a_20;
  wire f_s_dadda_pg_rca32_and_20_20_b_20;
  wire f_s_dadda_pg_rca32_and_20_20_y0;
  wire f_s_dadda_pg_rca32_and_19_21_a_19;
  wire f_s_dadda_pg_rca32_and_19_21_b_21;
  wire f_s_dadda_pg_rca32_and_19_21_y0;
  wire f_s_dadda_pg_rca32_and_18_22_a_18;
  wire f_s_dadda_pg_rca32_and_18_22_b_22;
  wire f_s_dadda_pg_rca32_and_18_22_y0;
  wire f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_20_20_y0;
  wire f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_19_21_y0;
  wire f_s_dadda_pg_rca32_fa515_y0;
  wire f_s_dadda_pg_rca32_fa515_y1;
  wire f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_18_22_y0;
  wire f_s_dadda_pg_rca32_fa515_y2;
  wire f_s_dadda_pg_rca32_fa515_y3;
  wire f_s_dadda_pg_rca32_fa515_y4;
  wire f_s_dadda_pg_rca32_and_17_23_a_17;
  wire f_s_dadda_pg_rca32_and_17_23_b_23;
  wire f_s_dadda_pg_rca32_and_17_23_y0;
  wire f_s_dadda_pg_rca32_and_16_24_a_16;
  wire f_s_dadda_pg_rca32_and_16_24_b_24;
  wire f_s_dadda_pg_rca32_and_16_24_y0;
  wire f_s_dadda_pg_rca32_and_15_25_a_15;
  wire f_s_dadda_pg_rca32_and_15_25_b_25;
  wire f_s_dadda_pg_rca32_and_15_25_y0;
  wire f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_17_23_y0;
  wire f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_16_24_y0;
  wire f_s_dadda_pg_rca32_fa516_y0;
  wire f_s_dadda_pg_rca32_fa516_y1;
  wire f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_15_25_y0;
  wire f_s_dadda_pg_rca32_fa516_y2;
  wire f_s_dadda_pg_rca32_fa516_y3;
  wire f_s_dadda_pg_rca32_fa516_y4;
  wire f_s_dadda_pg_rca32_and_14_26_a_14;
  wire f_s_dadda_pg_rca32_and_14_26_b_26;
  wire f_s_dadda_pg_rca32_and_14_26_y0;
  wire f_s_dadda_pg_rca32_and_13_27_a_13;
  wire f_s_dadda_pg_rca32_and_13_27_b_27;
  wire f_s_dadda_pg_rca32_and_13_27_y0;
  wire f_s_dadda_pg_rca32_and_12_28_a_12;
  wire f_s_dadda_pg_rca32_and_12_28_b_28;
  wire f_s_dadda_pg_rca32_and_12_28_y0;
  wire f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_14_26_y0;
  wire f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_13_27_y0;
  wire f_s_dadda_pg_rca32_fa517_y0;
  wire f_s_dadda_pg_rca32_fa517_y1;
  wire f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_12_28_y0;
  wire f_s_dadda_pg_rca32_fa517_y2;
  wire f_s_dadda_pg_rca32_fa517_y3;
  wire f_s_dadda_pg_rca32_fa517_y4;
  wire f_s_dadda_pg_rca32_and_11_29_a_11;
  wire f_s_dadda_pg_rca32_and_11_29_b_29;
  wire f_s_dadda_pg_rca32_and_11_29_y0;
  wire f_s_dadda_pg_rca32_and_10_30_a_10;
  wire f_s_dadda_pg_rca32_and_10_30_b_30;
  wire f_s_dadda_pg_rca32_and_10_30_y0;
  wire f_s_dadda_pg_rca32_nand_9_31_a_9;
  wire f_s_dadda_pg_rca32_nand_9_31_b_31;
  wire f_s_dadda_pg_rca32_nand_9_31_y0;
  wire f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_and_11_29_y0;
  wire f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_and_10_30_y0;
  wire f_s_dadda_pg_rca32_fa518_y0;
  wire f_s_dadda_pg_rca32_fa518_y1;
  wire f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_nand_9_31_y0;
  wire f_s_dadda_pg_rca32_fa518_y2;
  wire f_s_dadda_pg_rca32_fa518_y3;
  wire f_s_dadda_pg_rca32_fa518_y4;
  wire f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa505_y2;
  wire f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa506_y2;
  wire f_s_dadda_pg_rca32_fa519_y0;
  wire f_s_dadda_pg_rca32_fa519_y1;
  wire f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa507_y2;
  wire f_s_dadda_pg_rca32_fa519_y2;
  wire f_s_dadda_pg_rca32_fa519_y3;
  wire f_s_dadda_pg_rca32_fa519_y4;
  wire f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa508_y2;
  wire f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa509_y2;
  wire f_s_dadda_pg_rca32_fa520_y0;
  wire f_s_dadda_pg_rca32_fa520_y1;
  wire f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa510_y2;
  wire f_s_dadda_pg_rca32_fa520_y2;
  wire f_s_dadda_pg_rca32_fa520_y3;
  wire f_s_dadda_pg_rca32_fa520_y4;
  wire f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa511_y2;
  wire f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa512_y2;
  wire f_s_dadda_pg_rca32_fa521_y0;
  wire f_s_dadda_pg_rca32_fa521_y1;
  wire f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa513_y2;
  wire f_s_dadda_pg_rca32_fa521_y2;
  wire f_s_dadda_pg_rca32_fa521_y3;
  wire f_s_dadda_pg_rca32_fa521_y4;
  wire f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa514_y2;
  wire f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa515_y2;
  wire f_s_dadda_pg_rca32_fa522_y0;
  wire f_s_dadda_pg_rca32_fa522_y1;
  wire f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa516_y2;
  wire f_s_dadda_pg_rca32_fa522_y2;
  wire f_s_dadda_pg_rca32_fa522_y3;
  wire f_s_dadda_pg_rca32_fa522_y4;
  wire f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa522_y4;
  wire f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa521_y4;
  wire f_s_dadda_pg_rca32_fa523_y0;
  wire f_s_dadda_pg_rca32_fa523_y1;
  wire f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa520_y4;
  wire f_s_dadda_pg_rca32_fa523_y2;
  wire f_s_dadda_pg_rca32_fa523_y3;
  wire f_s_dadda_pg_rca32_fa523_y4;
  wire f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa519_y4;
  wire f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa518_y4;
  wire f_s_dadda_pg_rca32_fa524_y0;
  wire f_s_dadda_pg_rca32_fa524_y1;
  wire f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa517_y4;
  wire f_s_dadda_pg_rca32_fa524_y2;
  wire f_s_dadda_pg_rca32_fa524_y3;
  wire f_s_dadda_pg_rca32_fa524_y4;
  wire f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa516_y4;
  wire f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa515_y4;
  wire f_s_dadda_pg_rca32_fa525_y0;
  wire f_s_dadda_pg_rca32_fa525_y1;
  wire f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa514_y4;
  wire f_s_dadda_pg_rca32_fa525_y2;
  wire f_s_dadda_pg_rca32_fa525_y3;
  wire f_s_dadda_pg_rca32_fa525_y4;
  wire f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa513_y4;
  wire f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa512_y4;
  wire f_s_dadda_pg_rca32_fa526_y0;
  wire f_s_dadda_pg_rca32_fa526_y1;
  wire f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa511_y4;
  wire f_s_dadda_pg_rca32_fa526_y2;
  wire f_s_dadda_pg_rca32_fa526_y3;
  wire f_s_dadda_pg_rca32_fa526_y4;
  wire f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa510_y4;
  wire f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa509_y4;
  wire f_s_dadda_pg_rca32_fa527_y0;
  wire f_s_dadda_pg_rca32_fa527_y1;
  wire f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa508_y4;
  wire f_s_dadda_pg_rca32_fa527_y2;
  wire f_s_dadda_pg_rca32_fa527_y3;
  wire f_s_dadda_pg_rca32_fa527_y4;
  wire f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa507_y4;
  wire f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa506_y4;
  wire f_s_dadda_pg_rca32_fa528_y0;
  wire f_s_dadda_pg_rca32_fa528_y1;
  wire f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa505_y4;
  wire f_s_dadda_pg_rca32_fa528_y2;
  wire f_s_dadda_pg_rca32_fa528_y3;
  wire f_s_dadda_pg_rca32_fa528_y4;
  wire f_s_dadda_pg_rca32_nand_31_10_a_31;
  wire f_s_dadda_pg_rca32_nand_31_10_b_10;
  wire f_s_dadda_pg_rca32_nand_31_10_y0;
  wire f_s_dadda_pg_rca32_and_30_11_a_30;
  wire f_s_dadda_pg_rca32_and_30_11_b_11;
  wire f_s_dadda_pg_rca32_and_30_11_y0;
  wire f_s_dadda_pg_rca32_and_29_12_a_29;
  wire f_s_dadda_pg_rca32_and_29_12_b_12;
  wire f_s_dadda_pg_rca32_and_29_12_y0;
  wire f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_nand_31_10_y0;
  wire f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_and_30_11_y0;
  wire f_s_dadda_pg_rca32_fa529_y0;
  wire f_s_dadda_pg_rca32_fa529_y1;
  wire f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_and_29_12_y0;
  wire f_s_dadda_pg_rca32_fa529_y2;
  wire f_s_dadda_pg_rca32_fa529_y3;
  wire f_s_dadda_pg_rca32_fa529_y4;
  wire f_s_dadda_pg_rca32_and_28_13_a_28;
  wire f_s_dadda_pg_rca32_and_28_13_b_13;
  wire f_s_dadda_pg_rca32_and_28_13_y0;
  wire f_s_dadda_pg_rca32_and_27_14_a_27;
  wire f_s_dadda_pg_rca32_and_27_14_b_14;
  wire f_s_dadda_pg_rca32_and_27_14_y0;
  wire f_s_dadda_pg_rca32_and_26_15_a_26;
  wire f_s_dadda_pg_rca32_and_26_15_b_15;
  wire f_s_dadda_pg_rca32_and_26_15_y0;
  wire f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_28_13_y0;
  wire f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_27_14_y0;
  wire f_s_dadda_pg_rca32_fa530_y0;
  wire f_s_dadda_pg_rca32_fa530_y1;
  wire f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_26_15_y0;
  wire f_s_dadda_pg_rca32_fa530_y2;
  wire f_s_dadda_pg_rca32_fa530_y3;
  wire f_s_dadda_pg_rca32_fa530_y4;
  wire f_s_dadda_pg_rca32_and_25_16_a_25;
  wire f_s_dadda_pg_rca32_and_25_16_b_16;
  wire f_s_dadda_pg_rca32_and_25_16_y0;
  wire f_s_dadda_pg_rca32_and_24_17_a_24;
  wire f_s_dadda_pg_rca32_and_24_17_b_17;
  wire f_s_dadda_pg_rca32_and_24_17_y0;
  wire f_s_dadda_pg_rca32_and_23_18_a_23;
  wire f_s_dadda_pg_rca32_and_23_18_b_18;
  wire f_s_dadda_pg_rca32_and_23_18_y0;
  wire f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_25_16_y0;
  wire f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_24_17_y0;
  wire f_s_dadda_pg_rca32_fa531_y0;
  wire f_s_dadda_pg_rca32_fa531_y1;
  wire f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_23_18_y0;
  wire f_s_dadda_pg_rca32_fa531_y2;
  wire f_s_dadda_pg_rca32_fa531_y3;
  wire f_s_dadda_pg_rca32_fa531_y4;
  wire f_s_dadda_pg_rca32_and_22_19_a_22;
  wire f_s_dadda_pg_rca32_and_22_19_b_19;
  wire f_s_dadda_pg_rca32_and_22_19_y0;
  wire f_s_dadda_pg_rca32_and_21_20_a_21;
  wire f_s_dadda_pg_rca32_and_21_20_b_20;
  wire f_s_dadda_pg_rca32_and_21_20_y0;
  wire f_s_dadda_pg_rca32_and_20_21_a_20;
  wire f_s_dadda_pg_rca32_and_20_21_b_21;
  wire f_s_dadda_pg_rca32_and_20_21_y0;
  wire f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_22_19_y0;
  wire f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_21_20_y0;
  wire f_s_dadda_pg_rca32_fa532_y0;
  wire f_s_dadda_pg_rca32_fa532_y1;
  wire f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_20_21_y0;
  wire f_s_dadda_pg_rca32_fa532_y2;
  wire f_s_dadda_pg_rca32_fa532_y3;
  wire f_s_dadda_pg_rca32_fa532_y4;
  wire f_s_dadda_pg_rca32_and_19_22_a_19;
  wire f_s_dadda_pg_rca32_and_19_22_b_22;
  wire f_s_dadda_pg_rca32_and_19_22_y0;
  wire f_s_dadda_pg_rca32_and_18_23_a_18;
  wire f_s_dadda_pg_rca32_and_18_23_b_23;
  wire f_s_dadda_pg_rca32_and_18_23_y0;
  wire f_s_dadda_pg_rca32_and_17_24_a_17;
  wire f_s_dadda_pg_rca32_and_17_24_b_24;
  wire f_s_dadda_pg_rca32_and_17_24_y0;
  wire f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_19_22_y0;
  wire f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_18_23_y0;
  wire f_s_dadda_pg_rca32_fa533_y0;
  wire f_s_dadda_pg_rca32_fa533_y1;
  wire f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_17_24_y0;
  wire f_s_dadda_pg_rca32_fa533_y2;
  wire f_s_dadda_pg_rca32_fa533_y3;
  wire f_s_dadda_pg_rca32_fa533_y4;
  wire f_s_dadda_pg_rca32_and_16_25_a_16;
  wire f_s_dadda_pg_rca32_and_16_25_b_25;
  wire f_s_dadda_pg_rca32_and_16_25_y0;
  wire f_s_dadda_pg_rca32_and_15_26_a_15;
  wire f_s_dadda_pg_rca32_and_15_26_b_26;
  wire f_s_dadda_pg_rca32_and_15_26_y0;
  wire f_s_dadda_pg_rca32_and_14_27_a_14;
  wire f_s_dadda_pg_rca32_and_14_27_b_27;
  wire f_s_dadda_pg_rca32_and_14_27_y0;
  wire f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_16_25_y0;
  wire f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_15_26_y0;
  wire f_s_dadda_pg_rca32_fa534_y0;
  wire f_s_dadda_pg_rca32_fa534_y1;
  wire f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_14_27_y0;
  wire f_s_dadda_pg_rca32_fa534_y2;
  wire f_s_dadda_pg_rca32_fa534_y3;
  wire f_s_dadda_pg_rca32_fa534_y4;
  wire f_s_dadda_pg_rca32_and_13_28_a_13;
  wire f_s_dadda_pg_rca32_and_13_28_b_28;
  wire f_s_dadda_pg_rca32_and_13_28_y0;
  wire f_s_dadda_pg_rca32_and_12_29_a_12;
  wire f_s_dadda_pg_rca32_and_12_29_b_29;
  wire f_s_dadda_pg_rca32_and_12_29_y0;
  wire f_s_dadda_pg_rca32_and_11_30_a_11;
  wire f_s_dadda_pg_rca32_and_11_30_b_30;
  wire f_s_dadda_pg_rca32_and_11_30_y0;
  wire f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_13_28_y0;
  wire f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_12_29_y0;
  wire f_s_dadda_pg_rca32_fa535_y0;
  wire f_s_dadda_pg_rca32_fa535_y1;
  wire f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_11_30_y0;
  wire f_s_dadda_pg_rca32_fa535_y2;
  wire f_s_dadda_pg_rca32_fa535_y3;
  wire f_s_dadda_pg_rca32_fa535_y4;
  wire f_s_dadda_pg_rca32_nand_10_31_a_10;
  wire f_s_dadda_pg_rca32_nand_10_31_b_31;
  wire f_s_dadda_pg_rca32_nand_10_31_y0;
  wire f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_nand_10_31_y0;
  wire f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_fa523_y2;
  wire f_s_dadda_pg_rca32_fa536_y0;
  wire f_s_dadda_pg_rca32_fa536_y1;
  wire f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_fa524_y2;
  wire f_s_dadda_pg_rca32_fa536_y2;
  wire f_s_dadda_pg_rca32_fa536_y3;
  wire f_s_dadda_pg_rca32_fa536_y4;
  wire f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa525_y2;
  wire f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa526_y2;
  wire f_s_dadda_pg_rca32_fa537_y0;
  wire f_s_dadda_pg_rca32_fa537_y1;
  wire f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa527_y2;
  wire f_s_dadda_pg_rca32_fa537_y2;
  wire f_s_dadda_pg_rca32_fa537_y3;
  wire f_s_dadda_pg_rca32_fa537_y4;
  wire f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa528_y2;
  wire f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa529_y2;
  wire f_s_dadda_pg_rca32_fa538_y0;
  wire f_s_dadda_pg_rca32_fa538_y1;
  wire f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa530_y2;
  wire f_s_dadda_pg_rca32_fa538_y2;
  wire f_s_dadda_pg_rca32_fa538_y3;
  wire f_s_dadda_pg_rca32_fa538_y4;
  wire f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa531_y2;
  wire f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa532_y2;
  wire f_s_dadda_pg_rca32_fa539_y0;
  wire f_s_dadda_pg_rca32_fa539_y1;
  wire f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa533_y2;
  wire f_s_dadda_pg_rca32_fa539_y2;
  wire f_s_dadda_pg_rca32_fa539_y3;
  wire f_s_dadda_pg_rca32_fa539_y4;
  wire f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa539_y4;
  wire f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa538_y4;
  wire f_s_dadda_pg_rca32_fa540_y0;
  wire f_s_dadda_pg_rca32_fa540_y1;
  wire f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa537_y4;
  wire f_s_dadda_pg_rca32_fa540_y2;
  wire f_s_dadda_pg_rca32_fa540_y3;
  wire f_s_dadda_pg_rca32_fa540_y4;
  wire f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa536_y4;
  wire f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa535_y4;
  wire f_s_dadda_pg_rca32_fa541_y0;
  wire f_s_dadda_pg_rca32_fa541_y1;
  wire f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa534_y4;
  wire f_s_dadda_pg_rca32_fa541_y2;
  wire f_s_dadda_pg_rca32_fa541_y3;
  wire f_s_dadda_pg_rca32_fa541_y4;
  wire f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa533_y4;
  wire f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa532_y4;
  wire f_s_dadda_pg_rca32_fa542_y0;
  wire f_s_dadda_pg_rca32_fa542_y1;
  wire f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa531_y4;
  wire f_s_dadda_pg_rca32_fa542_y2;
  wire f_s_dadda_pg_rca32_fa542_y3;
  wire f_s_dadda_pg_rca32_fa542_y4;
  wire f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa530_y4;
  wire f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa529_y4;
  wire f_s_dadda_pg_rca32_fa543_y0;
  wire f_s_dadda_pg_rca32_fa543_y1;
  wire f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa528_y4;
  wire f_s_dadda_pg_rca32_fa543_y2;
  wire f_s_dadda_pg_rca32_fa543_y3;
  wire f_s_dadda_pg_rca32_fa543_y4;
  wire f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa527_y4;
  wire f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa526_y4;
  wire f_s_dadda_pg_rca32_fa544_y0;
  wire f_s_dadda_pg_rca32_fa544_y1;
  wire f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa525_y4;
  wire f_s_dadda_pg_rca32_fa544_y2;
  wire f_s_dadda_pg_rca32_fa544_y3;
  wire f_s_dadda_pg_rca32_fa544_y4;
  wire f_s_dadda_pg_rca32_nand_31_11_a_31;
  wire f_s_dadda_pg_rca32_nand_31_11_b_11;
  wire f_s_dadda_pg_rca32_nand_31_11_y0;
  wire f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_fa524_y4;
  wire f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_fa523_y4;
  wire f_s_dadda_pg_rca32_fa545_y0;
  wire f_s_dadda_pg_rca32_fa545_y1;
  wire f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_nand_31_11_y0;
  wire f_s_dadda_pg_rca32_fa545_y2;
  wire f_s_dadda_pg_rca32_fa545_y3;
  wire f_s_dadda_pg_rca32_fa545_y4;
  wire f_s_dadda_pg_rca32_and_30_12_a_30;
  wire f_s_dadda_pg_rca32_and_30_12_b_12;
  wire f_s_dadda_pg_rca32_and_30_12_y0;
  wire f_s_dadda_pg_rca32_and_29_13_a_29;
  wire f_s_dadda_pg_rca32_and_29_13_b_13;
  wire f_s_dadda_pg_rca32_and_29_13_y0;
  wire f_s_dadda_pg_rca32_and_28_14_a_28;
  wire f_s_dadda_pg_rca32_and_28_14_b_14;
  wire f_s_dadda_pg_rca32_and_28_14_y0;
  wire f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_30_12_y0;
  wire f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_29_13_y0;
  wire f_s_dadda_pg_rca32_fa546_y0;
  wire f_s_dadda_pg_rca32_fa546_y1;
  wire f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_28_14_y0;
  wire f_s_dadda_pg_rca32_fa546_y2;
  wire f_s_dadda_pg_rca32_fa546_y3;
  wire f_s_dadda_pg_rca32_fa546_y4;
  wire f_s_dadda_pg_rca32_and_27_15_a_27;
  wire f_s_dadda_pg_rca32_and_27_15_b_15;
  wire f_s_dadda_pg_rca32_and_27_15_y0;
  wire f_s_dadda_pg_rca32_and_26_16_a_26;
  wire f_s_dadda_pg_rca32_and_26_16_b_16;
  wire f_s_dadda_pg_rca32_and_26_16_y0;
  wire f_s_dadda_pg_rca32_and_25_17_a_25;
  wire f_s_dadda_pg_rca32_and_25_17_b_17;
  wire f_s_dadda_pg_rca32_and_25_17_y0;
  wire f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_27_15_y0;
  wire f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_26_16_y0;
  wire f_s_dadda_pg_rca32_fa547_y0;
  wire f_s_dadda_pg_rca32_fa547_y1;
  wire f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_25_17_y0;
  wire f_s_dadda_pg_rca32_fa547_y2;
  wire f_s_dadda_pg_rca32_fa547_y3;
  wire f_s_dadda_pg_rca32_fa547_y4;
  wire f_s_dadda_pg_rca32_and_24_18_a_24;
  wire f_s_dadda_pg_rca32_and_24_18_b_18;
  wire f_s_dadda_pg_rca32_and_24_18_y0;
  wire f_s_dadda_pg_rca32_and_23_19_a_23;
  wire f_s_dadda_pg_rca32_and_23_19_b_19;
  wire f_s_dadda_pg_rca32_and_23_19_y0;
  wire f_s_dadda_pg_rca32_and_22_20_a_22;
  wire f_s_dadda_pg_rca32_and_22_20_b_20;
  wire f_s_dadda_pg_rca32_and_22_20_y0;
  wire f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_24_18_y0;
  wire f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_23_19_y0;
  wire f_s_dadda_pg_rca32_fa548_y0;
  wire f_s_dadda_pg_rca32_fa548_y1;
  wire f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_22_20_y0;
  wire f_s_dadda_pg_rca32_fa548_y2;
  wire f_s_dadda_pg_rca32_fa548_y3;
  wire f_s_dadda_pg_rca32_fa548_y4;
  wire f_s_dadda_pg_rca32_and_21_21_a_21;
  wire f_s_dadda_pg_rca32_and_21_21_b_21;
  wire f_s_dadda_pg_rca32_and_21_21_y0;
  wire f_s_dadda_pg_rca32_and_20_22_a_20;
  wire f_s_dadda_pg_rca32_and_20_22_b_22;
  wire f_s_dadda_pg_rca32_and_20_22_y0;
  wire f_s_dadda_pg_rca32_and_19_23_a_19;
  wire f_s_dadda_pg_rca32_and_19_23_b_23;
  wire f_s_dadda_pg_rca32_and_19_23_y0;
  wire f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_21_21_y0;
  wire f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_20_22_y0;
  wire f_s_dadda_pg_rca32_fa549_y0;
  wire f_s_dadda_pg_rca32_fa549_y1;
  wire f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_19_23_y0;
  wire f_s_dadda_pg_rca32_fa549_y2;
  wire f_s_dadda_pg_rca32_fa549_y3;
  wire f_s_dadda_pg_rca32_fa549_y4;
  wire f_s_dadda_pg_rca32_and_18_24_a_18;
  wire f_s_dadda_pg_rca32_and_18_24_b_24;
  wire f_s_dadda_pg_rca32_and_18_24_y0;
  wire f_s_dadda_pg_rca32_and_17_25_a_17;
  wire f_s_dadda_pg_rca32_and_17_25_b_25;
  wire f_s_dadda_pg_rca32_and_17_25_y0;
  wire f_s_dadda_pg_rca32_and_16_26_a_16;
  wire f_s_dadda_pg_rca32_and_16_26_b_26;
  wire f_s_dadda_pg_rca32_and_16_26_y0;
  wire f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_18_24_y0;
  wire f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_17_25_y0;
  wire f_s_dadda_pg_rca32_fa550_y0;
  wire f_s_dadda_pg_rca32_fa550_y1;
  wire f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_16_26_y0;
  wire f_s_dadda_pg_rca32_fa550_y2;
  wire f_s_dadda_pg_rca32_fa550_y3;
  wire f_s_dadda_pg_rca32_fa550_y4;
  wire f_s_dadda_pg_rca32_and_15_27_a_15;
  wire f_s_dadda_pg_rca32_and_15_27_b_27;
  wire f_s_dadda_pg_rca32_and_15_27_y0;
  wire f_s_dadda_pg_rca32_and_14_28_a_14;
  wire f_s_dadda_pg_rca32_and_14_28_b_28;
  wire f_s_dadda_pg_rca32_and_14_28_y0;
  wire f_s_dadda_pg_rca32_and_13_29_a_13;
  wire f_s_dadda_pg_rca32_and_13_29_b_29;
  wire f_s_dadda_pg_rca32_and_13_29_y0;
  wire f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_15_27_y0;
  wire f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_14_28_y0;
  wire f_s_dadda_pg_rca32_fa551_y0;
  wire f_s_dadda_pg_rca32_fa551_y1;
  wire f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_13_29_y0;
  wire f_s_dadda_pg_rca32_fa551_y2;
  wire f_s_dadda_pg_rca32_fa551_y3;
  wire f_s_dadda_pg_rca32_fa551_y4;
  wire f_s_dadda_pg_rca32_and_12_30_a_12;
  wire f_s_dadda_pg_rca32_and_12_30_b_30;
  wire f_s_dadda_pg_rca32_and_12_30_y0;
  wire f_s_dadda_pg_rca32_nand_11_31_a_11;
  wire f_s_dadda_pg_rca32_nand_11_31_b_31;
  wire f_s_dadda_pg_rca32_nand_11_31_y0;
  wire f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_and_12_30_y0;
  wire f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_nand_11_31_y0;
  wire f_s_dadda_pg_rca32_fa552_y0;
  wire f_s_dadda_pg_rca32_fa552_y1;
  wire f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_fa540_y2;
  wire f_s_dadda_pg_rca32_fa552_y2;
  wire f_s_dadda_pg_rca32_fa552_y3;
  wire f_s_dadda_pg_rca32_fa552_y4;
  wire f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa541_y2;
  wire f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa542_y2;
  wire f_s_dadda_pg_rca32_fa553_y0;
  wire f_s_dadda_pg_rca32_fa553_y1;
  wire f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa543_y2;
  wire f_s_dadda_pg_rca32_fa553_y2;
  wire f_s_dadda_pg_rca32_fa553_y3;
  wire f_s_dadda_pg_rca32_fa553_y4;
  wire f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa544_y2;
  wire f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa545_y2;
  wire f_s_dadda_pg_rca32_fa554_y0;
  wire f_s_dadda_pg_rca32_fa554_y1;
  wire f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa546_y2;
  wire f_s_dadda_pg_rca32_fa554_y2;
  wire f_s_dadda_pg_rca32_fa554_y3;
  wire f_s_dadda_pg_rca32_fa554_y4;
  wire f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa547_y2;
  wire f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa548_y2;
  wire f_s_dadda_pg_rca32_fa555_y0;
  wire f_s_dadda_pg_rca32_fa555_y1;
  wire f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa549_y2;
  wire f_s_dadda_pg_rca32_fa555_y2;
  wire f_s_dadda_pg_rca32_fa555_y3;
  wire f_s_dadda_pg_rca32_fa555_y4;
  wire f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa555_y4;
  wire f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa554_y4;
  wire f_s_dadda_pg_rca32_fa556_y0;
  wire f_s_dadda_pg_rca32_fa556_y1;
  wire f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa553_y4;
  wire f_s_dadda_pg_rca32_fa556_y2;
  wire f_s_dadda_pg_rca32_fa556_y3;
  wire f_s_dadda_pg_rca32_fa556_y4;
  wire f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa552_y4;
  wire f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa551_y4;
  wire f_s_dadda_pg_rca32_fa557_y0;
  wire f_s_dadda_pg_rca32_fa557_y1;
  wire f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa550_y4;
  wire f_s_dadda_pg_rca32_fa557_y2;
  wire f_s_dadda_pg_rca32_fa557_y3;
  wire f_s_dadda_pg_rca32_fa557_y4;
  wire f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa549_y4;
  wire f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa548_y4;
  wire f_s_dadda_pg_rca32_fa558_y0;
  wire f_s_dadda_pg_rca32_fa558_y1;
  wire f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa547_y4;
  wire f_s_dadda_pg_rca32_fa558_y2;
  wire f_s_dadda_pg_rca32_fa558_y3;
  wire f_s_dadda_pg_rca32_fa558_y4;
  wire f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa546_y4;
  wire f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa545_y4;
  wire f_s_dadda_pg_rca32_fa559_y0;
  wire f_s_dadda_pg_rca32_fa559_y1;
  wire f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa544_y4;
  wire f_s_dadda_pg_rca32_fa559_y2;
  wire f_s_dadda_pg_rca32_fa559_y3;
  wire f_s_dadda_pg_rca32_fa559_y4;
  wire f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa543_y4;
  wire f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa542_y4;
  wire f_s_dadda_pg_rca32_fa560_y0;
  wire f_s_dadda_pg_rca32_fa560_y1;
  wire f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa541_y4;
  wire f_s_dadda_pg_rca32_fa560_y2;
  wire f_s_dadda_pg_rca32_fa560_y3;
  wire f_s_dadda_pg_rca32_fa560_y4;
  wire f_s_dadda_pg_rca32_nand_31_12_a_31;
  wire f_s_dadda_pg_rca32_nand_31_12_b_12;
  wire f_s_dadda_pg_rca32_nand_31_12_y0;
  wire f_s_dadda_pg_rca32_and_30_13_a_30;
  wire f_s_dadda_pg_rca32_and_30_13_b_13;
  wire f_s_dadda_pg_rca32_and_30_13_y0;
  wire f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_fa540_y4;
  wire f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_nand_31_12_y0;
  wire f_s_dadda_pg_rca32_fa561_y0;
  wire f_s_dadda_pg_rca32_fa561_y1;
  wire f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_and_30_13_y0;
  wire f_s_dadda_pg_rca32_fa561_y2;
  wire f_s_dadda_pg_rca32_fa561_y3;
  wire f_s_dadda_pg_rca32_fa561_y4;
  wire f_s_dadda_pg_rca32_and_29_14_a_29;
  wire f_s_dadda_pg_rca32_and_29_14_b_14;
  wire f_s_dadda_pg_rca32_and_29_14_y0;
  wire f_s_dadda_pg_rca32_and_28_15_a_28;
  wire f_s_dadda_pg_rca32_and_28_15_b_15;
  wire f_s_dadda_pg_rca32_and_28_15_y0;
  wire f_s_dadda_pg_rca32_and_27_16_a_27;
  wire f_s_dadda_pg_rca32_and_27_16_b_16;
  wire f_s_dadda_pg_rca32_and_27_16_y0;
  wire f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_29_14_y0;
  wire f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_28_15_y0;
  wire f_s_dadda_pg_rca32_fa562_y0;
  wire f_s_dadda_pg_rca32_fa562_y1;
  wire f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_27_16_y0;
  wire f_s_dadda_pg_rca32_fa562_y2;
  wire f_s_dadda_pg_rca32_fa562_y3;
  wire f_s_dadda_pg_rca32_fa562_y4;
  wire f_s_dadda_pg_rca32_and_26_17_a_26;
  wire f_s_dadda_pg_rca32_and_26_17_b_17;
  wire f_s_dadda_pg_rca32_and_26_17_y0;
  wire f_s_dadda_pg_rca32_and_25_18_a_25;
  wire f_s_dadda_pg_rca32_and_25_18_b_18;
  wire f_s_dadda_pg_rca32_and_25_18_y0;
  wire f_s_dadda_pg_rca32_and_24_19_a_24;
  wire f_s_dadda_pg_rca32_and_24_19_b_19;
  wire f_s_dadda_pg_rca32_and_24_19_y0;
  wire f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_26_17_y0;
  wire f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_25_18_y0;
  wire f_s_dadda_pg_rca32_fa563_y0;
  wire f_s_dadda_pg_rca32_fa563_y1;
  wire f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_24_19_y0;
  wire f_s_dadda_pg_rca32_fa563_y2;
  wire f_s_dadda_pg_rca32_fa563_y3;
  wire f_s_dadda_pg_rca32_fa563_y4;
  wire f_s_dadda_pg_rca32_and_23_20_a_23;
  wire f_s_dadda_pg_rca32_and_23_20_b_20;
  wire f_s_dadda_pg_rca32_and_23_20_y0;
  wire f_s_dadda_pg_rca32_and_22_21_a_22;
  wire f_s_dadda_pg_rca32_and_22_21_b_21;
  wire f_s_dadda_pg_rca32_and_22_21_y0;
  wire f_s_dadda_pg_rca32_and_21_22_a_21;
  wire f_s_dadda_pg_rca32_and_21_22_b_22;
  wire f_s_dadda_pg_rca32_and_21_22_y0;
  wire f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_23_20_y0;
  wire f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_22_21_y0;
  wire f_s_dadda_pg_rca32_fa564_y0;
  wire f_s_dadda_pg_rca32_fa564_y1;
  wire f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_21_22_y0;
  wire f_s_dadda_pg_rca32_fa564_y2;
  wire f_s_dadda_pg_rca32_fa564_y3;
  wire f_s_dadda_pg_rca32_fa564_y4;
  wire f_s_dadda_pg_rca32_and_20_23_a_20;
  wire f_s_dadda_pg_rca32_and_20_23_b_23;
  wire f_s_dadda_pg_rca32_and_20_23_y0;
  wire f_s_dadda_pg_rca32_and_19_24_a_19;
  wire f_s_dadda_pg_rca32_and_19_24_b_24;
  wire f_s_dadda_pg_rca32_and_19_24_y0;
  wire f_s_dadda_pg_rca32_and_18_25_a_18;
  wire f_s_dadda_pg_rca32_and_18_25_b_25;
  wire f_s_dadda_pg_rca32_and_18_25_y0;
  wire f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_20_23_y0;
  wire f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_19_24_y0;
  wire f_s_dadda_pg_rca32_fa565_y0;
  wire f_s_dadda_pg_rca32_fa565_y1;
  wire f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_18_25_y0;
  wire f_s_dadda_pg_rca32_fa565_y2;
  wire f_s_dadda_pg_rca32_fa565_y3;
  wire f_s_dadda_pg_rca32_fa565_y4;
  wire f_s_dadda_pg_rca32_and_17_26_a_17;
  wire f_s_dadda_pg_rca32_and_17_26_b_26;
  wire f_s_dadda_pg_rca32_and_17_26_y0;
  wire f_s_dadda_pg_rca32_and_16_27_a_16;
  wire f_s_dadda_pg_rca32_and_16_27_b_27;
  wire f_s_dadda_pg_rca32_and_16_27_y0;
  wire f_s_dadda_pg_rca32_and_15_28_a_15;
  wire f_s_dadda_pg_rca32_and_15_28_b_28;
  wire f_s_dadda_pg_rca32_and_15_28_y0;
  wire f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_17_26_y0;
  wire f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_16_27_y0;
  wire f_s_dadda_pg_rca32_fa566_y0;
  wire f_s_dadda_pg_rca32_fa566_y1;
  wire f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_15_28_y0;
  wire f_s_dadda_pg_rca32_fa566_y2;
  wire f_s_dadda_pg_rca32_fa566_y3;
  wire f_s_dadda_pg_rca32_fa566_y4;
  wire f_s_dadda_pg_rca32_and_14_29_a_14;
  wire f_s_dadda_pg_rca32_and_14_29_b_29;
  wire f_s_dadda_pg_rca32_and_14_29_y0;
  wire f_s_dadda_pg_rca32_and_13_30_a_13;
  wire f_s_dadda_pg_rca32_and_13_30_b_30;
  wire f_s_dadda_pg_rca32_and_13_30_y0;
  wire f_s_dadda_pg_rca32_nand_12_31_a_12;
  wire f_s_dadda_pg_rca32_nand_12_31_b_31;
  wire f_s_dadda_pg_rca32_nand_12_31_y0;
  wire f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_and_14_29_y0;
  wire f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_and_13_30_y0;
  wire f_s_dadda_pg_rca32_fa567_y0;
  wire f_s_dadda_pg_rca32_fa567_y1;
  wire f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_nand_12_31_y0;
  wire f_s_dadda_pg_rca32_fa567_y2;
  wire f_s_dadda_pg_rca32_fa567_y3;
  wire f_s_dadda_pg_rca32_fa567_y4;
  wire f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa556_y2;
  wire f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa557_y2;
  wire f_s_dadda_pg_rca32_fa568_y0;
  wire f_s_dadda_pg_rca32_fa568_y1;
  wire f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa558_y2;
  wire f_s_dadda_pg_rca32_fa568_y2;
  wire f_s_dadda_pg_rca32_fa568_y3;
  wire f_s_dadda_pg_rca32_fa568_y4;
  wire f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa559_y2;
  wire f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa560_y2;
  wire f_s_dadda_pg_rca32_fa569_y0;
  wire f_s_dadda_pg_rca32_fa569_y1;
  wire f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa561_y2;
  wire f_s_dadda_pg_rca32_fa569_y2;
  wire f_s_dadda_pg_rca32_fa569_y3;
  wire f_s_dadda_pg_rca32_fa569_y4;
  wire f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa562_y2;
  wire f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa563_y2;
  wire f_s_dadda_pg_rca32_fa570_y0;
  wire f_s_dadda_pg_rca32_fa570_y1;
  wire f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa564_y2;
  wire f_s_dadda_pg_rca32_fa570_y2;
  wire f_s_dadda_pg_rca32_fa570_y3;
  wire f_s_dadda_pg_rca32_fa570_y4;
  wire f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa570_y4;
  wire f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa569_y4;
  wire f_s_dadda_pg_rca32_fa571_y0;
  wire f_s_dadda_pg_rca32_fa571_y1;
  wire f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa568_y4;
  wire f_s_dadda_pg_rca32_fa571_y2;
  wire f_s_dadda_pg_rca32_fa571_y3;
  wire f_s_dadda_pg_rca32_fa571_y4;
  wire f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa567_y4;
  wire f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa566_y4;
  wire f_s_dadda_pg_rca32_fa572_y0;
  wire f_s_dadda_pg_rca32_fa572_y1;
  wire f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa565_y4;
  wire f_s_dadda_pg_rca32_fa572_y2;
  wire f_s_dadda_pg_rca32_fa572_y3;
  wire f_s_dadda_pg_rca32_fa572_y4;
  wire f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa564_y4;
  wire f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa563_y4;
  wire f_s_dadda_pg_rca32_fa573_y0;
  wire f_s_dadda_pg_rca32_fa573_y1;
  wire f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa562_y4;
  wire f_s_dadda_pg_rca32_fa573_y2;
  wire f_s_dadda_pg_rca32_fa573_y3;
  wire f_s_dadda_pg_rca32_fa573_y4;
  wire f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa561_y4;
  wire f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa560_y4;
  wire f_s_dadda_pg_rca32_fa574_y0;
  wire f_s_dadda_pg_rca32_fa574_y1;
  wire f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa559_y4;
  wire f_s_dadda_pg_rca32_fa574_y2;
  wire f_s_dadda_pg_rca32_fa574_y3;
  wire f_s_dadda_pg_rca32_fa574_y4;
  wire f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa558_y4;
  wire f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa557_y4;
  wire f_s_dadda_pg_rca32_fa575_y0;
  wire f_s_dadda_pg_rca32_fa575_y1;
  wire f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa556_y4;
  wire f_s_dadda_pg_rca32_fa575_y2;
  wire f_s_dadda_pg_rca32_fa575_y3;
  wire f_s_dadda_pg_rca32_fa575_y4;
  wire f_s_dadda_pg_rca32_nand_31_13_a_31;
  wire f_s_dadda_pg_rca32_nand_31_13_b_13;
  wire f_s_dadda_pg_rca32_nand_31_13_y0;
  wire f_s_dadda_pg_rca32_and_30_14_a_30;
  wire f_s_dadda_pg_rca32_and_30_14_b_14;
  wire f_s_dadda_pg_rca32_and_30_14_y0;
  wire f_s_dadda_pg_rca32_and_29_15_a_29;
  wire f_s_dadda_pg_rca32_and_29_15_b_15;
  wire f_s_dadda_pg_rca32_and_29_15_y0;
  wire f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_nand_31_13_y0;
  wire f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_and_30_14_y0;
  wire f_s_dadda_pg_rca32_fa576_y0;
  wire f_s_dadda_pg_rca32_fa576_y1;
  wire f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_and_29_15_y0;
  wire f_s_dadda_pg_rca32_fa576_y2;
  wire f_s_dadda_pg_rca32_fa576_y3;
  wire f_s_dadda_pg_rca32_fa576_y4;
  wire f_s_dadda_pg_rca32_and_28_16_a_28;
  wire f_s_dadda_pg_rca32_and_28_16_b_16;
  wire f_s_dadda_pg_rca32_and_28_16_y0;
  wire f_s_dadda_pg_rca32_and_27_17_a_27;
  wire f_s_dadda_pg_rca32_and_27_17_b_17;
  wire f_s_dadda_pg_rca32_and_27_17_y0;
  wire f_s_dadda_pg_rca32_and_26_18_a_26;
  wire f_s_dadda_pg_rca32_and_26_18_b_18;
  wire f_s_dadda_pg_rca32_and_26_18_y0;
  wire f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_28_16_y0;
  wire f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_27_17_y0;
  wire f_s_dadda_pg_rca32_fa577_y0;
  wire f_s_dadda_pg_rca32_fa577_y1;
  wire f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_26_18_y0;
  wire f_s_dadda_pg_rca32_fa577_y2;
  wire f_s_dadda_pg_rca32_fa577_y3;
  wire f_s_dadda_pg_rca32_fa577_y4;
  wire f_s_dadda_pg_rca32_and_25_19_a_25;
  wire f_s_dadda_pg_rca32_and_25_19_b_19;
  wire f_s_dadda_pg_rca32_and_25_19_y0;
  wire f_s_dadda_pg_rca32_and_24_20_a_24;
  wire f_s_dadda_pg_rca32_and_24_20_b_20;
  wire f_s_dadda_pg_rca32_and_24_20_y0;
  wire f_s_dadda_pg_rca32_and_23_21_a_23;
  wire f_s_dadda_pg_rca32_and_23_21_b_21;
  wire f_s_dadda_pg_rca32_and_23_21_y0;
  wire f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_25_19_y0;
  wire f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_24_20_y0;
  wire f_s_dadda_pg_rca32_fa578_y0;
  wire f_s_dadda_pg_rca32_fa578_y1;
  wire f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_23_21_y0;
  wire f_s_dadda_pg_rca32_fa578_y2;
  wire f_s_dadda_pg_rca32_fa578_y3;
  wire f_s_dadda_pg_rca32_fa578_y4;
  wire f_s_dadda_pg_rca32_and_22_22_a_22;
  wire f_s_dadda_pg_rca32_and_22_22_b_22;
  wire f_s_dadda_pg_rca32_and_22_22_y0;
  wire f_s_dadda_pg_rca32_and_21_23_a_21;
  wire f_s_dadda_pg_rca32_and_21_23_b_23;
  wire f_s_dadda_pg_rca32_and_21_23_y0;
  wire f_s_dadda_pg_rca32_and_20_24_a_20;
  wire f_s_dadda_pg_rca32_and_20_24_b_24;
  wire f_s_dadda_pg_rca32_and_20_24_y0;
  wire f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_22_22_y0;
  wire f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_21_23_y0;
  wire f_s_dadda_pg_rca32_fa579_y0;
  wire f_s_dadda_pg_rca32_fa579_y1;
  wire f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_20_24_y0;
  wire f_s_dadda_pg_rca32_fa579_y2;
  wire f_s_dadda_pg_rca32_fa579_y3;
  wire f_s_dadda_pg_rca32_fa579_y4;
  wire f_s_dadda_pg_rca32_and_19_25_a_19;
  wire f_s_dadda_pg_rca32_and_19_25_b_25;
  wire f_s_dadda_pg_rca32_and_19_25_y0;
  wire f_s_dadda_pg_rca32_and_18_26_a_18;
  wire f_s_dadda_pg_rca32_and_18_26_b_26;
  wire f_s_dadda_pg_rca32_and_18_26_y0;
  wire f_s_dadda_pg_rca32_and_17_27_a_17;
  wire f_s_dadda_pg_rca32_and_17_27_b_27;
  wire f_s_dadda_pg_rca32_and_17_27_y0;
  wire f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_19_25_y0;
  wire f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_18_26_y0;
  wire f_s_dadda_pg_rca32_fa580_y0;
  wire f_s_dadda_pg_rca32_fa580_y1;
  wire f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_17_27_y0;
  wire f_s_dadda_pg_rca32_fa580_y2;
  wire f_s_dadda_pg_rca32_fa580_y3;
  wire f_s_dadda_pg_rca32_fa580_y4;
  wire f_s_dadda_pg_rca32_and_16_28_a_16;
  wire f_s_dadda_pg_rca32_and_16_28_b_28;
  wire f_s_dadda_pg_rca32_and_16_28_y0;
  wire f_s_dadda_pg_rca32_and_15_29_a_15;
  wire f_s_dadda_pg_rca32_and_15_29_b_29;
  wire f_s_dadda_pg_rca32_and_15_29_y0;
  wire f_s_dadda_pg_rca32_and_14_30_a_14;
  wire f_s_dadda_pg_rca32_and_14_30_b_30;
  wire f_s_dadda_pg_rca32_and_14_30_y0;
  wire f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_16_28_y0;
  wire f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_15_29_y0;
  wire f_s_dadda_pg_rca32_fa581_y0;
  wire f_s_dadda_pg_rca32_fa581_y1;
  wire f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_14_30_y0;
  wire f_s_dadda_pg_rca32_fa581_y2;
  wire f_s_dadda_pg_rca32_fa581_y3;
  wire f_s_dadda_pg_rca32_fa581_y4;
  wire f_s_dadda_pg_rca32_nand_13_31_a_13;
  wire f_s_dadda_pg_rca32_nand_13_31_b_31;
  wire f_s_dadda_pg_rca32_nand_13_31_y0;
  wire f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_nand_13_31_y0;
  wire f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_fa571_y2;
  wire f_s_dadda_pg_rca32_fa582_y0;
  wire f_s_dadda_pg_rca32_fa582_y1;
  wire f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_fa572_y2;
  wire f_s_dadda_pg_rca32_fa582_y2;
  wire f_s_dadda_pg_rca32_fa582_y3;
  wire f_s_dadda_pg_rca32_fa582_y4;
  wire f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa573_y2;
  wire f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa574_y2;
  wire f_s_dadda_pg_rca32_fa583_y0;
  wire f_s_dadda_pg_rca32_fa583_y1;
  wire f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa575_y2;
  wire f_s_dadda_pg_rca32_fa583_y2;
  wire f_s_dadda_pg_rca32_fa583_y3;
  wire f_s_dadda_pg_rca32_fa583_y4;
  wire f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa576_y2;
  wire f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa577_y2;
  wire f_s_dadda_pg_rca32_fa584_y0;
  wire f_s_dadda_pg_rca32_fa584_y1;
  wire f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa578_y2;
  wire f_s_dadda_pg_rca32_fa584_y2;
  wire f_s_dadda_pg_rca32_fa584_y3;
  wire f_s_dadda_pg_rca32_fa584_y4;
  wire f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa584_y4;
  wire f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa583_y4;
  wire f_s_dadda_pg_rca32_fa585_y0;
  wire f_s_dadda_pg_rca32_fa585_y1;
  wire f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa582_y4;
  wire f_s_dadda_pg_rca32_fa585_y2;
  wire f_s_dadda_pg_rca32_fa585_y3;
  wire f_s_dadda_pg_rca32_fa585_y4;
  wire f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa581_y4;
  wire f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa580_y4;
  wire f_s_dadda_pg_rca32_fa586_y0;
  wire f_s_dadda_pg_rca32_fa586_y1;
  wire f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa579_y4;
  wire f_s_dadda_pg_rca32_fa586_y2;
  wire f_s_dadda_pg_rca32_fa586_y3;
  wire f_s_dadda_pg_rca32_fa586_y4;
  wire f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa578_y4;
  wire f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa577_y4;
  wire f_s_dadda_pg_rca32_fa587_y0;
  wire f_s_dadda_pg_rca32_fa587_y1;
  wire f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa576_y4;
  wire f_s_dadda_pg_rca32_fa587_y2;
  wire f_s_dadda_pg_rca32_fa587_y3;
  wire f_s_dadda_pg_rca32_fa587_y4;
  wire f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa575_y4;
  wire f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa574_y4;
  wire f_s_dadda_pg_rca32_fa588_y0;
  wire f_s_dadda_pg_rca32_fa588_y1;
  wire f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa573_y4;
  wire f_s_dadda_pg_rca32_fa588_y2;
  wire f_s_dadda_pg_rca32_fa588_y3;
  wire f_s_dadda_pg_rca32_fa588_y4;
  wire f_s_dadda_pg_rca32_nand_31_14_a_31;
  wire f_s_dadda_pg_rca32_nand_31_14_b_14;
  wire f_s_dadda_pg_rca32_nand_31_14_y0;
  wire f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_fa572_y4;
  wire f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_fa571_y4;
  wire f_s_dadda_pg_rca32_fa589_y0;
  wire f_s_dadda_pg_rca32_fa589_y1;
  wire f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_nand_31_14_y0;
  wire f_s_dadda_pg_rca32_fa589_y2;
  wire f_s_dadda_pg_rca32_fa589_y3;
  wire f_s_dadda_pg_rca32_fa589_y4;
  wire f_s_dadda_pg_rca32_and_30_15_a_30;
  wire f_s_dadda_pg_rca32_and_30_15_b_15;
  wire f_s_dadda_pg_rca32_and_30_15_y0;
  wire f_s_dadda_pg_rca32_and_29_16_a_29;
  wire f_s_dadda_pg_rca32_and_29_16_b_16;
  wire f_s_dadda_pg_rca32_and_29_16_y0;
  wire f_s_dadda_pg_rca32_and_28_17_a_28;
  wire f_s_dadda_pg_rca32_and_28_17_b_17;
  wire f_s_dadda_pg_rca32_and_28_17_y0;
  wire f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_30_15_y0;
  wire f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_29_16_y0;
  wire f_s_dadda_pg_rca32_fa590_y0;
  wire f_s_dadda_pg_rca32_fa590_y1;
  wire f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_28_17_y0;
  wire f_s_dadda_pg_rca32_fa590_y2;
  wire f_s_dadda_pg_rca32_fa590_y3;
  wire f_s_dadda_pg_rca32_fa590_y4;
  wire f_s_dadda_pg_rca32_and_27_18_a_27;
  wire f_s_dadda_pg_rca32_and_27_18_b_18;
  wire f_s_dadda_pg_rca32_and_27_18_y0;
  wire f_s_dadda_pg_rca32_and_26_19_a_26;
  wire f_s_dadda_pg_rca32_and_26_19_b_19;
  wire f_s_dadda_pg_rca32_and_26_19_y0;
  wire f_s_dadda_pg_rca32_and_25_20_a_25;
  wire f_s_dadda_pg_rca32_and_25_20_b_20;
  wire f_s_dadda_pg_rca32_and_25_20_y0;
  wire f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_27_18_y0;
  wire f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_26_19_y0;
  wire f_s_dadda_pg_rca32_fa591_y0;
  wire f_s_dadda_pg_rca32_fa591_y1;
  wire f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_25_20_y0;
  wire f_s_dadda_pg_rca32_fa591_y2;
  wire f_s_dadda_pg_rca32_fa591_y3;
  wire f_s_dadda_pg_rca32_fa591_y4;
  wire f_s_dadda_pg_rca32_and_24_21_a_24;
  wire f_s_dadda_pg_rca32_and_24_21_b_21;
  wire f_s_dadda_pg_rca32_and_24_21_y0;
  wire f_s_dadda_pg_rca32_and_23_22_a_23;
  wire f_s_dadda_pg_rca32_and_23_22_b_22;
  wire f_s_dadda_pg_rca32_and_23_22_y0;
  wire f_s_dadda_pg_rca32_and_22_23_a_22;
  wire f_s_dadda_pg_rca32_and_22_23_b_23;
  wire f_s_dadda_pg_rca32_and_22_23_y0;
  wire f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_24_21_y0;
  wire f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_23_22_y0;
  wire f_s_dadda_pg_rca32_fa592_y0;
  wire f_s_dadda_pg_rca32_fa592_y1;
  wire f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_22_23_y0;
  wire f_s_dadda_pg_rca32_fa592_y2;
  wire f_s_dadda_pg_rca32_fa592_y3;
  wire f_s_dadda_pg_rca32_fa592_y4;
  wire f_s_dadda_pg_rca32_and_21_24_a_21;
  wire f_s_dadda_pg_rca32_and_21_24_b_24;
  wire f_s_dadda_pg_rca32_and_21_24_y0;
  wire f_s_dadda_pg_rca32_and_20_25_a_20;
  wire f_s_dadda_pg_rca32_and_20_25_b_25;
  wire f_s_dadda_pg_rca32_and_20_25_y0;
  wire f_s_dadda_pg_rca32_and_19_26_a_19;
  wire f_s_dadda_pg_rca32_and_19_26_b_26;
  wire f_s_dadda_pg_rca32_and_19_26_y0;
  wire f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_21_24_y0;
  wire f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_20_25_y0;
  wire f_s_dadda_pg_rca32_fa593_y0;
  wire f_s_dadda_pg_rca32_fa593_y1;
  wire f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_19_26_y0;
  wire f_s_dadda_pg_rca32_fa593_y2;
  wire f_s_dadda_pg_rca32_fa593_y3;
  wire f_s_dadda_pg_rca32_fa593_y4;
  wire f_s_dadda_pg_rca32_and_18_27_a_18;
  wire f_s_dadda_pg_rca32_and_18_27_b_27;
  wire f_s_dadda_pg_rca32_and_18_27_y0;
  wire f_s_dadda_pg_rca32_and_17_28_a_17;
  wire f_s_dadda_pg_rca32_and_17_28_b_28;
  wire f_s_dadda_pg_rca32_and_17_28_y0;
  wire f_s_dadda_pg_rca32_and_16_29_a_16;
  wire f_s_dadda_pg_rca32_and_16_29_b_29;
  wire f_s_dadda_pg_rca32_and_16_29_y0;
  wire f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_18_27_y0;
  wire f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_17_28_y0;
  wire f_s_dadda_pg_rca32_fa594_y0;
  wire f_s_dadda_pg_rca32_fa594_y1;
  wire f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_16_29_y0;
  wire f_s_dadda_pg_rca32_fa594_y2;
  wire f_s_dadda_pg_rca32_fa594_y3;
  wire f_s_dadda_pg_rca32_fa594_y4;
  wire f_s_dadda_pg_rca32_and_15_30_a_15;
  wire f_s_dadda_pg_rca32_and_15_30_b_30;
  wire f_s_dadda_pg_rca32_and_15_30_y0;
  wire f_s_dadda_pg_rca32_nand_14_31_a_14;
  wire f_s_dadda_pg_rca32_nand_14_31_b_31;
  wire f_s_dadda_pg_rca32_nand_14_31_y0;
  wire f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_and_15_30_y0;
  wire f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_nand_14_31_y0;
  wire f_s_dadda_pg_rca32_fa595_y0;
  wire f_s_dadda_pg_rca32_fa595_y1;
  wire f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_fa585_y2;
  wire f_s_dadda_pg_rca32_fa595_y2;
  wire f_s_dadda_pg_rca32_fa595_y3;
  wire f_s_dadda_pg_rca32_fa595_y4;
  wire f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa586_y2;
  wire f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa587_y2;
  wire f_s_dadda_pg_rca32_fa596_y0;
  wire f_s_dadda_pg_rca32_fa596_y1;
  wire f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa588_y2;
  wire f_s_dadda_pg_rca32_fa596_y2;
  wire f_s_dadda_pg_rca32_fa596_y3;
  wire f_s_dadda_pg_rca32_fa596_y4;
  wire f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa589_y2;
  wire f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa590_y2;
  wire f_s_dadda_pg_rca32_fa597_y0;
  wire f_s_dadda_pg_rca32_fa597_y1;
  wire f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa591_y2;
  wire f_s_dadda_pg_rca32_fa597_y2;
  wire f_s_dadda_pg_rca32_fa597_y3;
  wire f_s_dadda_pg_rca32_fa597_y4;
  wire f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa597_y4;
  wire f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa596_y4;
  wire f_s_dadda_pg_rca32_fa598_y0;
  wire f_s_dadda_pg_rca32_fa598_y1;
  wire f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa595_y4;
  wire f_s_dadda_pg_rca32_fa598_y2;
  wire f_s_dadda_pg_rca32_fa598_y3;
  wire f_s_dadda_pg_rca32_fa598_y4;
  wire f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa594_y4;
  wire f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa593_y4;
  wire f_s_dadda_pg_rca32_fa599_y0;
  wire f_s_dadda_pg_rca32_fa599_y1;
  wire f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa592_y4;
  wire f_s_dadda_pg_rca32_fa599_y2;
  wire f_s_dadda_pg_rca32_fa599_y3;
  wire f_s_dadda_pg_rca32_fa599_y4;
  wire f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa591_y4;
  wire f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa590_y4;
  wire f_s_dadda_pg_rca32_fa600_y0;
  wire f_s_dadda_pg_rca32_fa600_y1;
  wire f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa589_y4;
  wire f_s_dadda_pg_rca32_fa600_y2;
  wire f_s_dadda_pg_rca32_fa600_y3;
  wire f_s_dadda_pg_rca32_fa600_y4;
  wire f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa588_y4;
  wire f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa587_y4;
  wire f_s_dadda_pg_rca32_fa601_y0;
  wire f_s_dadda_pg_rca32_fa601_y1;
  wire f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa586_y4;
  wire f_s_dadda_pg_rca32_fa601_y2;
  wire f_s_dadda_pg_rca32_fa601_y3;
  wire f_s_dadda_pg_rca32_fa601_y4;
  wire f_s_dadda_pg_rca32_nand_31_15_a_31;
  wire f_s_dadda_pg_rca32_nand_31_15_b_15;
  wire f_s_dadda_pg_rca32_nand_31_15_y0;
  wire f_s_dadda_pg_rca32_and_30_16_a_30;
  wire f_s_dadda_pg_rca32_and_30_16_b_16;
  wire f_s_dadda_pg_rca32_and_30_16_y0;
  wire f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_fa585_y4;
  wire f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_nand_31_15_y0;
  wire f_s_dadda_pg_rca32_fa602_y0;
  wire f_s_dadda_pg_rca32_fa602_y1;
  wire f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_and_30_16_y0;
  wire f_s_dadda_pg_rca32_fa602_y2;
  wire f_s_dadda_pg_rca32_fa602_y3;
  wire f_s_dadda_pg_rca32_fa602_y4;
  wire f_s_dadda_pg_rca32_and_29_17_a_29;
  wire f_s_dadda_pg_rca32_and_29_17_b_17;
  wire f_s_dadda_pg_rca32_and_29_17_y0;
  wire f_s_dadda_pg_rca32_and_28_18_a_28;
  wire f_s_dadda_pg_rca32_and_28_18_b_18;
  wire f_s_dadda_pg_rca32_and_28_18_y0;
  wire f_s_dadda_pg_rca32_and_27_19_a_27;
  wire f_s_dadda_pg_rca32_and_27_19_b_19;
  wire f_s_dadda_pg_rca32_and_27_19_y0;
  wire f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_29_17_y0;
  wire f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_28_18_y0;
  wire f_s_dadda_pg_rca32_fa603_y0;
  wire f_s_dadda_pg_rca32_fa603_y1;
  wire f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_27_19_y0;
  wire f_s_dadda_pg_rca32_fa603_y2;
  wire f_s_dadda_pg_rca32_fa603_y3;
  wire f_s_dadda_pg_rca32_fa603_y4;
  wire f_s_dadda_pg_rca32_and_26_20_a_26;
  wire f_s_dadda_pg_rca32_and_26_20_b_20;
  wire f_s_dadda_pg_rca32_and_26_20_y0;
  wire f_s_dadda_pg_rca32_and_25_21_a_25;
  wire f_s_dadda_pg_rca32_and_25_21_b_21;
  wire f_s_dadda_pg_rca32_and_25_21_y0;
  wire f_s_dadda_pg_rca32_and_24_22_a_24;
  wire f_s_dadda_pg_rca32_and_24_22_b_22;
  wire f_s_dadda_pg_rca32_and_24_22_y0;
  wire f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_26_20_y0;
  wire f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_25_21_y0;
  wire f_s_dadda_pg_rca32_fa604_y0;
  wire f_s_dadda_pg_rca32_fa604_y1;
  wire f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_24_22_y0;
  wire f_s_dadda_pg_rca32_fa604_y2;
  wire f_s_dadda_pg_rca32_fa604_y3;
  wire f_s_dadda_pg_rca32_fa604_y4;
  wire f_s_dadda_pg_rca32_and_23_23_a_23;
  wire f_s_dadda_pg_rca32_and_23_23_b_23;
  wire f_s_dadda_pg_rca32_and_23_23_y0;
  wire f_s_dadda_pg_rca32_and_22_24_a_22;
  wire f_s_dadda_pg_rca32_and_22_24_b_24;
  wire f_s_dadda_pg_rca32_and_22_24_y0;
  wire f_s_dadda_pg_rca32_and_21_25_a_21;
  wire f_s_dadda_pg_rca32_and_21_25_b_25;
  wire f_s_dadda_pg_rca32_and_21_25_y0;
  wire f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_23_23_y0;
  wire f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_22_24_y0;
  wire f_s_dadda_pg_rca32_fa605_y0;
  wire f_s_dadda_pg_rca32_fa605_y1;
  wire f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_21_25_y0;
  wire f_s_dadda_pg_rca32_fa605_y2;
  wire f_s_dadda_pg_rca32_fa605_y3;
  wire f_s_dadda_pg_rca32_fa605_y4;
  wire f_s_dadda_pg_rca32_and_20_26_a_20;
  wire f_s_dadda_pg_rca32_and_20_26_b_26;
  wire f_s_dadda_pg_rca32_and_20_26_y0;
  wire f_s_dadda_pg_rca32_and_19_27_a_19;
  wire f_s_dadda_pg_rca32_and_19_27_b_27;
  wire f_s_dadda_pg_rca32_and_19_27_y0;
  wire f_s_dadda_pg_rca32_and_18_28_a_18;
  wire f_s_dadda_pg_rca32_and_18_28_b_28;
  wire f_s_dadda_pg_rca32_and_18_28_y0;
  wire f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_20_26_y0;
  wire f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_19_27_y0;
  wire f_s_dadda_pg_rca32_fa606_y0;
  wire f_s_dadda_pg_rca32_fa606_y1;
  wire f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_18_28_y0;
  wire f_s_dadda_pg_rca32_fa606_y2;
  wire f_s_dadda_pg_rca32_fa606_y3;
  wire f_s_dadda_pg_rca32_fa606_y4;
  wire f_s_dadda_pg_rca32_and_17_29_a_17;
  wire f_s_dadda_pg_rca32_and_17_29_b_29;
  wire f_s_dadda_pg_rca32_and_17_29_y0;
  wire f_s_dadda_pg_rca32_and_16_30_a_16;
  wire f_s_dadda_pg_rca32_and_16_30_b_30;
  wire f_s_dadda_pg_rca32_and_16_30_y0;
  wire f_s_dadda_pg_rca32_nand_15_31_a_15;
  wire f_s_dadda_pg_rca32_nand_15_31_b_31;
  wire f_s_dadda_pg_rca32_nand_15_31_y0;
  wire f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_and_17_29_y0;
  wire f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_and_16_30_y0;
  wire f_s_dadda_pg_rca32_fa607_y0;
  wire f_s_dadda_pg_rca32_fa607_y1;
  wire f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_nand_15_31_y0;
  wire f_s_dadda_pg_rca32_fa607_y2;
  wire f_s_dadda_pg_rca32_fa607_y3;
  wire f_s_dadda_pg_rca32_fa607_y4;
  wire f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa598_y2;
  wire f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa599_y2;
  wire f_s_dadda_pg_rca32_fa608_y0;
  wire f_s_dadda_pg_rca32_fa608_y1;
  wire f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa600_y2;
  wire f_s_dadda_pg_rca32_fa608_y2;
  wire f_s_dadda_pg_rca32_fa608_y3;
  wire f_s_dadda_pg_rca32_fa608_y4;
  wire f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa601_y2;
  wire f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa602_y2;
  wire f_s_dadda_pg_rca32_fa609_y0;
  wire f_s_dadda_pg_rca32_fa609_y1;
  wire f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa603_y2;
  wire f_s_dadda_pg_rca32_fa609_y2;
  wire f_s_dadda_pg_rca32_fa609_y3;
  wire f_s_dadda_pg_rca32_fa609_y4;
  wire f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa609_y4;
  wire f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa608_y4;
  wire f_s_dadda_pg_rca32_fa610_y0;
  wire f_s_dadda_pg_rca32_fa610_y1;
  wire f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa607_y4;
  wire f_s_dadda_pg_rca32_fa610_y2;
  wire f_s_dadda_pg_rca32_fa610_y3;
  wire f_s_dadda_pg_rca32_fa610_y4;
  wire f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa606_y4;
  wire f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa605_y4;
  wire f_s_dadda_pg_rca32_fa611_y0;
  wire f_s_dadda_pg_rca32_fa611_y1;
  wire f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa604_y4;
  wire f_s_dadda_pg_rca32_fa611_y2;
  wire f_s_dadda_pg_rca32_fa611_y3;
  wire f_s_dadda_pg_rca32_fa611_y4;
  wire f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa603_y4;
  wire f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa602_y4;
  wire f_s_dadda_pg_rca32_fa612_y0;
  wire f_s_dadda_pg_rca32_fa612_y1;
  wire f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa601_y4;
  wire f_s_dadda_pg_rca32_fa612_y2;
  wire f_s_dadda_pg_rca32_fa612_y3;
  wire f_s_dadda_pg_rca32_fa612_y4;
  wire f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa600_y4;
  wire f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa599_y4;
  wire f_s_dadda_pg_rca32_fa613_y0;
  wire f_s_dadda_pg_rca32_fa613_y1;
  wire f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa598_y4;
  wire f_s_dadda_pg_rca32_fa613_y2;
  wire f_s_dadda_pg_rca32_fa613_y3;
  wire f_s_dadda_pg_rca32_fa613_y4;
  wire f_s_dadda_pg_rca32_nand_31_16_a_31;
  wire f_s_dadda_pg_rca32_nand_31_16_b_16;
  wire f_s_dadda_pg_rca32_nand_31_16_y0;
  wire f_s_dadda_pg_rca32_and_30_17_a_30;
  wire f_s_dadda_pg_rca32_and_30_17_b_17;
  wire f_s_dadda_pg_rca32_and_30_17_y0;
  wire f_s_dadda_pg_rca32_and_29_18_a_29;
  wire f_s_dadda_pg_rca32_and_29_18_b_18;
  wire f_s_dadda_pg_rca32_and_29_18_y0;
  wire f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_nand_31_16_y0;
  wire f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_and_30_17_y0;
  wire f_s_dadda_pg_rca32_fa614_y0;
  wire f_s_dadda_pg_rca32_fa614_y1;
  wire f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_and_29_18_y0;
  wire f_s_dadda_pg_rca32_fa614_y2;
  wire f_s_dadda_pg_rca32_fa614_y3;
  wire f_s_dadda_pg_rca32_fa614_y4;
  wire f_s_dadda_pg_rca32_and_28_19_a_28;
  wire f_s_dadda_pg_rca32_and_28_19_b_19;
  wire f_s_dadda_pg_rca32_and_28_19_y0;
  wire f_s_dadda_pg_rca32_and_27_20_a_27;
  wire f_s_dadda_pg_rca32_and_27_20_b_20;
  wire f_s_dadda_pg_rca32_and_27_20_y0;
  wire f_s_dadda_pg_rca32_and_26_21_a_26;
  wire f_s_dadda_pg_rca32_and_26_21_b_21;
  wire f_s_dadda_pg_rca32_and_26_21_y0;
  wire f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_28_19_y0;
  wire f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_27_20_y0;
  wire f_s_dadda_pg_rca32_fa615_y0;
  wire f_s_dadda_pg_rca32_fa615_y1;
  wire f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_26_21_y0;
  wire f_s_dadda_pg_rca32_fa615_y2;
  wire f_s_dadda_pg_rca32_fa615_y3;
  wire f_s_dadda_pg_rca32_fa615_y4;
  wire f_s_dadda_pg_rca32_and_25_22_a_25;
  wire f_s_dadda_pg_rca32_and_25_22_b_22;
  wire f_s_dadda_pg_rca32_and_25_22_y0;
  wire f_s_dadda_pg_rca32_and_24_23_a_24;
  wire f_s_dadda_pg_rca32_and_24_23_b_23;
  wire f_s_dadda_pg_rca32_and_24_23_y0;
  wire f_s_dadda_pg_rca32_and_23_24_a_23;
  wire f_s_dadda_pg_rca32_and_23_24_b_24;
  wire f_s_dadda_pg_rca32_and_23_24_y0;
  wire f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_25_22_y0;
  wire f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_24_23_y0;
  wire f_s_dadda_pg_rca32_fa616_y0;
  wire f_s_dadda_pg_rca32_fa616_y1;
  wire f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_23_24_y0;
  wire f_s_dadda_pg_rca32_fa616_y2;
  wire f_s_dadda_pg_rca32_fa616_y3;
  wire f_s_dadda_pg_rca32_fa616_y4;
  wire f_s_dadda_pg_rca32_and_22_25_a_22;
  wire f_s_dadda_pg_rca32_and_22_25_b_25;
  wire f_s_dadda_pg_rca32_and_22_25_y0;
  wire f_s_dadda_pg_rca32_and_21_26_a_21;
  wire f_s_dadda_pg_rca32_and_21_26_b_26;
  wire f_s_dadda_pg_rca32_and_21_26_y0;
  wire f_s_dadda_pg_rca32_and_20_27_a_20;
  wire f_s_dadda_pg_rca32_and_20_27_b_27;
  wire f_s_dadda_pg_rca32_and_20_27_y0;
  wire f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_22_25_y0;
  wire f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_21_26_y0;
  wire f_s_dadda_pg_rca32_fa617_y0;
  wire f_s_dadda_pg_rca32_fa617_y1;
  wire f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_20_27_y0;
  wire f_s_dadda_pg_rca32_fa617_y2;
  wire f_s_dadda_pg_rca32_fa617_y3;
  wire f_s_dadda_pg_rca32_fa617_y4;
  wire f_s_dadda_pg_rca32_and_19_28_a_19;
  wire f_s_dadda_pg_rca32_and_19_28_b_28;
  wire f_s_dadda_pg_rca32_and_19_28_y0;
  wire f_s_dadda_pg_rca32_and_18_29_a_18;
  wire f_s_dadda_pg_rca32_and_18_29_b_29;
  wire f_s_dadda_pg_rca32_and_18_29_y0;
  wire f_s_dadda_pg_rca32_and_17_30_a_17;
  wire f_s_dadda_pg_rca32_and_17_30_b_30;
  wire f_s_dadda_pg_rca32_and_17_30_y0;
  wire f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_19_28_y0;
  wire f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_18_29_y0;
  wire f_s_dadda_pg_rca32_fa618_y0;
  wire f_s_dadda_pg_rca32_fa618_y1;
  wire f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_17_30_y0;
  wire f_s_dadda_pg_rca32_fa618_y2;
  wire f_s_dadda_pg_rca32_fa618_y3;
  wire f_s_dadda_pg_rca32_fa618_y4;
  wire f_s_dadda_pg_rca32_nand_16_31_a_16;
  wire f_s_dadda_pg_rca32_nand_16_31_b_31;
  wire f_s_dadda_pg_rca32_nand_16_31_y0;
  wire f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_nand_16_31_y0;
  wire f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_fa610_y2;
  wire f_s_dadda_pg_rca32_fa619_y0;
  wire f_s_dadda_pg_rca32_fa619_y1;
  wire f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_fa611_y2;
  wire f_s_dadda_pg_rca32_fa619_y2;
  wire f_s_dadda_pg_rca32_fa619_y3;
  wire f_s_dadda_pg_rca32_fa619_y4;
  wire f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa612_y2;
  wire f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa613_y2;
  wire f_s_dadda_pg_rca32_fa620_y0;
  wire f_s_dadda_pg_rca32_fa620_y1;
  wire f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa614_y2;
  wire f_s_dadda_pg_rca32_fa620_y2;
  wire f_s_dadda_pg_rca32_fa620_y3;
  wire f_s_dadda_pg_rca32_fa620_y4;
  wire f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa620_y4;
  wire f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa619_y4;
  wire f_s_dadda_pg_rca32_fa621_y0;
  wire f_s_dadda_pg_rca32_fa621_y1;
  wire f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa618_y4;
  wire f_s_dadda_pg_rca32_fa621_y2;
  wire f_s_dadda_pg_rca32_fa621_y3;
  wire f_s_dadda_pg_rca32_fa621_y4;
  wire f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa617_y4;
  wire f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa616_y4;
  wire f_s_dadda_pg_rca32_fa622_y0;
  wire f_s_dadda_pg_rca32_fa622_y1;
  wire f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa615_y4;
  wire f_s_dadda_pg_rca32_fa622_y2;
  wire f_s_dadda_pg_rca32_fa622_y3;
  wire f_s_dadda_pg_rca32_fa622_y4;
  wire f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa614_y4;
  wire f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa613_y4;
  wire f_s_dadda_pg_rca32_fa623_y0;
  wire f_s_dadda_pg_rca32_fa623_y1;
  wire f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa612_y4;
  wire f_s_dadda_pg_rca32_fa623_y2;
  wire f_s_dadda_pg_rca32_fa623_y3;
  wire f_s_dadda_pg_rca32_fa623_y4;
  wire f_s_dadda_pg_rca32_nand_31_17_a_31;
  wire f_s_dadda_pg_rca32_nand_31_17_b_17;
  wire f_s_dadda_pg_rca32_nand_31_17_y0;
  wire f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_fa611_y4;
  wire f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_fa610_y4;
  wire f_s_dadda_pg_rca32_fa624_y0;
  wire f_s_dadda_pg_rca32_fa624_y1;
  wire f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_nand_31_17_y0;
  wire f_s_dadda_pg_rca32_fa624_y2;
  wire f_s_dadda_pg_rca32_fa624_y3;
  wire f_s_dadda_pg_rca32_fa624_y4;
  wire f_s_dadda_pg_rca32_and_30_18_a_30;
  wire f_s_dadda_pg_rca32_and_30_18_b_18;
  wire f_s_dadda_pg_rca32_and_30_18_y0;
  wire f_s_dadda_pg_rca32_and_29_19_a_29;
  wire f_s_dadda_pg_rca32_and_29_19_b_19;
  wire f_s_dadda_pg_rca32_and_29_19_y0;
  wire f_s_dadda_pg_rca32_and_28_20_a_28;
  wire f_s_dadda_pg_rca32_and_28_20_b_20;
  wire f_s_dadda_pg_rca32_and_28_20_y0;
  wire f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_30_18_y0;
  wire f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_29_19_y0;
  wire f_s_dadda_pg_rca32_fa625_y0;
  wire f_s_dadda_pg_rca32_fa625_y1;
  wire f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_28_20_y0;
  wire f_s_dadda_pg_rca32_fa625_y2;
  wire f_s_dadda_pg_rca32_fa625_y3;
  wire f_s_dadda_pg_rca32_fa625_y4;
  wire f_s_dadda_pg_rca32_and_27_21_a_27;
  wire f_s_dadda_pg_rca32_and_27_21_b_21;
  wire f_s_dadda_pg_rca32_and_27_21_y0;
  wire f_s_dadda_pg_rca32_and_26_22_a_26;
  wire f_s_dadda_pg_rca32_and_26_22_b_22;
  wire f_s_dadda_pg_rca32_and_26_22_y0;
  wire f_s_dadda_pg_rca32_and_25_23_a_25;
  wire f_s_dadda_pg_rca32_and_25_23_b_23;
  wire f_s_dadda_pg_rca32_and_25_23_y0;
  wire f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_27_21_y0;
  wire f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_26_22_y0;
  wire f_s_dadda_pg_rca32_fa626_y0;
  wire f_s_dadda_pg_rca32_fa626_y1;
  wire f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_25_23_y0;
  wire f_s_dadda_pg_rca32_fa626_y2;
  wire f_s_dadda_pg_rca32_fa626_y3;
  wire f_s_dadda_pg_rca32_fa626_y4;
  wire f_s_dadda_pg_rca32_and_24_24_a_24;
  wire f_s_dadda_pg_rca32_and_24_24_b_24;
  wire f_s_dadda_pg_rca32_and_24_24_y0;
  wire f_s_dadda_pg_rca32_and_23_25_a_23;
  wire f_s_dadda_pg_rca32_and_23_25_b_25;
  wire f_s_dadda_pg_rca32_and_23_25_y0;
  wire f_s_dadda_pg_rca32_and_22_26_a_22;
  wire f_s_dadda_pg_rca32_and_22_26_b_26;
  wire f_s_dadda_pg_rca32_and_22_26_y0;
  wire f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_24_24_y0;
  wire f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_23_25_y0;
  wire f_s_dadda_pg_rca32_fa627_y0;
  wire f_s_dadda_pg_rca32_fa627_y1;
  wire f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_22_26_y0;
  wire f_s_dadda_pg_rca32_fa627_y2;
  wire f_s_dadda_pg_rca32_fa627_y3;
  wire f_s_dadda_pg_rca32_fa627_y4;
  wire f_s_dadda_pg_rca32_and_21_27_a_21;
  wire f_s_dadda_pg_rca32_and_21_27_b_27;
  wire f_s_dadda_pg_rca32_and_21_27_y0;
  wire f_s_dadda_pg_rca32_and_20_28_a_20;
  wire f_s_dadda_pg_rca32_and_20_28_b_28;
  wire f_s_dadda_pg_rca32_and_20_28_y0;
  wire f_s_dadda_pg_rca32_and_19_29_a_19;
  wire f_s_dadda_pg_rca32_and_19_29_b_29;
  wire f_s_dadda_pg_rca32_and_19_29_y0;
  wire f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_21_27_y0;
  wire f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_20_28_y0;
  wire f_s_dadda_pg_rca32_fa628_y0;
  wire f_s_dadda_pg_rca32_fa628_y1;
  wire f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_19_29_y0;
  wire f_s_dadda_pg_rca32_fa628_y2;
  wire f_s_dadda_pg_rca32_fa628_y3;
  wire f_s_dadda_pg_rca32_fa628_y4;
  wire f_s_dadda_pg_rca32_and_18_30_a_18;
  wire f_s_dadda_pg_rca32_and_18_30_b_30;
  wire f_s_dadda_pg_rca32_and_18_30_y0;
  wire f_s_dadda_pg_rca32_nand_17_31_a_17;
  wire f_s_dadda_pg_rca32_nand_17_31_b_31;
  wire f_s_dadda_pg_rca32_nand_17_31_y0;
  wire f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_and_18_30_y0;
  wire f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_nand_17_31_y0;
  wire f_s_dadda_pg_rca32_fa629_y0;
  wire f_s_dadda_pg_rca32_fa629_y1;
  wire f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_fa621_y2;
  wire f_s_dadda_pg_rca32_fa629_y2;
  wire f_s_dadda_pg_rca32_fa629_y3;
  wire f_s_dadda_pg_rca32_fa629_y4;
  wire f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa622_y2;
  wire f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa623_y2;
  wire f_s_dadda_pg_rca32_fa630_y0;
  wire f_s_dadda_pg_rca32_fa630_y1;
  wire f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa624_y2;
  wire f_s_dadda_pg_rca32_fa630_y2;
  wire f_s_dadda_pg_rca32_fa630_y3;
  wire f_s_dadda_pg_rca32_fa630_y4;
  wire f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa630_y4;
  wire f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa629_y4;
  wire f_s_dadda_pg_rca32_fa631_y0;
  wire f_s_dadda_pg_rca32_fa631_y1;
  wire f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa628_y4;
  wire f_s_dadda_pg_rca32_fa631_y2;
  wire f_s_dadda_pg_rca32_fa631_y3;
  wire f_s_dadda_pg_rca32_fa631_y4;
  wire f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa627_y4;
  wire f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa626_y4;
  wire f_s_dadda_pg_rca32_fa632_y0;
  wire f_s_dadda_pg_rca32_fa632_y1;
  wire f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa625_y4;
  wire f_s_dadda_pg_rca32_fa632_y2;
  wire f_s_dadda_pg_rca32_fa632_y3;
  wire f_s_dadda_pg_rca32_fa632_y4;
  wire f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa624_y4;
  wire f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa623_y4;
  wire f_s_dadda_pg_rca32_fa633_y0;
  wire f_s_dadda_pg_rca32_fa633_y1;
  wire f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa622_y4;
  wire f_s_dadda_pg_rca32_fa633_y2;
  wire f_s_dadda_pg_rca32_fa633_y3;
  wire f_s_dadda_pg_rca32_fa633_y4;
  wire f_s_dadda_pg_rca32_nand_31_18_a_31;
  wire f_s_dadda_pg_rca32_nand_31_18_b_18;
  wire f_s_dadda_pg_rca32_nand_31_18_y0;
  wire f_s_dadda_pg_rca32_and_30_19_a_30;
  wire f_s_dadda_pg_rca32_and_30_19_b_19;
  wire f_s_dadda_pg_rca32_and_30_19_y0;
  wire f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_fa621_y4;
  wire f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_nand_31_18_y0;
  wire f_s_dadda_pg_rca32_fa634_y0;
  wire f_s_dadda_pg_rca32_fa634_y1;
  wire f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_and_30_19_y0;
  wire f_s_dadda_pg_rca32_fa634_y2;
  wire f_s_dadda_pg_rca32_fa634_y3;
  wire f_s_dadda_pg_rca32_fa634_y4;
  wire f_s_dadda_pg_rca32_and_29_20_a_29;
  wire f_s_dadda_pg_rca32_and_29_20_b_20;
  wire f_s_dadda_pg_rca32_and_29_20_y0;
  wire f_s_dadda_pg_rca32_and_28_21_a_28;
  wire f_s_dadda_pg_rca32_and_28_21_b_21;
  wire f_s_dadda_pg_rca32_and_28_21_y0;
  wire f_s_dadda_pg_rca32_and_27_22_a_27;
  wire f_s_dadda_pg_rca32_and_27_22_b_22;
  wire f_s_dadda_pg_rca32_and_27_22_y0;
  wire f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_29_20_y0;
  wire f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_28_21_y0;
  wire f_s_dadda_pg_rca32_fa635_y0;
  wire f_s_dadda_pg_rca32_fa635_y1;
  wire f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_27_22_y0;
  wire f_s_dadda_pg_rca32_fa635_y2;
  wire f_s_dadda_pg_rca32_fa635_y3;
  wire f_s_dadda_pg_rca32_fa635_y4;
  wire f_s_dadda_pg_rca32_and_26_23_a_26;
  wire f_s_dadda_pg_rca32_and_26_23_b_23;
  wire f_s_dadda_pg_rca32_and_26_23_y0;
  wire f_s_dadda_pg_rca32_and_25_24_a_25;
  wire f_s_dadda_pg_rca32_and_25_24_b_24;
  wire f_s_dadda_pg_rca32_and_25_24_y0;
  wire f_s_dadda_pg_rca32_and_24_25_a_24;
  wire f_s_dadda_pg_rca32_and_24_25_b_25;
  wire f_s_dadda_pg_rca32_and_24_25_y0;
  wire f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_26_23_y0;
  wire f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_25_24_y0;
  wire f_s_dadda_pg_rca32_fa636_y0;
  wire f_s_dadda_pg_rca32_fa636_y1;
  wire f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_24_25_y0;
  wire f_s_dadda_pg_rca32_fa636_y2;
  wire f_s_dadda_pg_rca32_fa636_y3;
  wire f_s_dadda_pg_rca32_fa636_y4;
  wire f_s_dadda_pg_rca32_and_23_26_a_23;
  wire f_s_dadda_pg_rca32_and_23_26_b_26;
  wire f_s_dadda_pg_rca32_and_23_26_y0;
  wire f_s_dadda_pg_rca32_and_22_27_a_22;
  wire f_s_dadda_pg_rca32_and_22_27_b_27;
  wire f_s_dadda_pg_rca32_and_22_27_y0;
  wire f_s_dadda_pg_rca32_and_21_28_a_21;
  wire f_s_dadda_pg_rca32_and_21_28_b_28;
  wire f_s_dadda_pg_rca32_and_21_28_y0;
  wire f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_23_26_y0;
  wire f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_22_27_y0;
  wire f_s_dadda_pg_rca32_fa637_y0;
  wire f_s_dadda_pg_rca32_fa637_y1;
  wire f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_21_28_y0;
  wire f_s_dadda_pg_rca32_fa637_y2;
  wire f_s_dadda_pg_rca32_fa637_y3;
  wire f_s_dadda_pg_rca32_fa637_y4;
  wire f_s_dadda_pg_rca32_and_20_29_a_20;
  wire f_s_dadda_pg_rca32_and_20_29_b_29;
  wire f_s_dadda_pg_rca32_and_20_29_y0;
  wire f_s_dadda_pg_rca32_and_19_30_a_19;
  wire f_s_dadda_pg_rca32_and_19_30_b_30;
  wire f_s_dadda_pg_rca32_and_19_30_y0;
  wire f_s_dadda_pg_rca32_nand_18_31_a_18;
  wire f_s_dadda_pg_rca32_nand_18_31_b_31;
  wire f_s_dadda_pg_rca32_nand_18_31_y0;
  wire f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_and_20_29_y0;
  wire f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_and_19_30_y0;
  wire f_s_dadda_pg_rca32_fa638_y0;
  wire f_s_dadda_pg_rca32_fa638_y1;
  wire f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_nand_18_31_y0;
  wire f_s_dadda_pg_rca32_fa638_y2;
  wire f_s_dadda_pg_rca32_fa638_y3;
  wire f_s_dadda_pg_rca32_fa638_y4;
  wire f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa631_y2;
  wire f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa632_y2;
  wire f_s_dadda_pg_rca32_fa639_y0;
  wire f_s_dadda_pg_rca32_fa639_y1;
  wire f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa633_y2;
  wire f_s_dadda_pg_rca32_fa639_y2;
  wire f_s_dadda_pg_rca32_fa639_y3;
  wire f_s_dadda_pg_rca32_fa639_y4;
  wire f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa639_y4;
  wire f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa638_y4;
  wire f_s_dadda_pg_rca32_fa640_y0;
  wire f_s_dadda_pg_rca32_fa640_y1;
  wire f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa637_y4;
  wire f_s_dadda_pg_rca32_fa640_y2;
  wire f_s_dadda_pg_rca32_fa640_y3;
  wire f_s_dadda_pg_rca32_fa640_y4;
  wire f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa636_y4;
  wire f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa635_y4;
  wire f_s_dadda_pg_rca32_fa641_y0;
  wire f_s_dadda_pg_rca32_fa641_y1;
  wire f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa634_y4;
  wire f_s_dadda_pg_rca32_fa641_y2;
  wire f_s_dadda_pg_rca32_fa641_y3;
  wire f_s_dadda_pg_rca32_fa641_y4;
  wire f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa633_y4;
  wire f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa632_y4;
  wire f_s_dadda_pg_rca32_fa642_y0;
  wire f_s_dadda_pg_rca32_fa642_y1;
  wire f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa631_y4;
  wire f_s_dadda_pg_rca32_fa642_y2;
  wire f_s_dadda_pg_rca32_fa642_y3;
  wire f_s_dadda_pg_rca32_fa642_y4;
  wire f_s_dadda_pg_rca32_nand_31_19_a_31;
  wire f_s_dadda_pg_rca32_nand_31_19_b_19;
  wire f_s_dadda_pg_rca32_nand_31_19_y0;
  wire f_s_dadda_pg_rca32_and_30_20_a_30;
  wire f_s_dadda_pg_rca32_and_30_20_b_20;
  wire f_s_dadda_pg_rca32_and_30_20_y0;
  wire f_s_dadda_pg_rca32_and_29_21_a_29;
  wire f_s_dadda_pg_rca32_and_29_21_b_21;
  wire f_s_dadda_pg_rca32_and_29_21_y0;
  wire f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_nand_31_19_y0;
  wire f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_and_30_20_y0;
  wire f_s_dadda_pg_rca32_fa643_y0;
  wire f_s_dadda_pg_rca32_fa643_y1;
  wire f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_and_29_21_y0;
  wire f_s_dadda_pg_rca32_fa643_y2;
  wire f_s_dadda_pg_rca32_fa643_y3;
  wire f_s_dadda_pg_rca32_fa643_y4;
  wire f_s_dadda_pg_rca32_and_28_22_a_28;
  wire f_s_dadda_pg_rca32_and_28_22_b_22;
  wire f_s_dadda_pg_rca32_and_28_22_y0;
  wire f_s_dadda_pg_rca32_and_27_23_a_27;
  wire f_s_dadda_pg_rca32_and_27_23_b_23;
  wire f_s_dadda_pg_rca32_and_27_23_y0;
  wire f_s_dadda_pg_rca32_and_26_24_a_26;
  wire f_s_dadda_pg_rca32_and_26_24_b_24;
  wire f_s_dadda_pg_rca32_and_26_24_y0;
  wire f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_28_22_y0;
  wire f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_27_23_y0;
  wire f_s_dadda_pg_rca32_fa644_y0;
  wire f_s_dadda_pg_rca32_fa644_y1;
  wire f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_26_24_y0;
  wire f_s_dadda_pg_rca32_fa644_y2;
  wire f_s_dadda_pg_rca32_fa644_y3;
  wire f_s_dadda_pg_rca32_fa644_y4;
  wire f_s_dadda_pg_rca32_and_25_25_a_25;
  wire f_s_dadda_pg_rca32_and_25_25_b_25;
  wire f_s_dadda_pg_rca32_and_25_25_y0;
  wire f_s_dadda_pg_rca32_and_24_26_a_24;
  wire f_s_dadda_pg_rca32_and_24_26_b_26;
  wire f_s_dadda_pg_rca32_and_24_26_y0;
  wire f_s_dadda_pg_rca32_and_23_27_a_23;
  wire f_s_dadda_pg_rca32_and_23_27_b_27;
  wire f_s_dadda_pg_rca32_and_23_27_y0;
  wire f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_25_25_y0;
  wire f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_24_26_y0;
  wire f_s_dadda_pg_rca32_fa645_y0;
  wire f_s_dadda_pg_rca32_fa645_y1;
  wire f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_23_27_y0;
  wire f_s_dadda_pg_rca32_fa645_y2;
  wire f_s_dadda_pg_rca32_fa645_y3;
  wire f_s_dadda_pg_rca32_fa645_y4;
  wire f_s_dadda_pg_rca32_and_22_28_a_22;
  wire f_s_dadda_pg_rca32_and_22_28_b_28;
  wire f_s_dadda_pg_rca32_and_22_28_y0;
  wire f_s_dadda_pg_rca32_and_21_29_a_21;
  wire f_s_dadda_pg_rca32_and_21_29_b_29;
  wire f_s_dadda_pg_rca32_and_21_29_y0;
  wire f_s_dadda_pg_rca32_and_20_30_a_20;
  wire f_s_dadda_pg_rca32_and_20_30_b_30;
  wire f_s_dadda_pg_rca32_and_20_30_y0;
  wire f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_22_28_y0;
  wire f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_21_29_y0;
  wire f_s_dadda_pg_rca32_fa646_y0;
  wire f_s_dadda_pg_rca32_fa646_y1;
  wire f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_20_30_y0;
  wire f_s_dadda_pg_rca32_fa646_y2;
  wire f_s_dadda_pg_rca32_fa646_y3;
  wire f_s_dadda_pg_rca32_fa646_y4;
  wire f_s_dadda_pg_rca32_nand_19_31_a_19;
  wire f_s_dadda_pg_rca32_nand_19_31_b_31;
  wire f_s_dadda_pg_rca32_nand_19_31_y0;
  wire f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_nand_19_31_y0;
  wire f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_fa640_y2;
  wire f_s_dadda_pg_rca32_fa647_y0;
  wire f_s_dadda_pg_rca32_fa647_y1;
  wire f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_fa641_y2;
  wire f_s_dadda_pg_rca32_fa647_y2;
  wire f_s_dadda_pg_rca32_fa647_y3;
  wire f_s_dadda_pg_rca32_fa647_y4;
  wire f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa647_y4;
  wire f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa646_y4;
  wire f_s_dadda_pg_rca32_fa648_y0;
  wire f_s_dadda_pg_rca32_fa648_y1;
  wire f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa645_y4;
  wire f_s_dadda_pg_rca32_fa648_y2;
  wire f_s_dadda_pg_rca32_fa648_y3;
  wire f_s_dadda_pg_rca32_fa648_y4;
  wire f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa644_y4;
  wire f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa643_y4;
  wire f_s_dadda_pg_rca32_fa649_y0;
  wire f_s_dadda_pg_rca32_fa649_y1;
  wire f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa642_y4;
  wire f_s_dadda_pg_rca32_fa649_y2;
  wire f_s_dadda_pg_rca32_fa649_y3;
  wire f_s_dadda_pg_rca32_fa649_y4;
  wire f_s_dadda_pg_rca32_nand_31_20_a_31;
  wire f_s_dadda_pg_rca32_nand_31_20_b_20;
  wire f_s_dadda_pg_rca32_nand_31_20_y0;
  wire f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_fa641_y4;
  wire f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_fa640_y4;
  wire f_s_dadda_pg_rca32_fa650_y0;
  wire f_s_dadda_pg_rca32_fa650_y1;
  wire f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_nand_31_20_y0;
  wire f_s_dadda_pg_rca32_fa650_y2;
  wire f_s_dadda_pg_rca32_fa650_y3;
  wire f_s_dadda_pg_rca32_fa650_y4;
  wire f_s_dadda_pg_rca32_and_30_21_a_30;
  wire f_s_dadda_pg_rca32_and_30_21_b_21;
  wire f_s_dadda_pg_rca32_and_30_21_y0;
  wire f_s_dadda_pg_rca32_and_29_22_a_29;
  wire f_s_dadda_pg_rca32_and_29_22_b_22;
  wire f_s_dadda_pg_rca32_and_29_22_y0;
  wire f_s_dadda_pg_rca32_and_28_23_a_28;
  wire f_s_dadda_pg_rca32_and_28_23_b_23;
  wire f_s_dadda_pg_rca32_and_28_23_y0;
  wire f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_30_21_y0;
  wire f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_29_22_y0;
  wire f_s_dadda_pg_rca32_fa651_y0;
  wire f_s_dadda_pg_rca32_fa651_y1;
  wire f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_28_23_y0;
  wire f_s_dadda_pg_rca32_fa651_y2;
  wire f_s_dadda_pg_rca32_fa651_y3;
  wire f_s_dadda_pg_rca32_fa651_y4;
  wire f_s_dadda_pg_rca32_and_27_24_a_27;
  wire f_s_dadda_pg_rca32_and_27_24_b_24;
  wire f_s_dadda_pg_rca32_and_27_24_y0;
  wire f_s_dadda_pg_rca32_and_26_25_a_26;
  wire f_s_dadda_pg_rca32_and_26_25_b_25;
  wire f_s_dadda_pg_rca32_and_26_25_y0;
  wire f_s_dadda_pg_rca32_and_25_26_a_25;
  wire f_s_dadda_pg_rca32_and_25_26_b_26;
  wire f_s_dadda_pg_rca32_and_25_26_y0;
  wire f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_27_24_y0;
  wire f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_26_25_y0;
  wire f_s_dadda_pg_rca32_fa652_y0;
  wire f_s_dadda_pg_rca32_fa652_y1;
  wire f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_25_26_y0;
  wire f_s_dadda_pg_rca32_fa652_y2;
  wire f_s_dadda_pg_rca32_fa652_y3;
  wire f_s_dadda_pg_rca32_fa652_y4;
  wire f_s_dadda_pg_rca32_and_24_27_a_24;
  wire f_s_dadda_pg_rca32_and_24_27_b_27;
  wire f_s_dadda_pg_rca32_and_24_27_y0;
  wire f_s_dadda_pg_rca32_and_23_28_a_23;
  wire f_s_dadda_pg_rca32_and_23_28_b_28;
  wire f_s_dadda_pg_rca32_and_23_28_y0;
  wire f_s_dadda_pg_rca32_and_22_29_a_22;
  wire f_s_dadda_pg_rca32_and_22_29_b_29;
  wire f_s_dadda_pg_rca32_and_22_29_y0;
  wire f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_24_27_y0;
  wire f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_23_28_y0;
  wire f_s_dadda_pg_rca32_fa653_y0;
  wire f_s_dadda_pg_rca32_fa653_y1;
  wire f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_22_29_y0;
  wire f_s_dadda_pg_rca32_fa653_y2;
  wire f_s_dadda_pg_rca32_fa653_y3;
  wire f_s_dadda_pg_rca32_fa653_y4;
  wire f_s_dadda_pg_rca32_and_21_30_a_21;
  wire f_s_dadda_pg_rca32_and_21_30_b_30;
  wire f_s_dadda_pg_rca32_and_21_30_y0;
  wire f_s_dadda_pg_rca32_nand_20_31_a_20;
  wire f_s_dadda_pg_rca32_nand_20_31_b_31;
  wire f_s_dadda_pg_rca32_nand_20_31_y0;
  wire f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_and_21_30_y0;
  wire f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_nand_20_31_y0;
  wire f_s_dadda_pg_rca32_fa654_y0;
  wire f_s_dadda_pg_rca32_fa654_y1;
  wire f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_fa648_y2;
  wire f_s_dadda_pg_rca32_fa654_y2;
  wire f_s_dadda_pg_rca32_fa654_y3;
  wire f_s_dadda_pg_rca32_fa654_y4;
  wire f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa654_y4;
  wire f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa653_y4;
  wire f_s_dadda_pg_rca32_fa655_y0;
  wire f_s_dadda_pg_rca32_fa655_y1;
  wire f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa652_y4;
  wire f_s_dadda_pg_rca32_fa655_y2;
  wire f_s_dadda_pg_rca32_fa655_y3;
  wire f_s_dadda_pg_rca32_fa655_y4;
  wire f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa651_y4;
  wire f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa650_y4;
  wire f_s_dadda_pg_rca32_fa656_y0;
  wire f_s_dadda_pg_rca32_fa656_y1;
  wire f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa649_y4;
  wire f_s_dadda_pg_rca32_fa656_y2;
  wire f_s_dadda_pg_rca32_fa656_y3;
  wire f_s_dadda_pg_rca32_fa656_y4;
  wire f_s_dadda_pg_rca32_nand_31_21_a_31;
  wire f_s_dadda_pg_rca32_nand_31_21_b_21;
  wire f_s_dadda_pg_rca32_nand_31_21_y0;
  wire f_s_dadda_pg_rca32_and_30_22_a_30;
  wire f_s_dadda_pg_rca32_and_30_22_b_22;
  wire f_s_dadda_pg_rca32_and_30_22_y0;
  wire f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_fa648_y4;
  wire f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_nand_31_21_y0;
  wire f_s_dadda_pg_rca32_fa657_y0;
  wire f_s_dadda_pg_rca32_fa657_y1;
  wire f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_and_30_22_y0;
  wire f_s_dadda_pg_rca32_fa657_y2;
  wire f_s_dadda_pg_rca32_fa657_y3;
  wire f_s_dadda_pg_rca32_fa657_y4;
  wire f_s_dadda_pg_rca32_and_29_23_a_29;
  wire f_s_dadda_pg_rca32_and_29_23_b_23;
  wire f_s_dadda_pg_rca32_and_29_23_y0;
  wire f_s_dadda_pg_rca32_and_28_24_a_28;
  wire f_s_dadda_pg_rca32_and_28_24_b_24;
  wire f_s_dadda_pg_rca32_and_28_24_y0;
  wire f_s_dadda_pg_rca32_and_27_25_a_27;
  wire f_s_dadda_pg_rca32_and_27_25_b_25;
  wire f_s_dadda_pg_rca32_and_27_25_y0;
  wire f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_29_23_y0;
  wire f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_28_24_y0;
  wire f_s_dadda_pg_rca32_fa658_y0;
  wire f_s_dadda_pg_rca32_fa658_y1;
  wire f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_27_25_y0;
  wire f_s_dadda_pg_rca32_fa658_y2;
  wire f_s_dadda_pg_rca32_fa658_y3;
  wire f_s_dadda_pg_rca32_fa658_y4;
  wire f_s_dadda_pg_rca32_and_26_26_a_26;
  wire f_s_dadda_pg_rca32_and_26_26_b_26;
  wire f_s_dadda_pg_rca32_and_26_26_y0;
  wire f_s_dadda_pg_rca32_and_25_27_a_25;
  wire f_s_dadda_pg_rca32_and_25_27_b_27;
  wire f_s_dadda_pg_rca32_and_25_27_y0;
  wire f_s_dadda_pg_rca32_and_24_28_a_24;
  wire f_s_dadda_pg_rca32_and_24_28_b_28;
  wire f_s_dadda_pg_rca32_and_24_28_y0;
  wire f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_26_26_y0;
  wire f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_25_27_y0;
  wire f_s_dadda_pg_rca32_fa659_y0;
  wire f_s_dadda_pg_rca32_fa659_y1;
  wire f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_24_28_y0;
  wire f_s_dadda_pg_rca32_fa659_y2;
  wire f_s_dadda_pg_rca32_fa659_y3;
  wire f_s_dadda_pg_rca32_fa659_y4;
  wire f_s_dadda_pg_rca32_and_23_29_a_23;
  wire f_s_dadda_pg_rca32_and_23_29_b_29;
  wire f_s_dadda_pg_rca32_and_23_29_y0;
  wire f_s_dadda_pg_rca32_and_22_30_a_22;
  wire f_s_dadda_pg_rca32_and_22_30_b_30;
  wire f_s_dadda_pg_rca32_and_22_30_y0;
  wire f_s_dadda_pg_rca32_nand_21_31_a_21;
  wire f_s_dadda_pg_rca32_nand_21_31_b_31;
  wire f_s_dadda_pg_rca32_nand_21_31_y0;
  wire f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_and_23_29_y0;
  wire f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_and_22_30_y0;
  wire f_s_dadda_pg_rca32_fa660_y0;
  wire f_s_dadda_pg_rca32_fa660_y1;
  wire f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_nand_21_31_y0;
  wire f_s_dadda_pg_rca32_fa660_y2;
  wire f_s_dadda_pg_rca32_fa660_y3;
  wire f_s_dadda_pg_rca32_fa660_y4;
  wire f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa660_y4;
  wire f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa659_y4;
  wire f_s_dadda_pg_rca32_fa661_y0;
  wire f_s_dadda_pg_rca32_fa661_y1;
  wire f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa658_y4;
  wire f_s_dadda_pg_rca32_fa661_y2;
  wire f_s_dadda_pg_rca32_fa661_y3;
  wire f_s_dadda_pg_rca32_fa661_y4;
  wire f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa657_y4;
  wire f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa656_y4;
  wire f_s_dadda_pg_rca32_fa662_y0;
  wire f_s_dadda_pg_rca32_fa662_y1;
  wire f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa655_y4;
  wire f_s_dadda_pg_rca32_fa662_y2;
  wire f_s_dadda_pg_rca32_fa662_y3;
  wire f_s_dadda_pg_rca32_fa662_y4;
  wire f_s_dadda_pg_rca32_nand_31_22_a_31;
  wire f_s_dadda_pg_rca32_nand_31_22_b_22;
  wire f_s_dadda_pg_rca32_nand_31_22_y0;
  wire f_s_dadda_pg_rca32_and_30_23_a_30;
  wire f_s_dadda_pg_rca32_and_30_23_b_23;
  wire f_s_dadda_pg_rca32_and_30_23_y0;
  wire f_s_dadda_pg_rca32_and_29_24_a_29;
  wire f_s_dadda_pg_rca32_and_29_24_b_24;
  wire f_s_dadda_pg_rca32_and_29_24_y0;
  wire f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_nand_31_22_y0;
  wire f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_and_30_23_y0;
  wire f_s_dadda_pg_rca32_fa663_y0;
  wire f_s_dadda_pg_rca32_fa663_y1;
  wire f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_and_29_24_y0;
  wire f_s_dadda_pg_rca32_fa663_y2;
  wire f_s_dadda_pg_rca32_fa663_y3;
  wire f_s_dadda_pg_rca32_fa663_y4;
  wire f_s_dadda_pg_rca32_and_28_25_a_28;
  wire f_s_dadda_pg_rca32_and_28_25_b_25;
  wire f_s_dadda_pg_rca32_and_28_25_y0;
  wire f_s_dadda_pg_rca32_and_27_26_a_27;
  wire f_s_dadda_pg_rca32_and_27_26_b_26;
  wire f_s_dadda_pg_rca32_and_27_26_y0;
  wire f_s_dadda_pg_rca32_and_26_27_a_26;
  wire f_s_dadda_pg_rca32_and_26_27_b_27;
  wire f_s_dadda_pg_rca32_and_26_27_y0;
  wire f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_28_25_y0;
  wire f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_27_26_y0;
  wire f_s_dadda_pg_rca32_fa664_y0;
  wire f_s_dadda_pg_rca32_fa664_y1;
  wire f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_26_27_y0;
  wire f_s_dadda_pg_rca32_fa664_y2;
  wire f_s_dadda_pg_rca32_fa664_y3;
  wire f_s_dadda_pg_rca32_fa664_y4;
  wire f_s_dadda_pg_rca32_and_25_28_a_25;
  wire f_s_dadda_pg_rca32_and_25_28_b_28;
  wire f_s_dadda_pg_rca32_and_25_28_y0;
  wire f_s_dadda_pg_rca32_and_24_29_a_24;
  wire f_s_dadda_pg_rca32_and_24_29_b_29;
  wire f_s_dadda_pg_rca32_and_24_29_y0;
  wire f_s_dadda_pg_rca32_and_23_30_a_23;
  wire f_s_dadda_pg_rca32_and_23_30_b_30;
  wire f_s_dadda_pg_rca32_and_23_30_y0;
  wire f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_25_28_y0;
  wire f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_24_29_y0;
  wire f_s_dadda_pg_rca32_fa665_y0;
  wire f_s_dadda_pg_rca32_fa665_y1;
  wire f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_23_30_y0;
  wire f_s_dadda_pg_rca32_fa665_y2;
  wire f_s_dadda_pg_rca32_fa665_y3;
  wire f_s_dadda_pg_rca32_fa665_y4;
  wire f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa665_y4;
  wire f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa664_y4;
  wire f_s_dadda_pg_rca32_fa666_y0;
  wire f_s_dadda_pg_rca32_fa666_y1;
  wire f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa663_y4;
  wire f_s_dadda_pg_rca32_fa666_y2;
  wire f_s_dadda_pg_rca32_fa666_y3;
  wire f_s_dadda_pg_rca32_fa666_y4;
  wire f_s_dadda_pg_rca32_nand_31_23_a_31;
  wire f_s_dadda_pg_rca32_nand_31_23_b_23;
  wire f_s_dadda_pg_rca32_nand_31_23_y0;
  wire f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_fa662_y4;
  wire f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_fa661_y4;
  wire f_s_dadda_pg_rca32_fa667_y0;
  wire f_s_dadda_pg_rca32_fa667_y1;
  wire f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_nand_31_23_y0;
  wire f_s_dadda_pg_rca32_fa667_y2;
  wire f_s_dadda_pg_rca32_fa667_y3;
  wire f_s_dadda_pg_rca32_fa667_y4;
  wire f_s_dadda_pg_rca32_and_30_24_a_30;
  wire f_s_dadda_pg_rca32_and_30_24_b_24;
  wire f_s_dadda_pg_rca32_and_30_24_y0;
  wire f_s_dadda_pg_rca32_and_29_25_a_29;
  wire f_s_dadda_pg_rca32_and_29_25_b_25;
  wire f_s_dadda_pg_rca32_and_29_25_y0;
  wire f_s_dadda_pg_rca32_and_28_26_a_28;
  wire f_s_dadda_pg_rca32_and_28_26_b_26;
  wire f_s_dadda_pg_rca32_and_28_26_y0;
  wire f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_30_24_y0;
  wire f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_29_25_y0;
  wire f_s_dadda_pg_rca32_fa668_y0;
  wire f_s_dadda_pg_rca32_fa668_y1;
  wire f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_28_26_y0;
  wire f_s_dadda_pg_rca32_fa668_y2;
  wire f_s_dadda_pg_rca32_fa668_y3;
  wire f_s_dadda_pg_rca32_fa668_y4;
  wire f_s_dadda_pg_rca32_and_27_27_a_27;
  wire f_s_dadda_pg_rca32_and_27_27_b_27;
  wire f_s_dadda_pg_rca32_and_27_27_y0;
  wire f_s_dadda_pg_rca32_and_26_28_a_26;
  wire f_s_dadda_pg_rca32_and_26_28_b_28;
  wire f_s_dadda_pg_rca32_and_26_28_y0;
  wire f_s_dadda_pg_rca32_and_25_29_a_25;
  wire f_s_dadda_pg_rca32_and_25_29_b_29;
  wire f_s_dadda_pg_rca32_and_25_29_y0;
  wire f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_27_27_y0;
  wire f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_26_28_y0;
  wire f_s_dadda_pg_rca32_fa669_y0;
  wire f_s_dadda_pg_rca32_fa669_y1;
  wire f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_25_29_y0;
  wire f_s_dadda_pg_rca32_fa669_y2;
  wire f_s_dadda_pg_rca32_fa669_y3;
  wire f_s_dadda_pg_rca32_fa669_y4;
  wire f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa669_y4;
  wire f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa668_y4;
  wire f_s_dadda_pg_rca32_fa670_y0;
  wire f_s_dadda_pg_rca32_fa670_y1;
  wire f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa667_y4;
  wire f_s_dadda_pg_rca32_fa670_y2;
  wire f_s_dadda_pg_rca32_fa670_y3;
  wire f_s_dadda_pg_rca32_fa670_y4;
  wire f_s_dadda_pg_rca32_nand_31_24_a_31;
  wire f_s_dadda_pg_rca32_nand_31_24_b_24;
  wire f_s_dadda_pg_rca32_nand_31_24_y0;
  wire f_s_dadda_pg_rca32_and_30_25_a_30;
  wire f_s_dadda_pg_rca32_and_30_25_b_25;
  wire f_s_dadda_pg_rca32_and_30_25_y0;
  wire f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_fa666_y4;
  wire f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_nand_31_24_y0;
  wire f_s_dadda_pg_rca32_fa671_y0;
  wire f_s_dadda_pg_rca32_fa671_y1;
  wire f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_and_30_25_y0;
  wire f_s_dadda_pg_rca32_fa671_y2;
  wire f_s_dadda_pg_rca32_fa671_y3;
  wire f_s_dadda_pg_rca32_fa671_y4;
  wire f_s_dadda_pg_rca32_and_29_26_a_29;
  wire f_s_dadda_pg_rca32_and_29_26_b_26;
  wire f_s_dadda_pg_rca32_and_29_26_y0;
  wire f_s_dadda_pg_rca32_and_28_27_a_28;
  wire f_s_dadda_pg_rca32_and_28_27_b_27;
  wire f_s_dadda_pg_rca32_and_28_27_y0;
  wire f_s_dadda_pg_rca32_and_27_28_a_27;
  wire f_s_dadda_pg_rca32_and_27_28_b_28;
  wire f_s_dadda_pg_rca32_and_27_28_y0;
  wire f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_29_26_y0;
  wire f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_28_27_y0;
  wire f_s_dadda_pg_rca32_fa672_y0;
  wire f_s_dadda_pg_rca32_fa672_y1;
  wire f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_27_28_y0;
  wire f_s_dadda_pg_rca32_fa672_y2;
  wire f_s_dadda_pg_rca32_fa672_y3;
  wire f_s_dadda_pg_rca32_fa672_y4;
  wire f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa672_y4;
  wire f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa671_y4;
  wire f_s_dadda_pg_rca32_fa673_y0;
  wire f_s_dadda_pg_rca32_fa673_y1;
  wire f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa670_y4;
  wire f_s_dadda_pg_rca32_fa673_y2;
  wire f_s_dadda_pg_rca32_fa673_y3;
  wire f_s_dadda_pg_rca32_fa673_y4;
  wire f_s_dadda_pg_rca32_nand_31_25_a_31;
  wire f_s_dadda_pg_rca32_nand_31_25_b_25;
  wire f_s_dadda_pg_rca32_nand_31_25_y0;
  wire f_s_dadda_pg_rca32_and_30_26_a_30;
  wire f_s_dadda_pg_rca32_and_30_26_b_26;
  wire f_s_dadda_pg_rca32_and_30_26_y0;
  wire f_s_dadda_pg_rca32_and_29_27_a_29;
  wire f_s_dadda_pg_rca32_and_29_27_b_27;
  wire f_s_dadda_pg_rca32_and_29_27_y0;
  wire f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_nand_31_25_y0;
  wire f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_and_30_26_y0;
  wire f_s_dadda_pg_rca32_fa674_y0;
  wire f_s_dadda_pg_rca32_fa674_y1;
  wire f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_and_29_27_y0;
  wire f_s_dadda_pg_rca32_fa674_y2;
  wire f_s_dadda_pg_rca32_fa674_y3;
  wire f_s_dadda_pg_rca32_fa674_y4;
  wire f_s_dadda_pg_rca32_nand_31_26_a_31;
  wire f_s_dadda_pg_rca32_nand_31_26_b_26;
  wire f_s_dadda_pg_rca32_nand_31_26_y0;
  wire f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_fa674_y4;
  wire f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_fa673_y4;
  wire f_s_dadda_pg_rca32_fa675_y0;
  wire f_s_dadda_pg_rca32_fa675_y1;
  wire f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_nand_31_26_y0;
  wire f_s_dadda_pg_rca32_fa675_y2;
  wire f_s_dadda_pg_rca32_fa675_y3;
  wire f_s_dadda_pg_rca32_fa675_y4;
  wire f_s_dadda_pg_rca32_and_4_0_a_4;
  wire f_s_dadda_pg_rca32_and_4_0_b_0;
  wire f_s_dadda_pg_rca32_and_4_0_y0;
  wire f_s_dadda_pg_rca32_and_3_1_a_3;
  wire f_s_dadda_pg_rca32_and_3_1_b_1;
  wire f_s_dadda_pg_rca32_and_3_1_y0;
  wire f_s_dadda_pg_rca32_ha26_f_s_dadda_pg_rca32_and_4_0_y0;
  wire f_s_dadda_pg_rca32_ha26_f_s_dadda_pg_rca32_and_3_1_y0;
  wire f_s_dadda_pg_rca32_ha26_y0;
  wire f_s_dadda_pg_rca32_ha26_y1;
  wire f_s_dadda_pg_rca32_and_5_0_a_5;
  wire f_s_dadda_pg_rca32_and_5_0_b_0;
  wire f_s_dadda_pg_rca32_and_5_0_y0;
  wire f_s_dadda_pg_rca32_and_4_1_a_4;
  wire f_s_dadda_pg_rca32_and_4_1_b_1;
  wire f_s_dadda_pg_rca32_and_4_1_y0;
  wire f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_ha26_y1;
  wire f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_and_5_0_y0;
  wire f_s_dadda_pg_rca32_fa676_y0;
  wire f_s_dadda_pg_rca32_fa676_y1;
  wire f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_and_4_1_y0;
  wire f_s_dadda_pg_rca32_fa676_y2;
  wire f_s_dadda_pg_rca32_fa676_y3;
  wire f_s_dadda_pg_rca32_fa676_y4;
  wire f_s_dadda_pg_rca32_and_3_2_a_3;
  wire f_s_dadda_pg_rca32_and_3_2_b_2;
  wire f_s_dadda_pg_rca32_and_3_2_y0;
  wire f_s_dadda_pg_rca32_and_2_3_a_2;
  wire f_s_dadda_pg_rca32_and_2_3_b_3;
  wire f_s_dadda_pg_rca32_and_2_3_y0;
  wire f_s_dadda_pg_rca32_ha27_f_s_dadda_pg_rca32_and_3_2_y0;
  wire f_s_dadda_pg_rca32_ha27_f_s_dadda_pg_rca32_and_2_3_y0;
  wire f_s_dadda_pg_rca32_ha27_y0;
  wire f_s_dadda_pg_rca32_ha27_y1;
  wire f_s_dadda_pg_rca32_and_4_2_a_4;
  wire f_s_dadda_pg_rca32_and_4_2_b_2;
  wire f_s_dadda_pg_rca32_and_4_2_y0;
  wire f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_ha27_y1;
  wire f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_fa676_y4;
  wire f_s_dadda_pg_rca32_fa677_y0;
  wire f_s_dadda_pg_rca32_fa677_y1;
  wire f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_and_4_2_y0;
  wire f_s_dadda_pg_rca32_fa677_y2;
  wire f_s_dadda_pg_rca32_fa677_y3;
  wire f_s_dadda_pg_rca32_fa677_y4;
  wire f_s_dadda_pg_rca32_and_3_3_a_3;
  wire f_s_dadda_pg_rca32_and_3_3_b_3;
  wire f_s_dadda_pg_rca32_and_3_3_y0;
  wire f_s_dadda_pg_rca32_and_2_4_a_2;
  wire f_s_dadda_pg_rca32_and_2_4_b_4;
  wire f_s_dadda_pg_rca32_and_2_4_y0;
  wire f_s_dadda_pg_rca32_and_1_5_a_1;
  wire f_s_dadda_pg_rca32_and_1_5_b_5;
  wire f_s_dadda_pg_rca32_and_1_5_y0;
  wire f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_3_3_y0;
  wire f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_2_4_y0;
  wire f_s_dadda_pg_rca32_fa678_y0;
  wire f_s_dadda_pg_rca32_fa678_y1;
  wire f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_1_5_y0;
  wire f_s_dadda_pg_rca32_fa678_y2;
  wire f_s_dadda_pg_rca32_fa678_y3;
  wire f_s_dadda_pg_rca32_fa678_y4;
  wire f_s_dadda_pg_rca32_and_3_4_a_3;
  wire f_s_dadda_pg_rca32_and_3_4_b_4;
  wire f_s_dadda_pg_rca32_and_3_4_y0;
  wire f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_fa678_y4;
  wire f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_fa677_y4;
  wire f_s_dadda_pg_rca32_fa679_y0;
  wire f_s_dadda_pg_rca32_fa679_y1;
  wire f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_and_3_4_y0;
  wire f_s_dadda_pg_rca32_fa679_y2;
  wire f_s_dadda_pg_rca32_fa679_y3;
  wire f_s_dadda_pg_rca32_fa679_y4;
  wire f_s_dadda_pg_rca32_and_2_5_a_2;
  wire f_s_dadda_pg_rca32_and_2_5_b_5;
  wire f_s_dadda_pg_rca32_and_2_5_y0;
  wire f_s_dadda_pg_rca32_and_1_6_a_1;
  wire f_s_dadda_pg_rca32_and_1_6_b_6;
  wire f_s_dadda_pg_rca32_and_1_6_y0;
  wire f_s_dadda_pg_rca32_and_0_7_a_0;
  wire f_s_dadda_pg_rca32_and_0_7_b_7;
  wire f_s_dadda_pg_rca32_and_0_7_y0;
  wire f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_2_5_y0;
  wire f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_1_6_y0;
  wire f_s_dadda_pg_rca32_fa680_y0;
  wire f_s_dadda_pg_rca32_fa680_y1;
  wire f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_0_7_y0;
  wire f_s_dadda_pg_rca32_fa680_y2;
  wire f_s_dadda_pg_rca32_fa680_y3;
  wire f_s_dadda_pg_rca32_fa680_y4;
  wire f_s_dadda_pg_rca32_and_2_6_a_2;
  wire f_s_dadda_pg_rca32_and_2_6_b_6;
  wire f_s_dadda_pg_rca32_and_2_6_y0;
  wire f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_fa680_y4;
  wire f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_fa679_y4;
  wire f_s_dadda_pg_rca32_fa681_y0;
  wire f_s_dadda_pg_rca32_fa681_y1;
  wire f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_and_2_6_y0;
  wire f_s_dadda_pg_rca32_fa681_y2;
  wire f_s_dadda_pg_rca32_fa681_y3;
  wire f_s_dadda_pg_rca32_fa681_y4;
  wire f_s_dadda_pg_rca32_and_1_7_a_1;
  wire f_s_dadda_pg_rca32_and_1_7_b_7;
  wire f_s_dadda_pg_rca32_and_1_7_y0;
  wire f_s_dadda_pg_rca32_and_0_8_a_0;
  wire f_s_dadda_pg_rca32_and_0_8_b_8;
  wire f_s_dadda_pg_rca32_and_0_8_y0;
  wire f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_and_1_7_y0;
  wire f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_and_0_8_y0;
  wire f_s_dadda_pg_rca32_fa682_y0;
  wire f_s_dadda_pg_rca32_fa682_y1;
  wire f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_fa17_y2;
  wire f_s_dadda_pg_rca32_fa682_y2;
  wire f_s_dadda_pg_rca32_fa682_y3;
  wire f_s_dadda_pg_rca32_fa682_y4;
  wire f_s_dadda_pg_rca32_and_1_8_a_1;
  wire f_s_dadda_pg_rca32_and_1_8_b_8;
  wire f_s_dadda_pg_rca32_and_1_8_y0;
  wire f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_fa682_y4;
  wire f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_fa681_y4;
  wire f_s_dadda_pg_rca32_fa683_y0;
  wire f_s_dadda_pg_rca32_fa683_y1;
  wire f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_and_1_8_y0;
  wire f_s_dadda_pg_rca32_fa683_y2;
  wire f_s_dadda_pg_rca32_fa683_y3;
  wire f_s_dadda_pg_rca32_fa683_y4;
  wire f_s_dadda_pg_rca32_and_0_9_a_0;
  wire f_s_dadda_pg_rca32_and_0_9_b_9;
  wire f_s_dadda_pg_rca32_and_0_9_y0;
  wire f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_and_0_9_y0;
  wire f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_fa19_y2;
  wire f_s_dadda_pg_rca32_fa684_y0;
  wire f_s_dadda_pg_rca32_fa684_y1;
  wire f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_fa20_y2;
  wire f_s_dadda_pg_rca32_fa684_y2;
  wire f_s_dadda_pg_rca32_fa684_y3;
  wire f_s_dadda_pg_rca32_fa684_y4;
  wire f_s_dadda_pg_rca32_and_0_10_a_0;
  wire f_s_dadda_pg_rca32_and_0_10_b_10;
  wire f_s_dadda_pg_rca32_and_0_10_y0;
  wire f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_fa684_y4;
  wire f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_fa683_y4;
  wire f_s_dadda_pg_rca32_fa685_y0;
  wire f_s_dadda_pg_rca32_fa685_y1;
  wire f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_and_0_10_y0;
  wire f_s_dadda_pg_rca32_fa685_y2;
  wire f_s_dadda_pg_rca32_fa685_y3;
  wire f_s_dadda_pg_rca32_fa685_y4;
  wire f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa22_y2;
  wire f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa23_y2;
  wire f_s_dadda_pg_rca32_fa686_y0;
  wire f_s_dadda_pg_rca32_fa686_y1;
  wire f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa24_y2;
  wire f_s_dadda_pg_rca32_fa686_y2;
  wire f_s_dadda_pg_rca32_fa686_y3;
  wire f_s_dadda_pg_rca32_fa686_y4;
  wire f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa686_y4;
  wire f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa685_y4;
  wire f_s_dadda_pg_rca32_fa687_y0;
  wire f_s_dadda_pg_rca32_fa687_y1;
  wire f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa26_y2;
  wire f_s_dadda_pg_rca32_fa687_y2;
  wire f_s_dadda_pg_rca32_fa687_y3;
  wire f_s_dadda_pg_rca32_fa687_y4;
  wire f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa27_y2;
  wire f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa28_y2;
  wire f_s_dadda_pg_rca32_fa688_y0;
  wire f_s_dadda_pg_rca32_fa688_y1;
  wire f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa29_y2;
  wire f_s_dadda_pg_rca32_fa688_y2;
  wire f_s_dadda_pg_rca32_fa688_y3;
  wire f_s_dadda_pg_rca32_fa688_y4;
  wire f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa688_y4;
  wire f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa687_y4;
  wire f_s_dadda_pg_rca32_fa689_y0;
  wire f_s_dadda_pg_rca32_fa689_y1;
  wire f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa32_y2;
  wire f_s_dadda_pg_rca32_fa689_y2;
  wire f_s_dadda_pg_rca32_fa689_y3;
  wire f_s_dadda_pg_rca32_fa689_y4;
  wire f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa33_y2;
  wire f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa34_y2;
  wire f_s_dadda_pg_rca32_fa690_y0;
  wire f_s_dadda_pg_rca32_fa690_y1;
  wire f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa35_y2;
  wire f_s_dadda_pg_rca32_fa690_y2;
  wire f_s_dadda_pg_rca32_fa690_y3;
  wire f_s_dadda_pg_rca32_fa690_y4;
  wire f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa690_y4;
  wire f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa689_y4;
  wire f_s_dadda_pg_rca32_fa691_y0;
  wire f_s_dadda_pg_rca32_fa691_y1;
  wire f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa39_y2;
  wire f_s_dadda_pg_rca32_fa691_y2;
  wire f_s_dadda_pg_rca32_fa691_y3;
  wire f_s_dadda_pg_rca32_fa691_y4;
  wire f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa40_y2;
  wire f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa41_y2;
  wire f_s_dadda_pg_rca32_fa692_y0;
  wire f_s_dadda_pg_rca32_fa692_y1;
  wire f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa42_y2;
  wire f_s_dadda_pg_rca32_fa692_y2;
  wire f_s_dadda_pg_rca32_fa692_y3;
  wire f_s_dadda_pg_rca32_fa692_y4;
  wire f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa692_y4;
  wire f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa691_y4;
  wire f_s_dadda_pg_rca32_fa693_y0;
  wire f_s_dadda_pg_rca32_fa693_y1;
  wire f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa47_y2;
  wire f_s_dadda_pg_rca32_fa693_y2;
  wire f_s_dadda_pg_rca32_fa693_y3;
  wire f_s_dadda_pg_rca32_fa693_y4;
  wire f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa48_y2;
  wire f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa49_y2;
  wire f_s_dadda_pg_rca32_fa694_y0;
  wire f_s_dadda_pg_rca32_fa694_y1;
  wire f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa50_y2;
  wire f_s_dadda_pg_rca32_fa694_y2;
  wire f_s_dadda_pg_rca32_fa694_y3;
  wire f_s_dadda_pg_rca32_fa694_y4;
  wire f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa694_y4;
  wire f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa693_y4;
  wire f_s_dadda_pg_rca32_fa695_y0;
  wire f_s_dadda_pg_rca32_fa695_y1;
  wire f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa56_y2;
  wire f_s_dadda_pg_rca32_fa695_y2;
  wire f_s_dadda_pg_rca32_fa695_y3;
  wire f_s_dadda_pg_rca32_fa695_y4;
  wire f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa57_y2;
  wire f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa58_y2;
  wire f_s_dadda_pg_rca32_fa696_y0;
  wire f_s_dadda_pg_rca32_fa696_y1;
  wire f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa59_y2;
  wire f_s_dadda_pg_rca32_fa696_y2;
  wire f_s_dadda_pg_rca32_fa696_y3;
  wire f_s_dadda_pg_rca32_fa696_y4;
  wire f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa696_y4;
  wire f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa695_y4;
  wire f_s_dadda_pg_rca32_fa697_y0;
  wire f_s_dadda_pg_rca32_fa697_y1;
  wire f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa66_y2;
  wire f_s_dadda_pg_rca32_fa697_y2;
  wire f_s_dadda_pg_rca32_fa697_y3;
  wire f_s_dadda_pg_rca32_fa697_y4;
  wire f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa67_y2;
  wire f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa68_y2;
  wire f_s_dadda_pg_rca32_fa698_y0;
  wire f_s_dadda_pg_rca32_fa698_y1;
  wire f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa69_y2;
  wire f_s_dadda_pg_rca32_fa698_y2;
  wire f_s_dadda_pg_rca32_fa698_y3;
  wire f_s_dadda_pg_rca32_fa698_y4;
  wire f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa698_y4;
  wire f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa697_y4;
  wire f_s_dadda_pg_rca32_fa699_y0;
  wire f_s_dadda_pg_rca32_fa699_y1;
  wire f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa77_y2;
  wire f_s_dadda_pg_rca32_fa699_y2;
  wire f_s_dadda_pg_rca32_fa699_y3;
  wire f_s_dadda_pg_rca32_fa699_y4;
  wire f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa78_y2;
  wire f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa79_y2;
  wire f_s_dadda_pg_rca32_fa700_y0;
  wire f_s_dadda_pg_rca32_fa700_y1;
  wire f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa80_y2;
  wire f_s_dadda_pg_rca32_fa700_y2;
  wire f_s_dadda_pg_rca32_fa700_y3;
  wire f_s_dadda_pg_rca32_fa700_y4;
  wire f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa700_y4;
  wire f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa699_y4;
  wire f_s_dadda_pg_rca32_fa701_y0;
  wire f_s_dadda_pg_rca32_fa701_y1;
  wire f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa89_y2;
  wire f_s_dadda_pg_rca32_fa701_y2;
  wire f_s_dadda_pg_rca32_fa701_y3;
  wire f_s_dadda_pg_rca32_fa701_y4;
  wire f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa90_y2;
  wire f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa91_y2;
  wire f_s_dadda_pg_rca32_fa702_y0;
  wire f_s_dadda_pg_rca32_fa702_y1;
  wire f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa92_y2;
  wire f_s_dadda_pg_rca32_fa702_y2;
  wire f_s_dadda_pg_rca32_fa702_y3;
  wire f_s_dadda_pg_rca32_fa702_y4;
  wire f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa702_y4;
  wire f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa701_y4;
  wire f_s_dadda_pg_rca32_fa703_y0;
  wire f_s_dadda_pg_rca32_fa703_y1;
  wire f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa102_y2;
  wire f_s_dadda_pg_rca32_fa703_y2;
  wire f_s_dadda_pg_rca32_fa703_y3;
  wire f_s_dadda_pg_rca32_fa703_y4;
  wire f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa103_y2;
  wire f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa104_y2;
  wire f_s_dadda_pg_rca32_fa704_y0;
  wire f_s_dadda_pg_rca32_fa704_y1;
  wire f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa105_y2;
  wire f_s_dadda_pg_rca32_fa704_y2;
  wire f_s_dadda_pg_rca32_fa704_y3;
  wire f_s_dadda_pg_rca32_fa704_y4;
  wire f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa704_y4;
  wire f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa703_y4;
  wire f_s_dadda_pg_rca32_fa705_y0;
  wire f_s_dadda_pg_rca32_fa705_y1;
  wire f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa116_y2;
  wire f_s_dadda_pg_rca32_fa705_y2;
  wire f_s_dadda_pg_rca32_fa705_y3;
  wire f_s_dadda_pg_rca32_fa705_y4;
  wire f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa117_y2;
  wire f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa118_y2;
  wire f_s_dadda_pg_rca32_fa706_y0;
  wire f_s_dadda_pg_rca32_fa706_y1;
  wire f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa119_y2;
  wire f_s_dadda_pg_rca32_fa706_y2;
  wire f_s_dadda_pg_rca32_fa706_y3;
  wire f_s_dadda_pg_rca32_fa706_y4;
  wire f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa706_y4;
  wire f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa705_y4;
  wire f_s_dadda_pg_rca32_fa707_y0;
  wire f_s_dadda_pg_rca32_fa707_y1;
  wire f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa131_y2;
  wire f_s_dadda_pg_rca32_fa707_y2;
  wire f_s_dadda_pg_rca32_fa707_y3;
  wire f_s_dadda_pg_rca32_fa707_y4;
  wire f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa132_y2;
  wire f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa133_y2;
  wire f_s_dadda_pg_rca32_fa708_y0;
  wire f_s_dadda_pg_rca32_fa708_y1;
  wire f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa134_y2;
  wire f_s_dadda_pg_rca32_fa708_y2;
  wire f_s_dadda_pg_rca32_fa708_y3;
  wire f_s_dadda_pg_rca32_fa708_y4;
  wire f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa708_y4;
  wire f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa707_y4;
  wire f_s_dadda_pg_rca32_fa709_y0;
  wire f_s_dadda_pg_rca32_fa709_y1;
  wire f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa147_y2;
  wire f_s_dadda_pg_rca32_fa709_y2;
  wire f_s_dadda_pg_rca32_fa709_y3;
  wire f_s_dadda_pg_rca32_fa709_y4;
  wire f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa148_y2;
  wire f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa149_y2;
  wire f_s_dadda_pg_rca32_fa710_y0;
  wire f_s_dadda_pg_rca32_fa710_y1;
  wire f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa150_y2;
  wire f_s_dadda_pg_rca32_fa710_y2;
  wire f_s_dadda_pg_rca32_fa710_y3;
  wire f_s_dadda_pg_rca32_fa710_y4;
  wire f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa710_y4;
  wire f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa709_y4;
  wire f_s_dadda_pg_rca32_fa711_y0;
  wire f_s_dadda_pg_rca32_fa711_y1;
  wire f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa164_y2;
  wire f_s_dadda_pg_rca32_fa711_y2;
  wire f_s_dadda_pg_rca32_fa711_y3;
  wire f_s_dadda_pg_rca32_fa711_y4;
  wire f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa165_y2;
  wire f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa166_y2;
  wire f_s_dadda_pg_rca32_fa712_y0;
  wire f_s_dadda_pg_rca32_fa712_y1;
  wire f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa167_y2;
  wire f_s_dadda_pg_rca32_fa712_y2;
  wire f_s_dadda_pg_rca32_fa712_y3;
  wire f_s_dadda_pg_rca32_fa712_y4;
  wire f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa712_y4;
  wire f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa711_y4;
  wire f_s_dadda_pg_rca32_fa713_y0;
  wire f_s_dadda_pg_rca32_fa713_y1;
  wire f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa182_y2;
  wire f_s_dadda_pg_rca32_fa713_y2;
  wire f_s_dadda_pg_rca32_fa713_y3;
  wire f_s_dadda_pg_rca32_fa713_y4;
  wire f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa183_y2;
  wire f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa184_y2;
  wire f_s_dadda_pg_rca32_fa714_y0;
  wire f_s_dadda_pg_rca32_fa714_y1;
  wire f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa185_y2;
  wire f_s_dadda_pg_rca32_fa714_y2;
  wire f_s_dadda_pg_rca32_fa714_y3;
  wire f_s_dadda_pg_rca32_fa714_y4;
  wire f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa714_y4;
  wire f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa713_y4;
  wire f_s_dadda_pg_rca32_fa715_y0;
  wire f_s_dadda_pg_rca32_fa715_y1;
  wire f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa201_y2;
  wire f_s_dadda_pg_rca32_fa715_y2;
  wire f_s_dadda_pg_rca32_fa715_y3;
  wire f_s_dadda_pg_rca32_fa715_y4;
  wire f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa202_y2;
  wire f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa203_y2;
  wire f_s_dadda_pg_rca32_fa716_y0;
  wire f_s_dadda_pg_rca32_fa716_y1;
  wire f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa204_y2;
  wire f_s_dadda_pg_rca32_fa716_y2;
  wire f_s_dadda_pg_rca32_fa716_y3;
  wire f_s_dadda_pg_rca32_fa716_y4;
  wire f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa716_y4;
  wire f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa715_y4;
  wire f_s_dadda_pg_rca32_fa717_y0;
  wire f_s_dadda_pg_rca32_fa717_y1;
  wire f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa221_y2;
  wire f_s_dadda_pg_rca32_fa717_y2;
  wire f_s_dadda_pg_rca32_fa717_y3;
  wire f_s_dadda_pg_rca32_fa717_y4;
  wire f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa222_y2;
  wire f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa223_y2;
  wire f_s_dadda_pg_rca32_fa718_y0;
  wire f_s_dadda_pg_rca32_fa718_y1;
  wire f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa224_y2;
  wire f_s_dadda_pg_rca32_fa718_y2;
  wire f_s_dadda_pg_rca32_fa718_y3;
  wire f_s_dadda_pg_rca32_fa718_y4;
  wire f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa718_y4;
  wire f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa717_y4;
  wire f_s_dadda_pg_rca32_fa719_y0;
  wire f_s_dadda_pg_rca32_fa719_y1;
  wire f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa242_y2;
  wire f_s_dadda_pg_rca32_fa719_y2;
  wire f_s_dadda_pg_rca32_fa719_y3;
  wire f_s_dadda_pg_rca32_fa719_y4;
  wire f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa243_y2;
  wire f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa244_y2;
  wire f_s_dadda_pg_rca32_fa720_y0;
  wire f_s_dadda_pg_rca32_fa720_y1;
  wire f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa245_y2;
  wire f_s_dadda_pg_rca32_fa720_y2;
  wire f_s_dadda_pg_rca32_fa720_y3;
  wire f_s_dadda_pg_rca32_fa720_y4;
  wire f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa720_y4;
  wire f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa719_y4;
  wire f_s_dadda_pg_rca32_fa721_y0;
  wire f_s_dadda_pg_rca32_fa721_y1;
  wire f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa263_y2;
  wire f_s_dadda_pg_rca32_fa721_y2;
  wire f_s_dadda_pg_rca32_fa721_y3;
  wire f_s_dadda_pg_rca32_fa721_y4;
  wire f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa264_y2;
  wire f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa265_y2;
  wire f_s_dadda_pg_rca32_fa722_y0;
  wire f_s_dadda_pg_rca32_fa722_y1;
  wire f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa266_y2;
  wire f_s_dadda_pg_rca32_fa722_y2;
  wire f_s_dadda_pg_rca32_fa722_y3;
  wire f_s_dadda_pg_rca32_fa722_y4;
  wire f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa722_y4;
  wire f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa721_y4;
  wire f_s_dadda_pg_rca32_fa723_y0;
  wire f_s_dadda_pg_rca32_fa723_y1;
  wire f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa285_y2;
  wire f_s_dadda_pg_rca32_fa723_y2;
  wire f_s_dadda_pg_rca32_fa723_y3;
  wire f_s_dadda_pg_rca32_fa723_y4;
  wire f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa286_y2;
  wire f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa287_y2;
  wire f_s_dadda_pg_rca32_fa724_y0;
  wire f_s_dadda_pg_rca32_fa724_y1;
  wire f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa288_y2;
  wire f_s_dadda_pg_rca32_fa724_y2;
  wire f_s_dadda_pg_rca32_fa724_y3;
  wire f_s_dadda_pg_rca32_fa724_y4;
  wire f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa724_y4;
  wire f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa723_y4;
  wire f_s_dadda_pg_rca32_fa725_y0;
  wire f_s_dadda_pg_rca32_fa725_y1;
  wire f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa307_y2;
  wire f_s_dadda_pg_rca32_fa725_y2;
  wire f_s_dadda_pg_rca32_fa725_y3;
  wire f_s_dadda_pg_rca32_fa725_y4;
  wire f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa308_y2;
  wire f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa309_y2;
  wire f_s_dadda_pg_rca32_fa726_y0;
  wire f_s_dadda_pg_rca32_fa726_y1;
  wire f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa310_y2;
  wire f_s_dadda_pg_rca32_fa726_y2;
  wire f_s_dadda_pg_rca32_fa726_y3;
  wire f_s_dadda_pg_rca32_fa726_y4;
  wire f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa726_y4;
  wire f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa725_y4;
  wire f_s_dadda_pg_rca32_fa727_y0;
  wire f_s_dadda_pg_rca32_fa727_y1;
  wire f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa329_y2;
  wire f_s_dadda_pg_rca32_fa727_y2;
  wire f_s_dadda_pg_rca32_fa727_y3;
  wire f_s_dadda_pg_rca32_fa727_y4;
  wire f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa330_y2;
  wire f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa331_y2;
  wire f_s_dadda_pg_rca32_fa728_y0;
  wire f_s_dadda_pg_rca32_fa728_y1;
  wire f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa332_y2;
  wire f_s_dadda_pg_rca32_fa728_y2;
  wire f_s_dadda_pg_rca32_fa728_y3;
  wire f_s_dadda_pg_rca32_fa728_y4;
  wire f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa728_y4;
  wire f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa727_y4;
  wire f_s_dadda_pg_rca32_fa729_y0;
  wire f_s_dadda_pg_rca32_fa729_y1;
  wire f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa351_y2;
  wire f_s_dadda_pg_rca32_fa729_y2;
  wire f_s_dadda_pg_rca32_fa729_y3;
  wire f_s_dadda_pg_rca32_fa729_y4;
  wire f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa352_y2;
  wire f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa353_y2;
  wire f_s_dadda_pg_rca32_fa730_y0;
  wire f_s_dadda_pg_rca32_fa730_y1;
  wire f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa354_y2;
  wire f_s_dadda_pg_rca32_fa730_y2;
  wire f_s_dadda_pg_rca32_fa730_y3;
  wire f_s_dadda_pg_rca32_fa730_y4;
  wire f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa730_y4;
  wire f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa729_y4;
  wire f_s_dadda_pg_rca32_fa731_y0;
  wire f_s_dadda_pg_rca32_fa731_y1;
  wire f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa373_y2;
  wire f_s_dadda_pg_rca32_fa731_y2;
  wire f_s_dadda_pg_rca32_fa731_y3;
  wire f_s_dadda_pg_rca32_fa731_y4;
  wire f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa374_y2;
  wire f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa375_y2;
  wire f_s_dadda_pg_rca32_fa732_y0;
  wire f_s_dadda_pg_rca32_fa732_y1;
  wire f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa376_y2;
  wire f_s_dadda_pg_rca32_fa732_y2;
  wire f_s_dadda_pg_rca32_fa732_y3;
  wire f_s_dadda_pg_rca32_fa732_y4;
  wire f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa732_y4;
  wire f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa731_y4;
  wire f_s_dadda_pg_rca32_fa733_y0;
  wire f_s_dadda_pg_rca32_fa733_y1;
  wire f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa395_y2;
  wire f_s_dadda_pg_rca32_fa733_y2;
  wire f_s_dadda_pg_rca32_fa733_y3;
  wire f_s_dadda_pg_rca32_fa733_y4;
  wire f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa396_y2;
  wire f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa397_y2;
  wire f_s_dadda_pg_rca32_fa734_y0;
  wire f_s_dadda_pg_rca32_fa734_y1;
  wire f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa398_y2;
  wire f_s_dadda_pg_rca32_fa734_y2;
  wire f_s_dadda_pg_rca32_fa734_y3;
  wire f_s_dadda_pg_rca32_fa734_y4;
  wire f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa734_y4;
  wire f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa733_y4;
  wire f_s_dadda_pg_rca32_fa735_y0;
  wire f_s_dadda_pg_rca32_fa735_y1;
  wire f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa417_y2;
  wire f_s_dadda_pg_rca32_fa735_y2;
  wire f_s_dadda_pg_rca32_fa735_y3;
  wire f_s_dadda_pg_rca32_fa735_y4;
  wire f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa418_y2;
  wire f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa419_y2;
  wire f_s_dadda_pg_rca32_fa736_y0;
  wire f_s_dadda_pg_rca32_fa736_y1;
  wire f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa420_y2;
  wire f_s_dadda_pg_rca32_fa736_y2;
  wire f_s_dadda_pg_rca32_fa736_y3;
  wire f_s_dadda_pg_rca32_fa736_y4;
  wire f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa736_y4;
  wire f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa735_y4;
  wire f_s_dadda_pg_rca32_fa737_y0;
  wire f_s_dadda_pg_rca32_fa737_y1;
  wire f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa439_y2;
  wire f_s_dadda_pg_rca32_fa737_y2;
  wire f_s_dadda_pg_rca32_fa737_y3;
  wire f_s_dadda_pg_rca32_fa737_y4;
  wire f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa440_y2;
  wire f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa441_y2;
  wire f_s_dadda_pg_rca32_fa738_y0;
  wire f_s_dadda_pg_rca32_fa738_y1;
  wire f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa442_y2;
  wire f_s_dadda_pg_rca32_fa738_y2;
  wire f_s_dadda_pg_rca32_fa738_y3;
  wire f_s_dadda_pg_rca32_fa738_y4;
  wire f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa738_y4;
  wire f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa737_y4;
  wire f_s_dadda_pg_rca32_fa739_y0;
  wire f_s_dadda_pg_rca32_fa739_y1;
  wire f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa460_y2;
  wire f_s_dadda_pg_rca32_fa739_y2;
  wire f_s_dadda_pg_rca32_fa739_y3;
  wire f_s_dadda_pg_rca32_fa739_y4;
  wire f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa461_y2;
  wire f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa462_y2;
  wire f_s_dadda_pg_rca32_fa740_y0;
  wire f_s_dadda_pg_rca32_fa740_y1;
  wire f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa463_y2;
  wire f_s_dadda_pg_rca32_fa740_y2;
  wire f_s_dadda_pg_rca32_fa740_y3;
  wire f_s_dadda_pg_rca32_fa740_y4;
  wire f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa740_y4;
  wire f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa739_y4;
  wire f_s_dadda_pg_rca32_fa741_y0;
  wire f_s_dadda_pg_rca32_fa741_y1;
  wire f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa480_y2;
  wire f_s_dadda_pg_rca32_fa741_y2;
  wire f_s_dadda_pg_rca32_fa741_y3;
  wire f_s_dadda_pg_rca32_fa741_y4;
  wire f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa481_y2;
  wire f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa482_y2;
  wire f_s_dadda_pg_rca32_fa742_y0;
  wire f_s_dadda_pg_rca32_fa742_y1;
  wire f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa483_y2;
  wire f_s_dadda_pg_rca32_fa742_y2;
  wire f_s_dadda_pg_rca32_fa742_y3;
  wire f_s_dadda_pg_rca32_fa742_y4;
  wire f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa742_y4;
  wire f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa741_y4;
  wire f_s_dadda_pg_rca32_fa743_y0;
  wire f_s_dadda_pg_rca32_fa743_y1;
  wire f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa499_y2;
  wire f_s_dadda_pg_rca32_fa743_y2;
  wire f_s_dadda_pg_rca32_fa743_y3;
  wire f_s_dadda_pg_rca32_fa743_y4;
  wire f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa500_y2;
  wire f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa501_y2;
  wire f_s_dadda_pg_rca32_fa744_y0;
  wire f_s_dadda_pg_rca32_fa744_y1;
  wire f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa502_y2;
  wire f_s_dadda_pg_rca32_fa744_y2;
  wire f_s_dadda_pg_rca32_fa744_y3;
  wire f_s_dadda_pg_rca32_fa744_y4;
  wire f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa744_y4;
  wire f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa743_y4;
  wire f_s_dadda_pg_rca32_fa745_y0;
  wire f_s_dadda_pg_rca32_fa745_y1;
  wire f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa517_y2;
  wire f_s_dadda_pg_rca32_fa745_y2;
  wire f_s_dadda_pg_rca32_fa745_y3;
  wire f_s_dadda_pg_rca32_fa745_y4;
  wire f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa518_y2;
  wire f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa519_y2;
  wire f_s_dadda_pg_rca32_fa746_y0;
  wire f_s_dadda_pg_rca32_fa746_y1;
  wire f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa520_y2;
  wire f_s_dadda_pg_rca32_fa746_y2;
  wire f_s_dadda_pg_rca32_fa746_y3;
  wire f_s_dadda_pg_rca32_fa746_y4;
  wire f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa746_y4;
  wire f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa745_y4;
  wire f_s_dadda_pg_rca32_fa747_y0;
  wire f_s_dadda_pg_rca32_fa747_y1;
  wire f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa534_y2;
  wire f_s_dadda_pg_rca32_fa747_y2;
  wire f_s_dadda_pg_rca32_fa747_y3;
  wire f_s_dadda_pg_rca32_fa747_y4;
  wire f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa535_y2;
  wire f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa536_y2;
  wire f_s_dadda_pg_rca32_fa748_y0;
  wire f_s_dadda_pg_rca32_fa748_y1;
  wire f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa537_y2;
  wire f_s_dadda_pg_rca32_fa748_y2;
  wire f_s_dadda_pg_rca32_fa748_y3;
  wire f_s_dadda_pg_rca32_fa748_y4;
  wire f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa748_y4;
  wire f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa747_y4;
  wire f_s_dadda_pg_rca32_fa749_y0;
  wire f_s_dadda_pg_rca32_fa749_y1;
  wire f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa550_y2;
  wire f_s_dadda_pg_rca32_fa749_y2;
  wire f_s_dadda_pg_rca32_fa749_y3;
  wire f_s_dadda_pg_rca32_fa749_y4;
  wire f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa551_y2;
  wire f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa552_y2;
  wire f_s_dadda_pg_rca32_fa750_y0;
  wire f_s_dadda_pg_rca32_fa750_y1;
  wire f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa553_y2;
  wire f_s_dadda_pg_rca32_fa750_y2;
  wire f_s_dadda_pg_rca32_fa750_y3;
  wire f_s_dadda_pg_rca32_fa750_y4;
  wire f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa750_y4;
  wire f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa749_y4;
  wire f_s_dadda_pg_rca32_fa751_y0;
  wire f_s_dadda_pg_rca32_fa751_y1;
  wire f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa565_y2;
  wire f_s_dadda_pg_rca32_fa751_y2;
  wire f_s_dadda_pg_rca32_fa751_y3;
  wire f_s_dadda_pg_rca32_fa751_y4;
  wire f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa566_y2;
  wire f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa567_y2;
  wire f_s_dadda_pg_rca32_fa752_y0;
  wire f_s_dadda_pg_rca32_fa752_y1;
  wire f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa568_y2;
  wire f_s_dadda_pg_rca32_fa752_y2;
  wire f_s_dadda_pg_rca32_fa752_y3;
  wire f_s_dadda_pg_rca32_fa752_y4;
  wire f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa752_y4;
  wire f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa751_y4;
  wire f_s_dadda_pg_rca32_fa753_y0;
  wire f_s_dadda_pg_rca32_fa753_y1;
  wire f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa579_y2;
  wire f_s_dadda_pg_rca32_fa753_y2;
  wire f_s_dadda_pg_rca32_fa753_y3;
  wire f_s_dadda_pg_rca32_fa753_y4;
  wire f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa580_y2;
  wire f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa581_y2;
  wire f_s_dadda_pg_rca32_fa754_y0;
  wire f_s_dadda_pg_rca32_fa754_y1;
  wire f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa582_y2;
  wire f_s_dadda_pg_rca32_fa754_y2;
  wire f_s_dadda_pg_rca32_fa754_y3;
  wire f_s_dadda_pg_rca32_fa754_y4;
  wire f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa754_y4;
  wire f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa753_y4;
  wire f_s_dadda_pg_rca32_fa755_y0;
  wire f_s_dadda_pg_rca32_fa755_y1;
  wire f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa592_y2;
  wire f_s_dadda_pg_rca32_fa755_y2;
  wire f_s_dadda_pg_rca32_fa755_y3;
  wire f_s_dadda_pg_rca32_fa755_y4;
  wire f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa593_y2;
  wire f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa594_y2;
  wire f_s_dadda_pg_rca32_fa756_y0;
  wire f_s_dadda_pg_rca32_fa756_y1;
  wire f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa595_y2;
  wire f_s_dadda_pg_rca32_fa756_y2;
  wire f_s_dadda_pg_rca32_fa756_y3;
  wire f_s_dadda_pg_rca32_fa756_y4;
  wire f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa756_y4;
  wire f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa755_y4;
  wire f_s_dadda_pg_rca32_fa757_y0;
  wire f_s_dadda_pg_rca32_fa757_y1;
  wire f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa604_y2;
  wire f_s_dadda_pg_rca32_fa757_y2;
  wire f_s_dadda_pg_rca32_fa757_y3;
  wire f_s_dadda_pg_rca32_fa757_y4;
  wire f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa605_y2;
  wire f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa606_y2;
  wire f_s_dadda_pg_rca32_fa758_y0;
  wire f_s_dadda_pg_rca32_fa758_y1;
  wire f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa607_y2;
  wire f_s_dadda_pg_rca32_fa758_y2;
  wire f_s_dadda_pg_rca32_fa758_y3;
  wire f_s_dadda_pg_rca32_fa758_y4;
  wire f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa758_y4;
  wire f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa757_y4;
  wire f_s_dadda_pg_rca32_fa759_y0;
  wire f_s_dadda_pg_rca32_fa759_y1;
  wire f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa615_y2;
  wire f_s_dadda_pg_rca32_fa759_y2;
  wire f_s_dadda_pg_rca32_fa759_y3;
  wire f_s_dadda_pg_rca32_fa759_y4;
  wire f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa616_y2;
  wire f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa617_y2;
  wire f_s_dadda_pg_rca32_fa760_y0;
  wire f_s_dadda_pg_rca32_fa760_y1;
  wire f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa618_y2;
  wire f_s_dadda_pg_rca32_fa760_y2;
  wire f_s_dadda_pg_rca32_fa760_y3;
  wire f_s_dadda_pg_rca32_fa760_y4;
  wire f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa760_y4;
  wire f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa759_y4;
  wire f_s_dadda_pg_rca32_fa761_y0;
  wire f_s_dadda_pg_rca32_fa761_y1;
  wire f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa625_y2;
  wire f_s_dadda_pg_rca32_fa761_y2;
  wire f_s_dadda_pg_rca32_fa761_y3;
  wire f_s_dadda_pg_rca32_fa761_y4;
  wire f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa626_y2;
  wire f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa627_y2;
  wire f_s_dadda_pg_rca32_fa762_y0;
  wire f_s_dadda_pg_rca32_fa762_y1;
  wire f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa628_y2;
  wire f_s_dadda_pg_rca32_fa762_y2;
  wire f_s_dadda_pg_rca32_fa762_y3;
  wire f_s_dadda_pg_rca32_fa762_y4;
  wire f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa762_y4;
  wire f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa761_y4;
  wire f_s_dadda_pg_rca32_fa763_y0;
  wire f_s_dadda_pg_rca32_fa763_y1;
  wire f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa634_y2;
  wire f_s_dadda_pg_rca32_fa763_y2;
  wire f_s_dadda_pg_rca32_fa763_y3;
  wire f_s_dadda_pg_rca32_fa763_y4;
  wire f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa635_y2;
  wire f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa636_y2;
  wire f_s_dadda_pg_rca32_fa764_y0;
  wire f_s_dadda_pg_rca32_fa764_y1;
  wire f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa637_y2;
  wire f_s_dadda_pg_rca32_fa764_y2;
  wire f_s_dadda_pg_rca32_fa764_y3;
  wire f_s_dadda_pg_rca32_fa764_y4;
  wire f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa764_y4;
  wire f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa763_y4;
  wire f_s_dadda_pg_rca32_fa765_y0;
  wire f_s_dadda_pg_rca32_fa765_y1;
  wire f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa642_y2;
  wire f_s_dadda_pg_rca32_fa765_y2;
  wire f_s_dadda_pg_rca32_fa765_y3;
  wire f_s_dadda_pg_rca32_fa765_y4;
  wire f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa643_y2;
  wire f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa644_y2;
  wire f_s_dadda_pg_rca32_fa766_y0;
  wire f_s_dadda_pg_rca32_fa766_y1;
  wire f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa645_y2;
  wire f_s_dadda_pg_rca32_fa766_y2;
  wire f_s_dadda_pg_rca32_fa766_y3;
  wire f_s_dadda_pg_rca32_fa766_y4;
  wire f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa766_y4;
  wire f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa765_y4;
  wire f_s_dadda_pg_rca32_fa767_y0;
  wire f_s_dadda_pg_rca32_fa767_y1;
  wire f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa649_y2;
  wire f_s_dadda_pg_rca32_fa767_y2;
  wire f_s_dadda_pg_rca32_fa767_y3;
  wire f_s_dadda_pg_rca32_fa767_y4;
  wire f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa650_y2;
  wire f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa651_y2;
  wire f_s_dadda_pg_rca32_fa768_y0;
  wire f_s_dadda_pg_rca32_fa768_y1;
  wire f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa652_y2;
  wire f_s_dadda_pg_rca32_fa768_y2;
  wire f_s_dadda_pg_rca32_fa768_y3;
  wire f_s_dadda_pg_rca32_fa768_y4;
  wire f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa768_y4;
  wire f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa767_y4;
  wire f_s_dadda_pg_rca32_fa769_y0;
  wire f_s_dadda_pg_rca32_fa769_y1;
  wire f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa655_y2;
  wire f_s_dadda_pg_rca32_fa769_y2;
  wire f_s_dadda_pg_rca32_fa769_y3;
  wire f_s_dadda_pg_rca32_fa769_y4;
  wire f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa656_y2;
  wire f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa657_y2;
  wire f_s_dadda_pg_rca32_fa770_y0;
  wire f_s_dadda_pg_rca32_fa770_y1;
  wire f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa658_y2;
  wire f_s_dadda_pg_rca32_fa770_y2;
  wire f_s_dadda_pg_rca32_fa770_y3;
  wire f_s_dadda_pg_rca32_fa770_y4;
  wire f_s_dadda_pg_rca32_nand_22_31_a_22;
  wire f_s_dadda_pg_rca32_nand_22_31_b_31;
  wire f_s_dadda_pg_rca32_nand_22_31_y0;
  wire f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_fa770_y4;
  wire f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_fa769_y4;
  wire f_s_dadda_pg_rca32_fa771_y0;
  wire f_s_dadda_pg_rca32_fa771_y1;
  wire f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_nand_22_31_y0;
  wire f_s_dadda_pg_rca32_fa771_y2;
  wire f_s_dadda_pg_rca32_fa771_y3;
  wire f_s_dadda_pg_rca32_fa771_y4;
  wire f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa661_y2;
  wire f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa662_y2;
  wire f_s_dadda_pg_rca32_fa772_y0;
  wire f_s_dadda_pg_rca32_fa772_y1;
  wire f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa663_y2;
  wire f_s_dadda_pg_rca32_fa772_y2;
  wire f_s_dadda_pg_rca32_fa772_y3;
  wire f_s_dadda_pg_rca32_fa772_y4;
  wire f_s_dadda_pg_rca32_and_24_30_a_24;
  wire f_s_dadda_pg_rca32_and_24_30_b_30;
  wire f_s_dadda_pg_rca32_and_24_30_y0;
  wire f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_fa772_y4;
  wire f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_fa771_y4;
  wire f_s_dadda_pg_rca32_fa773_y0;
  wire f_s_dadda_pg_rca32_fa773_y1;
  wire f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_and_24_30_y0;
  wire f_s_dadda_pg_rca32_fa773_y2;
  wire f_s_dadda_pg_rca32_fa773_y3;
  wire f_s_dadda_pg_rca32_fa773_y4;
  wire f_s_dadda_pg_rca32_nand_23_31_a_23;
  wire f_s_dadda_pg_rca32_nand_23_31_b_31;
  wire f_s_dadda_pg_rca32_nand_23_31_y0;
  wire f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_nand_23_31_y0;
  wire f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_fa666_y2;
  wire f_s_dadda_pg_rca32_fa774_y0;
  wire f_s_dadda_pg_rca32_fa774_y1;
  wire f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_fa667_y2;
  wire f_s_dadda_pg_rca32_fa774_y2;
  wire f_s_dadda_pg_rca32_fa774_y3;
  wire f_s_dadda_pg_rca32_fa774_y4;
  wire f_s_dadda_pg_rca32_and_26_29_a_26;
  wire f_s_dadda_pg_rca32_and_26_29_b_29;
  wire f_s_dadda_pg_rca32_and_26_29_y0;
  wire f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_fa774_y4;
  wire f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_fa773_y4;
  wire f_s_dadda_pg_rca32_fa775_y0;
  wire f_s_dadda_pg_rca32_fa775_y1;
  wire f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_and_26_29_y0;
  wire f_s_dadda_pg_rca32_fa775_y2;
  wire f_s_dadda_pg_rca32_fa775_y3;
  wire f_s_dadda_pg_rca32_fa775_y4;
  wire f_s_dadda_pg_rca32_and_25_30_a_25;
  wire f_s_dadda_pg_rca32_and_25_30_b_30;
  wire f_s_dadda_pg_rca32_and_25_30_y0;
  wire f_s_dadda_pg_rca32_nand_24_31_a_24;
  wire f_s_dadda_pg_rca32_nand_24_31_b_31;
  wire f_s_dadda_pg_rca32_nand_24_31_y0;
  wire f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_and_25_30_y0;
  wire f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_nand_24_31_y0;
  wire f_s_dadda_pg_rca32_fa776_y0;
  wire f_s_dadda_pg_rca32_fa776_y1;
  wire f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_fa670_y2;
  wire f_s_dadda_pg_rca32_fa776_y2;
  wire f_s_dadda_pg_rca32_fa776_y3;
  wire f_s_dadda_pg_rca32_fa776_y4;
  wire f_s_dadda_pg_rca32_and_28_28_a_28;
  wire f_s_dadda_pg_rca32_and_28_28_b_28;
  wire f_s_dadda_pg_rca32_and_28_28_y0;
  wire f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_fa776_y4;
  wire f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_fa775_y4;
  wire f_s_dadda_pg_rca32_fa777_y0;
  wire f_s_dadda_pg_rca32_fa777_y1;
  wire f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_and_28_28_y0;
  wire f_s_dadda_pg_rca32_fa777_y2;
  wire f_s_dadda_pg_rca32_fa777_y3;
  wire f_s_dadda_pg_rca32_fa777_y4;
  wire f_s_dadda_pg_rca32_and_27_29_a_27;
  wire f_s_dadda_pg_rca32_and_27_29_b_29;
  wire f_s_dadda_pg_rca32_and_27_29_y0;
  wire f_s_dadda_pg_rca32_and_26_30_a_26;
  wire f_s_dadda_pg_rca32_and_26_30_b_30;
  wire f_s_dadda_pg_rca32_and_26_30_y0;
  wire f_s_dadda_pg_rca32_nand_25_31_a_25;
  wire f_s_dadda_pg_rca32_nand_25_31_b_31;
  wire f_s_dadda_pg_rca32_nand_25_31_y0;
  wire f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_and_27_29_y0;
  wire f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_and_26_30_y0;
  wire f_s_dadda_pg_rca32_fa778_y0;
  wire f_s_dadda_pg_rca32_fa778_y1;
  wire f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_nand_25_31_y0;
  wire f_s_dadda_pg_rca32_fa778_y2;
  wire f_s_dadda_pg_rca32_fa778_y3;
  wire f_s_dadda_pg_rca32_fa778_y4;
  wire f_s_dadda_pg_rca32_and_30_27_a_30;
  wire f_s_dadda_pg_rca32_and_30_27_b_27;
  wire f_s_dadda_pg_rca32_and_30_27_y0;
  wire f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_fa778_y4;
  wire f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_fa777_y4;
  wire f_s_dadda_pg_rca32_fa779_y0;
  wire f_s_dadda_pg_rca32_fa779_y1;
  wire f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_and_30_27_y0;
  wire f_s_dadda_pg_rca32_fa779_y2;
  wire f_s_dadda_pg_rca32_fa779_y3;
  wire f_s_dadda_pg_rca32_fa779_y4;
  wire f_s_dadda_pg_rca32_and_29_28_a_29;
  wire f_s_dadda_pg_rca32_and_29_28_b_28;
  wire f_s_dadda_pg_rca32_and_29_28_y0;
  wire f_s_dadda_pg_rca32_and_28_29_a_28;
  wire f_s_dadda_pg_rca32_and_28_29_b_29;
  wire f_s_dadda_pg_rca32_and_28_29_y0;
  wire f_s_dadda_pg_rca32_and_27_30_a_27;
  wire f_s_dadda_pg_rca32_and_27_30_b_30;
  wire f_s_dadda_pg_rca32_and_27_30_y0;
  wire f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_29_28_y0;
  wire f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_28_29_y0;
  wire f_s_dadda_pg_rca32_fa780_y0;
  wire f_s_dadda_pg_rca32_fa780_y1;
  wire f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_27_30_y0;
  wire f_s_dadda_pg_rca32_fa780_y2;
  wire f_s_dadda_pg_rca32_fa780_y3;
  wire f_s_dadda_pg_rca32_fa780_y4;
  wire f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa780_y4;
  wire f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa779_y4;
  wire f_s_dadda_pg_rca32_fa781_y0;
  wire f_s_dadda_pg_rca32_fa781_y1;
  wire f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa675_y4;
  wire f_s_dadda_pg_rca32_fa781_y2;
  wire f_s_dadda_pg_rca32_fa781_y3;
  wire f_s_dadda_pg_rca32_fa781_y4;
  wire f_s_dadda_pg_rca32_nand_31_27_a_31;
  wire f_s_dadda_pg_rca32_nand_31_27_b_27;
  wire f_s_dadda_pg_rca32_nand_31_27_y0;
  wire f_s_dadda_pg_rca32_and_30_28_a_30;
  wire f_s_dadda_pg_rca32_and_30_28_b_28;
  wire f_s_dadda_pg_rca32_and_30_28_y0;
  wire f_s_dadda_pg_rca32_and_29_29_a_29;
  wire f_s_dadda_pg_rca32_and_29_29_b_29;
  wire f_s_dadda_pg_rca32_and_29_29_y0;
  wire f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_nand_31_27_y0;
  wire f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_and_30_28_y0;
  wire f_s_dadda_pg_rca32_fa782_y0;
  wire f_s_dadda_pg_rca32_fa782_y1;
  wire f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_and_29_29_y0;
  wire f_s_dadda_pg_rca32_fa782_y2;
  wire f_s_dadda_pg_rca32_fa782_y3;
  wire f_s_dadda_pg_rca32_fa782_y4;
  wire f_s_dadda_pg_rca32_nand_31_28_a_31;
  wire f_s_dadda_pg_rca32_nand_31_28_b_28;
  wire f_s_dadda_pg_rca32_nand_31_28_y0;
  wire f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_fa782_y4;
  wire f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_fa781_y4;
  wire f_s_dadda_pg_rca32_fa783_y0;
  wire f_s_dadda_pg_rca32_fa783_y1;
  wire f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_nand_31_28_y0;
  wire f_s_dadda_pg_rca32_fa783_y2;
  wire f_s_dadda_pg_rca32_fa783_y3;
  wire f_s_dadda_pg_rca32_fa783_y4;
  wire f_s_dadda_pg_rca32_and_3_0_a_3;
  wire f_s_dadda_pg_rca32_and_3_0_b_0;
  wire f_s_dadda_pg_rca32_and_3_0_y0;
  wire f_s_dadda_pg_rca32_and_2_1_a_2;
  wire f_s_dadda_pg_rca32_and_2_1_b_1;
  wire f_s_dadda_pg_rca32_and_2_1_y0;
  wire f_s_dadda_pg_rca32_ha28_f_s_dadda_pg_rca32_and_3_0_y0;
  wire f_s_dadda_pg_rca32_ha28_f_s_dadda_pg_rca32_and_2_1_y0;
  wire f_s_dadda_pg_rca32_ha28_y0;
  wire f_s_dadda_pg_rca32_ha28_y1;
  wire f_s_dadda_pg_rca32_and_2_2_a_2;
  wire f_s_dadda_pg_rca32_and_2_2_b_2;
  wire f_s_dadda_pg_rca32_and_2_2_y0;
  wire f_s_dadda_pg_rca32_and_1_3_a_1;
  wire f_s_dadda_pg_rca32_and_1_3_b_3;
  wire f_s_dadda_pg_rca32_and_1_3_y0;
  wire f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_ha28_y1;
  wire f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_and_2_2_y0;
  wire f_s_dadda_pg_rca32_fa784_y0;
  wire f_s_dadda_pg_rca32_fa784_y1;
  wire f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_and_1_3_y0;
  wire f_s_dadda_pg_rca32_fa784_y2;
  wire f_s_dadda_pg_rca32_fa784_y3;
  wire f_s_dadda_pg_rca32_fa784_y4;
  wire f_s_dadda_pg_rca32_and_1_4_a_1;
  wire f_s_dadda_pg_rca32_and_1_4_b_4;
  wire f_s_dadda_pg_rca32_and_1_4_y0;
  wire f_s_dadda_pg_rca32_and_0_5_a_0;
  wire f_s_dadda_pg_rca32_and_0_5_b_5;
  wire f_s_dadda_pg_rca32_and_0_5_y0;
  wire f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_fa784_y4;
  wire f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_and_1_4_y0;
  wire f_s_dadda_pg_rca32_fa785_y0;
  wire f_s_dadda_pg_rca32_fa785_y1;
  wire f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_and_0_5_y0;
  wire f_s_dadda_pg_rca32_fa785_y2;
  wire f_s_dadda_pg_rca32_fa785_y3;
  wire f_s_dadda_pg_rca32_fa785_y4;
  wire f_s_dadda_pg_rca32_and_0_6_a_0;
  wire f_s_dadda_pg_rca32_and_0_6_b_6;
  wire f_s_dadda_pg_rca32_and_0_6_y0;
  wire f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_fa785_y4;
  wire f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_and_0_6_y0;
  wire f_s_dadda_pg_rca32_fa786_y0;
  wire f_s_dadda_pg_rca32_fa786_y1;
  wire f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_ha4_y0;
  wire f_s_dadda_pg_rca32_fa786_y2;
  wire f_s_dadda_pg_rca32_fa786_y3;
  wire f_s_dadda_pg_rca32_fa786_y4;
  wire f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_fa786_y4;
  wire f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_fa16_y2;
  wire f_s_dadda_pg_rca32_fa787_y0;
  wire f_s_dadda_pg_rca32_fa787_y1;
  wire f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_ha5_y0;
  wire f_s_dadda_pg_rca32_fa787_y2;
  wire f_s_dadda_pg_rca32_fa787_y3;
  wire f_s_dadda_pg_rca32_fa787_y4;
  wire f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_fa787_y4;
  wire f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_fa18_y2;
  wire f_s_dadda_pg_rca32_fa788_y0;
  wire f_s_dadda_pg_rca32_fa788_y1;
  wire f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_ha6_y0;
  wire f_s_dadda_pg_rca32_fa788_y2;
  wire f_s_dadda_pg_rca32_fa788_y3;
  wire f_s_dadda_pg_rca32_fa788_y4;
  wire f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_fa788_y4;
  wire f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_fa21_y2;
  wire f_s_dadda_pg_rca32_fa789_y0;
  wire f_s_dadda_pg_rca32_fa789_y1;
  wire f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_ha7_y0;
  wire f_s_dadda_pg_rca32_fa789_y2;
  wire f_s_dadda_pg_rca32_fa789_y3;
  wire f_s_dadda_pg_rca32_fa789_y4;
  wire f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_fa789_y4;
  wire f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_fa25_y2;
  wire f_s_dadda_pg_rca32_fa790_y0;
  wire f_s_dadda_pg_rca32_fa790_y1;
  wire f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_ha8_y0;
  wire f_s_dadda_pg_rca32_fa790_y2;
  wire f_s_dadda_pg_rca32_fa790_y3;
  wire f_s_dadda_pg_rca32_fa790_y4;
  wire f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_fa790_y4;
  wire f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_fa30_y2;
  wire f_s_dadda_pg_rca32_fa791_y0;
  wire f_s_dadda_pg_rca32_fa791_y1;
  wire f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_ha9_y0;
  wire f_s_dadda_pg_rca32_fa791_y2;
  wire f_s_dadda_pg_rca32_fa791_y3;
  wire f_s_dadda_pg_rca32_fa791_y4;
  wire f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_fa791_y4;
  wire f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_fa36_y2;
  wire f_s_dadda_pg_rca32_fa792_y0;
  wire f_s_dadda_pg_rca32_fa792_y1;
  wire f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_ha10_y0;
  wire f_s_dadda_pg_rca32_fa792_y2;
  wire f_s_dadda_pg_rca32_fa792_y3;
  wire f_s_dadda_pg_rca32_fa792_y4;
  wire f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_fa792_y4;
  wire f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_fa43_y2;
  wire f_s_dadda_pg_rca32_fa793_y0;
  wire f_s_dadda_pg_rca32_fa793_y1;
  wire f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_ha11_y0;
  wire f_s_dadda_pg_rca32_fa793_y2;
  wire f_s_dadda_pg_rca32_fa793_y3;
  wire f_s_dadda_pg_rca32_fa793_y4;
  wire f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_fa793_y4;
  wire f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_fa51_y2;
  wire f_s_dadda_pg_rca32_fa794_y0;
  wire f_s_dadda_pg_rca32_fa794_y1;
  wire f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_ha12_y0;
  wire f_s_dadda_pg_rca32_fa794_y2;
  wire f_s_dadda_pg_rca32_fa794_y3;
  wire f_s_dadda_pg_rca32_fa794_y4;
  wire f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_fa794_y4;
  wire f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_fa60_y2;
  wire f_s_dadda_pg_rca32_fa795_y0;
  wire f_s_dadda_pg_rca32_fa795_y1;
  wire f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_ha13_y0;
  wire f_s_dadda_pg_rca32_fa795_y2;
  wire f_s_dadda_pg_rca32_fa795_y3;
  wire f_s_dadda_pg_rca32_fa795_y4;
  wire f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_fa795_y4;
  wire f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_fa70_y2;
  wire f_s_dadda_pg_rca32_fa796_y0;
  wire f_s_dadda_pg_rca32_fa796_y1;
  wire f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_ha14_y0;
  wire f_s_dadda_pg_rca32_fa796_y2;
  wire f_s_dadda_pg_rca32_fa796_y3;
  wire f_s_dadda_pg_rca32_fa796_y4;
  wire f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_fa796_y4;
  wire f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_fa81_y2;
  wire f_s_dadda_pg_rca32_fa797_y0;
  wire f_s_dadda_pg_rca32_fa797_y1;
  wire f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_ha15_y0;
  wire f_s_dadda_pg_rca32_fa797_y2;
  wire f_s_dadda_pg_rca32_fa797_y3;
  wire f_s_dadda_pg_rca32_fa797_y4;
  wire f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_fa797_y4;
  wire f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_fa93_y2;
  wire f_s_dadda_pg_rca32_fa798_y0;
  wire f_s_dadda_pg_rca32_fa798_y1;
  wire f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_ha16_y0;
  wire f_s_dadda_pg_rca32_fa798_y2;
  wire f_s_dadda_pg_rca32_fa798_y3;
  wire f_s_dadda_pg_rca32_fa798_y4;
  wire f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_fa798_y4;
  wire f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_fa106_y2;
  wire f_s_dadda_pg_rca32_fa799_y0;
  wire f_s_dadda_pg_rca32_fa799_y1;
  wire f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_ha17_y0;
  wire f_s_dadda_pg_rca32_fa799_y2;
  wire f_s_dadda_pg_rca32_fa799_y3;
  wire f_s_dadda_pg_rca32_fa799_y4;
  wire f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_fa799_y4;
  wire f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_fa120_y2;
  wire f_s_dadda_pg_rca32_fa800_y0;
  wire f_s_dadda_pg_rca32_fa800_y1;
  wire f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_ha18_y0;
  wire f_s_dadda_pg_rca32_fa800_y2;
  wire f_s_dadda_pg_rca32_fa800_y3;
  wire f_s_dadda_pg_rca32_fa800_y4;
  wire f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_fa800_y4;
  wire f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_fa135_y2;
  wire f_s_dadda_pg_rca32_fa801_y0;
  wire f_s_dadda_pg_rca32_fa801_y1;
  wire f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_ha19_y0;
  wire f_s_dadda_pg_rca32_fa801_y2;
  wire f_s_dadda_pg_rca32_fa801_y3;
  wire f_s_dadda_pg_rca32_fa801_y4;
  wire f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_fa801_y4;
  wire f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_fa151_y2;
  wire f_s_dadda_pg_rca32_fa802_y0;
  wire f_s_dadda_pg_rca32_fa802_y1;
  wire f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_ha20_y0;
  wire f_s_dadda_pg_rca32_fa802_y2;
  wire f_s_dadda_pg_rca32_fa802_y3;
  wire f_s_dadda_pg_rca32_fa802_y4;
  wire f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_fa802_y4;
  wire f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_fa168_y2;
  wire f_s_dadda_pg_rca32_fa803_y0;
  wire f_s_dadda_pg_rca32_fa803_y1;
  wire f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_ha21_y0;
  wire f_s_dadda_pg_rca32_fa803_y2;
  wire f_s_dadda_pg_rca32_fa803_y3;
  wire f_s_dadda_pg_rca32_fa803_y4;
  wire f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_fa803_y4;
  wire f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_fa186_y2;
  wire f_s_dadda_pg_rca32_fa804_y0;
  wire f_s_dadda_pg_rca32_fa804_y1;
  wire f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_ha22_y0;
  wire f_s_dadda_pg_rca32_fa804_y2;
  wire f_s_dadda_pg_rca32_fa804_y3;
  wire f_s_dadda_pg_rca32_fa804_y4;
  wire f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_fa804_y4;
  wire f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_fa205_y2;
  wire f_s_dadda_pg_rca32_fa805_y0;
  wire f_s_dadda_pg_rca32_fa805_y1;
  wire f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_ha23_y0;
  wire f_s_dadda_pg_rca32_fa805_y2;
  wire f_s_dadda_pg_rca32_fa805_y3;
  wire f_s_dadda_pg_rca32_fa805_y4;
  wire f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_fa805_y4;
  wire f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_fa225_y2;
  wire f_s_dadda_pg_rca32_fa806_y0;
  wire f_s_dadda_pg_rca32_fa806_y1;
  wire f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_ha24_y0;
  wire f_s_dadda_pg_rca32_fa806_y2;
  wire f_s_dadda_pg_rca32_fa806_y3;
  wire f_s_dadda_pg_rca32_fa806_y4;
  wire f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_fa806_y4;
  wire f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_fa246_y2;
  wire f_s_dadda_pg_rca32_fa807_y0;
  wire f_s_dadda_pg_rca32_fa807_y1;
  wire f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_ha25_y0;
  wire f_s_dadda_pg_rca32_fa807_y2;
  wire f_s_dadda_pg_rca32_fa807_y3;
  wire f_s_dadda_pg_rca32_fa807_y4;
  wire f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa807_y4;
  wire f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa267_y2;
  wire f_s_dadda_pg_rca32_fa808_y0;
  wire f_s_dadda_pg_rca32_fa808_y1;
  wire f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa268_y2;
  wire f_s_dadda_pg_rca32_fa808_y2;
  wire f_s_dadda_pg_rca32_fa808_y3;
  wire f_s_dadda_pg_rca32_fa808_y4;
  wire f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa808_y4;
  wire f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa289_y2;
  wire f_s_dadda_pg_rca32_fa809_y0;
  wire f_s_dadda_pg_rca32_fa809_y1;
  wire f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa290_y2;
  wire f_s_dadda_pg_rca32_fa809_y2;
  wire f_s_dadda_pg_rca32_fa809_y3;
  wire f_s_dadda_pg_rca32_fa809_y4;
  wire f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa809_y4;
  wire f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa311_y2;
  wire f_s_dadda_pg_rca32_fa810_y0;
  wire f_s_dadda_pg_rca32_fa810_y1;
  wire f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa312_y2;
  wire f_s_dadda_pg_rca32_fa810_y2;
  wire f_s_dadda_pg_rca32_fa810_y3;
  wire f_s_dadda_pg_rca32_fa810_y4;
  wire f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa810_y4;
  wire f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa333_y2;
  wire f_s_dadda_pg_rca32_fa811_y0;
  wire f_s_dadda_pg_rca32_fa811_y1;
  wire f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa334_y2;
  wire f_s_dadda_pg_rca32_fa811_y2;
  wire f_s_dadda_pg_rca32_fa811_y3;
  wire f_s_dadda_pg_rca32_fa811_y4;
  wire f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa811_y4;
  wire f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa355_y2;
  wire f_s_dadda_pg_rca32_fa812_y0;
  wire f_s_dadda_pg_rca32_fa812_y1;
  wire f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa356_y2;
  wire f_s_dadda_pg_rca32_fa812_y2;
  wire f_s_dadda_pg_rca32_fa812_y3;
  wire f_s_dadda_pg_rca32_fa812_y4;
  wire f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa812_y4;
  wire f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa377_y2;
  wire f_s_dadda_pg_rca32_fa813_y0;
  wire f_s_dadda_pg_rca32_fa813_y1;
  wire f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa378_y2;
  wire f_s_dadda_pg_rca32_fa813_y2;
  wire f_s_dadda_pg_rca32_fa813_y3;
  wire f_s_dadda_pg_rca32_fa813_y4;
  wire f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa813_y4;
  wire f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa399_y2;
  wire f_s_dadda_pg_rca32_fa814_y0;
  wire f_s_dadda_pg_rca32_fa814_y1;
  wire f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa400_y2;
  wire f_s_dadda_pg_rca32_fa814_y2;
  wire f_s_dadda_pg_rca32_fa814_y3;
  wire f_s_dadda_pg_rca32_fa814_y4;
  wire f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa814_y4;
  wire f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa421_y2;
  wire f_s_dadda_pg_rca32_fa815_y0;
  wire f_s_dadda_pg_rca32_fa815_y1;
  wire f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa422_y2;
  wire f_s_dadda_pg_rca32_fa815_y2;
  wire f_s_dadda_pg_rca32_fa815_y3;
  wire f_s_dadda_pg_rca32_fa815_y4;
  wire f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa815_y4;
  wire f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa443_y2;
  wire f_s_dadda_pg_rca32_fa816_y0;
  wire f_s_dadda_pg_rca32_fa816_y1;
  wire f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa444_y2;
  wire f_s_dadda_pg_rca32_fa816_y2;
  wire f_s_dadda_pg_rca32_fa816_y3;
  wire f_s_dadda_pg_rca32_fa816_y4;
  wire f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa816_y4;
  wire f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa464_y2;
  wire f_s_dadda_pg_rca32_fa817_y0;
  wire f_s_dadda_pg_rca32_fa817_y1;
  wire f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa465_y2;
  wire f_s_dadda_pg_rca32_fa817_y2;
  wire f_s_dadda_pg_rca32_fa817_y3;
  wire f_s_dadda_pg_rca32_fa817_y4;
  wire f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa817_y4;
  wire f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa484_y2;
  wire f_s_dadda_pg_rca32_fa818_y0;
  wire f_s_dadda_pg_rca32_fa818_y1;
  wire f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa485_y2;
  wire f_s_dadda_pg_rca32_fa818_y2;
  wire f_s_dadda_pg_rca32_fa818_y3;
  wire f_s_dadda_pg_rca32_fa818_y4;
  wire f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa818_y4;
  wire f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa503_y2;
  wire f_s_dadda_pg_rca32_fa819_y0;
  wire f_s_dadda_pg_rca32_fa819_y1;
  wire f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa504_y2;
  wire f_s_dadda_pg_rca32_fa819_y2;
  wire f_s_dadda_pg_rca32_fa819_y3;
  wire f_s_dadda_pg_rca32_fa819_y4;
  wire f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa819_y4;
  wire f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa521_y2;
  wire f_s_dadda_pg_rca32_fa820_y0;
  wire f_s_dadda_pg_rca32_fa820_y1;
  wire f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa522_y2;
  wire f_s_dadda_pg_rca32_fa820_y2;
  wire f_s_dadda_pg_rca32_fa820_y3;
  wire f_s_dadda_pg_rca32_fa820_y4;
  wire f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa820_y4;
  wire f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa538_y2;
  wire f_s_dadda_pg_rca32_fa821_y0;
  wire f_s_dadda_pg_rca32_fa821_y1;
  wire f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa539_y2;
  wire f_s_dadda_pg_rca32_fa821_y2;
  wire f_s_dadda_pg_rca32_fa821_y3;
  wire f_s_dadda_pg_rca32_fa821_y4;
  wire f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa821_y4;
  wire f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa554_y2;
  wire f_s_dadda_pg_rca32_fa822_y0;
  wire f_s_dadda_pg_rca32_fa822_y1;
  wire f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa555_y2;
  wire f_s_dadda_pg_rca32_fa822_y2;
  wire f_s_dadda_pg_rca32_fa822_y3;
  wire f_s_dadda_pg_rca32_fa822_y4;
  wire f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa822_y4;
  wire f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa569_y2;
  wire f_s_dadda_pg_rca32_fa823_y0;
  wire f_s_dadda_pg_rca32_fa823_y1;
  wire f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa570_y2;
  wire f_s_dadda_pg_rca32_fa823_y2;
  wire f_s_dadda_pg_rca32_fa823_y3;
  wire f_s_dadda_pg_rca32_fa823_y4;
  wire f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa823_y4;
  wire f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa583_y2;
  wire f_s_dadda_pg_rca32_fa824_y0;
  wire f_s_dadda_pg_rca32_fa824_y1;
  wire f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa584_y2;
  wire f_s_dadda_pg_rca32_fa824_y2;
  wire f_s_dadda_pg_rca32_fa824_y3;
  wire f_s_dadda_pg_rca32_fa824_y4;
  wire f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa824_y4;
  wire f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa596_y2;
  wire f_s_dadda_pg_rca32_fa825_y0;
  wire f_s_dadda_pg_rca32_fa825_y1;
  wire f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa597_y2;
  wire f_s_dadda_pg_rca32_fa825_y2;
  wire f_s_dadda_pg_rca32_fa825_y3;
  wire f_s_dadda_pg_rca32_fa825_y4;
  wire f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa825_y4;
  wire f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa608_y2;
  wire f_s_dadda_pg_rca32_fa826_y0;
  wire f_s_dadda_pg_rca32_fa826_y1;
  wire f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa609_y2;
  wire f_s_dadda_pg_rca32_fa826_y2;
  wire f_s_dadda_pg_rca32_fa826_y3;
  wire f_s_dadda_pg_rca32_fa826_y4;
  wire f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa826_y4;
  wire f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa619_y2;
  wire f_s_dadda_pg_rca32_fa827_y0;
  wire f_s_dadda_pg_rca32_fa827_y1;
  wire f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa620_y2;
  wire f_s_dadda_pg_rca32_fa827_y2;
  wire f_s_dadda_pg_rca32_fa827_y3;
  wire f_s_dadda_pg_rca32_fa827_y4;
  wire f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa827_y4;
  wire f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa629_y2;
  wire f_s_dadda_pg_rca32_fa828_y0;
  wire f_s_dadda_pg_rca32_fa828_y1;
  wire f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa630_y2;
  wire f_s_dadda_pg_rca32_fa828_y2;
  wire f_s_dadda_pg_rca32_fa828_y3;
  wire f_s_dadda_pg_rca32_fa828_y4;
  wire f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa828_y4;
  wire f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa638_y2;
  wire f_s_dadda_pg_rca32_fa829_y0;
  wire f_s_dadda_pg_rca32_fa829_y1;
  wire f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa639_y2;
  wire f_s_dadda_pg_rca32_fa829_y2;
  wire f_s_dadda_pg_rca32_fa829_y3;
  wire f_s_dadda_pg_rca32_fa829_y4;
  wire f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa829_y4;
  wire f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa646_y2;
  wire f_s_dadda_pg_rca32_fa830_y0;
  wire f_s_dadda_pg_rca32_fa830_y1;
  wire f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa647_y2;
  wire f_s_dadda_pg_rca32_fa830_y2;
  wire f_s_dadda_pg_rca32_fa830_y3;
  wire f_s_dadda_pg_rca32_fa830_y4;
  wire f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa830_y4;
  wire f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa653_y2;
  wire f_s_dadda_pg_rca32_fa831_y0;
  wire f_s_dadda_pg_rca32_fa831_y1;
  wire f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa654_y2;
  wire f_s_dadda_pg_rca32_fa831_y2;
  wire f_s_dadda_pg_rca32_fa831_y3;
  wire f_s_dadda_pg_rca32_fa831_y4;
  wire f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa831_y4;
  wire f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa659_y2;
  wire f_s_dadda_pg_rca32_fa832_y0;
  wire f_s_dadda_pg_rca32_fa832_y1;
  wire f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa660_y2;
  wire f_s_dadda_pg_rca32_fa832_y2;
  wire f_s_dadda_pg_rca32_fa832_y3;
  wire f_s_dadda_pg_rca32_fa832_y4;
  wire f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa832_y4;
  wire f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa664_y2;
  wire f_s_dadda_pg_rca32_fa833_y0;
  wire f_s_dadda_pg_rca32_fa833_y1;
  wire f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa665_y2;
  wire f_s_dadda_pg_rca32_fa833_y2;
  wire f_s_dadda_pg_rca32_fa833_y3;
  wire f_s_dadda_pg_rca32_fa833_y4;
  wire f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa833_y4;
  wire f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa668_y2;
  wire f_s_dadda_pg_rca32_fa834_y0;
  wire f_s_dadda_pg_rca32_fa834_y1;
  wire f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa669_y2;
  wire f_s_dadda_pg_rca32_fa834_y2;
  wire f_s_dadda_pg_rca32_fa834_y3;
  wire f_s_dadda_pg_rca32_fa834_y4;
  wire f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa834_y4;
  wire f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa671_y2;
  wire f_s_dadda_pg_rca32_fa835_y0;
  wire f_s_dadda_pg_rca32_fa835_y1;
  wire f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa672_y2;
  wire f_s_dadda_pg_rca32_fa835_y2;
  wire f_s_dadda_pg_rca32_fa835_y3;
  wire f_s_dadda_pg_rca32_fa835_y4;
  wire f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa835_y4;
  wire f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa673_y2;
  wire f_s_dadda_pg_rca32_fa836_y0;
  wire f_s_dadda_pg_rca32_fa836_y1;
  wire f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa674_y2;
  wire f_s_dadda_pg_rca32_fa836_y2;
  wire f_s_dadda_pg_rca32_fa836_y3;
  wire f_s_dadda_pg_rca32_fa836_y4;
  wire f_s_dadda_pg_rca32_nand_26_31_a_26;
  wire f_s_dadda_pg_rca32_nand_26_31_b_31;
  wire f_s_dadda_pg_rca32_nand_26_31_y0;
  wire f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_fa836_y4;
  wire f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_nand_26_31_y0;
  wire f_s_dadda_pg_rca32_fa837_y0;
  wire f_s_dadda_pg_rca32_fa837_y1;
  wire f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_fa675_y2;
  wire f_s_dadda_pg_rca32_fa837_y2;
  wire f_s_dadda_pg_rca32_fa837_y3;
  wire f_s_dadda_pg_rca32_fa837_y4;
  wire f_s_dadda_pg_rca32_and_28_30_a_28;
  wire f_s_dadda_pg_rca32_and_28_30_b_30;
  wire f_s_dadda_pg_rca32_and_28_30_y0;
  wire f_s_dadda_pg_rca32_nand_27_31_a_27;
  wire f_s_dadda_pg_rca32_nand_27_31_b_31;
  wire f_s_dadda_pg_rca32_nand_27_31_y0;
  wire f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_fa837_y4;
  wire f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_and_28_30_y0;
  wire f_s_dadda_pg_rca32_fa838_y0;
  wire f_s_dadda_pg_rca32_fa838_y1;
  wire f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_nand_27_31_y0;
  wire f_s_dadda_pg_rca32_fa838_y2;
  wire f_s_dadda_pg_rca32_fa838_y3;
  wire f_s_dadda_pg_rca32_fa838_y4;
  wire f_s_dadda_pg_rca32_and_30_29_a_30;
  wire f_s_dadda_pg_rca32_and_30_29_b_29;
  wire f_s_dadda_pg_rca32_and_30_29_y0;
  wire f_s_dadda_pg_rca32_and_29_30_a_29;
  wire f_s_dadda_pg_rca32_and_29_30_b_30;
  wire f_s_dadda_pg_rca32_and_29_30_y0;
  wire f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_fa838_y4;
  wire f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_and_30_29_y0;
  wire f_s_dadda_pg_rca32_fa839_y0;
  wire f_s_dadda_pg_rca32_fa839_y1;
  wire f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_and_29_30_y0;
  wire f_s_dadda_pg_rca32_fa839_y2;
  wire f_s_dadda_pg_rca32_fa839_y3;
  wire f_s_dadda_pg_rca32_fa839_y4;
  wire f_s_dadda_pg_rca32_nand_31_29_a_31;
  wire f_s_dadda_pg_rca32_nand_31_29_b_29;
  wire f_s_dadda_pg_rca32_nand_31_29_y0;
  wire f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_fa839_y4;
  wire f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_fa783_y4;
  wire f_s_dadda_pg_rca32_fa840_y0;
  wire f_s_dadda_pg_rca32_fa840_y1;
  wire f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_nand_31_29_y0;
  wire f_s_dadda_pg_rca32_fa840_y2;
  wire f_s_dadda_pg_rca32_fa840_y3;
  wire f_s_dadda_pg_rca32_fa840_y4;
  wire f_s_dadda_pg_rca32_and_2_0_a_2;
  wire f_s_dadda_pg_rca32_and_2_0_b_0;
  wire f_s_dadda_pg_rca32_and_2_0_y0;
  wire f_s_dadda_pg_rca32_and_1_1_a_1;
  wire f_s_dadda_pg_rca32_and_1_1_b_1;
  wire f_s_dadda_pg_rca32_and_1_1_y0;
  wire f_s_dadda_pg_rca32_ha29_f_s_dadda_pg_rca32_and_2_0_y0;
  wire f_s_dadda_pg_rca32_ha29_f_s_dadda_pg_rca32_and_1_1_y0;
  wire f_s_dadda_pg_rca32_ha29_y0;
  wire f_s_dadda_pg_rca32_ha29_y1;
  wire f_s_dadda_pg_rca32_and_1_2_a_1;
  wire f_s_dadda_pg_rca32_and_1_2_b_2;
  wire f_s_dadda_pg_rca32_and_1_2_y0;
  wire f_s_dadda_pg_rca32_and_0_3_a_0;
  wire f_s_dadda_pg_rca32_and_0_3_b_3;
  wire f_s_dadda_pg_rca32_and_0_3_y0;
  wire f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_ha29_y1;
  wire f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_and_1_2_y0;
  wire f_s_dadda_pg_rca32_fa841_y0;
  wire f_s_dadda_pg_rca32_fa841_y1;
  wire f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_and_0_3_y0;
  wire f_s_dadda_pg_rca32_fa841_y2;
  wire f_s_dadda_pg_rca32_fa841_y3;
  wire f_s_dadda_pg_rca32_fa841_y4;
  wire f_s_dadda_pg_rca32_and_0_4_a_0;
  wire f_s_dadda_pg_rca32_and_0_4_b_4;
  wire f_s_dadda_pg_rca32_and_0_4_y0;
  wire f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_fa841_y4;
  wire f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_and_0_4_y0;
  wire f_s_dadda_pg_rca32_fa842_y0;
  wire f_s_dadda_pg_rca32_fa842_y1;
  wire f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_ha26_y0;
  wire f_s_dadda_pg_rca32_fa842_y2;
  wire f_s_dadda_pg_rca32_fa842_y3;
  wire f_s_dadda_pg_rca32_fa842_y4;
  wire f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_fa842_y4;
  wire f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_fa676_y2;
  wire f_s_dadda_pg_rca32_fa843_y0;
  wire f_s_dadda_pg_rca32_fa843_y1;
  wire f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_ha27_y0;
  wire f_s_dadda_pg_rca32_fa843_y2;
  wire f_s_dadda_pg_rca32_fa843_y3;
  wire f_s_dadda_pg_rca32_fa843_y4;
  wire f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa843_y4;
  wire f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa677_y2;
  wire f_s_dadda_pg_rca32_fa844_y0;
  wire f_s_dadda_pg_rca32_fa844_y1;
  wire f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa678_y2;
  wire f_s_dadda_pg_rca32_fa844_y2;
  wire f_s_dadda_pg_rca32_fa844_y3;
  wire f_s_dadda_pg_rca32_fa844_y4;
  wire f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa844_y4;
  wire f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa679_y2;
  wire f_s_dadda_pg_rca32_fa845_y0;
  wire f_s_dadda_pg_rca32_fa845_y1;
  wire f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa680_y2;
  wire f_s_dadda_pg_rca32_fa845_y2;
  wire f_s_dadda_pg_rca32_fa845_y3;
  wire f_s_dadda_pg_rca32_fa845_y4;
  wire f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa845_y4;
  wire f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa681_y2;
  wire f_s_dadda_pg_rca32_fa846_y0;
  wire f_s_dadda_pg_rca32_fa846_y1;
  wire f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa682_y2;
  wire f_s_dadda_pg_rca32_fa846_y2;
  wire f_s_dadda_pg_rca32_fa846_y3;
  wire f_s_dadda_pg_rca32_fa846_y4;
  wire f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa846_y4;
  wire f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa683_y2;
  wire f_s_dadda_pg_rca32_fa847_y0;
  wire f_s_dadda_pg_rca32_fa847_y1;
  wire f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa684_y2;
  wire f_s_dadda_pg_rca32_fa847_y2;
  wire f_s_dadda_pg_rca32_fa847_y3;
  wire f_s_dadda_pg_rca32_fa847_y4;
  wire f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa847_y4;
  wire f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa685_y2;
  wire f_s_dadda_pg_rca32_fa848_y0;
  wire f_s_dadda_pg_rca32_fa848_y1;
  wire f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa686_y2;
  wire f_s_dadda_pg_rca32_fa848_y2;
  wire f_s_dadda_pg_rca32_fa848_y3;
  wire f_s_dadda_pg_rca32_fa848_y4;
  wire f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa848_y4;
  wire f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa687_y2;
  wire f_s_dadda_pg_rca32_fa849_y0;
  wire f_s_dadda_pg_rca32_fa849_y1;
  wire f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa688_y2;
  wire f_s_dadda_pg_rca32_fa849_y2;
  wire f_s_dadda_pg_rca32_fa849_y3;
  wire f_s_dadda_pg_rca32_fa849_y4;
  wire f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa849_y4;
  wire f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa689_y2;
  wire f_s_dadda_pg_rca32_fa850_y0;
  wire f_s_dadda_pg_rca32_fa850_y1;
  wire f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa690_y2;
  wire f_s_dadda_pg_rca32_fa850_y2;
  wire f_s_dadda_pg_rca32_fa850_y3;
  wire f_s_dadda_pg_rca32_fa850_y4;
  wire f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa850_y4;
  wire f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa691_y2;
  wire f_s_dadda_pg_rca32_fa851_y0;
  wire f_s_dadda_pg_rca32_fa851_y1;
  wire f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa692_y2;
  wire f_s_dadda_pg_rca32_fa851_y2;
  wire f_s_dadda_pg_rca32_fa851_y3;
  wire f_s_dadda_pg_rca32_fa851_y4;
  wire f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa851_y4;
  wire f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa693_y2;
  wire f_s_dadda_pg_rca32_fa852_y0;
  wire f_s_dadda_pg_rca32_fa852_y1;
  wire f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa694_y2;
  wire f_s_dadda_pg_rca32_fa852_y2;
  wire f_s_dadda_pg_rca32_fa852_y3;
  wire f_s_dadda_pg_rca32_fa852_y4;
  wire f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa852_y4;
  wire f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa695_y2;
  wire f_s_dadda_pg_rca32_fa853_y0;
  wire f_s_dadda_pg_rca32_fa853_y1;
  wire f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa696_y2;
  wire f_s_dadda_pg_rca32_fa853_y2;
  wire f_s_dadda_pg_rca32_fa853_y3;
  wire f_s_dadda_pg_rca32_fa853_y4;
  wire f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa853_y4;
  wire f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa697_y2;
  wire f_s_dadda_pg_rca32_fa854_y0;
  wire f_s_dadda_pg_rca32_fa854_y1;
  wire f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa698_y2;
  wire f_s_dadda_pg_rca32_fa854_y2;
  wire f_s_dadda_pg_rca32_fa854_y3;
  wire f_s_dadda_pg_rca32_fa854_y4;
  wire f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa854_y4;
  wire f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa699_y2;
  wire f_s_dadda_pg_rca32_fa855_y0;
  wire f_s_dadda_pg_rca32_fa855_y1;
  wire f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa700_y2;
  wire f_s_dadda_pg_rca32_fa855_y2;
  wire f_s_dadda_pg_rca32_fa855_y3;
  wire f_s_dadda_pg_rca32_fa855_y4;
  wire f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa855_y4;
  wire f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa701_y2;
  wire f_s_dadda_pg_rca32_fa856_y0;
  wire f_s_dadda_pg_rca32_fa856_y1;
  wire f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa702_y2;
  wire f_s_dadda_pg_rca32_fa856_y2;
  wire f_s_dadda_pg_rca32_fa856_y3;
  wire f_s_dadda_pg_rca32_fa856_y4;
  wire f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa856_y4;
  wire f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa703_y2;
  wire f_s_dadda_pg_rca32_fa857_y0;
  wire f_s_dadda_pg_rca32_fa857_y1;
  wire f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa704_y2;
  wire f_s_dadda_pg_rca32_fa857_y2;
  wire f_s_dadda_pg_rca32_fa857_y3;
  wire f_s_dadda_pg_rca32_fa857_y4;
  wire f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa857_y4;
  wire f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa705_y2;
  wire f_s_dadda_pg_rca32_fa858_y0;
  wire f_s_dadda_pg_rca32_fa858_y1;
  wire f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa706_y2;
  wire f_s_dadda_pg_rca32_fa858_y2;
  wire f_s_dadda_pg_rca32_fa858_y3;
  wire f_s_dadda_pg_rca32_fa858_y4;
  wire f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa858_y4;
  wire f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa707_y2;
  wire f_s_dadda_pg_rca32_fa859_y0;
  wire f_s_dadda_pg_rca32_fa859_y1;
  wire f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa708_y2;
  wire f_s_dadda_pg_rca32_fa859_y2;
  wire f_s_dadda_pg_rca32_fa859_y3;
  wire f_s_dadda_pg_rca32_fa859_y4;
  wire f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa859_y4;
  wire f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa709_y2;
  wire f_s_dadda_pg_rca32_fa860_y0;
  wire f_s_dadda_pg_rca32_fa860_y1;
  wire f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa710_y2;
  wire f_s_dadda_pg_rca32_fa860_y2;
  wire f_s_dadda_pg_rca32_fa860_y3;
  wire f_s_dadda_pg_rca32_fa860_y4;
  wire f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa860_y4;
  wire f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa711_y2;
  wire f_s_dadda_pg_rca32_fa861_y0;
  wire f_s_dadda_pg_rca32_fa861_y1;
  wire f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa712_y2;
  wire f_s_dadda_pg_rca32_fa861_y2;
  wire f_s_dadda_pg_rca32_fa861_y3;
  wire f_s_dadda_pg_rca32_fa861_y4;
  wire f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa861_y4;
  wire f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa713_y2;
  wire f_s_dadda_pg_rca32_fa862_y0;
  wire f_s_dadda_pg_rca32_fa862_y1;
  wire f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa714_y2;
  wire f_s_dadda_pg_rca32_fa862_y2;
  wire f_s_dadda_pg_rca32_fa862_y3;
  wire f_s_dadda_pg_rca32_fa862_y4;
  wire f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa862_y4;
  wire f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa715_y2;
  wire f_s_dadda_pg_rca32_fa863_y0;
  wire f_s_dadda_pg_rca32_fa863_y1;
  wire f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa716_y2;
  wire f_s_dadda_pg_rca32_fa863_y2;
  wire f_s_dadda_pg_rca32_fa863_y3;
  wire f_s_dadda_pg_rca32_fa863_y4;
  wire f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa863_y4;
  wire f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa717_y2;
  wire f_s_dadda_pg_rca32_fa864_y0;
  wire f_s_dadda_pg_rca32_fa864_y1;
  wire f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa718_y2;
  wire f_s_dadda_pg_rca32_fa864_y2;
  wire f_s_dadda_pg_rca32_fa864_y3;
  wire f_s_dadda_pg_rca32_fa864_y4;
  wire f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa864_y4;
  wire f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa719_y2;
  wire f_s_dadda_pg_rca32_fa865_y0;
  wire f_s_dadda_pg_rca32_fa865_y1;
  wire f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa720_y2;
  wire f_s_dadda_pg_rca32_fa865_y2;
  wire f_s_dadda_pg_rca32_fa865_y3;
  wire f_s_dadda_pg_rca32_fa865_y4;
  wire f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa865_y4;
  wire f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa721_y2;
  wire f_s_dadda_pg_rca32_fa866_y0;
  wire f_s_dadda_pg_rca32_fa866_y1;
  wire f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa722_y2;
  wire f_s_dadda_pg_rca32_fa866_y2;
  wire f_s_dadda_pg_rca32_fa866_y3;
  wire f_s_dadda_pg_rca32_fa866_y4;
  wire f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa866_y4;
  wire f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa723_y2;
  wire f_s_dadda_pg_rca32_fa867_y0;
  wire f_s_dadda_pg_rca32_fa867_y1;
  wire f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa724_y2;
  wire f_s_dadda_pg_rca32_fa867_y2;
  wire f_s_dadda_pg_rca32_fa867_y3;
  wire f_s_dadda_pg_rca32_fa867_y4;
  wire f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa867_y4;
  wire f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa725_y2;
  wire f_s_dadda_pg_rca32_fa868_y0;
  wire f_s_dadda_pg_rca32_fa868_y1;
  wire f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa726_y2;
  wire f_s_dadda_pg_rca32_fa868_y2;
  wire f_s_dadda_pg_rca32_fa868_y3;
  wire f_s_dadda_pg_rca32_fa868_y4;
  wire f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa868_y4;
  wire f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa727_y2;
  wire f_s_dadda_pg_rca32_fa869_y0;
  wire f_s_dadda_pg_rca32_fa869_y1;
  wire f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa728_y2;
  wire f_s_dadda_pg_rca32_fa869_y2;
  wire f_s_dadda_pg_rca32_fa869_y3;
  wire f_s_dadda_pg_rca32_fa869_y4;
  wire f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa869_y4;
  wire f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa729_y2;
  wire f_s_dadda_pg_rca32_fa870_y0;
  wire f_s_dadda_pg_rca32_fa870_y1;
  wire f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa730_y2;
  wire f_s_dadda_pg_rca32_fa870_y2;
  wire f_s_dadda_pg_rca32_fa870_y3;
  wire f_s_dadda_pg_rca32_fa870_y4;
  wire f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa870_y4;
  wire f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa731_y2;
  wire f_s_dadda_pg_rca32_fa871_y0;
  wire f_s_dadda_pg_rca32_fa871_y1;
  wire f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa732_y2;
  wire f_s_dadda_pg_rca32_fa871_y2;
  wire f_s_dadda_pg_rca32_fa871_y3;
  wire f_s_dadda_pg_rca32_fa871_y4;
  wire f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa871_y4;
  wire f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa733_y2;
  wire f_s_dadda_pg_rca32_fa872_y0;
  wire f_s_dadda_pg_rca32_fa872_y1;
  wire f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa734_y2;
  wire f_s_dadda_pg_rca32_fa872_y2;
  wire f_s_dadda_pg_rca32_fa872_y3;
  wire f_s_dadda_pg_rca32_fa872_y4;
  wire f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa872_y4;
  wire f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa735_y2;
  wire f_s_dadda_pg_rca32_fa873_y0;
  wire f_s_dadda_pg_rca32_fa873_y1;
  wire f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa736_y2;
  wire f_s_dadda_pg_rca32_fa873_y2;
  wire f_s_dadda_pg_rca32_fa873_y3;
  wire f_s_dadda_pg_rca32_fa873_y4;
  wire f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa873_y4;
  wire f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa737_y2;
  wire f_s_dadda_pg_rca32_fa874_y0;
  wire f_s_dadda_pg_rca32_fa874_y1;
  wire f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa738_y2;
  wire f_s_dadda_pg_rca32_fa874_y2;
  wire f_s_dadda_pg_rca32_fa874_y3;
  wire f_s_dadda_pg_rca32_fa874_y4;
  wire f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa874_y4;
  wire f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa739_y2;
  wire f_s_dadda_pg_rca32_fa875_y0;
  wire f_s_dadda_pg_rca32_fa875_y1;
  wire f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa740_y2;
  wire f_s_dadda_pg_rca32_fa875_y2;
  wire f_s_dadda_pg_rca32_fa875_y3;
  wire f_s_dadda_pg_rca32_fa875_y4;
  wire f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa875_y4;
  wire f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa741_y2;
  wire f_s_dadda_pg_rca32_fa876_y0;
  wire f_s_dadda_pg_rca32_fa876_y1;
  wire f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa742_y2;
  wire f_s_dadda_pg_rca32_fa876_y2;
  wire f_s_dadda_pg_rca32_fa876_y3;
  wire f_s_dadda_pg_rca32_fa876_y4;
  wire f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa876_y4;
  wire f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa743_y2;
  wire f_s_dadda_pg_rca32_fa877_y0;
  wire f_s_dadda_pg_rca32_fa877_y1;
  wire f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa744_y2;
  wire f_s_dadda_pg_rca32_fa877_y2;
  wire f_s_dadda_pg_rca32_fa877_y3;
  wire f_s_dadda_pg_rca32_fa877_y4;
  wire f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa877_y4;
  wire f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa745_y2;
  wire f_s_dadda_pg_rca32_fa878_y0;
  wire f_s_dadda_pg_rca32_fa878_y1;
  wire f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa746_y2;
  wire f_s_dadda_pg_rca32_fa878_y2;
  wire f_s_dadda_pg_rca32_fa878_y3;
  wire f_s_dadda_pg_rca32_fa878_y4;
  wire f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa878_y4;
  wire f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa747_y2;
  wire f_s_dadda_pg_rca32_fa879_y0;
  wire f_s_dadda_pg_rca32_fa879_y1;
  wire f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa748_y2;
  wire f_s_dadda_pg_rca32_fa879_y2;
  wire f_s_dadda_pg_rca32_fa879_y3;
  wire f_s_dadda_pg_rca32_fa879_y4;
  wire f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa879_y4;
  wire f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa749_y2;
  wire f_s_dadda_pg_rca32_fa880_y0;
  wire f_s_dadda_pg_rca32_fa880_y1;
  wire f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa750_y2;
  wire f_s_dadda_pg_rca32_fa880_y2;
  wire f_s_dadda_pg_rca32_fa880_y3;
  wire f_s_dadda_pg_rca32_fa880_y4;
  wire f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa880_y4;
  wire f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa751_y2;
  wire f_s_dadda_pg_rca32_fa881_y0;
  wire f_s_dadda_pg_rca32_fa881_y1;
  wire f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa752_y2;
  wire f_s_dadda_pg_rca32_fa881_y2;
  wire f_s_dadda_pg_rca32_fa881_y3;
  wire f_s_dadda_pg_rca32_fa881_y4;
  wire f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa881_y4;
  wire f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa753_y2;
  wire f_s_dadda_pg_rca32_fa882_y0;
  wire f_s_dadda_pg_rca32_fa882_y1;
  wire f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa754_y2;
  wire f_s_dadda_pg_rca32_fa882_y2;
  wire f_s_dadda_pg_rca32_fa882_y3;
  wire f_s_dadda_pg_rca32_fa882_y4;
  wire f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa882_y4;
  wire f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa755_y2;
  wire f_s_dadda_pg_rca32_fa883_y0;
  wire f_s_dadda_pg_rca32_fa883_y1;
  wire f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa756_y2;
  wire f_s_dadda_pg_rca32_fa883_y2;
  wire f_s_dadda_pg_rca32_fa883_y3;
  wire f_s_dadda_pg_rca32_fa883_y4;
  wire f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa883_y4;
  wire f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa757_y2;
  wire f_s_dadda_pg_rca32_fa884_y0;
  wire f_s_dadda_pg_rca32_fa884_y1;
  wire f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa758_y2;
  wire f_s_dadda_pg_rca32_fa884_y2;
  wire f_s_dadda_pg_rca32_fa884_y3;
  wire f_s_dadda_pg_rca32_fa884_y4;
  wire f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa884_y4;
  wire f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa759_y2;
  wire f_s_dadda_pg_rca32_fa885_y0;
  wire f_s_dadda_pg_rca32_fa885_y1;
  wire f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa760_y2;
  wire f_s_dadda_pg_rca32_fa885_y2;
  wire f_s_dadda_pg_rca32_fa885_y3;
  wire f_s_dadda_pg_rca32_fa885_y4;
  wire f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa885_y4;
  wire f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa761_y2;
  wire f_s_dadda_pg_rca32_fa886_y0;
  wire f_s_dadda_pg_rca32_fa886_y1;
  wire f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa762_y2;
  wire f_s_dadda_pg_rca32_fa886_y2;
  wire f_s_dadda_pg_rca32_fa886_y3;
  wire f_s_dadda_pg_rca32_fa886_y4;
  wire f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa886_y4;
  wire f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa763_y2;
  wire f_s_dadda_pg_rca32_fa887_y0;
  wire f_s_dadda_pg_rca32_fa887_y1;
  wire f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa764_y2;
  wire f_s_dadda_pg_rca32_fa887_y2;
  wire f_s_dadda_pg_rca32_fa887_y3;
  wire f_s_dadda_pg_rca32_fa887_y4;
  wire f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa887_y4;
  wire f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa765_y2;
  wire f_s_dadda_pg_rca32_fa888_y0;
  wire f_s_dadda_pg_rca32_fa888_y1;
  wire f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa766_y2;
  wire f_s_dadda_pg_rca32_fa888_y2;
  wire f_s_dadda_pg_rca32_fa888_y3;
  wire f_s_dadda_pg_rca32_fa888_y4;
  wire f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa888_y4;
  wire f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa767_y2;
  wire f_s_dadda_pg_rca32_fa889_y0;
  wire f_s_dadda_pg_rca32_fa889_y1;
  wire f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa768_y2;
  wire f_s_dadda_pg_rca32_fa889_y2;
  wire f_s_dadda_pg_rca32_fa889_y3;
  wire f_s_dadda_pg_rca32_fa889_y4;
  wire f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa889_y4;
  wire f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa769_y2;
  wire f_s_dadda_pg_rca32_fa890_y0;
  wire f_s_dadda_pg_rca32_fa890_y1;
  wire f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa770_y2;
  wire f_s_dadda_pg_rca32_fa890_y2;
  wire f_s_dadda_pg_rca32_fa890_y3;
  wire f_s_dadda_pg_rca32_fa890_y4;
  wire f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa890_y4;
  wire f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa771_y2;
  wire f_s_dadda_pg_rca32_fa891_y0;
  wire f_s_dadda_pg_rca32_fa891_y1;
  wire f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa772_y2;
  wire f_s_dadda_pg_rca32_fa891_y2;
  wire f_s_dadda_pg_rca32_fa891_y3;
  wire f_s_dadda_pg_rca32_fa891_y4;
  wire f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa891_y4;
  wire f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa773_y2;
  wire f_s_dadda_pg_rca32_fa892_y0;
  wire f_s_dadda_pg_rca32_fa892_y1;
  wire f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa774_y2;
  wire f_s_dadda_pg_rca32_fa892_y2;
  wire f_s_dadda_pg_rca32_fa892_y3;
  wire f_s_dadda_pg_rca32_fa892_y4;
  wire f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa892_y4;
  wire f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa775_y2;
  wire f_s_dadda_pg_rca32_fa893_y0;
  wire f_s_dadda_pg_rca32_fa893_y1;
  wire f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa776_y2;
  wire f_s_dadda_pg_rca32_fa893_y2;
  wire f_s_dadda_pg_rca32_fa893_y3;
  wire f_s_dadda_pg_rca32_fa893_y4;
  wire f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa893_y4;
  wire f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa777_y2;
  wire f_s_dadda_pg_rca32_fa894_y0;
  wire f_s_dadda_pg_rca32_fa894_y1;
  wire f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa778_y2;
  wire f_s_dadda_pg_rca32_fa894_y2;
  wire f_s_dadda_pg_rca32_fa894_y3;
  wire f_s_dadda_pg_rca32_fa894_y4;
  wire f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa894_y4;
  wire f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa779_y2;
  wire f_s_dadda_pg_rca32_fa895_y0;
  wire f_s_dadda_pg_rca32_fa895_y1;
  wire f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa780_y2;
  wire f_s_dadda_pg_rca32_fa895_y2;
  wire f_s_dadda_pg_rca32_fa895_y3;
  wire f_s_dadda_pg_rca32_fa895_y4;
  wire f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa895_y4;
  wire f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa781_y2;
  wire f_s_dadda_pg_rca32_fa896_y0;
  wire f_s_dadda_pg_rca32_fa896_y1;
  wire f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa782_y2;
  wire f_s_dadda_pg_rca32_fa896_y2;
  wire f_s_dadda_pg_rca32_fa896_y3;
  wire f_s_dadda_pg_rca32_fa896_y4;
  wire f_s_dadda_pg_rca32_nand_28_31_a_28;
  wire f_s_dadda_pg_rca32_nand_28_31_b_31;
  wire f_s_dadda_pg_rca32_nand_28_31_y0;
  wire f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_fa896_y4;
  wire f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_nand_28_31_y0;
  wire f_s_dadda_pg_rca32_fa897_y0;
  wire f_s_dadda_pg_rca32_fa897_y1;
  wire f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_fa783_y2;
  wire f_s_dadda_pg_rca32_fa897_y2;
  wire f_s_dadda_pg_rca32_fa897_y3;
  wire f_s_dadda_pg_rca32_fa897_y4;
  wire f_s_dadda_pg_rca32_and_30_30_a_30;
  wire f_s_dadda_pg_rca32_and_30_30_b_30;
  wire f_s_dadda_pg_rca32_and_30_30_y0;
  wire f_s_dadda_pg_rca32_nand_29_31_a_29;
  wire f_s_dadda_pg_rca32_nand_29_31_b_31;
  wire f_s_dadda_pg_rca32_nand_29_31_y0;
  wire f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_fa897_y4;
  wire f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_and_30_30_y0;
  wire f_s_dadda_pg_rca32_fa898_y0;
  wire f_s_dadda_pg_rca32_fa898_y1;
  wire f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_nand_29_31_y0;
  wire f_s_dadda_pg_rca32_fa898_y2;
  wire f_s_dadda_pg_rca32_fa898_y3;
  wire f_s_dadda_pg_rca32_fa898_y4;
  wire f_s_dadda_pg_rca32_nand_31_30_a_31;
  wire f_s_dadda_pg_rca32_nand_31_30_b_30;
  wire f_s_dadda_pg_rca32_nand_31_30_y0;
  wire f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_fa898_y4;
  wire f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_fa840_y4;
  wire f_s_dadda_pg_rca32_fa899_y0;
  wire f_s_dadda_pg_rca32_fa899_y1;
  wire f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_nand_31_30_y0;
  wire f_s_dadda_pg_rca32_fa899_y2;
  wire f_s_dadda_pg_rca32_fa899_y3;
  wire f_s_dadda_pg_rca32_fa899_y4;
  wire f_s_dadda_pg_rca32_and_0_0_a_0;
  wire f_s_dadda_pg_rca32_and_0_0_b_0;
  wire f_s_dadda_pg_rca32_and_0_0_y0;
  wire f_s_dadda_pg_rca32_and_1_0_a_1;
  wire f_s_dadda_pg_rca32_and_1_0_b_0;
  wire f_s_dadda_pg_rca32_and_1_0_y0;
  wire f_s_dadda_pg_rca32_and_0_2_a_0;
  wire f_s_dadda_pg_rca32_and_0_2_b_2;
  wire f_s_dadda_pg_rca32_and_0_2_y0;
  wire f_s_dadda_pg_rca32_nand_30_31_a_30;
  wire f_s_dadda_pg_rca32_nand_30_31_b_31;
  wire f_s_dadda_pg_rca32_nand_30_31_y0;
  wire f_s_dadda_pg_rca32_and_0_1_a_0;
  wire f_s_dadda_pg_rca32_and_0_1_b_1;
  wire f_s_dadda_pg_rca32_and_0_1_y0;
  wire f_s_dadda_pg_rca32_and_31_31_a_31;
  wire f_s_dadda_pg_rca32_and_31_31_b_31;
  wire f_s_dadda_pg_rca32_and_31_31_y0;
  wire constant_wire_value_0_f_s_dadda_pg_rca32_and_1_0_y0;
  wire constant_wire_value_0_f_s_dadda_pg_rca32_and_0_1_y0;
  wire constant_wire_value_0_y0;
  wire constant_wire_value_0_y1;
  wire constant_wire_0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa0_f_s_dadda_pg_rca32_and_1_0_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa0_f_s_dadda_pg_rca32_and_0_1_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa0_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa0_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa0_constant_wire_0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa0_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and0_constant_wire_0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and0_f_s_dadda_pg_rca32_u_pg_rca_fa0_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and0_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or0_f_s_dadda_pg_rca32_u_pg_rca_and0_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or0_f_s_dadda_pg_rca32_u_pg_rca_fa0_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or0_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_and_0_2_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_ha29_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa1_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa1_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_u_pg_rca_or0_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa1_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and1_f_s_dadda_pg_rca32_u_pg_rca_or0_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and1_f_s_dadda_pg_rca32_u_pg_rca_fa1_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and1_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or1_f_s_dadda_pg_rca32_u_pg_rca_and1_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or1_f_s_dadda_pg_rca32_u_pg_rca_fa1_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or1_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_ha28_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_fa841_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa2_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa2_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_u_pg_rca_or1_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa2_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and2_f_s_dadda_pg_rca32_u_pg_rca_or1_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and2_f_s_dadda_pg_rca32_u_pg_rca_fa2_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and2_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or2_f_s_dadda_pg_rca32_u_pg_rca_and2_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or2_f_s_dadda_pg_rca32_u_pg_rca_fa2_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or2_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_fa784_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_fa842_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa3_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa3_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_u_pg_rca_or2_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa3_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and3_f_s_dadda_pg_rca32_u_pg_rca_or2_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and3_f_s_dadda_pg_rca32_u_pg_rca_fa3_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and3_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or3_f_s_dadda_pg_rca32_u_pg_rca_and3_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or3_f_s_dadda_pg_rca32_u_pg_rca_fa3_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or3_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_fa785_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_fa843_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa4_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa4_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_u_pg_rca_or3_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa4_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and4_f_s_dadda_pg_rca32_u_pg_rca_or3_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and4_f_s_dadda_pg_rca32_u_pg_rca_fa4_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and4_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or4_f_s_dadda_pg_rca32_u_pg_rca_and4_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or4_f_s_dadda_pg_rca32_u_pg_rca_fa4_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or4_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_fa786_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_fa844_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa5_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa5_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_u_pg_rca_or4_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa5_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and5_f_s_dadda_pg_rca32_u_pg_rca_or4_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and5_f_s_dadda_pg_rca32_u_pg_rca_fa5_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and5_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or5_f_s_dadda_pg_rca32_u_pg_rca_and5_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or5_f_s_dadda_pg_rca32_u_pg_rca_fa5_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or5_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_fa787_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_fa845_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa6_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa6_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_u_pg_rca_or5_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa6_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and6_f_s_dadda_pg_rca32_u_pg_rca_or5_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and6_f_s_dadda_pg_rca32_u_pg_rca_fa6_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and6_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or6_f_s_dadda_pg_rca32_u_pg_rca_and6_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or6_f_s_dadda_pg_rca32_u_pg_rca_fa6_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or6_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_fa788_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_fa846_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa7_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa7_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_u_pg_rca_or6_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa7_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and7_f_s_dadda_pg_rca32_u_pg_rca_or6_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and7_f_s_dadda_pg_rca32_u_pg_rca_fa7_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and7_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or7_f_s_dadda_pg_rca32_u_pg_rca_and7_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or7_f_s_dadda_pg_rca32_u_pg_rca_fa7_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or7_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_fa789_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_fa847_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa8_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa8_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_u_pg_rca_or7_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa8_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and8_f_s_dadda_pg_rca32_u_pg_rca_or7_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and8_f_s_dadda_pg_rca32_u_pg_rca_fa8_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and8_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or8_f_s_dadda_pg_rca32_u_pg_rca_and8_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or8_f_s_dadda_pg_rca32_u_pg_rca_fa8_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or8_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_fa790_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_fa848_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa9_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa9_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_u_pg_rca_or8_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa9_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and9_f_s_dadda_pg_rca32_u_pg_rca_or8_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and9_f_s_dadda_pg_rca32_u_pg_rca_fa9_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and9_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or9_f_s_dadda_pg_rca32_u_pg_rca_and9_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or9_f_s_dadda_pg_rca32_u_pg_rca_fa9_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or9_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_fa791_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_fa849_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa10_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa10_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_u_pg_rca_or9_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa10_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and10_f_s_dadda_pg_rca32_u_pg_rca_or9_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and10_f_s_dadda_pg_rca32_u_pg_rca_fa10_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and10_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or10_f_s_dadda_pg_rca32_u_pg_rca_and10_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or10_f_s_dadda_pg_rca32_u_pg_rca_fa10_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or10_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_fa792_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_fa850_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa11_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa11_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_u_pg_rca_or10_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa11_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and11_f_s_dadda_pg_rca32_u_pg_rca_or10_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and11_f_s_dadda_pg_rca32_u_pg_rca_fa11_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and11_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or11_f_s_dadda_pg_rca32_u_pg_rca_and11_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or11_f_s_dadda_pg_rca32_u_pg_rca_fa11_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or11_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_fa793_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_fa851_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa12_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa12_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_u_pg_rca_or11_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa12_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and12_f_s_dadda_pg_rca32_u_pg_rca_or11_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and12_f_s_dadda_pg_rca32_u_pg_rca_fa12_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and12_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or12_f_s_dadda_pg_rca32_u_pg_rca_and12_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or12_f_s_dadda_pg_rca32_u_pg_rca_fa12_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or12_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_fa794_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_fa852_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa13_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa13_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_u_pg_rca_or12_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa13_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and13_f_s_dadda_pg_rca32_u_pg_rca_or12_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and13_f_s_dadda_pg_rca32_u_pg_rca_fa13_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and13_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or13_f_s_dadda_pg_rca32_u_pg_rca_and13_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or13_f_s_dadda_pg_rca32_u_pg_rca_fa13_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or13_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_fa795_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_fa853_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa14_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa14_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_u_pg_rca_or13_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa14_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and14_f_s_dadda_pg_rca32_u_pg_rca_or13_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and14_f_s_dadda_pg_rca32_u_pg_rca_fa14_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and14_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or14_f_s_dadda_pg_rca32_u_pg_rca_and14_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or14_f_s_dadda_pg_rca32_u_pg_rca_fa14_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or14_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_fa796_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_fa854_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa15_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa15_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_u_pg_rca_or14_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa15_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and15_f_s_dadda_pg_rca32_u_pg_rca_or14_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and15_f_s_dadda_pg_rca32_u_pg_rca_fa15_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and15_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or15_f_s_dadda_pg_rca32_u_pg_rca_and15_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or15_f_s_dadda_pg_rca32_u_pg_rca_fa15_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or15_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_fa797_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_fa855_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa16_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa16_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_u_pg_rca_or15_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa16_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and16_f_s_dadda_pg_rca32_u_pg_rca_or15_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and16_f_s_dadda_pg_rca32_u_pg_rca_fa16_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and16_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or16_f_s_dadda_pg_rca32_u_pg_rca_and16_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or16_f_s_dadda_pg_rca32_u_pg_rca_fa16_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or16_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_fa798_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_fa856_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa17_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa17_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_u_pg_rca_or16_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa17_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and17_f_s_dadda_pg_rca32_u_pg_rca_or16_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and17_f_s_dadda_pg_rca32_u_pg_rca_fa17_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and17_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or17_f_s_dadda_pg_rca32_u_pg_rca_and17_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or17_f_s_dadda_pg_rca32_u_pg_rca_fa17_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or17_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_fa799_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_fa857_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa18_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa18_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_u_pg_rca_or17_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa18_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and18_f_s_dadda_pg_rca32_u_pg_rca_or17_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and18_f_s_dadda_pg_rca32_u_pg_rca_fa18_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and18_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or18_f_s_dadda_pg_rca32_u_pg_rca_and18_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or18_f_s_dadda_pg_rca32_u_pg_rca_fa18_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or18_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_fa800_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_fa858_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa19_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa19_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_u_pg_rca_or18_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa19_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and19_f_s_dadda_pg_rca32_u_pg_rca_or18_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and19_f_s_dadda_pg_rca32_u_pg_rca_fa19_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and19_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or19_f_s_dadda_pg_rca32_u_pg_rca_and19_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or19_f_s_dadda_pg_rca32_u_pg_rca_fa19_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or19_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_fa801_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_fa859_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa20_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa20_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_u_pg_rca_or19_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa20_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and20_f_s_dadda_pg_rca32_u_pg_rca_or19_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and20_f_s_dadda_pg_rca32_u_pg_rca_fa20_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and20_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or20_f_s_dadda_pg_rca32_u_pg_rca_and20_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or20_f_s_dadda_pg_rca32_u_pg_rca_fa20_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or20_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_fa802_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_fa860_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa21_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa21_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_u_pg_rca_or20_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa21_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and21_f_s_dadda_pg_rca32_u_pg_rca_or20_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and21_f_s_dadda_pg_rca32_u_pg_rca_fa21_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and21_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or21_f_s_dadda_pg_rca32_u_pg_rca_and21_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or21_f_s_dadda_pg_rca32_u_pg_rca_fa21_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or21_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_fa803_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_fa861_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa22_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa22_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_u_pg_rca_or21_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa22_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and22_f_s_dadda_pg_rca32_u_pg_rca_or21_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and22_f_s_dadda_pg_rca32_u_pg_rca_fa22_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and22_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or22_f_s_dadda_pg_rca32_u_pg_rca_and22_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or22_f_s_dadda_pg_rca32_u_pg_rca_fa22_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or22_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_fa804_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_fa862_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa23_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa23_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_u_pg_rca_or22_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa23_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and23_f_s_dadda_pg_rca32_u_pg_rca_or22_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and23_f_s_dadda_pg_rca32_u_pg_rca_fa23_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and23_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or23_f_s_dadda_pg_rca32_u_pg_rca_and23_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or23_f_s_dadda_pg_rca32_u_pg_rca_fa23_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or23_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_fa805_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_fa863_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa24_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa24_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_u_pg_rca_or23_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa24_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and24_f_s_dadda_pg_rca32_u_pg_rca_or23_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and24_f_s_dadda_pg_rca32_u_pg_rca_fa24_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and24_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or24_f_s_dadda_pg_rca32_u_pg_rca_and24_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or24_f_s_dadda_pg_rca32_u_pg_rca_fa24_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or24_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_fa806_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_fa864_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa25_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa25_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_u_pg_rca_or24_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa25_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and25_f_s_dadda_pg_rca32_u_pg_rca_or24_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and25_f_s_dadda_pg_rca32_u_pg_rca_fa25_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and25_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or25_f_s_dadda_pg_rca32_u_pg_rca_and25_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or25_f_s_dadda_pg_rca32_u_pg_rca_fa25_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or25_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_fa807_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_fa865_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa26_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa26_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_u_pg_rca_or25_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa26_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and26_f_s_dadda_pg_rca32_u_pg_rca_or25_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and26_f_s_dadda_pg_rca32_u_pg_rca_fa26_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and26_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or26_f_s_dadda_pg_rca32_u_pg_rca_and26_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or26_f_s_dadda_pg_rca32_u_pg_rca_fa26_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or26_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_fa808_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_fa866_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa27_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa27_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_u_pg_rca_or26_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa27_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and27_f_s_dadda_pg_rca32_u_pg_rca_or26_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and27_f_s_dadda_pg_rca32_u_pg_rca_fa27_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and27_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or27_f_s_dadda_pg_rca32_u_pg_rca_and27_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or27_f_s_dadda_pg_rca32_u_pg_rca_fa27_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or27_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_fa809_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_fa867_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa28_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa28_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_u_pg_rca_or27_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa28_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and28_f_s_dadda_pg_rca32_u_pg_rca_or27_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and28_f_s_dadda_pg_rca32_u_pg_rca_fa28_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and28_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or28_f_s_dadda_pg_rca32_u_pg_rca_and28_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or28_f_s_dadda_pg_rca32_u_pg_rca_fa28_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or28_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_fa810_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_fa868_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa29_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa29_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_u_pg_rca_or28_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa29_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and29_f_s_dadda_pg_rca32_u_pg_rca_or28_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and29_f_s_dadda_pg_rca32_u_pg_rca_fa29_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and29_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or29_f_s_dadda_pg_rca32_u_pg_rca_and29_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or29_f_s_dadda_pg_rca32_u_pg_rca_fa29_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or29_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_fa811_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_fa869_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa30_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa30_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_u_pg_rca_or29_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa30_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and30_f_s_dadda_pg_rca32_u_pg_rca_or29_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and30_f_s_dadda_pg_rca32_u_pg_rca_fa30_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and30_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or30_f_s_dadda_pg_rca32_u_pg_rca_and30_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or30_f_s_dadda_pg_rca32_u_pg_rca_fa30_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or30_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_fa812_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_fa870_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa31_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_u_pg_rca_or30_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa31_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and31_f_s_dadda_pg_rca32_u_pg_rca_or30_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and31_f_s_dadda_pg_rca32_u_pg_rca_fa31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or31_f_s_dadda_pg_rca32_u_pg_rca_and31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or31_f_s_dadda_pg_rca32_u_pg_rca_fa31_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_fa813_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_fa871_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa32_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa32_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_u_pg_rca_or31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa32_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and32_f_s_dadda_pg_rca32_u_pg_rca_or31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and32_f_s_dadda_pg_rca32_u_pg_rca_fa32_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and32_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or32_f_s_dadda_pg_rca32_u_pg_rca_and32_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or32_f_s_dadda_pg_rca32_u_pg_rca_fa32_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or32_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_fa814_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_fa872_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa33_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa33_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_u_pg_rca_or32_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa33_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and33_f_s_dadda_pg_rca32_u_pg_rca_or32_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and33_f_s_dadda_pg_rca32_u_pg_rca_fa33_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and33_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or33_f_s_dadda_pg_rca32_u_pg_rca_and33_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or33_f_s_dadda_pg_rca32_u_pg_rca_fa33_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or33_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_fa815_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_fa873_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa34_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa34_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_u_pg_rca_or33_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa34_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and34_f_s_dadda_pg_rca32_u_pg_rca_or33_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and34_f_s_dadda_pg_rca32_u_pg_rca_fa34_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and34_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or34_f_s_dadda_pg_rca32_u_pg_rca_and34_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or34_f_s_dadda_pg_rca32_u_pg_rca_fa34_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or34_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_fa816_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_fa874_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa35_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa35_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_u_pg_rca_or34_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa35_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and35_f_s_dadda_pg_rca32_u_pg_rca_or34_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and35_f_s_dadda_pg_rca32_u_pg_rca_fa35_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and35_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or35_f_s_dadda_pg_rca32_u_pg_rca_and35_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or35_f_s_dadda_pg_rca32_u_pg_rca_fa35_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or35_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_fa817_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_fa875_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa36_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa36_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_u_pg_rca_or35_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa36_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and36_f_s_dadda_pg_rca32_u_pg_rca_or35_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and36_f_s_dadda_pg_rca32_u_pg_rca_fa36_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and36_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or36_f_s_dadda_pg_rca32_u_pg_rca_and36_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or36_f_s_dadda_pg_rca32_u_pg_rca_fa36_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or36_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_fa818_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_fa876_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa37_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa37_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_u_pg_rca_or36_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa37_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and37_f_s_dadda_pg_rca32_u_pg_rca_or36_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and37_f_s_dadda_pg_rca32_u_pg_rca_fa37_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and37_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or37_f_s_dadda_pg_rca32_u_pg_rca_and37_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or37_f_s_dadda_pg_rca32_u_pg_rca_fa37_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or37_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_fa819_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_fa877_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa38_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa38_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_u_pg_rca_or37_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa38_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and38_f_s_dadda_pg_rca32_u_pg_rca_or37_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and38_f_s_dadda_pg_rca32_u_pg_rca_fa38_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and38_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or38_f_s_dadda_pg_rca32_u_pg_rca_and38_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or38_f_s_dadda_pg_rca32_u_pg_rca_fa38_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or38_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_fa820_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_fa878_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa39_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa39_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_u_pg_rca_or38_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa39_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and39_f_s_dadda_pg_rca32_u_pg_rca_or38_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and39_f_s_dadda_pg_rca32_u_pg_rca_fa39_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and39_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or39_f_s_dadda_pg_rca32_u_pg_rca_and39_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or39_f_s_dadda_pg_rca32_u_pg_rca_fa39_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or39_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_fa821_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_fa879_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa40_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa40_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_u_pg_rca_or39_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa40_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and40_f_s_dadda_pg_rca32_u_pg_rca_or39_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and40_f_s_dadda_pg_rca32_u_pg_rca_fa40_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and40_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or40_f_s_dadda_pg_rca32_u_pg_rca_and40_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or40_f_s_dadda_pg_rca32_u_pg_rca_fa40_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or40_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_fa822_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_fa880_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa41_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa41_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_u_pg_rca_or40_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa41_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and41_f_s_dadda_pg_rca32_u_pg_rca_or40_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and41_f_s_dadda_pg_rca32_u_pg_rca_fa41_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and41_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or41_f_s_dadda_pg_rca32_u_pg_rca_and41_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or41_f_s_dadda_pg_rca32_u_pg_rca_fa41_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or41_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_fa823_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_fa881_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa42_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa42_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_u_pg_rca_or41_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa42_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and42_f_s_dadda_pg_rca32_u_pg_rca_or41_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and42_f_s_dadda_pg_rca32_u_pg_rca_fa42_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and42_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or42_f_s_dadda_pg_rca32_u_pg_rca_and42_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or42_f_s_dadda_pg_rca32_u_pg_rca_fa42_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or42_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_fa824_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_fa882_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa43_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa43_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_u_pg_rca_or42_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa43_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and43_f_s_dadda_pg_rca32_u_pg_rca_or42_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and43_f_s_dadda_pg_rca32_u_pg_rca_fa43_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and43_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or43_f_s_dadda_pg_rca32_u_pg_rca_and43_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or43_f_s_dadda_pg_rca32_u_pg_rca_fa43_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or43_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_fa825_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_fa883_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa44_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa44_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_u_pg_rca_or43_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa44_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and44_f_s_dadda_pg_rca32_u_pg_rca_or43_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and44_f_s_dadda_pg_rca32_u_pg_rca_fa44_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and44_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or44_f_s_dadda_pg_rca32_u_pg_rca_and44_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or44_f_s_dadda_pg_rca32_u_pg_rca_fa44_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or44_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_fa826_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_fa884_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa45_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa45_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_u_pg_rca_or44_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa45_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and45_f_s_dadda_pg_rca32_u_pg_rca_or44_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and45_f_s_dadda_pg_rca32_u_pg_rca_fa45_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and45_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or45_f_s_dadda_pg_rca32_u_pg_rca_and45_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or45_f_s_dadda_pg_rca32_u_pg_rca_fa45_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or45_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_fa827_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_fa885_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa46_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa46_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_u_pg_rca_or45_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa46_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and46_f_s_dadda_pg_rca32_u_pg_rca_or45_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and46_f_s_dadda_pg_rca32_u_pg_rca_fa46_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and46_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or46_f_s_dadda_pg_rca32_u_pg_rca_and46_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or46_f_s_dadda_pg_rca32_u_pg_rca_fa46_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or46_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_fa828_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_fa886_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa47_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa47_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_u_pg_rca_or46_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa47_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and47_f_s_dadda_pg_rca32_u_pg_rca_or46_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and47_f_s_dadda_pg_rca32_u_pg_rca_fa47_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and47_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or47_f_s_dadda_pg_rca32_u_pg_rca_and47_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or47_f_s_dadda_pg_rca32_u_pg_rca_fa47_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or47_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_fa829_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_fa887_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa48_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa48_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_u_pg_rca_or47_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa48_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and48_f_s_dadda_pg_rca32_u_pg_rca_or47_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and48_f_s_dadda_pg_rca32_u_pg_rca_fa48_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and48_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or48_f_s_dadda_pg_rca32_u_pg_rca_and48_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or48_f_s_dadda_pg_rca32_u_pg_rca_fa48_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or48_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_fa830_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_fa888_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa49_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa49_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_u_pg_rca_or48_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa49_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and49_f_s_dadda_pg_rca32_u_pg_rca_or48_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and49_f_s_dadda_pg_rca32_u_pg_rca_fa49_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and49_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or49_f_s_dadda_pg_rca32_u_pg_rca_and49_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or49_f_s_dadda_pg_rca32_u_pg_rca_fa49_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or49_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_fa831_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_fa889_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa50_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa50_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_u_pg_rca_or49_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa50_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and50_f_s_dadda_pg_rca32_u_pg_rca_or49_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and50_f_s_dadda_pg_rca32_u_pg_rca_fa50_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and50_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or50_f_s_dadda_pg_rca32_u_pg_rca_and50_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or50_f_s_dadda_pg_rca32_u_pg_rca_fa50_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or50_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_fa832_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_fa890_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa51_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa51_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_u_pg_rca_or50_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa51_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and51_f_s_dadda_pg_rca32_u_pg_rca_or50_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and51_f_s_dadda_pg_rca32_u_pg_rca_fa51_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and51_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or51_f_s_dadda_pg_rca32_u_pg_rca_and51_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or51_f_s_dadda_pg_rca32_u_pg_rca_fa51_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or51_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_fa833_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_fa891_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa52_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa52_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_u_pg_rca_or51_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa52_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and52_f_s_dadda_pg_rca32_u_pg_rca_or51_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and52_f_s_dadda_pg_rca32_u_pg_rca_fa52_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and52_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or52_f_s_dadda_pg_rca32_u_pg_rca_and52_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or52_f_s_dadda_pg_rca32_u_pg_rca_fa52_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or52_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_fa834_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_fa892_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa53_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa53_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_u_pg_rca_or52_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa53_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and53_f_s_dadda_pg_rca32_u_pg_rca_or52_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and53_f_s_dadda_pg_rca32_u_pg_rca_fa53_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and53_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or53_f_s_dadda_pg_rca32_u_pg_rca_and53_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or53_f_s_dadda_pg_rca32_u_pg_rca_fa53_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or53_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_fa835_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_fa893_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa54_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa54_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_u_pg_rca_or53_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa54_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and54_f_s_dadda_pg_rca32_u_pg_rca_or53_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and54_f_s_dadda_pg_rca32_u_pg_rca_fa54_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and54_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or54_f_s_dadda_pg_rca32_u_pg_rca_and54_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or54_f_s_dadda_pg_rca32_u_pg_rca_fa54_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or54_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_fa836_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_fa894_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa55_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa55_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_u_pg_rca_or54_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa55_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and55_f_s_dadda_pg_rca32_u_pg_rca_or54_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and55_f_s_dadda_pg_rca32_u_pg_rca_fa55_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and55_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or55_f_s_dadda_pg_rca32_u_pg_rca_and55_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or55_f_s_dadda_pg_rca32_u_pg_rca_fa55_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or55_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_fa837_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_fa895_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa56_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa56_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_u_pg_rca_or55_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa56_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and56_f_s_dadda_pg_rca32_u_pg_rca_or55_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and56_f_s_dadda_pg_rca32_u_pg_rca_fa56_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and56_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or56_f_s_dadda_pg_rca32_u_pg_rca_and56_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or56_f_s_dadda_pg_rca32_u_pg_rca_fa56_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or56_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_fa838_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_fa896_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa57_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa57_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_u_pg_rca_or56_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa57_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and57_f_s_dadda_pg_rca32_u_pg_rca_or56_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and57_f_s_dadda_pg_rca32_u_pg_rca_fa57_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and57_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or57_f_s_dadda_pg_rca32_u_pg_rca_and57_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or57_f_s_dadda_pg_rca32_u_pg_rca_fa57_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or57_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_fa839_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_fa897_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa58_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa58_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_u_pg_rca_or57_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa58_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and58_f_s_dadda_pg_rca32_u_pg_rca_or57_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and58_f_s_dadda_pg_rca32_u_pg_rca_fa58_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and58_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or58_f_s_dadda_pg_rca32_u_pg_rca_and58_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or58_f_s_dadda_pg_rca32_u_pg_rca_fa58_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or58_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_fa840_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_fa898_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa59_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa59_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_u_pg_rca_or58_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa59_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and59_f_s_dadda_pg_rca32_u_pg_rca_or58_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and59_f_s_dadda_pg_rca32_u_pg_rca_fa59_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and59_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or59_f_s_dadda_pg_rca32_u_pg_rca_and59_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or59_f_s_dadda_pg_rca32_u_pg_rca_fa59_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or59_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_nand_30_31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_fa899_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa60_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa60_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_u_pg_rca_or59_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa60_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and60_f_s_dadda_pg_rca32_u_pg_rca_or59_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and60_f_s_dadda_pg_rca32_u_pg_rca_fa60_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and60_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or60_f_s_dadda_pg_rca32_u_pg_rca_and60_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or60_f_s_dadda_pg_rca32_u_pg_rca_fa60_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or60_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_fa899_y4;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_and_31_31_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa61_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa61_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_u_pg_rca_or60_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_fa61_y2;
  wire f_s_dadda_pg_rca32_u_pg_rca_and61_f_s_dadda_pg_rca32_u_pg_rca_or60_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and61_f_s_dadda_pg_rca32_u_pg_rca_fa61_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_and61_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or61_f_s_dadda_pg_rca32_u_pg_rca_and61_y0;
  wire f_s_dadda_pg_rca32_u_pg_rca_or61_f_s_dadda_pg_rca32_u_pg_rca_fa61_y1;
  wire f_s_dadda_pg_rca32_u_pg_rca_or61_y0;
  wire f_s_dadda_pg_rca32_xor0_constant_wire_1;
  wire f_s_dadda_pg_rca32_xor0_f_s_dadda_pg_rca32_u_pg_rca_or61_y0;
  wire f_s_dadda_pg_rca32_xor0_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign a_24 = a[24];
  assign a_25 = a[25];
  assign a_26 = a[26];
  assign a_27 = a[27];
  assign a_28 = a[28];
  assign a_29 = a[29];
  assign a_30 = a[30];
  assign a_31 = a[31];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign b_24 = b[24];
  assign b_25 = b[25];
  assign b_26 = b[26];
  assign b_27 = b[27];
  assign b_28 = b[28];
  assign b_29 = b[29];
  assign b_30 = b[30];
  assign b_31 = b[31];
  assign constant_wire_value_1_a_0 = a_0;
  assign constant_wire_value_1_b_0 = b_0;
  assign constant_wire_value_1_y0 = constant_wire_value_1_a_0 ^ constant_wire_value_1_b_0;
  assign constant_wire_value_1_y1 = ~(constant_wire_value_1_a_0 ^ constant_wire_value_1_b_0);
  assign constant_wire_1 = constant_wire_value_1_y0 | constant_wire_value_1_y1;
  assign f_s_dadda_pg_rca32_and_28_0_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_28_0_y0 = f_s_dadda_pg_rca32_and_28_0_a_28 & f_s_dadda_pg_rca32_and_28_0_b_0;
  assign f_s_dadda_pg_rca32_and_27_1_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_27_1_y0 = f_s_dadda_pg_rca32_and_27_1_a_27 & f_s_dadda_pg_rca32_and_27_1_b_1;
  assign f_s_dadda_pg_rca32_ha0_f_s_dadda_pg_rca32_and_28_0_y0 = f_s_dadda_pg_rca32_and_28_0_y0;
  assign f_s_dadda_pg_rca32_ha0_f_s_dadda_pg_rca32_and_27_1_y0 = f_s_dadda_pg_rca32_and_27_1_y0;
  assign f_s_dadda_pg_rca32_ha0_y0 = f_s_dadda_pg_rca32_ha0_f_s_dadda_pg_rca32_and_28_0_y0 ^ f_s_dadda_pg_rca32_ha0_f_s_dadda_pg_rca32_and_27_1_y0;
  assign f_s_dadda_pg_rca32_ha0_y1 = f_s_dadda_pg_rca32_ha0_f_s_dadda_pg_rca32_and_28_0_y0 & f_s_dadda_pg_rca32_ha0_f_s_dadda_pg_rca32_and_27_1_y0;
  assign f_s_dadda_pg_rca32_and_29_0_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_29_0_y0 = f_s_dadda_pg_rca32_and_29_0_a_29 & f_s_dadda_pg_rca32_and_29_0_b_0;
  assign f_s_dadda_pg_rca32_and_28_1_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_28_1_y0 = f_s_dadda_pg_rca32_and_28_1_a_28 & f_s_dadda_pg_rca32_and_28_1_b_1;
  assign f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_ha0_y1 = f_s_dadda_pg_rca32_ha0_y1;
  assign f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_and_29_0_y0 = f_s_dadda_pg_rca32_and_29_0_y0;
  assign f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_and_28_1_y0 = f_s_dadda_pg_rca32_and_28_1_y0;
  assign f_s_dadda_pg_rca32_fa0_y0 = f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_ha0_y1 ^ f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_and_29_0_y0;
  assign f_s_dadda_pg_rca32_fa0_y1 = f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_ha0_y1 & f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_and_29_0_y0;
  assign f_s_dadda_pg_rca32_fa0_y2 = f_s_dadda_pg_rca32_fa0_y0 ^ f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_and_28_1_y0;
  assign f_s_dadda_pg_rca32_fa0_y3 = f_s_dadda_pg_rca32_fa0_y0 & f_s_dadda_pg_rca32_fa0_f_s_dadda_pg_rca32_and_28_1_y0;
  assign f_s_dadda_pg_rca32_fa0_y4 = f_s_dadda_pg_rca32_fa0_y1 | f_s_dadda_pg_rca32_fa0_y3;
  assign f_s_dadda_pg_rca32_and_27_2_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_27_2_y0 = f_s_dadda_pg_rca32_and_27_2_a_27 & f_s_dadda_pg_rca32_and_27_2_b_2;
  assign f_s_dadda_pg_rca32_and_26_3_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_26_3_y0 = f_s_dadda_pg_rca32_and_26_3_a_26 & f_s_dadda_pg_rca32_and_26_3_b_3;
  assign f_s_dadda_pg_rca32_ha1_f_s_dadda_pg_rca32_and_27_2_y0 = f_s_dadda_pg_rca32_and_27_2_y0;
  assign f_s_dadda_pg_rca32_ha1_f_s_dadda_pg_rca32_and_26_3_y0 = f_s_dadda_pg_rca32_and_26_3_y0;
  assign f_s_dadda_pg_rca32_ha1_y0 = f_s_dadda_pg_rca32_ha1_f_s_dadda_pg_rca32_and_27_2_y0 ^ f_s_dadda_pg_rca32_ha1_f_s_dadda_pg_rca32_and_26_3_y0;
  assign f_s_dadda_pg_rca32_ha1_y1 = f_s_dadda_pg_rca32_ha1_f_s_dadda_pg_rca32_and_27_2_y0 & f_s_dadda_pg_rca32_ha1_f_s_dadda_pg_rca32_and_26_3_y0;
  assign f_s_dadda_pg_rca32_and_30_0_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_30_0_y0 = f_s_dadda_pg_rca32_and_30_0_a_30 & f_s_dadda_pg_rca32_and_30_0_b_0;
  assign f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_ha1_y1 = f_s_dadda_pg_rca32_ha1_y1;
  assign f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_fa0_y4 = f_s_dadda_pg_rca32_fa0_y4;
  assign f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_and_30_0_y0 = f_s_dadda_pg_rca32_and_30_0_y0;
  assign f_s_dadda_pg_rca32_fa1_y0 = f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_ha1_y1 ^ f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_fa0_y4;
  assign f_s_dadda_pg_rca32_fa1_y1 = f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_ha1_y1 & f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_fa0_y4;
  assign f_s_dadda_pg_rca32_fa1_y2 = f_s_dadda_pg_rca32_fa1_y0 ^ f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_and_30_0_y0;
  assign f_s_dadda_pg_rca32_fa1_y3 = f_s_dadda_pg_rca32_fa1_y0 & f_s_dadda_pg_rca32_fa1_f_s_dadda_pg_rca32_and_30_0_y0;
  assign f_s_dadda_pg_rca32_fa1_y4 = f_s_dadda_pg_rca32_fa1_y1 | f_s_dadda_pg_rca32_fa1_y3;
  assign f_s_dadda_pg_rca32_and_29_1_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_29_1_y0 = f_s_dadda_pg_rca32_and_29_1_a_29 & f_s_dadda_pg_rca32_and_29_1_b_1;
  assign f_s_dadda_pg_rca32_and_28_2_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_28_2_y0 = f_s_dadda_pg_rca32_and_28_2_a_28 & f_s_dadda_pg_rca32_and_28_2_b_2;
  assign f_s_dadda_pg_rca32_and_27_3_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_27_3_y0 = f_s_dadda_pg_rca32_and_27_3_a_27 & f_s_dadda_pg_rca32_and_27_3_b_3;
  assign f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_29_1_y0 = f_s_dadda_pg_rca32_and_29_1_y0;
  assign f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_28_2_y0 = f_s_dadda_pg_rca32_and_28_2_y0;
  assign f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_27_3_y0 = f_s_dadda_pg_rca32_and_27_3_y0;
  assign f_s_dadda_pg_rca32_fa2_y0 = f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_29_1_y0 ^ f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_28_2_y0;
  assign f_s_dadda_pg_rca32_fa2_y1 = f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_29_1_y0 & f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_28_2_y0;
  assign f_s_dadda_pg_rca32_fa2_y2 = f_s_dadda_pg_rca32_fa2_y0 ^ f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_27_3_y0;
  assign f_s_dadda_pg_rca32_fa2_y3 = f_s_dadda_pg_rca32_fa2_y0 & f_s_dadda_pg_rca32_fa2_f_s_dadda_pg_rca32_and_27_3_y0;
  assign f_s_dadda_pg_rca32_fa2_y4 = f_s_dadda_pg_rca32_fa2_y1 | f_s_dadda_pg_rca32_fa2_y3;
  assign f_s_dadda_pg_rca32_and_26_4_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_26_4_y0 = f_s_dadda_pg_rca32_and_26_4_a_26 & f_s_dadda_pg_rca32_and_26_4_b_4;
  assign f_s_dadda_pg_rca32_and_25_5_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_25_5_y0 = f_s_dadda_pg_rca32_and_25_5_a_25 & f_s_dadda_pg_rca32_and_25_5_b_5;
  assign f_s_dadda_pg_rca32_ha2_f_s_dadda_pg_rca32_and_26_4_y0 = f_s_dadda_pg_rca32_and_26_4_y0;
  assign f_s_dadda_pg_rca32_ha2_f_s_dadda_pg_rca32_and_25_5_y0 = f_s_dadda_pg_rca32_and_25_5_y0;
  assign f_s_dadda_pg_rca32_ha2_y0 = f_s_dadda_pg_rca32_ha2_f_s_dadda_pg_rca32_and_26_4_y0 ^ f_s_dadda_pg_rca32_ha2_f_s_dadda_pg_rca32_and_25_5_y0;
  assign f_s_dadda_pg_rca32_ha2_y1 = f_s_dadda_pg_rca32_ha2_f_s_dadda_pg_rca32_and_26_4_y0 & f_s_dadda_pg_rca32_ha2_f_s_dadda_pg_rca32_and_25_5_y0;
  assign f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_ha2_y1 = f_s_dadda_pg_rca32_ha2_y1;
  assign f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_fa2_y4 = f_s_dadda_pg_rca32_fa2_y4;
  assign f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_fa1_y4 = f_s_dadda_pg_rca32_fa1_y4;
  assign f_s_dadda_pg_rca32_fa3_y0 = f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_ha2_y1 ^ f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_fa2_y4;
  assign f_s_dadda_pg_rca32_fa3_y1 = f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_ha2_y1 & f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_fa2_y4;
  assign f_s_dadda_pg_rca32_fa3_y2 = f_s_dadda_pg_rca32_fa3_y0 ^ f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_fa1_y4;
  assign f_s_dadda_pg_rca32_fa3_y3 = f_s_dadda_pg_rca32_fa3_y0 & f_s_dadda_pg_rca32_fa3_f_s_dadda_pg_rca32_fa1_y4;
  assign f_s_dadda_pg_rca32_fa3_y4 = f_s_dadda_pg_rca32_fa3_y1 | f_s_dadda_pg_rca32_fa3_y3;
  assign f_s_dadda_pg_rca32_nand_31_0_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_nand_31_0_y0 = ~(f_s_dadda_pg_rca32_nand_31_0_a_31 & f_s_dadda_pg_rca32_nand_31_0_b_0);
  assign f_s_dadda_pg_rca32_and_30_1_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_30_1_y0 = f_s_dadda_pg_rca32_and_30_1_a_30 & f_s_dadda_pg_rca32_and_30_1_b_1;
  assign f_s_dadda_pg_rca32_and_29_2_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_29_2_y0 = f_s_dadda_pg_rca32_and_29_2_a_29 & f_s_dadda_pg_rca32_and_29_2_b_2;
  assign f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_nand_31_0_y0 = f_s_dadda_pg_rca32_nand_31_0_y0;
  assign f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_and_30_1_y0 = f_s_dadda_pg_rca32_and_30_1_y0;
  assign f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_and_29_2_y0 = f_s_dadda_pg_rca32_and_29_2_y0;
  assign f_s_dadda_pg_rca32_fa4_y0 = f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_nand_31_0_y0 ^ f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_and_30_1_y0;
  assign f_s_dadda_pg_rca32_fa4_y1 = f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_nand_31_0_y0 & f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_and_30_1_y0;
  assign f_s_dadda_pg_rca32_fa4_y2 = f_s_dadda_pg_rca32_fa4_y0 ^ f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_and_29_2_y0;
  assign f_s_dadda_pg_rca32_fa4_y3 = f_s_dadda_pg_rca32_fa4_y0 & f_s_dadda_pg_rca32_fa4_f_s_dadda_pg_rca32_and_29_2_y0;
  assign f_s_dadda_pg_rca32_fa4_y4 = f_s_dadda_pg_rca32_fa4_y1 | f_s_dadda_pg_rca32_fa4_y3;
  assign f_s_dadda_pg_rca32_and_28_3_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_28_3_y0 = f_s_dadda_pg_rca32_and_28_3_a_28 & f_s_dadda_pg_rca32_and_28_3_b_3;
  assign f_s_dadda_pg_rca32_and_27_4_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_27_4_y0 = f_s_dadda_pg_rca32_and_27_4_a_27 & f_s_dadda_pg_rca32_and_27_4_b_4;
  assign f_s_dadda_pg_rca32_and_26_5_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_26_5_y0 = f_s_dadda_pg_rca32_and_26_5_a_26 & f_s_dadda_pg_rca32_and_26_5_b_5;
  assign f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_28_3_y0 = f_s_dadda_pg_rca32_and_28_3_y0;
  assign f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_27_4_y0 = f_s_dadda_pg_rca32_and_27_4_y0;
  assign f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_26_5_y0 = f_s_dadda_pg_rca32_and_26_5_y0;
  assign f_s_dadda_pg_rca32_fa5_y0 = f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_28_3_y0 ^ f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_27_4_y0;
  assign f_s_dadda_pg_rca32_fa5_y1 = f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_28_3_y0 & f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_27_4_y0;
  assign f_s_dadda_pg_rca32_fa5_y2 = f_s_dadda_pg_rca32_fa5_y0 ^ f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_26_5_y0;
  assign f_s_dadda_pg_rca32_fa5_y3 = f_s_dadda_pg_rca32_fa5_y0 & f_s_dadda_pg_rca32_fa5_f_s_dadda_pg_rca32_and_26_5_y0;
  assign f_s_dadda_pg_rca32_fa5_y4 = f_s_dadda_pg_rca32_fa5_y1 | f_s_dadda_pg_rca32_fa5_y3;
  assign f_s_dadda_pg_rca32_and_25_6_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_25_6_y0 = f_s_dadda_pg_rca32_and_25_6_a_25 & f_s_dadda_pg_rca32_and_25_6_b_6;
  assign f_s_dadda_pg_rca32_and_24_7_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_24_7_y0 = f_s_dadda_pg_rca32_and_24_7_a_24 & f_s_dadda_pg_rca32_and_24_7_b_7;
  assign f_s_dadda_pg_rca32_ha3_f_s_dadda_pg_rca32_and_25_6_y0 = f_s_dadda_pg_rca32_and_25_6_y0;
  assign f_s_dadda_pg_rca32_ha3_f_s_dadda_pg_rca32_and_24_7_y0 = f_s_dadda_pg_rca32_and_24_7_y0;
  assign f_s_dadda_pg_rca32_ha3_y0 = f_s_dadda_pg_rca32_ha3_f_s_dadda_pg_rca32_and_25_6_y0 ^ f_s_dadda_pg_rca32_ha3_f_s_dadda_pg_rca32_and_24_7_y0;
  assign f_s_dadda_pg_rca32_ha3_y1 = f_s_dadda_pg_rca32_ha3_f_s_dadda_pg_rca32_and_25_6_y0 & f_s_dadda_pg_rca32_ha3_f_s_dadda_pg_rca32_and_24_7_y0;
  assign f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_ha3_y1 = f_s_dadda_pg_rca32_ha3_y1;
  assign f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_fa5_y4 = f_s_dadda_pg_rca32_fa5_y4;
  assign f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_fa4_y4 = f_s_dadda_pg_rca32_fa4_y4;
  assign f_s_dadda_pg_rca32_fa6_y0 = f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_ha3_y1 ^ f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_fa5_y4;
  assign f_s_dadda_pg_rca32_fa6_y1 = f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_ha3_y1 & f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_fa5_y4;
  assign f_s_dadda_pg_rca32_fa6_y2 = f_s_dadda_pg_rca32_fa6_y0 ^ f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_fa4_y4;
  assign f_s_dadda_pg_rca32_fa6_y3 = f_s_dadda_pg_rca32_fa6_y0 & f_s_dadda_pg_rca32_fa6_f_s_dadda_pg_rca32_fa4_y4;
  assign f_s_dadda_pg_rca32_fa6_y4 = f_s_dadda_pg_rca32_fa6_y1 | f_s_dadda_pg_rca32_fa6_y3;
  assign f_s_dadda_pg_rca32_nand_31_1_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_nand_31_1_y0 = ~(f_s_dadda_pg_rca32_nand_31_1_a_31 & f_s_dadda_pg_rca32_nand_31_1_b_1);
  assign f_s_dadda_pg_rca32_fa7_f_s_dadda_pg_rca32_fa3_y4 = f_s_dadda_pg_rca32_fa3_y4;
  assign f_s_dadda_pg_rca32_fa7_constant_wire_1 = constant_wire_1;
  assign f_s_dadda_pg_rca32_fa7_f_s_dadda_pg_rca32_nand_31_1_y0 = f_s_dadda_pg_rca32_nand_31_1_y0;
  assign f_s_dadda_pg_rca32_fa7_y0 = f_s_dadda_pg_rca32_fa7_f_s_dadda_pg_rca32_fa3_y4 ^ f_s_dadda_pg_rca32_fa7_constant_wire_1;
  assign f_s_dadda_pg_rca32_fa7_y1 = f_s_dadda_pg_rca32_fa7_f_s_dadda_pg_rca32_fa3_y4 & f_s_dadda_pg_rca32_fa7_constant_wire_1;
  assign f_s_dadda_pg_rca32_fa7_y2 = f_s_dadda_pg_rca32_fa7_y0 ^ f_s_dadda_pg_rca32_fa7_f_s_dadda_pg_rca32_nand_31_1_y0;
  assign f_s_dadda_pg_rca32_fa7_y3 = f_s_dadda_pg_rca32_fa7_y0 & f_s_dadda_pg_rca32_fa7_f_s_dadda_pg_rca32_nand_31_1_y0;
  assign f_s_dadda_pg_rca32_fa7_y4 = f_s_dadda_pg_rca32_fa7_y1 | f_s_dadda_pg_rca32_fa7_y3;
  assign f_s_dadda_pg_rca32_and_30_2_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_30_2_y0 = f_s_dadda_pg_rca32_and_30_2_a_30 & f_s_dadda_pg_rca32_and_30_2_b_2;
  assign f_s_dadda_pg_rca32_and_29_3_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_29_3_y0 = f_s_dadda_pg_rca32_and_29_3_a_29 & f_s_dadda_pg_rca32_and_29_3_b_3;
  assign f_s_dadda_pg_rca32_and_28_4_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_28_4_y0 = f_s_dadda_pg_rca32_and_28_4_a_28 & f_s_dadda_pg_rca32_and_28_4_b_4;
  assign f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_30_2_y0 = f_s_dadda_pg_rca32_and_30_2_y0;
  assign f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_29_3_y0 = f_s_dadda_pg_rca32_and_29_3_y0;
  assign f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_28_4_y0 = f_s_dadda_pg_rca32_and_28_4_y0;
  assign f_s_dadda_pg_rca32_fa8_y0 = f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_30_2_y0 ^ f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_29_3_y0;
  assign f_s_dadda_pg_rca32_fa8_y1 = f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_30_2_y0 & f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_29_3_y0;
  assign f_s_dadda_pg_rca32_fa8_y2 = f_s_dadda_pg_rca32_fa8_y0 ^ f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_28_4_y0;
  assign f_s_dadda_pg_rca32_fa8_y3 = f_s_dadda_pg_rca32_fa8_y0 & f_s_dadda_pg_rca32_fa8_f_s_dadda_pg_rca32_and_28_4_y0;
  assign f_s_dadda_pg_rca32_fa8_y4 = f_s_dadda_pg_rca32_fa8_y1 | f_s_dadda_pg_rca32_fa8_y3;
  assign f_s_dadda_pg_rca32_and_27_5_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_27_5_y0 = f_s_dadda_pg_rca32_and_27_5_a_27 & f_s_dadda_pg_rca32_and_27_5_b_5;
  assign f_s_dadda_pg_rca32_and_26_6_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_26_6_y0 = f_s_dadda_pg_rca32_and_26_6_a_26 & f_s_dadda_pg_rca32_and_26_6_b_6;
  assign f_s_dadda_pg_rca32_and_25_7_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_25_7_y0 = f_s_dadda_pg_rca32_and_25_7_a_25 & f_s_dadda_pg_rca32_and_25_7_b_7;
  assign f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_27_5_y0 = f_s_dadda_pg_rca32_and_27_5_y0;
  assign f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_26_6_y0 = f_s_dadda_pg_rca32_and_26_6_y0;
  assign f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_25_7_y0 = f_s_dadda_pg_rca32_and_25_7_y0;
  assign f_s_dadda_pg_rca32_fa9_y0 = f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_27_5_y0 ^ f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_26_6_y0;
  assign f_s_dadda_pg_rca32_fa9_y1 = f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_27_5_y0 & f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_26_6_y0;
  assign f_s_dadda_pg_rca32_fa9_y2 = f_s_dadda_pg_rca32_fa9_y0 ^ f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_25_7_y0;
  assign f_s_dadda_pg_rca32_fa9_y3 = f_s_dadda_pg_rca32_fa9_y0 & f_s_dadda_pg_rca32_fa9_f_s_dadda_pg_rca32_and_25_7_y0;
  assign f_s_dadda_pg_rca32_fa9_y4 = f_s_dadda_pg_rca32_fa9_y1 | f_s_dadda_pg_rca32_fa9_y3;
  assign f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa9_y4 = f_s_dadda_pg_rca32_fa9_y4;
  assign f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa8_y4 = f_s_dadda_pg_rca32_fa8_y4;
  assign f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa7_y4 = f_s_dadda_pg_rca32_fa7_y4;
  assign f_s_dadda_pg_rca32_fa10_y0 = f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa9_y4 ^ f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa8_y4;
  assign f_s_dadda_pg_rca32_fa10_y1 = f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa9_y4 & f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa8_y4;
  assign f_s_dadda_pg_rca32_fa10_y2 = f_s_dadda_pg_rca32_fa10_y0 ^ f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa7_y4;
  assign f_s_dadda_pg_rca32_fa10_y3 = f_s_dadda_pg_rca32_fa10_y0 & f_s_dadda_pg_rca32_fa10_f_s_dadda_pg_rca32_fa7_y4;
  assign f_s_dadda_pg_rca32_fa10_y4 = f_s_dadda_pg_rca32_fa10_y1 | f_s_dadda_pg_rca32_fa10_y3;
  assign f_s_dadda_pg_rca32_nand_31_2_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_nand_31_2_y0 = ~(f_s_dadda_pg_rca32_nand_31_2_a_31 & f_s_dadda_pg_rca32_nand_31_2_b_2);
  assign f_s_dadda_pg_rca32_and_30_3_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_30_3_y0 = f_s_dadda_pg_rca32_and_30_3_a_30 & f_s_dadda_pg_rca32_and_30_3_b_3;
  assign f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_fa6_y4 = f_s_dadda_pg_rca32_fa6_y4;
  assign f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_nand_31_2_y0 = f_s_dadda_pg_rca32_nand_31_2_y0;
  assign f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_and_30_3_y0 = f_s_dadda_pg_rca32_and_30_3_y0;
  assign f_s_dadda_pg_rca32_fa11_y0 = f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_fa6_y4 ^ f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_nand_31_2_y0;
  assign f_s_dadda_pg_rca32_fa11_y1 = f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_fa6_y4 & f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_nand_31_2_y0;
  assign f_s_dadda_pg_rca32_fa11_y2 = f_s_dadda_pg_rca32_fa11_y0 ^ f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_and_30_3_y0;
  assign f_s_dadda_pg_rca32_fa11_y3 = f_s_dadda_pg_rca32_fa11_y0 & f_s_dadda_pg_rca32_fa11_f_s_dadda_pg_rca32_and_30_3_y0;
  assign f_s_dadda_pg_rca32_fa11_y4 = f_s_dadda_pg_rca32_fa11_y1 | f_s_dadda_pg_rca32_fa11_y3;
  assign f_s_dadda_pg_rca32_and_29_4_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_29_4_y0 = f_s_dadda_pg_rca32_and_29_4_a_29 & f_s_dadda_pg_rca32_and_29_4_b_4;
  assign f_s_dadda_pg_rca32_and_28_5_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_28_5_y0 = f_s_dadda_pg_rca32_and_28_5_a_28 & f_s_dadda_pg_rca32_and_28_5_b_5;
  assign f_s_dadda_pg_rca32_and_27_6_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_27_6_y0 = f_s_dadda_pg_rca32_and_27_6_a_27 & f_s_dadda_pg_rca32_and_27_6_b_6;
  assign f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_29_4_y0 = f_s_dadda_pg_rca32_and_29_4_y0;
  assign f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_28_5_y0 = f_s_dadda_pg_rca32_and_28_5_y0;
  assign f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_27_6_y0 = f_s_dadda_pg_rca32_and_27_6_y0;
  assign f_s_dadda_pg_rca32_fa12_y0 = f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_29_4_y0 ^ f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_28_5_y0;
  assign f_s_dadda_pg_rca32_fa12_y1 = f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_29_4_y0 & f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_28_5_y0;
  assign f_s_dadda_pg_rca32_fa12_y2 = f_s_dadda_pg_rca32_fa12_y0 ^ f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_27_6_y0;
  assign f_s_dadda_pg_rca32_fa12_y3 = f_s_dadda_pg_rca32_fa12_y0 & f_s_dadda_pg_rca32_fa12_f_s_dadda_pg_rca32_and_27_6_y0;
  assign f_s_dadda_pg_rca32_fa12_y4 = f_s_dadda_pg_rca32_fa12_y1 | f_s_dadda_pg_rca32_fa12_y3;
  assign f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa12_y4 = f_s_dadda_pg_rca32_fa12_y4;
  assign f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa11_y4 = f_s_dadda_pg_rca32_fa11_y4;
  assign f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa10_y4 = f_s_dadda_pg_rca32_fa10_y4;
  assign f_s_dadda_pg_rca32_fa13_y0 = f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa12_y4 ^ f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa11_y4;
  assign f_s_dadda_pg_rca32_fa13_y1 = f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa12_y4 & f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa11_y4;
  assign f_s_dadda_pg_rca32_fa13_y2 = f_s_dadda_pg_rca32_fa13_y0 ^ f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa10_y4;
  assign f_s_dadda_pg_rca32_fa13_y3 = f_s_dadda_pg_rca32_fa13_y0 & f_s_dadda_pg_rca32_fa13_f_s_dadda_pg_rca32_fa10_y4;
  assign f_s_dadda_pg_rca32_fa13_y4 = f_s_dadda_pg_rca32_fa13_y1 | f_s_dadda_pg_rca32_fa13_y3;
  assign f_s_dadda_pg_rca32_nand_31_3_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_nand_31_3_y0 = ~(f_s_dadda_pg_rca32_nand_31_3_a_31 & f_s_dadda_pg_rca32_nand_31_3_b_3);
  assign f_s_dadda_pg_rca32_and_30_4_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_30_4_y0 = f_s_dadda_pg_rca32_and_30_4_a_30 & f_s_dadda_pg_rca32_and_30_4_b_4;
  assign f_s_dadda_pg_rca32_and_29_5_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_29_5_y0 = f_s_dadda_pg_rca32_and_29_5_a_29 & f_s_dadda_pg_rca32_and_29_5_b_5;
  assign f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_nand_31_3_y0 = f_s_dadda_pg_rca32_nand_31_3_y0;
  assign f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_and_30_4_y0 = f_s_dadda_pg_rca32_and_30_4_y0;
  assign f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_and_29_5_y0 = f_s_dadda_pg_rca32_and_29_5_y0;
  assign f_s_dadda_pg_rca32_fa14_y0 = f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_nand_31_3_y0 ^ f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_and_30_4_y0;
  assign f_s_dadda_pg_rca32_fa14_y1 = f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_nand_31_3_y0 & f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_and_30_4_y0;
  assign f_s_dadda_pg_rca32_fa14_y2 = f_s_dadda_pg_rca32_fa14_y0 ^ f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_and_29_5_y0;
  assign f_s_dadda_pg_rca32_fa14_y3 = f_s_dadda_pg_rca32_fa14_y0 & f_s_dadda_pg_rca32_fa14_f_s_dadda_pg_rca32_and_29_5_y0;
  assign f_s_dadda_pg_rca32_fa14_y4 = f_s_dadda_pg_rca32_fa14_y1 | f_s_dadda_pg_rca32_fa14_y3;
  assign f_s_dadda_pg_rca32_nand_31_4_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_nand_31_4_y0 = ~(f_s_dadda_pg_rca32_nand_31_4_a_31 & f_s_dadda_pg_rca32_nand_31_4_b_4);
  assign f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_fa14_y4 = f_s_dadda_pg_rca32_fa14_y4;
  assign f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_fa13_y4 = f_s_dadda_pg_rca32_fa13_y4;
  assign f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_nand_31_4_y0 = f_s_dadda_pg_rca32_nand_31_4_y0;
  assign f_s_dadda_pg_rca32_fa15_y0 = f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_fa14_y4 ^ f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_fa13_y4;
  assign f_s_dadda_pg_rca32_fa15_y1 = f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_fa14_y4 & f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_fa13_y4;
  assign f_s_dadda_pg_rca32_fa15_y2 = f_s_dadda_pg_rca32_fa15_y0 ^ f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_nand_31_4_y0;
  assign f_s_dadda_pg_rca32_fa15_y3 = f_s_dadda_pg_rca32_fa15_y0 & f_s_dadda_pg_rca32_fa15_f_s_dadda_pg_rca32_nand_31_4_y0;
  assign f_s_dadda_pg_rca32_fa15_y4 = f_s_dadda_pg_rca32_fa15_y1 | f_s_dadda_pg_rca32_fa15_y3;
  assign f_s_dadda_pg_rca32_and_6_0_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_6_0_y0 = f_s_dadda_pg_rca32_and_6_0_a_6 & f_s_dadda_pg_rca32_and_6_0_b_0;
  assign f_s_dadda_pg_rca32_and_5_1_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_5_1_y0 = f_s_dadda_pg_rca32_and_5_1_a_5 & f_s_dadda_pg_rca32_and_5_1_b_1;
  assign f_s_dadda_pg_rca32_ha4_f_s_dadda_pg_rca32_and_6_0_y0 = f_s_dadda_pg_rca32_and_6_0_y0;
  assign f_s_dadda_pg_rca32_ha4_f_s_dadda_pg_rca32_and_5_1_y0 = f_s_dadda_pg_rca32_and_5_1_y0;
  assign f_s_dadda_pg_rca32_ha4_y0 = f_s_dadda_pg_rca32_ha4_f_s_dadda_pg_rca32_and_6_0_y0 ^ f_s_dadda_pg_rca32_ha4_f_s_dadda_pg_rca32_and_5_1_y0;
  assign f_s_dadda_pg_rca32_ha4_y1 = f_s_dadda_pg_rca32_ha4_f_s_dadda_pg_rca32_and_6_0_y0 & f_s_dadda_pg_rca32_ha4_f_s_dadda_pg_rca32_and_5_1_y0;
  assign f_s_dadda_pg_rca32_and_7_0_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_7_0_y0 = f_s_dadda_pg_rca32_and_7_0_a_7 & f_s_dadda_pg_rca32_and_7_0_b_0;
  assign f_s_dadda_pg_rca32_and_6_1_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_6_1_y0 = f_s_dadda_pg_rca32_and_6_1_a_6 & f_s_dadda_pg_rca32_and_6_1_b_1;
  assign f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_ha4_y1 = f_s_dadda_pg_rca32_ha4_y1;
  assign f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_and_7_0_y0 = f_s_dadda_pg_rca32_and_7_0_y0;
  assign f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_and_6_1_y0 = f_s_dadda_pg_rca32_and_6_1_y0;
  assign f_s_dadda_pg_rca32_fa16_y0 = f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_ha4_y1 ^ f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_and_7_0_y0;
  assign f_s_dadda_pg_rca32_fa16_y1 = f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_ha4_y1 & f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_and_7_0_y0;
  assign f_s_dadda_pg_rca32_fa16_y2 = f_s_dadda_pg_rca32_fa16_y0 ^ f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_and_6_1_y0;
  assign f_s_dadda_pg_rca32_fa16_y3 = f_s_dadda_pg_rca32_fa16_y0 & f_s_dadda_pg_rca32_fa16_f_s_dadda_pg_rca32_and_6_1_y0;
  assign f_s_dadda_pg_rca32_fa16_y4 = f_s_dadda_pg_rca32_fa16_y1 | f_s_dadda_pg_rca32_fa16_y3;
  assign f_s_dadda_pg_rca32_and_5_2_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_5_2_y0 = f_s_dadda_pg_rca32_and_5_2_a_5 & f_s_dadda_pg_rca32_and_5_2_b_2;
  assign f_s_dadda_pg_rca32_and_4_3_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_4_3_y0 = f_s_dadda_pg_rca32_and_4_3_a_4 & f_s_dadda_pg_rca32_and_4_3_b_3;
  assign f_s_dadda_pg_rca32_ha5_f_s_dadda_pg_rca32_and_5_2_y0 = f_s_dadda_pg_rca32_and_5_2_y0;
  assign f_s_dadda_pg_rca32_ha5_f_s_dadda_pg_rca32_and_4_3_y0 = f_s_dadda_pg_rca32_and_4_3_y0;
  assign f_s_dadda_pg_rca32_ha5_y0 = f_s_dadda_pg_rca32_ha5_f_s_dadda_pg_rca32_and_5_2_y0 ^ f_s_dadda_pg_rca32_ha5_f_s_dadda_pg_rca32_and_4_3_y0;
  assign f_s_dadda_pg_rca32_ha5_y1 = f_s_dadda_pg_rca32_ha5_f_s_dadda_pg_rca32_and_5_2_y0 & f_s_dadda_pg_rca32_ha5_f_s_dadda_pg_rca32_and_4_3_y0;
  assign f_s_dadda_pg_rca32_and_8_0_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_8_0_y0 = f_s_dadda_pg_rca32_and_8_0_a_8 & f_s_dadda_pg_rca32_and_8_0_b_0;
  assign f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_ha5_y1 = f_s_dadda_pg_rca32_ha5_y1;
  assign f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_fa16_y4 = f_s_dadda_pg_rca32_fa16_y4;
  assign f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_and_8_0_y0 = f_s_dadda_pg_rca32_and_8_0_y0;
  assign f_s_dadda_pg_rca32_fa17_y0 = f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_ha5_y1 ^ f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_fa16_y4;
  assign f_s_dadda_pg_rca32_fa17_y1 = f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_ha5_y1 & f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_fa16_y4;
  assign f_s_dadda_pg_rca32_fa17_y2 = f_s_dadda_pg_rca32_fa17_y0 ^ f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_and_8_0_y0;
  assign f_s_dadda_pg_rca32_fa17_y3 = f_s_dadda_pg_rca32_fa17_y0 & f_s_dadda_pg_rca32_fa17_f_s_dadda_pg_rca32_and_8_0_y0;
  assign f_s_dadda_pg_rca32_fa17_y4 = f_s_dadda_pg_rca32_fa17_y1 | f_s_dadda_pg_rca32_fa17_y3;
  assign f_s_dadda_pg_rca32_and_7_1_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_7_1_y0 = f_s_dadda_pg_rca32_and_7_1_a_7 & f_s_dadda_pg_rca32_and_7_1_b_1;
  assign f_s_dadda_pg_rca32_and_6_2_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_6_2_y0 = f_s_dadda_pg_rca32_and_6_2_a_6 & f_s_dadda_pg_rca32_and_6_2_b_2;
  assign f_s_dadda_pg_rca32_and_5_3_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_5_3_y0 = f_s_dadda_pg_rca32_and_5_3_a_5 & f_s_dadda_pg_rca32_and_5_3_b_3;
  assign f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_7_1_y0 = f_s_dadda_pg_rca32_and_7_1_y0;
  assign f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_6_2_y0 = f_s_dadda_pg_rca32_and_6_2_y0;
  assign f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_5_3_y0 = f_s_dadda_pg_rca32_and_5_3_y0;
  assign f_s_dadda_pg_rca32_fa18_y0 = f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_7_1_y0 ^ f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_6_2_y0;
  assign f_s_dadda_pg_rca32_fa18_y1 = f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_7_1_y0 & f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_6_2_y0;
  assign f_s_dadda_pg_rca32_fa18_y2 = f_s_dadda_pg_rca32_fa18_y0 ^ f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_5_3_y0;
  assign f_s_dadda_pg_rca32_fa18_y3 = f_s_dadda_pg_rca32_fa18_y0 & f_s_dadda_pg_rca32_fa18_f_s_dadda_pg_rca32_and_5_3_y0;
  assign f_s_dadda_pg_rca32_fa18_y4 = f_s_dadda_pg_rca32_fa18_y1 | f_s_dadda_pg_rca32_fa18_y3;
  assign f_s_dadda_pg_rca32_and_4_4_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_4_4_y0 = f_s_dadda_pg_rca32_and_4_4_a_4 & f_s_dadda_pg_rca32_and_4_4_b_4;
  assign f_s_dadda_pg_rca32_and_3_5_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_3_5_y0 = f_s_dadda_pg_rca32_and_3_5_a_3 & f_s_dadda_pg_rca32_and_3_5_b_5;
  assign f_s_dadda_pg_rca32_ha6_f_s_dadda_pg_rca32_and_4_4_y0 = f_s_dadda_pg_rca32_and_4_4_y0;
  assign f_s_dadda_pg_rca32_ha6_f_s_dadda_pg_rca32_and_3_5_y0 = f_s_dadda_pg_rca32_and_3_5_y0;
  assign f_s_dadda_pg_rca32_ha6_y0 = f_s_dadda_pg_rca32_ha6_f_s_dadda_pg_rca32_and_4_4_y0 ^ f_s_dadda_pg_rca32_ha6_f_s_dadda_pg_rca32_and_3_5_y0;
  assign f_s_dadda_pg_rca32_ha6_y1 = f_s_dadda_pg_rca32_ha6_f_s_dadda_pg_rca32_and_4_4_y0 & f_s_dadda_pg_rca32_ha6_f_s_dadda_pg_rca32_and_3_5_y0;
  assign f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_ha6_y1 = f_s_dadda_pg_rca32_ha6_y1;
  assign f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_fa18_y4 = f_s_dadda_pg_rca32_fa18_y4;
  assign f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_fa17_y4 = f_s_dadda_pg_rca32_fa17_y4;
  assign f_s_dadda_pg_rca32_fa19_y0 = f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_ha6_y1 ^ f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_fa18_y4;
  assign f_s_dadda_pg_rca32_fa19_y1 = f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_ha6_y1 & f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_fa18_y4;
  assign f_s_dadda_pg_rca32_fa19_y2 = f_s_dadda_pg_rca32_fa19_y0 ^ f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_fa17_y4;
  assign f_s_dadda_pg_rca32_fa19_y3 = f_s_dadda_pg_rca32_fa19_y0 & f_s_dadda_pg_rca32_fa19_f_s_dadda_pg_rca32_fa17_y4;
  assign f_s_dadda_pg_rca32_fa19_y4 = f_s_dadda_pg_rca32_fa19_y1 | f_s_dadda_pg_rca32_fa19_y3;
  assign f_s_dadda_pg_rca32_and_9_0_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_9_0_y0 = f_s_dadda_pg_rca32_and_9_0_a_9 & f_s_dadda_pg_rca32_and_9_0_b_0;
  assign f_s_dadda_pg_rca32_and_8_1_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_8_1_y0 = f_s_dadda_pg_rca32_and_8_1_a_8 & f_s_dadda_pg_rca32_and_8_1_b_1;
  assign f_s_dadda_pg_rca32_and_7_2_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_7_2_y0 = f_s_dadda_pg_rca32_and_7_2_a_7 & f_s_dadda_pg_rca32_and_7_2_b_2;
  assign f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_9_0_y0 = f_s_dadda_pg_rca32_and_9_0_y0;
  assign f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_8_1_y0 = f_s_dadda_pg_rca32_and_8_1_y0;
  assign f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_7_2_y0 = f_s_dadda_pg_rca32_and_7_2_y0;
  assign f_s_dadda_pg_rca32_fa20_y0 = f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_9_0_y0 ^ f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_8_1_y0;
  assign f_s_dadda_pg_rca32_fa20_y1 = f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_9_0_y0 & f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_8_1_y0;
  assign f_s_dadda_pg_rca32_fa20_y2 = f_s_dadda_pg_rca32_fa20_y0 ^ f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_7_2_y0;
  assign f_s_dadda_pg_rca32_fa20_y3 = f_s_dadda_pg_rca32_fa20_y0 & f_s_dadda_pg_rca32_fa20_f_s_dadda_pg_rca32_and_7_2_y0;
  assign f_s_dadda_pg_rca32_fa20_y4 = f_s_dadda_pg_rca32_fa20_y1 | f_s_dadda_pg_rca32_fa20_y3;
  assign f_s_dadda_pg_rca32_and_6_3_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_6_3_y0 = f_s_dadda_pg_rca32_and_6_3_a_6 & f_s_dadda_pg_rca32_and_6_3_b_3;
  assign f_s_dadda_pg_rca32_and_5_4_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_5_4_y0 = f_s_dadda_pg_rca32_and_5_4_a_5 & f_s_dadda_pg_rca32_and_5_4_b_4;
  assign f_s_dadda_pg_rca32_and_4_5_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_4_5_y0 = f_s_dadda_pg_rca32_and_4_5_a_4 & f_s_dadda_pg_rca32_and_4_5_b_5;
  assign f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_6_3_y0 = f_s_dadda_pg_rca32_and_6_3_y0;
  assign f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_5_4_y0 = f_s_dadda_pg_rca32_and_5_4_y0;
  assign f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_4_5_y0 = f_s_dadda_pg_rca32_and_4_5_y0;
  assign f_s_dadda_pg_rca32_fa21_y0 = f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_6_3_y0 ^ f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_5_4_y0;
  assign f_s_dadda_pg_rca32_fa21_y1 = f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_6_3_y0 & f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_5_4_y0;
  assign f_s_dadda_pg_rca32_fa21_y2 = f_s_dadda_pg_rca32_fa21_y0 ^ f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_4_5_y0;
  assign f_s_dadda_pg_rca32_fa21_y3 = f_s_dadda_pg_rca32_fa21_y0 & f_s_dadda_pg_rca32_fa21_f_s_dadda_pg_rca32_and_4_5_y0;
  assign f_s_dadda_pg_rca32_fa21_y4 = f_s_dadda_pg_rca32_fa21_y1 | f_s_dadda_pg_rca32_fa21_y3;
  assign f_s_dadda_pg_rca32_and_3_6_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_3_6_y0 = f_s_dadda_pg_rca32_and_3_6_a_3 & f_s_dadda_pg_rca32_and_3_6_b_6;
  assign f_s_dadda_pg_rca32_and_2_7_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_2_7_y0 = f_s_dadda_pg_rca32_and_2_7_a_2 & f_s_dadda_pg_rca32_and_2_7_b_7;
  assign f_s_dadda_pg_rca32_ha7_f_s_dadda_pg_rca32_and_3_6_y0 = f_s_dadda_pg_rca32_and_3_6_y0;
  assign f_s_dadda_pg_rca32_ha7_f_s_dadda_pg_rca32_and_2_7_y0 = f_s_dadda_pg_rca32_and_2_7_y0;
  assign f_s_dadda_pg_rca32_ha7_y0 = f_s_dadda_pg_rca32_ha7_f_s_dadda_pg_rca32_and_3_6_y0 ^ f_s_dadda_pg_rca32_ha7_f_s_dadda_pg_rca32_and_2_7_y0;
  assign f_s_dadda_pg_rca32_ha7_y1 = f_s_dadda_pg_rca32_ha7_f_s_dadda_pg_rca32_and_3_6_y0 & f_s_dadda_pg_rca32_ha7_f_s_dadda_pg_rca32_and_2_7_y0;
  assign f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_ha7_y1 = f_s_dadda_pg_rca32_ha7_y1;
  assign f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_fa21_y4 = f_s_dadda_pg_rca32_fa21_y4;
  assign f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_fa20_y4 = f_s_dadda_pg_rca32_fa20_y4;
  assign f_s_dadda_pg_rca32_fa22_y0 = f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_ha7_y1 ^ f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_fa21_y4;
  assign f_s_dadda_pg_rca32_fa22_y1 = f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_ha7_y1 & f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_fa21_y4;
  assign f_s_dadda_pg_rca32_fa22_y2 = f_s_dadda_pg_rca32_fa22_y0 ^ f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_fa20_y4;
  assign f_s_dadda_pg_rca32_fa22_y3 = f_s_dadda_pg_rca32_fa22_y0 & f_s_dadda_pg_rca32_fa22_f_s_dadda_pg_rca32_fa20_y4;
  assign f_s_dadda_pg_rca32_fa22_y4 = f_s_dadda_pg_rca32_fa22_y1 | f_s_dadda_pg_rca32_fa22_y3;
  assign f_s_dadda_pg_rca32_and_10_0_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_10_0_y0 = f_s_dadda_pg_rca32_and_10_0_a_10 & f_s_dadda_pg_rca32_and_10_0_b_0;
  assign f_s_dadda_pg_rca32_and_9_1_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_9_1_y0 = f_s_dadda_pg_rca32_and_9_1_a_9 & f_s_dadda_pg_rca32_and_9_1_b_1;
  assign f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_fa19_y4 = f_s_dadda_pg_rca32_fa19_y4;
  assign f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_and_10_0_y0 = f_s_dadda_pg_rca32_and_10_0_y0;
  assign f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_and_9_1_y0 = f_s_dadda_pg_rca32_and_9_1_y0;
  assign f_s_dadda_pg_rca32_fa23_y0 = f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_fa19_y4 ^ f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_and_10_0_y0;
  assign f_s_dadda_pg_rca32_fa23_y1 = f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_fa19_y4 & f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_and_10_0_y0;
  assign f_s_dadda_pg_rca32_fa23_y2 = f_s_dadda_pg_rca32_fa23_y0 ^ f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_and_9_1_y0;
  assign f_s_dadda_pg_rca32_fa23_y3 = f_s_dadda_pg_rca32_fa23_y0 & f_s_dadda_pg_rca32_fa23_f_s_dadda_pg_rca32_and_9_1_y0;
  assign f_s_dadda_pg_rca32_fa23_y4 = f_s_dadda_pg_rca32_fa23_y1 | f_s_dadda_pg_rca32_fa23_y3;
  assign f_s_dadda_pg_rca32_and_8_2_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_8_2_y0 = f_s_dadda_pg_rca32_and_8_2_a_8 & f_s_dadda_pg_rca32_and_8_2_b_2;
  assign f_s_dadda_pg_rca32_and_7_3_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_7_3_y0 = f_s_dadda_pg_rca32_and_7_3_a_7 & f_s_dadda_pg_rca32_and_7_3_b_3;
  assign f_s_dadda_pg_rca32_and_6_4_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_6_4_y0 = f_s_dadda_pg_rca32_and_6_4_a_6 & f_s_dadda_pg_rca32_and_6_4_b_4;
  assign f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_8_2_y0 = f_s_dadda_pg_rca32_and_8_2_y0;
  assign f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_7_3_y0 = f_s_dadda_pg_rca32_and_7_3_y0;
  assign f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_6_4_y0 = f_s_dadda_pg_rca32_and_6_4_y0;
  assign f_s_dadda_pg_rca32_fa24_y0 = f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_8_2_y0 ^ f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_7_3_y0;
  assign f_s_dadda_pg_rca32_fa24_y1 = f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_8_2_y0 & f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_7_3_y0;
  assign f_s_dadda_pg_rca32_fa24_y2 = f_s_dadda_pg_rca32_fa24_y0 ^ f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_6_4_y0;
  assign f_s_dadda_pg_rca32_fa24_y3 = f_s_dadda_pg_rca32_fa24_y0 & f_s_dadda_pg_rca32_fa24_f_s_dadda_pg_rca32_and_6_4_y0;
  assign f_s_dadda_pg_rca32_fa24_y4 = f_s_dadda_pg_rca32_fa24_y1 | f_s_dadda_pg_rca32_fa24_y3;
  assign f_s_dadda_pg_rca32_and_5_5_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_5_5_y0 = f_s_dadda_pg_rca32_and_5_5_a_5 & f_s_dadda_pg_rca32_and_5_5_b_5;
  assign f_s_dadda_pg_rca32_and_4_6_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_4_6_y0 = f_s_dadda_pg_rca32_and_4_6_a_4 & f_s_dadda_pg_rca32_and_4_6_b_6;
  assign f_s_dadda_pg_rca32_and_3_7_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_3_7_y0 = f_s_dadda_pg_rca32_and_3_7_a_3 & f_s_dadda_pg_rca32_and_3_7_b_7;
  assign f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_5_5_y0 = f_s_dadda_pg_rca32_and_5_5_y0;
  assign f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_4_6_y0 = f_s_dadda_pg_rca32_and_4_6_y0;
  assign f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_3_7_y0 = f_s_dadda_pg_rca32_and_3_7_y0;
  assign f_s_dadda_pg_rca32_fa25_y0 = f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_5_5_y0 ^ f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_4_6_y0;
  assign f_s_dadda_pg_rca32_fa25_y1 = f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_5_5_y0 & f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_4_6_y0;
  assign f_s_dadda_pg_rca32_fa25_y2 = f_s_dadda_pg_rca32_fa25_y0 ^ f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_3_7_y0;
  assign f_s_dadda_pg_rca32_fa25_y3 = f_s_dadda_pg_rca32_fa25_y0 & f_s_dadda_pg_rca32_fa25_f_s_dadda_pg_rca32_and_3_7_y0;
  assign f_s_dadda_pg_rca32_fa25_y4 = f_s_dadda_pg_rca32_fa25_y1 | f_s_dadda_pg_rca32_fa25_y3;
  assign f_s_dadda_pg_rca32_and_2_8_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_2_8_y0 = f_s_dadda_pg_rca32_and_2_8_a_2 & f_s_dadda_pg_rca32_and_2_8_b_8;
  assign f_s_dadda_pg_rca32_and_1_9_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_1_9_y0 = f_s_dadda_pg_rca32_and_1_9_a_1 & f_s_dadda_pg_rca32_and_1_9_b_9;
  assign f_s_dadda_pg_rca32_ha8_f_s_dadda_pg_rca32_and_2_8_y0 = f_s_dadda_pg_rca32_and_2_8_y0;
  assign f_s_dadda_pg_rca32_ha8_f_s_dadda_pg_rca32_and_1_9_y0 = f_s_dadda_pg_rca32_and_1_9_y0;
  assign f_s_dadda_pg_rca32_ha8_y0 = f_s_dadda_pg_rca32_ha8_f_s_dadda_pg_rca32_and_2_8_y0 ^ f_s_dadda_pg_rca32_ha8_f_s_dadda_pg_rca32_and_1_9_y0;
  assign f_s_dadda_pg_rca32_ha8_y1 = f_s_dadda_pg_rca32_ha8_f_s_dadda_pg_rca32_and_2_8_y0 & f_s_dadda_pg_rca32_ha8_f_s_dadda_pg_rca32_and_1_9_y0;
  assign f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_ha8_y1 = f_s_dadda_pg_rca32_ha8_y1;
  assign f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_fa25_y4 = f_s_dadda_pg_rca32_fa25_y4;
  assign f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_fa24_y4 = f_s_dadda_pg_rca32_fa24_y4;
  assign f_s_dadda_pg_rca32_fa26_y0 = f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_ha8_y1 ^ f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_fa25_y4;
  assign f_s_dadda_pg_rca32_fa26_y1 = f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_ha8_y1 & f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_fa25_y4;
  assign f_s_dadda_pg_rca32_fa26_y2 = f_s_dadda_pg_rca32_fa26_y0 ^ f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_fa24_y4;
  assign f_s_dadda_pg_rca32_fa26_y3 = f_s_dadda_pg_rca32_fa26_y0 & f_s_dadda_pg_rca32_fa26_f_s_dadda_pg_rca32_fa24_y4;
  assign f_s_dadda_pg_rca32_fa26_y4 = f_s_dadda_pg_rca32_fa26_y1 | f_s_dadda_pg_rca32_fa26_y3;
  assign f_s_dadda_pg_rca32_and_11_0_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_11_0_y0 = f_s_dadda_pg_rca32_and_11_0_a_11 & f_s_dadda_pg_rca32_and_11_0_b_0;
  assign f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_fa23_y4 = f_s_dadda_pg_rca32_fa23_y4;
  assign f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_fa22_y4 = f_s_dadda_pg_rca32_fa22_y4;
  assign f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_and_11_0_y0 = f_s_dadda_pg_rca32_and_11_0_y0;
  assign f_s_dadda_pg_rca32_fa27_y0 = f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_fa23_y4 ^ f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_fa22_y4;
  assign f_s_dadda_pg_rca32_fa27_y1 = f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_fa23_y4 & f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_fa22_y4;
  assign f_s_dadda_pg_rca32_fa27_y2 = f_s_dadda_pg_rca32_fa27_y0 ^ f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_and_11_0_y0;
  assign f_s_dadda_pg_rca32_fa27_y3 = f_s_dadda_pg_rca32_fa27_y0 & f_s_dadda_pg_rca32_fa27_f_s_dadda_pg_rca32_and_11_0_y0;
  assign f_s_dadda_pg_rca32_fa27_y4 = f_s_dadda_pg_rca32_fa27_y1 | f_s_dadda_pg_rca32_fa27_y3;
  assign f_s_dadda_pg_rca32_and_10_1_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_10_1_y0 = f_s_dadda_pg_rca32_and_10_1_a_10 & f_s_dadda_pg_rca32_and_10_1_b_1;
  assign f_s_dadda_pg_rca32_and_9_2_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_9_2_y0 = f_s_dadda_pg_rca32_and_9_2_a_9 & f_s_dadda_pg_rca32_and_9_2_b_2;
  assign f_s_dadda_pg_rca32_and_8_3_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_8_3_y0 = f_s_dadda_pg_rca32_and_8_3_a_8 & f_s_dadda_pg_rca32_and_8_3_b_3;
  assign f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_10_1_y0 = f_s_dadda_pg_rca32_and_10_1_y0;
  assign f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_9_2_y0 = f_s_dadda_pg_rca32_and_9_2_y0;
  assign f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_8_3_y0 = f_s_dadda_pg_rca32_and_8_3_y0;
  assign f_s_dadda_pg_rca32_fa28_y0 = f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_10_1_y0 ^ f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_9_2_y0;
  assign f_s_dadda_pg_rca32_fa28_y1 = f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_10_1_y0 & f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_9_2_y0;
  assign f_s_dadda_pg_rca32_fa28_y2 = f_s_dadda_pg_rca32_fa28_y0 ^ f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_8_3_y0;
  assign f_s_dadda_pg_rca32_fa28_y3 = f_s_dadda_pg_rca32_fa28_y0 & f_s_dadda_pg_rca32_fa28_f_s_dadda_pg_rca32_and_8_3_y0;
  assign f_s_dadda_pg_rca32_fa28_y4 = f_s_dadda_pg_rca32_fa28_y1 | f_s_dadda_pg_rca32_fa28_y3;
  assign f_s_dadda_pg_rca32_and_7_4_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_7_4_y0 = f_s_dadda_pg_rca32_and_7_4_a_7 & f_s_dadda_pg_rca32_and_7_4_b_4;
  assign f_s_dadda_pg_rca32_and_6_5_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_6_5_y0 = f_s_dadda_pg_rca32_and_6_5_a_6 & f_s_dadda_pg_rca32_and_6_5_b_5;
  assign f_s_dadda_pg_rca32_and_5_6_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_5_6_y0 = f_s_dadda_pg_rca32_and_5_6_a_5 & f_s_dadda_pg_rca32_and_5_6_b_6;
  assign f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_7_4_y0 = f_s_dadda_pg_rca32_and_7_4_y0;
  assign f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_6_5_y0 = f_s_dadda_pg_rca32_and_6_5_y0;
  assign f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_5_6_y0 = f_s_dadda_pg_rca32_and_5_6_y0;
  assign f_s_dadda_pg_rca32_fa29_y0 = f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_7_4_y0 ^ f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_6_5_y0;
  assign f_s_dadda_pg_rca32_fa29_y1 = f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_7_4_y0 & f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_6_5_y0;
  assign f_s_dadda_pg_rca32_fa29_y2 = f_s_dadda_pg_rca32_fa29_y0 ^ f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_5_6_y0;
  assign f_s_dadda_pg_rca32_fa29_y3 = f_s_dadda_pg_rca32_fa29_y0 & f_s_dadda_pg_rca32_fa29_f_s_dadda_pg_rca32_and_5_6_y0;
  assign f_s_dadda_pg_rca32_fa29_y4 = f_s_dadda_pg_rca32_fa29_y1 | f_s_dadda_pg_rca32_fa29_y3;
  assign f_s_dadda_pg_rca32_and_4_7_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_4_7_y0 = f_s_dadda_pg_rca32_and_4_7_a_4 & f_s_dadda_pg_rca32_and_4_7_b_7;
  assign f_s_dadda_pg_rca32_and_3_8_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_3_8_y0 = f_s_dadda_pg_rca32_and_3_8_a_3 & f_s_dadda_pg_rca32_and_3_8_b_8;
  assign f_s_dadda_pg_rca32_and_2_9_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_2_9_y0 = f_s_dadda_pg_rca32_and_2_9_a_2 & f_s_dadda_pg_rca32_and_2_9_b_9;
  assign f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_4_7_y0 = f_s_dadda_pg_rca32_and_4_7_y0;
  assign f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_3_8_y0 = f_s_dadda_pg_rca32_and_3_8_y0;
  assign f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_2_9_y0 = f_s_dadda_pg_rca32_and_2_9_y0;
  assign f_s_dadda_pg_rca32_fa30_y0 = f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_4_7_y0 ^ f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_3_8_y0;
  assign f_s_dadda_pg_rca32_fa30_y1 = f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_4_7_y0 & f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_3_8_y0;
  assign f_s_dadda_pg_rca32_fa30_y2 = f_s_dadda_pg_rca32_fa30_y0 ^ f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_2_9_y0;
  assign f_s_dadda_pg_rca32_fa30_y3 = f_s_dadda_pg_rca32_fa30_y0 & f_s_dadda_pg_rca32_fa30_f_s_dadda_pg_rca32_and_2_9_y0;
  assign f_s_dadda_pg_rca32_fa30_y4 = f_s_dadda_pg_rca32_fa30_y1 | f_s_dadda_pg_rca32_fa30_y3;
  assign f_s_dadda_pg_rca32_and_1_10_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_1_10_y0 = f_s_dadda_pg_rca32_and_1_10_a_1 & f_s_dadda_pg_rca32_and_1_10_b_10;
  assign f_s_dadda_pg_rca32_and_0_11_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_0_11_y0 = f_s_dadda_pg_rca32_and_0_11_a_0 & f_s_dadda_pg_rca32_and_0_11_b_11;
  assign f_s_dadda_pg_rca32_ha9_f_s_dadda_pg_rca32_and_1_10_y0 = f_s_dadda_pg_rca32_and_1_10_y0;
  assign f_s_dadda_pg_rca32_ha9_f_s_dadda_pg_rca32_and_0_11_y0 = f_s_dadda_pg_rca32_and_0_11_y0;
  assign f_s_dadda_pg_rca32_ha9_y0 = f_s_dadda_pg_rca32_ha9_f_s_dadda_pg_rca32_and_1_10_y0 ^ f_s_dadda_pg_rca32_ha9_f_s_dadda_pg_rca32_and_0_11_y0;
  assign f_s_dadda_pg_rca32_ha9_y1 = f_s_dadda_pg_rca32_ha9_f_s_dadda_pg_rca32_and_1_10_y0 & f_s_dadda_pg_rca32_ha9_f_s_dadda_pg_rca32_and_0_11_y0;
  assign f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_ha9_y1 = f_s_dadda_pg_rca32_ha9_y1;
  assign f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_fa30_y4 = f_s_dadda_pg_rca32_fa30_y4;
  assign f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_fa29_y4 = f_s_dadda_pg_rca32_fa29_y4;
  assign f_s_dadda_pg_rca32_fa31_y0 = f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_ha9_y1 ^ f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_fa30_y4;
  assign f_s_dadda_pg_rca32_fa31_y1 = f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_ha9_y1 & f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_fa30_y4;
  assign f_s_dadda_pg_rca32_fa31_y2 = f_s_dadda_pg_rca32_fa31_y0 ^ f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_fa29_y4;
  assign f_s_dadda_pg_rca32_fa31_y3 = f_s_dadda_pg_rca32_fa31_y0 & f_s_dadda_pg_rca32_fa31_f_s_dadda_pg_rca32_fa29_y4;
  assign f_s_dadda_pg_rca32_fa31_y4 = f_s_dadda_pg_rca32_fa31_y1 | f_s_dadda_pg_rca32_fa31_y3;
  assign f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa28_y4 = f_s_dadda_pg_rca32_fa28_y4;
  assign f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa27_y4 = f_s_dadda_pg_rca32_fa27_y4;
  assign f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa26_y4 = f_s_dadda_pg_rca32_fa26_y4;
  assign f_s_dadda_pg_rca32_fa32_y0 = f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa28_y4 ^ f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa27_y4;
  assign f_s_dadda_pg_rca32_fa32_y1 = f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa28_y4 & f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa27_y4;
  assign f_s_dadda_pg_rca32_fa32_y2 = f_s_dadda_pg_rca32_fa32_y0 ^ f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa26_y4;
  assign f_s_dadda_pg_rca32_fa32_y3 = f_s_dadda_pg_rca32_fa32_y0 & f_s_dadda_pg_rca32_fa32_f_s_dadda_pg_rca32_fa26_y4;
  assign f_s_dadda_pg_rca32_fa32_y4 = f_s_dadda_pg_rca32_fa32_y1 | f_s_dadda_pg_rca32_fa32_y3;
  assign f_s_dadda_pg_rca32_and_12_0_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_12_0_y0 = f_s_dadda_pg_rca32_and_12_0_a_12 & f_s_dadda_pg_rca32_and_12_0_b_0;
  assign f_s_dadda_pg_rca32_and_11_1_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_11_1_y0 = f_s_dadda_pg_rca32_and_11_1_a_11 & f_s_dadda_pg_rca32_and_11_1_b_1;
  assign f_s_dadda_pg_rca32_and_10_2_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_10_2_y0 = f_s_dadda_pg_rca32_and_10_2_a_10 & f_s_dadda_pg_rca32_and_10_2_b_2;
  assign f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_12_0_y0 = f_s_dadda_pg_rca32_and_12_0_y0;
  assign f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_11_1_y0 = f_s_dadda_pg_rca32_and_11_1_y0;
  assign f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_10_2_y0 = f_s_dadda_pg_rca32_and_10_2_y0;
  assign f_s_dadda_pg_rca32_fa33_y0 = f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_12_0_y0 ^ f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_11_1_y0;
  assign f_s_dadda_pg_rca32_fa33_y1 = f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_12_0_y0 & f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_11_1_y0;
  assign f_s_dadda_pg_rca32_fa33_y2 = f_s_dadda_pg_rca32_fa33_y0 ^ f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_10_2_y0;
  assign f_s_dadda_pg_rca32_fa33_y3 = f_s_dadda_pg_rca32_fa33_y0 & f_s_dadda_pg_rca32_fa33_f_s_dadda_pg_rca32_and_10_2_y0;
  assign f_s_dadda_pg_rca32_fa33_y4 = f_s_dadda_pg_rca32_fa33_y1 | f_s_dadda_pg_rca32_fa33_y3;
  assign f_s_dadda_pg_rca32_and_9_3_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_9_3_y0 = f_s_dadda_pg_rca32_and_9_3_a_9 & f_s_dadda_pg_rca32_and_9_3_b_3;
  assign f_s_dadda_pg_rca32_and_8_4_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_8_4_y0 = f_s_dadda_pg_rca32_and_8_4_a_8 & f_s_dadda_pg_rca32_and_8_4_b_4;
  assign f_s_dadda_pg_rca32_and_7_5_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_7_5_y0 = f_s_dadda_pg_rca32_and_7_5_a_7 & f_s_dadda_pg_rca32_and_7_5_b_5;
  assign f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_9_3_y0 = f_s_dadda_pg_rca32_and_9_3_y0;
  assign f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_8_4_y0 = f_s_dadda_pg_rca32_and_8_4_y0;
  assign f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_7_5_y0 = f_s_dadda_pg_rca32_and_7_5_y0;
  assign f_s_dadda_pg_rca32_fa34_y0 = f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_9_3_y0 ^ f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_8_4_y0;
  assign f_s_dadda_pg_rca32_fa34_y1 = f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_9_3_y0 & f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_8_4_y0;
  assign f_s_dadda_pg_rca32_fa34_y2 = f_s_dadda_pg_rca32_fa34_y0 ^ f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_7_5_y0;
  assign f_s_dadda_pg_rca32_fa34_y3 = f_s_dadda_pg_rca32_fa34_y0 & f_s_dadda_pg_rca32_fa34_f_s_dadda_pg_rca32_and_7_5_y0;
  assign f_s_dadda_pg_rca32_fa34_y4 = f_s_dadda_pg_rca32_fa34_y1 | f_s_dadda_pg_rca32_fa34_y3;
  assign f_s_dadda_pg_rca32_and_6_6_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_6_6_y0 = f_s_dadda_pg_rca32_and_6_6_a_6 & f_s_dadda_pg_rca32_and_6_6_b_6;
  assign f_s_dadda_pg_rca32_and_5_7_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_5_7_y0 = f_s_dadda_pg_rca32_and_5_7_a_5 & f_s_dadda_pg_rca32_and_5_7_b_7;
  assign f_s_dadda_pg_rca32_and_4_8_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_4_8_y0 = f_s_dadda_pg_rca32_and_4_8_a_4 & f_s_dadda_pg_rca32_and_4_8_b_8;
  assign f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_6_6_y0 = f_s_dadda_pg_rca32_and_6_6_y0;
  assign f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_5_7_y0 = f_s_dadda_pg_rca32_and_5_7_y0;
  assign f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_4_8_y0 = f_s_dadda_pg_rca32_and_4_8_y0;
  assign f_s_dadda_pg_rca32_fa35_y0 = f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_6_6_y0 ^ f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_5_7_y0;
  assign f_s_dadda_pg_rca32_fa35_y1 = f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_6_6_y0 & f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_5_7_y0;
  assign f_s_dadda_pg_rca32_fa35_y2 = f_s_dadda_pg_rca32_fa35_y0 ^ f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_4_8_y0;
  assign f_s_dadda_pg_rca32_fa35_y3 = f_s_dadda_pg_rca32_fa35_y0 & f_s_dadda_pg_rca32_fa35_f_s_dadda_pg_rca32_and_4_8_y0;
  assign f_s_dadda_pg_rca32_fa35_y4 = f_s_dadda_pg_rca32_fa35_y1 | f_s_dadda_pg_rca32_fa35_y3;
  assign f_s_dadda_pg_rca32_and_3_9_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_3_9_y0 = f_s_dadda_pg_rca32_and_3_9_a_3 & f_s_dadda_pg_rca32_and_3_9_b_9;
  assign f_s_dadda_pg_rca32_and_2_10_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_2_10_y0 = f_s_dadda_pg_rca32_and_2_10_a_2 & f_s_dadda_pg_rca32_and_2_10_b_10;
  assign f_s_dadda_pg_rca32_and_1_11_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_1_11_y0 = f_s_dadda_pg_rca32_and_1_11_a_1 & f_s_dadda_pg_rca32_and_1_11_b_11;
  assign f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_3_9_y0 = f_s_dadda_pg_rca32_and_3_9_y0;
  assign f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_2_10_y0 = f_s_dadda_pg_rca32_and_2_10_y0;
  assign f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_1_11_y0 = f_s_dadda_pg_rca32_and_1_11_y0;
  assign f_s_dadda_pg_rca32_fa36_y0 = f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_3_9_y0 ^ f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_2_10_y0;
  assign f_s_dadda_pg_rca32_fa36_y1 = f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_3_9_y0 & f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_2_10_y0;
  assign f_s_dadda_pg_rca32_fa36_y2 = f_s_dadda_pg_rca32_fa36_y0 ^ f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_1_11_y0;
  assign f_s_dadda_pg_rca32_fa36_y3 = f_s_dadda_pg_rca32_fa36_y0 & f_s_dadda_pg_rca32_fa36_f_s_dadda_pg_rca32_and_1_11_y0;
  assign f_s_dadda_pg_rca32_fa36_y4 = f_s_dadda_pg_rca32_fa36_y1 | f_s_dadda_pg_rca32_fa36_y3;
  assign f_s_dadda_pg_rca32_and_0_12_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_0_12_y0 = f_s_dadda_pg_rca32_and_0_12_a_0 & f_s_dadda_pg_rca32_and_0_12_b_12;
  assign f_s_dadda_pg_rca32_ha10_f_s_dadda_pg_rca32_and_0_12_y0 = f_s_dadda_pg_rca32_and_0_12_y0;
  assign f_s_dadda_pg_rca32_ha10_f_s_dadda_pg_rca32_fa31_y2 = f_s_dadda_pg_rca32_fa31_y2;
  assign f_s_dadda_pg_rca32_ha10_y0 = f_s_dadda_pg_rca32_ha10_f_s_dadda_pg_rca32_and_0_12_y0 ^ f_s_dadda_pg_rca32_ha10_f_s_dadda_pg_rca32_fa31_y2;
  assign f_s_dadda_pg_rca32_ha10_y1 = f_s_dadda_pg_rca32_ha10_f_s_dadda_pg_rca32_and_0_12_y0 & f_s_dadda_pg_rca32_ha10_f_s_dadda_pg_rca32_fa31_y2;
  assign f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_ha10_y1 = f_s_dadda_pg_rca32_ha10_y1;
  assign f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_fa36_y4 = f_s_dadda_pg_rca32_fa36_y4;
  assign f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_fa35_y4 = f_s_dadda_pg_rca32_fa35_y4;
  assign f_s_dadda_pg_rca32_fa37_y0 = f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_ha10_y1 ^ f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_fa36_y4;
  assign f_s_dadda_pg_rca32_fa37_y1 = f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_ha10_y1 & f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_fa36_y4;
  assign f_s_dadda_pg_rca32_fa37_y2 = f_s_dadda_pg_rca32_fa37_y0 ^ f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_fa35_y4;
  assign f_s_dadda_pg_rca32_fa37_y3 = f_s_dadda_pg_rca32_fa37_y0 & f_s_dadda_pg_rca32_fa37_f_s_dadda_pg_rca32_fa35_y4;
  assign f_s_dadda_pg_rca32_fa37_y4 = f_s_dadda_pg_rca32_fa37_y1 | f_s_dadda_pg_rca32_fa37_y3;
  assign f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa34_y4 = f_s_dadda_pg_rca32_fa34_y4;
  assign f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa33_y4 = f_s_dadda_pg_rca32_fa33_y4;
  assign f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa32_y4 = f_s_dadda_pg_rca32_fa32_y4;
  assign f_s_dadda_pg_rca32_fa38_y0 = f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa34_y4 ^ f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa33_y4;
  assign f_s_dadda_pg_rca32_fa38_y1 = f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa34_y4 & f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa33_y4;
  assign f_s_dadda_pg_rca32_fa38_y2 = f_s_dadda_pg_rca32_fa38_y0 ^ f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa32_y4;
  assign f_s_dadda_pg_rca32_fa38_y3 = f_s_dadda_pg_rca32_fa38_y0 & f_s_dadda_pg_rca32_fa38_f_s_dadda_pg_rca32_fa32_y4;
  assign f_s_dadda_pg_rca32_fa38_y4 = f_s_dadda_pg_rca32_fa38_y1 | f_s_dadda_pg_rca32_fa38_y3;
  assign f_s_dadda_pg_rca32_and_13_0_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_13_0_y0 = f_s_dadda_pg_rca32_and_13_0_a_13 & f_s_dadda_pg_rca32_and_13_0_b_0;
  assign f_s_dadda_pg_rca32_and_12_1_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_12_1_y0 = f_s_dadda_pg_rca32_and_12_1_a_12 & f_s_dadda_pg_rca32_and_12_1_b_1;
  assign f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_fa31_y4 = f_s_dadda_pg_rca32_fa31_y4;
  assign f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_and_13_0_y0 = f_s_dadda_pg_rca32_and_13_0_y0;
  assign f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_and_12_1_y0 = f_s_dadda_pg_rca32_and_12_1_y0;
  assign f_s_dadda_pg_rca32_fa39_y0 = f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_fa31_y4 ^ f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_and_13_0_y0;
  assign f_s_dadda_pg_rca32_fa39_y1 = f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_fa31_y4 & f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_and_13_0_y0;
  assign f_s_dadda_pg_rca32_fa39_y2 = f_s_dadda_pg_rca32_fa39_y0 ^ f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_and_12_1_y0;
  assign f_s_dadda_pg_rca32_fa39_y3 = f_s_dadda_pg_rca32_fa39_y0 & f_s_dadda_pg_rca32_fa39_f_s_dadda_pg_rca32_and_12_1_y0;
  assign f_s_dadda_pg_rca32_fa39_y4 = f_s_dadda_pg_rca32_fa39_y1 | f_s_dadda_pg_rca32_fa39_y3;
  assign f_s_dadda_pg_rca32_and_11_2_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_11_2_y0 = f_s_dadda_pg_rca32_and_11_2_a_11 & f_s_dadda_pg_rca32_and_11_2_b_2;
  assign f_s_dadda_pg_rca32_and_10_3_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_10_3_y0 = f_s_dadda_pg_rca32_and_10_3_a_10 & f_s_dadda_pg_rca32_and_10_3_b_3;
  assign f_s_dadda_pg_rca32_and_9_4_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_9_4_y0 = f_s_dadda_pg_rca32_and_9_4_a_9 & f_s_dadda_pg_rca32_and_9_4_b_4;
  assign f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_11_2_y0 = f_s_dadda_pg_rca32_and_11_2_y0;
  assign f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_10_3_y0 = f_s_dadda_pg_rca32_and_10_3_y0;
  assign f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_9_4_y0 = f_s_dadda_pg_rca32_and_9_4_y0;
  assign f_s_dadda_pg_rca32_fa40_y0 = f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_11_2_y0 ^ f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_10_3_y0;
  assign f_s_dadda_pg_rca32_fa40_y1 = f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_11_2_y0 & f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_10_3_y0;
  assign f_s_dadda_pg_rca32_fa40_y2 = f_s_dadda_pg_rca32_fa40_y0 ^ f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_9_4_y0;
  assign f_s_dadda_pg_rca32_fa40_y3 = f_s_dadda_pg_rca32_fa40_y0 & f_s_dadda_pg_rca32_fa40_f_s_dadda_pg_rca32_and_9_4_y0;
  assign f_s_dadda_pg_rca32_fa40_y4 = f_s_dadda_pg_rca32_fa40_y1 | f_s_dadda_pg_rca32_fa40_y3;
  assign f_s_dadda_pg_rca32_and_8_5_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_8_5_y0 = f_s_dadda_pg_rca32_and_8_5_a_8 & f_s_dadda_pg_rca32_and_8_5_b_5;
  assign f_s_dadda_pg_rca32_and_7_6_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_7_6_y0 = f_s_dadda_pg_rca32_and_7_6_a_7 & f_s_dadda_pg_rca32_and_7_6_b_6;
  assign f_s_dadda_pg_rca32_and_6_7_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_6_7_y0 = f_s_dadda_pg_rca32_and_6_7_a_6 & f_s_dadda_pg_rca32_and_6_7_b_7;
  assign f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_8_5_y0 = f_s_dadda_pg_rca32_and_8_5_y0;
  assign f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_7_6_y0 = f_s_dadda_pg_rca32_and_7_6_y0;
  assign f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_6_7_y0 = f_s_dadda_pg_rca32_and_6_7_y0;
  assign f_s_dadda_pg_rca32_fa41_y0 = f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_8_5_y0 ^ f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_7_6_y0;
  assign f_s_dadda_pg_rca32_fa41_y1 = f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_8_5_y0 & f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_7_6_y0;
  assign f_s_dadda_pg_rca32_fa41_y2 = f_s_dadda_pg_rca32_fa41_y0 ^ f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_6_7_y0;
  assign f_s_dadda_pg_rca32_fa41_y3 = f_s_dadda_pg_rca32_fa41_y0 & f_s_dadda_pg_rca32_fa41_f_s_dadda_pg_rca32_and_6_7_y0;
  assign f_s_dadda_pg_rca32_fa41_y4 = f_s_dadda_pg_rca32_fa41_y1 | f_s_dadda_pg_rca32_fa41_y3;
  assign f_s_dadda_pg_rca32_and_5_8_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_5_8_y0 = f_s_dadda_pg_rca32_and_5_8_a_5 & f_s_dadda_pg_rca32_and_5_8_b_8;
  assign f_s_dadda_pg_rca32_and_4_9_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_4_9_y0 = f_s_dadda_pg_rca32_and_4_9_a_4 & f_s_dadda_pg_rca32_and_4_9_b_9;
  assign f_s_dadda_pg_rca32_and_3_10_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_3_10_y0 = f_s_dadda_pg_rca32_and_3_10_a_3 & f_s_dadda_pg_rca32_and_3_10_b_10;
  assign f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_5_8_y0 = f_s_dadda_pg_rca32_and_5_8_y0;
  assign f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_4_9_y0 = f_s_dadda_pg_rca32_and_4_9_y0;
  assign f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_3_10_y0 = f_s_dadda_pg_rca32_and_3_10_y0;
  assign f_s_dadda_pg_rca32_fa42_y0 = f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_5_8_y0 ^ f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_4_9_y0;
  assign f_s_dadda_pg_rca32_fa42_y1 = f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_5_8_y0 & f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_4_9_y0;
  assign f_s_dadda_pg_rca32_fa42_y2 = f_s_dadda_pg_rca32_fa42_y0 ^ f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_3_10_y0;
  assign f_s_dadda_pg_rca32_fa42_y3 = f_s_dadda_pg_rca32_fa42_y0 & f_s_dadda_pg_rca32_fa42_f_s_dadda_pg_rca32_and_3_10_y0;
  assign f_s_dadda_pg_rca32_fa42_y4 = f_s_dadda_pg_rca32_fa42_y1 | f_s_dadda_pg_rca32_fa42_y3;
  assign f_s_dadda_pg_rca32_and_2_11_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_2_11_y0 = f_s_dadda_pg_rca32_and_2_11_a_2 & f_s_dadda_pg_rca32_and_2_11_b_11;
  assign f_s_dadda_pg_rca32_and_1_12_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_1_12_y0 = f_s_dadda_pg_rca32_and_1_12_a_1 & f_s_dadda_pg_rca32_and_1_12_b_12;
  assign f_s_dadda_pg_rca32_and_0_13_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_0_13_y0 = f_s_dadda_pg_rca32_and_0_13_a_0 & f_s_dadda_pg_rca32_and_0_13_b_13;
  assign f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_2_11_y0 = f_s_dadda_pg_rca32_and_2_11_y0;
  assign f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_1_12_y0 = f_s_dadda_pg_rca32_and_1_12_y0;
  assign f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_0_13_y0 = f_s_dadda_pg_rca32_and_0_13_y0;
  assign f_s_dadda_pg_rca32_fa43_y0 = f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_2_11_y0 ^ f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_1_12_y0;
  assign f_s_dadda_pg_rca32_fa43_y1 = f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_2_11_y0 & f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_1_12_y0;
  assign f_s_dadda_pg_rca32_fa43_y2 = f_s_dadda_pg_rca32_fa43_y0 ^ f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_0_13_y0;
  assign f_s_dadda_pg_rca32_fa43_y3 = f_s_dadda_pg_rca32_fa43_y0 & f_s_dadda_pg_rca32_fa43_f_s_dadda_pg_rca32_and_0_13_y0;
  assign f_s_dadda_pg_rca32_fa43_y4 = f_s_dadda_pg_rca32_fa43_y1 | f_s_dadda_pg_rca32_fa43_y3;
  assign f_s_dadda_pg_rca32_ha11_f_s_dadda_pg_rca32_fa37_y2 = f_s_dadda_pg_rca32_fa37_y2;
  assign f_s_dadda_pg_rca32_ha11_f_s_dadda_pg_rca32_fa38_y2 = f_s_dadda_pg_rca32_fa38_y2;
  assign f_s_dadda_pg_rca32_ha11_y0 = f_s_dadda_pg_rca32_ha11_f_s_dadda_pg_rca32_fa37_y2 ^ f_s_dadda_pg_rca32_ha11_f_s_dadda_pg_rca32_fa38_y2;
  assign f_s_dadda_pg_rca32_ha11_y1 = f_s_dadda_pg_rca32_ha11_f_s_dadda_pg_rca32_fa37_y2 & f_s_dadda_pg_rca32_ha11_f_s_dadda_pg_rca32_fa38_y2;
  assign f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_ha11_y1 = f_s_dadda_pg_rca32_ha11_y1;
  assign f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_fa43_y4 = f_s_dadda_pg_rca32_fa43_y4;
  assign f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_fa42_y4 = f_s_dadda_pg_rca32_fa42_y4;
  assign f_s_dadda_pg_rca32_fa44_y0 = f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_ha11_y1 ^ f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_fa43_y4;
  assign f_s_dadda_pg_rca32_fa44_y1 = f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_ha11_y1 & f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_fa43_y4;
  assign f_s_dadda_pg_rca32_fa44_y2 = f_s_dadda_pg_rca32_fa44_y0 ^ f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_fa42_y4;
  assign f_s_dadda_pg_rca32_fa44_y3 = f_s_dadda_pg_rca32_fa44_y0 & f_s_dadda_pg_rca32_fa44_f_s_dadda_pg_rca32_fa42_y4;
  assign f_s_dadda_pg_rca32_fa44_y4 = f_s_dadda_pg_rca32_fa44_y1 | f_s_dadda_pg_rca32_fa44_y3;
  assign f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa41_y4 = f_s_dadda_pg_rca32_fa41_y4;
  assign f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa40_y4 = f_s_dadda_pg_rca32_fa40_y4;
  assign f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa39_y4 = f_s_dadda_pg_rca32_fa39_y4;
  assign f_s_dadda_pg_rca32_fa45_y0 = f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa41_y4 ^ f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa40_y4;
  assign f_s_dadda_pg_rca32_fa45_y1 = f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa41_y4 & f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa40_y4;
  assign f_s_dadda_pg_rca32_fa45_y2 = f_s_dadda_pg_rca32_fa45_y0 ^ f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa39_y4;
  assign f_s_dadda_pg_rca32_fa45_y3 = f_s_dadda_pg_rca32_fa45_y0 & f_s_dadda_pg_rca32_fa45_f_s_dadda_pg_rca32_fa39_y4;
  assign f_s_dadda_pg_rca32_fa45_y4 = f_s_dadda_pg_rca32_fa45_y1 | f_s_dadda_pg_rca32_fa45_y3;
  assign f_s_dadda_pg_rca32_and_14_0_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_14_0_y0 = f_s_dadda_pg_rca32_and_14_0_a_14 & f_s_dadda_pg_rca32_and_14_0_b_0;
  assign f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_fa38_y4 = f_s_dadda_pg_rca32_fa38_y4;
  assign f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_fa37_y4 = f_s_dadda_pg_rca32_fa37_y4;
  assign f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_and_14_0_y0 = f_s_dadda_pg_rca32_and_14_0_y0;
  assign f_s_dadda_pg_rca32_fa46_y0 = f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_fa38_y4 ^ f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_fa37_y4;
  assign f_s_dadda_pg_rca32_fa46_y1 = f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_fa38_y4 & f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_fa37_y4;
  assign f_s_dadda_pg_rca32_fa46_y2 = f_s_dadda_pg_rca32_fa46_y0 ^ f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_and_14_0_y0;
  assign f_s_dadda_pg_rca32_fa46_y3 = f_s_dadda_pg_rca32_fa46_y0 & f_s_dadda_pg_rca32_fa46_f_s_dadda_pg_rca32_and_14_0_y0;
  assign f_s_dadda_pg_rca32_fa46_y4 = f_s_dadda_pg_rca32_fa46_y1 | f_s_dadda_pg_rca32_fa46_y3;
  assign f_s_dadda_pg_rca32_and_13_1_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_13_1_y0 = f_s_dadda_pg_rca32_and_13_1_a_13 & f_s_dadda_pg_rca32_and_13_1_b_1;
  assign f_s_dadda_pg_rca32_and_12_2_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_12_2_y0 = f_s_dadda_pg_rca32_and_12_2_a_12 & f_s_dadda_pg_rca32_and_12_2_b_2;
  assign f_s_dadda_pg_rca32_and_11_3_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_11_3_y0 = f_s_dadda_pg_rca32_and_11_3_a_11 & f_s_dadda_pg_rca32_and_11_3_b_3;
  assign f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_13_1_y0 = f_s_dadda_pg_rca32_and_13_1_y0;
  assign f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_12_2_y0 = f_s_dadda_pg_rca32_and_12_2_y0;
  assign f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_11_3_y0 = f_s_dadda_pg_rca32_and_11_3_y0;
  assign f_s_dadda_pg_rca32_fa47_y0 = f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_13_1_y0 ^ f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_12_2_y0;
  assign f_s_dadda_pg_rca32_fa47_y1 = f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_13_1_y0 & f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_12_2_y0;
  assign f_s_dadda_pg_rca32_fa47_y2 = f_s_dadda_pg_rca32_fa47_y0 ^ f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_11_3_y0;
  assign f_s_dadda_pg_rca32_fa47_y3 = f_s_dadda_pg_rca32_fa47_y0 & f_s_dadda_pg_rca32_fa47_f_s_dadda_pg_rca32_and_11_3_y0;
  assign f_s_dadda_pg_rca32_fa47_y4 = f_s_dadda_pg_rca32_fa47_y1 | f_s_dadda_pg_rca32_fa47_y3;
  assign f_s_dadda_pg_rca32_and_10_4_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_10_4_y0 = f_s_dadda_pg_rca32_and_10_4_a_10 & f_s_dadda_pg_rca32_and_10_4_b_4;
  assign f_s_dadda_pg_rca32_and_9_5_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_9_5_y0 = f_s_dadda_pg_rca32_and_9_5_a_9 & f_s_dadda_pg_rca32_and_9_5_b_5;
  assign f_s_dadda_pg_rca32_and_8_6_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_8_6_y0 = f_s_dadda_pg_rca32_and_8_6_a_8 & f_s_dadda_pg_rca32_and_8_6_b_6;
  assign f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_10_4_y0 = f_s_dadda_pg_rca32_and_10_4_y0;
  assign f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_9_5_y0 = f_s_dadda_pg_rca32_and_9_5_y0;
  assign f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_8_6_y0 = f_s_dadda_pg_rca32_and_8_6_y0;
  assign f_s_dadda_pg_rca32_fa48_y0 = f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_10_4_y0 ^ f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_9_5_y0;
  assign f_s_dadda_pg_rca32_fa48_y1 = f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_10_4_y0 & f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_9_5_y0;
  assign f_s_dadda_pg_rca32_fa48_y2 = f_s_dadda_pg_rca32_fa48_y0 ^ f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_8_6_y0;
  assign f_s_dadda_pg_rca32_fa48_y3 = f_s_dadda_pg_rca32_fa48_y0 & f_s_dadda_pg_rca32_fa48_f_s_dadda_pg_rca32_and_8_6_y0;
  assign f_s_dadda_pg_rca32_fa48_y4 = f_s_dadda_pg_rca32_fa48_y1 | f_s_dadda_pg_rca32_fa48_y3;
  assign f_s_dadda_pg_rca32_and_7_7_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_7_7_y0 = f_s_dadda_pg_rca32_and_7_7_a_7 & f_s_dadda_pg_rca32_and_7_7_b_7;
  assign f_s_dadda_pg_rca32_and_6_8_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_6_8_y0 = f_s_dadda_pg_rca32_and_6_8_a_6 & f_s_dadda_pg_rca32_and_6_8_b_8;
  assign f_s_dadda_pg_rca32_and_5_9_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_5_9_y0 = f_s_dadda_pg_rca32_and_5_9_a_5 & f_s_dadda_pg_rca32_and_5_9_b_9;
  assign f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_7_7_y0 = f_s_dadda_pg_rca32_and_7_7_y0;
  assign f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_6_8_y0 = f_s_dadda_pg_rca32_and_6_8_y0;
  assign f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_5_9_y0 = f_s_dadda_pg_rca32_and_5_9_y0;
  assign f_s_dadda_pg_rca32_fa49_y0 = f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_7_7_y0 ^ f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_6_8_y0;
  assign f_s_dadda_pg_rca32_fa49_y1 = f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_7_7_y0 & f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_6_8_y0;
  assign f_s_dadda_pg_rca32_fa49_y2 = f_s_dadda_pg_rca32_fa49_y0 ^ f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_5_9_y0;
  assign f_s_dadda_pg_rca32_fa49_y3 = f_s_dadda_pg_rca32_fa49_y0 & f_s_dadda_pg_rca32_fa49_f_s_dadda_pg_rca32_and_5_9_y0;
  assign f_s_dadda_pg_rca32_fa49_y4 = f_s_dadda_pg_rca32_fa49_y1 | f_s_dadda_pg_rca32_fa49_y3;
  assign f_s_dadda_pg_rca32_and_4_10_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_4_10_y0 = f_s_dadda_pg_rca32_and_4_10_a_4 & f_s_dadda_pg_rca32_and_4_10_b_10;
  assign f_s_dadda_pg_rca32_and_3_11_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_3_11_y0 = f_s_dadda_pg_rca32_and_3_11_a_3 & f_s_dadda_pg_rca32_and_3_11_b_11;
  assign f_s_dadda_pg_rca32_and_2_12_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_2_12_y0 = f_s_dadda_pg_rca32_and_2_12_a_2 & f_s_dadda_pg_rca32_and_2_12_b_12;
  assign f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_4_10_y0 = f_s_dadda_pg_rca32_and_4_10_y0;
  assign f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_3_11_y0 = f_s_dadda_pg_rca32_and_3_11_y0;
  assign f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_2_12_y0 = f_s_dadda_pg_rca32_and_2_12_y0;
  assign f_s_dadda_pg_rca32_fa50_y0 = f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_4_10_y0 ^ f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_3_11_y0;
  assign f_s_dadda_pg_rca32_fa50_y1 = f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_4_10_y0 & f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_3_11_y0;
  assign f_s_dadda_pg_rca32_fa50_y2 = f_s_dadda_pg_rca32_fa50_y0 ^ f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_2_12_y0;
  assign f_s_dadda_pg_rca32_fa50_y3 = f_s_dadda_pg_rca32_fa50_y0 & f_s_dadda_pg_rca32_fa50_f_s_dadda_pg_rca32_and_2_12_y0;
  assign f_s_dadda_pg_rca32_fa50_y4 = f_s_dadda_pg_rca32_fa50_y1 | f_s_dadda_pg_rca32_fa50_y3;
  assign f_s_dadda_pg_rca32_and_1_13_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_1_13_y0 = f_s_dadda_pg_rca32_and_1_13_a_1 & f_s_dadda_pg_rca32_and_1_13_b_13;
  assign f_s_dadda_pg_rca32_and_0_14_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_0_14_y0 = f_s_dadda_pg_rca32_and_0_14_a_0 & f_s_dadda_pg_rca32_and_0_14_b_14;
  assign f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_and_1_13_y0 = f_s_dadda_pg_rca32_and_1_13_y0;
  assign f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_and_0_14_y0 = f_s_dadda_pg_rca32_and_0_14_y0;
  assign f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_fa44_y2 = f_s_dadda_pg_rca32_fa44_y2;
  assign f_s_dadda_pg_rca32_fa51_y0 = f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_and_1_13_y0 ^ f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_and_0_14_y0;
  assign f_s_dadda_pg_rca32_fa51_y1 = f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_and_1_13_y0 & f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_and_0_14_y0;
  assign f_s_dadda_pg_rca32_fa51_y2 = f_s_dadda_pg_rca32_fa51_y0 ^ f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_fa44_y2;
  assign f_s_dadda_pg_rca32_fa51_y3 = f_s_dadda_pg_rca32_fa51_y0 & f_s_dadda_pg_rca32_fa51_f_s_dadda_pg_rca32_fa44_y2;
  assign f_s_dadda_pg_rca32_fa51_y4 = f_s_dadda_pg_rca32_fa51_y1 | f_s_dadda_pg_rca32_fa51_y3;
  assign f_s_dadda_pg_rca32_ha12_f_s_dadda_pg_rca32_fa45_y2 = f_s_dadda_pg_rca32_fa45_y2;
  assign f_s_dadda_pg_rca32_ha12_f_s_dadda_pg_rca32_fa46_y2 = f_s_dadda_pg_rca32_fa46_y2;
  assign f_s_dadda_pg_rca32_ha12_y0 = f_s_dadda_pg_rca32_ha12_f_s_dadda_pg_rca32_fa45_y2 ^ f_s_dadda_pg_rca32_ha12_f_s_dadda_pg_rca32_fa46_y2;
  assign f_s_dadda_pg_rca32_ha12_y1 = f_s_dadda_pg_rca32_ha12_f_s_dadda_pg_rca32_fa45_y2 & f_s_dadda_pg_rca32_ha12_f_s_dadda_pg_rca32_fa46_y2;
  assign f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_ha12_y1 = f_s_dadda_pg_rca32_ha12_y1;
  assign f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_fa51_y4 = f_s_dadda_pg_rca32_fa51_y4;
  assign f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_fa50_y4 = f_s_dadda_pg_rca32_fa50_y4;
  assign f_s_dadda_pg_rca32_fa52_y0 = f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_ha12_y1 ^ f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_fa51_y4;
  assign f_s_dadda_pg_rca32_fa52_y1 = f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_ha12_y1 & f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_fa51_y4;
  assign f_s_dadda_pg_rca32_fa52_y2 = f_s_dadda_pg_rca32_fa52_y0 ^ f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_fa50_y4;
  assign f_s_dadda_pg_rca32_fa52_y3 = f_s_dadda_pg_rca32_fa52_y0 & f_s_dadda_pg_rca32_fa52_f_s_dadda_pg_rca32_fa50_y4;
  assign f_s_dadda_pg_rca32_fa52_y4 = f_s_dadda_pg_rca32_fa52_y1 | f_s_dadda_pg_rca32_fa52_y3;
  assign f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa49_y4 = f_s_dadda_pg_rca32_fa49_y4;
  assign f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa48_y4 = f_s_dadda_pg_rca32_fa48_y4;
  assign f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa47_y4 = f_s_dadda_pg_rca32_fa47_y4;
  assign f_s_dadda_pg_rca32_fa53_y0 = f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa49_y4 ^ f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa48_y4;
  assign f_s_dadda_pg_rca32_fa53_y1 = f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa49_y4 & f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa48_y4;
  assign f_s_dadda_pg_rca32_fa53_y2 = f_s_dadda_pg_rca32_fa53_y0 ^ f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa47_y4;
  assign f_s_dadda_pg_rca32_fa53_y3 = f_s_dadda_pg_rca32_fa53_y0 & f_s_dadda_pg_rca32_fa53_f_s_dadda_pg_rca32_fa47_y4;
  assign f_s_dadda_pg_rca32_fa53_y4 = f_s_dadda_pg_rca32_fa53_y1 | f_s_dadda_pg_rca32_fa53_y3;
  assign f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa46_y4 = f_s_dadda_pg_rca32_fa46_y4;
  assign f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa45_y4 = f_s_dadda_pg_rca32_fa45_y4;
  assign f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa44_y4 = f_s_dadda_pg_rca32_fa44_y4;
  assign f_s_dadda_pg_rca32_fa54_y0 = f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa46_y4 ^ f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa45_y4;
  assign f_s_dadda_pg_rca32_fa54_y1 = f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa46_y4 & f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa45_y4;
  assign f_s_dadda_pg_rca32_fa54_y2 = f_s_dadda_pg_rca32_fa54_y0 ^ f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa44_y4;
  assign f_s_dadda_pg_rca32_fa54_y3 = f_s_dadda_pg_rca32_fa54_y0 & f_s_dadda_pg_rca32_fa54_f_s_dadda_pg_rca32_fa44_y4;
  assign f_s_dadda_pg_rca32_fa54_y4 = f_s_dadda_pg_rca32_fa54_y1 | f_s_dadda_pg_rca32_fa54_y3;
  assign f_s_dadda_pg_rca32_and_15_0_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_15_0_y0 = f_s_dadda_pg_rca32_and_15_0_a_15 & f_s_dadda_pg_rca32_and_15_0_b_0;
  assign f_s_dadda_pg_rca32_and_14_1_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_14_1_y0 = f_s_dadda_pg_rca32_and_14_1_a_14 & f_s_dadda_pg_rca32_and_14_1_b_1;
  assign f_s_dadda_pg_rca32_and_13_2_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_13_2_y0 = f_s_dadda_pg_rca32_and_13_2_a_13 & f_s_dadda_pg_rca32_and_13_2_b_2;
  assign f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_15_0_y0 = f_s_dadda_pg_rca32_and_15_0_y0;
  assign f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_14_1_y0 = f_s_dadda_pg_rca32_and_14_1_y0;
  assign f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_13_2_y0 = f_s_dadda_pg_rca32_and_13_2_y0;
  assign f_s_dadda_pg_rca32_fa55_y0 = f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_15_0_y0 ^ f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_14_1_y0;
  assign f_s_dadda_pg_rca32_fa55_y1 = f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_15_0_y0 & f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_14_1_y0;
  assign f_s_dadda_pg_rca32_fa55_y2 = f_s_dadda_pg_rca32_fa55_y0 ^ f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_13_2_y0;
  assign f_s_dadda_pg_rca32_fa55_y3 = f_s_dadda_pg_rca32_fa55_y0 & f_s_dadda_pg_rca32_fa55_f_s_dadda_pg_rca32_and_13_2_y0;
  assign f_s_dadda_pg_rca32_fa55_y4 = f_s_dadda_pg_rca32_fa55_y1 | f_s_dadda_pg_rca32_fa55_y3;
  assign f_s_dadda_pg_rca32_and_12_3_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_12_3_y0 = f_s_dadda_pg_rca32_and_12_3_a_12 & f_s_dadda_pg_rca32_and_12_3_b_3;
  assign f_s_dadda_pg_rca32_and_11_4_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_11_4_y0 = f_s_dadda_pg_rca32_and_11_4_a_11 & f_s_dadda_pg_rca32_and_11_4_b_4;
  assign f_s_dadda_pg_rca32_and_10_5_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_10_5_y0 = f_s_dadda_pg_rca32_and_10_5_a_10 & f_s_dadda_pg_rca32_and_10_5_b_5;
  assign f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_12_3_y0 = f_s_dadda_pg_rca32_and_12_3_y0;
  assign f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_11_4_y0 = f_s_dadda_pg_rca32_and_11_4_y0;
  assign f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_10_5_y0 = f_s_dadda_pg_rca32_and_10_5_y0;
  assign f_s_dadda_pg_rca32_fa56_y0 = f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_12_3_y0 ^ f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_11_4_y0;
  assign f_s_dadda_pg_rca32_fa56_y1 = f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_12_3_y0 & f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_11_4_y0;
  assign f_s_dadda_pg_rca32_fa56_y2 = f_s_dadda_pg_rca32_fa56_y0 ^ f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_10_5_y0;
  assign f_s_dadda_pg_rca32_fa56_y3 = f_s_dadda_pg_rca32_fa56_y0 & f_s_dadda_pg_rca32_fa56_f_s_dadda_pg_rca32_and_10_5_y0;
  assign f_s_dadda_pg_rca32_fa56_y4 = f_s_dadda_pg_rca32_fa56_y1 | f_s_dadda_pg_rca32_fa56_y3;
  assign f_s_dadda_pg_rca32_and_9_6_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_9_6_y0 = f_s_dadda_pg_rca32_and_9_6_a_9 & f_s_dadda_pg_rca32_and_9_6_b_6;
  assign f_s_dadda_pg_rca32_and_8_7_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_8_7_y0 = f_s_dadda_pg_rca32_and_8_7_a_8 & f_s_dadda_pg_rca32_and_8_7_b_7;
  assign f_s_dadda_pg_rca32_and_7_8_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_7_8_y0 = f_s_dadda_pg_rca32_and_7_8_a_7 & f_s_dadda_pg_rca32_and_7_8_b_8;
  assign f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_9_6_y0 = f_s_dadda_pg_rca32_and_9_6_y0;
  assign f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_8_7_y0 = f_s_dadda_pg_rca32_and_8_7_y0;
  assign f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_7_8_y0 = f_s_dadda_pg_rca32_and_7_8_y0;
  assign f_s_dadda_pg_rca32_fa57_y0 = f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_9_6_y0 ^ f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_8_7_y0;
  assign f_s_dadda_pg_rca32_fa57_y1 = f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_9_6_y0 & f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_8_7_y0;
  assign f_s_dadda_pg_rca32_fa57_y2 = f_s_dadda_pg_rca32_fa57_y0 ^ f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_7_8_y0;
  assign f_s_dadda_pg_rca32_fa57_y3 = f_s_dadda_pg_rca32_fa57_y0 & f_s_dadda_pg_rca32_fa57_f_s_dadda_pg_rca32_and_7_8_y0;
  assign f_s_dadda_pg_rca32_fa57_y4 = f_s_dadda_pg_rca32_fa57_y1 | f_s_dadda_pg_rca32_fa57_y3;
  assign f_s_dadda_pg_rca32_and_6_9_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_6_9_y0 = f_s_dadda_pg_rca32_and_6_9_a_6 & f_s_dadda_pg_rca32_and_6_9_b_9;
  assign f_s_dadda_pg_rca32_and_5_10_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_5_10_y0 = f_s_dadda_pg_rca32_and_5_10_a_5 & f_s_dadda_pg_rca32_and_5_10_b_10;
  assign f_s_dadda_pg_rca32_and_4_11_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_4_11_y0 = f_s_dadda_pg_rca32_and_4_11_a_4 & f_s_dadda_pg_rca32_and_4_11_b_11;
  assign f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_6_9_y0 = f_s_dadda_pg_rca32_and_6_9_y0;
  assign f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_5_10_y0 = f_s_dadda_pg_rca32_and_5_10_y0;
  assign f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_4_11_y0 = f_s_dadda_pg_rca32_and_4_11_y0;
  assign f_s_dadda_pg_rca32_fa58_y0 = f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_6_9_y0 ^ f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_5_10_y0;
  assign f_s_dadda_pg_rca32_fa58_y1 = f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_6_9_y0 & f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_5_10_y0;
  assign f_s_dadda_pg_rca32_fa58_y2 = f_s_dadda_pg_rca32_fa58_y0 ^ f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_4_11_y0;
  assign f_s_dadda_pg_rca32_fa58_y3 = f_s_dadda_pg_rca32_fa58_y0 & f_s_dadda_pg_rca32_fa58_f_s_dadda_pg_rca32_and_4_11_y0;
  assign f_s_dadda_pg_rca32_fa58_y4 = f_s_dadda_pg_rca32_fa58_y1 | f_s_dadda_pg_rca32_fa58_y3;
  assign f_s_dadda_pg_rca32_and_3_12_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_3_12_y0 = f_s_dadda_pg_rca32_and_3_12_a_3 & f_s_dadda_pg_rca32_and_3_12_b_12;
  assign f_s_dadda_pg_rca32_and_2_13_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_2_13_y0 = f_s_dadda_pg_rca32_and_2_13_a_2 & f_s_dadda_pg_rca32_and_2_13_b_13;
  assign f_s_dadda_pg_rca32_and_1_14_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_1_14_y0 = f_s_dadda_pg_rca32_and_1_14_a_1 & f_s_dadda_pg_rca32_and_1_14_b_14;
  assign f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_3_12_y0 = f_s_dadda_pg_rca32_and_3_12_y0;
  assign f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_2_13_y0 = f_s_dadda_pg_rca32_and_2_13_y0;
  assign f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_1_14_y0 = f_s_dadda_pg_rca32_and_1_14_y0;
  assign f_s_dadda_pg_rca32_fa59_y0 = f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_3_12_y0 ^ f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_2_13_y0;
  assign f_s_dadda_pg_rca32_fa59_y1 = f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_3_12_y0 & f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_2_13_y0;
  assign f_s_dadda_pg_rca32_fa59_y2 = f_s_dadda_pg_rca32_fa59_y0 ^ f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_1_14_y0;
  assign f_s_dadda_pg_rca32_fa59_y3 = f_s_dadda_pg_rca32_fa59_y0 & f_s_dadda_pg_rca32_fa59_f_s_dadda_pg_rca32_and_1_14_y0;
  assign f_s_dadda_pg_rca32_fa59_y4 = f_s_dadda_pg_rca32_fa59_y1 | f_s_dadda_pg_rca32_fa59_y3;
  assign f_s_dadda_pg_rca32_and_0_15_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_0_15_y0 = f_s_dadda_pg_rca32_and_0_15_a_0 & f_s_dadda_pg_rca32_and_0_15_b_15;
  assign f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_and_0_15_y0 = f_s_dadda_pg_rca32_and_0_15_y0;
  assign f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_fa52_y2 = f_s_dadda_pg_rca32_fa52_y2;
  assign f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_fa53_y2 = f_s_dadda_pg_rca32_fa53_y2;
  assign f_s_dadda_pg_rca32_fa60_y0 = f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_and_0_15_y0 ^ f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_fa52_y2;
  assign f_s_dadda_pg_rca32_fa60_y1 = f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_and_0_15_y0 & f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_fa52_y2;
  assign f_s_dadda_pg_rca32_fa60_y2 = f_s_dadda_pg_rca32_fa60_y0 ^ f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_fa53_y2;
  assign f_s_dadda_pg_rca32_fa60_y3 = f_s_dadda_pg_rca32_fa60_y0 & f_s_dadda_pg_rca32_fa60_f_s_dadda_pg_rca32_fa53_y2;
  assign f_s_dadda_pg_rca32_fa60_y4 = f_s_dadda_pg_rca32_fa60_y1 | f_s_dadda_pg_rca32_fa60_y3;
  assign f_s_dadda_pg_rca32_ha13_f_s_dadda_pg_rca32_fa54_y2 = f_s_dadda_pg_rca32_fa54_y2;
  assign f_s_dadda_pg_rca32_ha13_f_s_dadda_pg_rca32_fa55_y2 = f_s_dadda_pg_rca32_fa55_y2;
  assign f_s_dadda_pg_rca32_ha13_y0 = f_s_dadda_pg_rca32_ha13_f_s_dadda_pg_rca32_fa54_y2 ^ f_s_dadda_pg_rca32_ha13_f_s_dadda_pg_rca32_fa55_y2;
  assign f_s_dadda_pg_rca32_ha13_y1 = f_s_dadda_pg_rca32_ha13_f_s_dadda_pg_rca32_fa54_y2 & f_s_dadda_pg_rca32_ha13_f_s_dadda_pg_rca32_fa55_y2;
  assign f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_ha13_y1 = f_s_dadda_pg_rca32_ha13_y1;
  assign f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_fa60_y4 = f_s_dadda_pg_rca32_fa60_y4;
  assign f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_fa59_y4 = f_s_dadda_pg_rca32_fa59_y4;
  assign f_s_dadda_pg_rca32_fa61_y0 = f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_ha13_y1 ^ f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_fa60_y4;
  assign f_s_dadda_pg_rca32_fa61_y1 = f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_ha13_y1 & f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_fa60_y4;
  assign f_s_dadda_pg_rca32_fa61_y2 = f_s_dadda_pg_rca32_fa61_y0 ^ f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_fa59_y4;
  assign f_s_dadda_pg_rca32_fa61_y3 = f_s_dadda_pg_rca32_fa61_y0 & f_s_dadda_pg_rca32_fa61_f_s_dadda_pg_rca32_fa59_y4;
  assign f_s_dadda_pg_rca32_fa61_y4 = f_s_dadda_pg_rca32_fa61_y1 | f_s_dadda_pg_rca32_fa61_y3;
  assign f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa58_y4 = f_s_dadda_pg_rca32_fa58_y4;
  assign f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa57_y4 = f_s_dadda_pg_rca32_fa57_y4;
  assign f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa56_y4 = f_s_dadda_pg_rca32_fa56_y4;
  assign f_s_dadda_pg_rca32_fa62_y0 = f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa58_y4 ^ f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa57_y4;
  assign f_s_dadda_pg_rca32_fa62_y1 = f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa58_y4 & f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa57_y4;
  assign f_s_dadda_pg_rca32_fa62_y2 = f_s_dadda_pg_rca32_fa62_y0 ^ f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa56_y4;
  assign f_s_dadda_pg_rca32_fa62_y3 = f_s_dadda_pg_rca32_fa62_y0 & f_s_dadda_pg_rca32_fa62_f_s_dadda_pg_rca32_fa56_y4;
  assign f_s_dadda_pg_rca32_fa62_y4 = f_s_dadda_pg_rca32_fa62_y1 | f_s_dadda_pg_rca32_fa62_y3;
  assign f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa55_y4 = f_s_dadda_pg_rca32_fa55_y4;
  assign f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa54_y4 = f_s_dadda_pg_rca32_fa54_y4;
  assign f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa53_y4 = f_s_dadda_pg_rca32_fa53_y4;
  assign f_s_dadda_pg_rca32_fa63_y0 = f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa55_y4 ^ f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa54_y4;
  assign f_s_dadda_pg_rca32_fa63_y1 = f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa55_y4 & f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa54_y4;
  assign f_s_dadda_pg_rca32_fa63_y2 = f_s_dadda_pg_rca32_fa63_y0 ^ f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa53_y4;
  assign f_s_dadda_pg_rca32_fa63_y3 = f_s_dadda_pg_rca32_fa63_y0 & f_s_dadda_pg_rca32_fa63_f_s_dadda_pg_rca32_fa53_y4;
  assign f_s_dadda_pg_rca32_fa63_y4 = f_s_dadda_pg_rca32_fa63_y1 | f_s_dadda_pg_rca32_fa63_y3;
  assign f_s_dadda_pg_rca32_and_16_0_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_16_0_y0 = f_s_dadda_pg_rca32_and_16_0_a_16 & f_s_dadda_pg_rca32_and_16_0_b_0;
  assign f_s_dadda_pg_rca32_and_15_1_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_15_1_y0 = f_s_dadda_pg_rca32_and_15_1_a_15 & f_s_dadda_pg_rca32_and_15_1_b_1;
  assign f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_fa52_y4 = f_s_dadda_pg_rca32_fa52_y4;
  assign f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_and_16_0_y0 = f_s_dadda_pg_rca32_and_16_0_y0;
  assign f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_and_15_1_y0 = f_s_dadda_pg_rca32_and_15_1_y0;
  assign f_s_dadda_pg_rca32_fa64_y0 = f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_fa52_y4 ^ f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_and_16_0_y0;
  assign f_s_dadda_pg_rca32_fa64_y1 = f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_fa52_y4 & f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_and_16_0_y0;
  assign f_s_dadda_pg_rca32_fa64_y2 = f_s_dadda_pg_rca32_fa64_y0 ^ f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_and_15_1_y0;
  assign f_s_dadda_pg_rca32_fa64_y3 = f_s_dadda_pg_rca32_fa64_y0 & f_s_dadda_pg_rca32_fa64_f_s_dadda_pg_rca32_and_15_1_y0;
  assign f_s_dadda_pg_rca32_fa64_y4 = f_s_dadda_pg_rca32_fa64_y1 | f_s_dadda_pg_rca32_fa64_y3;
  assign f_s_dadda_pg_rca32_and_14_2_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_14_2_y0 = f_s_dadda_pg_rca32_and_14_2_a_14 & f_s_dadda_pg_rca32_and_14_2_b_2;
  assign f_s_dadda_pg_rca32_and_13_3_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_13_3_y0 = f_s_dadda_pg_rca32_and_13_3_a_13 & f_s_dadda_pg_rca32_and_13_3_b_3;
  assign f_s_dadda_pg_rca32_and_12_4_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_12_4_y0 = f_s_dadda_pg_rca32_and_12_4_a_12 & f_s_dadda_pg_rca32_and_12_4_b_4;
  assign f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_14_2_y0 = f_s_dadda_pg_rca32_and_14_2_y0;
  assign f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_13_3_y0 = f_s_dadda_pg_rca32_and_13_3_y0;
  assign f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_12_4_y0 = f_s_dadda_pg_rca32_and_12_4_y0;
  assign f_s_dadda_pg_rca32_fa65_y0 = f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_14_2_y0 ^ f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_13_3_y0;
  assign f_s_dadda_pg_rca32_fa65_y1 = f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_14_2_y0 & f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_13_3_y0;
  assign f_s_dadda_pg_rca32_fa65_y2 = f_s_dadda_pg_rca32_fa65_y0 ^ f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_12_4_y0;
  assign f_s_dadda_pg_rca32_fa65_y3 = f_s_dadda_pg_rca32_fa65_y0 & f_s_dadda_pg_rca32_fa65_f_s_dadda_pg_rca32_and_12_4_y0;
  assign f_s_dadda_pg_rca32_fa65_y4 = f_s_dadda_pg_rca32_fa65_y1 | f_s_dadda_pg_rca32_fa65_y3;
  assign f_s_dadda_pg_rca32_and_11_5_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_11_5_y0 = f_s_dadda_pg_rca32_and_11_5_a_11 & f_s_dadda_pg_rca32_and_11_5_b_5;
  assign f_s_dadda_pg_rca32_and_10_6_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_10_6_y0 = f_s_dadda_pg_rca32_and_10_6_a_10 & f_s_dadda_pg_rca32_and_10_6_b_6;
  assign f_s_dadda_pg_rca32_and_9_7_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_9_7_y0 = f_s_dadda_pg_rca32_and_9_7_a_9 & f_s_dadda_pg_rca32_and_9_7_b_7;
  assign f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_11_5_y0 = f_s_dadda_pg_rca32_and_11_5_y0;
  assign f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_10_6_y0 = f_s_dadda_pg_rca32_and_10_6_y0;
  assign f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_9_7_y0 = f_s_dadda_pg_rca32_and_9_7_y0;
  assign f_s_dadda_pg_rca32_fa66_y0 = f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_11_5_y0 ^ f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_10_6_y0;
  assign f_s_dadda_pg_rca32_fa66_y1 = f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_11_5_y0 & f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_10_6_y0;
  assign f_s_dadda_pg_rca32_fa66_y2 = f_s_dadda_pg_rca32_fa66_y0 ^ f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_9_7_y0;
  assign f_s_dadda_pg_rca32_fa66_y3 = f_s_dadda_pg_rca32_fa66_y0 & f_s_dadda_pg_rca32_fa66_f_s_dadda_pg_rca32_and_9_7_y0;
  assign f_s_dadda_pg_rca32_fa66_y4 = f_s_dadda_pg_rca32_fa66_y1 | f_s_dadda_pg_rca32_fa66_y3;
  assign f_s_dadda_pg_rca32_and_8_8_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_8_8_y0 = f_s_dadda_pg_rca32_and_8_8_a_8 & f_s_dadda_pg_rca32_and_8_8_b_8;
  assign f_s_dadda_pg_rca32_and_7_9_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_7_9_y0 = f_s_dadda_pg_rca32_and_7_9_a_7 & f_s_dadda_pg_rca32_and_7_9_b_9;
  assign f_s_dadda_pg_rca32_and_6_10_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_6_10_y0 = f_s_dadda_pg_rca32_and_6_10_a_6 & f_s_dadda_pg_rca32_and_6_10_b_10;
  assign f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_8_8_y0 = f_s_dadda_pg_rca32_and_8_8_y0;
  assign f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_7_9_y0 = f_s_dadda_pg_rca32_and_7_9_y0;
  assign f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_6_10_y0 = f_s_dadda_pg_rca32_and_6_10_y0;
  assign f_s_dadda_pg_rca32_fa67_y0 = f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_8_8_y0 ^ f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_7_9_y0;
  assign f_s_dadda_pg_rca32_fa67_y1 = f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_8_8_y0 & f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_7_9_y0;
  assign f_s_dadda_pg_rca32_fa67_y2 = f_s_dadda_pg_rca32_fa67_y0 ^ f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_6_10_y0;
  assign f_s_dadda_pg_rca32_fa67_y3 = f_s_dadda_pg_rca32_fa67_y0 & f_s_dadda_pg_rca32_fa67_f_s_dadda_pg_rca32_and_6_10_y0;
  assign f_s_dadda_pg_rca32_fa67_y4 = f_s_dadda_pg_rca32_fa67_y1 | f_s_dadda_pg_rca32_fa67_y3;
  assign f_s_dadda_pg_rca32_and_5_11_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_5_11_y0 = f_s_dadda_pg_rca32_and_5_11_a_5 & f_s_dadda_pg_rca32_and_5_11_b_11;
  assign f_s_dadda_pg_rca32_and_4_12_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_4_12_y0 = f_s_dadda_pg_rca32_and_4_12_a_4 & f_s_dadda_pg_rca32_and_4_12_b_12;
  assign f_s_dadda_pg_rca32_and_3_13_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_3_13_y0 = f_s_dadda_pg_rca32_and_3_13_a_3 & f_s_dadda_pg_rca32_and_3_13_b_13;
  assign f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_5_11_y0 = f_s_dadda_pg_rca32_and_5_11_y0;
  assign f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_4_12_y0 = f_s_dadda_pg_rca32_and_4_12_y0;
  assign f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_3_13_y0 = f_s_dadda_pg_rca32_and_3_13_y0;
  assign f_s_dadda_pg_rca32_fa68_y0 = f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_5_11_y0 ^ f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_4_12_y0;
  assign f_s_dadda_pg_rca32_fa68_y1 = f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_5_11_y0 & f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_4_12_y0;
  assign f_s_dadda_pg_rca32_fa68_y2 = f_s_dadda_pg_rca32_fa68_y0 ^ f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_3_13_y0;
  assign f_s_dadda_pg_rca32_fa68_y3 = f_s_dadda_pg_rca32_fa68_y0 & f_s_dadda_pg_rca32_fa68_f_s_dadda_pg_rca32_and_3_13_y0;
  assign f_s_dadda_pg_rca32_fa68_y4 = f_s_dadda_pg_rca32_fa68_y1 | f_s_dadda_pg_rca32_fa68_y3;
  assign f_s_dadda_pg_rca32_and_2_14_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_2_14_y0 = f_s_dadda_pg_rca32_and_2_14_a_2 & f_s_dadda_pg_rca32_and_2_14_b_14;
  assign f_s_dadda_pg_rca32_and_1_15_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_1_15_y0 = f_s_dadda_pg_rca32_and_1_15_a_1 & f_s_dadda_pg_rca32_and_1_15_b_15;
  assign f_s_dadda_pg_rca32_and_0_16_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_0_16_y0 = f_s_dadda_pg_rca32_and_0_16_a_0 & f_s_dadda_pg_rca32_and_0_16_b_16;
  assign f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_2_14_y0 = f_s_dadda_pg_rca32_and_2_14_y0;
  assign f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_1_15_y0 = f_s_dadda_pg_rca32_and_1_15_y0;
  assign f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_0_16_y0 = f_s_dadda_pg_rca32_and_0_16_y0;
  assign f_s_dadda_pg_rca32_fa69_y0 = f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_2_14_y0 ^ f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_1_15_y0;
  assign f_s_dadda_pg_rca32_fa69_y1 = f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_2_14_y0 & f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_1_15_y0;
  assign f_s_dadda_pg_rca32_fa69_y2 = f_s_dadda_pg_rca32_fa69_y0 ^ f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_0_16_y0;
  assign f_s_dadda_pg_rca32_fa69_y3 = f_s_dadda_pg_rca32_fa69_y0 & f_s_dadda_pg_rca32_fa69_f_s_dadda_pg_rca32_and_0_16_y0;
  assign f_s_dadda_pg_rca32_fa69_y4 = f_s_dadda_pg_rca32_fa69_y1 | f_s_dadda_pg_rca32_fa69_y3;
  assign f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa61_y2 = f_s_dadda_pg_rca32_fa61_y2;
  assign f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa62_y2 = f_s_dadda_pg_rca32_fa62_y2;
  assign f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa63_y2 = f_s_dadda_pg_rca32_fa63_y2;
  assign f_s_dadda_pg_rca32_fa70_y0 = f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa61_y2 ^ f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa62_y2;
  assign f_s_dadda_pg_rca32_fa70_y1 = f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa61_y2 & f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa62_y2;
  assign f_s_dadda_pg_rca32_fa70_y2 = f_s_dadda_pg_rca32_fa70_y0 ^ f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa63_y2;
  assign f_s_dadda_pg_rca32_fa70_y3 = f_s_dadda_pg_rca32_fa70_y0 & f_s_dadda_pg_rca32_fa70_f_s_dadda_pg_rca32_fa63_y2;
  assign f_s_dadda_pg_rca32_fa70_y4 = f_s_dadda_pg_rca32_fa70_y1 | f_s_dadda_pg_rca32_fa70_y3;
  assign f_s_dadda_pg_rca32_ha14_f_s_dadda_pg_rca32_fa64_y2 = f_s_dadda_pg_rca32_fa64_y2;
  assign f_s_dadda_pg_rca32_ha14_f_s_dadda_pg_rca32_fa65_y2 = f_s_dadda_pg_rca32_fa65_y2;
  assign f_s_dadda_pg_rca32_ha14_y0 = f_s_dadda_pg_rca32_ha14_f_s_dadda_pg_rca32_fa64_y2 ^ f_s_dadda_pg_rca32_ha14_f_s_dadda_pg_rca32_fa65_y2;
  assign f_s_dadda_pg_rca32_ha14_y1 = f_s_dadda_pg_rca32_ha14_f_s_dadda_pg_rca32_fa64_y2 & f_s_dadda_pg_rca32_ha14_f_s_dadda_pg_rca32_fa65_y2;
  assign f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_ha14_y1 = f_s_dadda_pg_rca32_ha14_y1;
  assign f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_fa70_y4 = f_s_dadda_pg_rca32_fa70_y4;
  assign f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_fa69_y4 = f_s_dadda_pg_rca32_fa69_y4;
  assign f_s_dadda_pg_rca32_fa71_y0 = f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_ha14_y1 ^ f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_fa70_y4;
  assign f_s_dadda_pg_rca32_fa71_y1 = f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_ha14_y1 & f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_fa70_y4;
  assign f_s_dadda_pg_rca32_fa71_y2 = f_s_dadda_pg_rca32_fa71_y0 ^ f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_fa69_y4;
  assign f_s_dadda_pg_rca32_fa71_y3 = f_s_dadda_pg_rca32_fa71_y0 & f_s_dadda_pg_rca32_fa71_f_s_dadda_pg_rca32_fa69_y4;
  assign f_s_dadda_pg_rca32_fa71_y4 = f_s_dadda_pg_rca32_fa71_y1 | f_s_dadda_pg_rca32_fa71_y3;
  assign f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa68_y4 = f_s_dadda_pg_rca32_fa68_y4;
  assign f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa67_y4 = f_s_dadda_pg_rca32_fa67_y4;
  assign f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa66_y4 = f_s_dadda_pg_rca32_fa66_y4;
  assign f_s_dadda_pg_rca32_fa72_y0 = f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa68_y4 ^ f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa67_y4;
  assign f_s_dadda_pg_rca32_fa72_y1 = f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa68_y4 & f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa67_y4;
  assign f_s_dadda_pg_rca32_fa72_y2 = f_s_dadda_pg_rca32_fa72_y0 ^ f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa66_y4;
  assign f_s_dadda_pg_rca32_fa72_y3 = f_s_dadda_pg_rca32_fa72_y0 & f_s_dadda_pg_rca32_fa72_f_s_dadda_pg_rca32_fa66_y4;
  assign f_s_dadda_pg_rca32_fa72_y4 = f_s_dadda_pg_rca32_fa72_y1 | f_s_dadda_pg_rca32_fa72_y3;
  assign f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa65_y4 = f_s_dadda_pg_rca32_fa65_y4;
  assign f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa64_y4 = f_s_dadda_pg_rca32_fa64_y4;
  assign f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa63_y4 = f_s_dadda_pg_rca32_fa63_y4;
  assign f_s_dadda_pg_rca32_fa73_y0 = f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa65_y4 ^ f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa64_y4;
  assign f_s_dadda_pg_rca32_fa73_y1 = f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa65_y4 & f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa64_y4;
  assign f_s_dadda_pg_rca32_fa73_y2 = f_s_dadda_pg_rca32_fa73_y0 ^ f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa63_y4;
  assign f_s_dadda_pg_rca32_fa73_y3 = f_s_dadda_pg_rca32_fa73_y0 & f_s_dadda_pg_rca32_fa73_f_s_dadda_pg_rca32_fa63_y4;
  assign f_s_dadda_pg_rca32_fa73_y4 = f_s_dadda_pg_rca32_fa73_y1 | f_s_dadda_pg_rca32_fa73_y3;
  assign f_s_dadda_pg_rca32_and_17_0_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_17_0_y0 = f_s_dadda_pg_rca32_and_17_0_a_17 & f_s_dadda_pg_rca32_and_17_0_b_0;
  assign f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_fa62_y4 = f_s_dadda_pg_rca32_fa62_y4;
  assign f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_fa61_y4 = f_s_dadda_pg_rca32_fa61_y4;
  assign f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_and_17_0_y0 = f_s_dadda_pg_rca32_and_17_0_y0;
  assign f_s_dadda_pg_rca32_fa74_y0 = f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_fa62_y4 ^ f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_fa61_y4;
  assign f_s_dadda_pg_rca32_fa74_y1 = f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_fa62_y4 & f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_fa61_y4;
  assign f_s_dadda_pg_rca32_fa74_y2 = f_s_dadda_pg_rca32_fa74_y0 ^ f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_and_17_0_y0;
  assign f_s_dadda_pg_rca32_fa74_y3 = f_s_dadda_pg_rca32_fa74_y0 & f_s_dadda_pg_rca32_fa74_f_s_dadda_pg_rca32_and_17_0_y0;
  assign f_s_dadda_pg_rca32_fa74_y4 = f_s_dadda_pg_rca32_fa74_y1 | f_s_dadda_pg_rca32_fa74_y3;
  assign f_s_dadda_pg_rca32_and_16_1_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_16_1_y0 = f_s_dadda_pg_rca32_and_16_1_a_16 & f_s_dadda_pg_rca32_and_16_1_b_1;
  assign f_s_dadda_pg_rca32_and_15_2_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_15_2_y0 = f_s_dadda_pg_rca32_and_15_2_a_15 & f_s_dadda_pg_rca32_and_15_2_b_2;
  assign f_s_dadda_pg_rca32_and_14_3_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_14_3_y0 = f_s_dadda_pg_rca32_and_14_3_a_14 & f_s_dadda_pg_rca32_and_14_3_b_3;
  assign f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_16_1_y0 = f_s_dadda_pg_rca32_and_16_1_y0;
  assign f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_15_2_y0 = f_s_dadda_pg_rca32_and_15_2_y0;
  assign f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_14_3_y0 = f_s_dadda_pg_rca32_and_14_3_y0;
  assign f_s_dadda_pg_rca32_fa75_y0 = f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_16_1_y0 ^ f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_15_2_y0;
  assign f_s_dadda_pg_rca32_fa75_y1 = f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_16_1_y0 & f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_15_2_y0;
  assign f_s_dadda_pg_rca32_fa75_y2 = f_s_dadda_pg_rca32_fa75_y0 ^ f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_14_3_y0;
  assign f_s_dadda_pg_rca32_fa75_y3 = f_s_dadda_pg_rca32_fa75_y0 & f_s_dadda_pg_rca32_fa75_f_s_dadda_pg_rca32_and_14_3_y0;
  assign f_s_dadda_pg_rca32_fa75_y4 = f_s_dadda_pg_rca32_fa75_y1 | f_s_dadda_pg_rca32_fa75_y3;
  assign f_s_dadda_pg_rca32_and_13_4_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_13_4_y0 = f_s_dadda_pg_rca32_and_13_4_a_13 & f_s_dadda_pg_rca32_and_13_4_b_4;
  assign f_s_dadda_pg_rca32_and_12_5_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_12_5_y0 = f_s_dadda_pg_rca32_and_12_5_a_12 & f_s_dadda_pg_rca32_and_12_5_b_5;
  assign f_s_dadda_pg_rca32_and_11_6_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_11_6_y0 = f_s_dadda_pg_rca32_and_11_6_a_11 & f_s_dadda_pg_rca32_and_11_6_b_6;
  assign f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_13_4_y0 = f_s_dadda_pg_rca32_and_13_4_y0;
  assign f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_12_5_y0 = f_s_dadda_pg_rca32_and_12_5_y0;
  assign f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_11_6_y0 = f_s_dadda_pg_rca32_and_11_6_y0;
  assign f_s_dadda_pg_rca32_fa76_y0 = f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_13_4_y0 ^ f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_12_5_y0;
  assign f_s_dadda_pg_rca32_fa76_y1 = f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_13_4_y0 & f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_12_5_y0;
  assign f_s_dadda_pg_rca32_fa76_y2 = f_s_dadda_pg_rca32_fa76_y0 ^ f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_11_6_y0;
  assign f_s_dadda_pg_rca32_fa76_y3 = f_s_dadda_pg_rca32_fa76_y0 & f_s_dadda_pg_rca32_fa76_f_s_dadda_pg_rca32_and_11_6_y0;
  assign f_s_dadda_pg_rca32_fa76_y4 = f_s_dadda_pg_rca32_fa76_y1 | f_s_dadda_pg_rca32_fa76_y3;
  assign f_s_dadda_pg_rca32_and_10_7_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_10_7_y0 = f_s_dadda_pg_rca32_and_10_7_a_10 & f_s_dadda_pg_rca32_and_10_7_b_7;
  assign f_s_dadda_pg_rca32_and_9_8_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_9_8_y0 = f_s_dadda_pg_rca32_and_9_8_a_9 & f_s_dadda_pg_rca32_and_9_8_b_8;
  assign f_s_dadda_pg_rca32_and_8_9_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_8_9_y0 = f_s_dadda_pg_rca32_and_8_9_a_8 & f_s_dadda_pg_rca32_and_8_9_b_9;
  assign f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_10_7_y0 = f_s_dadda_pg_rca32_and_10_7_y0;
  assign f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_9_8_y0 = f_s_dadda_pg_rca32_and_9_8_y0;
  assign f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_8_9_y0 = f_s_dadda_pg_rca32_and_8_9_y0;
  assign f_s_dadda_pg_rca32_fa77_y0 = f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_10_7_y0 ^ f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_9_8_y0;
  assign f_s_dadda_pg_rca32_fa77_y1 = f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_10_7_y0 & f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_9_8_y0;
  assign f_s_dadda_pg_rca32_fa77_y2 = f_s_dadda_pg_rca32_fa77_y0 ^ f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_8_9_y0;
  assign f_s_dadda_pg_rca32_fa77_y3 = f_s_dadda_pg_rca32_fa77_y0 & f_s_dadda_pg_rca32_fa77_f_s_dadda_pg_rca32_and_8_9_y0;
  assign f_s_dadda_pg_rca32_fa77_y4 = f_s_dadda_pg_rca32_fa77_y1 | f_s_dadda_pg_rca32_fa77_y3;
  assign f_s_dadda_pg_rca32_and_7_10_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_7_10_y0 = f_s_dadda_pg_rca32_and_7_10_a_7 & f_s_dadda_pg_rca32_and_7_10_b_10;
  assign f_s_dadda_pg_rca32_and_6_11_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_6_11_y0 = f_s_dadda_pg_rca32_and_6_11_a_6 & f_s_dadda_pg_rca32_and_6_11_b_11;
  assign f_s_dadda_pg_rca32_and_5_12_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_5_12_y0 = f_s_dadda_pg_rca32_and_5_12_a_5 & f_s_dadda_pg_rca32_and_5_12_b_12;
  assign f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_7_10_y0 = f_s_dadda_pg_rca32_and_7_10_y0;
  assign f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_6_11_y0 = f_s_dadda_pg_rca32_and_6_11_y0;
  assign f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_5_12_y0 = f_s_dadda_pg_rca32_and_5_12_y0;
  assign f_s_dadda_pg_rca32_fa78_y0 = f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_7_10_y0 ^ f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_6_11_y0;
  assign f_s_dadda_pg_rca32_fa78_y1 = f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_7_10_y0 & f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_6_11_y0;
  assign f_s_dadda_pg_rca32_fa78_y2 = f_s_dadda_pg_rca32_fa78_y0 ^ f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_5_12_y0;
  assign f_s_dadda_pg_rca32_fa78_y3 = f_s_dadda_pg_rca32_fa78_y0 & f_s_dadda_pg_rca32_fa78_f_s_dadda_pg_rca32_and_5_12_y0;
  assign f_s_dadda_pg_rca32_fa78_y4 = f_s_dadda_pg_rca32_fa78_y1 | f_s_dadda_pg_rca32_fa78_y3;
  assign f_s_dadda_pg_rca32_and_4_13_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_4_13_y0 = f_s_dadda_pg_rca32_and_4_13_a_4 & f_s_dadda_pg_rca32_and_4_13_b_13;
  assign f_s_dadda_pg_rca32_and_3_14_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_3_14_y0 = f_s_dadda_pg_rca32_and_3_14_a_3 & f_s_dadda_pg_rca32_and_3_14_b_14;
  assign f_s_dadda_pg_rca32_and_2_15_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_2_15_y0 = f_s_dadda_pg_rca32_and_2_15_a_2 & f_s_dadda_pg_rca32_and_2_15_b_15;
  assign f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_4_13_y0 = f_s_dadda_pg_rca32_and_4_13_y0;
  assign f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_3_14_y0 = f_s_dadda_pg_rca32_and_3_14_y0;
  assign f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_2_15_y0 = f_s_dadda_pg_rca32_and_2_15_y0;
  assign f_s_dadda_pg_rca32_fa79_y0 = f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_4_13_y0 ^ f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_3_14_y0;
  assign f_s_dadda_pg_rca32_fa79_y1 = f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_4_13_y0 & f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_3_14_y0;
  assign f_s_dadda_pg_rca32_fa79_y2 = f_s_dadda_pg_rca32_fa79_y0 ^ f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_2_15_y0;
  assign f_s_dadda_pg_rca32_fa79_y3 = f_s_dadda_pg_rca32_fa79_y0 & f_s_dadda_pg_rca32_fa79_f_s_dadda_pg_rca32_and_2_15_y0;
  assign f_s_dadda_pg_rca32_fa79_y4 = f_s_dadda_pg_rca32_fa79_y1 | f_s_dadda_pg_rca32_fa79_y3;
  assign f_s_dadda_pg_rca32_and_1_16_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_1_16_y0 = f_s_dadda_pg_rca32_and_1_16_a_1 & f_s_dadda_pg_rca32_and_1_16_b_16;
  assign f_s_dadda_pg_rca32_and_0_17_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_0_17_y0 = f_s_dadda_pg_rca32_and_0_17_a_0 & f_s_dadda_pg_rca32_and_0_17_b_17;
  assign f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_and_1_16_y0 = f_s_dadda_pg_rca32_and_1_16_y0;
  assign f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_and_0_17_y0 = f_s_dadda_pg_rca32_and_0_17_y0;
  assign f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_fa71_y2 = f_s_dadda_pg_rca32_fa71_y2;
  assign f_s_dadda_pg_rca32_fa80_y0 = f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_and_1_16_y0 ^ f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_and_0_17_y0;
  assign f_s_dadda_pg_rca32_fa80_y1 = f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_and_1_16_y0 & f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_and_0_17_y0;
  assign f_s_dadda_pg_rca32_fa80_y2 = f_s_dadda_pg_rca32_fa80_y0 ^ f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_fa71_y2;
  assign f_s_dadda_pg_rca32_fa80_y3 = f_s_dadda_pg_rca32_fa80_y0 & f_s_dadda_pg_rca32_fa80_f_s_dadda_pg_rca32_fa71_y2;
  assign f_s_dadda_pg_rca32_fa80_y4 = f_s_dadda_pg_rca32_fa80_y1 | f_s_dadda_pg_rca32_fa80_y3;
  assign f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa72_y2 = f_s_dadda_pg_rca32_fa72_y2;
  assign f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa73_y2 = f_s_dadda_pg_rca32_fa73_y2;
  assign f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa74_y2 = f_s_dadda_pg_rca32_fa74_y2;
  assign f_s_dadda_pg_rca32_fa81_y0 = f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa72_y2 ^ f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa73_y2;
  assign f_s_dadda_pg_rca32_fa81_y1 = f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa72_y2 & f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa73_y2;
  assign f_s_dadda_pg_rca32_fa81_y2 = f_s_dadda_pg_rca32_fa81_y0 ^ f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa74_y2;
  assign f_s_dadda_pg_rca32_fa81_y3 = f_s_dadda_pg_rca32_fa81_y0 & f_s_dadda_pg_rca32_fa81_f_s_dadda_pg_rca32_fa74_y2;
  assign f_s_dadda_pg_rca32_fa81_y4 = f_s_dadda_pg_rca32_fa81_y1 | f_s_dadda_pg_rca32_fa81_y3;
  assign f_s_dadda_pg_rca32_ha15_f_s_dadda_pg_rca32_fa75_y2 = f_s_dadda_pg_rca32_fa75_y2;
  assign f_s_dadda_pg_rca32_ha15_f_s_dadda_pg_rca32_fa76_y2 = f_s_dadda_pg_rca32_fa76_y2;
  assign f_s_dadda_pg_rca32_ha15_y0 = f_s_dadda_pg_rca32_ha15_f_s_dadda_pg_rca32_fa75_y2 ^ f_s_dadda_pg_rca32_ha15_f_s_dadda_pg_rca32_fa76_y2;
  assign f_s_dadda_pg_rca32_ha15_y1 = f_s_dadda_pg_rca32_ha15_f_s_dadda_pg_rca32_fa75_y2 & f_s_dadda_pg_rca32_ha15_f_s_dadda_pg_rca32_fa76_y2;
  assign f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_ha15_y1 = f_s_dadda_pg_rca32_ha15_y1;
  assign f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_fa81_y4 = f_s_dadda_pg_rca32_fa81_y4;
  assign f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_fa80_y4 = f_s_dadda_pg_rca32_fa80_y4;
  assign f_s_dadda_pg_rca32_fa82_y0 = f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_ha15_y1 ^ f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_fa81_y4;
  assign f_s_dadda_pg_rca32_fa82_y1 = f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_ha15_y1 & f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_fa81_y4;
  assign f_s_dadda_pg_rca32_fa82_y2 = f_s_dadda_pg_rca32_fa82_y0 ^ f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_fa80_y4;
  assign f_s_dadda_pg_rca32_fa82_y3 = f_s_dadda_pg_rca32_fa82_y0 & f_s_dadda_pg_rca32_fa82_f_s_dadda_pg_rca32_fa80_y4;
  assign f_s_dadda_pg_rca32_fa82_y4 = f_s_dadda_pg_rca32_fa82_y1 | f_s_dadda_pg_rca32_fa82_y3;
  assign f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa79_y4 = f_s_dadda_pg_rca32_fa79_y4;
  assign f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa78_y4 = f_s_dadda_pg_rca32_fa78_y4;
  assign f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa77_y4 = f_s_dadda_pg_rca32_fa77_y4;
  assign f_s_dadda_pg_rca32_fa83_y0 = f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa79_y4 ^ f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa78_y4;
  assign f_s_dadda_pg_rca32_fa83_y1 = f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa79_y4 & f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa78_y4;
  assign f_s_dadda_pg_rca32_fa83_y2 = f_s_dadda_pg_rca32_fa83_y0 ^ f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa77_y4;
  assign f_s_dadda_pg_rca32_fa83_y3 = f_s_dadda_pg_rca32_fa83_y0 & f_s_dadda_pg_rca32_fa83_f_s_dadda_pg_rca32_fa77_y4;
  assign f_s_dadda_pg_rca32_fa83_y4 = f_s_dadda_pg_rca32_fa83_y1 | f_s_dadda_pg_rca32_fa83_y3;
  assign f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa76_y4 = f_s_dadda_pg_rca32_fa76_y4;
  assign f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa75_y4 = f_s_dadda_pg_rca32_fa75_y4;
  assign f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa74_y4 = f_s_dadda_pg_rca32_fa74_y4;
  assign f_s_dadda_pg_rca32_fa84_y0 = f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa76_y4 ^ f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa75_y4;
  assign f_s_dadda_pg_rca32_fa84_y1 = f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa76_y4 & f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa75_y4;
  assign f_s_dadda_pg_rca32_fa84_y2 = f_s_dadda_pg_rca32_fa84_y0 ^ f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa74_y4;
  assign f_s_dadda_pg_rca32_fa84_y3 = f_s_dadda_pg_rca32_fa84_y0 & f_s_dadda_pg_rca32_fa84_f_s_dadda_pg_rca32_fa74_y4;
  assign f_s_dadda_pg_rca32_fa84_y4 = f_s_dadda_pg_rca32_fa84_y1 | f_s_dadda_pg_rca32_fa84_y3;
  assign f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa73_y4 = f_s_dadda_pg_rca32_fa73_y4;
  assign f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa72_y4 = f_s_dadda_pg_rca32_fa72_y4;
  assign f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa71_y4 = f_s_dadda_pg_rca32_fa71_y4;
  assign f_s_dadda_pg_rca32_fa85_y0 = f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa73_y4 ^ f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa72_y4;
  assign f_s_dadda_pg_rca32_fa85_y1 = f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa73_y4 & f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa72_y4;
  assign f_s_dadda_pg_rca32_fa85_y2 = f_s_dadda_pg_rca32_fa85_y0 ^ f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa71_y4;
  assign f_s_dadda_pg_rca32_fa85_y3 = f_s_dadda_pg_rca32_fa85_y0 & f_s_dadda_pg_rca32_fa85_f_s_dadda_pg_rca32_fa71_y4;
  assign f_s_dadda_pg_rca32_fa85_y4 = f_s_dadda_pg_rca32_fa85_y1 | f_s_dadda_pg_rca32_fa85_y3;
  assign f_s_dadda_pg_rca32_and_18_0_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_18_0_y0 = f_s_dadda_pg_rca32_and_18_0_a_18 & f_s_dadda_pg_rca32_and_18_0_b_0;
  assign f_s_dadda_pg_rca32_and_17_1_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_17_1_y0 = f_s_dadda_pg_rca32_and_17_1_a_17 & f_s_dadda_pg_rca32_and_17_1_b_1;
  assign f_s_dadda_pg_rca32_and_16_2_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_16_2_y0 = f_s_dadda_pg_rca32_and_16_2_a_16 & f_s_dadda_pg_rca32_and_16_2_b_2;
  assign f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_18_0_y0 = f_s_dadda_pg_rca32_and_18_0_y0;
  assign f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_17_1_y0 = f_s_dadda_pg_rca32_and_17_1_y0;
  assign f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_16_2_y0 = f_s_dadda_pg_rca32_and_16_2_y0;
  assign f_s_dadda_pg_rca32_fa86_y0 = f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_18_0_y0 ^ f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_17_1_y0;
  assign f_s_dadda_pg_rca32_fa86_y1 = f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_18_0_y0 & f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_17_1_y0;
  assign f_s_dadda_pg_rca32_fa86_y2 = f_s_dadda_pg_rca32_fa86_y0 ^ f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_16_2_y0;
  assign f_s_dadda_pg_rca32_fa86_y3 = f_s_dadda_pg_rca32_fa86_y0 & f_s_dadda_pg_rca32_fa86_f_s_dadda_pg_rca32_and_16_2_y0;
  assign f_s_dadda_pg_rca32_fa86_y4 = f_s_dadda_pg_rca32_fa86_y1 | f_s_dadda_pg_rca32_fa86_y3;
  assign f_s_dadda_pg_rca32_and_15_3_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_15_3_y0 = f_s_dadda_pg_rca32_and_15_3_a_15 & f_s_dadda_pg_rca32_and_15_3_b_3;
  assign f_s_dadda_pg_rca32_and_14_4_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_14_4_y0 = f_s_dadda_pg_rca32_and_14_4_a_14 & f_s_dadda_pg_rca32_and_14_4_b_4;
  assign f_s_dadda_pg_rca32_and_13_5_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_13_5_y0 = f_s_dadda_pg_rca32_and_13_5_a_13 & f_s_dadda_pg_rca32_and_13_5_b_5;
  assign f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_15_3_y0 = f_s_dadda_pg_rca32_and_15_3_y0;
  assign f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_14_4_y0 = f_s_dadda_pg_rca32_and_14_4_y0;
  assign f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_13_5_y0 = f_s_dadda_pg_rca32_and_13_5_y0;
  assign f_s_dadda_pg_rca32_fa87_y0 = f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_15_3_y0 ^ f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_14_4_y0;
  assign f_s_dadda_pg_rca32_fa87_y1 = f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_15_3_y0 & f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_14_4_y0;
  assign f_s_dadda_pg_rca32_fa87_y2 = f_s_dadda_pg_rca32_fa87_y0 ^ f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_13_5_y0;
  assign f_s_dadda_pg_rca32_fa87_y3 = f_s_dadda_pg_rca32_fa87_y0 & f_s_dadda_pg_rca32_fa87_f_s_dadda_pg_rca32_and_13_5_y0;
  assign f_s_dadda_pg_rca32_fa87_y4 = f_s_dadda_pg_rca32_fa87_y1 | f_s_dadda_pg_rca32_fa87_y3;
  assign f_s_dadda_pg_rca32_and_12_6_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_12_6_y0 = f_s_dadda_pg_rca32_and_12_6_a_12 & f_s_dadda_pg_rca32_and_12_6_b_6;
  assign f_s_dadda_pg_rca32_and_11_7_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_11_7_y0 = f_s_dadda_pg_rca32_and_11_7_a_11 & f_s_dadda_pg_rca32_and_11_7_b_7;
  assign f_s_dadda_pg_rca32_and_10_8_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_10_8_y0 = f_s_dadda_pg_rca32_and_10_8_a_10 & f_s_dadda_pg_rca32_and_10_8_b_8;
  assign f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_12_6_y0 = f_s_dadda_pg_rca32_and_12_6_y0;
  assign f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_11_7_y0 = f_s_dadda_pg_rca32_and_11_7_y0;
  assign f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_10_8_y0 = f_s_dadda_pg_rca32_and_10_8_y0;
  assign f_s_dadda_pg_rca32_fa88_y0 = f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_12_6_y0 ^ f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_11_7_y0;
  assign f_s_dadda_pg_rca32_fa88_y1 = f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_12_6_y0 & f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_11_7_y0;
  assign f_s_dadda_pg_rca32_fa88_y2 = f_s_dadda_pg_rca32_fa88_y0 ^ f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_10_8_y0;
  assign f_s_dadda_pg_rca32_fa88_y3 = f_s_dadda_pg_rca32_fa88_y0 & f_s_dadda_pg_rca32_fa88_f_s_dadda_pg_rca32_and_10_8_y0;
  assign f_s_dadda_pg_rca32_fa88_y4 = f_s_dadda_pg_rca32_fa88_y1 | f_s_dadda_pg_rca32_fa88_y3;
  assign f_s_dadda_pg_rca32_and_9_9_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_9_9_y0 = f_s_dadda_pg_rca32_and_9_9_a_9 & f_s_dadda_pg_rca32_and_9_9_b_9;
  assign f_s_dadda_pg_rca32_and_8_10_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_8_10_y0 = f_s_dadda_pg_rca32_and_8_10_a_8 & f_s_dadda_pg_rca32_and_8_10_b_10;
  assign f_s_dadda_pg_rca32_and_7_11_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_7_11_y0 = f_s_dadda_pg_rca32_and_7_11_a_7 & f_s_dadda_pg_rca32_and_7_11_b_11;
  assign f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_9_9_y0 = f_s_dadda_pg_rca32_and_9_9_y0;
  assign f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_8_10_y0 = f_s_dadda_pg_rca32_and_8_10_y0;
  assign f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_7_11_y0 = f_s_dadda_pg_rca32_and_7_11_y0;
  assign f_s_dadda_pg_rca32_fa89_y0 = f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_9_9_y0 ^ f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_8_10_y0;
  assign f_s_dadda_pg_rca32_fa89_y1 = f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_9_9_y0 & f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_8_10_y0;
  assign f_s_dadda_pg_rca32_fa89_y2 = f_s_dadda_pg_rca32_fa89_y0 ^ f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_7_11_y0;
  assign f_s_dadda_pg_rca32_fa89_y3 = f_s_dadda_pg_rca32_fa89_y0 & f_s_dadda_pg_rca32_fa89_f_s_dadda_pg_rca32_and_7_11_y0;
  assign f_s_dadda_pg_rca32_fa89_y4 = f_s_dadda_pg_rca32_fa89_y1 | f_s_dadda_pg_rca32_fa89_y3;
  assign f_s_dadda_pg_rca32_and_6_12_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_6_12_y0 = f_s_dadda_pg_rca32_and_6_12_a_6 & f_s_dadda_pg_rca32_and_6_12_b_12;
  assign f_s_dadda_pg_rca32_and_5_13_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_5_13_y0 = f_s_dadda_pg_rca32_and_5_13_a_5 & f_s_dadda_pg_rca32_and_5_13_b_13;
  assign f_s_dadda_pg_rca32_and_4_14_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_4_14_y0 = f_s_dadda_pg_rca32_and_4_14_a_4 & f_s_dadda_pg_rca32_and_4_14_b_14;
  assign f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_6_12_y0 = f_s_dadda_pg_rca32_and_6_12_y0;
  assign f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_5_13_y0 = f_s_dadda_pg_rca32_and_5_13_y0;
  assign f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_4_14_y0 = f_s_dadda_pg_rca32_and_4_14_y0;
  assign f_s_dadda_pg_rca32_fa90_y0 = f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_6_12_y0 ^ f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_5_13_y0;
  assign f_s_dadda_pg_rca32_fa90_y1 = f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_6_12_y0 & f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_5_13_y0;
  assign f_s_dadda_pg_rca32_fa90_y2 = f_s_dadda_pg_rca32_fa90_y0 ^ f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_4_14_y0;
  assign f_s_dadda_pg_rca32_fa90_y3 = f_s_dadda_pg_rca32_fa90_y0 & f_s_dadda_pg_rca32_fa90_f_s_dadda_pg_rca32_and_4_14_y0;
  assign f_s_dadda_pg_rca32_fa90_y4 = f_s_dadda_pg_rca32_fa90_y1 | f_s_dadda_pg_rca32_fa90_y3;
  assign f_s_dadda_pg_rca32_and_3_15_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_3_15_y0 = f_s_dadda_pg_rca32_and_3_15_a_3 & f_s_dadda_pg_rca32_and_3_15_b_15;
  assign f_s_dadda_pg_rca32_and_2_16_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_2_16_y0 = f_s_dadda_pg_rca32_and_2_16_a_2 & f_s_dadda_pg_rca32_and_2_16_b_16;
  assign f_s_dadda_pg_rca32_and_1_17_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_1_17_y0 = f_s_dadda_pg_rca32_and_1_17_a_1 & f_s_dadda_pg_rca32_and_1_17_b_17;
  assign f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_3_15_y0 = f_s_dadda_pg_rca32_and_3_15_y0;
  assign f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_2_16_y0 = f_s_dadda_pg_rca32_and_2_16_y0;
  assign f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_1_17_y0 = f_s_dadda_pg_rca32_and_1_17_y0;
  assign f_s_dadda_pg_rca32_fa91_y0 = f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_3_15_y0 ^ f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_2_16_y0;
  assign f_s_dadda_pg_rca32_fa91_y1 = f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_3_15_y0 & f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_2_16_y0;
  assign f_s_dadda_pg_rca32_fa91_y2 = f_s_dadda_pg_rca32_fa91_y0 ^ f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_1_17_y0;
  assign f_s_dadda_pg_rca32_fa91_y3 = f_s_dadda_pg_rca32_fa91_y0 & f_s_dadda_pg_rca32_fa91_f_s_dadda_pg_rca32_and_1_17_y0;
  assign f_s_dadda_pg_rca32_fa91_y4 = f_s_dadda_pg_rca32_fa91_y1 | f_s_dadda_pg_rca32_fa91_y3;
  assign f_s_dadda_pg_rca32_and_0_18_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_0_18_y0 = f_s_dadda_pg_rca32_and_0_18_a_0 & f_s_dadda_pg_rca32_and_0_18_b_18;
  assign f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_and_0_18_y0 = f_s_dadda_pg_rca32_and_0_18_y0;
  assign f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_fa82_y2 = f_s_dadda_pg_rca32_fa82_y2;
  assign f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_fa83_y2 = f_s_dadda_pg_rca32_fa83_y2;
  assign f_s_dadda_pg_rca32_fa92_y0 = f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_and_0_18_y0 ^ f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_fa82_y2;
  assign f_s_dadda_pg_rca32_fa92_y1 = f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_and_0_18_y0 & f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_fa82_y2;
  assign f_s_dadda_pg_rca32_fa92_y2 = f_s_dadda_pg_rca32_fa92_y0 ^ f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_fa83_y2;
  assign f_s_dadda_pg_rca32_fa92_y3 = f_s_dadda_pg_rca32_fa92_y0 & f_s_dadda_pg_rca32_fa92_f_s_dadda_pg_rca32_fa83_y2;
  assign f_s_dadda_pg_rca32_fa92_y4 = f_s_dadda_pg_rca32_fa92_y1 | f_s_dadda_pg_rca32_fa92_y3;
  assign f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa84_y2 = f_s_dadda_pg_rca32_fa84_y2;
  assign f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa85_y2 = f_s_dadda_pg_rca32_fa85_y2;
  assign f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa86_y2 = f_s_dadda_pg_rca32_fa86_y2;
  assign f_s_dadda_pg_rca32_fa93_y0 = f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa84_y2 ^ f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa85_y2;
  assign f_s_dadda_pg_rca32_fa93_y1 = f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa84_y2 & f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa85_y2;
  assign f_s_dadda_pg_rca32_fa93_y2 = f_s_dadda_pg_rca32_fa93_y0 ^ f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa86_y2;
  assign f_s_dadda_pg_rca32_fa93_y3 = f_s_dadda_pg_rca32_fa93_y0 & f_s_dadda_pg_rca32_fa93_f_s_dadda_pg_rca32_fa86_y2;
  assign f_s_dadda_pg_rca32_fa93_y4 = f_s_dadda_pg_rca32_fa93_y1 | f_s_dadda_pg_rca32_fa93_y3;
  assign f_s_dadda_pg_rca32_ha16_f_s_dadda_pg_rca32_fa87_y2 = f_s_dadda_pg_rca32_fa87_y2;
  assign f_s_dadda_pg_rca32_ha16_f_s_dadda_pg_rca32_fa88_y2 = f_s_dadda_pg_rca32_fa88_y2;
  assign f_s_dadda_pg_rca32_ha16_y0 = f_s_dadda_pg_rca32_ha16_f_s_dadda_pg_rca32_fa87_y2 ^ f_s_dadda_pg_rca32_ha16_f_s_dadda_pg_rca32_fa88_y2;
  assign f_s_dadda_pg_rca32_ha16_y1 = f_s_dadda_pg_rca32_ha16_f_s_dadda_pg_rca32_fa87_y2 & f_s_dadda_pg_rca32_ha16_f_s_dadda_pg_rca32_fa88_y2;
  assign f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_ha16_y1 = f_s_dadda_pg_rca32_ha16_y1;
  assign f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_fa93_y4 = f_s_dadda_pg_rca32_fa93_y4;
  assign f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_fa92_y4 = f_s_dadda_pg_rca32_fa92_y4;
  assign f_s_dadda_pg_rca32_fa94_y0 = f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_ha16_y1 ^ f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_fa93_y4;
  assign f_s_dadda_pg_rca32_fa94_y1 = f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_ha16_y1 & f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_fa93_y4;
  assign f_s_dadda_pg_rca32_fa94_y2 = f_s_dadda_pg_rca32_fa94_y0 ^ f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_fa92_y4;
  assign f_s_dadda_pg_rca32_fa94_y3 = f_s_dadda_pg_rca32_fa94_y0 & f_s_dadda_pg_rca32_fa94_f_s_dadda_pg_rca32_fa92_y4;
  assign f_s_dadda_pg_rca32_fa94_y4 = f_s_dadda_pg_rca32_fa94_y1 | f_s_dadda_pg_rca32_fa94_y3;
  assign f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa91_y4 = f_s_dadda_pg_rca32_fa91_y4;
  assign f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa90_y4 = f_s_dadda_pg_rca32_fa90_y4;
  assign f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa89_y4 = f_s_dadda_pg_rca32_fa89_y4;
  assign f_s_dadda_pg_rca32_fa95_y0 = f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa91_y4 ^ f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa90_y4;
  assign f_s_dadda_pg_rca32_fa95_y1 = f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa91_y4 & f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa90_y4;
  assign f_s_dadda_pg_rca32_fa95_y2 = f_s_dadda_pg_rca32_fa95_y0 ^ f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa89_y4;
  assign f_s_dadda_pg_rca32_fa95_y3 = f_s_dadda_pg_rca32_fa95_y0 & f_s_dadda_pg_rca32_fa95_f_s_dadda_pg_rca32_fa89_y4;
  assign f_s_dadda_pg_rca32_fa95_y4 = f_s_dadda_pg_rca32_fa95_y1 | f_s_dadda_pg_rca32_fa95_y3;
  assign f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa88_y4 = f_s_dadda_pg_rca32_fa88_y4;
  assign f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa87_y4 = f_s_dadda_pg_rca32_fa87_y4;
  assign f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa86_y4 = f_s_dadda_pg_rca32_fa86_y4;
  assign f_s_dadda_pg_rca32_fa96_y0 = f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa88_y4 ^ f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa87_y4;
  assign f_s_dadda_pg_rca32_fa96_y1 = f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa88_y4 & f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa87_y4;
  assign f_s_dadda_pg_rca32_fa96_y2 = f_s_dadda_pg_rca32_fa96_y0 ^ f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa86_y4;
  assign f_s_dadda_pg_rca32_fa96_y3 = f_s_dadda_pg_rca32_fa96_y0 & f_s_dadda_pg_rca32_fa96_f_s_dadda_pg_rca32_fa86_y4;
  assign f_s_dadda_pg_rca32_fa96_y4 = f_s_dadda_pg_rca32_fa96_y1 | f_s_dadda_pg_rca32_fa96_y3;
  assign f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa85_y4 = f_s_dadda_pg_rca32_fa85_y4;
  assign f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa84_y4 = f_s_dadda_pg_rca32_fa84_y4;
  assign f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa83_y4 = f_s_dadda_pg_rca32_fa83_y4;
  assign f_s_dadda_pg_rca32_fa97_y0 = f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa85_y4 ^ f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa84_y4;
  assign f_s_dadda_pg_rca32_fa97_y1 = f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa85_y4 & f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa84_y4;
  assign f_s_dadda_pg_rca32_fa97_y2 = f_s_dadda_pg_rca32_fa97_y0 ^ f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa83_y4;
  assign f_s_dadda_pg_rca32_fa97_y3 = f_s_dadda_pg_rca32_fa97_y0 & f_s_dadda_pg_rca32_fa97_f_s_dadda_pg_rca32_fa83_y4;
  assign f_s_dadda_pg_rca32_fa97_y4 = f_s_dadda_pg_rca32_fa97_y1 | f_s_dadda_pg_rca32_fa97_y3;
  assign f_s_dadda_pg_rca32_and_19_0_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_19_0_y0 = f_s_dadda_pg_rca32_and_19_0_a_19 & f_s_dadda_pg_rca32_and_19_0_b_0;
  assign f_s_dadda_pg_rca32_and_18_1_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_18_1_y0 = f_s_dadda_pg_rca32_and_18_1_a_18 & f_s_dadda_pg_rca32_and_18_1_b_1;
  assign f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_fa82_y4 = f_s_dadda_pg_rca32_fa82_y4;
  assign f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_and_19_0_y0 = f_s_dadda_pg_rca32_and_19_0_y0;
  assign f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_and_18_1_y0 = f_s_dadda_pg_rca32_and_18_1_y0;
  assign f_s_dadda_pg_rca32_fa98_y0 = f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_fa82_y4 ^ f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_and_19_0_y0;
  assign f_s_dadda_pg_rca32_fa98_y1 = f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_fa82_y4 & f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_and_19_0_y0;
  assign f_s_dadda_pg_rca32_fa98_y2 = f_s_dadda_pg_rca32_fa98_y0 ^ f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_and_18_1_y0;
  assign f_s_dadda_pg_rca32_fa98_y3 = f_s_dadda_pg_rca32_fa98_y0 & f_s_dadda_pg_rca32_fa98_f_s_dadda_pg_rca32_and_18_1_y0;
  assign f_s_dadda_pg_rca32_fa98_y4 = f_s_dadda_pg_rca32_fa98_y1 | f_s_dadda_pg_rca32_fa98_y3;
  assign f_s_dadda_pg_rca32_and_17_2_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_17_2_y0 = f_s_dadda_pg_rca32_and_17_2_a_17 & f_s_dadda_pg_rca32_and_17_2_b_2;
  assign f_s_dadda_pg_rca32_and_16_3_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_16_3_y0 = f_s_dadda_pg_rca32_and_16_3_a_16 & f_s_dadda_pg_rca32_and_16_3_b_3;
  assign f_s_dadda_pg_rca32_and_15_4_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_15_4_y0 = f_s_dadda_pg_rca32_and_15_4_a_15 & f_s_dadda_pg_rca32_and_15_4_b_4;
  assign f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_17_2_y0 = f_s_dadda_pg_rca32_and_17_2_y0;
  assign f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_16_3_y0 = f_s_dadda_pg_rca32_and_16_3_y0;
  assign f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_15_4_y0 = f_s_dadda_pg_rca32_and_15_4_y0;
  assign f_s_dadda_pg_rca32_fa99_y0 = f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_17_2_y0 ^ f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_16_3_y0;
  assign f_s_dadda_pg_rca32_fa99_y1 = f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_17_2_y0 & f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_16_3_y0;
  assign f_s_dadda_pg_rca32_fa99_y2 = f_s_dadda_pg_rca32_fa99_y0 ^ f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_15_4_y0;
  assign f_s_dadda_pg_rca32_fa99_y3 = f_s_dadda_pg_rca32_fa99_y0 & f_s_dadda_pg_rca32_fa99_f_s_dadda_pg_rca32_and_15_4_y0;
  assign f_s_dadda_pg_rca32_fa99_y4 = f_s_dadda_pg_rca32_fa99_y1 | f_s_dadda_pg_rca32_fa99_y3;
  assign f_s_dadda_pg_rca32_and_14_5_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_14_5_y0 = f_s_dadda_pg_rca32_and_14_5_a_14 & f_s_dadda_pg_rca32_and_14_5_b_5;
  assign f_s_dadda_pg_rca32_and_13_6_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_13_6_y0 = f_s_dadda_pg_rca32_and_13_6_a_13 & f_s_dadda_pg_rca32_and_13_6_b_6;
  assign f_s_dadda_pg_rca32_and_12_7_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_12_7_y0 = f_s_dadda_pg_rca32_and_12_7_a_12 & f_s_dadda_pg_rca32_and_12_7_b_7;
  assign f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_14_5_y0 = f_s_dadda_pg_rca32_and_14_5_y0;
  assign f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_13_6_y0 = f_s_dadda_pg_rca32_and_13_6_y0;
  assign f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_12_7_y0 = f_s_dadda_pg_rca32_and_12_7_y0;
  assign f_s_dadda_pg_rca32_fa100_y0 = f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_14_5_y0 ^ f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_13_6_y0;
  assign f_s_dadda_pg_rca32_fa100_y1 = f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_14_5_y0 & f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_13_6_y0;
  assign f_s_dadda_pg_rca32_fa100_y2 = f_s_dadda_pg_rca32_fa100_y0 ^ f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_12_7_y0;
  assign f_s_dadda_pg_rca32_fa100_y3 = f_s_dadda_pg_rca32_fa100_y0 & f_s_dadda_pg_rca32_fa100_f_s_dadda_pg_rca32_and_12_7_y0;
  assign f_s_dadda_pg_rca32_fa100_y4 = f_s_dadda_pg_rca32_fa100_y1 | f_s_dadda_pg_rca32_fa100_y3;
  assign f_s_dadda_pg_rca32_and_11_8_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_11_8_y0 = f_s_dadda_pg_rca32_and_11_8_a_11 & f_s_dadda_pg_rca32_and_11_8_b_8;
  assign f_s_dadda_pg_rca32_and_10_9_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_10_9_y0 = f_s_dadda_pg_rca32_and_10_9_a_10 & f_s_dadda_pg_rca32_and_10_9_b_9;
  assign f_s_dadda_pg_rca32_and_9_10_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_9_10_y0 = f_s_dadda_pg_rca32_and_9_10_a_9 & f_s_dadda_pg_rca32_and_9_10_b_10;
  assign f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_11_8_y0 = f_s_dadda_pg_rca32_and_11_8_y0;
  assign f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_10_9_y0 = f_s_dadda_pg_rca32_and_10_9_y0;
  assign f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_9_10_y0 = f_s_dadda_pg_rca32_and_9_10_y0;
  assign f_s_dadda_pg_rca32_fa101_y0 = f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_11_8_y0 ^ f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_10_9_y0;
  assign f_s_dadda_pg_rca32_fa101_y1 = f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_11_8_y0 & f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_10_9_y0;
  assign f_s_dadda_pg_rca32_fa101_y2 = f_s_dadda_pg_rca32_fa101_y0 ^ f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_9_10_y0;
  assign f_s_dadda_pg_rca32_fa101_y3 = f_s_dadda_pg_rca32_fa101_y0 & f_s_dadda_pg_rca32_fa101_f_s_dadda_pg_rca32_and_9_10_y0;
  assign f_s_dadda_pg_rca32_fa101_y4 = f_s_dadda_pg_rca32_fa101_y1 | f_s_dadda_pg_rca32_fa101_y3;
  assign f_s_dadda_pg_rca32_and_8_11_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_8_11_y0 = f_s_dadda_pg_rca32_and_8_11_a_8 & f_s_dadda_pg_rca32_and_8_11_b_11;
  assign f_s_dadda_pg_rca32_and_7_12_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_7_12_y0 = f_s_dadda_pg_rca32_and_7_12_a_7 & f_s_dadda_pg_rca32_and_7_12_b_12;
  assign f_s_dadda_pg_rca32_and_6_13_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_6_13_y0 = f_s_dadda_pg_rca32_and_6_13_a_6 & f_s_dadda_pg_rca32_and_6_13_b_13;
  assign f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_8_11_y0 = f_s_dadda_pg_rca32_and_8_11_y0;
  assign f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_7_12_y0 = f_s_dadda_pg_rca32_and_7_12_y0;
  assign f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_6_13_y0 = f_s_dadda_pg_rca32_and_6_13_y0;
  assign f_s_dadda_pg_rca32_fa102_y0 = f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_8_11_y0 ^ f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_7_12_y0;
  assign f_s_dadda_pg_rca32_fa102_y1 = f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_8_11_y0 & f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_7_12_y0;
  assign f_s_dadda_pg_rca32_fa102_y2 = f_s_dadda_pg_rca32_fa102_y0 ^ f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_6_13_y0;
  assign f_s_dadda_pg_rca32_fa102_y3 = f_s_dadda_pg_rca32_fa102_y0 & f_s_dadda_pg_rca32_fa102_f_s_dadda_pg_rca32_and_6_13_y0;
  assign f_s_dadda_pg_rca32_fa102_y4 = f_s_dadda_pg_rca32_fa102_y1 | f_s_dadda_pg_rca32_fa102_y3;
  assign f_s_dadda_pg_rca32_and_5_14_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_5_14_y0 = f_s_dadda_pg_rca32_and_5_14_a_5 & f_s_dadda_pg_rca32_and_5_14_b_14;
  assign f_s_dadda_pg_rca32_and_4_15_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_4_15_y0 = f_s_dadda_pg_rca32_and_4_15_a_4 & f_s_dadda_pg_rca32_and_4_15_b_15;
  assign f_s_dadda_pg_rca32_and_3_16_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_3_16_y0 = f_s_dadda_pg_rca32_and_3_16_a_3 & f_s_dadda_pg_rca32_and_3_16_b_16;
  assign f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_5_14_y0 = f_s_dadda_pg_rca32_and_5_14_y0;
  assign f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_4_15_y0 = f_s_dadda_pg_rca32_and_4_15_y0;
  assign f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_3_16_y0 = f_s_dadda_pg_rca32_and_3_16_y0;
  assign f_s_dadda_pg_rca32_fa103_y0 = f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_5_14_y0 ^ f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_4_15_y0;
  assign f_s_dadda_pg_rca32_fa103_y1 = f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_5_14_y0 & f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_4_15_y0;
  assign f_s_dadda_pg_rca32_fa103_y2 = f_s_dadda_pg_rca32_fa103_y0 ^ f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_3_16_y0;
  assign f_s_dadda_pg_rca32_fa103_y3 = f_s_dadda_pg_rca32_fa103_y0 & f_s_dadda_pg_rca32_fa103_f_s_dadda_pg_rca32_and_3_16_y0;
  assign f_s_dadda_pg_rca32_fa103_y4 = f_s_dadda_pg_rca32_fa103_y1 | f_s_dadda_pg_rca32_fa103_y3;
  assign f_s_dadda_pg_rca32_and_2_17_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_2_17_y0 = f_s_dadda_pg_rca32_and_2_17_a_2 & f_s_dadda_pg_rca32_and_2_17_b_17;
  assign f_s_dadda_pg_rca32_and_1_18_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_1_18_y0 = f_s_dadda_pg_rca32_and_1_18_a_1 & f_s_dadda_pg_rca32_and_1_18_b_18;
  assign f_s_dadda_pg_rca32_and_0_19_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_0_19_y0 = f_s_dadda_pg_rca32_and_0_19_a_0 & f_s_dadda_pg_rca32_and_0_19_b_19;
  assign f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_2_17_y0 = f_s_dadda_pg_rca32_and_2_17_y0;
  assign f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_1_18_y0 = f_s_dadda_pg_rca32_and_1_18_y0;
  assign f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_0_19_y0 = f_s_dadda_pg_rca32_and_0_19_y0;
  assign f_s_dadda_pg_rca32_fa104_y0 = f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_2_17_y0 ^ f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_1_18_y0;
  assign f_s_dadda_pg_rca32_fa104_y1 = f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_2_17_y0 & f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_1_18_y0;
  assign f_s_dadda_pg_rca32_fa104_y2 = f_s_dadda_pg_rca32_fa104_y0 ^ f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_0_19_y0;
  assign f_s_dadda_pg_rca32_fa104_y3 = f_s_dadda_pg_rca32_fa104_y0 & f_s_dadda_pg_rca32_fa104_f_s_dadda_pg_rca32_and_0_19_y0;
  assign f_s_dadda_pg_rca32_fa104_y4 = f_s_dadda_pg_rca32_fa104_y1 | f_s_dadda_pg_rca32_fa104_y3;
  assign f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa94_y2 = f_s_dadda_pg_rca32_fa94_y2;
  assign f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa95_y2 = f_s_dadda_pg_rca32_fa95_y2;
  assign f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa96_y2 = f_s_dadda_pg_rca32_fa96_y2;
  assign f_s_dadda_pg_rca32_fa105_y0 = f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa94_y2 ^ f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa95_y2;
  assign f_s_dadda_pg_rca32_fa105_y1 = f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa94_y2 & f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa95_y2;
  assign f_s_dadda_pg_rca32_fa105_y2 = f_s_dadda_pg_rca32_fa105_y0 ^ f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa96_y2;
  assign f_s_dadda_pg_rca32_fa105_y3 = f_s_dadda_pg_rca32_fa105_y0 & f_s_dadda_pg_rca32_fa105_f_s_dadda_pg_rca32_fa96_y2;
  assign f_s_dadda_pg_rca32_fa105_y4 = f_s_dadda_pg_rca32_fa105_y1 | f_s_dadda_pg_rca32_fa105_y3;
  assign f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa97_y2 = f_s_dadda_pg_rca32_fa97_y2;
  assign f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa98_y2 = f_s_dadda_pg_rca32_fa98_y2;
  assign f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa99_y2 = f_s_dadda_pg_rca32_fa99_y2;
  assign f_s_dadda_pg_rca32_fa106_y0 = f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa97_y2 ^ f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa98_y2;
  assign f_s_dadda_pg_rca32_fa106_y1 = f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa97_y2 & f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa98_y2;
  assign f_s_dadda_pg_rca32_fa106_y2 = f_s_dadda_pg_rca32_fa106_y0 ^ f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa99_y2;
  assign f_s_dadda_pg_rca32_fa106_y3 = f_s_dadda_pg_rca32_fa106_y0 & f_s_dadda_pg_rca32_fa106_f_s_dadda_pg_rca32_fa99_y2;
  assign f_s_dadda_pg_rca32_fa106_y4 = f_s_dadda_pg_rca32_fa106_y1 | f_s_dadda_pg_rca32_fa106_y3;
  assign f_s_dadda_pg_rca32_ha17_f_s_dadda_pg_rca32_fa100_y2 = f_s_dadda_pg_rca32_fa100_y2;
  assign f_s_dadda_pg_rca32_ha17_f_s_dadda_pg_rca32_fa101_y2 = f_s_dadda_pg_rca32_fa101_y2;
  assign f_s_dadda_pg_rca32_ha17_y0 = f_s_dadda_pg_rca32_ha17_f_s_dadda_pg_rca32_fa100_y2 ^ f_s_dadda_pg_rca32_ha17_f_s_dadda_pg_rca32_fa101_y2;
  assign f_s_dadda_pg_rca32_ha17_y1 = f_s_dadda_pg_rca32_ha17_f_s_dadda_pg_rca32_fa100_y2 & f_s_dadda_pg_rca32_ha17_f_s_dadda_pg_rca32_fa101_y2;
  assign f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_ha17_y1 = f_s_dadda_pg_rca32_ha17_y1;
  assign f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_fa106_y4 = f_s_dadda_pg_rca32_fa106_y4;
  assign f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_fa105_y4 = f_s_dadda_pg_rca32_fa105_y4;
  assign f_s_dadda_pg_rca32_fa107_y0 = f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_ha17_y1 ^ f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_fa106_y4;
  assign f_s_dadda_pg_rca32_fa107_y1 = f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_ha17_y1 & f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_fa106_y4;
  assign f_s_dadda_pg_rca32_fa107_y2 = f_s_dadda_pg_rca32_fa107_y0 ^ f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_fa105_y4;
  assign f_s_dadda_pg_rca32_fa107_y3 = f_s_dadda_pg_rca32_fa107_y0 & f_s_dadda_pg_rca32_fa107_f_s_dadda_pg_rca32_fa105_y4;
  assign f_s_dadda_pg_rca32_fa107_y4 = f_s_dadda_pg_rca32_fa107_y1 | f_s_dadda_pg_rca32_fa107_y3;
  assign f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa104_y4 = f_s_dadda_pg_rca32_fa104_y4;
  assign f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa103_y4 = f_s_dadda_pg_rca32_fa103_y4;
  assign f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa102_y4 = f_s_dadda_pg_rca32_fa102_y4;
  assign f_s_dadda_pg_rca32_fa108_y0 = f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa104_y4 ^ f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa103_y4;
  assign f_s_dadda_pg_rca32_fa108_y1 = f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa104_y4 & f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa103_y4;
  assign f_s_dadda_pg_rca32_fa108_y2 = f_s_dadda_pg_rca32_fa108_y0 ^ f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa102_y4;
  assign f_s_dadda_pg_rca32_fa108_y3 = f_s_dadda_pg_rca32_fa108_y0 & f_s_dadda_pg_rca32_fa108_f_s_dadda_pg_rca32_fa102_y4;
  assign f_s_dadda_pg_rca32_fa108_y4 = f_s_dadda_pg_rca32_fa108_y1 | f_s_dadda_pg_rca32_fa108_y3;
  assign f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa101_y4 = f_s_dadda_pg_rca32_fa101_y4;
  assign f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa100_y4 = f_s_dadda_pg_rca32_fa100_y4;
  assign f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa99_y4 = f_s_dadda_pg_rca32_fa99_y4;
  assign f_s_dadda_pg_rca32_fa109_y0 = f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa101_y4 ^ f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa100_y4;
  assign f_s_dadda_pg_rca32_fa109_y1 = f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa101_y4 & f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa100_y4;
  assign f_s_dadda_pg_rca32_fa109_y2 = f_s_dadda_pg_rca32_fa109_y0 ^ f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa99_y4;
  assign f_s_dadda_pg_rca32_fa109_y3 = f_s_dadda_pg_rca32_fa109_y0 & f_s_dadda_pg_rca32_fa109_f_s_dadda_pg_rca32_fa99_y4;
  assign f_s_dadda_pg_rca32_fa109_y4 = f_s_dadda_pg_rca32_fa109_y1 | f_s_dadda_pg_rca32_fa109_y3;
  assign f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa98_y4 = f_s_dadda_pg_rca32_fa98_y4;
  assign f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa97_y4 = f_s_dadda_pg_rca32_fa97_y4;
  assign f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa96_y4 = f_s_dadda_pg_rca32_fa96_y4;
  assign f_s_dadda_pg_rca32_fa110_y0 = f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa98_y4 ^ f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa97_y4;
  assign f_s_dadda_pg_rca32_fa110_y1 = f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa98_y4 & f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa97_y4;
  assign f_s_dadda_pg_rca32_fa110_y2 = f_s_dadda_pg_rca32_fa110_y0 ^ f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa96_y4;
  assign f_s_dadda_pg_rca32_fa110_y3 = f_s_dadda_pg_rca32_fa110_y0 & f_s_dadda_pg_rca32_fa110_f_s_dadda_pg_rca32_fa96_y4;
  assign f_s_dadda_pg_rca32_fa110_y4 = f_s_dadda_pg_rca32_fa110_y1 | f_s_dadda_pg_rca32_fa110_y3;
  assign f_s_dadda_pg_rca32_and_20_0_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_20_0_y0 = f_s_dadda_pg_rca32_and_20_0_a_20 & f_s_dadda_pg_rca32_and_20_0_b_0;
  assign f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_fa95_y4 = f_s_dadda_pg_rca32_fa95_y4;
  assign f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_fa94_y4 = f_s_dadda_pg_rca32_fa94_y4;
  assign f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_and_20_0_y0 = f_s_dadda_pg_rca32_and_20_0_y0;
  assign f_s_dadda_pg_rca32_fa111_y0 = f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_fa95_y4 ^ f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_fa94_y4;
  assign f_s_dadda_pg_rca32_fa111_y1 = f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_fa95_y4 & f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_fa94_y4;
  assign f_s_dadda_pg_rca32_fa111_y2 = f_s_dadda_pg_rca32_fa111_y0 ^ f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_and_20_0_y0;
  assign f_s_dadda_pg_rca32_fa111_y3 = f_s_dadda_pg_rca32_fa111_y0 & f_s_dadda_pg_rca32_fa111_f_s_dadda_pg_rca32_and_20_0_y0;
  assign f_s_dadda_pg_rca32_fa111_y4 = f_s_dadda_pg_rca32_fa111_y1 | f_s_dadda_pg_rca32_fa111_y3;
  assign f_s_dadda_pg_rca32_and_19_1_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_19_1_y0 = f_s_dadda_pg_rca32_and_19_1_a_19 & f_s_dadda_pg_rca32_and_19_1_b_1;
  assign f_s_dadda_pg_rca32_and_18_2_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_18_2_y0 = f_s_dadda_pg_rca32_and_18_2_a_18 & f_s_dadda_pg_rca32_and_18_2_b_2;
  assign f_s_dadda_pg_rca32_and_17_3_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_17_3_y0 = f_s_dadda_pg_rca32_and_17_3_a_17 & f_s_dadda_pg_rca32_and_17_3_b_3;
  assign f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_19_1_y0 = f_s_dadda_pg_rca32_and_19_1_y0;
  assign f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_18_2_y0 = f_s_dadda_pg_rca32_and_18_2_y0;
  assign f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_17_3_y0 = f_s_dadda_pg_rca32_and_17_3_y0;
  assign f_s_dadda_pg_rca32_fa112_y0 = f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_19_1_y0 ^ f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_18_2_y0;
  assign f_s_dadda_pg_rca32_fa112_y1 = f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_19_1_y0 & f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_18_2_y0;
  assign f_s_dadda_pg_rca32_fa112_y2 = f_s_dadda_pg_rca32_fa112_y0 ^ f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_17_3_y0;
  assign f_s_dadda_pg_rca32_fa112_y3 = f_s_dadda_pg_rca32_fa112_y0 & f_s_dadda_pg_rca32_fa112_f_s_dadda_pg_rca32_and_17_3_y0;
  assign f_s_dadda_pg_rca32_fa112_y4 = f_s_dadda_pg_rca32_fa112_y1 | f_s_dadda_pg_rca32_fa112_y3;
  assign f_s_dadda_pg_rca32_and_16_4_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_16_4_y0 = f_s_dadda_pg_rca32_and_16_4_a_16 & f_s_dadda_pg_rca32_and_16_4_b_4;
  assign f_s_dadda_pg_rca32_and_15_5_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_15_5_y0 = f_s_dadda_pg_rca32_and_15_5_a_15 & f_s_dadda_pg_rca32_and_15_5_b_5;
  assign f_s_dadda_pg_rca32_and_14_6_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_14_6_y0 = f_s_dadda_pg_rca32_and_14_6_a_14 & f_s_dadda_pg_rca32_and_14_6_b_6;
  assign f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_16_4_y0 = f_s_dadda_pg_rca32_and_16_4_y0;
  assign f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_15_5_y0 = f_s_dadda_pg_rca32_and_15_5_y0;
  assign f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_14_6_y0 = f_s_dadda_pg_rca32_and_14_6_y0;
  assign f_s_dadda_pg_rca32_fa113_y0 = f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_16_4_y0 ^ f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_15_5_y0;
  assign f_s_dadda_pg_rca32_fa113_y1 = f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_16_4_y0 & f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_15_5_y0;
  assign f_s_dadda_pg_rca32_fa113_y2 = f_s_dadda_pg_rca32_fa113_y0 ^ f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_14_6_y0;
  assign f_s_dadda_pg_rca32_fa113_y3 = f_s_dadda_pg_rca32_fa113_y0 & f_s_dadda_pg_rca32_fa113_f_s_dadda_pg_rca32_and_14_6_y0;
  assign f_s_dadda_pg_rca32_fa113_y4 = f_s_dadda_pg_rca32_fa113_y1 | f_s_dadda_pg_rca32_fa113_y3;
  assign f_s_dadda_pg_rca32_and_13_7_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_13_7_y0 = f_s_dadda_pg_rca32_and_13_7_a_13 & f_s_dadda_pg_rca32_and_13_7_b_7;
  assign f_s_dadda_pg_rca32_and_12_8_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_12_8_y0 = f_s_dadda_pg_rca32_and_12_8_a_12 & f_s_dadda_pg_rca32_and_12_8_b_8;
  assign f_s_dadda_pg_rca32_and_11_9_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_11_9_y0 = f_s_dadda_pg_rca32_and_11_9_a_11 & f_s_dadda_pg_rca32_and_11_9_b_9;
  assign f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_13_7_y0 = f_s_dadda_pg_rca32_and_13_7_y0;
  assign f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_12_8_y0 = f_s_dadda_pg_rca32_and_12_8_y0;
  assign f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_11_9_y0 = f_s_dadda_pg_rca32_and_11_9_y0;
  assign f_s_dadda_pg_rca32_fa114_y0 = f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_13_7_y0 ^ f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_12_8_y0;
  assign f_s_dadda_pg_rca32_fa114_y1 = f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_13_7_y0 & f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_12_8_y0;
  assign f_s_dadda_pg_rca32_fa114_y2 = f_s_dadda_pg_rca32_fa114_y0 ^ f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_11_9_y0;
  assign f_s_dadda_pg_rca32_fa114_y3 = f_s_dadda_pg_rca32_fa114_y0 & f_s_dadda_pg_rca32_fa114_f_s_dadda_pg_rca32_and_11_9_y0;
  assign f_s_dadda_pg_rca32_fa114_y4 = f_s_dadda_pg_rca32_fa114_y1 | f_s_dadda_pg_rca32_fa114_y3;
  assign f_s_dadda_pg_rca32_and_10_10_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_10_10_y0 = f_s_dadda_pg_rca32_and_10_10_a_10 & f_s_dadda_pg_rca32_and_10_10_b_10;
  assign f_s_dadda_pg_rca32_and_9_11_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_9_11_y0 = f_s_dadda_pg_rca32_and_9_11_a_9 & f_s_dadda_pg_rca32_and_9_11_b_11;
  assign f_s_dadda_pg_rca32_and_8_12_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_8_12_y0 = f_s_dadda_pg_rca32_and_8_12_a_8 & f_s_dadda_pg_rca32_and_8_12_b_12;
  assign f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_10_10_y0 = f_s_dadda_pg_rca32_and_10_10_y0;
  assign f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_9_11_y0 = f_s_dadda_pg_rca32_and_9_11_y0;
  assign f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_8_12_y0 = f_s_dadda_pg_rca32_and_8_12_y0;
  assign f_s_dadda_pg_rca32_fa115_y0 = f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_10_10_y0 ^ f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_9_11_y0;
  assign f_s_dadda_pg_rca32_fa115_y1 = f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_10_10_y0 & f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_9_11_y0;
  assign f_s_dadda_pg_rca32_fa115_y2 = f_s_dadda_pg_rca32_fa115_y0 ^ f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_8_12_y0;
  assign f_s_dadda_pg_rca32_fa115_y3 = f_s_dadda_pg_rca32_fa115_y0 & f_s_dadda_pg_rca32_fa115_f_s_dadda_pg_rca32_and_8_12_y0;
  assign f_s_dadda_pg_rca32_fa115_y4 = f_s_dadda_pg_rca32_fa115_y1 | f_s_dadda_pg_rca32_fa115_y3;
  assign f_s_dadda_pg_rca32_and_7_13_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_7_13_y0 = f_s_dadda_pg_rca32_and_7_13_a_7 & f_s_dadda_pg_rca32_and_7_13_b_13;
  assign f_s_dadda_pg_rca32_and_6_14_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_6_14_y0 = f_s_dadda_pg_rca32_and_6_14_a_6 & f_s_dadda_pg_rca32_and_6_14_b_14;
  assign f_s_dadda_pg_rca32_and_5_15_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_5_15_y0 = f_s_dadda_pg_rca32_and_5_15_a_5 & f_s_dadda_pg_rca32_and_5_15_b_15;
  assign f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_7_13_y0 = f_s_dadda_pg_rca32_and_7_13_y0;
  assign f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_6_14_y0 = f_s_dadda_pg_rca32_and_6_14_y0;
  assign f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_5_15_y0 = f_s_dadda_pg_rca32_and_5_15_y0;
  assign f_s_dadda_pg_rca32_fa116_y0 = f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_7_13_y0 ^ f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_6_14_y0;
  assign f_s_dadda_pg_rca32_fa116_y1 = f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_7_13_y0 & f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_6_14_y0;
  assign f_s_dadda_pg_rca32_fa116_y2 = f_s_dadda_pg_rca32_fa116_y0 ^ f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_5_15_y0;
  assign f_s_dadda_pg_rca32_fa116_y3 = f_s_dadda_pg_rca32_fa116_y0 & f_s_dadda_pg_rca32_fa116_f_s_dadda_pg_rca32_and_5_15_y0;
  assign f_s_dadda_pg_rca32_fa116_y4 = f_s_dadda_pg_rca32_fa116_y1 | f_s_dadda_pg_rca32_fa116_y3;
  assign f_s_dadda_pg_rca32_and_4_16_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_4_16_y0 = f_s_dadda_pg_rca32_and_4_16_a_4 & f_s_dadda_pg_rca32_and_4_16_b_16;
  assign f_s_dadda_pg_rca32_and_3_17_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_3_17_y0 = f_s_dadda_pg_rca32_and_3_17_a_3 & f_s_dadda_pg_rca32_and_3_17_b_17;
  assign f_s_dadda_pg_rca32_and_2_18_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_2_18_y0 = f_s_dadda_pg_rca32_and_2_18_a_2 & f_s_dadda_pg_rca32_and_2_18_b_18;
  assign f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_4_16_y0 = f_s_dadda_pg_rca32_and_4_16_y0;
  assign f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_3_17_y0 = f_s_dadda_pg_rca32_and_3_17_y0;
  assign f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_2_18_y0 = f_s_dadda_pg_rca32_and_2_18_y0;
  assign f_s_dadda_pg_rca32_fa117_y0 = f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_4_16_y0 ^ f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_3_17_y0;
  assign f_s_dadda_pg_rca32_fa117_y1 = f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_4_16_y0 & f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_3_17_y0;
  assign f_s_dadda_pg_rca32_fa117_y2 = f_s_dadda_pg_rca32_fa117_y0 ^ f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_2_18_y0;
  assign f_s_dadda_pg_rca32_fa117_y3 = f_s_dadda_pg_rca32_fa117_y0 & f_s_dadda_pg_rca32_fa117_f_s_dadda_pg_rca32_and_2_18_y0;
  assign f_s_dadda_pg_rca32_fa117_y4 = f_s_dadda_pg_rca32_fa117_y1 | f_s_dadda_pg_rca32_fa117_y3;
  assign f_s_dadda_pg_rca32_and_1_19_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_1_19_y0 = f_s_dadda_pg_rca32_and_1_19_a_1 & f_s_dadda_pg_rca32_and_1_19_b_19;
  assign f_s_dadda_pg_rca32_and_0_20_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_0_20_y0 = f_s_dadda_pg_rca32_and_0_20_a_0 & f_s_dadda_pg_rca32_and_0_20_b_20;
  assign f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_and_1_19_y0 = f_s_dadda_pg_rca32_and_1_19_y0;
  assign f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_and_0_20_y0 = f_s_dadda_pg_rca32_and_0_20_y0;
  assign f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_fa107_y2 = f_s_dadda_pg_rca32_fa107_y2;
  assign f_s_dadda_pg_rca32_fa118_y0 = f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_and_1_19_y0 ^ f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_and_0_20_y0;
  assign f_s_dadda_pg_rca32_fa118_y1 = f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_and_1_19_y0 & f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_and_0_20_y0;
  assign f_s_dadda_pg_rca32_fa118_y2 = f_s_dadda_pg_rca32_fa118_y0 ^ f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_fa107_y2;
  assign f_s_dadda_pg_rca32_fa118_y3 = f_s_dadda_pg_rca32_fa118_y0 & f_s_dadda_pg_rca32_fa118_f_s_dadda_pg_rca32_fa107_y2;
  assign f_s_dadda_pg_rca32_fa118_y4 = f_s_dadda_pg_rca32_fa118_y1 | f_s_dadda_pg_rca32_fa118_y3;
  assign f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa108_y2 = f_s_dadda_pg_rca32_fa108_y2;
  assign f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa109_y2 = f_s_dadda_pg_rca32_fa109_y2;
  assign f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa110_y2 = f_s_dadda_pg_rca32_fa110_y2;
  assign f_s_dadda_pg_rca32_fa119_y0 = f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa108_y2 ^ f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa109_y2;
  assign f_s_dadda_pg_rca32_fa119_y1 = f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa108_y2 & f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa109_y2;
  assign f_s_dadda_pg_rca32_fa119_y2 = f_s_dadda_pg_rca32_fa119_y0 ^ f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa110_y2;
  assign f_s_dadda_pg_rca32_fa119_y3 = f_s_dadda_pg_rca32_fa119_y0 & f_s_dadda_pg_rca32_fa119_f_s_dadda_pg_rca32_fa110_y2;
  assign f_s_dadda_pg_rca32_fa119_y4 = f_s_dadda_pg_rca32_fa119_y1 | f_s_dadda_pg_rca32_fa119_y3;
  assign f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa111_y2 = f_s_dadda_pg_rca32_fa111_y2;
  assign f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa112_y2 = f_s_dadda_pg_rca32_fa112_y2;
  assign f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa113_y2 = f_s_dadda_pg_rca32_fa113_y2;
  assign f_s_dadda_pg_rca32_fa120_y0 = f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa111_y2 ^ f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa112_y2;
  assign f_s_dadda_pg_rca32_fa120_y1 = f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa111_y2 & f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa112_y2;
  assign f_s_dadda_pg_rca32_fa120_y2 = f_s_dadda_pg_rca32_fa120_y0 ^ f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa113_y2;
  assign f_s_dadda_pg_rca32_fa120_y3 = f_s_dadda_pg_rca32_fa120_y0 & f_s_dadda_pg_rca32_fa120_f_s_dadda_pg_rca32_fa113_y2;
  assign f_s_dadda_pg_rca32_fa120_y4 = f_s_dadda_pg_rca32_fa120_y1 | f_s_dadda_pg_rca32_fa120_y3;
  assign f_s_dadda_pg_rca32_ha18_f_s_dadda_pg_rca32_fa114_y2 = f_s_dadda_pg_rca32_fa114_y2;
  assign f_s_dadda_pg_rca32_ha18_f_s_dadda_pg_rca32_fa115_y2 = f_s_dadda_pg_rca32_fa115_y2;
  assign f_s_dadda_pg_rca32_ha18_y0 = f_s_dadda_pg_rca32_ha18_f_s_dadda_pg_rca32_fa114_y2 ^ f_s_dadda_pg_rca32_ha18_f_s_dadda_pg_rca32_fa115_y2;
  assign f_s_dadda_pg_rca32_ha18_y1 = f_s_dadda_pg_rca32_ha18_f_s_dadda_pg_rca32_fa114_y2 & f_s_dadda_pg_rca32_ha18_f_s_dadda_pg_rca32_fa115_y2;
  assign f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_ha18_y1 = f_s_dadda_pg_rca32_ha18_y1;
  assign f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_fa120_y4 = f_s_dadda_pg_rca32_fa120_y4;
  assign f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_fa119_y4 = f_s_dadda_pg_rca32_fa119_y4;
  assign f_s_dadda_pg_rca32_fa121_y0 = f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_ha18_y1 ^ f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_fa120_y4;
  assign f_s_dadda_pg_rca32_fa121_y1 = f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_ha18_y1 & f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_fa120_y4;
  assign f_s_dadda_pg_rca32_fa121_y2 = f_s_dadda_pg_rca32_fa121_y0 ^ f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_fa119_y4;
  assign f_s_dadda_pg_rca32_fa121_y3 = f_s_dadda_pg_rca32_fa121_y0 & f_s_dadda_pg_rca32_fa121_f_s_dadda_pg_rca32_fa119_y4;
  assign f_s_dadda_pg_rca32_fa121_y4 = f_s_dadda_pg_rca32_fa121_y1 | f_s_dadda_pg_rca32_fa121_y3;
  assign f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa118_y4 = f_s_dadda_pg_rca32_fa118_y4;
  assign f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa117_y4 = f_s_dadda_pg_rca32_fa117_y4;
  assign f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa116_y4 = f_s_dadda_pg_rca32_fa116_y4;
  assign f_s_dadda_pg_rca32_fa122_y0 = f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa118_y4 ^ f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa117_y4;
  assign f_s_dadda_pg_rca32_fa122_y1 = f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa118_y4 & f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa117_y4;
  assign f_s_dadda_pg_rca32_fa122_y2 = f_s_dadda_pg_rca32_fa122_y0 ^ f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa116_y4;
  assign f_s_dadda_pg_rca32_fa122_y3 = f_s_dadda_pg_rca32_fa122_y0 & f_s_dadda_pg_rca32_fa122_f_s_dadda_pg_rca32_fa116_y4;
  assign f_s_dadda_pg_rca32_fa122_y4 = f_s_dadda_pg_rca32_fa122_y1 | f_s_dadda_pg_rca32_fa122_y3;
  assign f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa115_y4 = f_s_dadda_pg_rca32_fa115_y4;
  assign f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa114_y4 = f_s_dadda_pg_rca32_fa114_y4;
  assign f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa113_y4 = f_s_dadda_pg_rca32_fa113_y4;
  assign f_s_dadda_pg_rca32_fa123_y0 = f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa115_y4 ^ f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa114_y4;
  assign f_s_dadda_pg_rca32_fa123_y1 = f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa115_y4 & f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa114_y4;
  assign f_s_dadda_pg_rca32_fa123_y2 = f_s_dadda_pg_rca32_fa123_y0 ^ f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa113_y4;
  assign f_s_dadda_pg_rca32_fa123_y3 = f_s_dadda_pg_rca32_fa123_y0 & f_s_dadda_pg_rca32_fa123_f_s_dadda_pg_rca32_fa113_y4;
  assign f_s_dadda_pg_rca32_fa123_y4 = f_s_dadda_pg_rca32_fa123_y1 | f_s_dadda_pg_rca32_fa123_y3;
  assign f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa112_y4 = f_s_dadda_pg_rca32_fa112_y4;
  assign f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa111_y4 = f_s_dadda_pg_rca32_fa111_y4;
  assign f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa110_y4 = f_s_dadda_pg_rca32_fa110_y4;
  assign f_s_dadda_pg_rca32_fa124_y0 = f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa112_y4 ^ f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa111_y4;
  assign f_s_dadda_pg_rca32_fa124_y1 = f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa112_y4 & f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa111_y4;
  assign f_s_dadda_pg_rca32_fa124_y2 = f_s_dadda_pg_rca32_fa124_y0 ^ f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa110_y4;
  assign f_s_dadda_pg_rca32_fa124_y3 = f_s_dadda_pg_rca32_fa124_y0 & f_s_dadda_pg_rca32_fa124_f_s_dadda_pg_rca32_fa110_y4;
  assign f_s_dadda_pg_rca32_fa124_y4 = f_s_dadda_pg_rca32_fa124_y1 | f_s_dadda_pg_rca32_fa124_y3;
  assign f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa109_y4 = f_s_dadda_pg_rca32_fa109_y4;
  assign f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa108_y4 = f_s_dadda_pg_rca32_fa108_y4;
  assign f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa107_y4 = f_s_dadda_pg_rca32_fa107_y4;
  assign f_s_dadda_pg_rca32_fa125_y0 = f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa109_y4 ^ f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa108_y4;
  assign f_s_dadda_pg_rca32_fa125_y1 = f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa109_y4 & f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa108_y4;
  assign f_s_dadda_pg_rca32_fa125_y2 = f_s_dadda_pg_rca32_fa125_y0 ^ f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa107_y4;
  assign f_s_dadda_pg_rca32_fa125_y3 = f_s_dadda_pg_rca32_fa125_y0 & f_s_dadda_pg_rca32_fa125_f_s_dadda_pg_rca32_fa107_y4;
  assign f_s_dadda_pg_rca32_fa125_y4 = f_s_dadda_pg_rca32_fa125_y1 | f_s_dadda_pg_rca32_fa125_y3;
  assign f_s_dadda_pg_rca32_and_21_0_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_21_0_y0 = f_s_dadda_pg_rca32_and_21_0_a_21 & f_s_dadda_pg_rca32_and_21_0_b_0;
  assign f_s_dadda_pg_rca32_and_20_1_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_20_1_y0 = f_s_dadda_pg_rca32_and_20_1_a_20 & f_s_dadda_pg_rca32_and_20_1_b_1;
  assign f_s_dadda_pg_rca32_and_19_2_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_19_2_y0 = f_s_dadda_pg_rca32_and_19_2_a_19 & f_s_dadda_pg_rca32_and_19_2_b_2;
  assign f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_21_0_y0 = f_s_dadda_pg_rca32_and_21_0_y0;
  assign f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_20_1_y0 = f_s_dadda_pg_rca32_and_20_1_y0;
  assign f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_19_2_y0 = f_s_dadda_pg_rca32_and_19_2_y0;
  assign f_s_dadda_pg_rca32_fa126_y0 = f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_21_0_y0 ^ f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_20_1_y0;
  assign f_s_dadda_pg_rca32_fa126_y1 = f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_21_0_y0 & f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_20_1_y0;
  assign f_s_dadda_pg_rca32_fa126_y2 = f_s_dadda_pg_rca32_fa126_y0 ^ f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_19_2_y0;
  assign f_s_dadda_pg_rca32_fa126_y3 = f_s_dadda_pg_rca32_fa126_y0 & f_s_dadda_pg_rca32_fa126_f_s_dadda_pg_rca32_and_19_2_y0;
  assign f_s_dadda_pg_rca32_fa126_y4 = f_s_dadda_pg_rca32_fa126_y1 | f_s_dadda_pg_rca32_fa126_y3;
  assign f_s_dadda_pg_rca32_and_18_3_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_18_3_y0 = f_s_dadda_pg_rca32_and_18_3_a_18 & f_s_dadda_pg_rca32_and_18_3_b_3;
  assign f_s_dadda_pg_rca32_and_17_4_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_17_4_y0 = f_s_dadda_pg_rca32_and_17_4_a_17 & f_s_dadda_pg_rca32_and_17_4_b_4;
  assign f_s_dadda_pg_rca32_and_16_5_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_16_5_y0 = f_s_dadda_pg_rca32_and_16_5_a_16 & f_s_dadda_pg_rca32_and_16_5_b_5;
  assign f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_18_3_y0 = f_s_dadda_pg_rca32_and_18_3_y0;
  assign f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_17_4_y0 = f_s_dadda_pg_rca32_and_17_4_y0;
  assign f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_16_5_y0 = f_s_dadda_pg_rca32_and_16_5_y0;
  assign f_s_dadda_pg_rca32_fa127_y0 = f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_18_3_y0 ^ f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_17_4_y0;
  assign f_s_dadda_pg_rca32_fa127_y1 = f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_18_3_y0 & f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_17_4_y0;
  assign f_s_dadda_pg_rca32_fa127_y2 = f_s_dadda_pg_rca32_fa127_y0 ^ f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_16_5_y0;
  assign f_s_dadda_pg_rca32_fa127_y3 = f_s_dadda_pg_rca32_fa127_y0 & f_s_dadda_pg_rca32_fa127_f_s_dadda_pg_rca32_and_16_5_y0;
  assign f_s_dadda_pg_rca32_fa127_y4 = f_s_dadda_pg_rca32_fa127_y1 | f_s_dadda_pg_rca32_fa127_y3;
  assign f_s_dadda_pg_rca32_and_15_6_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_15_6_y0 = f_s_dadda_pg_rca32_and_15_6_a_15 & f_s_dadda_pg_rca32_and_15_6_b_6;
  assign f_s_dadda_pg_rca32_and_14_7_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_14_7_y0 = f_s_dadda_pg_rca32_and_14_7_a_14 & f_s_dadda_pg_rca32_and_14_7_b_7;
  assign f_s_dadda_pg_rca32_and_13_8_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_13_8_y0 = f_s_dadda_pg_rca32_and_13_8_a_13 & f_s_dadda_pg_rca32_and_13_8_b_8;
  assign f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_15_6_y0 = f_s_dadda_pg_rca32_and_15_6_y0;
  assign f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_14_7_y0 = f_s_dadda_pg_rca32_and_14_7_y0;
  assign f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_13_8_y0 = f_s_dadda_pg_rca32_and_13_8_y0;
  assign f_s_dadda_pg_rca32_fa128_y0 = f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_15_6_y0 ^ f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_14_7_y0;
  assign f_s_dadda_pg_rca32_fa128_y1 = f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_15_6_y0 & f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_14_7_y0;
  assign f_s_dadda_pg_rca32_fa128_y2 = f_s_dadda_pg_rca32_fa128_y0 ^ f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_13_8_y0;
  assign f_s_dadda_pg_rca32_fa128_y3 = f_s_dadda_pg_rca32_fa128_y0 & f_s_dadda_pg_rca32_fa128_f_s_dadda_pg_rca32_and_13_8_y0;
  assign f_s_dadda_pg_rca32_fa128_y4 = f_s_dadda_pg_rca32_fa128_y1 | f_s_dadda_pg_rca32_fa128_y3;
  assign f_s_dadda_pg_rca32_and_12_9_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_12_9_y0 = f_s_dadda_pg_rca32_and_12_9_a_12 & f_s_dadda_pg_rca32_and_12_9_b_9;
  assign f_s_dadda_pg_rca32_and_11_10_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_11_10_y0 = f_s_dadda_pg_rca32_and_11_10_a_11 & f_s_dadda_pg_rca32_and_11_10_b_10;
  assign f_s_dadda_pg_rca32_and_10_11_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_10_11_y0 = f_s_dadda_pg_rca32_and_10_11_a_10 & f_s_dadda_pg_rca32_and_10_11_b_11;
  assign f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_12_9_y0 = f_s_dadda_pg_rca32_and_12_9_y0;
  assign f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_11_10_y0 = f_s_dadda_pg_rca32_and_11_10_y0;
  assign f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_10_11_y0 = f_s_dadda_pg_rca32_and_10_11_y0;
  assign f_s_dadda_pg_rca32_fa129_y0 = f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_12_9_y0 ^ f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_11_10_y0;
  assign f_s_dadda_pg_rca32_fa129_y1 = f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_12_9_y0 & f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_11_10_y0;
  assign f_s_dadda_pg_rca32_fa129_y2 = f_s_dadda_pg_rca32_fa129_y0 ^ f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_10_11_y0;
  assign f_s_dadda_pg_rca32_fa129_y3 = f_s_dadda_pg_rca32_fa129_y0 & f_s_dadda_pg_rca32_fa129_f_s_dadda_pg_rca32_and_10_11_y0;
  assign f_s_dadda_pg_rca32_fa129_y4 = f_s_dadda_pg_rca32_fa129_y1 | f_s_dadda_pg_rca32_fa129_y3;
  assign f_s_dadda_pg_rca32_and_9_12_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_9_12_y0 = f_s_dadda_pg_rca32_and_9_12_a_9 & f_s_dadda_pg_rca32_and_9_12_b_12;
  assign f_s_dadda_pg_rca32_and_8_13_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_8_13_y0 = f_s_dadda_pg_rca32_and_8_13_a_8 & f_s_dadda_pg_rca32_and_8_13_b_13;
  assign f_s_dadda_pg_rca32_and_7_14_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_7_14_y0 = f_s_dadda_pg_rca32_and_7_14_a_7 & f_s_dadda_pg_rca32_and_7_14_b_14;
  assign f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_9_12_y0 = f_s_dadda_pg_rca32_and_9_12_y0;
  assign f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_8_13_y0 = f_s_dadda_pg_rca32_and_8_13_y0;
  assign f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_7_14_y0 = f_s_dadda_pg_rca32_and_7_14_y0;
  assign f_s_dadda_pg_rca32_fa130_y0 = f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_9_12_y0 ^ f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_8_13_y0;
  assign f_s_dadda_pg_rca32_fa130_y1 = f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_9_12_y0 & f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_8_13_y0;
  assign f_s_dadda_pg_rca32_fa130_y2 = f_s_dadda_pg_rca32_fa130_y0 ^ f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_7_14_y0;
  assign f_s_dadda_pg_rca32_fa130_y3 = f_s_dadda_pg_rca32_fa130_y0 & f_s_dadda_pg_rca32_fa130_f_s_dadda_pg_rca32_and_7_14_y0;
  assign f_s_dadda_pg_rca32_fa130_y4 = f_s_dadda_pg_rca32_fa130_y1 | f_s_dadda_pg_rca32_fa130_y3;
  assign f_s_dadda_pg_rca32_and_6_15_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_6_15_y0 = f_s_dadda_pg_rca32_and_6_15_a_6 & f_s_dadda_pg_rca32_and_6_15_b_15;
  assign f_s_dadda_pg_rca32_and_5_16_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_5_16_y0 = f_s_dadda_pg_rca32_and_5_16_a_5 & f_s_dadda_pg_rca32_and_5_16_b_16;
  assign f_s_dadda_pg_rca32_and_4_17_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_4_17_y0 = f_s_dadda_pg_rca32_and_4_17_a_4 & f_s_dadda_pg_rca32_and_4_17_b_17;
  assign f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_6_15_y0 = f_s_dadda_pg_rca32_and_6_15_y0;
  assign f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_5_16_y0 = f_s_dadda_pg_rca32_and_5_16_y0;
  assign f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_4_17_y0 = f_s_dadda_pg_rca32_and_4_17_y0;
  assign f_s_dadda_pg_rca32_fa131_y0 = f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_6_15_y0 ^ f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_5_16_y0;
  assign f_s_dadda_pg_rca32_fa131_y1 = f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_6_15_y0 & f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_5_16_y0;
  assign f_s_dadda_pg_rca32_fa131_y2 = f_s_dadda_pg_rca32_fa131_y0 ^ f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_4_17_y0;
  assign f_s_dadda_pg_rca32_fa131_y3 = f_s_dadda_pg_rca32_fa131_y0 & f_s_dadda_pg_rca32_fa131_f_s_dadda_pg_rca32_and_4_17_y0;
  assign f_s_dadda_pg_rca32_fa131_y4 = f_s_dadda_pg_rca32_fa131_y1 | f_s_dadda_pg_rca32_fa131_y3;
  assign f_s_dadda_pg_rca32_and_3_18_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_3_18_y0 = f_s_dadda_pg_rca32_and_3_18_a_3 & f_s_dadda_pg_rca32_and_3_18_b_18;
  assign f_s_dadda_pg_rca32_and_2_19_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_2_19_y0 = f_s_dadda_pg_rca32_and_2_19_a_2 & f_s_dadda_pg_rca32_and_2_19_b_19;
  assign f_s_dadda_pg_rca32_and_1_20_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_1_20_y0 = f_s_dadda_pg_rca32_and_1_20_a_1 & f_s_dadda_pg_rca32_and_1_20_b_20;
  assign f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_3_18_y0 = f_s_dadda_pg_rca32_and_3_18_y0;
  assign f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_2_19_y0 = f_s_dadda_pg_rca32_and_2_19_y0;
  assign f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_1_20_y0 = f_s_dadda_pg_rca32_and_1_20_y0;
  assign f_s_dadda_pg_rca32_fa132_y0 = f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_3_18_y0 ^ f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_2_19_y0;
  assign f_s_dadda_pg_rca32_fa132_y1 = f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_3_18_y0 & f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_2_19_y0;
  assign f_s_dadda_pg_rca32_fa132_y2 = f_s_dadda_pg_rca32_fa132_y0 ^ f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_1_20_y0;
  assign f_s_dadda_pg_rca32_fa132_y3 = f_s_dadda_pg_rca32_fa132_y0 & f_s_dadda_pg_rca32_fa132_f_s_dadda_pg_rca32_and_1_20_y0;
  assign f_s_dadda_pg_rca32_fa132_y4 = f_s_dadda_pg_rca32_fa132_y1 | f_s_dadda_pg_rca32_fa132_y3;
  assign f_s_dadda_pg_rca32_and_0_21_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_0_21_y0 = f_s_dadda_pg_rca32_and_0_21_a_0 & f_s_dadda_pg_rca32_and_0_21_b_21;
  assign f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_and_0_21_y0 = f_s_dadda_pg_rca32_and_0_21_y0;
  assign f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_fa121_y2 = f_s_dadda_pg_rca32_fa121_y2;
  assign f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_fa122_y2 = f_s_dadda_pg_rca32_fa122_y2;
  assign f_s_dadda_pg_rca32_fa133_y0 = f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_and_0_21_y0 ^ f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_fa121_y2;
  assign f_s_dadda_pg_rca32_fa133_y1 = f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_and_0_21_y0 & f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_fa121_y2;
  assign f_s_dadda_pg_rca32_fa133_y2 = f_s_dadda_pg_rca32_fa133_y0 ^ f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_fa122_y2;
  assign f_s_dadda_pg_rca32_fa133_y3 = f_s_dadda_pg_rca32_fa133_y0 & f_s_dadda_pg_rca32_fa133_f_s_dadda_pg_rca32_fa122_y2;
  assign f_s_dadda_pg_rca32_fa133_y4 = f_s_dadda_pg_rca32_fa133_y1 | f_s_dadda_pg_rca32_fa133_y3;
  assign f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa123_y2 = f_s_dadda_pg_rca32_fa123_y2;
  assign f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa124_y2 = f_s_dadda_pg_rca32_fa124_y2;
  assign f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa125_y2 = f_s_dadda_pg_rca32_fa125_y2;
  assign f_s_dadda_pg_rca32_fa134_y0 = f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa123_y2 ^ f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa124_y2;
  assign f_s_dadda_pg_rca32_fa134_y1 = f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa123_y2 & f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa124_y2;
  assign f_s_dadda_pg_rca32_fa134_y2 = f_s_dadda_pg_rca32_fa134_y0 ^ f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa125_y2;
  assign f_s_dadda_pg_rca32_fa134_y3 = f_s_dadda_pg_rca32_fa134_y0 & f_s_dadda_pg_rca32_fa134_f_s_dadda_pg_rca32_fa125_y2;
  assign f_s_dadda_pg_rca32_fa134_y4 = f_s_dadda_pg_rca32_fa134_y1 | f_s_dadda_pg_rca32_fa134_y3;
  assign f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa126_y2 = f_s_dadda_pg_rca32_fa126_y2;
  assign f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa127_y2 = f_s_dadda_pg_rca32_fa127_y2;
  assign f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa128_y2 = f_s_dadda_pg_rca32_fa128_y2;
  assign f_s_dadda_pg_rca32_fa135_y0 = f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa126_y2 ^ f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa127_y2;
  assign f_s_dadda_pg_rca32_fa135_y1 = f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa126_y2 & f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa127_y2;
  assign f_s_dadda_pg_rca32_fa135_y2 = f_s_dadda_pg_rca32_fa135_y0 ^ f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa128_y2;
  assign f_s_dadda_pg_rca32_fa135_y3 = f_s_dadda_pg_rca32_fa135_y0 & f_s_dadda_pg_rca32_fa135_f_s_dadda_pg_rca32_fa128_y2;
  assign f_s_dadda_pg_rca32_fa135_y4 = f_s_dadda_pg_rca32_fa135_y1 | f_s_dadda_pg_rca32_fa135_y3;
  assign f_s_dadda_pg_rca32_ha19_f_s_dadda_pg_rca32_fa129_y2 = f_s_dadda_pg_rca32_fa129_y2;
  assign f_s_dadda_pg_rca32_ha19_f_s_dadda_pg_rca32_fa130_y2 = f_s_dadda_pg_rca32_fa130_y2;
  assign f_s_dadda_pg_rca32_ha19_y0 = f_s_dadda_pg_rca32_ha19_f_s_dadda_pg_rca32_fa129_y2 ^ f_s_dadda_pg_rca32_ha19_f_s_dadda_pg_rca32_fa130_y2;
  assign f_s_dadda_pg_rca32_ha19_y1 = f_s_dadda_pg_rca32_ha19_f_s_dadda_pg_rca32_fa129_y2 & f_s_dadda_pg_rca32_ha19_f_s_dadda_pg_rca32_fa130_y2;
  assign f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_ha19_y1 = f_s_dadda_pg_rca32_ha19_y1;
  assign f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_fa135_y4 = f_s_dadda_pg_rca32_fa135_y4;
  assign f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_fa134_y4 = f_s_dadda_pg_rca32_fa134_y4;
  assign f_s_dadda_pg_rca32_fa136_y0 = f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_ha19_y1 ^ f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_fa135_y4;
  assign f_s_dadda_pg_rca32_fa136_y1 = f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_ha19_y1 & f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_fa135_y4;
  assign f_s_dadda_pg_rca32_fa136_y2 = f_s_dadda_pg_rca32_fa136_y0 ^ f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_fa134_y4;
  assign f_s_dadda_pg_rca32_fa136_y3 = f_s_dadda_pg_rca32_fa136_y0 & f_s_dadda_pg_rca32_fa136_f_s_dadda_pg_rca32_fa134_y4;
  assign f_s_dadda_pg_rca32_fa136_y4 = f_s_dadda_pg_rca32_fa136_y1 | f_s_dadda_pg_rca32_fa136_y3;
  assign f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa133_y4 = f_s_dadda_pg_rca32_fa133_y4;
  assign f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa132_y4 = f_s_dadda_pg_rca32_fa132_y4;
  assign f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa131_y4 = f_s_dadda_pg_rca32_fa131_y4;
  assign f_s_dadda_pg_rca32_fa137_y0 = f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa133_y4 ^ f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa132_y4;
  assign f_s_dadda_pg_rca32_fa137_y1 = f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa133_y4 & f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa132_y4;
  assign f_s_dadda_pg_rca32_fa137_y2 = f_s_dadda_pg_rca32_fa137_y0 ^ f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa131_y4;
  assign f_s_dadda_pg_rca32_fa137_y3 = f_s_dadda_pg_rca32_fa137_y0 & f_s_dadda_pg_rca32_fa137_f_s_dadda_pg_rca32_fa131_y4;
  assign f_s_dadda_pg_rca32_fa137_y4 = f_s_dadda_pg_rca32_fa137_y1 | f_s_dadda_pg_rca32_fa137_y3;
  assign f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa130_y4 = f_s_dadda_pg_rca32_fa130_y4;
  assign f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa129_y4 = f_s_dadda_pg_rca32_fa129_y4;
  assign f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa128_y4 = f_s_dadda_pg_rca32_fa128_y4;
  assign f_s_dadda_pg_rca32_fa138_y0 = f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa130_y4 ^ f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa129_y4;
  assign f_s_dadda_pg_rca32_fa138_y1 = f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa130_y4 & f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa129_y4;
  assign f_s_dadda_pg_rca32_fa138_y2 = f_s_dadda_pg_rca32_fa138_y0 ^ f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa128_y4;
  assign f_s_dadda_pg_rca32_fa138_y3 = f_s_dadda_pg_rca32_fa138_y0 & f_s_dadda_pg_rca32_fa138_f_s_dadda_pg_rca32_fa128_y4;
  assign f_s_dadda_pg_rca32_fa138_y4 = f_s_dadda_pg_rca32_fa138_y1 | f_s_dadda_pg_rca32_fa138_y3;
  assign f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa127_y4 = f_s_dadda_pg_rca32_fa127_y4;
  assign f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa126_y4 = f_s_dadda_pg_rca32_fa126_y4;
  assign f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa125_y4 = f_s_dadda_pg_rca32_fa125_y4;
  assign f_s_dadda_pg_rca32_fa139_y0 = f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa127_y4 ^ f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa126_y4;
  assign f_s_dadda_pg_rca32_fa139_y1 = f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa127_y4 & f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa126_y4;
  assign f_s_dadda_pg_rca32_fa139_y2 = f_s_dadda_pg_rca32_fa139_y0 ^ f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa125_y4;
  assign f_s_dadda_pg_rca32_fa139_y3 = f_s_dadda_pg_rca32_fa139_y0 & f_s_dadda_pg_rca32_fa139_f_s_dadda_pg_rca32_fa125_y4;
  assign f_s_dadda_pg_rca32_fa139_y4 = f_s_dadda_pg_rca32_fa139_y1 | f_s_dadda_pg_rca32_fa139_y3;
  assign f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa124_y4 = f_s_dadda_pg_rca32_fa124_y4;
  assign f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa123_y4 = f_s_dadda_pg_rca32_fa123_y4;
  assign f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa122_y4 = f_s_dadda_pg_rca32_fa122_y4;
  assign f_s_dadda_pg_rca32_fa140_y0 = f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa124_y4 ^ f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa123_y4;
  assign f_s_dadda_pg_rca32_fa140_y1 = f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa124_y4 & f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa123_y4;
  assign f_s_dadda_pg_rca32_fa140_y2 = f_s_dadda_pg_rca32_fa140_y0 ^ f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa122_y4;
  assign f_s_dadda_pg_rca32_fa140_y3 = f_s_dadda_pg_rca32_fa140_y0 & f_s_dadda_pg_rca32_fa140_f_s_dadda_pg_rca32_fa122_y4;
  assign f_s_dadda_pg_rca32_fa140_y4 = f_s_dadda_pg_rca32_fa140_y1 | f_s_dadda_pg_rca32_fa140_y3;
  assign f_s_dadda_pg_rca32_and_22_0_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_22_0_y0 = f_s_dadda_pg_rca32_and_22_0_a_22 & f_s_dadda_pg_rca32_and_22_0_b_0;
  assign f_s_dadda_pg_rca32_and_21_1_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_21_1_y0 = f_s_dadda_pg_rca32_and_21_1_a_21 & f_s_dadda_pg_rca32_and_21_1_b_1;
  assign f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_fa121_y4 = f_s_dadda_pg_rca32_fa121_y4;
  assign f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_and_22_0_y0 = f_s_dadda_pg_rca32_and_22_0_y0;
  assign f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_and_21_1_y0 = f_s_dadda_pg_rca32_and_21_1_y0;
  assign f_s_dadda_pg_rca32_fa141_y0 = f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_fa121_y4 ^ f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_and_22_0_y0;
  assign f_s_dadda_pg_rca32_fa141_y1 = f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_fa121_y4 & f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_and_22_0_y0;
  assign f_s_dadda_pg_rca32_fa141_y2 = f_s_dadda_pg_rca32_fa141_y0 ^ f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_and_21_1_y0;
  assign f_s_dadda_pg_rca32_fa141_y3 = f_s_dadda_pg_rca32_fa141_y0 & f_s_dadda_pg_rca32_fa141_f_s_dadda_pg_rca32_and_21_1_y0;
  assign f_s_dadda_pg_rca32_fa141_y4 = f_s_dadda_pg_rca32_fa141_y1 | f_s_dadda_pg_rca32_fa141_y3;
  assign f_s_dadda_pg_rca32_and_20_2_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_20_2_y0 = f_s_dadda_pg_rca32_and_20_2_a_20 & f_s_dadda_pg_rca32_and_20_2_b_2;
  assign f_s_dadda_pg_rca32_and_19_3_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_19_3_y0 = f_s_dadda_pg_rca32_and_19_3_a_19 & f_s_dadda_pg_rca32_and_19_3_b_3;
  assign f_s_dadda_pg_rca32_and_18_4_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_18_4_y0 = f_s_dadda_pg_rca32_and_18_4_a_18 & f_s_dadda_pg_rca32_and_18_4_b_4;
  assign f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_20_2_y0 = f_s_dadda_pg_rca32_and_20_2_y0;
  assign f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_19_3_y0 = f_s_dadda_pg_rca32_and_19_3_y0;
  assign f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_18_4_y0 = f_s_dadda_pg_rca32_and_18_4_y0;
  assign f_s_dadda_pg_rca32_fa142_y0 = f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_20_2_y0 ^ f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_19_3_y0;
  assign f_s_dadda_pg_rca32_fa142_y1 = f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_20_2_y0 & f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_19_3_y0;
  assign f_s_dadda_pg_rca32_fa142_y2 = f_s_dadda_pg_rca32_fa142_y0 ^ f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_18_4_y0;
  assign f_s_dadda_pg_rca32_fa142_y3 = f_s_dadda_pg_rca32_fa142_y0 & f_s_dadda_pg_rca32_fa142_f_s_dadda_pg_rca32_and_18_4_y0;
  assign f_s_dadda_pg_rca32_fa142_y4 = f_s_dadda_pg_rca32_fa142_y1 | f_s_dadda_pg_rca32_fa142_y3;
  assign f_s_dadda_pg_rca32_and_17_5_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_17_5_y0 = f_s_dadda_pg_rca32_and_17_5_a_17 & f_s_dadda_pg_rca32_and_17_5_b_5;
  assign f_s_dadda_pg_rca32_and_16_6_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_16_6_y0 = f_s_dadda_pg_rca32_and_16_6_a_16 & f_s_dadda_pg_rca32_and_16_6_b_6;
  assign f_s_dadda_pg_rca32_and_15_7_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_15_7_y0 = f_s_dadda_pg_rca32_and_15_7_a_15 & f_s_dadda_pg_rca32_and_15_7_b_7;
  assign f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_17_5_y0 = f_s_dadda_pg_rca32_and_17_5_y0;
  assign f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_16_6_y0 = f_s_dadda_pg_rca32_and_16_6_y0;
  assign f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_15_7_y0 = f_s_dadda_pg_rca32_and_15_7_y0;
  assign f_s_dadda_pg_rca32_fa143_y0 = f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_17_5_y0 ^ f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_16_6_y0;
  assign f_s_dadda_pg_rca32_fa143_y1 = f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_17_5_y0 & f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_16_6_y0;
  assign f_s_dadda_pg_rca32_fa143_y2 = f_s_dadda_pg_rca32_fa143_y0 ^ f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_15_7_y0;
  assign f_s_dadda_pg_rca32_fa143_y3 = f_s_dadda_pg_rca32_fa143_y0 & f_s_dadda_pg_rca32_fa143_f_s_dadda_pg_rca32_and_15_7_y0;
  assign f_s_dadda_pg_rca32_fa143_y4 = f_s_dadda_pg_rca32_fa143_y1 | f_s_dadda_pg_rca32_fa143_y3;
  assign f_s_dadda_pg_rca32_and_14_8_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_14_8_y0 = f_s_dadda_pg_rca32_and_14_8_a_14 & f_s_dadda_pg_rca32_and_14_8_b_8;
  assign f_s_dadda_pg_rca32_and_13_9_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_13_9_y0 = f_s_dadda_pg_rca32_and_13_9_a_13 & f_s_dadda_pg_rca32_and_13_9_b_9;
  assign f_s_dadda_pg_rca32_and_12_10_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_12_10_y0 = f_s_dadda_pg_rca32_and_12_10_a_12 & f_s_dadda_pg_rca32_and_12_10_b_10;
  assign f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_14_8_y0 = f_s_dadda_pg_rca32_and_14_8_y0;
  assign f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_13_9_y0 = f_s_dadda_pg_rca32_and_13_9_y0;
  assign f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_12_10_y0 = f_s_dadda_pg_rca32_and_12_10_y0;
  assign f_s_dadda_pg_rca32_fa144_y0 = f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_14_8_y0 ^ f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_13_9_y0;
  assign f_s_dadda_pg_rca32_fa144_y1 = f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_14_8_y0 & f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_13_9_y0;
  assign f_s_dadda_pg_rca32_fa144_y2 = f_s_dadda_pg_rca32_fa144_y0 ^ f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_12_10_y0;
  assign f_s_dadda_pg_rca32_fa144_y3 = f_s_dadda_pg_rca32_fa144_y0 & f_s_dadda_pg_rca32_fa144_f_s_dadda_pg_rca32_and_12_10_y0;
  assign f_s_dadda_pg_rca32_fa144_y4 = f_s_dadda_pg_rca32_fa144_y1 | f_s_dadda_pg_rca32_fa144_y3;
  assign f_s_dadda_pg_rca32_and_11_11_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_11_11_y0 = f_s_dadda_pg_rca32_and_11_11_a_11 & f_s_dadda_pg_rca32_and_11_11_b_11;
  assign f_s_dadda_pg_rca32_and_10_12_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_10_12_y0 = f_s_dadda_pg_rca32_and_10_12_a_10 & f_s_dadda_pg_rca32_and_10_12_b_12;
  assign f_s_dadda_pg_rca32_and_9_13_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_9_13_y0 = f_s_dadda_pg_rca32_and_9_13_a_9 & f_s_dadda_pg_rca32_and_9_13_b_13;
  assign f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_11_11_y0 = f_s_dadda_pg_rca32_and_11_11_y0;
  assign f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_10_12_y0 = f_s_dadda_pg_rca32_and_10_12_y0;
  assign f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_9_13_y0 = f_s_dadda_pg_rca32_and_9_13_y0;
  assign f_s_dadda_pg_rca32_fa145_y0 = f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_11_11_y0 ^ f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_10_12_y0;
  assign f_s_dadda_pg_rca32_fa145_y1 = f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_11_11_y0 & f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_10_12_y0;
  assign f_s_dadda_pg_rca32_fa145_y2 = f_s_dadda_pg_rca32_fa145_y0 ^ f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_9_13_y0;
  assign f_s_dadda_pg_rca32_fa145_y3 = f_s_dadda_pg_rca32_fa145_y0 & f_s_dadda_pg_rca32_fa145_f_s_dadda_pg_rca32_and_9_13_y0;
  assign f_s_dadda_pg_rca32_fa145_y4 = f_s_dadda_pg_rca32_fa145_y1 | f_s_dadda_pg_rca32_fa145_y3;
  assign f_s_dadda_pg_rca32_and_8_14_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_8_14_y0 = f_s_dadda_pg_rca32_and_8_14_a_8 & f_s_dadda_pg_rca32_and_8_14_b_14;
  assign f_s_dadda_pg_rca32_and_7_15_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_7_15_y0 = f_s_dadda_pg_rca32_and_7_15_a_7 & f_s_dadda_pg_rca32_and_7_15_b_15;
  assign f_s_dadda_pg_rca32_and_6_16_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_6_16_y0 = f_s_dadda_pg_rca32_and_6_16_a_6 & f_s_dadda_pg_rca32_and_6_16_b_16;
  assign f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_8_14_y0 = f_s_dadda_pg_rca32_and_8_14_y0;
  assign f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_7_15_y0 = f_s_dadda_pg_rca32_and_7_15_y0;
  assign f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_6_16_y0 = f_s_dadda_pg_rca32_and_6_16_y0;
  assign f_s_dadda_pg_rca32_fa146_y0 = f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_8_14_y0 ^ f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_7_15_y0;
  assign f_s_dadda_pg_rca32_fa146_y1 = f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_8_14_y0 & f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_7_15_y0;
  assign f_s_dadda_pg_rca32_fa146_y2 = f_s_dadda_pg_rca32_fa146_y0 ^ f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_6_16_y0;
  assign f_s_dadda_pg_rca32_fa146_y3 = f_s_dadda_pg_rca32_fa146_y0 & f_s_dadda_pg_rca32_fa146_f_s_dadda_pg_rca32_and_6_16_y0;
  assign f_s_dadda_pg_rca32_fa146_y4 = f_s_dadda_pg_rca32_fa146_y1 | f_s_dadda_pg_rca32_fa146_y3;
  assign f_s_dadda_pg_rca32_and_5_17_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_5_17_y0 = f_s_dadda_pg_rca32_and_5_17_a_5 & f_s_dadda_pg_rca32_and_5_17_b_17;
  assign f_s_dadda_pg_rca32_and_4_18_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_4_18_y0 = f_s_dadda_pg_rca32_and_4_18_a_4 & f_s_dadda_pg_rca32_and_4_18_b_18;
  assign f_s_dadda_pg_rca32_and_3_19_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_3_19_y0 = f_s_dadda_pg_rca32_and_3_19_a_3 & f_s_dadda_pg_rca32_and_3_19_b_19;
  assign f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_5_17_y0 = f_s_dadda_pg_rca32_and_5_17_y0;
  assign f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_4_18_y0 = f_s_dadda_pg_rca32_and_4_18_y0;
  assign f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_3_19_y0 = f_s_dadda_pg_rca32_and_3_19_y0;
  assign f_s_dadda_pg_rca32_fa147_y0 = f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_5_17_y0 ^ f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_4_18_y0;
  assign f_s_dadda_pg_rca32_fa147_y1 = f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_5_17_y0 & f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_4_18_y0;
  assign f_s_dadda_pg_rca32_fa147_y2 = f_s_dadda_pg_rca32_fa147_y0 ^ f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_3_19_y0;
  assign f_s_dadda_pg_rca32_fa147_y3 = f_s_dadda_pg_rca32_fa147_y0 & f_s_dadda_pg_rca32_fa147_f_s_dadda_pg_rca32_and_3_19_y0;
  assign f_s_dadda_pg_rca32_fa147_y4 = f_s_dadda_pg_rca32_fa147_y1 | f_s_dadda_pg_rca32_fa147_y3;
  assign f_s_dadda_pg_rca32_and_2_20_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_2_20_y0 = f_s_dadda_pg_rca32_and_2_20_a_2 & f_s_dadda_pg_rca32_and_2_20_b_20;
  assign f_s_dadda_pg_rca32_and_1_21_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_1_21_y0 = f_s_dadda_pg_rca32_and_1_21_a_1 & f_s_dadda_pg_rca32_and_1_21_b_21;
  assign f_s_dadda_pg_rca32_and_0_22_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_0_22_y0 = f_s_dadda_pg_rca32_and_0_22_a_0 & f_s_dadda_pg_rca32_and_0_22_b_22;
  assign f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_2_20_y0 = f_s_dadda_pg_rca32_and_2_20_y0;
  assign f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_1_21_y0 = f_s_dadda_pg_rca32_and_1_21_y0;
  assign f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_0_22_y0 = f_s_dadda_pg_rca32_and_0_22_y0;
  assign f_s_dadda_pg_rca32_fa148_y0 = f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_2_20_y0 ^ f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_1_21_y0;
  assign f_s_dadda_pg_rca32_fa148_y1 = f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_2_20_y0 & f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_1_21_y0;
  assign f_s_dadda_pg_rca32_fa148_y2 = f_s_dadda_pg_rca32_fa148_y0 ^ f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_0_22_y0;
  assign f_s_dadda_pg_rca32_fa148_y3 = f_s_dadda_pg_rca32_fa148_y0 & f_s_dadda_pg_rca32_fa148_f_s_dadda_pg_rca32_and_0_22_y0;
  assign f_s_dadda_pg_rca32_fa148_y4 = f_s_dadda_pg_rca32_fa148_y1 | f_s_dadda_pg_rca32_fa148_y3;
  assign f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa136_y2 = f_s_dadda_pg_rca32_fa136_y2;
  assign f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa137_y2 = f_s_dadda_pg_rca32_fa137_y2;
  assign f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa138_y2 = f_s_dadda_pg_rca32_fa138_y2;
  assign f_s_dadda_pg_rca32_fa149_y0 = f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa136_y2 ^ f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa137_y2;
  assign f_s_dadda_pg_rca32_fa149_y1 = f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa136_y2 & f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa137_y2;
  assign f_s_dadda_pg_rca32_fa149_y2 = f_s_dadda_pg_rca32_fa149_y0 ^ f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa138_y2;
  assign f_s_dadda_pg_rca32_fa149_y3 = f_s_dadda_pg_rca32_fa149_y0 & f_s_dadda_pg_rca32_fa149_f_s_dadda_pg_rca32_fa138_y2;
  assign f_s_dadda_pg_rca32_fa149_y4 = f_s_dadda_pg_rca32_fa149_y1 | f_s_dadda_pg_rca32_fa149_y3;
  assign f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa139_y2 = f_s_dadda_pg_rca32_fa139_y2;
  assign f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa140_y2 = f_s_dadda_pg_rca32_fa140_y2;
  assign f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa141_y2 = f_s_dadda_pg_rca32_fa141_y2;
  assign f_s_dadda_pg_rca32_fa150_y0 = f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa139_y2 ^ f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa140_y2;
  assign f_s_dadda_pg_rca32_fa150_y1 = f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa139_y2 & f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa140_y2;
  assign f_s_dadda_pg_rca32_fa150_y2 = f_s_dadda_pg_rca32_fa150_y0 ^ f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa141_y2;
  assign f_s_dadda_pg_rca32_fa150_y3 = f_s_dadda_pg_rca32_fa150_y0 & f_s_dadda_pg_rca32_fa150_f_s_dadda_pg_rca32_fa141_y2;
  assign f_s_dadda_pg_rca32_fa150_y4 = f_s_dadda_pg_rca32_fa150_y1 | f_s_dadda_pg_rca32_fa150_y3;
  assign f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa142_y2 = f_s_dadda_pg_rca32_fa142_y2;
  assign f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa143_y2 = f_s_dadda_pg_rca32_fa143_y2;
  assign f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa144_y2 = f_s_dadda_pg_rca32_fa144_y2;
  assign f_s_dadda_pg_rca32_fa151_y0 = f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa142_y2 ^ f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa143_y2;
  assign f_s_dadda_pg_rca32_fa151_y1 = f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa142_y2 & f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa143_y2;
  assign f_s_dadda_pg_rca32_fa151_y2 = f_s_dadda_pg_rca32_fa151_y0 ^ f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa144_y2;
  assign f_s_dadda_pg_rca32_fa151_y3 = f_s_dadda_pg_rca32_fa151_y0 & f_s_dadda_pg_rca32_fa151_f_s_dadda_pg_rca32_fa144_y2;
  assign f_s_dadda_pg_rca32_fa151_y4 = f_s_dadda_pg_rca32_fa151_y1 | f_s_dadda_pg_rca32_fa151_y3;
  assign f_s_dadda_pg_rca32_ha20_f_s_dadda_pg_rca32_fa145_y2 = f_s_dadda_pg_rca32_fa145_y2;
  assign f_s_dadda_pg_rca32_ha20_f_s_dadda_pg_rca32_fa146_y2 = f_s_dadda_pg_rca32_fa146_y2;
  assign f_s_dadda_pg_rca32_ha20_y0 = f_s_dadda_pg_rca32_ha20_f_s_dadda_pg_rca32_fa145_y2 ^ f_s_dadda_pg_rca32_ha20_f_s_dadda_pg_rca32_fa146_y2;
  assign f_s_dadda_pg_rca32_ha20_y1 = f_s_dadda_pg_rca32_ha20_f_s_dadda_pg_rca32_fa145_y2 & f_s_dadda_pg_rca32_ha20_f_s_dadda_pg_rca32_fa146_y2;
  assign f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_ha20_y1 = f_s_dadda_pg_rca32_ha20_y1;
  assign f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_fa151_y4 = f_s_dadda_pg_rca32_fa151_y4;
  assign f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_fa150_y4 = f_s_dadda_pg_rca32_fa150_y4;
  assign f_s_dadda_pg_rca32_fa152_y0 = f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_ha20_y1 ^ f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_fa151_y4;
  assign f_s_dadda_pg_rca32_fa152_y1 = f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_ha20_y1 & f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_fa151_y4;
  assign f_s_dadda_pg_rca32_fa152_y2 = f_s_dadda_pg_rca32_fa152_y0 ^ f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_fa150_y4;
  assign f_s_dadda_pg_rca32_fa152_y3 = f_s_dadda_pg_rca32_fa152_y0 & f_s_dadda_pg_rca32_fa152_f_s_dadda_pg_rca32_fa150_y4;
  assign f_s_dadda_pg_rca32_fa152_y4 = f_s_dadda_pg_rca32_fa152_y1 | f_s_dadda_pg_rca32_fa152_y3;
  assign f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa149_y4 = f_s_dadda_pg_rca32_fa149_y4;
  assign f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa148_y4 = f_s_dadda_pg_rca32_fa148_y4;
  assign f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa147_y4 = f_s_dadda_pg_rca32_fa147_y4;
  assign f_s_dadda_pg_rca32_fa153_y0 = f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa149_y4 ^ f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa148_y4;
  assign f_s_dadda_pg_rca32_fa153_y1 = f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa149_y4 & f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa148_y4;
  assign f_s_dadda_pg_rca32_fa153_y2 = f_s_dadda_pg_rca32_fa153_y0 ^ f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa147_y4;
  assign f_s_dadda_pg_rca32_fa153_y3 = f_s_dadda_pg_rca32_fa153_y0 & f_s_dadda_pg_rca32_fa153_f_s_dadda_pg_rca32_fa147_y4;
  assign f_s_dadda_pg_rca32_fa153_y4 = f_s_dadda_pg_rca32_fa153_y1 | f_s_dadda_pg_rca32_fa153_y3;
  assign f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa146_y4 = f_s_dadda_pg_rca32_fa146_y4;
  assign f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa145_y4 = f_s_dadda_pg_rca32_fa145_y4;
  assign f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa144_y4 = f_s_dadda_pg_rca32_fa144_y4;
  assign f_s_dadda_pg_rca32_fa154_y0 = f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa146_y4 ^ f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa145_y4;
  assign f_s_dadda_pg_rca32_fa154_y1 = f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa146_y4 & f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa145_y4;
  assign f_s_dadda_pg_rca32_fa154_y2 = f_s_dadda_pg_rca32_fa154_y0 ^ f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa144_y4;
  assign f_s_dadda_pg_rca32_fa154_y3 = f_s_dadda_pg_rca32_fa154_y0 & f_s_dadda_pg_rca32_fa154_f_s_dadda_pg_rca32_fa144_y4;
  assign f_s_dadda_pg_rca32_fa154_y4 = f_s_dadda_pg_rca32_fa154_y1 | f_s_dadda_pg_rca32_fa154_y3;
  assign f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa143_y4 = f_s_dadda_pg_rca32_fa143_y4;
  assign f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa142_y4 = f_s_dadda_pg_rca32_fa142_y4;
  assign f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa141_y4 = f_s_dadda_pg_rca32_fa141_y4;
  assign f_s_dadda_pg_rca32_fa155_y0 = f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa143_y4 ^ f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa142_y4;
  assign f_s_dadda_pg_rca32_fa155_y1 = f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa143_y4 & f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa142_y4;
  assign f_s_dadda_pg_rca32_fa155_y2 = f_s_dadda_pg_rca32_fa155_y0 ^ f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa141_y4;
  assign f_s_dadda_pg_rca32_fa155_y3 = f_s_dadda_pg_rca32_fa155_y0 & f_s_dadda_pg_rca32_fa155_f_s_dadda_pg_rca32_fa141_y4;
  assign f_s_dadda_pg_rca32_fa155_y4 = f_s_dadda_pg_rca32_fa155_y1 | f_s_dadda_pg_rca32_fa155_y3;
  assign f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa140_y4 = f_s_dadda_pg_rca32_fa140_y4;
  assign f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa139_y4 = f_s_dadda_pg_rca32_fa139_y4;
  assign f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa138_y4 = f_s_dadda_pg_rca32_fa138_y4;
  assign f_s_dadda_pg_rca32_fa156_y0 = f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa140_y4 ^ f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa139_y4;
  assign f_s_dadda_pg_rca32_fa156_y1 = f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa140_y4 & f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa139_y4;
  assign f_s_dadda_pg_rca32_fa156_y2 = f_s_dadda_pg_rca32_fa156_y0 ^ f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa138_y4;
  assign f_s_dadda_pg_rca32_fa156_y3 = f_s_dadda_pg_rca32_fa156_y0 & f_s_dadda_pg_rca32_fa156_f_s_dadda_pg_rca32_fa138_y4;
  assign f_s_dadda_pg_rca32_fa156_y4 = f_s_dadda_pg_rca32_fa156_y1 | f_s_dadda_pg_rca32_fa156_y3;
  assign f_s_dadda_pg_rca32_and_23_0_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_23_0_y0 = f_s_dadda_pg_rca32_and_23_0_a_23 & f_s_dadda_pg_rca32_and_23_0_b_0;
  assign f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_fa137_y4 = f_s_dadda_pg_rca32_fa137_y4;
  assign f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_fa136_y4 = f_s_dadda_pg_rca32_fa136_y4;
  assign f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_and_23_0_y0 = f_s_dadda_pg_rca32_and_23_0_y0;
  assign f_s_dadda_pg_rca32_fa157_y0 = f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_fa137_y4 ^ f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_fa136_y4;
  assign f_s_dadda_pg_rca32_fa157_y1 = f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_fa137_y4 & f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_fa136_y4;
  assign f_s_dadda_pg_rca32_fa157_y2 = f_s_dadda_pg_rca32_fa157_y0 ^ f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_and_23_0_y0;
  assign f_s_dadda_pg_rca32_fa157_y3 = f_s_dadda_pg_rca32_fa157_y0 & f_s_dadda_pg_rca32_fa157_f_s_dadda_pg_rca32_and_23_0_y0;
  assign f_s_dadda_pg_rca32_fa157_y4 = f_s_dadda_pg_rca32_fa157_y1 | f_s_dadda_pg_rca32_fa157_y3;
  assign f_s_dadda_pg_rca32_and_22_1_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_22_1_y0 = f_s_dadda_pg_rca32_and_22_1_a_22 & f_s_dadda_pg_rca32_and_22_1_b_1;
  assign f_s_dadda_pg_rca32_and_21_2_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_21_2_y0 = f_s_dadda_pg_rca32_and_21_2_a_21 & f_s_dadda_pg_rca32_and_21_2_b_2;
  assign f_s_dadda_pg_rca32_and_20_3_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_20_3_y0 = f_s_dadda_pg_rca32_and_20_3_a_20 & f_s_dadda_pg_rca32_and_20_3_b_3;
  assign f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_22_1_y0 = f_s_dadda_pg_rca32_and_22_1_y0;
  assign f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_21_2_y0 = f_s_dadda_pg_rca32_and_21_2_y0;
  assign f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_20_3_y0 = f_s_dadda_pg_rca32_and_20_3_y0;
  assign f_s_dadda_pg_rca32_fa158_y0 = f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_22_1_y0 ^ f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_21_2_y0;
  assign f_s_dadda_pg_rca32_fa158_y1 = f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_22_1_y0 & f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_21_2_y0;
  assign f_s_dadda_pg_rca32_fa158_y2 = f_s_dadda_pg_rca32_fa158_y0 ^ f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_20_3_y0;
  assign f_s_dadda_pg_rca32_fa158_y3 = f_s_dadda_pg_rca32_fa158_y0 & f_s_dadda_pg_rca32_fa158_f_s_dadda_pg_rca32_and_20_3_y0;
  assign f_s_dadda_pg_rca32_fa158_y4 = f_s_dadda_pg_rca32_fa158_y1 | f_s_dadda_pg_rca32_fa158_y3;
  assign f_s_dadda_pg_rca32_and_19_4_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_19_4_y0 = f_s_dadda_pg_rca32_and_19_4_a_19 & f_s_dadda_pg_rca32_and_19_4_b_4;
  assign f_s_dadda_pg_rca32_and_18_5_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_18_5_y0 = f_s_dadda_pg_rca32_and_18_5_a_18 & f_s_dadda_pg_rca32_and_18_5_b_5;
  assign f_s_dadda_pg_rca32_and_17_6_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_17_6_y0 = f_s_dadda_pg_rca32_and_17_6_a_17 & f_s_dadda_pg_rca32_and_17_6_b_6;
  assign f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_19_4_y0 = f_s_dadda_pg_rca32_and_19_4_y0;
  assign f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_18_5_y0 = f_s_dadda_pg_rca32_and_18_5_y0;
  assign f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_17_6_y0 = f_s_dadda_pg_rca32_and_17_6_y0;
  assign f_s_dadda_pg_rca32_fa159_y0 = f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_19_4_y0 ^ f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_18_5_y0;
  assign f_s_dadda_pg_rca32_fa159_y1 = f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_19_4_y0 & f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_18_5_y0;
  assign f_s_dadda_pg_rca32_fa159_y2 = f_s_dadda_pg_rca32_fa159_y0 ^ f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_17_6_y0;
  assign f_s_dadda_pg_rca32_fa159_y3 = f_s_dadda_pg_rca32_fa159_y0 & f_s_dadda_pg_rca32_fa159_f_s_dadda_pg_rca32_and_17_6_y0;
  assign f_s_dadda_pg_rca32_fa159_y4 = f_s_dadda_pg_rca32_fa159_y1 | f_s_dadda_pg_rca32_fa159_y3;
  assign f_s_dadda_pg_rca32_and_16_7_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_16_7_y0 = f_s_dadda_pg_rca32_and_16_7_a_16 & f_s_dadda_pg_rca32_and_16_7_b_7;
  assign f_s_dadda_pg_rca32_and_15_8_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_15_8_y0 = f_s_dadda_pg_rca32_and_15_8_a_15 & f_s_dadda_pg_rca32_and_15_8_b_8;
  assign f_s_dadda_pg_rca32_and_14_9_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_14_9_y0 = f_s_dadda_pg_rca32_and_14_9_a_14 & f_s_dadda_pg_rca32_and_14_9_b_9;
  assign f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_16_7_y0 = f_s_dadda_pg_rca32_and_16_7_y0;
  assign f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_15_8_y0 = f_s_dadda_pg_rca32_and_15_8_y0;
  assign f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_14_9_y0 = f_s_dadda_pg_rca32_and_14_9_y0;
  assign f_s_dadda_pg_rca32_fa160_y0 = f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_16_7_y0 ^ f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_15_8_y0;
  assign f_s_dadda_pg_rca32_fa160_y1 = f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_16_7_y0 & f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_15_8_y0;
  assign f_s_dadda_pg_rca32_fa160_y2 = f_s_dadda_pg_rca32_fa160_y0 ^ f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_14_9_y0;
  assign f_s_dadda_pg_rca32_fa160_y3 = f_s_dadda_pg_rca32_fa160_y0 & f_s_dadda_pg_rca32_fa160_f_s_dadda_pg_rca32_and_14_9_y0;
  assign f_s_dadda_pg_rca32_fa160_y4 = f_s_dadda_pg_rca32_fa160_y1 | f_s_dadda_pg_rca32_fa160_y3;
  assign f_s_dadda_pg_rca32_and_13_10_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_13_10_y0 = f_s_dadda_pg_rca32_and_13_10_a_13 & f_s_dadda_pg_rca32_and_13_10_b_10;
  assign f_s_dadda_pg_rca32_and_12_11_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_12_11_y0 = f_s_dadda_pg_rca32_and_12_11_a_12 & f_s_dadda_pg_rca32_and_12_11_b_11;
  assign f_s_dadda_pg_rca32_and_11_12_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_11_12_y0 = f_s_dadda_pg_rca32_and_11_12_a_11 & f_s_dadda_pg_rca32_and_11_12_b_12;
  assign f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_13_10_y0 = f_s_dadda_pg_rca32_and_13_10_y0;
  assign f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_12_11_y0 = f_s_dadda_pg_rca32_and_12_11_y0;
  assign f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_11_12_y0 = f_s_dadda_pg_rca32_and_11_12_y0;
  assign f_s_dadda_pg_rca32_fa161_y0 = f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_13_10_y0 ^ f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_12_11_y0;
  assign f_s_dadda_pg_rca32_fa161_y1 = f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_13_10_y0 & f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_12_11_y0;
  assign f_s_dadda_pg_rca32_fa161_y2 = f_s_dadda_pg_rca32_fa161_y0 ^ f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_11_12_y0;
  assign f_s_dadda_pg_rca32_fa161_y3 = f_s_dadda_pg_rca32_fa161_y0 & f_s_dadda_pg_rca32_fa161_f_s_dadda_pg_rca32_and_11_12_y0;
  assign f_s_dadda_pg_rca32_fa161_y4 = f_s_dadda_pg_rca32_fa161_y1 | f_s_dadda_pg_rca32_fa161_y3;
  assign f_s_dadda_pg_rca32_and_10_13_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_10_13_y0 = f_s_dadda_pg_rca32_and_10_13_a_10 & f_s_dadda_pg_rca32_and_10_13_b_13;
  assign f_s_dadda_pg_rca32_and_9_14_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_9_14_y0 = f_s_dadda_pg_rca32_and_9_14_a_9 & f_s_dadda_pg_rca32_and_9_14_b_14;
  assign f_s_dadda_pg_rca32_and_8_15_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_8_15_y0 = f_s_dadda_pg_rca32_and_8_15_a_8 & f_s_dadda_pg_rca32_and_8_15_b_15;
  assign f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_10_13_y0 = f_s_dadda_pg_rca32_and_10_13_y0;
  assign f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_9_14_y0 = f_s_dadda_pg_rca32_and_9_14_y0;
  assign f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_8_15_y0 = f_s_dadda_pg_rca32_and_8_15_y0;
  assign f_s_dadda_pg_rca32_fa162_y0 = f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_10_13_y0 ^ f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_9_14_y0;
  assign f_s_dadda_pg_rca32_fa162_y1 = f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_10_13_y0 & f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_9_14_y0;
  assign f_s_dadda_pg_rca32_fa162_y2 = f_s_dadda_pg_rca32_fa162_y0 ^ f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_8_15_y0;
  assign f_s_dadda_pg_rca32_fa162_y3 = f_s_dadda_pg_rca32_fa162_y0 & f_s_dadda_pg_rca32_fa162_f_s_dadda_pg_rca32_and_8_15_y0;
  assign f_s_dadda_pg_rca32_fa162_y4 = f_s_dadda_pg_rca32_fa162_y1 | f_s_dadda_pg_rca32_fa162_y3;
  assign f_s_dadda_pg_rca32_and_7_16_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_7_16_y0 = f_s_dadda_pg_rca32_and_7_16_a_7 & f_s_dadda_pg_rca32_and_7_16_b_16;
  assign f_s_dadda_pg_rca32_and_6_17_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_6_17_y0 = f_s_dadda_pg_rca32_and_6_17_a_6 & f_s_dadda_pg_rca32_and_6_17_b_17;
  assign f_s_dadda_pg_rca32_and_5_18_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_5_18_y0 = f_s_dadda_pg_rca32_and_5_18_a_5 & f_s_dadda_pg_rca32_and_5_18_b_18;
  assign f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_7_16_y0 = f_s_dadda_pg_rca32_and_7_16_y0;
  assign f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_6_17_y0 = f_s_dadda_pg_rca32_and_6_17_y0;
  assign f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_5_18_y0 = f_s_dadda_pg_rca32_and_5_18_y0;
  assign f_s_dadda_pg_rca32_fa163_y0 = f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_7_16_y0 ^ f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_6_17_y0;
  assign f_s_dadda_pg_rca32_fa163_y1 = f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_7_16_y0 & f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_6_17_y0;
  assign f_s_dadda_pg_rca32_fa163_y2 = f_s_dadda_pg_rca32_fa163_y0 ^ f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_5_18_y0;
  assign f_s_dadda_pg_rca32_fa163_y3 = f_s_dadda_pg_rca32_fa163_y0 & f_s_dadda_pg_rca32_fa163_f_s_dadda_pg_rca32_and_5_18_y0;
  assign f_s_dadda_pg_rca32_fa163_y4 = f_s_dadda_pg_rca32_fa163_y1 | f_s_dadda_pg_rca32_fa163_y3;
  assign f_s_dadda_pg_rca32_and_4_19_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_4_19_y0 = f_s_dadda_pg_rca32_and_4_19_a_4 & f_s_dadda_pg_rca32_and_4_19_b_19;
  assign f_s_dadda_pg_rca32_and_3_20_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_3_20_y0 = f_s_dadda_pg_rca32_and_3_20_a_3 & f_s_dadda_pg_rca32_and_3_20_b_20;
  assign f_s_dadda_pg_rca32_and_2_21_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_2_21_y0 = f_s_dadda_pg_rca32_and_2_21_a_2 & f_s_dadda_pg_rca32_and_2_21_b_21;
  assign f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_4_19_y0 = f_s_dadda_pg_rca32_and_4_19_y0;
  assign f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_3_20_y0 = f_s_dadda_pg_rca32_and_3_20_y0;
  assign f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_2_21_y0 = f_s_dadda_pg_rca32_and_2_21_y0;
  assign f_s_dadda_pg_rca32_fa164_y0 = f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_4_19_y0 ^ f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_3_20_y0;
  assign f_s_dadda_pg_rca32_fa164_y1 = f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_4_19_y0 & f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_3_20_y0;
  assign f_s_dadda_pg_rca32_fa164_y2 = f_s_dadda_pg_rca32_fa164_y0 ^ f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_2_21_y0;
  assign f_s_dadda_pg_rca32_fa164_y3 = f_s_dadda_pg_rca32_fa164_y0 & f_s_dadda_pg_rca32_fa164_f_s_dadda_pg_rca32_and_2_21_y0;
  assign f_s_dadda_pg_rca32_fa164_y4 = f_s_dadda_pg_rca32_fa164_y1 | f_s_dadda_pg_rca32_fa164_y3;
  assign f_s_dadda_pg_rca32_and_1_22_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_1_22_y0 = f_s_dadda_pg_rca32_and_1_22_a_1 & f_s_dadda_pg_rca32_and_1_22_b_22;
  assign f_s_dadda_pg_rca32_and_0_23_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_0_23_y0 = f_s_dadda_pg_rca32_and_0_23_a_0 & f_s_dadda_pg_rca32_and_0_23_b_23;
  assign f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_and_1_22_y0 = f_s_dadda_pg_rca32_and_1_22_y0;
  assign f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_and_0_23_y0 = f_s_dadda_pg_rca32_and_0_23_y0;
  assign f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_fa152_y2 = f_s_dadda_pg_rca32_fa152_y2;
  assign f_s_dadda_pg_rca32_fa165_y0 = f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_and_1_22_y0 ^ f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_and_0_23_y0;
  assign f_s_dadda_pg_rca32_fa165_y1 = f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_and_1_22_y0 & f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_and_0_23_y0;
  assign f_s_dadda_pg_rca32_fa165_y2 = f_s_dadda_pg_rca32_fa165_y0 ^ f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_fa152_y2;
  assign f_s_dadda_pg_rca32_fa165_y3 = f_s_dadda_pg_rca32_fa165_y0 & f_s_dadda_pg_rca32_fa165_f_s_dadda_pg_rca32_fa152_y2;
  assign f_s_dadda_pg_rca32_fa165_y4 = f_s_dadda_pg_rca32_fa165_y1 | f_s_dadda_pg_rca32_fa165_y3;
  assign f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa153_y2 = f_s_dadda_pg_rca32_fa153_y2;
  assign f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa154_y2 = f_s_dadda_pg_rca32_fa154_y2;
  assign f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa155_y2 = f_s_dadda_pg_rca32_fa155_y2;
  assign f_s_dadda_pg_rca32_fa166_y0 = f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa153_y2 ^ f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa154_y2;
  assign f_s_dadda_pg_rca32_fa166_y1 = f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa153_y2 & f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa154_y2;
  assign f_s_dadda_pg_rca32_fa166_y2 = f_s_dadda_pg_rca32_fa166_y0 ^ f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa155_y2;
  assign f_s_dadda_pg_rca32_fa166_y3 = f_s_dadda_pg_rca32_fa166_y0 & f_s_dadda_pg_rca32_fa166_f_s_dadda_pg_rca32_fa155_y2;
  assign f_s_dadda_pg_rca32_fa166_y4 = f_s_dadda_pg_rca32_fa166_y1 | f_s_dadda_pg_rca32_fa166_y3;
  assign f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa156_y2 = f_s_dadda_pg_rca32_fa156_y2;
  assign f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa157_y2 = f_s_dadda_pg_rca32_fa157_y2;
  assign f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa158_y2 = f_s_dadda_pg_rca32_fa158_y2;
  assign f_s_dadda_pg_rca32_fa167_y0 = f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa156_y2 ^ f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa157_y2;
  assign f_s_dadda_pg_rca32_fa167_y1 = f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa156_y2 & f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa157_y2;
  assign f_s_dadda_pg_rca32_fa167_y2 = f_s_dadda_pg_rca32_fa167_y0 ^ f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa158_y2;
  assign f_s_dadda_pg_rca32_fa167_y3 = f_s_dadda_pg_rca32_fa167_y0 & f_s_dadda_pg_rca32_fa167_f_s_dadda_pg_rca32_fa158_y2;
  assign f_s_dadda_pg_rca32_fa167_y4 = f_s_dadda_pg_rca32_fa167_y1 | f_s_dadda_pg_rca32_fa167_y3;
  assign f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa159_y2 = f_s_dadda_pg_rca32_fa159_y2;
  assign f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa160_y2 = f_s_dadda_pg_rca32_fa160_y2;
  assign f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa161_y2 = f_s_dadda_pg_rca32_fa161_y2;
  assign f_s_dadda_pg_rca32_fa168_y0 = f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa159_y2 ^ f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa160_y2;
  assign f_s_dadda_pg_rca32_fa168_y1 = f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa159_y2 & f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa160_y2;
  assign f_s_dadda_pg_rca32_fa168_y2 = f_s_dadda_pg_rca32_fa168_y0 ^ f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa161_y2;
  assign f_s_dadda_pg_rca32_fa168_y3 = f_s_dadda_pg_rca32_fa168_y0 & f_s_dadda_pg_rca32_fa168_f_s_dadda_pg_rca32_fa161_y2;
  assign f_s_dadda_pg_rca32_fa168_y4 = f_s_dadda_pg_rca32_fa168_y1 | f_s_dadda_pg_rca32_fa168_y3;
  assign f_s_dadda_pg_rca32_ha21_f_s_dadda_pg_rca32_fa162_y2 = f_s_dadda_pg_rca32_fa162_y2;
  assign f_s_dadda_pg_rca32_ha21_f_s_dadda_pg_rca32_fa163_y2 = f_s_dadda_pg_rca32_fa163_y2;
  assign f_s_dadda_pg_rca32_ha21_y0 = f_s_dadda_pg_rca32_ha21_f_s_dadda_pg_rca32_fa162_y2 ^ f_s_dadda_pg_rca32_ha21_f_s_dadda_pg_rca32_fa163_y2;
  assign f_s_dadda_pg_rca32_ha21_y1 = f_s_dadda_pg_rca32_ha21_f_s_dadda_pg_rca32_fa162_y2 & f_s_dadda_pg_rca32_ha21_f_s_dadda_pg_rca32_fa163_y2;
  assign f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_ha21_y1 = f_s_dadda_pg_rca32_ha21_y1;
  assign f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_fa168_y4 = f_s_dadda_pg_rca32_fa168_y4;
  assign f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_fa167_y4 = f_s_dadda_pg_rca32_fa167_y4;
  assign f_s_dadda_pg_rca32_fa169_y0 = f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_ha21_y1 ^ f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_fa168_y4;
  assign f_s_dadda_pg_rca32_fa169_y1 = f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_ha21_y1 & f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_fa168_y4;
  assign f_s_dadda_pg_rca32_fa169_y2 = f_s_dadda_pg_rca32_fa169_y0 ^ f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_fa167_y4;
  assign f_s_dadda_pg_rca32_fa169_y3 = f_s_dadda_pg_rca32_fa169_y0 & f_s_dadda_pg_rca32_fa169_f_s_dadda_pg_rca32_fa167_y4;
  assign f_s_dadda_pg_rca32_fa169_y4 = f_s_dadda_pg_rca32_fa169_y1 | f_s_dadda_pg_rca32_fa169_y3;
  assign f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa166_y4 = f_s_dadda_pg_rca32_fa166_y4;
  assign f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa165_y4 = f_s_dadda_pg_rca32_fa165_y4;
  assign f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa164_y4 = f_s_dadda_pg_rca32_fa164_y4;
  assign f_s_dadda_pg_rca32_fa170_y0 = f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa166_y4 ^ f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa165_y4;
  assign f_s_dadda_pg_rca32_fa170_y1 = f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa166_y4 & f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa165_y4;
  assign f_s_dadda_pg_rca32_fa170_y2 = f_s_dadda_pg_rca32_fa170_y0 ^ f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa164_y4;
  assign f_s_dadda_pg_rca32_fa170_y3 = f_s_dadda_pg_rca32_fa170_y0 & f_s_dadda_pg_rca32_fa170_f_s_dadda_pg_rca32_fa164_y4;
  assign f_s_dadda_pg_rca32_fa170_y4 = f_s_dadda_pg_rca32_fa170_y1 | f_s_dadda_pg_rca32_fa170_y3;
  assign f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa163_y4 = f_s_dadda_pg_rca32_fa163_y4;
  assign f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa162_y4 = f_s_dadda_pg_rca32_fa162_y4;
  assign f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa161_y4 = f_s_dadda_pg_rca32_fa161_y4;
  assign f_s_dadda_pg_rca32_fa171_y0 = f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa163_y4 ^ f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa162_y4;
  assign f_s_dadda_pg_rca32_fa171_y1 = f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa163_y4 & f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa162_y4;
  assign f_s_dadda_pg_rca32_fa171_y2 = f_s_dadda_pg_rca32_fa171_y0 ^ f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa161_y4;
  assign f_s_dadda_pg_rca32_fa171_y3 = f_s_dadda_pg_rca32_fa171_y0 & f_s_dadda_pg_rca32_fa171_f_s_dadda_pg_rca32_fa161_y4;
  assign f_s_dadda_pg_rca32_fa171_y4 = f_s_dadda_pg_rca32_fa171_y1 | f_s_dadda_pg_rca32_fa171_y3;
  assign f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa160_y4 = f_s_dadda_pg_rca32_fa160_y4;
  assign f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa159_y4 = f_s_dadda_pg_rca32_fa159_y4;
  assign f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa158_y4 = f_s_dadda_pg_rca32_fa158_y4;
  assign f_s_dadda_pg_rca32_fa172_y0 = f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa160_y4 ^ f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa159_y4;
  assign f_s_dadda_pg_rca32_fa172_y1 = f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa160_y4 & f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa159_y4;
  assign f_s_dadda_pg_rca32_fa172_y2 = f_s_dadda_pg_rca32_fa172_y0 ^ f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa158_y4;
  assign f_s_dadda_pg_rca32_fa172_y3 = f_s_dadda_pg_rca32_fa172_y0 & f_s_dadda_pg_rca32_fa172_f_s_dadda_pg_rca32_fa158_y4;
  assign f_s_dadda_pg_rca32_fa172_y4 = f_s_dadda_pg_rca32_fa172_y1 | f_s_dadda_pg_rca32_fa172_y3;
  assign f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa157_y4 = f_s_dadda_pg_rca32_fa157_y4;
  assign f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa156_y4 = f_s_dadda_pg_rca32_fa156_y4;
  assign f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa155_y4 = f_s_dadda_pg_rca32_fa155_y4;
  assign f_s_dadda_pg_rca32_fa173_y0 = f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa157_y4 ^ f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa156_y4;
  assign f_s_dadda_pg_rca32_fa173_y1 = f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa157_y4 & f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa156_y4;
  assign f_s_dadda_pg_rca32_fa173_y2 = f_s_dadda_pg_rca32_fa173_y0 ^ f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa155_y4;
  assign f_s_dadda_pg_rca32_fa173_y3 = f_s_dadda_pg_rca32_fa173_y0 & f_s_dadda_pg_rca32_fa173_f_s_dadda_pg_rca32_fa155_y4;
  assign f_s_dadda_pg_rca32_fa173_y4 = f_s_dadda_pg_rca32_fa173_y1 | f_s_dadda_pg_rca32_fa173_y3;
  assign f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa154_y4 = f_s_dadda_pg_rca32_fa154_y4;
  assign f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa153_y4 = f_s_dadda_pg_rca32_fa153_y4;
  assign f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa152_y4 = f_s_dadda_pg_rca32_fa152_y4;
  assign f_s_dadda_pg_rca32_fa174_y0 = f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa154_y4 ^ f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa153_y4;
  assign f_s_dadda_pg_rca32_fa174_y1 = f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa154_y4 & f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa153_y4;
  assign f_s_dadda_pg_rca32_fa174_y2 = f_s_dadda_pg_rca32_fa174_y0 ^ f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa152_y4;
  assign f_s_dadda_pg_rca32_fa174_y3 = f_s_dadda_pg_rca32_fa174_y0 & f_s_dadda_pg_rca32_fa174_f_s_dadda_pg_rca32_fa152_y4;
  assign f_s_dadda_pg_rca32_fa174_y4 = f_s_dadda_pg_rca32_fa174_y1 | f_s_dadda_pg_rca32_fa174_y3;
  assign f_s_dadda_pg_rca32_and_24_0_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_24_0_y0 = f_s_dadda_pg_rca32_and_24_0_a_24 & f_s_dadda_pg_rca32_and_24_0_b_0;
  assign f_s_dadda_pg_rca32_and_23_1_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_23_1_y0 = f_s_dadda_pg_rca32_and_23_1_a_23 & f_s_dadda_pg_rca32_and_23_1_b_1;
  assign f_s_dadda_pg_rca32_and_22_2_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_22_2_y0 = f_s_dadda_pg_rca32_and_22_2_a_22 & f_s_dadda_pg_rca32_and_22_2_b_2;
  assign f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_24_0_y0 = f_s_dadda_pg_rca32_and_24_0_y0;
  assign f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_23_1_y0 = f_s_dadda_pg_rca32_and_23_1_y0;
  assign f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_22_2_y0 = f_s_dadda_pg_rca32_and_22_2_y0;
  assign f_s_dadda_pg_rca32_fa175_y0 = f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_24_0_y0 ^ f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_23_1_y0;
  assign f_s_dadda_pg_rca32_fa175_y1 = f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_24_0_y0 & f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_23_1_y0;
  assign f_s_dadda_pg_rca32_fa175_y2 = f_s_dadda_pg_rca32_fa175_y0 ^ f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_22_2_y0;
  assign f_s_dadda_pg_rca32_fa175_y3 = f_s_dadda_pg_rca32_fa175_y0 & f_s_dadda_pg_rca32_fa175_f_s_dadda_pg_rca32_and_22_2_y0;
  assign f_s_dadda_pg_rca32_fa175_y4 = f_s_dadda_pg_rca32_fa175_y1 | f_s_dadda_pg_rca32_fa175_y3;
  assign f_s_dadda_pg_rca32_and_21_3_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_21_3_y0 = f_s_dadda_pg_rca32_and_21_3_a_21 & f_s_dadda_pg_rca32_and_21_3_b_3;
  assign f_s_dadda_pg_rca32_and_20_4_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_20_4_y0 = f_s_dadda_pg_rca32_and_20_4_a_20 & f_s_dadda_pg_rca32_and_20_4_b_4;
  assign f_s_dadda_pg_rca32_and_19_5_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_19_5_y0 = f_s_dadda_pg_rca32_and_19_5_a_19 & f_s_dadda_pg_rca32_and_19_5_b_5;
  assign f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_21_3_y0 = f_s_dadda_pg_rca32_and_21_3_y0;
  assign f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_20_4_y0 = f_s_dadda_pg_rca32_and_20_4_y0;
  assign f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_19_5_y0 = f_s_dadda_pg_rca32_and_19_5_y0;
  assign f_s_dadda_pg_rca32_fa176_y0 = f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_21_3_y0 ^ f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_20_4_y0;
  assign f_s_dadda_pg_rca32_fa176_y1 = f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_21_3_y0 & f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_20_4_y0;
  assign f_s_dadda_pg_rca32_fa176_y2 = f_s_dadda_pg_rca32_fa176_y0 ^ f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_19_5_y0;
  assign f_s_dadda_pg_rca32_fa176_y3 = f_s_dadda_pg_rca32_fa176_y0 & f_s_dadda_pg_rca32_fa176_f_s_dadda_pg_rca32_and_19_5_y0;
  assign f_s_dadda_pg_rca32_fa176_y4 = f_s_dadda_pg_rca32_fa176_y1 | f_s_dadda_pg_rca32_fa176_y3;
  assign f_s_dadda_pg_rca32_and_18_6_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_18_6_y0 = f_s_dadda_pg_rca32_and_18_6_a_18 & f_s_dadda_pg_rca32_and_18_6_b_6;
  assign f_s_dadda_pg_rca32_and_17_7_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_17_7_y0 = f_s_dadda_pg_rca32_and_17_7_a_17 & f_s_dadda_pg_rca32_and_17_7_b_7;
  assign f_s_dadda_pg_rca32_and_16_8_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_16_8_y0 = f_s_dadda_pg_rca32_and_16_8_a_16 & f_s_dadda_pg_rca32_and_16_8_b_8;
  assign f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_18_6_y0 = f_s_dadda_pg_rca32_and_18_6_y0;
  assign f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_17_7_y0 = f_s_dadda_pg_rca32_and_17_7_y0;
  assign f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_16_8_y0 = f_s_dadda_pg_rca32_and_16_8_y0;
  assign f_s_dadda_pg_rca32_fa177_y0 = f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_18_6_y0 ^ f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_17_7_y0;
  assign f_s_dadda_pg_rca32_fa177_y1 = f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_18_6_y0 & f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_17_7_y0;
  assign f_s_dadda_pg_rca32_fa177_y2 = f_s_dadda_pg_rca32_fa177_y0 ^ f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_16_8_y0;
  assign f_s_dadda_pg_rca32_fa177_y3 = f_s_dadda_pg_rca32_fa177_y0 & f_s_dadda_pg_rca32_fa177_f_s_dadda_pg_rca32_and_16_8_y0;
  assign f_s_dadda_pg_rca32_fa177_y4 = f_s_dadda_pg_rca32_fa177_y1 | f_s_dadda_pg_rca32_fa177_y3;
  assign f_s_dadda_pg_rca32_and_15_9_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_15_9_y0 = f_s_dadda_pg_rca32_and_15_9_a_15 & f_s_dadda_pg_rca32_and_15_9_b_9;
  assign f_s_dadda_pg_rca32_and_14_10_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_14_10_y0 = f_s_dadda_pg_rca32_and_14_10_a_14 & f_s_dadda_pg_rca32_and_14_10_b_10;
  assign f_s_dadda_pg_rca32_and_13_11_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_13_11_y0 = f_s_dadda_pg_rca32_and_13_11_a_13 & f_s_dadda_pg_rca32_and_13_11_b_11;
  assign f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_15_9_y0 = f_s_dadda_pg_rca32_and_15_9_y0;
  assign f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_14_10_y0 = f_s_dadda_pg_rca32_and_14_10_y0;
  assign f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_13_11_y0 = f_s_dadda_pg_rca32_and_13_11_y0;
  assign f_s_dadda_pg_rca32_fa178_y0 = f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_15_9_y0 ^ f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_14_10_y0;
  assign f_s_dadda_pg_rca32_fa178_y1 = f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_15_9_y0 & f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_14_10_y0;
  assign f_s_dadda_pg_rca32_fa178_y2 = f_s_dadda_pg_rca32_fa178_y0 ^ f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_13_11_y0;
  assign f_s_dadda_pg_rca32_fa178_y3 = f_s_dadda_pg_rca32_fa178_y0 & f_s_dadda_pg_rca32_fa178_f_s_dadda_pg_rca32_and_13_11_y0;
  assign f_s_dadda_pg_rca32_fa178_y4 = f_s_dadda_pg_rca32_fa178_y1 | f_s_dadda_pg_rca32_fa178_y3;
  assign f_s_dadda_pg_rca32_and_12_12_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_12_12_y0 = f_s_dadda_pg_rca32_and_12_12_a_12 & f_s_dadda_pg_rca32_and_12_12_b_12;
  assign f_s_dadda_pg_rca32_and_11_13_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_11_13_y0 = f_s_dadda_pg_rca32_and_11_13_a_11 & f_s_dadda_pg_rca32_and_11_13_b_13;
  assign f_s_dadda_pg_rca32_and_10_14_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_10_14_y0 = f_s_dadda_pg_rca32_and_10_14_a_10 & f_s_dadda_pg_rca32_and_10_14_b_14;
  assign f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_12_12_y0 = f_s_dadda_pg_rca32_and_12_12_y0;
  assign f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_11_13_y0 = f_s_dadda_pg_rca32_and_11_13_y0;
  assign f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_10_14_y0 = f_s_dadda_pg_rca32_and_10_14_y0;
  assign f_s_dadda_pg_rca32_fa179_y0 = f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_12_12_y0 ^ f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_11_13_y0;
  assign f_s_dadda_pg_rca32_fa179_y1 = f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_12_12_y0 & f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_11_13_y0;
  assign f_s_dadda_pg_rca32_fa179_y2 = f_s_dadda_pg_rca32_fa179_y0 ^ f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_10_14_y0;
  assign f_s_dadda_pg_rca32_fa179_y3 = f_s_dadda_pg_rca32_fa179_y0 & f_s_dadda_pg_rca32_fa179_f_s_dadda_pg_rca32_and_10_14_y0;
  assign f_s_dadda_pg_rca32_fa179_y4 = f_s_dadda_pg_rca32_fa179_y1 | f_s_dadda_pg_rca32_fa179_y3;
  assign f_s_dadda_pg_rca32_and_9_15_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_9_15_y0 = f_s_dadda_pg_rca32_and_9_15_a_9 & f_s_dadda_pg_rca32_and_9_15_b_15;
  assign f_s_dadda_pg_rca32_and_8_16_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_8_16_y0 = f_s_dadda_pg_rca32_and_8_16_a_8 & f_s_dadda_pg_rca32_and_8_16_b_16;
  assign f_s_dadda_pg_rca32_and_7_17_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_7_17_y0 = f_s_dadda_pg_rca32_and_7_17_a_7 & f_s_dadda_pg_rca32_and_7_17_b_17;
  assign f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_9_15_y0 = f_s_dadda_pg_rca32_and_9_15_y0;
  assign f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_8_16_y0 = f_s_dadda_pg_rca32_and_8_16_y0;
  assign f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_7_17_y0 = f_s_dadda_pg_rca32_and_7_17_y0;
  assign f_s_dadda_pg_rca32_fa180_y0 = f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_9_15_y0 ^ f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_8_16_y0;
  assign f_s_dadda_pg_rca32_fa180_y1 = f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_9_15_y0 & f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_8_16_y0;
  assign f_s_dadda_pg_rca32_fa180_y2 = f_s_dadda_pg_rca32_fa180_y0 ^ f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_7_17_y0;
  assign f_s_dadda_pg_rca32_fa180_y3 = f_s_dadda_pg_rca32_fa180_y0 & f_s_dadda_pg_rca32_fa180_f_s_dadda_pg_rca32_and_7_17_y0;
  assign f_s_dadda_pg_rca32_fa180_y4 = f_s_dadda_pg_rca32_fa180_y1 | f_s_dadda_pg_rca32_fa180_y3;
  assign f_s_dadda_pg_rca32_and_6_18_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_6_18_y0 = f_s_dadda_pg_rca32_and_6_18_a_6 & f_s_dadda_pg_rca32_and_6_18_b_18;
  assign f_s_dadda_pg_rca32_and_5_19_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_5_19_y0 = f_s_dadda_pg_rca32_and_5_19_a_5 & f_s_dadda_pg_rca32_and_5_19_b_19;
  assign f_s_dadda_pg_rca32_and_4_20_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_4_20_y0 = f_s_dadda_pg_rca32_and_4_20_a_4 & f_s_dadda_pg_rca32_and_4_20_b_20;
  assign f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_6_18_y0 = f_s_dadda_pg_rca32_and_6_18_y0;
  assign f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_5_19_y0 = f_s_dadda_pg_rca32_and_5_19_y0;
  assign f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_4_20_y0 = f_s_dadda_pg_rca32_and_4_20_y0;
  assign f_s_dadda_pg_rca32_fa181_y0 = f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_6_18_y0 ^ f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_5_19_y0;
  assign f_s_dadda_pg_rca32_fa181_y1 = f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_6_18_y0 & f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_5_19_y0;
  assign f_s_dadda_pg_rca32_fa181_y2 = f_s_dadda_pg_rca32_fa181_y0 ^ f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_4_20_y0;
  assign f_s_dadda_pg_rca32_fa181_y3 = f_s_dadda_pg_rca32_fa181_y0 & f_s_dadda_pg_rca32_fa181_f_s_dadda_pg_rca32_and_4_20_y0;
  assign f_s_dadda_pg_rca32_fa181_y4 = f_s_dadda_pg_rca32_fa181_y1 | f_s_dadda_pg_rca32_fa181_y3;
  assign f_s_dadda_pg_rca32_and_3_21_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_3_21_y0 = f_s_dadda_pg_rca32_and_3_21_a_3 & f_s_dadda_pg_rca32_and_3_21_b_21;
  assign f_s_dadda_pg_rca32_and_2_22_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_2_22_y0 = f_s_dadda_pg_rca32_and_2_22_a_2 & f_s_dadda_pg_rca32_and_2_22_b_22;
  assign f_s_dadda_pg_rca32_and_1_23_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_1_23_y0 = f_s_dadda_pg_rca32_and_1_23_a_1 & f_s_dadda_pg_rca32_and_1_23_b_23;
  assign f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_3_21_y0 = f_s_dadda_pg_rca32_and_3_21_y0;
  assign f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_2_22_y0 = f_s_dadda_pg_rca32_and_2_22_y0;
  assign f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_1_23_y0 = f_s_dadda_pg_rca32_and_1_23_y0;
  assign f_s_dadda_pg_rca32_fa182_y0 = f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_3_21_y0 ^ f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_2_22_y0;
  assign f_s_dadda_pg_rca32_fa182_y1 = f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_3_21_y0 & f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_2_22_y0;
  assign f_s_dadda_pg_rca32_fa182_y2 = f_s_dadda_pg_rca32_fa182_y0 ^ f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_1_23_y0;
  assign f_s_dadda_pg_rca32_fa182_y3 = f_s_dadda_pg_rca32_fa182_y0 & f_s_dadda_pg_rca32_fa182_f_s_dadda_pg_rca32_and_1_23_y0;
  assign f_s_dadda_pg_rca32_fa182_y4 = f_s_dadda_pg_rca32_fa182_y1 | f_s_dadda_pg_rca32_fa182_y3;
  assign f_s_dadda_pg_rca32_and_0_24_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_0_24_y0 = f_s_dadda_pg_rca32_and_0_24_a_0 & f_s_dadda_pg_rca32_and_0_24_b_24;
  assign f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_and_0_24_y0 = f_s_dadda_pg_rca32_and_0_24_y0;
  assign f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_fa169_y2 = f_s_dadda_pg_rca32_fa169_y2;
  assign f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_fa170_y2 = f_s_dadda_pg_rca32_fa170_y2;
  assign f_s_dadda_pg_rca32_fa183_y0 = f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_and_0_24_y0 ^ f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_fa169_y2;
  assign f_s_dadda_pg_rca32_fa183_y1 = f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_and_0_24_y0 & f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_fa169_y2;
  assign f_s_dadda_pg_rca32_fa183_y2 = f_s_dadda_pg_rca32_fa183_y0 ^ f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_fa170_y2;
  assign f_s_dadda_pg_rca32_fa183_y3 = f_s_dadda_pg_rca32_fa183_y0 & f_s_dadda_pg_rca32_fa183_f_s_dadda_pg_rca32_fa170_y2;
  assign f_s_dadda_pg_rca32_fa183_y4 = f_s_dadda_pg_rca32_fa183_y1 | f_s_dadda_pg_rca32_fa183_y3;
  assign f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa171_y2 = f_s_dadda_pg_rca32_fa171_y2;
  assign f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa172_y2 = f_s_dadda_pg_rca32_fa172_y2;
  assign f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa173_y2 = f_s_dadda_pg_rca32_fa173_y2;
  assign f_s_dadda_pg_rca32_fa184_y0 = f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa171_y2 ^ f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa172_y2;
  assign f_s_dadda_pg_rca32_fa184_y1 = f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa171_y2 & f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa172_y2;
  assign f_s_dadda_pg_rca32_fa184_y2 = f_s_dadda_pg_rca32_fa184_y0 ^ f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa173_y2;
  assign f_s_dadda_pg_rca32_fa184_y3 = f_s_dadda_pg_rca32_fa184_y0 & f_s_dadda_pg_rca32_fa184_f_s_dadda_pg_rca32_fa173_y2;
  assign f_s_dadda_pg_rca32_fa184_y4 = f_s_dadda_pg_rca32_fa184_y1 | f_s_dadda_pg_rca32_fa184_y3;
  assign f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa174_y2 = f_s_dadda_pg_rca32_fa174_y2;
  assign f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa175_y2 = f_s_dadda_pg_rca32_fa175_y2;
  assign f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa176_y2 = f_s_dadda_pg_rca32_fa176_y2;
  assign f_s_dadda_pg_rca32_fa185_y0 = f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa174_y2 ^ f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa175_y2;
  assign f_s_dadda_pg_rca32_fa185_y1 = f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa174_y2 & f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa175_y2;
  assign f_s_dadda_pg_rca32_fa185_y2 = f_s_dadda_pg_rca32_fa185_y0 ^ f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa176_y2;
  assign f_s_dadda_pg_rca32_fa185_y3 = f_s_dadda_pg_rca32_fa185_y0 & f_s_dadda_pg_rca32_fa185_f_s_dadda_pg_rca32_fa176_y2;
  assign f_s_dadda_pg_rca32_fa185_y4 = f_s_dadda_pg_rca32_fa185_y1 | f_s_dadda_pg_rca32_fa185_y3;
  assign f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa177_y2 = f_s_dadda_pg_rca32_fa177_y2;
  assign f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa178_y2 = f_s_dadda_pg_rca32_fa178_y2;
  assign f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa179_y2 = f_s_dadda_pg_rca32_fa179_y2;
  assign f_s_dadda_pg_rca32_fa186_y0 = f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa177_y2 ^ f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa178_y2;
  assign f_s_dadda_pg_rca32_fa186_y1 = f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa177_y2 & f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa178_y2;
  assign f_s_dadda_pg_rca32_fa186_y2 = f_s_dadda_pg_rca32_fa186_y0 ^ f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa179_y2;
  assign f_s_dadda_pg_rca32_fa186_y3 = f_s_dadda_pg_rca32_fa186_y0 & f_s_dadda_pg_rca32_fa186_f_s_dadda_pg_rca32_fa179_y2;
  assign f_s_dadda_pg_rca32_fa186_y4 = f_s_dadda_pg_rca32_fa186_y1 | f_s_dadda_pg_rca32_fa186_y3;
  assign f_s_dadda_pg_rca32_ha22_f_s_dadda_pg_rca32_fa180_y2 = f_s_dadda_pg_rca32_fa180_y2;
  assign f_s_dadda_pg_rca32_ha22_f_s_dadda_pg_rca32_fa181_y2 = f_s_dadda_pg_rca32_fa181_y2;
  assign f_s_dadda_pg_rca32_ha22_y0 = f_s_dadda_pg_rca32_ha22_f_s_dadda_pg_rca32_fa180_y2 ^ f_s_dadda_pg_rca32_ha22_f_s_dadda_pg_rca32_fa181_y2;
  assign f_s_dadda_pg_rca32_ha22_y1 = f_s_dadda_pg_rca32_ha22_f_s_dadda_pg_rca32_fa180_y2 & f_s_dadda_pg_rca32_ha22_f_s_dadda_pg_rca32_fa181_y2;
  assign f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_ha22_y1 = f_s_dadda_pg_rca32_ha22_y1;
  assign f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_fa186_y4 = f_s_dadda_pg_rca32_fa186_y4;
  assign f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_fa185_y4 = f_s_dadda_pg_rca32_fa185_y4;
  assign f_s_dadda_pg_rca32_fa187_y0 = f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_ha22_y1 ^ f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_fa186_y4;
  assign f_s_dadda_pg_rca32_fa187_y1 = f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_ha22_y1 & f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_fa186_y4;
  assign f_s_dadda_pg_rca32_fa187_y2 = f_s_dadda_pg_rca32_fa187_y0 ^ f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_fa185_y4;
  assign f_s_dadda_pg_rca32_fa187_y3 = f_s_dadda_pg_rca32_fa187_y0 & f_s_dadda_pg_rca32_fa187_f_s_dadda_pg_rca32_fa185_y4;
  assign f_s_dadda_pg_rca32_fa187_y4 = f_s_dadda_pg_rca32_fa187_y1 | f_s_dadda_pg_rca32_fa187_y3;
  assign f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa184_y4 = f_s_dadda_pg_rca32_fa184_y4;
  assign f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa183_y4 = f_s_dadda_pg_rca32_fa183_y4;
  assign f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa182_y4 = f_s_dadda_pg_rca32_fa182_y4;
  assign f_s_dadda_pg_rca32_fa188_y0 = f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa184_y4 ^ f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa183_y4;
  assign f_s_dadda_pg_rca32_fa188_y1 = f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa184_y4 & f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa183_y4;
  assign f_s_dadda_pg_rca32_fa188_y2 = f_s_dadda_pg_rca32_fa188_y0 ^ f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa182_y4;
  assign f_s_dadda_pg_rca32_fa188_y3 = f_s_dadda_pg_rca32_fa188_y0 & f_s_dadda_pg_rca32_fa188_f_s_dadda_pg_rca32_fa182_y4;
  assign f_s_dadda_pg_rca32_fa188_y4 = f_s_dadda_pg_rca32_fa188_y1 | f_s_dadda_pg_rca32_fa188_y3;
  assign f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa181_y4 = f_s_dadda_pg_rca32_fa181_y4;
  assign f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa180_y4 = f_s_dadda_pg_rca32_fa180_y4;
  assign f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa179_y4 = f_s_dadda_pg_rca32_fa179_y4;
  assign f_s_dadda_pg_rca32_fa189_y0 = f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa181_y4 ^ f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa180_y4;
  assign f_s_dadda_pg_rca32_fa189_y1 = f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa181_y4 & f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa180_y4;
  assign f_s_dadda_pg_rca32_fa189_y2 = f_s_dadda_pg_rca32_fa189_y0 ^ f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa179_y4;
  assign f_s_dadda_pg_rca32_fa189_y3 = f_s_dadda_pg_rca32_fa189_y0 & f_s_dadda_pg_rca32_fa189_f_s_dadda_pg_rca32_fa179_y4;
  assign f_s_dadda_pg_rca32_fa189_y4 = f_s_dadda_pg_rca32_fa189_y1 | f_s_dadda_pg_rca32_fa189_y3;
  assign f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa178_y4 = f_s_dadda_pg_rca32_fa178_y4;
  assign f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa177_y4 = f_s_dadda_pg_rca32_fa177_y4;
  assign f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa176_y4 = f_s_dadda_pg_rca32_fa176_y4;
  assign f_s_dadda_pg_rca32_fa190_y0 = f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa178_y4 ^ f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa177_y4;
  assign f_s_dadda_pg_rca32_fa190_y1 = f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa178_y4 & f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa177_y4;
  assign f_s_dadda_pg_rca32_fa190_y2 = f_s_dadda_pg_rca32_fa190_y0 ^ f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa176_y4;
  assign f_s_dadda_pg_rca32_fa190_y3 = f_s_dadda_pg_rca32_fa190_y0 & f_s_dadda_pg_rca32_fa190_f_s_dadda_pg_rca32_fa176_y4;
  assign f_s_dadda_pg_rca32_fa190_y4 = f_s_dadda_pg_rca32_fa190_y1 | f_s_dadda_pg_rca32_fa190_y3;
  assign f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa175_y4 = f_s_dadda_pg_rca32_fa175_y4;
  assign f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa174_y4 = f_s_dadda_pg_rca32_fa174_y4;
  assign f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa173_y4 = f_s_dadda_pg_rca32_fa173_y4;
  assign f_s_dadda_pg_rca32_fa191_y0 = f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa175_y4 ^ f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa174_y4;
  assign f_s_dadda_pg_rca32_fa191_y1 = f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa175_y4 & f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa174_y4;
  assign f_s_dadda_pg_rca32_fa191_y2 = f_s_dadda_pg_rca32_fa191_y0 ^ f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa173_y4;
  assign f_s_dadda_pg_rca32_fa191_y3 = f_s_dadda_pg_rca32_fa191_y0 & f_s_dadda_pg_rca32_fa191_f_s_dadda_pg_rca32_fa173_y4;
  assign f_s_dadda_pg_rca32_fa191_y4 = f_s_dadda_pg_rca32_fa191_y1 | f_s_dadda_pg_rca32_fa191_y3;
  assign f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa172_y4 = f_s_dadda_pg_rca32_fa172_y4;
  assign f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa171_y4 = f_s_dadda_pg_rca32_fa171_y4;
  assign f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa170_y4 = f_s_dadda_pg_rca32_fa170_y4;
  assign f_s_dadda_pg_rca32_fa192_y0 = f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa172_y4 ^ f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa171_y4;
  assign f_s_dadda_pg_rca32_fa192_y1 = f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa172_y4 & f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa171_y4;
  assign f_s_dadda_pg_rca32_fa192_y2 = f_s_dadda_pg_rca32_fa192_y0 ^ f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa170_y4;
  assign f_s_dadda_pg_rca32_fa192_y3 = f_s_dadda_pg_rca32_fa192_y0 & f_s_dadda_pg_rca32_fa192_f_s_dadda_pg_rca32_fa170_y4;
  assign f_s_dadda_pg_rca32_fa192_y4 = f_s_dadda_pg_rca32_fa192_y1 | f_s_dadda_pg_rca32_fa192_y3;
  assign f_s_dadda_pg_rca32_and_25_0_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_25_0_y0 = f_s_dadda_pg_rca32_and_25_0_a_25 & f_s_dadda_pg_rca32_and_25_0_b_0;
  assign f_s_dadda_pg_rca32_and_24_1_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_24_1_y0 = f_s_dadda_pg_rca32_and_24_1_a_24 & f_s_dadda_pg_rca32_and_24_1_b_1;
  assign f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_fa169_y4 = f_s_dadda_pg_rca32_fa169_y4;
  assign f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_and_25_0_y0 = f_s_dadda_pg_rca32_and_25_0_y0;
  assign f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_and_24_1_y0 = f_s_dadda_pg_rca32_and_24_1_y0;
  assign f_s_dadda_pg_rca32_fa193_y0 = f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_fa169_y4 ^ f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_and_25_0_y0;
  assign f_s_dadda_pg_rca32_fa193_y1 = f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_fa169_y4 & f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_and_25_0_y0;
  assign f_s_dadda_pg_rca32_fa193_y2 = f_s_dadda_pg_rca32_fa193_y0 ^ f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_and_24_1_y0;
  assign f_s_dadda_pg_rca32_fa193_y3 = f_s_dadda_pg_rca32_fa193_y0 & f_s_dadda_pg_rca32_fa193_f_s_dadda_pg_rca32_and_24_1_y0;
  assign f_s_dadda_pg_rca32_fa193_y4 = f_s_dadda_pg_rca32_fa193_y1 | f_s_dadda_pg_rca32_fa193_y3;
  assign f_s_dadda_pg_rca32_and_23_2_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_23_2_y0 = f_s_dadda_pg_rca32_and_23_2_a_23 & f_s_dadda_pg_rca32_and_23_2_b_2;
  assign f_s_dadda_pg_rca32_and_22_3_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_22_3_y0 = f_s_dadda_pg_rca32_and_22_3_a_22 & f_s_dadda_pg_rca32_and_22_3_b_3;
  assign f_s_dadda_pg_rca32_and_21_4_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_21_4_y0 = f_s_dadda_pg_rca32_and_21_4_a_21 & f_s_dadda_pg_rca32_and_21_4_b_4;
  assign f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_23_2_y0 = f_s_dadda_pg_rca32_and_23_2_y0;
  assign f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_22_3_y0 = f_s_dadda_pg_rca32_and_22_3_y0;
  assign f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_21_4_y0 = f_s_dadda_pg_rca32_and_21_4_y0;
  assign f_s_dadda_pg_rca32_fa194_y0 = f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_23_2_y0 ^ f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_22_3_y0;
  assign f_s_dadda_pg_rca32_fa194_y1 = f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_23_2_y0 & f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_22_3_y0;
  assign f_s_dadda_pg_rca32_fa194_y2 = f_s_dadda_pg_rca32_fa194_y0 ^ f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_21_4_y0;
  assign f_s_dadda_pg_rca32_fa194_y3 = f_s_dadda_pg_rca32_fa194_y0 & f_s_dadda_pg_rca32_fa194_f_s_dadda_pg_rca32_and_21_4_y0;
  assign f_s_dadda_pg_rca32_fa194_y4 = f_s_dadda_pg_rca32_fa194_y1 | f_s_dadda_pg_rca32_fa194_y3;
  assign f_s_dadda_pg_rca32_and_20_5_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_20_5_y0 = f_s_dadda_pg_rca32_and_20_5_a_20 & f_s_dadda_pg_rca32_and_20_5_b_5;
  assign f_s_dadda_pg_rca32_and_19_6_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_19_6_y0 = f_s_dadda_pg_rca32_and_19_6_a_19 & f_s_dadda_pg_rca32_and_19_6_b_6;
  assign f_s_dadda_pg_rca32_and_18_7_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_18_7_y0 = f_s_dadda_pg_rca32_and_18_7_a_18 & f_s_dadda_pg_rca32_and_18_7_b_7;
  assign f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_20_5_y0 = f_s_dadda_pg_rca32_and_20_5_y0;
  assign f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_19_6_y0 = f_s_dadda_pg_rca32_and_19_6_y0;
  assign f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_18_7_y0 = f_s_dadda_pg_rca32_and_18_7_y0;
  assign f_s_dadda_pg_rca32_fa195_y0 = f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_20_5_y0 ^ f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_19_6_y0;
  assign f_s_dadda_pg_rca32_fa195_y1 = f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_20_5_y0 & f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_19_6_y0;
  assign f_s_dadda_pg_rca32_fa195_y2 = f_s_dadda_pg_rca32_fa195_y0 ^ f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_18_7_y0;
  assign f_s_dadda_pg_rca32_fa195_y3 = f_s_dadda_pg_rca32_fa195_y0 & f_s_dadda_pg_rca32_fa195_f_s_dadda_pg_rca32_and_18_7_y0;
  assign f_s_dadda_pg_rca32_fa195_y4 = f_s_dadda_pg_rca32_fa195_y1 | f_s_dadda_pg_rca32_fa195_y3;
  assign f_s_dadda_pg_rca32_and_17_8_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_17_8_y0 = f_s_dadda_pg_rca32_and_17_8_a_17 & f_s_dadda_pg_rca32_and_17_8_b_8;
  assign f_s_dadda_pg_rca32_and_16_9_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_16_9_y0 = f_s_dadda_pg_rca32_and_16_9_a_16 & f_s_dadda_pg_rca32_and_16_9_b_9;
  assign f_s_dadda_pg_rca32_and_15_10_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_15_10_y0 = f_s_dadda_pg_rca32_and_15_10_a_15 & f_s_dadda_pg_rca32_and_15_10_b_10;
  assign f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_17_8_y0 = f_s_dadda_pg_rca32_and_17_8_y0;
  assign f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_16_9_y0 = f_s_dadda_pg_rca32_and_16_9_y0;
  assign f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_15_10_y0 = f_s_dadda_pg_rca32_and_15_10_y0;
  assign f_s_dadda_pg_rca32_fa196_y0 = f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_17_8_y0 ^ f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_16_9_y0;
  assign f_s_dadda_pg_rca32_fa196_y1 = f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_17_8_y0 & f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_16_9_y0;
  assign f_s_dadda_pg_rca32_fa196_y2 = f_s_dadda_pg_rca32_fa196_y0 ^ f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_15_10_y0;
  assign f_s_dadda_pg_rca32_fa196_y3 = f_s_dadda_pg_rca32_fa196_y0 & f_s_dadda_pg_rca32_fa196_f_s_dadda_pg_rca32_and_15_10_y0;
  assign f_s_dadda_pg_rca32_fa196_y4 = f_s_dadda_pg_rca32_fa196_y1 | f_s_dadda_pg_rca32_fa196_y3;
  assign f_s_dadda_pg_rca32_and_14_11_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_14_11_y0 = f_s_dadda_pg_rca32_and_14_11_a_14 & f_s_dadda_pg_rca32_and_14_11_b_11;
  assign f_s_dadda_pg_rca32_and_13_12_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_13_12_y0 = f_s_dadda_pg_rca32_and_13_12_a_13 & f_s_dadda_pg_rca32_and_13_12_b_12;
  assign f_s_dadda_pg_rca32_and_12_13_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_12_13_y0 = f_s_dadda_pg_rca32_and_12_13_a_12 & f_s_dadda_pg_rca32_and_12_13_b_13;
  assign f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_14_11_y0 = f_s_dadda_pg_rca32_and_14_11_y0;
  assign f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_13_12_y0 = f_s_dadda_pg_rca32_and_13_12_y0;
  assign f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_12_13_y0 = f_s_dadda_pg_rca32_and_12_13_y0;
  assign f_s_dadda_pg_rca32_fa197_y0 = f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_14_11_y0 ^ f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_13_12_y0;
  assign f_s_dadda_pg_rca32_fa197_y1 = f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_14_11_y0 & f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_13_12_y0;
  assign f_s_dadda_pg_rca32_fa197_y2 = f_s_dadda_pg_rca32_fa197_y0 ^ f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_12_13_y0;
  assign f_s_dadda_pg_rca32_fa197_y3 = f_s_dadda_pg_rca32_fa197_y0 & f_s_dadda_pg_rca32_fa197_f_s_dadda_pg_rca32_and_12_13_y0;
  assign f_s_dadda_pg_rca32_fa197_y4 = f_s_dadda_pg_rca32_fa197_y1 | f_s_dadda_pg_rca32_fa197_y3;
  assign f_s_dadda_pg_rca32_and_11_14_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_11_14_y0 = f_s_dadda_pg_rca32_and_11_14_a_11 & f_s_dadda_pg_rca32_and_11_14_b_14;
  assign f_s_dadda_pg_rca32_and_10_15_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_10_15_y0 = f_s_dadda_pg_rca32_and_10_15_a_10 & f_s_dadda_pg_rca32_and_10_15_b_15;
  assign f_s_dadda_pg_rca32_and_9_16_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_9_16_y0 = f_s_dadda_pg_rca32_and_9_16_a_9 & f_s_dadda_pg_rca32_and_9_16_b_16;
  assign f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_11_14_y0 = f_s_dadda_pg_rca32_and_11_14_y0;
  assign f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_10_15_y0 = f_s_dadda_pg_rca32_and_10_15_y0;
  assign f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_9_16_y0 = f_s_dadda_pg_rca32_and_9_16_y0;
  assign f_s_dadda_pg_rca32_fa198_y0 = f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_11_14_y0 ^ f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_10_15_y0;
  assign f_s_dadda_pg_rca32_fa198_y1 = f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_11_14_y0 & f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_10_15_y0;
  assign f_s_dadda_pg_rca32_fa198_y2 = f_s_dadda_pg_rca32_fa198_y0 ^ f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_9_16_y0;
  assign f_s_dadda_pg_rca32_fa198_y3 = f_s_dadda_pg_rca32_fa198_y0 & f_s_dadda_pg_rca32_fa198_f_s_dadda_pg_rca32_and_9_16_y0;
  assign f_s_dadda_pg_rca32_fa198_y4 = f_s_dadda_pg_rca32_fa198_y1 | f_s_dadda_pg_rca32_fa198_y3;
  assign f_s_dadda_pg_rca32_and_8_17_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_8_17_y0 = f_s_dadda_pg_rca32_and_8_17_a_8 & f_s_dadda_pg_rca32_and_8_17_b_17;
  assign f_s_dadda_pg_rca32_and_7_18_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_7_18_y0 = f_s_dadda_pg_rca32_and_7_18_a_7 & f_s_dadda_pg_rca32_and_7_18_b_18;
  assign f_s_dadda_pg_rca32_and_6_19_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_6_19_y0 = f_s_dadda_pg_rca32_and_6_19_a_6 & f_s_dadda_pg_rca32_and_6_19_b_19;
  assign f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_8_17_y0 = f_s_dadda_pg_rca32_and_8_17_y0;
  assign f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_7_18_y0 = f_s_dadda_pg_rca32_and_7_18_y0;
  assign f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_6_19_y0 = f_s_dadda_pg_rca32_and_6_19_y0;
  assign f_s_dadda_pg_rca32_fa199_y0 = f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_8_17_y0 ^ f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_7_18_y0;
  assign f_s_dadda_pg_rca32_fa199_y1 = f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_8_17_y0 & f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_7_18_y0;
  assign f_s_dadda_pg_rca32_fa199_y2 = f_s_dadda_pg_rca32_fa199_y0 ^ f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_6_19_y0;
  assign f_s_dadda_pg_rca32_fa199_y3 = f_s_dadda_pg_rca32_fa199_y0 & f_s_dadda_pg_rca32_fa199_f_s_dadda_pg_rca32_and_6_19_y0;
  assign f_s_dadda_pg_rca32_fa199_y4 = f_s_dadda_pg_rca32_fa199_y1 | f_s_dadda_pg_rca32_fa199_y3;
  assign f_s_dadda_pg_rca32_and_5_20_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_5_20_y0 = f_s_dadda_pg_rca32_and_5_20_a_5 & f_s_dadda_pg_rca32_and_5_20_b_20;
  assign f_s_dadda_pg_rca32_and_4_21_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_4_21_y0 = f_s_dadda_pg_rca32_and_4_21_a_4 & f_s_dadda_pg_rca32_and_4_21_b_21;
  assign f_s_dadda_pg_rca32_and_3_22_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_3_22_y0 = f_s_dadda_pg_rca32_and_3_22_a_3 & f_s_dadda_pg_rca32_and_3_22_b_22;
  assign f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_5_20_y0 = f_s_dadda_pg_rca32_and_5_20_y0;
  assign f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_4_21_y0 = f_s_dadda_pg_rca32_and_4_21_y0;
  assign f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_3_22_y0 = f_s_dadda_pg_rca32_and_3_22_y0;
  assign f_s_dadda_pg_rca32_fa200_y0 = f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_5_20_y0 ^ f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_4_21_y0;
  assign f_s_dadda_pg_rca32_fa200_y1 = f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_5_20_y0 & f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_4_21_y0;
  assign f_s_dadda_pg_rca32_fa200_y2 = f_s_dadda_pg_rca32_fa200_y0 ^ f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_3_22_y0;
  assign f_s_dadda_pg_rca32_fa200_y3 = f_s_dadda_pg_rca32_fa200_y0 & f_s_dadda_pg_rca32_fa200_f_s_dadda_pg_rca32_and_3_22_y0;
  assign f_s_dadda_pg_rca32_fa200_y4 = f_s_dadda_pg_rca32_fa200_y1 | f_s_dadda_pg_rca32_fa200_y3;
  assign f_s_dadda_pg_rca32_and_2_23_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_2_23_y0 = f_s_dadda_pg_rca32_and_2_23_a_2 & f_s_dadda_pg_rca32_and_2_23_b_23;
  assign f_s_dadda_pg_rca32_and_1_24_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_1_24_y0 = f_s_dadda_pg_rca32_and_1_24_a_1 & f_s_dadda_pg_rca32_and_1_24_b_24;
  assign f_s_dadda_pg_rca32_and_0_25_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_0_25_y0 = f_s_dadda_pg_rca32_and_0_25_a_0 & f_s_dadda_pg_rca32_and_0_25_b_25;
  assign f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_2_23_y0 = f_s_dadda_pg_rca32_and_2_23_y0;
  assign f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_1_24_y0 = f_s_dadda_pg_rca32_and_1_24_y0;
  assign f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_0_25_y0 = f_s_dadda_pg_rca32_and_0_25_y0;
  assign f_s_dadda_pg_rca32_fa201_y0 = f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_2_23_y0 ^ f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_1_24_y0;
  assign f_s_dadda_pg_rca32_fa201_y1 = f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_2_23_y0 & f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_1_24_y0;
  assign f_s_dadda_pg_rca32_fa201_y2 = f_s_dadda_pg_rca32_fa201_y0 ^ f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_0_25_y0;
  assign f_s_dadda_pg_rca32_fa201_y3 = f_s_dadda_pg_rca32_fa201_y0 & f_s_dadda_pg_rca32_fa201_f_s_dadda_pg_rca32_and_0_25_y0;
  assign f_s_dadda_pg_rca32_fa201_y4 = f_s_dadda_pg_rca32_fa201_y1 | f_s_dadda_pg_rca32_fa201_y3;
  assign f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa187_y2 = f_s_dadda_pg_rca32_fa187_y2;
  assign f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa188_y2 = f_s_dadda_pg_rca32_fa188_y2;
  assign f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa189_y2 = f_s_dadda_pg_rca32_fa189_y2;
  assign f_s_dadda_pg_rca32_fa202_y0 = f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa187_y2 ^ f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa188_y2;
  assign f_s_dadda_pg_rca32_fa202_y1 = f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa187_y2 & f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa188_y2;
  assign f_s_dadda_pg_rca32_fa202_y2 = f_s_dadda_pg_rca32_fa202_y0 ^ f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa189_y2;
  assign f_s_dadda_pg_rca32_fa202_y3 = f_s_dadda_pg_rca32_fa202_y0 & f_s_dadda_pg_rca32_fa202_f_s_dadda_pg_rca32_fa189_y2;
  assign f_s_dadda_pg_rca32_fa202_y4 = f_s_dadda_pg_rca32_fa202_y1 | f_s_dadda_pg_rca32_fa202_y3;
  assign f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa190_y2 = f_s_dadda_pg_rca32_fa190_y2;
  assign f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa191_y2 = f_s_dadda_pg_rca32_fa191_y2;
  assign f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa192_y2 = f_s_dadda_pg_rca32_fa192_y2;
  assign f_s_dadda_pg_rca32_fa203_y0 = f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa190_y2 ^ f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa191_y2;
  assign f_s_dadda_pg_rca32_fa203_y1 = f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa190_y2 & f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa191_y2;
  assign f_s_dadda_pg_rca32_fa203_y2 = f_s_dadda_pg_rca32_fa203_y0 ^ f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa192_y2;
  assign f_s_dadda_pg_rca32_fa203_y3 = f_s_dadda_pg_rca32_fa203_y0 & f_s_dadda_pg_rca32_fa203_f_s_dadda_pg_rca32_fa192_y2;
  assign f_s_dadda_pg_rca32_fa203_y4 = f_s_dadda_pg_rca32_fa203_y1 | f_s_dadda_pg_rca32_fa203_y3;
  assign f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa193_y2 = f_s_dadda_pg_rca32_fa193_y2;
  assign f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa194_y2 = f_s_dadda_pg_rca32_fa194_y2;
  assign f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa195_y2 = f_s_dadda_pg_rca32_fa195_y2;
  assign f_s_dadda_pg_rca32_fa204_y0 = f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa193_y2 ^ f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa194_y2;
  assign f_s_dadda_pg_rca32_fa204_y1 = f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa193_y2 & f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa194_y2;
  assign f_s_dadda_pg_rca32_fa204_y2 = f_s_dadda_pg_rca32_fa204_y0 ^ f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa195_y2;
  assign f_s_dadda_pg_rca32_fa204_y3 = f_s_dadda_pg_rca32_fa204_y0 & f_s_dadda_pg_rca32_fa204_f_s_dadda_pg_rca32_fa195_y2;
  assign f_s_dadda_pg_rca32_fa204_y4 = f_s_dadda_pg_rca32_fa204_y1 | f_s_dadda_pg_rca32_fa204_y3;
  assign f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa196_y2 = f_s_dadda_pg_rca32_fa196_y2;
  assign f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa197_y2 = f_s_dadda_pg_rca32_fa197_y2;
  assign f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa198_y2 = f_s_dadda_pg_rca32_fa198_y2;
  assign f_s_dadda_pg_rca32_fa205_y0 = f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa196_y2 ^ f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa197_y2;
  assign f_s_dadda_pg_rca32_fa205_y1 = f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa196_y2 & f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa197_y2;
  assign f_s_dadda_pg_rca32_fa205_y2 = f_s_dadda_pg_rca32_fa205_y0 ^ f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa198_y2;
  assign f_s_dadda_pg_rca32_fa205_y3 = f_s_dadda_pg_rca32_fa205_y0 & f_s_dadda_pg_rca32_fa205_f_s_dadda_pg_rca32_fa198_y2;
  assign f_s_dadda_pg_rca32_fa205_y4 = f_s_dadda_pg_rca32_fa205_y1 | f_s_dadda_pg_rca32_fa205_y3;
  assign f_s_dadda_pg_rca32_ha23_f_s_dadda_pg_rca32_fa199_y2 = f_s_dadda_pg_rca32_fa199_y2;
  assign f_s_dadda_pg_rca32_ha23_f_s_dadda_pg_rca32_fa200_y2 = f_s_dadda_pg_rca32_fa200_y2;
  assign f_s_dadda_pg_rca32_ha23_y0 = f_s_dadda_pg_rca32_ha23_f_s_dadda_pg_rca32_fa199_y2 ^ f_s_dadda_pg_rca32_ha23_f_s_dadda_pg_rca32_fa200_y2;
  assign f_s_dadda_pg_rca32_ha23_y1 = f_s_dadda_pg_rca32_ha23_f_s_dadda_pg_rca32_fa199_y2 & f_s_dadda_pg_rca32_ha23_f_s_dadda_pg_rca32_fa200_y2;
  assign f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_ha23_y1 = f_s_dadda_pg_rca32_ha23_y1;
  assign f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_fa205_y4 = f_s_dadda_pg_rca32_fa205_y4;
  assign f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_fa204_y4 = f_s_dadda_pg_rca32_fa204_y4;
  assign f_s_dadda_pg_rca32_fa206_y0 = f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_ha23_y1 ^ f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_fa205_y4;
  assign f_s_dadda_pg_rca32_fa206_y1 = f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_ha23_y1 & f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_fa205_y4;
  assign f_s_dadda_pg_rca32_fa206_y2 = f_s_dadda_pg_rca32_fa206_y0 ^ f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_fa204_y4;
  assign f_s_dadda_pg_rca32_fa206_y3 = f_s_dadda_pg_rca32_fa206_y0 & f_s_dadda_pg_rca32_fa206_f_s_dadda_pg_rca32_fa204_y4;
  assign f_s_dadda_pg_rca32_fa206_y4 = f_s_dadda_pg_rca32_fa206_y1 | f_s_dadda_pg_rca32_fa206_y3;
  assign f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa203_y4 = f_s_dadda_pg_rca32_fa203_y4;
  assign f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa202_y4 = f_s_dadda_pg_rca32_fa202_y4;
  assign f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa201_y4 = f_s_dadda_pg_rca32_fa201_y4;
  assign f_s_dadda_pg_rca32_fa207_y0 = f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa203_y4 ^ f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa202_y4;
  assign f_s_dadda_pg_rca32_fa207_y1 = f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa203_y4 & f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa202_y4;
  assign f_s_dadda_pg_rca32_fa207_y2 = f_s_dadda_pg_rca32_fa207_y0 ^ f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa201_y4;
  assign f_s_dadda_pg_rca32_fa207_y3 = f_s_dadda_pg_rca32_fa207_y0 & f_s_dadda_pg_rca32_fa207_f_s_dadda_pg_rca32_fa201_y4;
  assign f_s_dadda_pg_rca32_fa207_y4 = f_s_dadda_pg_rca32_fa207_y1 | f_s_dadda_pg_rca32_fa207_y3;
  assign f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa200_y4 = f_s_dadda_pg_rca32_fa200_y4;
  assign f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa199_y4 = f_s_dadda_pg_rca32_fa199_y4;
  assign f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa198_y4 = f_s_dadda_pg_rca32_fa198_y4;
  assign f_s_dadda_pg_rca32_fa208_y0 = f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa200_y4 ^ f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa199_y4;
  assign f_s_dadda_pg_rca32_fa208_y1 = f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa200_y4 & f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa199_y4;
  assign f_s_dadda_pg_rca32_fa208_y2 = f_s_dadda_pg_rca32_fa208_y0 ^ f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa198_y4;
  assign f_s_dadda_pg_rca32_fa208_y3 = f_s_dadda_pg_rca32_fa208_y0 & f_s_dadda_pg_rca32_fa208_f_s_dadda_pg_rca32_fa198_y4;
  assign f_s_dadda_pg_rca32_fa208_y4 = f_s_dadda_pg_rca32_fa208_y1 | f_s_dadda_pg_rca32_fa208_y3;
  assign f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa197_y4 = f_s_dadda_pg_rca32_fa197_y4;
  assign f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa196_y4 = f_s_dadda_pg_rca32_fa196_y4;
  assign f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa195_y4 = f_s_dadda_pg_rca32_fa195_y4;
  assign f_s_dadda_pg_rca32_fa209_y0 = f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa197_y4 ^ f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa196_y4;
  assign f_s_dadda_pg_rca32_fa209_y1 = f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa197_y4 & f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa196_y4;
  assign f_s_dadda_pg_rca32_fa209_y2 = f_s_dadda_pg_rca32_fa209_y0 ^ f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa195_y4;
  assign f_s_dadda_pg_rca32_fa209_y3 = f_s_dadda_pg_rca32_fa209_y0 & f_s_dadda_pg_rca32_fa209_f_s_dadda_pg_rca32_fa195_y4;
  assign f_s_dadda_pg_rca32_fa209_y4 = f_s_dadda_pg_rca32_fa209_y1 | f_s_dadda_pg_rca32_fa209_y3;
  assign f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa194_y4 = f_s_dadda_pg_rca32_fa194_y4;
  assign f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa193_y4 = f_s_dadda_pg_rca32_fa193_y4;
  assign f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa192_y4 = f_s_dadda_pg_rca32_fa192_y4;
  assign f_s_dadda_pg_rca32_fa210_y0 = f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa194_y4 ^ f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa193_y4;
  assign f_s_dadda_pg_rca32_fa210_y1 = f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa194_y4 & f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa193_y4;
  assign f_s_dadda_pg_rca32_fa210_y2 = f_s_dadda_pg_rca32_fa210_y0 ^ f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa192_y4;
  assign f_s_dadda_pg_rca32_fa210_y3 = f_s_dadda_pg_rca32_fa210_y0 & f_s_dadda_pg_rca32_fa210_f_s_dadda_pg_rca32_fa192_y4;
  assign f_s_dadda_pg_rca32_fa210_y4 = f_s_dadda_pg_rca32_fa210_y1 | f_s_dadda_pg_rca32_fa210_y3;
  assign f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa191_y4 = f_s_dadda_pg_rca32_fa191_y4;
  assign f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa190_y4 = f_s_dadda_pg_rca32_fa190_y4;
  assign f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa189_y4 = f_s_dadda_pg_rca32_fa189_y4;
  assign f_s_dadda_pg_rca32_fa211_y0 = f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa191_y4 ^ f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa190_y4;
  assign f_s_dadda_pg_rca32_fa211_y1 = f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa191_y4 & f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa190_y4;
  assign f_s_dadda_pg_rca32_fa211_y2 = f_s_dadda_pg_rca32_fa211_y0 ^ f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa189_y4;
  assign f_s_dadda_pg_rca32_fa211_y3 = f_s_dadda_pg_rca32_fa211_y0 & f_s_dadda_pg_rca32_fa211_f_s_dadda_pg_rca32_fa189_y4;
  assign f_s_dadda_pg_rca32_fa211_y4 = f_s_dadda_pg_rca32_fa211_y1 | f_s_dadda_pg_rca32_fa211_y3;
  assign f_s_dadda_pg_rca32_and_26_0_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_26_0_y0 = f_s_dadda_pg_rca32_and_26_0_a_26 & f_s_dadda_pg_rca32_and_26_0_b_0;
  assign f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_fa188_y4 = f_s_dadda_pg_rca32_fa188_y4;
  assign f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_fa187_y4 = f_s_dadda_pg_rca32_fa187_y4;
  assign f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_and_26_0_y0 = f_s_dadda_pg_rca32_and_26_0_y0;
  assign f_s_dadda_pg_rca32_fa212_y0 = f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_fa188_y4 ^ f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_fa187_y4;
  assign f_s_dadda_pg_rca32_fa212_y1 = f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_fa188_y4 & f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_fa187_y4;
  assign f_s_dadda_pg_rca32_fa212_y2 = f_s_dadda_pg_rca32_fa212_y0 ^ f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_and_26_0_y0;
  assign f_s_dadda_pg_rca32_fa212_y3 = f_s_dadda_pg_rca32_fa212_y0 & f_s_dadda_pg_rca32_fa212_f_s_dadda_pg_rca32_and_26_0_y0;
  assign f_s_dadda_pg_rca32_fa212_y4 = f_s_dadda_pg_rca32_fa212_y1 | f_s_dadda_pg_rca32_fa212_y3;
  assign f_s_dadda_pg_rca32_and_25_1_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_25_1_y0 = f_s_dadda_pg_rca32_and_25_1_a_25 & f_s_dadda_pg_rca32_and_25_1_b_1;
  assign f_s_dadda_pg_rca32_and_24_2_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_24_2_y0 = f_s_dadda_pg_rca32_and_24_2_a_24 & f_s_dadda_pg_rca32_and_24_2_b_2;
  assign f_s_dadda_pg_rca32_and_23_3_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_23_3_y0 = f_s_dadda_pg_rca32_and_23_3_a_23 & f_s_dadda_pg_rca32_and_23_3_b_3;
  assign f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_25_1_y0 = f_s_dadda_pg_rca32_and_25_1_y0;
  assign f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_24_2_y0 = f_s_dadda_pg_rca32_and_24_2_y0;
  assign f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_23_3_y0 = f_s_dadda_pg_rca32_and_23_3_y0;
  assign f_s_dadda_pg_rca32_fa213_y0 = f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_25_1_y0 ^ f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_24_2_y0;
  assign f_s_dadda_pg_rca32_fa213_y1 = f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_25_1_y0 & f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_24_2_y0;
  assign f_s_dadda_pg_rca32_fa213_y2 = f_s_dadda_pg_rca32_fa213_y0 ^ f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_23_3_y0;
  assign f_s_dadda_pg_rca32_fa213_y3 = f_s_dadda_pg_rca32_fa213_y0 & f_s_dadda_pg_rca32_fa213_f_s_dadda_pg_rca32_and_23_3_y0;
  assign f_s_dadda_pg_rca32_fa213_y4 = f_s_dadda_pg_rca32_fa213_y1 | f_s_dadda_pg_rca32_fa213_y3;
  assign f_s_dadda_pg_rca32_and_22_4_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_22_4_y0 = f_s_dadda_pg_rca32_and_22_4_a_22 & f_s_dadda_pg_rca32_and_22_4_b_4;
  assign f_s_dadda_pg_rca32_and_21_5_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_21_5_y0 = f_s_dadda_pg_rca32_and_21_5_a_21 & f_s_dadda_pg_rca32_and_21_5_b_5;
  assign f_s_dadda_pg_rca32_and_20_6_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_20_6_y0 = f_s_dadda_pg_rca32_and_20_6_a_20 & f_s_dadda_pg_rca32_and_20_6_b_6;
  assign f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_22_4_y0 = f_s_dadda_pg_rca32_and_22_4_y0;
  assign f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_21_5_y0 = f_s_dadda_pg_rca32_and_21_5_y0;
  assign f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_20_6_y0 = f_s_dadda_pg_rca32_and_20_6_y0;
  assign f_s_dadda_pg_rca32_fa214_y0 = f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_22_4_y0 ^ f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_21_5_y0;
  assign f_s_dadda_pg_rca32_fa214_y1 = f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_22_4_y0 & f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_21_5_y0;
  assign f_s_dadda_pg_rca32_fa214_y2 = f_s_dadda_pg_rca32_fa214_y0 ^ f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_20_6_y0;
  assign f_s_dadda_pg_rca32_fa214_y3 = f_s_dadda_pg_rca32_fa214_y0 & f_s_dadda_pg_rca32_fa214_f_s_dadda_pg_rca32_and_20_6_y0;
  assign f_s_dadda_pg_rca32_fa214_y4 = f_s_dadda_pg_rca32_fa214_y1 | f_s_dadda_pg_rca32_fa214_y3;
  assign f_s_dadda_pg_rca32_and_19_7_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_19_7_y0 = f_s_dadda_pg_rca32_and_19_7_a_19 & f_s_dadda_pg_rca32_and_19_7_b_7;
  assign f_s_dadda_pg_rca32_and_18_8_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_18_8_y0 = f_s_dadda_pg_rca32_and_18_8_a_18 & f_s_dadda_pg_rca32_and_18_8_b_8;
  assign f_s_dadda_pg_rca32_and_17_9_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_17_9_y0 = f_s_dadda_pg_rca32_and_17_9_a_17 & f_s_dadda_pg_rca32_and_17_9_b_9;
  assign f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_19_7_y0 = f_s_dadda_pg_rca32_and_19_7_y0;
  assign f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_18_8_y0 = f_s_dadda_pg_rca32_and_18_8_y0;
  assign f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_17_9_y0 = f_s_dadda_pg_rca32_and_17_9_y0;
  assign f_s_dadda_pg_rca32_fa215_y0 = f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_19_7_y0 ^ f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_18_8_y0;
  assign f_s_dadda_pg_rca32_fa215_y1 = f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_19_7_y0 & f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_18_8_y0;
  assign f_s_dadda_pg_rca32_fa215_y2 = f_s_dadda_pg_rca32_fa215_y0 ^ f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_17_9_y0;
  assign f_s_dadda_pg_rca32_fa215_y3 = f_s_dadda_pg_rca32_fa215_y0 & f_s_dadda_pg_rca32_fa215_f_s_dadda_pg_rca32_and_17_9_y0;
  assign f_s_dadda_pg_rca32_fa215_y4 = f_s_dadda_pg_rca32_fa215_y1 | f_s_dadda_pg_rca32_fa215_y3;
  assign f_s_dadda_pg_rca32_and_16_10_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_16_10_y0 = f_s_dadda_pg_rca32_and_16_10_a_16 & f_s_dadda_pg_rca32_and_16_10_b_10;
  assign f_s_dadda_pg_rca32_and_15_11_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_15_11_y0 = f_s_dadda_pg_rca32_and_15_11_a_15 & f_s_dadda_pg_rca32_and_15_11_b_11;
  assign f_s_dadda_pg_rca32_and_14_12_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_14_12_y0 = f_s_dadda_pg_rca32_and_14_12_a_14 & f_s_dadda_pg_rca32_and_14_12_b_12;
  assign f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_16_10_y0 = f_s_dadda_pg_rca32_and_16_10_y0;
  assign f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_15_11_y0 = f_s_dadda_pg_rca32_and_15_11_y0;
  assign f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_14_12_y0 = f_s_dadda_pg_rca32_and_14_12_y0;
  assign f_s_dadda_pg_rca32_fa216_y0 = f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_16_10_y0 ^ f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_15_11_y0;
  assign f_s_dadda_pg_rca32_fa216_y1 = f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_16_10_y0 & f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_15_11_y0;
  assign f_s_dadda_pg_rca32_fa216_y2 = f_s_dadda_pg_rca32_fa216_y0 ^ f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_14_12_y0;
  assign f_s_dadda_pg_rca32_fa216_y3 = f_s_dadda_pg_rca32_fa216_y0 & f_s_dadda_pg_rca32_fa216_f_s_dadda_pg_rca32_and_14_12_y0;
  assign f_s_dadda_pg_rca32_fa216_y4 = f_s_dadda_pg_rca32_fa216_y1 | f_s_dadda_pg_rca32_fa216_y3;
  assign f_s_dadda_pg_rca32_and_13_13_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_13_13_y0 = f_s_dadda_pg_rca32_and_13_13_a_13 & f_s_dadda_pg_rca32_and_13_13_b_13;
  assign f_s_dadda_pg_rca32_and_12_14_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_12_14_y0 = f_s_dadda_pg_rca32_and_12_14_a_12 & f_s_dadda_pg_rca32_and_12_14_b_14;
  assign f_s_dadda_pg_rca32_and_11_15_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_11_15_y0 = f_s_dadda_pg_rca32_and_11_15_a_11 & f_s_dadda_pg_rca32_and_11_15_b_15;
  assign f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_13_13_y0 = f_s_dadda_pg_rca32_and_13_13_y0;
  assign f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_12_14_y0 = f_s_dadda_pg_rca32_and_12_14_y0;
  assign f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_11_15_y0 = f_s_dadda_pg_rca32_and_11_15_y0;
  assign f_s_dadda_pg_rca32_fa217_y0 = f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_13_13_y0 ^ f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_12_14_y0;
  assign f_s_dadda_pg_rca32_fa217_y1 = f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_13_13_y0 & f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_12_14_y0;
  assign f_s_dadda_pg_rca32_fa217_y2 = f_s_dadda_pg_rca32_fa217_y0 ^ f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_11_15_y0;
  assign f_s_dadda_pg_rca32_fa217_y3 = f_s_dadda_pg_rca32_fa217_y0 & f_s_dadda_pg_rca32_fa217_f_s_dadda_pg_rca32_and_11_15_y0;
  assign f_s_dadda_pg_rca32_fa217_y4 = f_s_dadda_pg_rca32_fa217_y1 | f_s_dadda_pg_rca32_fa217_y3;
  assign f_s_dadda_pg_rca32_and_10_16_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_10_16_y0 = f_s_dadda_pg_rca32_and_10_16_a_10 & f_s_dadda_pg_rca32_and_10_16_b_16;
  assign f_s_dadda_pg_rca32_and_9_17_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_9_17_y0 = f_s_dadda_pg_rca32_and_9_17_a_9 & f_s_dadda_pg_rca32_and_9_17_b_17;
  assign f_s_dadda_pg_rca32_and_8_18_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_8_18_y0 = f_s_dadda_pg_rca32_and_8_18_a_8 & f_s_dadda_pg_rca32_and_8_18_b_18;
  assign f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_10_16_y0 = f_s_dadda_pg_rca32_and_10_16_y0;
  assign f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_9_17_y0 = f_s_dadda_pg_rca32_and_9_17_y0;
  assign f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_8_18_y0 = f_s_dadda_pg_rca32_and_8_18_y0;
  assign f_s_dadda_pg_rca32_fa218_y0 = f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_10_16_y0 ^ f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_9_17_y0;
  assign f_s_dadda_pg_rca32_fa218_y1 = f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_10_16_y0 & f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_9_17_y0;
  assign f_s_dadda_pg_rca32_fa218_y2 = f_s_dadda_pg_rca32_fa218_y0 ^ f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_8_18_y0;
  assign f_s_dadda_pg_rca32_fa218_y3 = f_s_dadda_pg_rca32_fa218_y0 & f_s_dadda_pg_rca32_fa218_f_s_dadda_pg_rca32_and_8_18_y0;
  assign f_s_dadda_pg_rca32_fa218_y4 = f_s_dadda_pg_rca32_fa218_y1 | f_s_dadda_pg_rca32_fa218_y3;
  assign f_s_dadda_pg_rca32_and_7_19_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_7_19_y0 = f_s_dadda_pg_rca32_and_7_19_a_7 & f_s_dadda_pg_rca32_and_7_19_b_19;
  assign f_s_dadda_pg_rca32_and_6_20_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_6_20_y0 = f_s_dadda_pg_rca32_and_6_20_a_6 & f_s_dadda_pg_rca32_and_6_20_b_20;
  assign f_s_dadda_pg_rca32_and_5_21_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_5_21_y0 = f_s_dadda_pg_rca32_and_5_21_a_5 & f_s_dadda_pg_rca32_and_5_21_b_21;
  assign f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_7_19_y0 = f_s_dadda_pg_rca32_and_7_19_y0;
  assign f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_6_20_y0 = f_s_dadda_pg_rca32_and_6_20_y0;
  assign f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_5_21_y0 = f_s_dadda_pg_rca32_and_5_21_y0;
  assign f_s_dadda_pg_rca32_fa219_y0 = f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_7_19_y0 ^ f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_6_20_y0;
  assign f_s_dadda_pg_rca32_fa219_y1 = f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_7_19_y0 & f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_6_20_y0;
  assign f_s_dadda_pg_rca32_fa219_y2 = f_s_dadda_pg_rca32_fa219_y0 ^ f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_5_21_y0;
  assign f_s_dadda_pg_rca32_fa219_y3 = f_s_dadda_pg_rca32_fa219_y0 & f_s_dadda_pg_rca32_fa219_f_s_dadda_pg_rca32_and_5_21_y0;
  assign f_s_dadda_pg_rca32_fa219_y4 = f_s_dadda_pg_rca32_fa219_y1 | f_s_dadda_pg_rca32_fa219_y3;
  assign f_s_dadda_pg_rca32_and_4_22_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_4_22_y0 = f_s_dadda_pg_rca32_and_4_22_a_4 & f_s_dadda_pg_rca32_and_4_22_b_22;
  assign f_s_dadda_pg_rca32_and_3_23_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_3_23_y0 = f_s_dadda_pg_rca32_and_3_23_a_3 & f_s_dadda_pg_rca32_and_3_23_b_23;
  assign f_s_dadda_pg_rca32_and_2_24_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_2_24_y0 = f_s_dadda_pg_rca32_and_2_24_a_2 & f_s_dadda_pg_rca32_and_2_24_b_24;
  assign f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_4_22_y0 = f_s_dadda_pg_rca32_and_4_22_y0;
  assign f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_3_23_y0 = f_s_dadda_pg_rca32_and_3_23_y0;
  assign f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_2_24_y0 = f_s_dadda_pg_rca32_and_2_24_y0;
  assign f_s_dadda_pg_rca32_fa220_y0 = f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_4_22_y0 ^ f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_3_23_y0;
  assign f_s_dadda_pg_rca32_fa220_y1 = f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_4_22_y0 & f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_3_23_y0;
  assign f_s_dadda_pg_rca32_fa220_y2 = f_s_dadda_pg_rca32_fa220_y0 ^ f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_2_24_y0;
  assign f_s_dadda_pg_rca32_fa220_y3 = f_s_dadda_pg_rca32_fa220_y0 & f_s_dadda_pg_rca32_fa220_f_s_dadda_pg_rca32_and_2_24_y0;
  assign f_s_dadda_pg_rca32_fa220_y4 = f_s_dadda_pg_rca32_fa220_y1 | f_s_dadda_pg_rca32_fa220_y3;
  assign f_s_dadda_pg_rca32_and_1_25_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_1_25_y0 = f_s_dadda_pg_rca32_and_1_25_a_1 & f_s_dadda_pg_rca32_and_1_25_b_25;
  assign f_s_dadda_pg_rca32_and_0_26_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_0_26_y0 = f_s_dadda_pg_rca32_and_0_26_a_0 & f_s_dadda_pg_rca32_and_0_26_b_26;
  assign f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_and_1_25_y0 = f_s_dadda_pg_rca32_and_1_25_y0;
  assign f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_and_0_26_y0 = f_s_dadda_pg_rca32_and_0_26_y0;
  assign f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_fa206_y2 = f_s_dadda_pg_rca32_fa206_y2;
  assign f_s_dadda_pg_rca32_fa221_y0 = f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_and_1_25_y0 ^ f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_and_0_26_y0;
  assign f_s_dadda_pg_rca32_fa221_y1 = f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_and_1_25_y0 & f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_and_0_26_y0;
  assign f_s_dadda_pg_rca32_fa221_y2 = f_s_dadda_pg_rca32_fa221_y0 ^ f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_fa206_y2;
  assign f_s_dadda_pg_rca32_fa221_y3 = f_s_dadda_pg_rca32_fa221_y0 & f_s_dadda_pg_rca32_fa221_f_s_dadda_pg_rca32_fa206_y2;
  assign f_s_dadda_pg_rca32_fa221_y4 = f_s_dadda_pg_rca32_fa221_y1 | f_s_dadda_pg_rca32_fa221_y3;
  assign f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa207_y2 = f_s_dadda_pg_rca32_fa207_y2;
  assign f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa208_y2 = f_s_dadda_pg_rca32_fa208_y2;
  assign f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa209_y2 = f_s_dadda_pg_rca32_fa209_y2;
  assign f_s_dadda_pg_rca32_fa222_y0 = f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa207_y2 ^ f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa208_y2;
  assign f_s_dadda_pg_rca32_fa222_y1 = f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa207_y2 & f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa208_y2;
  assign f_s_dadda_pg_rca32_fa222_y2 = f_s_dadda_pg_rca32_fa222_y0 ^ f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa209_y2;
  assign f_s_dadda_pg_rca32_fa222_y3 = f_s_dadda_pg_rca32_fa222_y0 & f_s_dadda_pg_rca32_fa222_f_s_dadda_pg_rca32_fa209_y2;
  assign f_s_dadda_pg_rca32_fa222_y4 = f_s_dadda_pg_rca32_fa222_y1 | f_s_dadda_pg_rca32_fa222_y3;
  assign f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa210_y2 = f_s_dadda_pg_rca32_fa210_y2;
  assign f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa211_y2 = f_s_dadda_pg_rca32_fa211_y2;
  assign f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa212_y2 = f_s_dadda_pg_rca32_fa212_y2;
  assign f_s_dadda_pg_rca32_fa223_y0 = f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa210_y2 ^ f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa211_y2;
  assign f_s_dadda_pg_rca32_fa223_y1 = f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa210_y2 & f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa211_y2;
  assign f_s_dadda_pg_rca32_fa223_y2 = f_s_dadda_pg_rca32_fa223_y0 ^ f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa212_y2;
  assign f_s_dadda_pg_rca32_fa223_y3 = f_s_dadda_pg_rca32_fa223_y0 & f_s_dadda_pg_rca32_fa223_f_s_dadda_pg_rca32_fa212_y2;
  assign f_s_dadda_pg_rca32_fa223_y4 = f_s_dadda_pg_rca32_fa223_y1 | f_s_dadda_pg_rca32_fa223_y3;
  assign f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa213_y2 = f_s_dadda_pg_rca32_fa213_y2;
  assign f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa214_y2 = f_s_dadda_pg_rca32_fa214_y2;
  assign f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa215_y2 = f_s_dadda_pg_rca32_fa215_y2;
  assign f_s_dadda_pg_rca32_fa224_y0 = f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa213_y2 ^ f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa214_y2;
  assign f_s_dadda_pg_rca32_fa224_y1 = f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa213_y2 & f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa214_y2;
  assign f_s_dadda_pg_rca32_fa224_y2 = f_s_dadda_pg_rca32_fa224_y0 ^ f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa215_y2;
  assign f_s_dadda_pg_rca32_fa224_y3 = f_s_dadda_pg_rca32_fa224_y0 & f_s_dadda_pg_rca32_fa224_f_s_dadda_pg_rca32_fa215_y2;
  assign f_s_dadda_pg_rca32_fa224_y4 = f_s_dadda_pg_rca32_fa224_y1 | f_s_dadda_pg_rca32_fa224_y3;
  assign f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa216_y2 = f_s_dadda_pg_rca32_fa216_y2;
  assign f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa217_y2 = f_s_dadda_pg_rca32_fa217_y2;
  assign f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa218_y2 = f_s_dadda_pg_rca32_fa218_y2;
  assign f_s_dadda_pg_rca32_fa225_y0 = f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa216_y2 ^ f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa217_y2;
  assign f_s_dadda_pg_rca32_fa225_y1 = f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa216_y2 & f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa217_y2;
  assign f_s_dadda_pg_rca32_fa225_y2 = f_s_dadda_pg_rca32_fa225_y0 ^ f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa218_y2;
  assign f_s_dadda_pg_rca32_fa225_y3 = f_s_dadda_pg_rca32_fa225_y0 & f_s_dadda_pg_rca32_fa225_f_s_dadda_pg_rca32_fa218_y2;
  assign f_s_dadda_pg_rca32_fa225_y4 = f_s_dadda_pg_rca32_fa225_y1 | f_s_dadda_pg_rca32_fa225_y3;
  assign f_s_dadda_pg_rca32_ha24_f_s_dadda_pg_rca32_fa219_y2 = f_s_dadda_pg_rca32_fa219_y2;
  assign f_s_dadda_pg_rca32_ha24_f_s_dadda_pg_rca32_fa220_y2 = f_s_dadda_pg_rca32_fa220_y2;
  assign f_s_dadda_pg_rca32_ha24_y0 = f_s_dadda_pg_rca32_ha24_f_s_dadda_pg_rca32_fa219_y2 ^ f_s_dadda_pg_rca32_ha24_f_s_dadda_pg_rca32_fa220_y2;
  assign f_s_dadda_pg_rca32_ha24_y1 = f_s_dadda_pg_rca32_ha24_f_s_dadda_pg_rca32_fa219_y2 & f_s_dadda_pg_rca32_ha24_f_s_dadda_pg_rca32_fa220_y2;
  assign f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_ha24_y1 = f_s_dadda_pg_rca32_ha24_y1;
  assign f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_fa225_y4 = f_s_dadda_pg_rca32_fa225_y4;
  assign f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_fa224_y4 = f_s_dadda_pg_rca32_fa224_y4;
  assign f_s_dadda_pg_rca32_fa226_y0 = f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_ha24_y1 ^ f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_fa225_y4;
  assign f_s_dadda_pg_rca32_fa226_y1 = f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_ha24_y1 & f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_fa225_y4;
  assign f_s_dadda_pg_rca32_fa226_y2 = f_s_dadda_pg_rca32_fa226_y0 ^ f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_fa224_y4;
  assign f_s_dadda_pg_rca32_fa226_y3 = f_s_dadda_pg_rca32_fa226_y0 & f_s_dadda_pg_rca32_fa226_f_s_dadda_pg_rca32_fa224_y4;
  assign f_s_dadda_pg_rca32_fa226_y4 = f_s_dadda_pg_rca32_fa226_y1 | f_s_dadda_pg_rca32_fa226_y3;
  assign f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa223_y4 = f_s_dadda_pg_rca32_fa223_y4;
  assign f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa222_y4 = f_s_dadda_pg_rca32_fa222_y4;
  assign f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa221_y4 = f_s_dadda_pg_rca32_fa221_y4;
  assign f_s_dadda_pg_rca32_fa227_y0 = f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa223_y4 ^ f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa222_y4;
  assign f_s_dadda_pg_rca32_fa227_y1 = f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa223_y4 & f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa222_y4;
  assign f_s_dadda_pg_rca32_fa227_y2 = f_s_dadda_pg_rca32_fa227_y0 ^ f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa221_y4;
  assign f_s_dadda_pg_rca32_fa227_y3 = f_s_dadda_pg_rca32_fa227_y0 & f_s_dadda_pg_rca32_fa227_f_s_dadda_pg_rca32_fa221_y4;
  assign f_s_dadda_pg_rca32_fa227_y4 = f_s_dadda_pg_rca32_fa227_y1 | f_s_dadda_pg_rca32_fa227_y3;
  assign f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa220_y4 = f_s_dadda_pg_rca32_fa220_y4;
  assign f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa219_y4 = f_s_dadda_pg_rca32_fa219_y4;
  assign f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa218_y4 = f_s_dadda_pg_rca32_fa218_y4;
  assign f_s_dadda_pg_rca32_fa228_y0 = f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa220_y4 ^ f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa219_y4;
  assign f_s_dadda_pg_rca32_fa228_y1 = f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa220_y4 & f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa219_y4;
  assign f_s_dadda_pg_rca32_fa228_y2 = f_s_dadda_pg_rca32_fa228_y0 ^ f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa218_y4;
  assign f_s_dadda_pg_rca32_fa228_y3 = f_s_dadda_pg_rca32_fa228_y0 & f_s_dadda_pg_rca32_fa228_f_s_dadda_pg_rca32_fa218_y4;
  assign f_s_dadda_pg_rca32_fa228_y4 = f_s_dadda_pg_rca32_fa228_y1 | f_s_dadda_pg_rca32_fa228_y3;
  assign f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa217_y4 = f_s_dadda_pg_rca32_fa217_y4;
  assign f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa216_y4 = f_s_dadda_pg_rca32_fa216_y4;
  assign f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa215_y4 = f_s_dadda_pg_rca32_fa215_y4;
  assign f_s_dadda_pg_rca32_fa229_y0 = f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa217_y4 ^ f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa216_y4;
  assign f_s_dadda_pg_rca32_fa229_y1 = f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa217_y4 & f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa216_y4;
  assign f_s_dadda_pg_rca32_fa229_y2 = f_s_dadda_pg_rca32_fa229_y0 ^ f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa215_y4;
  assign f_s_dadda_pg_rca32_fa229_y3 = f_s_dadda_pg_rca32_fa229_y0 & f_s_dadda_pg_rca32_fa229_f_s_dadda_pg_rca32_fa215_y4;
  assign f_s_dadda_pg_rca32_fa229_y4 = f_s_dadda_pg_rca32_fa229_y1 | f_s_dadda_pg_rca32_fa229_y3;
  assign f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa214_y4 = f_s_dadda_pg_rca32_fa214_y4;
  assign f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa213_y4 = f_s_dadda_pg_rca32_fa213_y4;
  assign f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa212_y4 = f_s_dadda_pg_rca32_fa212_y4;
  assign f_s_dadda_pg_rca32_fa230_y0 = f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa214_y4 ^ f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa213_y4;
  assign f_s_dadda_pg_rca32_fa230_y1 = f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa214_y4 & f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa213_y4;
  assign f_s_dadda_pg_rca32_fa230_y2 = f_s_dadda_pg_rca32_fa230_y0 ^ f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa212_y4;
  assign f_s_dadda_pg_rca32_fa230_y3 = f_s_dadda_pg_rca32_fa230_y0 & f_s_dadda_pg_rca32_fa230_f_s_dadda_pg_rca32_fa212_y4;
  assign f_s_dadda_pg_rca32_fa230_y4 = f_s_dadda_pg_rca32_fa230_y1 | f_s_dadda_pg_rca32_fa230_y3;
  assign f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa211_y4 = f_s_dadda_pg_rca32_fa211_y4;
  assign f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa210_y4 = f_s_dadda_pg_rca32_fa210_y4;
  assign f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa209_y4 = f_s_dadda_pg_rca32_fa209_y4;
  assign f_s_dadda_pg_rca32_fa231_y0 = f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa211_y4 ^ f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa210_y4;
  assign f_s_dadda_pg_rca32_fa231_y1 = f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa211_y4 & f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa210_y4;
  assign f_s_dadda_pg_rca32_fa231_y2 = f_s_dadda_pg_rca32_fa231_y0 ^ f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa209_y4;
  assign f_s_dadda_pg_rca32_fa231_y3 = f_s_dadda_pg_rca32_fa231_y0 & f_s_dadda_pg_rca32_fa231_f_s_dadda_pg_rca32_fa209_y4;
  assign f_s_dadda_pg_rca32_fa231_y4 = f_s_dadda_pg_rca32_fa231_y1 | f_s_dadda_pg_rca32_fa231_y3;
  assign f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa208_y4 = f_s_dadda_pg_rca32_fa208_y4;
  assign f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa207_y4 = f_s_dadda_pg_rca32_fa207_y4;
  assign f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa206_y4 = f_s_dadda_pg_rca32_fa206_y4;
  assign f_s_dadda_pg_rca32_fa232_y0 = f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa208_y4 ^ f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa207_y4;
  assign f_s_dadda_pg_rca32_fa232_y1 = f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa208_y4 & f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa207_y4;
  assign f_s_dadda_pg_rca32_fa232_y2 = f_s_dadda_pg_rca32_fa232_y0 ^ f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa206_y4;
  assign f_s_dadda_pg_rca32_fa232_y3 = f_s_dadda_pg_rca32_fa232_y0 & f_s_dadda_pg_rca32_fa232_f_s_dadda_pg_rca32_fa206_y4;
  assign f_s_dadda_pg_rca32_fa232_y4 = f_s_dadda_pg_rca32_fa232_y1 | f_s_dadda_pg_rca32_fa232_y3;
  assign f_s_dadda_pg_rca32_and_27_0_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_27_0_y0 = f_s_dadda_pg_rca32_and_27_0_a_27 & f_s_dadda_pg_rca32_and_27_0_b_0;
  assign f_s_dadda_pg_rca32_and_26_1_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_26_1_y0 = f_s_dadda_pg_rca32_and_26_1_a_26 & f_s_dadda_pg_rca32_and_26_1_b_1;
  assign f_s_dadda_pg_rca32_and_25_2_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_25_2_y0 = f_s_dadda_pg_rca32_and_25_2_a_25 & f_s_dadda_pg_rca32_and_25_2_b_2;
  assign f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_27_0_y0 = f_s_dadda_pg_rca32_and_27_0_y0;
  assign f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_26_1_y0 = f_s_dadda_pg_rca32_and_26_1_y0;
  assign f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_25_2_y0 = f_s_dadda_pg_rca32_and_25_2_y0;
  assign f_s_dadda_pg_rca32_fa233_y0 = f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_27_0_y0 ^ f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_26_1_y0;
  assign f_s_dadda_pg_rca32_fa233_y1 = f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_27_0_y0 & f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_26_1_y0;
  assign f_s_dadda_pg_rca32_fa233_y2 = f_s_dadda_pg_rca32_fa233_y0 ^ f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_25_2_y0;
  assign f_s_dadda_pg_rca32_fa233_y3 = f_s_dadda_pg_rca32_fa233_y0 & f_s_dadda_pg_rca32_fa233_f_s_dadda_pg_rca32_and_25_2_y0;
  assign f_s_dadda_pg_rca32_fa233_y4 = f_s_dadda_pg_rca32_fa233_y1 | f_s_dadda_pg_rca32_fa233_y3;
  assign f_s_dadda_pg_rca32_and_24_3_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_24_3_y0 = f_s_dadda_pg_rca32_and_24_3_a_24 & f_s_dadda_pg_rca32_and_24_3_b_3;
  assign f_s_dadda_pg_rca32_and_23_4_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_23_4_y0 = f_s_dadda_pg_rca32_and_23_4_a_23 & f_s_dadda_pg_rca32_and_23_4_b_4;
  assign f_s_dadda_pg_rca32_and_22_5_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_22_5_y0 = f_s_dadda_pg_rca32_and_22_5_a_22 & f_s_dadda_pg_rca32_and_22_5_b_5;
  assign f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_24_3_y0 = f_s_dadda_pg_rca32_and_24_3_y0;
  assign f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_23_4_y0 = f_s_dadda_pg_rca32_and_23_4_y0;
  assign f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_22_5_y0 = f_s_dadda_pg_rca32_and_22_5_y0;
  assign f_s_dadda_pg_rca32_fa234_y0 = f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_24_3_y0 ^ f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_23_4_y0;
  assign f_s_dadda_pg_rca32_fa234_y1 = f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_24_3_y0 & f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_23_4_y0;
  assign f_s_dadda_pg_rca32_fa234_y2 = f_s_dadda_pg_rca32_fa234_y0 ^ f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_22_5_y0;
  assign f_s_dadda_pg_rca32_fa234_y3 = f_s_dadda_pg_rca32_fa234_y0 & f_s_dadda_pg_rca32_fa234_f_s_dadda_pg_rca32_and_22_5_y0;
  assign f_s_dadda_pg_rca32_fa234_y4 = f_s_dadda_pg_rca32_fa234_y1 | f_s_dadda_pg_rca32_fa234_y3;
  assign f_s_dadda_pg_rca32_and_21_6_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_21_6_y0 = f_s_dadda_pg_rca32_and_21_6_a_21 & f_s_dadda_pg_rca32_and_21_6_b_6;
  assign f_s_dadda_pg_rca32_and_20_7_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_20_7_y0 = f_s_dadda_pg_rca32_and_20_7_a_20 & f_s_dadda_pg_rca32_and_20_7_b_7;
  assign f_s_dadda_pg_rca32_and_19_8_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_19_8_y0 = f_s_dadda_pg_rca32_and_19_8_a_19 & f_s_dadda_pg_rca32_and_19_8_b_8;
  assign f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_21_6_y0 = f_s_dadda_pg_rca32_and_21_6_y0;
  assign f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_20_7_y0 = f_s_dadda_pg_rca32_and_20_7_y0;
  assign f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_19_8_y0 = f_s_dadda_pg_rca32_and_19_8_y0;
  assign f_s_dadda_pg_rca32_fa235_y0 = f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_21_6_y0 ^ f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_20_7_y0;
  assign f_s_dadda_pg_rca32_fa235_y1 = f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_21_6_y0 & f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_20_7_y0;
  assign f_s_dadda_pg_rca32_fa235_y2 = f_s_dadda_pg_rca32_fa235_y0 ^ f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_19_8_y0;
  assign f_s_dadda_pg_rca32_fa235_y3 = f_s_dadda_pg_rca32_fa235_y0 & f_s_dadda_pg_rca32_fa235_f_s_dadda_pg_rca32_and_19_8_y0;
  assign f_s_dadda_pg_rca32_fa235_y4 = f_s_dadda_pg_rca32_fa235_y1 | f_s_dadda_pg_rca32_fa235_y3;
  assign f_s_dadda_pg_rca32_and_18_9_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_18_9_y0 = f_s_dadda_pg_rca32_and_18_9_a_18 & f_s_dadda_pg_rca32_and_18_9_b_9;
  assign f_s_dadda_pg_rca32_and_17_10_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_17_10_y0 = f_s_dadda_pg_rca32_and_17_10_a_17 & f_s_dadda_pg_rca32_and_17_10_b_10;
  assign f_s_dadda_pg_rca32_and_16_11_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_16_11_y0 = f_s_dadda_pg_rca32_and_16_11_a_16 & f_s_dadda_pg_rca32_and_16_11_b_11;
  assign f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_18_9_y0 = f_s_dadda_pg_rca32_and_18_9_y0;
  assign f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_17_10_y0 = f_s_dadda_pg_rca32_and_17_10_y0;
  assign f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_16_11_y0 = f_s_dadda_pg_rca32_and_16_11_y0;
  assign f_s_dadda_pg_rca32_fa236_y0 = f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_18_9_y0 ^ f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_17_10_y0;
  assign f_s_dadda_pg_rca32_fa236_y1 = f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_18_9_y0 & f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_17_10_y0;
  assign f_s_dadda_pg_rca32_fa236_y2 = f_s_dadda_pg_rca32_fa236_y0 ^ f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_16_11_y0;
  assign f_s_dadda_pg_rca32_fa236_y3 = f_s_dadda_pg_rca32_fa236_y0 & f_s_dadda_pg_rca32_fa236_f_s_dadda_pg_rca32_and_16_11_y0;
  assign f_s_dadda_pg_rca32_fa236_y4 = f_s_dadda_pg_rca32_fa236_y1 | f_s_dadda_pg_rca32_fa236_y3;
  assign f_s_dadda_pg_rca32_and_15_12_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_15_12_y0 = f_s_dadda_pg_rca32_and_15_12_a_15 & f_s_dadda_pg_rca32_and_15_12_b_12;
  assign f_s_dadda_pg_rca32_and_14_13_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_14_13_y0 = f_s_dadda_pg_rca32_and_14_13_a_14 & f_s_dadda_pg_rca32_and_14_13_b_13;
  assign f_s_dadda_pg_rca32_and_13_14_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_13_14_y0 = f_s_dadda_pg_rca32_and_13_14_a_13 & f_s_dadda_pg_rca32_and_13_14_b_14;
  assign f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_15_12_y0 = f_s_dadda_pg_rca32_and_15_12_y0;
  assign f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_14_13_y0 = f_s_dadda_pg_rca32_and_14_13_y0;
  assign f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_13_14_y0 = f_s_dadda_pg_rca32_and_13_14_y0;
  assign f_s_dadda_pg_rca32_fa237_y0 = f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_15_12_y0 ^ f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_14_13_y0;
  assign f_s_dadda_pg_rca32_fa237_y1 = f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_15_12_y0 & f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_14_13_y0;
  assign f_s_dadda_pg_rca32_fa237_y2 = f_s_dadda_pg_rca32_fa237_y0 ^ f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_13_14_y0;
  assign f_s_dadda_pg_rca32_fa237_y3 = f_s_dadda_pg_rca32_fa237_y0 & f_s_dadda_pg_rca32_fa237_f_s_dadda_pg_rca32_and_13_14_y0;
  assign f_s_dadda_pg_rca32_fa237_y4 = f_s_dadda_pg_rca32_fa237_y1 | f_s_dadda_pg_rca32_fa237_y3;
  assign f_s_dadda_pg_rca32_and_12_15_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_12_15_y0 = f_s_dadda_pg_rca32_and_12_15_a_12 & f_s_dadda_pg_rca32_and_12_15_b_15;
  assign f_s_dadda_pg_rca32_and_11_16_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_11_16_y0 = f_s_dadda_pg_rca32_and_11_16_a_11 & f_s_dadda_pg_rca32_and_11_16_b_16;
  assign f_s_dadda_pg_rca32_and_10_17_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_10_17_y0 = f_s_dadda_pg_rca32_and_10_17_a_10 & f_s_dadda_pg_rca32_and_10_17_b_17;
  assign f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_12_15_y0 = f_s_dadda_pg_rca32_and_12_15_y0;
  assign f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_11_16_y0 = f_s_dadda_pg_rca32_and_11_16_y0;
  assign f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_10_17_y0 = f_s_dadda_pg_rca32_and_10_17_y0;
  assign f_s_dadda_pg_rca32_fa238_y0 = f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_12_15_y0 ^ f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_11_16_y0;
  assign f_s_dadda_pg_rca32_fa238_y1 = f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_12_15_y0 & f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_11_16_y0;
  assign f_s_dadda_pg_rca32_fa238_y2 = f_s_dadda_pg_rca32_fa238_y0 ^ f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_10_17_y0;
  assign f_s_dadda_pg_rca32_fa238_y3 = f_s_dadda_pg_rca32_fa238_y0 & f_s_dadda_pg_rca32_fa238_f_s_dadda_pg_rca32_and_10_17_y0;
  assign f_s_dadda_pg_rca32_fa238_y4 = f_s_dadda_pg_rca32_fa238_y1 | f_s_dadda_pg_rca32_fa238_y3;
  assign f_s_dadda_pg_rca32_and_9_18_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_9_18_y0 = f_s_dadda_pg_rca32_and_9_18_a_9 & f_s_dadda_pg_rca32_and_9_18_b_18;
  assign f_s_dadda_pg_rca32_and_8_19_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_8_19_y0 = f_s_dadda_pg_rca32_and_8_19_a_8 & f_s_dadda_pg_rca32_and_8_19_b_19;
  assign f_s_dadda_pg_rca32_and_7_20_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_7_20_y0 = f_s_dadda_pg_rca32_and_7_20_a_7 & f_s_dadda_pg_rca32_and_7_20_b_20;
  assign f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_9_18_y0 = f_s_dadda_pg_rca32_and_9_18_y0;
  assign f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_8_19_y0 = f_s_dadda_pg_rca32_and_8_19_y0;
  assign f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_7_20_y0 = f_s_dadda_pg_rca32_and_7_20_y0;
  assign f_s_dadda_pg_rca32_fa239_y0 = f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_9_18_y0 ^ f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_8_19_y0;
  assign f_s_dadda_pg_rca32_fa239_y1 = f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_9_18_y0 & f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_8_19_y0;
  assign f_s_dadda_pg_rca32_fa239_y2 = f_s_dadda_pg_rca32_fa239_y0 ^ f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_7_20_y0;
  assign f_s_dadda_pg_rca32_fa239_y3 = f_s_dadda_pg_rca32_fa239_y0 & f_s_dadda_pg_rca32_fa239_f_s_dadda_pg_rca32_and_7_20_y0;
  assign f_s_dadda_pg_rca32_fa239_y4 = f_s_dadda_pg_rca32_fa239_y1 | f_s_dadda_pg_rca32_fa239_y3;
  assign f_s_dadda_pg_rca32_and_6_21_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_6_21_y0 = f_s_dadda_pg_rca32_and_6_21_a_6 & f_s_dadda_pg_rca32_and_6_21_b_21;
  assign f_s_dadda_pg_rca32_and_5_22_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_5_22_y0 = f_s_dadda_pg_rca32_and_5_22_a_5 & f_s_dadda_pg_rca32_and_5_22_b_22;
  assign f_s_dadda_pg_rca32_and_4_23_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_4_23_y0 = f_s_dadda_pg_rca32_and_4_23_a_4 & f_s_dadda_pg_rca32_and_4_23_b_23;
  assign f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_6_21_y0 = f_s_dadda_pg_rca32_and_6_21_y0;
  assign f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_5_22_y0 = f_s_dadda_pg_rca32_and_5_22_y0;
  assign f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_4_23_y0 = f_s_dadda_pg_rca32_and_4_23_y0;
  assign f_s_dadda_pg_rca32_fa240_y0 = f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_6_21_y0 ^ f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_5_22_y0;
  assign f_s_dadda_pg_rca32_fa240_y1 = f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_6_21_y0 & f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_5_22_y0;
  assign f_s_dadda_pg_rca32_fa240_y2 = f_s_dadda_pg_rca32_fa240_y0 ^ f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_4_23_y0;
  assign f_s_dadda_pg_rca32_fa240_y3 = f_s_dadda_pg_rca32_fa240_y0 & f_s_dadda_pg_rca32_fa240_f_s_dadda_pg_rca32_and_4_23_y0;
  assign f_s_dadda_pg_rca32_fa240_y4 = f_s_dadda_pg_rca32_fa240_y1 | f_s_dadda_pg_rca32_fa240_y3;
  assign f_s_dadda_pg_rca32_and_3_24_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_3_24_y0 = f_s_dadda_pg_rca32_and_3_24_a_3 & f_s_dadda_pg_rca32_and_3_24_b_24;
  assign f_s_dadda_pg_rca32_and_2_25_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_2_25_y0 = f_s_dadda_pg_rca32_and_2_25_a_2 & f_s_dadda_pg_rca32_and_2_25_b_25;
  assign f_s_dadda_pg_rca32_and_1_26_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_1_26_y0 = f_s_dadda_pg_rca32_and_1_26_a_1 & f_s_dadda_pg_rca32_and_1_26_b_26;
  assign f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_3_24_y0 = f_s_dadda_pg_rca32_and_3_24_y0;
  assign f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_2_25_y0 = f_s_dadda_pg_rca32_and_2_25_y0;
  assign f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_1_26_y0 = f_s_dadda_pg_rca32_and_1_26_y0;
  assign f_s_dadda_pg_rca32_fa241_y0 = f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_3_24_y0 ^ f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_2_25_y0;
  assign f_s_dadda_pg_rca32_fa241_y1 = f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_3_24_y0 & f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_2_25_y0;
  assign f_s_dadda_pg_rca32_fa241_y2 = f_s_dadda_pg_rca32_fa241_y0 ^ f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_1_26_y0;
  assign f_s_dadda_pg_rca32_fa241_y3 = f_s_dadda_pg_rca32_fa241_y0 & f_s_dadda_pg_rca32_fa241_f_s_dadda_pg_rca32_and_1_26_y0;
  assign f_s_dadda_pg_rca32_fa241_y4 = f_s_dadda_pg_rca32_fa241_y1 | f_s_dadda_pg_rca32_fa241_y3;
  assign f_s_dadda_pg_rca32_and_0_27_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_0_27_y0 = f_s_dadda_pg_rca32_and_0_27_a_0 & f_s_dadda_pg_rca32_and_0_27_b_27;
  assign f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_and_0_27_y0 = f_s_dadda_pg_rca32_and_0_27_y0;
  assign f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_fa226_y2 = f_s_dadda_pg_rca32_fa226_y2;
  assign f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_fa227_y2 = f_s_dadda_pg_rca32_fa227_y2;
  assign f_s_dadda_pg_rca32_fa242_y0 = f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_and_0_27_y0 ^ f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_fa226_y2;
  assign f_s_dadda_pg_rca32_fa242_y1 = f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_and_0_27_y0 & f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_fa226_y2;
  assign f_s_dadda_pg_rca32_fa242_y2 = f_s_dadda_pg_rca32_fa242_y0 ^ f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_fa227_y2;
  assign f_s_dadda_pg_rca32_fa242_y3 = f_s_dadda_pg_rca32_fa242_y0 & f_s_dadda_pg_rca32_fa242_f_s_dadda_pg_rca32_fa227_y2;
  assign f_s_dadda_pg_rca32_fa242_y4 = f_s_dadda_pg_rca32_fa242_y1 | f_s_dadda_pg_rca32_fa242_y3;
  assign f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa228_y2 = f_s_dadda_pg_rca32_fa228_y2;
  assign f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa229_y2 = f_s_dadda_pg_rca32_fa229_y2;
  assign f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa230_y2 = f_s_dadda_pg_rca32_fa230_y2;
  assign f_s_dadda_pg_rca32_fa243_y0 = f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa228_y2 ^ f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa229_y2;
  assign f_s_dadda_pg_rca32_fa243_y1 = f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa228_y2 & f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa229_y2;
  assign f_s_dadda_pg_rca32_fa243_y2 = f_s_dadda_pg_rca32_fa243_y0 ^ f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa230_y2;
  assign f_s_dadda_pg_rca32_fa243_y3 = f_s_dadda_pg_rca32_fa243_y0 & f_s_dadda_pg_rca32_fa243_f_s_dadda_pg_rca32_fa230_y2;
  assign f_s_dadda_pg_rca32_fa243_y4 = f_s_dadda_pg_rca32_fa243_y1 | f_s_dadda_pg_rca32_fa243_y3;
  assign f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa231_y2 = f_s_dadda_pg_rca32_fa231_y2;
  assign f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa232_y2 = f_s_dadda_pg_rca32_fa232_y2;
  assign f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa233_y2 = f_s_dadda_pg_rca32_fa233_y2;
  assign f_s_dadda_pg_rca32_fa244_y0 = f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa231_y2 ^ f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa232_y2;
  assign f_s_dadda_pg_rca32_fa244_y1 = f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa231_y2 & f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa232_y2;
  assign f_s_dadda_pg_rca32_fa244_y2 = f_s_dadda_pg_rca32_fa244_y0 ^ f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa233_y2;
  assign f_s_dadda_pg_rca32_fa244_y3 = f_s_dadda_pg_rca32_fa244_y0 & f_s_dadda_pg_rca32_fa244_f_s_dadda_pg_rca32_fa233_y2;
  assign f_s_dadda_pg_rca32_fa244_y4 = f_s_dadda_pg_rca32_fa244_y1 | f_s_dadda_pg_rca32_fa244_y3;
  assign f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa234_y2 = f_s_dadda_pg_rca32_fa234_y2;
  assign f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa235_y2 = f_s_dadda_pg_rca32_fa235_y2;
  assign f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa236_y2 = f_s_dadda_pg_rca32_fa236_y2;
  assign f_s_dadda_pg_rca32_fa245_y0 = f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa234_y2 ^ f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa235_y2;
  assign f_s_dadda_pg_rca32_fa245_y1 = f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa234_y2 & f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa235_y2;
  assign f_s_dadda_pg_rca32_fa245_y2 = f_s_dadda_pg_rca32_fa245_y0 ^ f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa236_y2;
  assign f_s_dadda_pg_rca32_fa245_y3 = f_s_dadda_pg_rca32_fa245_y0 & f_s_dadda_pg_rca32_fa245_f_s_dadda_pg_rca32_fa236_y2;
  assign f_s_dadda_pg_rca32_fa245_y4 = f_s_dadda_pg_rca32_fa245_y1 | f_s_dadda_pg_rca32_fa245_y3;
  assign f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa237_y2 = f_s_dadda_pg_rca32_fa237_y2;
  assign f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa238_y2 = f_s_dadda_pg_rca32_fa238_y2;
  assign f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa239_y2 = f_s_dadda_pg_rca32_fa239_y2;
  assign f_s_dadda_pg_rca32_fa246_y0 = f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa237_y2 ^ f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa238_y2;
  assign f_s_dadda_pg_rca32_fa246_y1 = f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa237_y2 & f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa238_y2;
  assign f_s_dadda_pg_rca32_fa246_y2 = f_s_dadda_pg_rca32_fa246_y0 ^ f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa239_y2;
  assign f_s_dadda_pg_rca32_fa246_y3 = f_s_dadda_pg_rca32_fa246_y0 & f_s_dadda_pg_rca32_fa246_f_s_dadda_pg_rca32_fa239_y2;
  assign f_s_dadda_pg_rca32_fa246_y4 = f_s_dadda_pg_rca32_fa246_y1 | f_s_dadda_pg_rca32_fa246_y3;
  assign f_s_dadda_pg_rca32_ha25_f_s_dadda_pg_rca32_fa240_y2 = f_s_dadda_pg_rca32_fa240_y2;
  assign f_s_dadda_pg_rca32_ha25_f_s_dadda_pg_rca32_fa241_y2 = f_s_dadda_pg_rca32_fa241_y2;
  assign f_s_dadda_pg_rca32_ha25_y0 = f_s_dadda_pg_rca32_ha25_f_s_dadda_pg_rca32_fa240_y2 ^ f_s_dadda_pg_rca32_ha25_f_s_dadda_pg_rca32_fa241_y2;
  assign f_s_dadda_pg_rca32_ha25_y1 = f_s_dadda_pg_rca32_ha25_f_s_dadda_pg_rca32_fa240_y2 & f_s_dadda_pg_rca32_ha25_f_s_dadda_pg_rca32_fa241_y2;
  assign f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_ha25_y1 = f_s_dadda_pg_rca32_ha25_y1;
  assign f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_fa246_y4 = f_s_dadda_pg_rca32_fa246_y4;
  assign f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_fa245_y4 = f_s_dadda_pg_rca32_fa245_y4;
  assign f_s_dadda_pg_rca32_fa247_y0 = f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_ha25_y1 ^ f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_fa246_y4;
  assign f_s_dadda_pg_rca32_fa247_y1 = f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_ha25_y1 & f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_fa246_y4;
  assign f_s_dadda_pg_rca32_fa247_y2 = f_s_dadda_pg_rca32_fa247_y0 ^ f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_fa245_y4;
  assign f_s_dadda_pg_rca32_fa247_y3 = f_s_dadda_pg_rca32_fa247_y0 & f_s_dadda_pg_rca32_fa247_f_s_dadda_pg_rca32_fa245_y4;
  assign f_s_dadda_pg_rca32_fa247_y4 = f_s_dadda_pg_rca32_fa247_y1 | f_s_dadda_pg_rca32_fa247_y3;
  assign f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa244_y4 = f_s_dadda_pg_rca32_fa244_y4;
  assign f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa243_y4 = f_s_dadda_pg_rca32_fa243_y4;
  assign f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa242_y4 = f_s_dadda_pg_rca32_fa242_y4;
  assign f_s_dadda_pg_rca32_fa248_y0 = f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa244_y4 ^ f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa243_y4;
  assign f_s_dadda_pg_rca32_fa248_y1 = f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa244_y4 & f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa243_y4;
  assign f_s_dadda_pg_rca32_fa248_y2 = f_s_dadda_pg_rca32_fa248_y0 ^ f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa242_y4;
  assign f_s_dadda_pg_rca32_fa248_y3 = f_s_dadda_pg_rca32_fa248_y0 & f_s_dadda_pg_rca32_fa248_f_s_dadda_pg_rca32_fa242_y4;
  assign f_s_dadda_pg_rca32_fa248_y4 = f_s_dadda_pg_rca32_fa248_y1 | f_s_dadda_pg_rca32_fa248_y3;
  assign f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa241_y4 = f_s_dadda_pg_rca32_fa241_y4;
  assign f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa240_y4 = f_s_dadda_pg_rca32_fa240_y4;
  assign f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa239_y4 = f_s_dadda_pg_rca32_fa239_y4;
  assign f_s_dadda_pg_rca32_fa249_y0 = f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa241_y4 ^ f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa240_y4;
  assign f_s_dadda_pg_rca32_fa249_y1 = f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa241_y4 & f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa240_y4;
  assign f_s_dadda_pg_rca32_fa249_y2 = f_s_dadda_pg_rca32_fa249_y0 ^ f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa239_y4;
  assign f_s_dadda_pg_rca32_fa249_y3 = f_s_dadda_pg_rca32_fa249_y0 & f_s_dadda_pg_rca32_fa249_f_s_dadda_pg_rca32_fa239_y4;
  assign f_s_dadda_pg_rca32_fa249_y4 = f_s_dadda_pg_rca32_fa249_y1 | f_s_dadda_pg_rca32_fa249_y3;
  assign f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa238_y4 = f_s_dadda_pg_rca32_fa238_y4;
  assign f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa237_y4 = f_s_dadda_pg_rca32_fa237_y4;
  assign f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa236_y4 = f_s_dadda_pg_rca32_fa236_y4;
  assign f_s_dadda_pg_rca32_fa250_y0 = f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa238_y4 ^ f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa237_y4;
  assign f_s_dadda_pg_rca32_fa250_y1 = f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa238_y4 & f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa237_y4;
  assign f_s_dadda_pg_rca32_fa250_y2 = f_s_dadda_pg_rca32_fa250_y0 ^ f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa236_y4;
  assign f_s_dadda_pg_rca32_fa250_y3 = f_s_dadda_pg_rca32_fa250_y0 & f_s_dadda_pg_rca32_fa250_f_s_dadda_pg_rca32_fa236_y4;
  assign f_s_dadda_pg_rca32_fa250_y4 = f_s_dadda_pg_rca32_fa250_y1 | f_s_dadda_pg_rca32_fa250_y3;
  assign f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa235_y4 = f_s_dadda_pg_rca32_fa235_y4;
  assign f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa234_y4 = f_s_dadda_pg_rca32_fa234_y4;
  assign f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa233_y4 = f_s_dadda_pg_rca32_fa233_y4;
  assign f_s_dadda_pg_rca32_fa251_y0 = f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa235_y4 ^ f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa234_y4;
  assign f_s_dadda_pg_rca32_fa251_y1 = f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa235_y4 & f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa234_y4;
  assign f_s_dadda_pg_rca32_fa251_y2 = f_s_dadda_pg_rca32_fa251_y0 ^ f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa233_y4;
  assign f_s_dadda_pg_rca32_fa251_y3 = f_s_dadda_pg_rca32_fa251_y0 & f_s_dadda_pg_rca32_fa251_f_s_dadda_pg_rca32_fa233_y4;
  assign f_s_dadda_pg_rca32_fa251_y4 = f_s_dadda_pg_rca32_fa251_y1 | f_s_dadda_pg_rca32_fa251_y3;
  assign f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa232_y4 = f_s_dadda_pg_rca32_fa232_y4;
  assign f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa231_y4 = f_s_dadda_pg_rca32_fa231_y4;
  assign f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa230_y4 = f_s_dadda_pg_rca32_fa230_y4;
  assign f_s_dadda_pg_rca32_fa252_y0 = f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa232_y4 ^ f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa231_y4;
  assign f_s_dadda_pg_rca32_fa252_y1 = f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa232_y4 & f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa231_y4;
  assign f_s_dadda_pg_rca32_fa252_y2 = f_s_dadda_pg_rca32_fa252_y0 ^ f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa230_y4;
  assign f_s_dadda_pg_rca32_fa252_y3 = f_s_dadda_pg_rca32_fa252_y0 & f_s_dadda_pg_rca32_fa252_f_s_dadda_pg_rca32_fa230_y4;
  assign f_s_dadda_pg_rca32_fa252_y4 = f_s_dadda_pg_rca32_fa252_y1 | f_s_dadda_pg_rca32_fa252_y3;
  assign f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa229_y4 = f_s_dadda_pg_rca32_fa229_y4;
  assign f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa228_y4 = f_s_dadda_pg_rca32_fa228_y4;
  assign f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa227_y4 = f_s_dadda_pg_rca32_fa227_y4;
  assign f_s_dadda_pg_rca32_fa253_y0 = f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa229_y4 ^ f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa228_y4;
  assign f_s_dadda_pg_rca32_fa253_y1 = f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa229_y4 & f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa228_y4;
  assign f_s_dadda_pg_rca32_fa253_y2 = f_s_dadda_pg_rca32_fa253_y0 ^ f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa227_y4;
  assign f_s_dadda_pg_rca32_fa253_y3 = f_s_dadda_pg_rca32_fa253_y0 & f_s_dadda_pg_rca32_fa253_f_s_dadda_pg_rca32_fa227_y4;
  assign f_s_dadda_pg_rca32_fa253_y4 = f_s_dadda_pg_rca32_fa253_y1 | f_s_dadda_pg_rca32_fa253_y3;
  assign f_s_dadda_pg_rca32_and_26_2_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_26_2_y0 = f_s_dadda_pg_rca32_and_26_2_a_26 & f_s_dadda_pg_rca32_and_26_2_b_2;
  assign f_s_dadda_pg_rca32_and_25_3_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_25_3_y0 = f_s_dadda_pg_rca32_and_25_3_a_25 & f_s_dadda_pg_rca32_and_25_3_b_3;
  assign f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_fa226_y4 = f_s_dadda_pg_rca32_fa226_y4;
  assign f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_and_26_2_y0 = f_s_dadda_pg_rca32_and_26_2_y0;
  assign f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_and_25_3_y0 = f_s_dadda_pg_rca32_and_25_3_y0;
  assign f_s_dadda_pg_rca32_fa254_y0 = f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_fa226_y4 ^ f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_and_26_2_y0;
  assign f_s_dadda_pg_rca32_fa254_y1 = f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_fa226_y4 & f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_and_26_2_y0;
  assign f_s_dadda_pg_rca32_fa254_y2 = f_s_dadda_pg_rca32_fa254_y0 ^ f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_and_25_3_y0;
  assign f_s_dadda_pg_rca32_fa254_y3 = f_s_dadda_pg_rca32_fa254_y0 & f_s_dadda_pg_rca32_fa254_f_s_dadda_pg_rca32_and_25_3_y0;
  assign f_s_dadda_pg_rca32_fa254_y4 = f_s_dadda_pg_rca32_fa254_y1 | f_s_dadda_pg_rca32_fa254_y3;
  assign f_s_dadda_pg_rca32_and_24_4_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_24_4_y0 = f_s_dadda_pg_rca32_and_24_4_a_24 & f_s_dadda_pg_rca32_and_24_4_b_4;
  assign f_s_dadda_pg_rca32_and_23_5_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_23_5_y0 = f_s_dadda_pg_rca32_and_23_5_a_23 & f_s_dadda_pg_rca32_and_23_5_b_5;
  assign f_s_dadda_pg_rca32_and_22_6_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_22_6_y0 = f_s_dadda_pg_rca32_and_22_6_a_22 & f_s_dadda_pg_rca32_and_22_6_b_6;
  assign f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_24_4_y0 = f_s_dadda_pg_rca32_and_24_4_y0;
  assign f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_23_5_y0 = f_s_dadda_pg_rca32_and_23_5_y0;
  assign f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_22_6_y0 = f_s_dadda_pg_rca32_and_22_6_y0;
  assign f_s_dadda_pg_rca32_fa255_y0 = f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_24_4_y0 ^ f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_23_5_y0;
  assign f_s_dadda_pg_rca32_fa255_y1 = f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_24_4_y0 & f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_23_5_y0;
  assign f_s_dadda_pg_rca32_fa255_y2 = f_s_dadda_pg_rca32_fa255_y0 ^ f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_22_6_y0;
  assign f_s_dadda_pg_rca32_fa255_y3 = f_s_dadda_pg_rca32_fa255_y0 & f_s_dadda_pg_rca32_fa255_f_s_dadda_pg_rca32_and_22_6_y0;
  assign f_s_dadda_pg_rca32_fa255_y4 = f_s_dadda_pg_rca32_fa255_y1 | f_s_dadda_pg_rca32_fa255_y3;
  assign f_s_dadda_pg_rca32_and_21_7_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_21_7_y0 = f_s_dadda_pg_rca32_and_21_7_a_21 & f_s_dadda_pg_rca32_and_21_7_b_7;
  assign f_s_dadda_pg_rca32_and_20_8_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_20_8_y0 = f_s_dadda_pg_rca32_and_20_8_a_20 & f_s_dadda_pg_rca32_and_20_8_b_8;
  assign f_s_dadda_pg_rca32_and_19_9_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_19_9_y0 = f_s_dadda_pg_rca32_and_19_9_a_19 & f_s_dadda_pg_rca32_and_19_9_b_9;
  assign f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_21_7_y0 = f_s_dadda_pg_rca32_and_21_7_y0;
  assign f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_20_8_y0 = f_s_dadda_pg_rca32_and_20_8_y0;
  assign f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_19_9_y0 = f_s_dadda_pg_rca32_and_19_9_y0;
  assign f_s_dadda_pg_rca32_fa256_y0 = f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_21_7_y0 ^ f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_20_8_y0;
  assign f_s_dadda_pg_rca32_fa256_y1 = f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_21_7_y0 & f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_20_8_y0;
  assign f_s_dadda_pg_rca32_fa256_y2 = f_s_dadda_pg_rca32_fa256_y0 ^ f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_19_9_y0;
  assign f_s_dadda_pg_rca32_fa256_y3 = f_s_dadda_pg_rca32_fa256_y0 & f_s_dadda_pg_rca32_fa256_f_s_dadda_pg_rca32_and_19_9_y0;
  assign f_s_dadda_pg_rca32_fa256_y4 = f_s_dadda_pg_rca32_fa256_y1 | f_s_dadda_pg_rca32_fa256_y3;
  assign f_s_dadda_pg_rca32_and_18_10_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_18_10_y0 = f_s_dadda_pg_rca32_and_18_10_a_18 & f_s_dadda_pg_rca32_and_18_10_b_10;
  assign f_s_dadda_pg_rca32_and_17_11_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_17_11_y0 = f_s_dadda_pg_rca32_and_17_11_a_17 & f_s_dadda_pg_rca32_and_17_11_b_11;
  assign f_s_dadda_pg_rca32_and_16_12_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_16_12_y0 = f_s_dadda_pg_rca32_and_16_12_a_16 & f_s_dadda_pg_rca32_and_16_12_b_12;
  assign f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_18_10_y0 = f_s_dadda_pg_rca32_and_18_10_y0;
  assign f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_17_11_y0 = f_s_dadda_pg_rca32_and_17_11_y0;
  assign f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_16_12_y0 = f_s_dadda_pg_rca32_and_16_12_y0;
  assign f_s_dadda_pg_rca32_fa257_y0 = f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_18_10_y0 ^ f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_17_11_y0;
  assign f_s_dadda_pg_rca32_fa257_y1 = f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_18_10_y0 & f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_17_11_y0;
  assign f_s_dadda_pg_rca32_fa257_y2 = f_s_dadda_pg_rca32_fa257_y0 ^ f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_16_12_y0;
  assign f_s_dadda_pg_rca32_fa257_y3 = f_s_dadda_pg_rca32_fa257_y0 & f_s_dadda_pg_rca32_fa257_f_s_dadda_pg_rca32_and_16_12_y0;
  assign f_s_dadda_pg_rca32_fa257_y4 = f_s_dadda_pg_rca32_fa257_y1 | f_s_dadda_pg_rca32_fa257_y3;
  assign f_s_dadda_pg_rca32_and_15_13_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_15_13_y0 = f_s_dadda_pg_rca32_and_15_13_a_15 & f_s_dadda_pg_rca32_and_15_13_b_13;
  assign f_s_dadda_pg_rca32_and_14_14_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_14_14_y0 = f_s_dadda_pg_rca32_and_14_14_a_14 & f_s_dadda_pg_rca32_and_14_14_b_14;
  assign f_s_dadda_pg_rca32_and_13_15_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_13_15_y0 = f_s_dadda_pg_rca32_and_13_15_a_13 & f_s_dadda_pg_rca32_and_13_15_b_15;
  assign f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_15_13_y0 = f_s_dadda_pg_rca32_and_15_13_y0;
  assign f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_14_14_y0 = f_s_dadda_pg_rca32_and_14_14_y0;
  assign f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_13_15_y0 = f_s_dadda_pg_rca32_and_13_15_y0;
  assign f_s_dadda_pg_rca32_fa258_y0 = f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_15_13_y0 ^ f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_14_14_y0;
  assign f_s_dadda_pg_rca32_fa258_y1 = f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_15_13_y0 & f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_14_14_y0;
  assign f_s_dadda_pg_rca32_fa258_y2 = f_s_dadda_pg_rca32_fa258_y0 ^ f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_13_15_y0;
  assign f_s_dadda_pg_rca32_fa258_y3 = f_s_dadda_pg_rca32_fa258_y0 & f_s_dadda_pg_rca32_fa258_f_s_dadda_pg_rca32_and_13_15_y0;
  assign f_s_dadda_pg_rca32_fa258_y4 = f_s_dadda_pg_rca32_fa258_y1 | f_s_dadda_pg_rca32_fa258_y3;
  assign f_s_dadda_pg_rca32_and_12_16_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_12_16_y0 = f_s_dadda_pg_rca32_and_12_16_a_12 & f_s_dadda_pg_rca32_and_12_16_b_16;
  assign f_s_dadda_pg_rca32_and_11_17_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_11_17_y0 = f_s_dadda_pg_rca32_and_11_17_a_11 & f_s_dadda_pg_rca32_and_11_17_b_17;
  assign f_s_dadda_pg_rca32_and_10_18_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_10_18_y0 = f_s_dadda_pg_rca32_and_10_18_a_10 & f_s_dadda_pg_rca32_and_10_18_b_18;
  assign f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_12_16_y0 = f_s_dadda_pg_rca32_and_12_16_y0;
  assign f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_11_17_y0 = f_s_dadda_pg_rca32_and_11_17_y0;
  assign f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_10_18_y0 = f_s_dadda_pg_rca32_and_10_18_y0;
  assign f_s_dadda_pg_rca32_fa259_y0 = f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_12_16_y0 ^ f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_11_17_y0;
  assign f_s_dadda_pg_rca32_fa259_y1 = f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_12_16_y0 & f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_11_17_y0;
  assign f_s_dadda_pg_rca32_fa259_y2 = f_s_dadda_pg_rca32_fa259_y0 ^ f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_10_18_y0;
  assign f_s_dadda_pg_rca32_fa259_y3 = f_s_dadda_pg_rca32_fa259_y0 & f_s_dadda_pg_rca32_fa259_f_s_dadda_pg_rca32_and_10_18_y0;
  assign f_s_dadda_pg_rca32_fa259_y4 = f_s_dadda_pg_rca32_fa259_y1 | f_s_dadda_pg_rca32_fa259_y3;
  assign f_s_dadda_pg_rca32_and_9_19_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_9_19_y0 = f_s_dadda_pg_rca32_and_9_19_a_9 & f_s_dadda_pg_rca32_and_9_19_b_19;
  assign f_s_dadda_pg_rca32_and_8_20_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_8_20_y0 = f_s_dadda_pg_rca32_and_8_20_a_8 & f_s_dadda_pg_rca32_and_8_20_b_20;
  assign f_s_dadda_pg_rca32_and_7_21_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_7_21_y0 = f_s_dadda_pg_rca32_and_7_21_a_7 & f_s_dadda_pg_rca32_and_7_21_b_21;
  assign f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_9_19_y0 = f_s_dadda_pg_rca32_and_9_19_y0;
  assign f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_8_20_y0 = f_s_dadda_pg_rca32_and_8_20_y0;
  assign f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_7_21_y0 = f_s_dadda_pg_rca32_and_7_21_y0;
  assign f_s_dadda_pg_rca32_fa260_y0 = f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_9_19_y0 ^ f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_8_20_y0;
  assign f_s_dadda_pg_rca32_fa260_y1 = f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_9_19_y0 & f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_8_20_y0;
  assign f_s_dadda_pg_rca32_fa260_y2 = f_s_dadda_pg_rca32_fa260_y0 ^ f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_7_21_y0;
  assign f_s_dadda_pg_rca32_fa260_y3 = f_s_dadda_pg_rca32_fa260_y0 & f_s_dadda_pg_rca32_fa260_f_s_dadda_pg_rca32_and_7_21_y0;
  assign f_s_dadda_pg_rca32_fa260_y4 = f_s_dadda_pg_rca32_fa260_y1 | f_s_dadda_pg_rca32_fa260_y3;
  assign f_s_dadda_pg_rca32_and_6_22_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_6_22_y0 = f_s_dadda_pg_rca32_and_6_22_a_6 & f_s_dadda_pg_rca32_and_6_22_b_22;
  assign f_s_dadda_pg_rca32_and_5_23_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_5_23_y0 = f_s_dadda_pg_rca32_and_5_23_a_5 & f_s_dadda_pg_rca32_and_5_23_b_23;
  assign f_s_dadda_pg_rca32_and_4_24_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_4_24_y0 = f_s_dadda_pg_rca32_and_4_24_a_4 & f_s_dadda_pg_rca32_and_4_24_b_24;
  assign f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_6_22_y0 = f_s_dadda_pg_rca32_and_6_22_y0;
  assign f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_5_23_y0 = f_s_dadda_pg_rca32_and_5_23_y0;
  assign f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_4_24_y0 = f_s_dadda_pg_rca32_and_4_24_y0;
  assign f_s_dadda_pg_rca32_fa261_y0 = f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_6_22_y0 ^ f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_5_23_y0;
  assign f_s_dadda_pg_rca32_fa261_y1 = f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_6_22_y0 & f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_5_23_y0;
  assign f_s_dadda_pg_rca32_fa261_y2 = f_s_dadda_pg_rca32_fa261_y0 ^ f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_4_24_y0;
  assign f_s_dadda_pg_rca32_fa261_y3 = f_s_dadda_pg_rca32_fa261_y0 & f_s_dadda_pg_rca32_fa261_f_s_dadda_pg_rca32_and_4_24_y0;
  assign f_s_dadda_pg_rca32_fa261_y4 = f_s_dadda_pg_rca32_fa261_y1 | f_s_dadda_pg_rca32_fa261_y3;
  assign f_s_dadda_pg_rca32_and_3_25_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_3_25_y0 = f_s_dadda_pg_rca32_and_3_25_a_3 & f_s_dadda_pg_rca32_and_3_25_b_25;
  assign f_s_dadda_pg_rca32_and_2_26_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_2_26_y0 = f_s_dadda_pg_rca32_and_2_26_a_2 & f_s_dadda_pg_rca32_and_2_26_b_26;
  assign f_s_dadda_pg_rca32_and_1_27_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_1_27_y0 = f_s_dadda_pg_rca32_and_1_27_a_1 & f_s_dadda_pg_rca32_and_1_27_b_27;
  assign f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_3_25_y0 = f_s_dadda_pg_rca32_and_3_25_y0;
  assign f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_2_26_y0 = f_s_dadda_pg_rca32_and_2_26_y0;
  assign f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_1_27_y0 = f_s_dadda_pg_rca32_and_1_27_y0;
  assign f_s_dadda_pg_rca32_fa262_y0 = f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_3_25_y0 ^ f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_2_26_y0;
  assign f_s_dadda_pg_rca32_fa262_y1 = f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_3_25_y0 & f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_2_26_y0;
  assign f_s_dadda_pg_rca32_fa262_y2 = f_s_dadda_pg_rca32_fa262_y0 ^ f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_1_27_y0;
  assign f_s_dadda_pg_rca32_fa262_y3 = f_s_dadda_pg_rca32_fa262_y0 & f_s_dadda_pg_rca32_fa262_f_s_dadda_pg_rca32_and_1_27_y0;
  assign f_s_dadda_pg_rca32_fa262_y4 = f_s_dadda_pg_rca32_fa262_y1 | f_s_dadda_pg_rca32_fa262_y3;
  assign f_s_dadda_pg_rca32_and_0_28_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_0_28_y0 = f_s_dadda_pg_rca32_and_0_28_a_0 & f_s_dadda_pg_rca32_and_0_28_b_28;
  assign f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_and_0_28_y0 = f_s_dadda_pg_rca32_and_0_28_y0;
  assign f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_ha0_y0 = f_s_dadda_pg_rca32_ha0_y0;
  assign f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_fa247_y2 = f_s_dadda_pg_rca32_fa247_y2;
  assign f_s_dadda_pg_rca32_fa263_y0 = f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_and_0_28_y0 ^ f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_ha0_y0;
  assign f_s_dadda_pg_rca32_fa263_y1 = f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_and_0_28_y0 & f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_ha0_y0;
  assign f_s_dadda_pg_rca32_fa263_y2 = f_s_dadda_pg_rca32_fa263_y0 ^ f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_fa247_y2;
  assign f_s_dadda_pg_rca32_fa263_y3 = f_s_dadda_pg_rca32_fa263_y0 & f_s_dadda_pg_rca32_fa263_f_s_dadda_pg_rca32_fa247_y2;
  assign f_s_dadda_pg_rca32_fa263_y4 = f_s_dadda_pg_rca32_fa263_y1 | f_s_dadda_pg_rca32_fa263_y3;
  assign f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa248_y2 = f_s_dadda_pg_rca32_fa248_y2;
  assign f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa249_y2 = f_s_dadda_pg_rca32_fa249_y2;
  assign f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa250_y2 = f_s_dadda_pg_rca32_fa250_y2;
  assign f_s_dadda_pg_rca32_fa264_y0 = f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa248_y2 ^ f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa249_y2;
  assign f_s_dadda_pg_rca32_fa264_y1 = f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa248_y2 & f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa249_y2;
  assign f_s_dadda_pg_rca32_fa264_y2 = f_s_dadda_pg_rca32_fa264_y0 ^ f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa250_y2;
  assign f_s_dadda_pg_rca32_fa264_y3 = f_s_dadda_pg_rca32_fa264_y0 & f_s_dadda_pg_rca32_fa264_f_s_dadda_pg_rca32_fa250_y2;
  assign f_s_dadda_pg_rca32_fa264_y4 = f_s_dadda_pg_rca32_fa264_y1 | f_s_dadda_pg_rca32_fa264_y3;
  assign f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa251_y2 = f_s_dadda_pg_rca32_fa251_y2;
  assign f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa252_y2 = f_s_dadda_pg_rca32_fa252_y2;
  assign f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa253_y2 = f_s_dadda_pg_rca32_fa253_y2;
  assign f_s_dadda_pg_rca32_fa265_y0 = f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa251_y2 ^ f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa252_y2;
  assign f_s_dadda_pg_rca32_fa265_y1 = f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa251_y2 & f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa252_y2;
  assign f_s_dadda_pg_rca32_fa265_y2 = f_s_dadda_pg_rca32_fa265_y0 ^ f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa253_y2;
  assign f_s_dadda_pg_rca32_fa265_y3 = f_s_dadda_pg_rca32_fa265_y0 & f_s_dadda_pg_rca32_fa265_f_s_dadda_pg_rca32_fa253_y2;
  assign f_s_dadda_pg_rca32_fa265_y4 = f_s_dadda_pg_rca32_fa265_y1 | f_s_dadda_pg_rca32_fa265_y3;
  assign f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa254_y2 = f_s_dadda_pg_rca32_fa254_y2;
  assign f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa255_y2 = f_s_dadda_pg_rca32_fa255_y2;
  assign f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa256_y2 = f_s_dadda_pg_rca32_fa256_y2;
  assign f_s_dadda_pg_rca32_fa266_y0 = f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa254_y2 ^ f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa255_y2;
  assign f_s_dadda_pg_rca32_fa266_y1 = f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa254_y2 & f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa255_y2;
  assign f_s_dadda_pg_rca32_fa266_y2 = f_s_dadda_pg_rca32_fa266_y0 ^ f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa256_y2;
  assign f_s_dadda_pg_rca32_fa266_y3 = f_s_dadda_pg_rca32_fa266_y0 & f_s_dadda_pg_rca32_fa266_f_s_dadda_pg_rca32_fa256_y2;
  assign f_s_dadda_pg_rca32_fa266_y4 = f_s_dadda_pg_rca32_fa266_y1 | f_s_dadda_pg_rca32_fa266_y3;
  assign f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa257_y2 = f_s_dadda_pg_rca32_fa257_y2;
  assign f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa258_y2 = f_s_dadda_pg_rca32_fa258_y2;
  assign f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa259_y2 = f_s_dadda_pg_rca32_fa259_y2;
  assign f_s_dadda_pg_rca32_fa267_y0 = f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa257_y2 ^ f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa258_y2;
  assign f_s_dadda_pg_rca32_fa267_y1 = f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa257_y2 & f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa258_y2;
  assign f_s_dadda_pg_rca32_fa267_y2 = f_s_dadda_pg_rca32_fa267_y0 ^ f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa259_y2;
  assign f_s_dadda_pg_rca32_fa267_y3 = f_s_dadda_pg_rca32_fa267_y0 & f_s_dadda_pg_rca32_fa267_f_s_dadda_pg_rca32_fa259_y2;
  assign f_s_dadda_pg_rca32_fa267_y4 = f_s_dadda_pg_rca32_fa267_y1 | f_s_dadda_pg_rca32_fa267_y3;
  assign f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa260_y2 = f_s_dadda_pg_rca32_fa260_y2;
  assign f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa261_y2 = f_s_dadda_pg_rca32_fa261_y2;
  assign f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa262_y2 = f_s_dadda_pg_rca32_fa262_y2;
  assign f_s_dadda_pg_rca32_fa268_y0 = f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa260_y2 ^ f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa261_y2;
  assign f_s_dadda_pg_rca32_fa268_y1 = f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa260_y2 & f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa261_y2;
  assign f_s_dadda_pg_rca32_fa268_y2 = f_s_dadda_pg_rca32_fa268_y0 ^ f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa262_y2;
  assign f_s_dadda_pg_rca32_fa268_y3 = f_s_dadda_pg_rca32_fa268_y0 & f_s_dadda_pg_rca32_fa268_f_s_dadda_pg_rca32_fa262_y2;
  assign f_s_dadda_pg_rca32_fa268_y4 = f_s_dadda_pg_rca32_fa268_y1 | f_s_dadda_pg_rca32_fa268_y3;
  assign f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa268_y4 = f_s_dadda_pg_rca32_fa268_y4;
  assign f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa267_y4 = f_s_dadda_pg_rca32_fa267_y4;
  assign f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa266_y4 = f_s_dadda_pg_rca32_fa266_y4;
  assign f_s_dadda_pg_rca32_fa269_y0 = f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa268_y4 ^ f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa267_y4;
  assign f_s_dadda_pg_rca32_fa269_y1 = f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa268_y4 & f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa267_y4;
  assign f_s_dadda_pg_rca32_fa269_y2 = f_s_dadda_pg_rca32_fa269_y0 ^ f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa266_y4;
  assign f_s_dadda_pg_rca32_fa269_y3 = f_s_dadda_pg_rca32_fa269_y0 & f_s_dadda_pg_rca32_fa269_f_s_dadda_pg_rca32_fa266_y4;
  assign f_s_dadda_pg_rca32_fa269_y4 = f_s_dadda_pg_rca32_fa269_y1 | f_s_dadda_pg_rca32_fa269_y3;
  assign f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa265_y4 = f_s_dadda_pg_rca32_fa265_y4;
  assign f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa264_y4 = f_s_dadda_pg_rca32_fa264_y4;
  assign f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa263_y4 = f_s_dadda_pg_rca32_fa263_y4;
  assign f_s_dadda_pg_rca32_fa270_y0 = f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa265_y4 ^ f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa264_y4;
  assign f_s_dadda_pg_rca32_fa270_y1 = f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa265_y4 & f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa264_y4;
  assign f_s_dadda_pg_rca32_fa270_y2 = f_s_dadda_pg_rca32_fa270_y0 ^ f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa263_y4;
  assign f_s_dadda_pg_rca32_fa270_y3 = f_s_dadda_pg_rca32_fa270_y0 & f_s_dadda_pg_rca32_fa270_f_s_dadda_pg_rca32_fa263_y4;
  assign f_s_dadda_pg_rca32_fa270_y4 = f_s_dadda_pg_rca32_fa270_y1 | f_s_dadda_pg_rca32_fa270_y3;
  assign f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa262_y4 = f_s_dadda_pg_rca32_fa262_y4;
  assign f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa261_y4 = f_s_dadda_pg_rca32_fa261_y4;
  assign f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa260_y4 = f_s_dadda_pg_rca32_fa260_y4;
  assign f_s_dadda_pg_rca32_fa271_y0 = f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa262_y4 ^ f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa261_y4;
  assign f_s_dadda_pg_rca32_fa271_y1 = f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa262_y4 & f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa261_y4;
  assign f_s_dadda_pg_rca32_fa271_y2 = f_s_dadda_pg_rca32_fa271_y0 ^ f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa260_y4;
  assign f_s_dadda_pg_rca32_fa271_y3 = f_s_dadda_pg_rca32_fa271_y0 & f_s_dadda_pg_rca32_fa271_f_s_dadda_pg_rca32_fa260_y4;
  assign f_s_dadda_pg_rca32_fa271_y4 = f_s_dadda_pg_rca32_fa271_y1 | f_s_dadda_pg_rca32_fa271_y3;
  assign f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa259_y4 = f_s_dadda_pg_rca32_fa259_y4;
  assign f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa258_y4 = f_s_dadda_pg_rca32_fa258_y4;
  assign f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa257_y4 = f_s_dadda_pg_rca32_fa257_y4;
  assign f_s_dadda_pg_rca32_fa272_y0 = f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa259_y4 ^ f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa258_y4;
  assign f_s_dadda_pg_rca32_fa272_y1 = f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa259_y4 & f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa258_y4;
  assign f_s_dadda_pg_rca32_fa272_y2 = f_s_dadda_pg_rca32_fa272_y0 ^ f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa257_y4;
  assign f_s_dadda_pg_rca32_fa272_y3 = f_s_dadda_pg_rca32_fa272_y0 & f_s_dadda_pg_rca32_fa272_f_s_dadda_pg_rca32_fa257_y4;
  assign f_s_dadda_pg_rca32_fa272_y4 = f_s_dadda_pg_rca32_fa272_y1 | f_s_dadda_pg_rca32_fa272_y3;
  assign f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa256_y4 = f_s_dadda_pg_rca32_fa256_y4;
  assign f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa255_y4 = f_s_dadda_pg_rca32_fa255_y4;
  assign f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa254_y4 = f_s_dadda_pg_rca32_fa254_y4;
  assign f_s_dadda_pg_rca32_fa273_y0 = f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa256_y4 ^ f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa255_y4;
  assign f_s_dadda_pg_rca32_fa273_y1 = f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa256_y4 & f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa255_y4;
  assign f_s_dadda_pg_rca32_fa273_y2 = f_s_dadda_pg_rca32_fa273_y0 ^ f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa254_y4;
  assign f_s_dadda_pg_rca32_fa273_y3 = f_s_dadda_pg_rca32_fa273_y0 & f_s_dadda_pg_rca32_fa273_f_s_dadda_pg_rca32_fa254_y4;
  assign f_s_dadda_pg_rca32_fa273_y4 = f_s_dadda_pg_rca32_fa273_y1 | f_s_dadda_pg_rca32_fa273_y3;
  assign f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa253_y4 = f_s_dadda_pg_rca32_fa253_y4;
  assign f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa252_y4 = f_s_dadda_pg_rca32_fa252_y4;
  assign f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa251_y4 = f_s_dadda_pg_rca32_fa251_y4;
  assign f_s_dadda_pg_rca32_fa274_y0 = f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa253_y4 ^ f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa252_y4;
  assign f_s_dadda_pg_rca32_fa274_y1 = f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa253_y4 & f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa252_y4;
  assign f_s_dadda_pg_rca32_fa274_y2 = f_s_dadda_pg_rca32_fa274_y0 ^ f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa251_y4;
  assign f_s_dadda_pg_rca32_fa274_y3 = f_s_dadda_pg_rca32_fa274_y0 & f_s_dadda_pg_rca32_fa274_f_s_dadda_pg_rca32_fa251_y4;
  assign f_s_dadda_pg_rca32_fa274_y4 = f_s_dadda_pg_rca32_fa274_y1 | f_s_dadda_pg_rca32_fa274_y3;
  assign f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa250_y4 = f_s_dadda_pg_rca32_fa250_y4;
  assign f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa249_y4 = f_s_dadda_pg_rca32_fa249_y4;
  assign f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa248_y4 = f_s_dadda_pg_rca32_fa248_y4;
  assign f_s_dadda_pg_rca32_fa275_y0 = f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa250_y4 ^ f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa249_y4;
  assign f_s_dadda_pg_rca32_fa275_y1 = f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa250_y4 & f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa249_y4;
  assign f_s_dadda_pg_rca32_fa275_y2 = f_s_dadda_pg_rca32_fa275_y0 ^ f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa248_y4;
  assign f_s_dadda_pg_rca32_fa275_y3 = f_s_dadda_pg_rca32_fa275_y0 & f_s_dadda_pg_rca32_fa275_f_s_dadda_pg_rca32_fa248_y4;
  assign f_s_dadda_pg_rca32_fa275_y4 = f_s_dadda_pg_rca32_fa275_y1 | f_s_dadda_pg_rca32_fa275_y3;
  assign f_s_dadda_pg_rca32_and_25_4_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_25_4_y0 = f_s_dadda_pg_rca32_and_25_4_a_25 & f_s_dadda_pg_rca32_and_25_4_b_4;
  assign f_s_dadda_pg_rca32_and_24_5_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_24_5_y0 = f_s_dadda_pg_rca32_and_24_5_a_24 & f_s_dadda_pg_rca32_and_24_5_b_5;
  assign f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_fa247_y4 = f_s_dadda_pg_rca32_fa247_y4;
  assign f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_and_25_4_y0 = f_s_dadda_pg_rca32_and_25_4_y0;
  assign f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_and_24_5_y0 = f_s_dadda_pg_rca32_and_24_5_y0;
  assign f_s_dadda_pg_rca32_fa276_y0 = f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_fa247_y4 ^ f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_and_25_4_y0;
  assign f_s_dadda_pg_rca32_fa276_y1 = f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_fa247_y4 & f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_and_25_4_y0;
  assign f_s_dadda_pg_rca32_fa276_y2 = f_s_dadda_pg_rca32_fa276_y0 ^ f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_and_24_5_y0;
  assign f_s_dadda_pg_rca32_fa276_y3 = f_s_dadda_pg_rca32_fa276_y0 & f_s_dadda_pg_rca32_fa276_f_s_dadda_pg_rca32_and_24_5_y0;
  assign f_s_dadda_pg_rca32_fa276_y4 = f_s_dadda_pg_rca32_fa276_y1 | f_s_dadda_pg_rca32_fa276_y3;
  assign f_s_dadda_pg_rca32_and_23_6_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_23_6_y0 = f_s_dadda_pg_rca32_and_23_6_a_23 & f_s_dadda_pg_rca32_and_23_6_b_6;
  assign f_s_dadda_pg_rca32_and_22_7_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_22_7_y0 = f_s_dadda_pg_rca32_and_22_7_a_22 & f_s_dadda_pg_rca32_and_22_7_b_7;
  assign f_s_dadda_pg_rca32_and_21_8_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_21_8_y0 = f_s_dadda_pg_rca32_and_21_8_a_21 & f_s_dadda_pg_rca32_and_21_8_b_8;
  assign f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_23_6_y0 = f_s_dadda_pg_rca32_and_23_6_y0;
  assign f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_22_7_y0 = f_s_dadda_pg_rca32_and_22_7_y0;
  assign f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_21_8_y0 = f_s_dadda_pg_rca32_and_21_8_y0;
  assign f_s_dadda_pg_rca32_fa277_y0 = f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_23_6_y0 ^ f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_22_7_y0;
  assign f_s_dadda_pg_rca32_fa277_y1 = f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_23_6_y0 & f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_22_7_y0;
  assign f_s_dadda_pg_rca32_fa277_y2 = f_s_dadda_pg_rca32_fa277_y0 ^ f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_21_8_y0;
  assign f_s_dadda_pg_rca32_fa277_y3 = f_s_dadda_pg_rca32_fa277_y0 & f_s_dadda_pg_rca32_fa277_f_s_dadda_pg_rca32_and_21_8_y0;
  assign f_s_dadda_pg_rca32_fa277_y4 = f_s_dadda_pg_rca32_fa277_y1 | f_s_dadda_pg_rca32_fa277_y3;
  assign f_s_dadda_pg_rca32_and_20_9_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_20_9_y0 = f_s_dadda_pg_rca32_and_20_9_a_20 & f_s_dadda_pg_rca32_and_20_9_b_9;
  assign f_s_dadda_pg_rca32_and_19_10_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_19_10_y0 = f_s_dadda_pg_rca32_and_19_10_a_19 & f_s_dadda_pg_rca32_and_19_10_b_10;
  assign f_s_dadda_pg_rca32_and_18_11_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_18_11_y0 = f_s_dadda_pg_rca32_and_18_11_a_18 & f_s_dadda_pg_rca32_and_18_11_b_11;
  assign f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_20_9_y0 = f_s_dadda_pg_rca32_and_20_9_y0;
  assign f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_19_10_y0 = f_s_dadda_pg_rca32_and_19_10_y0;
  assign f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_18_11_y0 = f_s_dadda_pg_rca32_and_18_11_y0;
  assign f_s_dadda_pg_rca32_fa278_y0 = f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_20_9_y0 ^ f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_19_10_y0;
  assign f_s_dadda_pg_rca32_fa278_y1 = f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_20_9_y0 & f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_19_10_y0;
  assign f_s_dadda_pg_rca32_fa278_y2 = f_s_dadda_pg_rca32_fa278_y0 ^ f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_18_11_y0;
  assign f_s_dadda_pg_rca32_fa278_y3 = f_s_dadda_pg_rca32_fa278_y0 & f_s_dadda_pg_rca32_fa278_f_s_dadda_pg_rca32_and_18_11_y0;
  assign f_s_dadda_pg_rca32_fa278_y4 = f_s_dadda_pg_rca32_fa278_y1 | f_s_dadda_pg_rca32_fa278_y3;
  assign f_s_dadda_pg_rca32_and_17_12_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_17_12_y0 = f_s_dadda_pg_rca32_and_17_12_a_17 & f_s_dadda_pg_rca32_and_17_12_b_12;
  assign f_s_dadda_pg_rca32_and_16_13_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_16_13_y0 = f_s_dadda_pg_rca32_and_16_13_a_16 & f_s_dadda_pg_rca32_and_16_13_b_13;
  assign f_s_dadda_pg_rca32_and_15_14_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_15_14_y0 = f_s_dadda_pg_rca32_and_15_14_a_15 & f_s_dadda_pg_rca32_and_15_14_b_14;
  assign f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_17_12_y0 = f_s_dadda_pg_rca32_and_17_12_y0;
  assign f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_16_13_y0 = f_s_dadda_pg_rca32_and_16_13_y0;
  assign f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_15_14_y0 = f_s_dadda_pg_rca32_and_15_14_y0;
  assign f_s_dadda_pg_rca32_fa279_y0 = f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_17_12_y0 ^ f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_16_13_y0;
  assign f_s_dadda_pg_rca32_fa279_y1 = f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_17_12_y0 & f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_16_13_y0;
  assign f_s_dadda_pg_rca32_fa279_y2 = f_s_dadda_pg_rca32_fa279_y0 ^ f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_15_14_y0;
  assign f_s_dadda_pg_rca32_fa279_y3 = f_s_dadda_pg_rca32_fa279_y0 & f_s_dadda_pg_rca32_fa279_f_s_dadda_pg_rca32_and_15_14_y0;
  assign f_s_dadda_pg_rca32_fa279_y4 = f_s_dadda_pg_rca32_fa279_y1 | f_s_dadda_pg_rca32_fa279_y3;
  assign f_s_dadda_pg_rca32_and_14_15_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_14_15_y0 = f_s_dadda_pg_rca32_and_14_15_a_14 & f_s_dadda_pg_rca32_and_14_15_b_15;
  assign f_s_dadda_pg_rca32_and_13_16_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_13_16_y0 = f_s_dadda_pg_rca32_and_13_16_a_13 & f_s_dadda_pg_rca32_and_13_16_b_16;
  assign f_s_dadda_pg_rca32_and_12_17_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_12_17_y0 = f_s_dadda_pg_rca32_and_12_17_a_12 & f_s_dadda_pg_rca32_and_12_17_b_17;
  assign f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_14_15_y0 = f_s_dadda_pg_rca32_and_14_15_y0;
  assign f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_13_16_y0 = f_s_dadda_pg_rca32_and_13_16_y0;
  assign f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_12_17_y0 = f_s_dadda_pg_rca32_and_12_17_y0;
  assign f_s_dadda_pg_rca32_fa280_y0 = f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_14_15_y0 ^ f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_13_16_y0;
  assign f_s_dadda_pg_rca32_fa280_y1 = f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_14_15_y0 & f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_13_16_y0;
  assign f_s_dadda_pg_rca32_fa280_y2 = f_s_dadda_pg_rca32_fa280_y0 ^ f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_12_17_y0;
  assign f_s_dadda_pg_rca32_fa280_y3 = f_s_dadda_pg_rca32_fa280_y0 & f_s_dadda_pg_rca32_fa280_f_s_dadda_pg_rca32_and_12_17_y0;
  assign f_s_dadda_pg_rca32_fa280_y4 = f_s_dadda_pg_rca32_fa280_y1 | f_s_dadda_pg_rca32_fa280_y3;
  assign f_s_dadda_pg_rca32_and_11_18_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_11_18_y0 = f_s_dadda_pg_rca32_and_11_18_a_11 & f_s_dadda_pg_rca32_and_11_18_b_18;
  assign f_s_dadda_pg_rca32_and_10_19_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_10_19_y0 = f_s_dadda_pg_rca32_and_10_19_a_10 & f_s_dadda_pg_rca32_and_10_19_b_19;
  assign f_s_dadda_pg_rca32_and_9_20_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_9_20_y0 = f_s_dadda_pg_rca32_and_9_20_a_9 & f_s_dadda_pg_rca32_and_9_20_b_20;
  assign f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_11_18_y0 = f_s_dadda_pg_rca32_and_11_18_y0;
  assign f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_10_19_y0 = f_s_dadda_pg_rca32_and_10_19_y0;
  assign f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_9_20_y0 = f_s_dadda_pg_rca32_and_9_20_y0;
  assign f_s_dadda_pg_rca32_fa281_y0 = f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_11_18_y0 ^ f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_10_19_y0;
  assign f_s_dadda_pg_rca32_fa281_y1 = f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_11_18_y0 & f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_10_19_y0;
  assign f_s_dadda_pg_rca32_fa281_y2 = f_s_dadda_pg_rca32_fa281_y0 ^ f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_9_20_y0;
  assign f_s_dadda_pg_rca32_fa281_y3 = f_s_dadda_pg_rca32_fa281_y0 & f_s_dadda_pg_rca32_fa281_f_s_dadda_pg_rca32_and_9_20_y0;
  assign f_s_dadda_pg_rca32_fa281_y4 = f_s_dadda_pg_rca32_fa281_y1 | f_s_dadda_pg_rca32_fa281_y3;
  assign f_s_dadda_pg_rca32_and_8_21_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_8_21_y0 = f_s_dadda_pg_rca32_and_8_21_a_8 & f_s_dadda_pg_rca32_and_8_21_b_21;
  assign f_s_dadda_pg_rca32_and_7_22_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_7_22_y0 = f_s_dadda_pg_rca32_and_7_22_a_7 & f_s_dadda_pg_rca32_and_7_22_b_22;
  assign f_s_dadda_pg_rca32_and_6_23_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_6_23_y0 = f_s_dadda_pg_rca32_and_6_23_a_6 & f_s_dadda_pg_rca32_and_6_23_b_23;
  assign f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_8_21_y0 = f_s_dadda_pg_rca32_and_8_21_y0;
  assign f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_7_22_y0 = f_s_dadda_pg_rca32_and_7_22_y0;
  assign f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_6_23_y0 = f_s_dadda_pg_rca32_and_6_23_y0;
  assign f_s_dadda_pg_rca32_fa282_y0 = f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_8_21_y0 ^ f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_7_22_y0;
  assign f_s_dadda_pg_rca32_fa282_y1 = f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_8_21_y0 & f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_7_22_y0;
  assign f_s_dadda_pg_rca32_fa282_y2 = f_s_dadda_pg_rca32_fa282_y0 ^ f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_6_23_y0;
  assign f_s_dadda_pg_rca32_fa282_y3 = f_s_dadda_pg_rca32_fa282_y0 & f_s_dadda_pg_rca32_fa282_f_s_dadda_pg_rca32_and_6_23_y0;
  assign f_s_dadda_pg_rca32_fa282_y4 = f_s_dadda_pg_rca32_fa282_y1 | f_s_dadda_pg_rca32_fa282_y3;
  assign f_s_dadda_pg_rca32_and_5_24_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_5_24_y0 = f_s_dadda_pg_rca32_and_5_24_a_5 & f_s_dadda_pg_rca32_and_5_24_b_24;
  assign f_s_dadda_pg_rca32_and_4_25_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_4_25_y0 = f_s_dadda_pg_rca32_and_4_25_a_4 & f_s_dadda_pg_rca32_and_4_25_b_25;
  assign f_s_dadda_pg_rca32_and_3_26_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_3_26_y0 = f_s_dadda_pg_rca32_and_3_26_a_3 & f_s_dadda_pg_rca32_and_3_26_b_26;
  assign f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_5_24_y0 = f_s_dadda_pg_rca32_and_5_24_y0;
  assign f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_4_25_y0 = f_s_dadda_pg_rca32_and_4_25_y0;
  assign f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_3_26_y0 = f_s_dadda_pg_rca32_and_3_26_y0;
  assign f_s_dadda_pg_rca32_fa283_y0 = f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_5_24_y0 ^ f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_4_25_y0;
  assign f_s_dadda_pg_rca32_fa283_y1 = f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_5_24_y0 & f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_4_25_y0;
  assign f_s_dadda_pg_rca32_fa283_y2 = f_s_dadda_pg_rca32_fa283_y0 ^ f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_3_26_y0;
  assign f_s_dadda_pg_rca32_fa283_y3 = f_s_dadda_pg_rca32_fa283_y0 & f_s_dadda_pg_rca32_fa283_f_s_dadda_pg_rca32_and_3_26_y0;
  assign f_s_dadda_pg_rca32_fa283_y4 = f_s_dadda_pg_rca32_fa283_y1 | f_s_dadda_pg_rca32_fa283_y3;
  assign f_s_dadda_pg_rca32_and_2_27_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_2_27_y0 = f_s_dadda_pg_rca32_and_2_27_a_2 & f_s_dadda_pg_rca32_and_2_27_b_27;
  assign f_s_dadda_pg_rca32_and_1_28_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_1_28_y0 = f_s_dadda_pg_rca32_and_1_28_a_1 & f_s_dadda_pg_rca32_and_1_28_b_28;
  assign f_s_dadda_pg_rca32_and_0_29_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_0_29_y0 = f_s_dadda_pg_rca32_and_0_29_a_0 & f_s_dadda_pg_rca32_and_0_29_b_29;
  assign f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_2_27_y0 = f_s_dadda_pg_rca32_and_2_27_y0;
  assign f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_1_28_y0 = f_s_dadda_pg_rca32_and_1_28_y0;
  assign f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_0_29_y0 = f_s_dadda_pg_rca32_and_0_29_y0;
  assign f_s_dadda_pg_rca32_fa284_y0 = f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_2_27_y0 ^ f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_1_28_y0;
  assign f_s_dadda_pg_rca32_fa284_y1 = f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_2_27_y0 & f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_1_28_y0;
  assign f_s_dadda_pg_rca32_fa284_y2 = f_s_dadda_pg_rca32_fa284_y0 ^ f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_0_29_y0;
  assign f_s_dadda_pg_rca32_fa284_y3 = f_s_dadda_pg_rca32_fa284_y0 & f_s_dadda_pg_rca32_fa284_f_s_dadda_pg_rca32_and_0_29_y0;
  assign f_s_dadda_pg_rca32_fa284_y4 = f_s_dadda_pg_rca32_fa284_y1 | f_s_dadda_pg_rca32_fa284_y3;
  assign f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_fa0_y2 = f_s_dadda_pg_rca32_fa0_y2;
  assign f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_ha1_y0 = f_s_dadda_pg_rca32_ha1_y0;
  assign f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_fa269_y2 = f_s_dadda_pg_rca32_fa269_y2;
  assign f_s_dadda_pg_rca32_fa285_y0 = f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_fa0_y2 ^ f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_ha1_y0;
  assign f_s_dadda_pg_rca32_fa285_y1 = f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_fa0_y2 & f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_ha1_y0;
  assign f_s_dadda_pg_rca32_fa285_y2 = f_s_dadda_pg_rca32_fa285_y0 ^ f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_fa269_y2;
  assign f_s_dadda_pg_rca32_fa285_y3 = f_s_dadda_pg_rca32_fa285_y0 & f_s_dadda_pg_rca32_fa285_f_s_dadda_pg_rca32_fa269_y2;
  assign f_s_dadda_pg_rca32_fa285_y4 = f_s_dadda_pg_rca32_fa285_y1 | f_s_dadda_pg_rca32_fa285_y3;
  assign f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa270_y2 = f_s_dadda_pg_rca32_fa270_y2;
  assign f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa271_y2 = f_s_dadda_pg_rca32_fa271_y2;
  assign f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa272_y2 = f_s_dadda_pg_rca32_fa272_y2;
  assign f_s_dadda_pg_rca32_fa286_y0 = f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa270_y2 ^ f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa271_y2;
  assign f_s_dadda_pg_rca32_fa286_y1 = f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa270_y2 & f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa271_y2;
  assign f_s_dadda_pg_rca32_fa286_y2 = f_s_dadda_pg_rca32_fa286_y0 ^ f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa272_y2;
  assign f_s_dadda_pg_rca32_fa286_y3 = f_s_dadda_pg_rca32_fa286_y0 & f_s_dadda_pg_rca32_fa286_f_s_dadda_pg_rca32_fa272_y2;
  assign f_s_dadda_pg_rca32_fa286_y4 = f_s_dadda_pg_rca32_fa286_y1 | f_s_dadda_pg_rca32_fa286_y3;
  assign f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa273_y2 = f_s_dadda_pg_rca32_fa273_y2;
  assign f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa274_y2 = f_s_dadda_pg_rca32_fa274_y2;
  assign f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa275_y2 = f_s_dadda_pg_rca32_fa275_y2;
  assign f_s_dadda_pg_rca32_fa287_y0 = f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa273_y2 ^ f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa274_y2;
  assign f_s_dadda_pg_rca32_fa287_y1 = f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa273_y2 & f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa274_y2;
  assign f_s_dadda_pg_rca32_fa287_y2 = f_s_dadda_pg_rca32_fa287_y0 ^ f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa275_y2;
  assign f_s_dadda_pg_rca32_fa287_y3 = f_s_dadda_pg_rca32_fa287_y0 & f_s_dadda_pg_rca32_fa287_f_s_dadda_pg_rca32_fa275_y2;
  assign f_s_dadda_pg_rca32_fa287_y4 = f_s_dadda_pg_rca32_fa287_y1 | f_s_dadda_pg_rca32_fa287_y3;
  assign f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa276_y2 = f_s_dadda_pg_rca32_fa276_y2;
  assign f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa277_y2 = f_s_dadda_pg_rca32_fa277_y2;
  assign f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa278_y2 = f_s_dadda_pg_rca32_fa278_y2;
  assign f_s_dadda_pg_rca32_fa288_y0 = f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa276_y2 ^ f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa277_y2;
  assign f_s_dadda_pg_rca32_fa288_y1 = f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa276_y2 & f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa277_y2;
  assign f_s_dadda_pg_rca32_fa288_y2 = f_s_dadda_pg_rca32_fa288_y0 ^ f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa278_y2;
  assign f_s_dadda_pg_rca32_fa288_y3 = f_s_dadda_pg_rca32_fa288_y0 & f_s_dadda_pg_rca32_fa288_f_s_dadda_pg_rca32_fa278_y2;
  assign f_s_dadda_pg_rca32_fa288_y4 = f_s_dadda_pg_rca32_fa288_y1 | f_s_dadda_pg_rca32_fa288_y3;
  assign f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa279_y2 = f_s_dadda_pg_rca32_fa279_y2;
  assign f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa280_y2 = f_s_dadda_pg_rca32_fa280_y2;
  assign f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa281_y2 = f_s_dadda_pg_rca32_fa281_y2;
  assign f_s_dadda_pg_rca32_fa289_y0 = f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa279_y2 ^ f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa280_y2;
  assign f_s_dadda_pg_rca32_fa289_y1 = f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa279_y2 & f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa280_y2;
  assign f_s_dadda_pg_rca32_fa289_y2 = f_s_dadda_pg_rca32_fa289_y0 ^ f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa281_y2;
  assign f_s_dadda_pg_rca32_fa289_y3 = f_s_dadda_pg_rca32_fa289_y0 & f_s_dadda_pg_rca32_fa289_f_s_dadda_pg_rca32_fa281_y2;
  assign f_s_dadda_pg_rca32_fa289_y4 = f_s_dadda_pg_rca32_fa289_y1 | f_s_dadda_pg_rca32_fa289_y3;
  assign f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa282_y2 = f_s_dadda_pg_rca32_fa282_y2;
  assign f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa283_y2 = f_s_dadda_pg_rca32_fa283_y2;
  assign f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa284_y2 = f_s_dadda_pg_rca32_fa284_y2;
  assign f_s_dadda_pg_rca32_fa290_y0 = f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa282_y2 ^ f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa283_y2;
  assign f_s_dadda_pg_rca32_fa290_y1 = f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa282_y2 & f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa283_y2;
  assign f_s_dadda_pg_rca32_fa290_y2 = f_s_dadda_pg_rca32_fa290_y0 ^ f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa284_y2;
  assign f_s_dadda_pg_rca32_fa290_y3 = f_s_dadda_pg_rca32_fa290_y0 & f_s_dadda_pg_rca32_fa290_f_s_dadda_pg_rca32_fa284_y2;
  assign f_s_dadda_pg_rca32_fa290_y4 = f_s_dadda_pg_rca32_fa290_y1 | f_s_dadda_pg_rca32_fa290_y3;
  assign f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa290_y4 = f_s_dadda_pg_rca32_fa290_y4;
  assign f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa289_y4 = f_s_dadda_pg_rca32_fa289_y4;
  assign f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa288_y4 = f_s_dadda_pg_rca32_fa288_y4;
  assign f_s_dadda_pg_rca32_fa291_y0 = f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa290_y4 ^ f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa289_y4;
  assign f_s_dadda_pg_rca32_fa291_y1 = f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa290_y4 & f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa289_y4;
  assign f_s_dadda_pg_rca32_fa291_y2 = f_s_dadda_pg_rca32_fa291_y0 ^ f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa288_y4;
  assign f_s_dadda_pg_rca32_fa291_y3 = f_s_dadda_pg_rca32_fa291_y0 & f_s_dadda_pg_rca32_fa291_f_s_dadda_pg_rca32_fa288_y4;
  assign f_s_dadda_pg_rca32_fa291_y4 = f_s_dadda_pg_rca32_fa291_y1 | f_s_dadda_pg_rca32_fa291_y3;
  assign f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa287_y4 = f_s_dadda_pg_rca32_fa287_y4;
  assign f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa286_y4 = f_s_dadda_pg_rca32_fa286_y4;
  assign f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa285_y4 = f_s_dadda_pg_rca32_fa285_y4;
  assign f_s_dadda_pg_rca32_fa292_y0 = f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa287_y4 ^ f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa286_y4;
  assign f_s_dadda_pg_rca32_fa292_y1 = f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa287_y4 & f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa286_y4;
  assign f_s_dadda_pg_rca32_fa292_y2 = f_s_dadda_pg_rca32_fa292_y0 ^ f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa285_y4;
  assign f_s_dadda_pg_rca32_fa292_y3 = f_s_dadda_pg_rca32_fa292_y0 & f_s_dadda_pg_rca32_fa292_f_s_dadda_pg_rca32_fa285_y4;
  assign f_s_dadda_pg_rca32_fa292_y4 = f_s_dadda_pg_rca32_fa292_y1 | f_s_dadda_pg_rca32_fa292_y3;
  assign f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa284_y4 = f_s_dadda_pg_rca32_fa284_y4;
  assign f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa283_y4 = f_s_dadda_pg_rca32_fa283_y4;
  assign f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa282_y4 = f_s_dadda_pg_rca32_fa282_y4;
  assign f_s_dadda_pg_rca32_fa293_y0 = f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa284_y4 ^ f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa283_y4;
  assign f_s_dadda_pg_rca32_fa293_y1 = f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa284_y4 & f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa283_y4;
  assign f_s_dadda_pg_rca32_fa293_y2 = f_s_dadda_pg_rca32_fa293_y0 ^ f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa282_y4;
  assign f_s_dadda_pg_rca32_fa293_y3 = f_s_dadda_pg_rca32_fa293_y0 & f_s_dadda_pg_rca32_fa293_f_s_dadda_pg_rca32_fa282_y4;
  assign f_s_dadda_pg_rca32_fa293_y4 = f_s_dadda_pg_rca32_fa293_y1 | f_s_dadda_pg_rca32_fa293_y3;
  assign f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa281_y4 = f_s_dadda_pg_rca32_fa281_y4;
  assign f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa280_y4 = f_s_dadda_pg_rca32_fa280_y4;
  assign f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa279_y4 = f_s_dadda_pg_rca32_fa279_y4;
  assign f_s_dadda_pg_rca32_fa294_y0 = f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa281_y4 ^ f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa280_y4;
  assign f_s_dadda_pg_rca32_fa294_y1 = f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa281_y4 & f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa280_y4;
  assign f_s_dadda_pg_rca32_fa294_y2 = f_s_dadda_pg_rca32_fa294_y0 ^ f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa279_y4;
  assign f_s_dadda_pg_rca32_fa294_y3 = f_s_dadda_pg_rca32_fa294_y0 & f_s_dadda_pg_rca32_fa294_f_s_dadda_pg_rca32_fa279_y4;
  assign f_s_dadda_pg_rca32_fa294_y4 = f_s_dadda_pg_rca32_fa294_y1 | f_s_dadda_pg_rca32_fa294_y3;
  assign f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa278_y4 = f_s_dadda_pg_rca32_fa278_y4;
  assign f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa277_y4 = f_s_dadda_pg_rca32_fa277_y4;
  assign f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa276_y4 = f_s_dadda_pg_rca32_fa276_y4;
  assign f_s_dadda_pg_rca32_fa295_y0 = f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa278_y4 ^ f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa277_y4;
  assign f_s_dadda_pg_rca32_fa295_y1 = f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa278_y4 & f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa277_y4;
  assign f_s_dadda_pg_rca32_fa295_y2 = f_s_dadda_pg_rca32_fa295_y0 ^ f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa276_y4;
  assign f_s_dadda_pg_rca32_fa295_y3 = f_s_dadda_pg_rca32_fa295_y0 & f_s_dadda_pg_rca32_fa295_f_s_dadda_pg_rca32_fa276_y4;
  assign f_s_dadda_pg_rca32_fa295_y4 = f_s_dadda_pg_rca32_fa295_y1 | f_s_dadda_pg_rca32_fa295_y3;
  assign f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa275_y4 = f_s_dadda_pg_rca32_fa275_y4;
  assign f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa274_y4 = f_s_dadda_pg_rca32_fa274_y4;
  assign f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa273_y4 = f_s_dadda_pg_rca32_fa273_y4;
  assign f_s_dadda_pg_rca32_fa296_y0 = f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa275_y4 ^ f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa274_y4;
  assign f_s_dadda_pg_rca32_fa296_y1 = f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa275_y4 & f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa274_y4;
  assign f_s_dadda_pg_rca32_fa296_y2 = f_s_dadda_pg_rca32_fa296_y0 ^ f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa273_y4;
  assign f_s_dadda_pg_rca32_fa296_y3 = f_s_dadda_pg_rca32_fa296_y0 & f_s_dadda_pg_rca32_fa296_f_s_dadda_pg_rca32_fa273_y4;
  assign f_s_dadda_pg_rca32_fa296_y4 = f_s_dadda_pg_rca32_fa296_y1 | f_s_dadda_pg_rca32_fa296_y3;
  assign f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa272_y4 = f_s_dadda_pg_rca32_fa272_y4;
  assign f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa271_y4 = f_s_dadda_pg_rca32_fa271_y4;
  assign f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa270_y4 = f_s_dadda_pg_rca32_fa270_y4;
  assign f_s_dadda_pg_rca32_fa297_y0 = f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa272_y4 ^ f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa271_y4;
  assign f_s_dadda_pg_rca32_fa297_y1 = f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa272_y4 & f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa271_y4;
  assign f_s_dadda_pg_rca32_fa297_y2 = f_s_dadda_pg_rca32_fa297_y0 ^ f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa270_y4;
  assign f_s_dadda_pg_rca32_fa297_y3 = f_s_dadda_pg_rca32_fa297_y0 & f_s_dadda_pg_rca32_fa297_f_s_dadda_pg_rca32_fa270_y4;
  assign f_s_dadda_pg_rca32_fa297_y4 = f_s_dadda_pg_rca32_fa297_y1 | f_s_dadda_pg_rca32_fa297_y3;
  assign f_s_dadda_pg_rca32_and_24_6_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_24_6_y0 = f_s_dadda_pg_rca32_and_24_6_a_24 & f_s_dadda_pg_rca32_and_24_6_b_6;
  assign f_s_dadda_pg_rca32_and_23_7_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_23_7_y0 = f_s_dadda_pg_rca32_and_23_7_a_23 & f_s_dadda_pg_rca32_and_23_7_b_7;
  assign f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_fa269_y4 = f_s_dadda_pg_rca32_fa269_y4;
  assign f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_and_24_6_y0 = f_s_dadda_pg_rca32_and_24_6_y0;
  assign f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_and_23_7_y0 = f_s_dadda_pg_rca32_and_23_7_y0;
  assign f_s_dadda_pg_rca32_fa298_y0 = f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_fa269_y4 ^ f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_and_24_6_y0;
  assign f_s_dadda_pg_rca32_fa298_y1 = f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_fa269_y4 & f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_and_24_6_y0;
  assign f_s_dadda_pg_rca32_fa298_y2 = f_s_dadda_pg_rca32_fa298_y0 ^ f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_and_23_7_y0;
  assign f_s_dadda_pg_rca32_fa298_y3 = f_s_dadda_pg_rca32_fa298_y0 & f_s_dadda_pg_rca32_fa298_f_s_dadda_pg_rca32_and_23_7_y0;
  assign f_s_dadda_pg_rca32_fa298_y4 = f_s_dadda_pg_rca32_fa298_y1 | f_s_dadda_pg_rca32_fa298_y3;
  assign f_s_dadda_pg_rca32_and_22_8_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_22_8_y0 = f_s_dadda_pg_rca32_and_22_8_a_22 & f_s_dadda_pg_rca32_and_22_8_b_8;
  assign f_s_dadda_pg_rca32_and_21_9_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_21_9_y0 = f_s_dadda_pg_rca32_and_21_9_a_21 & f_s_dadda_pg_rca32_and_21_9_b_9;
  assign f_s_dadda_pg_rca32_and_20_10_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_20_10_y0 = f_s_dadda_pg_rca32_and_20_10_a_20 & f_s_dadda_pg_rca32_and_20_10_b_10;
  assign f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_22_8_y0 = f_s_dadda_pg_rca32_and_22_8_y0;
  assign f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_21_9_y0 = f_s_dadda_pg_rca32_and_21_9_y0;
  assign f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_20_10_y0 = f_s_dadda_pg_rca32_and_20_10_y0;
  assign f_s_dadda_pg_rca32_fa299_y0 = f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_22_8_y0 ^ f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_21_9_y0;
  assign f_s_dadda_pg_rca32_fa299_y1 = f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_22_8_y0 & f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_21_9_y0;
  assign f_s_dadda_pg_rca32_fa299_y2 = f_s_dadda_pg_rca32_fa299_y0 ^ f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_20_10_y0;
  assign f_s_dadda_pg_rca32_fa299_y3 = f_s_dadda_pg_rca32_fa299_y0 & f_s_dadda_pg_rca32_fa299_f_s_dadda_pg_rca32_and_20_10_y0;
  assign f_s_dadda_pg_rca32_fa299_y4 = f_s_dadda_pg_rca32_fa299_y1 | f_s_dadda_pg_rca32_fa299_y3;
  assign f_s_dadda_pg_rca32_and_19_11_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_19_11_y0 = f_s_dadda_pg_rca32_and_19_11_a_19 & f_s_dadda_pg_rca32_and_19_11_b_11;
  assign f_s_dadda_pg_rca32_and_18_12_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_18_12_y0 = f_s_dadda_pg_rca32_and_18_12_a_18 & f_s_dadda_pg_rca32_and_18_12_b_12;
  assign f_s_dadda_pg_rca32_and_17_13_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_17_13_y0 = f_s_dadda_pg_rca32_and_17_13_a_17 & f_s_dadda_pg_rca32_and_17_13_b_13;
  assign f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_19_11_y0 = f_s_dadda_pg_rca32_and_19_11_y0;
  assign f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_18_12_y0 = f_s_dadda_pg_rca32_and_18_12_y0;
  assign f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_17_13_y0 = f_s_dadda_pg_rca32_and_17_13_y0;
  assign f_s_dadda_pg_rca32_fa300_y0 = f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_19_11_y0 ^ f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_18_12_y0;
  assign f_s_dadda_pg_rca32_fa300_y1 = f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_19_11_y0 & f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_18_12_y0;
  assign f_s_dadda_pg_rca32_fa300_y2 = f_s_dadda_pg_rca32_fa300_y0 ^ f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_17_13_y0;
  assign f_s_dadda_pg_rca32_fa300_y3 = f_s_dadda_pg_rca32_fa300_y0 & f_s_dadda_pg_rca32_fa300_f_s_dadda_pg_rca32_and_17_13_y0;
  assign f_s_dadda_pg_rca32_fa300_y4 = f_s_dadda_pg_rca32_fa300_y1 | f_s_dadda_pg_rca32_fa300_y3;
  assign f_s_dadda_pg_rca32_and_16_14_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_16_14_y0 = f_s_dadda_pg_rca32_and_16_14_a_16 & f_s_dadda_pg_rca32_and_16_14_b_14;
  assign f_s_dadda_pg_rca32_and_15_15_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_15_15_y0 = f_s_dadda_pg_rca32_and_15_15_a_15 & f_s_dadda_pg_rca32_and_15_15_b_15;
  assign f_s_dadda_pg_rca32_and_14_16_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_14_16_y0 = f_s_dadda_pg_rca32_and_14_16_a_14 & f_s_dadda_pg_rca32_and_14_16_b_16;
  assign f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_16_14_y0 = f_s_dadda_pg_rca32_and_16_14_y0;
  assign f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_15_15_y0 = f_s_dadda_pg_rca32_and_15_15_y0;
  assign f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_14_16_y0 = f_s_dadda_pg_rca32_and_14_16_y0;
  assign f_s_dadda_pg_rca32_fa301_y0 = f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_16_14_y0 ^ f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_15_15_y0;
  assign f_s_dadda_pg_rca32_fa301_y1 = f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_16_14_y0 & f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_15_15_y0;
  assign f_s_dadda_pg_rca32_fa301_y2 = f_s_dadda_pg_rca32_fa301_y0 ^ f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_14_16_y0;
  assign f_s_dadda_pg_rca32_fa301_y3 = f_s_dadda_pg_rca32_fa301_y0 & f_s_dadda_pg_rca32_fa301_f_s_dadda_pg_rca32_and_14_16_y0;
  assign f_s_dadda_pg_rca32_fa301_y4 = f_s_dadda_pg_rca32_fa301_y1 | f_s_dadda_pg_rca32_fa301_y3;
  assign f_s_dadda_pg_rca32_and_13_17_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_13_17_y0 = f_s_dadda_pg_rca32_and_13_17_a_13 & f_s_dadda_pg_rca32_and_13_17_b_17;
  assign f_s_dadda_pg_rca32_and_12_18_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_12_18_y0 = f_s_dadda_pg_rca32_and_12_18_a_12 & f_s_dadda_pg_rca32_and_12_18_b_18;
  assign f_s_dadda_pg_rca32_and_11_19_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_11_19_y0 = f_s_dadda_pg_rca32_and_11_19_a_11 & f_s_dadda_pg_rca32_and_11_19_b_19;
  assign f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_13_17_y0 = f_s_dadda_pg_rca32_and_13_17_y0;
  assign f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_12_18_y0 = f_s_dadda_pg_rca32_and_12_18_y0;
  assign f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_11_19_y0 = f_s_dadda_pg_rca32_and_11_19_y0;
  assign f_s_dadda_pg_rca32_fa302_y0 = f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_13_17_y0 ^ f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_12_18_y0;
  assign f_s_dadda_pg_rca32_fa302_y1 = f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_13_17_y0 & f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_12_18_y0;
  assign f_s_dadda_pg_rca32_fa302_y2 = f_s_dadda_pg_rca32_fa302_y0 ^ f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_11_19_y0;
  assign f_s_dadda_pg_rca32_fa302_y3 = f_s_dadda_pg_rca32_fa302_y0 & f_s_dadda_pg_rca32_fa302_f_s_dadda_pg_rca32_and_11_19_y0;
  assign f_s_dadda_pg_rca32_fa302_y4 = f_s_dadda_pg_rca32_fa302_y1 | f_s_dadda_pg_rca32_fa302_y3;
  assign f_s_dadda_pg_rca32_and_10_20_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_10_20_y0 = f_s_dadda_pg_rca32_and_10_20_a_10 & f_s_dadda_pg_rca32_and_10_20_b_20;
  assign f_s_dadda_pg_rca32_and_9_21_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_9_21_y0 = f_s_dadda_pg_rca32_and_9_21_a_9 & f_s_dadda_pg_rca32_and_9_21_b_21;
  assign f_s_dadda_pg_rca32_and_8_22_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_8_22_y0 = f_s_dadda_pg_rca32_and_8_22_a_8 & f_s_dadda_pg_rca32_and_8_22_b_22;
  assign f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_10_20_y0 = f_s_dadda_pg_rca32_and_10_20_y0;
  assign f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_9_21_y0 = f_s_dadda_pg_rca32_and_9_21_y0;
  assign f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_8_22_y0 = f_s_dadda_pg_rca32_and_8_22_y0;
  assign f_s_dadda_pg_rca32_fa303_y0 = f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_10_20_y0 ^ f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_9_21_y0;
  assign f_s_dadda_pg_rca32_fa303_y1 = f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_10_20_y0 & f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_9_21_y0;
  assign f_s_dadda_pg_rca32_fa303_y2 = f_s_dadda_pg_rca32_fa303_y0 ^ f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_8_22_y0;
  assign f_s_dadda_pg_rca32_fa303_y3 = f_s_dadda_pg_rca32_fa303_y0 & f_s_dadda_pg_rca32_fa303_f_s_dadda_pg_rca32_and_8_22_y0;
  assign f_s_dadda_pg_rca32_fa303_y4 = f_s_dadda_pg_rca32_fa303_y1 | f_s_dadda_pg_rca32_fa303_y3;
  assign f_s_dadda_pg_rca32_and_7_23_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_7_23_y0 = f_s_dadda_pg_rca32_and_7_23_a_7 & f_s_dadda_pg_rca32_and_7_23_b_23;
  assign f_s_dadda_pg_rca32_and_6_24_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_6_24_y0 = f_s_dadda_pg_rca32_and_6_24_a_6 & f_s_dadda_pg_rca32_and_6_24_b_24;
  assign f_s_dadda_pg_rca32_and_5_25_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_5_25_y0 = f_s_dadda_pg_rca32_and_5_25_a_5 & f_s_dadda_pg_rca32_and_5_25_b_25;
  assign f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_7_23_y0 = f_s_dadda_pg_rca32_and_7_23_y0;
  assign f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_6_24_y0 = f_s_dadda_pg_rca32_and_6_24_y0;
  assign f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_5_25_y0 = f_s_dadda_pg_rca32_and_5_25_y0;
  assign f_s_dadda_pg_rca32_fa304_y0 = f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_7_23_y0 ^ f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_6_24_y0;
  assign f_s_dadda_pg_rca32_fa304_y1 = f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_7_23_y0 & f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_6_24_y0;
  assign f_s_dadda_pg_rca32_fa304_y2 = f_s_dadda_pg_rca32_fa304_y0 ^ f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_5_25_y0;
  assign f_s_dadda_pg_rca32_fa304_y3 = f_s_dadda_pg_rca32_fa304_y0 & f_s_dadda_pg_rca32_fa304_f_s_dadda_pg_rca32_and_5_25_y0;
  assign f_s_dadda_pg_rca32_fa304_y4 = f_s_dadda_pg_rca32_fa304_y1 | f_s_dadda_pg_rca32_fa304_y3;
  assign f_s_dadda_pg_rca32_and_4_26_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_4_26_y0 = f_s_dadda_pg_rca32_and_4_26_a_4 & f_s_dadda_pg_rca32_and_4_26_b_26;
  assign f_s_dadda_pg_rca32_and_3_27_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_3_27_y0 = f_s_dadda_pg_rca32_and_3_27_a_3 & f_s_dadda_pg_rca32_and_3_27_b_27;
  assign f_s_dadda_pg_rca32_and_2_28_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_2_28_y0 = f_s_dadda_pg_rca32_and_2_28_a_2 & f_s_dadda_pg_rca32_and_2_28_b_28;
  assign f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_4_26_y0 = f_s_dadda_pg_rca32_and_4_26_y0;
  assign f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_3_27_y0 = f_s_dadda_pg_rca32_and_3_27_y0;
  assign f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_2_28_y0 = f_s_dadda_pg_rca32_and_2_28_y0;
  assign f_s_dadda_pg_rca32_fa305_y0 = f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_4_26_y0 ^ f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_3_27_y0;
  assign f_s_dadda_pg_rca32_fa305_y1 = f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_4_26_y0 & f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_3_27_y0;
  assign f_s_dadda_pg_rca32_fa305_y2 = f_s_dadda_pg_rca32_fa305_y0 ^ f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_2_28_y0;
  assign f_s_dadda_pg_rca32_fa305_y3 = f_s_dadda_pg_rca32_fa305_y0 & f_s_dadda_pg_rca32_fa305_f_s_dadda_pg_rca32_and_2_28_y0;
  assign f_s_dadda_pg_rca32_fa305_y4 = f_s_dadda_pg_rca32_fa305_y1 | f_s_dadda_pg_rca32_fa305_y3;
  assign f_s_dadda_pg_rca32_and_1_29_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_1_29_y0 = f_s_dadda_pg_rca32_and_1_29_a_1 & f_s_dadda_pg_rca32_and_1_29_b_29;
  assign f_s_dadda_pg_rca32_and_0_30_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_0_30_y0 = f_s_dadda_pg_rca32_and_0_30_a_0 & f_s_dadda_pg_rca32_and_0_30_b_30;
  assign f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_and_1_29_y0 = f_s_dadda_pg_rca32_and_1_29_y0;
  assign f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_and_0_30_y0 = f_s_dadda_pg_rca32_and_0_30_y0;
  assign f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_fa1_y2 = f_s_dadda_pg_rca32_fa1_y2;
  assign f_s_dadda_pg_rca32_fa306_y0 = f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_and_1_29_y0 ^ f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_and_0_30_y0;
  assign f_s_dadda_pg_rca32_fa306_y1 = f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_and_1_29_y0 & f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_and_0_30_y0;
  assign f_s_dadda_pg_rca32_fa306_y2 = f_s_dadda_pg_rca32_fa306_y0 ^ f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_fa1_y2;
  assign f_s_dadda_pg_rca32_fa306_y3 = f_s_dadda_pg_rca32_fa306_y0 & f_s_dadda_pg_rca32_fa306_f_s_dadda_pg_rca32_fa1_y2;
  assign f_s_dadda_pg_rca32_fa306_y4 = f_s_dadda_pg_rca32_fa306_y1 | f_s_dadda_pg_rca32_fa306_y3;
  assign f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_fa2_y2 = f_s_dadda_pg_rca32_fa2_y2;
  assign f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_ha2_y0 = f_s_dadda_pg_rca32_ha2_y0;
  assign f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_fa291_y2 = f_s_dadda_pg_rca32_fa291_y2;
  assign f_s_dadda_pg_rca32_fa307_y0 = f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_fa2_y2 ^ f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_ha2_y0;
  assign f_s_dadda_pg_rca32_fa307_y1 = f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_fa2_y2 & f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_ha2_y0;
  assign f_s_dadda_pg_rca32_fa307_y2 = f_s_dadda_pg_rca32_fa307_y0 ^ f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_fa291_y2;
  assign f_s_dadda_pg_rca32_fa307_y3 = f_s_dadda_pg_rca32_fa307_y0 & f_s_dadda_pg_rca32_fa307_f_s_dadda_pg_rca32_fa291_y2;
  assign f_s_dadda_pg_rca32_fa307_y4 = f_s_dadda_pg_rca32_fa307_y1 | f_s_dadda_pg_rca32_fa307_y3;
  assign f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa292_y2 = f_s_dadda_pg_rca32_fa292_y2;
  assign f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa293_y2 = f_s_dadda_pg_rca32_fa293_y2;
  assign f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa294_y2 = f_s_dadda_pg_rca32_fa294_y2;
  assign f_s_dadda_pg_rca32_fa308_y0 = f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa292_y2 ^ f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa293_y2;
  assign f_s_dadda_pg_rca32_fa308_y1 = f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa292_y2 & f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa293_y2;
  assign f_s_dadda_pg_rca32_fa308_y2 = f_s_dadda_pg_rca32_fa308_y0 ^ f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa294_y2;
  assign f_s_dadda_pg_rca32_fa308_y3 = f_s_dadda_pg_rca32_fa308_y0 & f_s_dadda_pg_rca32_fa308_f_s_dadda_pg_rca32_fa294_y2;
  assign f_s_dadda_pg_rca32_fa308_y4 = f_s_dadda_pg_rca32_fa308_y1 | f_s_dadda_pg_rca32_fa308_y3;
  assign f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa295_y2 = f_s_dadda_pg_rca32_fa295_y2;
  assign f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa296_y2 = f_s_dadda_pg_rca32_fa296_y2;
  assign f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa297_y2 = f_s_dadda_pg_rca32_fa297_y2;
  assign f_s_dadda_pg_rca32_fa309_y0 = f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa295_y2 ^ f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa296_y2;
  assign f_s_dadda_pg_rca32_fa309_y1 = f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa295_y2 & f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa296_y2;
  assign f_s_dadda_pg_rca32_fa309_y2 = f_s_dadda_pg_rca32_fa309_y0 ^ f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa297_y2;
  assign f_s_dadda_pg_rca32_fa309_y3 = f_s_dadda_pg_rca32_fa309_y0 & f_s_dadda_pg_rca32_fa309_f_s_dadda_pg_rca32_fa297_y2;
  assign f_s_dadda_pg_rca32_fa309_y4 = f_s_dadda_pg_rca32_fa309_y1 | f_s_dadda_pg_rca32_fa309_y3;
  assign f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa298_y2 = f_s_dadda_pg_rca32_fa298_y2;
  assign f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa299_y2 = f_s_dadda_pg_rca32_fa299_y2;
  assign f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa300_y2 = f_s_dadda_pg_rca32_fa300_y2;
  assign f_s_dadda_pg_rca32_fa310_y0 = f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa298_y2 ^ f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa299_y2;
  assign f_s_dadda_pg_rca32_fa310_y1 = f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa298_y2 & f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa299_y2;
  assign f_s_dadda_pg_rca32_fa310_y2 = f_s_dadda_pg_rca32_fa310_y0 ^ f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa300_y2;
  assign f_s_dadda_pg_rca32_fa310_y3 = f_s_dadda_pg_rca32_fa310_y0 & f_s_dadda_pg_rca32_fa310_f_s_dadda_pg_rca32_fa300_y2;
  assign f_s_dadda_pg_rca32_fa310_y4 = f_s_dadda_pg_rca32_fa310_y1 | f_s_dadda_pg_rca32_fa310_y3;
  assign f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa301_y2 = f_s_dadda_pg_rca32_fa301_y2;
  assign f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa302_y2 = f_s_dadda_pg_rca32_fa302_y2;
  assign f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa303_y2 = f_s_dadda_pg_rca32_fa303_y2;
  assign f_s_dadda_pg_rca32_fa311_y0 = f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa301_y2 ^ f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa302_y2;
  assign f_s_dadda_pg_rca32_fa311_y1 = f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa301_y2 & f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa302_y2;
  assign f_s_dadda_pg_rca32_fa311_y2 = f_s_dadda_pg_rca32_fa311_y0 ^ f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa303_y2;
  assign f_s_dadda_pg_rca32_fa311_y3 = f_s_dadda_pg_rca32_fa311_y0 & f_s_dadda_pg_rca32_fa311_f_s_dadda_pg_rca32_fa303_y2;
  assign f_s_dadda_pg_rca32_fa311_y4 = f_s_dadda_pg_rca32_fa311_y1 | f_s_dadda_pg_rca32_fa311_y3;
  assign f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa304_y2 = f_s_dadda_pg_rca32_fa304_y2;
  assign f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa305_y2 = f_s_dadda_pg_rca32_fa305_y2;
  assign f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa306_y2 = f_s_dadda_pg_rca32_fa306_y2;
  assign f_s_dadda_pg_rca32_fa312_y0 = f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa304_y2 ^ f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa305_y2;
  assign f_s_dadda_pg_rca32_fa312_y1 = f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa304_y2 & f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa305_y2;
  assign f_s_dadda_pg_rca32_fa312_y2 = f_s_dadda_pg_rca32_fa312_y0 ^ f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa306_y2;
  assign f_s_dadda_pg_rca32_fa312_y3 = f_s_dadda_pg_rca32_fa312_y0 & f_s_dadda_pg_rca32_fa312_f_s_dadda_pg_rca32_fa306_y2;
  assign f_s_dadda_pg_rca32_fa312_y4 = f_s_dadda_pg_rca32_fa312_y1 | f_s_dadda_pg_rca32_fa312_y3;
  assign f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa312_y4 = f_s_dadda_pg_rca32_fa312_y4;
  assign f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa311_y4 = f_s_dadda_pg_rca32_fa311_y4;
  assign f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa310_y4 = f_s_dadda_pg_rca32_fa310_y4;
  assign f_s_dadda_pg_rca32_fa313_y0 = f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa312_y4 ^ f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa311_y4;
  assign f_s_dadda_pg_rca32_fa313_y1 = f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa312_y4 & f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa311_y4;
  assign f_s_dadda_pg_rca32_fa313_y2 = f_s_dadda_pg_rca32_fa313_y0 ^ f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa310_y4;
  assign f_s_dadda_pg_rca32_fa313_y3 = f_s_dadda_pg_rca32_fa313_y0 & f_s_dadda_pg_rca32_fa313_f_s_dadda_pg_rca32_fa310_y4;
  assign f_s_dadda_pg_rca32_fa313_y4 = f_s_dadda_pg_rca32_fa313_y1 | f_s_dadda_pg_rca32_fa313_y3;
  assign f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa309_y4 = f_s_dadda_pg_rca32_fa309_y4;
  assign f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa308_y4 = f_s_dadda_pg_rca32_fa308_y4;
  assign f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa307_y4 = f_s_dadda_pg_rca32_fa307_y4;
  assign f_s_dadda_pg_rca32_fa314_y0 = f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa309_y4 ^ f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa308_y4;
  assign f_s_dadda_pg_rca32_fa314_y1 = f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa309_y4 & f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa308_y4;
  assign f_s_dadda_pg_rca32_fa314_y2 = f_s_dadda_pg_rca32_fa314_y0 ^ f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa307_y4;
  assign f_s_dadda_pg_rca32_fa314_y3 = f_s_dadda_pg_rca32_fa314_y0 & f_s_dadda_pg_rca32_fa314_f_s_dadda_pg_rca32_fa307_y4;
  assign f_s_dadda_pg_rca32_fa314_y4 = f_s_dadda_pg_rca32_fa314_y1 | f_s_dadda_pg_rca32_fa314_y3;
  assign f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa306_y4 = f_s_dadda_pg_rca32_fa306_y4;
  assign f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa305_y4 = f_s_dadda_pg_rca32_fa305_y4;
  assign f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa304_y4 = f_s_dadda_pg_rca32_fa304_y4;
  assign f_s_dadda_pg_rca32_fa315_y0 = f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa306_y4 ^ f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa305_y4;
  assign f_s_dadda_pg_rca32_fa315_y1 = f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa306_y4 & f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa305_y4;
  assign f_s_dadda_pg_rca32_fa315_y2 = f_s_dadda_pg_rca32_fa315_y0 ^ f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa304_y4;
  assign f_s_dadda_pg_rca32_fa315_y3 = f_s_dadda_pg_rca32_fa315_y0 & f_s_dadda_pg_rca32_fa315_f_s_dadda_pg_rca32_fa304_y4;
  assign f_s_dadda_pg_rca32_fa315_y4 = f_s_dadda_pg_rca32_fa315_y1 | f_s_dadda_pg_rca32_fa315_y3;
  assign f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa303_y4 = f_s_dadda_pg_rca32_fa303_y4;
  assign f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa302_y4 = f_s_dadda_pg_rca32_fa302_y4;
  assign f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa301_y4 = f_s_dadda_pg_rca32_fa301_y4;
  assign f_s_dadda_pg_rca32_fa316_y0 = f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa303_y4 ^ f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa302_y4;
  assign f_s_dadda_pg_rca32_fa316_y1 = f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa303_y4 & f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa302_y4;
  assign f_s_dadda_pg_rca32_fa316_y2 = f_s_dadda_pg_rca32_fa316_y0 ^ f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa301_y4;
  assign f_s_dadda_pg_rca32_fa316_y3 = f_s_dadda_pg_rca32_fa316_y0 & f_s_dadda_pg_rca32_fa316_f_s_dadda_pg_rca32_fa301_y4;
  assign f_s_dadda_pg_rca32_fa316_y4 = f_s_dadda_pg_rca32_fa316_y1 | f_s_dadda_pg_rca32_fa316_y3;
  assign f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa300_y4 = f_s_dadda_pg_rca32_fa300_y4;
  assign f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa299_y4 = f_s_dadda_pg_rca32_fa299_y4;
  assign f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa298_y4 = f_s_dadda_pg_rca32_fa298_y4;
  assign f_s_dadda_pg_rca32_fa317_y0 = f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa300_y4 ^ f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa299_y4;
  assign f_s_dadda_pg_rca32_fa317_y1 = f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa300_y4 & f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa299_y4;
  assign f_s_dadda_pg_rca32_fa317_y2 = f_s_dadda_pg_rca32_fa317_y0 ^ f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa298_y4;
  assign f_s_dadda_pg_rca32_fa317_y3 = f_s_dadda_pg_rca32_fa317_y0 & f_s_dadda_pg_rca32_fa317_f_s_dadda_pg_rca32_fa298_y4;
  assign f_s_dadda_pg_rca32_fa317_y4 = f_s_dadda_pg_rca32_fa317_y1 | f_s_dadda_pg_rca32_fa317_y3;
  assign f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa297_y4 = f_s_dadda_pg_rca32_fa297_y4;
  assign f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa296_y4 = f_s_dadda_pg_rca32_fa296_y4;
  assign f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa295_y4 = f_s_dadda_pg_rca32_fa295_y4;
  assign f_s_dadda_pg_rca32_fa318_y0 = f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa297_y4 ^ f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa296_y4;
  assign f_s_dadda_pg_rca32_fa318_y1 = f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa297_y4 & f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa296_y4;
  assign f_s_dadda_pg_rca32_fa318_y2 = f_s_dadda_pg_rca32_fa318_y0 ^ f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa295_y4;
  assign f_s_dadda_pg_rca32_fa318_y3 = f_s_dadda_pg_rca32_fa318_y0 & f_s_dadda_pg_rca32_fa318_f_s_dadda_pg_rca32_fa295_y4;
  assign f_s_dadda_pg_rca32_fa318_y4 = f_s_dadda_pg_rca32_fa318_y1 | f_s_dadda_pg_rca32_fa318_y3;
  assign f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa294_y4 = f_s_dadda_pg_rca32_fa294_y4;
  assign f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa293_y4 = f_s_dadda_pg_rca32_fa293_y4;
  assign f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa292_y4 = f_s_dadda_pg_rca32_fa292_y4;
  assign f_s_dadda_pg_rca32_fa319_y0 = f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa294_y4 ^ f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa293_y4;
  assign f_s_dadda_pg_rca32_fa319_y1 = f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa294_y4 & f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa293_y4;
  assign f_s_dadda_pg_rca32_fa319_y2 = f_s_dadda_pg_rca32_fa319_y0 ^ f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa292_y4;
  assign f_s_dadda_pg_rca32_fa319_y3 = f_s_dadda_pg_rca32_fa319_y0 & f_s_dadda_pg_rca32_fa319_f_s_dadda_pg_rca32_fa292_y4;
  assign f_s_dadda_pg_rca32_fa319_y4 = f_s_dadda_pg_rca32_fa319_y1 | f_s_dadda_pg_rca32_fa319_y3;
  assign f_s_dadda_pg_rca32_and_23_8_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_23_8_y0 = f_s_dadda_pg_rca32_and_23_8_a_23 & f_s_dadda_pg_rca32_and_23_8_b_8;
  assign f_s_dadda_pg_rca32_and_22_9_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_22_9_y0 = f_s_dadda_pg_rca32_and_22_9_a_22 & f_s_dadda_pg_rca32_and_22_9_b_9;
  assign f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_fa291_y4 = f_s_dadda_pg_rca32_fa291_y4;
  assign f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_and_23_8_y0 = f_s_dadda_pg_rca32_and_23_8_y0;
  assign f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_and_22_9_y0 = f_s_dadda_pg_rca32_and_22_9_y0;
  assign f_s_dadda_pg_rca32_fa320_y0 = f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_fa291_y4 ^ f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_and_23_8_y0;
  assign f_s_dadda_pg_rca32_fa320_y1 = f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_fa291_y4 & f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_and_23_8_y0;
  assign f_s_dadda_pg_rca32_fa320_y2 = f_s_dadda_pg_rca32_fa320_y0 ^ f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_and_22_9_y0;
  assign f_s_dadda_pg_rca32_fa320_y3 = f_s_dadda_pg_rca32_fa320_y0 & f_s_dadda_pg_rca32_fa320_f_s_dadda_pg_rca32_and_22_9_y0;
  assign f_s_dadda_pg_rca32_fa320_y4 = f_s_dadda_pg_rca32_fa320_y1 | f_s_dadda_pg_rca32_fa320_y3;
  assign f_s_dadda_pg_rca32_and_21_10_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_21_10_y0 = f_s_dadda_pg_rca32_and_21_10_a_21 & f_s_dadda_pg_rca32_and_21_10_b_10;
  assign f_s_dadda_pg_rca32_and_20_11_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_20_11_y0 = f_s_dadda_pg_rca32_and_20_11_a_20 & f_s_dadda_pg_rca32_and_20_11_b_11;
  assign f_s_dadda_pg_rca32_and_19_12_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_19_12_y0 = f_s_dadda_pg_rca32_and_19_12_a_19 & f_s_dadda_pg_rca32_and_19_12_b_12;
  assign f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_21_10_y0 = f_s_dadda_pg_rca32_and_21_10_y0;
  assign f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_20_11_y0 = f_s_dadda_pg_rca32_and_20_11_y0;
  assign f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_19_12_y0 = f_s_dadda_pg_rca32_and_19_12_y0;
  assign f_s_dadda_pg_rca32_fa321_y0 = f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_21_10_y0 ^ f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_20_11_y0;
  assign f_s_dadda_pg_rca32_fa321_y1 = f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_21_10_y0 & f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_20_11_y0;
  assign f_s_dadda_pg_rca32_fa321_y2 = f_s_dadda_pg_rca32_fa321_y0 ^ f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_19_12_y0;
  assign f_s_dadda_pg_rca32_fa321_y3 = f_s_dadda_pg_rca32_fa321_y0 & f_s_dadda_pg_rca32_fa321_f_s_dadda_pg_rca32_and_19_12_y0;
  assign f_s_dadda_pg_rca32_fa321_y4 = f_s_dadda_pg_rca32_fa321_y1 | f_s_dadda_pg_rca32_fa321_y3;
  assign f_s_dadda_pg_rca32_and_18_13_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_18_13_y0 = f_s_dadda_pg_rca32_and_18_13_a_18 & f_s_dadda_pg_rca32_and_18_13_b_13;
  assign f_s_dadda_pg_rca32_and_17_14_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_17_14_y0 = f_s_dadda_pg_rca32_and_17_14_a_17 & f_s_dadda_pg_rca32_and_17_14_b_14;
  assign f_s_dadda_pg_rca32_and_16_15_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_16_15_y0 = f_s_dadda_pg_rca32_and_16_15_a_16 & f_s_dadda_pg_rca32_and_16_15_b_15;
  assign f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_18_13_y0 = f_s_dadda_pg_rca32_and_18_13_y0;
  assign f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_17_14_y0 = f_s_dadda_pg_rca32_and_17_14_y0;
  assign f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_16_15_y0 = f_s_dadda_pg_rca32_and_16_15_y0;
  assign f_s_dadda_pg_rca32_fa322_y0 = f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_18_13_y0 ^ f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_17_14_y0;
  assign f_s_dadda_pg_rca32_fa322_y1 = f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_18_13_y0 & f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_17_14_y0;
  assign f_s_dadda_pg_rca32_fa322_y2 = f_s_dadda_pg_rca32_fa322_y0 ^ f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_16_15_y0;
  assign f_s_dadda_pg_rca32_fa322_y3 = f_s_dadda_pg_rca32_fa322_y0 & f_s_dadda_pg_rca32_fa322_f_s_dadda_pg_rca32_and_16_15_y0;
  assign f_s_dadda_pg_rca32_fa322_y4 = f_s_dadda_pg_rca32_fa322_y1 | f_s_dadda_pg_rca32_fa322_y3;
  assign f_s_dadda_pg_rca32_and_15_16_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_15_16_y0 = f_s_dadda_pg_rca32_and_15_16_a_15 & f_s_dadda_pg_rca32_and_15_16_b_16;
  assign f_s_dadda_pg_rca32_and_14_17_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_14_17_y0 = f_s_dadda_pg_rca32_and_14_17_a_14 & f_s_dadda_pg_rca32_and_14_17_b_17;
  assign f_s_dadda_pg_rca32_and_13_18_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_13_18_y0 = f_s_dadda_pg_rca32_and_13_18_a_13 & f_s_dadda_pg_rca32_and_13_18_b_18;
  assign f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_15_16_y0 = f_s_dadda_pg_rca32_and_15_16_y0;
  assign f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_14_17_y0 = f_s_dadda_pg_rca32_and_14_17_y0;
  assign f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_13_18_y0 = f_s_dadda_pg_rca32_and_13_18_y0;
  assign f_s_dadda_pg_rca32_fa323_y0 = f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_15_16_y0 ^ f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_14_17_y0;
  assign f_s_dadda_pg_rca32_fa323_y1 = f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_15_16_y0 & f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_14_17_y0;
  assign f_s_dadda_pg_rca32_fa323_y2 = f_s_dadda_pg_rca32_fa323_y0 ^ f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_13_18_y0;
  assign f_s_dadda_pg_rca32_fa323_y3 = f_s_dadda_pg_rca32_fa323_y0 & f_s_dadda_pg_rca32_fa323_f_s_dadda_pg_rca32_and_13_18_y0;
  assign f_s_dadda_pg_rca32_fa323_y4 = f_s_dadda_pg_rca32_fa323_y1 | f_s_dadda_pg_rca32_fa323_y3;
  assign f_s_dadda_pg_rca32_and_12_19_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_12_19_y0 = f_s_dadda_pg_rca32_and_12_19_a_12 & f_s_dadda_pg_rca32_and_12_19_b_19;
  assign f_s_dadda_pg_rca32_and_11_20_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_11_20_y0 = f_s_dadda_pg_rca32_and_11_20_a_11 & f_s_dadda_pg_rca32_and_11_20_b_20;
  assign f_s_dadda_pg_rca32_and_10_21_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_10_21_y0 = f_s_dadda_pg_rca32_and_10_21_a_10 & f_s_dadda_pg_rca32_and_10_21_b_21;
  assign f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_12_19_y0 = f_s_dadda_pg_rca32_and_12_19_y0;
  assign f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_11_20_y0 = f_s_dadda_pg_rca32_and_11_20_y0;
  assign f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_10_21_y0 = f_s_dadda_pg_rca32_and_10_21_y0;
  assign f_s_dadda_pg_rca32_fa324_y0 = f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_12_19_y0 ^ f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_11_20_y0;
  assign f_s_dadda_pg_rca32_fa324_y1 = f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_12_19_y0 & f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_11_20_y0;
  assign f_s_dadda_pg_rca32_fa324_y2 = f_s_dadda_pg_rca32_fa324_y0 ^ f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_10_21_y0;
  assign f_s_dadda_pg_rca32_fa324_y3 = f_s_dadda_pg_rca32_fa324_y0 & f_s_dadda_pg_rca32_fa324_f_s_dadda_pg_rca32_and_10_21_y0;
  assign f_s_dadda_pg_rca32_fa324_y4 = f_s_dadda_pg_rca32_fa324_y1 | f_s_dadda_pg_rca32_fa324_y3;
  assign f_s_dadda_pg_rca32_and_9_22_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_9_22_y0 = f_s_dadda_pg_rca32_and_9_22_a_9 & f_s_dadda_pg_rca32_and_9_22_b_22;
  assign f_s_dadda_pg_rca32_and_8_23_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_8_23_y0 = f_s_dadda_pg_rca32_and_8_23_a_8 & f_s_dadda_pg_rca32_and_8_23_b_23;
  assign f_s_dadda_pg_rca32_and_7_24_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_7_24_y0 = f_s_dadda_pg_rca32_and_7_24_a_7 & f_s_dadda_pg_rca32_and_7_24_b_24;
  assign f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_9_22_y0 = f_s_dadda_pg_rca32_and_9_22_y0;
  assign f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_8_23_y0 = f_s_dadda_pg_rca32_and_8_23_y0;
  assign f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_7_24_y0 = f_s_dadda_pg_rca32_and_7_24_y0;
  assign f_s_dadda_pg_rca32_fa325_y0 = f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_9_22_y0 ^ f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_8_23_y0;
  assign f_s_dadda_pg_rca32_fa325_y1 = f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_9_22_y0 & f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_8_23_y0;
  assign f_s_dadda_pg_rca32_fa325_y2 = f_s_dadda_pg_rca32_fa325_y0 ^ f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_7_24_y0;
  assign f_s_dadda_pg_rca32_fa325_y3 = f_s_dadda_pg_rca32_fa325_y0 & f_s_dadda_pg_rca32_fa325_f_s_dadda_pg_rca32_and_7_24_y0;
  assign f_s_dadda_pg_rca32_fa325_y4 = f_s_dadda_pg_rca32_fa325_y1 | f_s_dadda_pg_rca32_fa325_y3;
  assign f_s_dadda_pg_rca32_and_6_25_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_6_25_y0 = f_s_dadda_pg_rca32_and_6_25_a_6 & f_s_dadda_pg_rca32_and_6_25_b_25;
  assign f_s_dadda_pg_rca32_and_5_26_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_5_26_y0 = f_s_dadda_pg_rca32_and_5_26_a_5 & f_s_dadda_pg_rca32_and_5_26_b_26;
  assign f_s_dadda_pg_rca32_and_4_27_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_4_27_y0 = f_s_dadda_pg_rca32_and_4_27_a_4 & f_s_dadda_pg_rca32_and_4_27_b_27;
  assign f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_6_25_y0 = f_s_dadda_pg_rca32_and_6_25_y0;
  assign f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_5_26_y0 = f_s_dadda_pg_rca32_and_5_26_y0;
  assign f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_4_27_y0 = f_s_dadda_pg_rca32_and_4_27_y0;
  assign f_s_dadda_pg_rca32_fa326_y0 = f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_6_25_y0 ^ f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_5_26_y0;
  assign f_s_dadda_pg_rca32_fa326_y1 = f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_6_25_y0 & f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_5_26_y0;
  assign f_s_dadda_pg_rca32_fa326_y2 = f_s_dadda_pg_rca32_fa326_y0 ^ f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_4_27_y0;
  assign f_s_dadda_pg_rca32_fa326_y3 = f_s_dadda_pg_rca32_fa326_y0 & f_s_dadda_pg_rca32_fa326_f_s_dadda_pg_rca32_and_4_27_y0;
  assign f_s_dadda_pg_rca32_fa326_y4 = f_s_dadda_pg_rca32_fa326_y1 | f_s_dadda_pg_rca32_fa326_y3;
  assign f_s_dadda_pg_rca32_and_3_28_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_3_28_y0 = f_s_dadda_pg_rca32_and_3_28_a_3 & f_s_dadda_pg_rca32_and_3_28_b_28;
  assign f_s_dadda_pg_rca32_and_2_29_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_2_29_y0 = f_s_dadda_pg_rca32_and_2_29_a_2 & f_s_dadda_pg_rca32_and_2_29_b_29;
  assign f_s_dadda_pg_rca32_and_1_30_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_1_30_y0 = f_s_dadda_pg_rca32_and_1_30_a_1 & f_s_dadda_pg_rca32_and_1_30_b_30;
  assign f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_3_28_y0 = f_s_dadda_pg_rca32_and_3_28_y0;
  assign f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_2_29_y0 = f_s_dadda_pg_rca32_and_2_29_y0;
  assign f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_1_30_y0 = f_s_dadda_pg_rca32_and_1_30_y0;
  assign f_s_dadda_pg_rca32_fa327_y0 = f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_3_28_y0 ^ f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_2_29_y0;
  assign f_s_dadda_pg_rca32_fa327_y1 = f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_3_28_y0 & f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_2_29_y0;
  assign f_s_dadda_pg_rca32_fa327_y2 = f_s_dadda_pg_rca32_fa327_y0 ^ f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_1_30_y0;
  assign f_s_dadda_pg_rca32_fa327_y3 = f_s_dadda_pg_rca32_fa327_y0 & f_s_dadda_pg_rca32_fa327_f_s_dadda_pg_rca32_and_1_30_y0;
  assign f_s_dadda_pg_rca32_fa327_y4 = f_s_dadda_pg_rca32_fa327_y1 | f_s_dadda_pg_rca32_fa327_y3;
  assign f_s_dadda_pg_rca32_nand_0_31_a_0 = a_0;
  assign f_s_dadda_pg_rca32_nand_0_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_0_31_y0 = ~(f_s_dadda_pg_rca32_nand_0_31_a_0 & f_s_dadda_pg_rca32_nand_0_31_b_31);
  assign f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_nand_0_31_y0 = f_s_dadda_pg_rca32_nand_0_31_y0;
  assign f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_fa3_y2 = f_s_dadda_pg_rca32_fa3_y2;
  assign f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_fa4_y2 = f_s_dadda_pg_rca32_fa4_y2;
  assign f_s_dadda_pg_rca32_fa328_y0 = f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_nand_0_31_y0 ^ f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_fa3_y2;
  assign f_s_dadda_pg_rca32_fa328_y1 = f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_nand_0_31_y0 & f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_fa3_y2;
  assign f_s_dadda_pg_rca32_fa328_y2 = f_s_dadda_pg_rca32_fa328_y0 ^ f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_fa4_y2;
  assign f_s_dadda_pg_rca32_fa328_y3 = f_s_dadda_pg_rca32_fa328_y0 & f_s_dadda_pg_rca32_fa328_f_s_dadda_pg_rca32_fa4_y2;
  assign f_s_dadda_pg_rca32_fa328_y4 = f_s_dadda_pg_rca32_fa328_y1 | f_s_dadda_pg_rca32_fa328_y3;
  assign f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_fa5_y2 = f_s_dadda_pg_rca32_fa5_y2;
  assign f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_ha3_y0 = f_s_dadda_pg_rca32_ha3_y0;
  assign f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_fa313_y2 = f_s_dadda_pg_rca32_fa313_y2;
  assign f_s_dadda_pg_rca32_fa329_y0 = f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_fa5_y2 ^ f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_ha3_y0;
  assign f_s_dadda_pg_rca32_fa329_y1 = f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_fa5_y2 & f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_ha3_y0;
  assign f_s_dadda_pg_rca32_fa329_y2 = f_s_dadda_pg_rca32_fa329_y0 ^ f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_fa313_y2;
  assign f_s_dadda_pg_rca32_fa329_y3 = f_s_dadda_pg_rca32_fa329_y0 & f_s_dadda_pg_rca32_fa329_f_s_dadda_pg_rca32_fa313_y2;
  assign f_s_dadda_pg_rca32_fa329_y4 = f_s_dadda_pg_rca32_fa329_y1 | f_s_dadda_pg_rca32_fa329_y3;
  assign f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa314_y2 = f_s_dadda_pg_rca32_fa314_y2;
  assign f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa315_y2 = f_s_dadda_pg_rca32_fa315_y2;
  assign f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa316_y2 = f_s_dadda_pg_rca32_fa316_y2;
  assign f_s_dadda_pg_rca32_fa330_y0 = f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa314_y2 ^ f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa315_y2;
  assign f_s_dadda_pg_rca32_fa330_y1 = f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa314_y2 & f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa315_y2;
  assign f_s_dadda_pg_rca32_fa330_y2 = f_s_dadda_pg_rca32_fa330_y0 ^ f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa316_y2;
  assign f_s_dadda_pg_rca32_fa330_y3 = f_s_dadda_pg_rca32_fa330_y0 & f_s_dadda_pg_rca32_fa330_f_s_dadda_pg_rca32_fa316_y2;
  assign f_s_dadda_pg_rca32_fa330_y4 = f_s_dadda_pg_rca32_fa330_y1 | f_s_dadda_pg_rca32_fa330_y3;
  assign f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa317_y2 = f_s_dadda_pg_rca32_fa317_y2;
  assign f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa318_y2 = f_s_dadda_pg_rca32_fa318_y2;
  assign f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa319_y2 = f_s_dadda_pg_rca32_fa319_y2;
  assign f_s_dadda_pg_rca32_fa331_y0 = f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa317_y2 ^ f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa318_y2;
  assign f_s_dadda_pg_rca32_fa331_y1 = f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa317_y2 & f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa318_y2;
  assign f_s_dadda_pg_rca32_fa331_y2 = f_s_dadda_pg_rca32_fa331_y0 ^ f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa319_y2;
  assign f_s_dadda_pg_rca32_fa331_y3 = f_s_dadda_pg_rca32_fa331_y0 & f_s_dadda_pg_rca32_fa331_f_s_dadda_pg_rca32_fa319_y2;
  assign f_s_dadda_pg_rca32_fa331_y4 = f_s_dadda_pg_rca32_fa331_y1 | f_s_dadda_pg_rca32_fa331_y3;
  assign f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa320_y2 = f_s_dadda_pg_rca32_fa320_y2;
  assign f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa321_y2 = f_s_dadda_pg_rca32_fa321_y2;
  assign f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa322_y2 = f_s_dadda_pg_rca32_fa322_y2;
  assign f_s_dadda_pg_rca32_fa332_y0 = f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa320_y2 ^ f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa321_y2;
  assign f_s_dadda_pg_rca32_fa332_y1 = f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa320_y2 & f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa321_y2;
  assign f_s_dadda_pg_rca32_fa332_y2 = f_s_dadda_pg_rca32_fa332_y0 ^ f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa322_y2;
  assign f_s_dadda_pg_rca32_fa332_y3 = f_s_dadda_pg_rca32_fa332_y0 & f_s_dadda_pg_rca32_fa332_f_s_dadda_pg_rca32_fa322_y2;
  assign f_s_dadda_pg_rca32_fa332_y4 = f_s_dadda_pg_rca32_fa332_y1 | f_s_dadda_pg_rca32_fa332_y3;
  assign f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa323_y2 = f_s_dadda_pg_rca32_fa323_y2;
  assign f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa324_y2 = f_s_dadda_pg_rca32_fa324_y2;
  assign f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa325_y2 = f_s_dadda_pg_rca32_fa325_y2;
  assign f_s_dadda_pg_rca32_fa333_y0 = f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa323_y2 ^ f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa324_y2;
  assign f_s_dadda_pg_rca32_fa333_y1 = f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa323_y2 & f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa324_y2;
  assign f_s_dadda_pg_rca32_fa333_y2 = f_s_dadda_pg_rca32_fa333_y0 ^ f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa325_y2;
  assign f_s_dadda_pg_rca32_fa333_y3 = f_s_dadda_pg_rca32_fa333_y0 & f_s_dadda_pg_rca32_fa333_f_s_dadda_pg_rca32_fa325_y2;
  assign f_s_dadda_pg_rca32_fa333_y4 = f_s_dadda_pg_rca32_fa333_y1 | f_s_dadda_pg_rca32_fa333_y3;
  assign f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa326_y2 = f_s_dadda_pg_rca32_fa326_y2;
  assign f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa327_y2 = f_s_dadda_pg_rca32_fa327_y2;
  assign f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa328_y2 = f_s_dadda_pg_rca32_fa328_y2;
  assign f_s_dadda_pg_rca32_fa334_y0 = f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa326_y2 ^ f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa327_y2;
  assign f_s_dadda_pg_rca32_fa334_y1 = f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa326_y2 & f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa327_y2;
  assign f_s_dadda_pg_rca32_fa334_y2 = f_s_dadda_pg_rca32_fa334_y0 ^ f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa328_y2;
  assign f_s_dadda_pg_rca32_fa334_y3 = f_s_dadda_pg_rca32_fa334_y0 & f_s_dadda_pg_rca32_fa334_f_s_dadda_pg_rca32_fa328_y2;
  assign f_s_dadda_pg_rca32_fa334_y4 = f_s_dadda_pg_rca32_fa334_y1 | f_s_dadda_pg_rca32_fa334_y3;
  assign f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa334_y4 = f_s_dadda_pg_rca32_fa334_y4;
  assign f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa333_y4 = f_s_dadda_pg_rca32_fa333_y4;
  assign f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa332_y4 = f_s_dadda_pg_rca32_fa332_y4;
  assign f_s_dadda_pg_rca32_fa335_y0 = f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa334_y4 ^ f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa333_y4;
  assign f_s_dadda_pg_rca32_fa335_y1 = f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa334_y4 & f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa333_y4;
  assign f_s_dadda_pg_rca32_fa335_y2 = f_s_dadda_pg_rca32_fa335_y0 ^ f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa332_y4;
  assign f_s_dadda_pg_rca32_fa335_y3 = f_s_dadda_pg_rca32_fa335_y0 & f_s_dadda_pg_rca32_fa335_f_s_dadda_pg_rca32_fa332_y4;
  assign f_s_dadda_pg_rca32_fa335_y4 = f_s_dadda_pg_rca32_fa335_y1 | f_s_dadda_pg_rca32_fa335_y3;
  assign f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa331_y4 = f_s_dadda_pg_rca32_fa331_y4;
  assign f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa330_y4 = f_s_dadda_pg_rca32_fa330_y4;
  assign f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa329_y4 = f_s_dadda_pg_rca32_fa329_y4;
  assign f_s_dadda_pg_rca32_fa336_y0 = f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa331_y4 ^ f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa330_y4;
  assign f_s_dadda_pg_rca32_fa336_y1 = f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa331_y4 & f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa330_y4;
  assign f_s_dadda_pg_rca32_fa336_y2 = f_s_dadda_pg_rca32_fa336_y0 ^ f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa329_y4;
  assign f_s_dadda_pg_rca32_fa336_y3 = f_s_dadda_pg_rca32_fa336_y0 & f_s_dadda_pg_rca32_fa336_f_s_dadda_pg_rca32_fa329_y4;
  assign f_s_dadda_pg_rca32_fa336_y4 = f_s_dadda_pg_rca32_fa336_y1 | f_s_dadda_pg_rca32_fa336_y3;
  assign f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa328_y4 = f_s_dadda_pg_rca32_fa328_y4;
  assign f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa327_y4 = f_s_dadda_pg_rca32_fa327_y4;
  assign f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa326_y4 = f_s_dadda_pg_rca32_fa326_y4;
  assign f_s_dadda_pg_rca32_fa337_y0 = f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa328_y4 ^ f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa327_y4;
  assign f_s_dadda_pg_rca32_fa337_y1 = f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa328_y4 & f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa327_y4;
  assign f_s_dadda_pg_rca32_fa337_y2 = f_s_dadda_pg_rca32_fa337_y0 ^ f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa326_y4;
  assign f_s_dadda_pg_rca32_fa337_y3 = f_s_dadda_pg_rca32_fa337_y0 & f_s_dadda_pg_rca32_fa337_f_s_dadda_pg_rca32_fa326_y4;
  assign f_s_dadda_pg_rca32_fa337_y4 = f_s_dadda_pg_rca32_fa337_y1 | f_s_dadda_pg_rca32_fa337_y3;
  assign f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa325_y4 = f_s_dadda_pg_rca32_fa325_y4;
  assign f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa324_y4 = f_s_dadda_pg_rca32_fa324_y4;
  assign f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa323_y4 = f_s_dadda_pg_rca32_fa323_y4;
  assign f_s_dadda_pg_rca32_fa338_y0 = f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa325_y4 ^ f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa324_y4;
  assign f_s_dadda_pg_rca32_fa338_y1 = f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa325_y4 & f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa324_y4;
  assign f_s_dadda_pg_rca32_fa338_y2 = f_s_dadda_pg_rca32_fa338_y0 ^ f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa323_y4;
  assign f_s_dadda_pg_rca32_fa338_y3 = f_s_dadda_pg_rca32_fa338_y0 & f_s_dadda_pg_rca32_fa338_f_s_dadda_pg_rca32_fa323_y4;
  assign f_s_dadda_pg_rca32_fa338_y4 = f_s_dadda_pg_rca32_fa338_y1 | f_s_dadda_pg_rca32_fa338_y3;
  assign f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa322_y4 = f_s_dadda_pg_rca32_fa322_y4;
  assign f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa321_y4 = f_s_dadda_pg_rca32_fa321_y4;
  assign f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa320_y4 = f_s_dadda_pg_rca32_fa320_y4;
  assign f_s_dadda_pg_rca32_fa339_y0 = f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa322_y4 ^ f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa321_y4;
  assign f_s_dadda_pg_rca32_fa339_y1 = f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa322_y4 & f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa321_y4;
  assign f_s_dadda_pg_rca32_fa339_y2 = f_s_dadda_pg_rca32_fa339_y0 ^ f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa320_y4;
  assign f_s_dadda_pg_rca32_fa339_y3 = f_s_dadda_pg_rca32_fa339_y0 & f_s_dadda_pg_rca32_fa339_f_s_dadda_pg_rca32_fa320_y4;
  assign f_s_dadda_pg_rca32_fa339_y4 = f_s_dadda_pg_rca32_fa339_y1 | f_s_dadda_pg_rca32_fa339_y3;
  assign f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa319_y4 = f_s_dadda_pg_rca32_fa319_y4;
  assign f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa318_y4 = f_s_dadda_pg_rca32_fa318_y4;
  assign f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa317_y4 = f_s_dadda_pg_rca32_fa317_y4;
  assign f_s_dadda_pg_rca32_fa340_y0 = f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa319_y4 ^ f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa318_y4;
  assign f_s_dadda_pg_rca32_fa340_y1 = f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa319_y4 & f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa318_y4;
  assign f_s_dadda_pg_rca32_fa340_y2 = f_s_dadda_pg_rca32_fa340_y0 ^ f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa317_y4;
  assign f_s_dadda_pg_rca32_fa340_y3 = f_s_dadda_pg_rca32_fa340_y0 & f_s_dadda_pg_rca32_fa340_f_s_dadda_pg_rca32_fa317_y4;
  assign f_s_dadda_pg_rca32_fa340_y4 = f_s_dadda_pg_rca32_fa340_y1 | f_s_dadda_pg_rca32_fa340_y3;
  assign f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa316_y4 = f_s_dadda_pg_rca32_fa316_y4;
  assign f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa315_y4 = f_s_dadda_pg_rca32_fa315_y4;
  assign f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa314_y4 = f_s_dadda_pg_rca32_fa314_y4;
  assign f_s_dadda_pg_rca32_fa341_y0 = f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa316_y4 ^ f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa315_y4;
  assign f_s_dadda_pg_rca32_fa341_y1 = f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa316_y4 & f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa315_y4;
  assign f_s_dadda_pg_rca32_fa341_y2 = f_s_dadda_pg_rca32_fa341_y0 ^ f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa314_y4;
  assign f_s_dadda_pg_rca32_fa341_y3 = f_s_dadda_pg_rca32_fa341_y0 & f_s_dadda_pg_rca32_fa341_f_s_dadda_pg_rca32_fa314_y4;
  assign f_s_dadda_pg_rca32_fa341_y4 = f_s_dadda_pg_rca32_fa341_y1 | f_s_dadda_pg_rca32_fa341_y3;
  assign f_s_dadda_pg_rca32_and_24_8_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_24_8_y0 = f_s_dadda_pg_rca32_and_24_8_a_24 & f_s_dadda_pg_rca32_and_24_8_b_8;
  assign f_s_dadda_pg_rca32_and_23_9_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_23_9_y0 = f_s_dadda_pg_rca32_and_23_9_a_23 & f_s_dadda_pg_rca32_and_23_9_b_9;
  assign f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_fa313_y4 = f_s_dadda_pg_rca32_fa313_y4;
  assign f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_and_24_8_y0 = f_s_dadda_pg_rca32_and_24_8_y0;
  assign f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_and_23_9_y0 = f_s_dadda_pg_rca32_and_23_9_y0;
  assign f_s_dadda_pg_rca32_fa342_y0 = f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_fa313_y4 ^ f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_and_24_8_y0;
  assign f_s_dadda_pg_rca32_fa342_y1 = f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_fa313_y4 & f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_and_24_8_y0;
  assign f_s_dadda_pg_rca32_fa342_y2 = f_s_dadda_pg_rca32_fa342_y0 ^ f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_and_23_9_y0;
  assign f_s_dadda_pg_rca32_fa342_y3 = f_s_dadda_pg_rca32_fa342_y0 & f_s_dadda_pg_rca32_fa342_f_s_dadda_pg_rca32_and_23_9_y0;
  assign f_s_dadda_pg_rca32_fa342_y4 = f_s_dadda_pg_rca32_fa342_y1 | f_s_dadda_pg_rca32_fa342_y3;
  assign f_s_dadda_pg_rca32_and_22_10_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_22_10_y0 = f_s_dadda_pg_rca32_and_22_10_a_22 & f_s_dadda_pg_rca32_and_22_10_b_10;
  assign f_s_dadda_pg_rca32_and_21_11_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_21_11_y0 = f_s_dadda_pg_rca32_and_21_11_a_21 & f_s_dadda_pg_rca32_and_21_11_b_11;
  assign f_s_dadda_pg_rca32_and_20_12_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_20_12_y0 = f_s_dadda_pg_rca32_and_20_12_a_20 & f_s_dadda_pg_rca32_and_20_12_b_12;
  assign f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_22_10_y0 = f_s_dadda_pg_rca32_and_22_10_y0;
  assign f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_21_11_y0 = f_s_dadda_pg_rca32_and_21_11_y0;
  assign f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_20_12_y0 = f_s_dadda_pg_rca32_and_20_12_y0;
  assign f_s_dadda_pg_rca32_fa343_y0 = f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_22_10_y0 ^ f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_21_11_y0;
  assign f_s_dadda_pg_rca32_fa343_y1 = f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_22_10_y0 & f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_21_11_y0;
  assign f_s_dadda_pg_rca32_fa343_y2 = f_s_dadda_pg_rca32_fa343_y0 ^ f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_20_12_y0;
  assign f_s_dadda_pg_rca32_fa343_y3 = f_s_dadda_pg_rca32_fa343_y0 & f_s_dadda_pg_rca32_fa343_f_s_dadda_pg_rca32_and_20_12_y0;
  assign f_s_dadda_pg_rca32_fa343_y4 = f_s_dadda_pg_rca32_fa343_y1 | f_s_dadda_pg_rca32_fa343_y3;
  assign f_s_dadda_pg_rca32_and_19_13_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_19_13_y0 = f_s_dadda_pg_rca32_and_19_13_a_19 & f_s_dadda_pg_rca32_and_19_13_b_13;
  assign f_s_dadda_pg_rca32_and_18_14_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_18_14_y0 = f_s_dadda_pg_rca32_and_18_14_a_18 & f_s_dadda_pg_rca32_and_18_14_b_14;
  assign f_s_dadda_pg_rca32_and_17_15_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_17_15_y0 = f_s_dadda_pg_rca32_and_17_15_a_17 & f_s_dadda_pg_rca32_and_17_15_b_15;
  assign f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_19_13_y0 = f_s_dadda_pg_rca32_and_19_13_y0;
  assign f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_18_14_y0 = f_s_dadda_pg_rca32_and_18_14_y0;
  assign f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_17_15_y0 = f_s_dadda_pg_rca32_and_17_15_y0;
  assign f_s_dadda_pg_rca32_fa344_y0 = f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_19_13_y0 ^ f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_18_14_y0;
  assign f_s_dadda_pg_rca32_fa344_y1 = f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_19_13_y0 & f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_18_14_y0;
  assign f_s_dadda_pg_rca32_fa344_y2 = f_s_dadda_pg_rca32_fa344_y0 ^ f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_17_15_y0;
  assign f_s_dadda_pg_rca32_fa344_y3 = f_s_dadda_pg_rca32_fa344_y0 & f_s_dadda_pg_rca32_fa344_f_s_dadda_pg_rca32_and_17_15_y0;
  assign f_s_dadda_pg_rca32_fa344_y4 = f_s_dadda_pg_rca32_fa344_y1 | f_s_dadda_pg_rca32_fa344_y3;
  assign f_s_dadda_pg_rca32_and_16_16_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_16_16_y0 = f_s_dadda_pg_rca32_and_16_16_a_16 & f_s_dadda_pg_rca32_and_16_16_b_16;
  assign f_s_dadda_pg_rca32_and_15_17_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_15_17_y0 = f_s_dadda_pg_rca32_and_15_17_a_15 & f_s_dadda_pg_rca32_and_15_17_b_17;
  assign f_s_dadda_pg_rca32_and_14_18_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_14_18_y0 = f_s_dadda_pg_rca32_and_14_18_a_14 & f_s_dadda_pg_rca32_and_14_18_b_18;
  assign f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_16_16_y0 = f_s_dadda_pg_rca32_and_16_16_y0;
  assign f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_15_17_y0 = f_s_dadda_pg_rca32_and_15_17_y0;
  assign f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_14_18_y0 = f_s_dadda_pg_rca32_and_14_18_y0;
  assign f_s_dadda_pg_rca32_fa345_y0 = f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_16_16_y0 ^ f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_15_17_y0;
  assign f_s_dadda_pg_rca32_fa345_y1 = f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_16_16_y0 & f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_15_17_y0;
  assign f_s_dadda_pg_rca32_fa345_y2 = f_s_dadda_pg_rca32_fa345_y0 ^ f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_14_18_y0;
  assign f_s_dadda_pg_rca32_fa345_y3 = f_s_dadda_pg_rca32_fa345_y0 & f_s_dadda_pg_rca32_fa345_f_s_dadda_pg_rca32_and_14_18_y0;
  assign f_s_dadda_pg_rca32_fa345_y4 = f_s_dadda_pg_rca32_fa345_y1 | f_s_dadda_pg_rca32_fa345_y3;
  assign f_s_dadda_pg_rca32_and_13_19_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_13_19_y0 = f_s_dadda_pg_rca32_and_13_19_a_13 & f_s_dadda_pg_rca32_and_13_19_b_19;
  assign f_s_dadda_pg_rca32_and_12_20_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_12_20_y0 = f_s_dadda_pg_rca32_and_12_20_a_12 & f_s_dadda_pg_rca32_and_12_20_b_20;
  assign f_s_dadda_pg_rca32_and_11_21_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_11_21_y0 = f_s_dadda_pg_rca32_and_11_21_a_11 & f_s_dadda_pg_rca32_and_11_21_b_21;
  assign f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_13_19_y0 = f_s_dadda_pg_rca32_and_13_19_y0;
  assign f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_12_20_y0 = f_s_dadda_pg_rca32_and_12_20_y0;
  assign f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_11_21_y0 = f_s_dadda_pg_rca32_and_11_21_y0;
  assign f_s_dadda_pg_rca32_fa346_y0 = f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_13_19_y0 ^ f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_12_20_y0;
  assign f_s_dadda_pg_rca32_fa346_y1 = f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_13_19_y0 & f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_12_20_y0;
  assign f_s_dadda_pg_rca32_fa346_y2 = f_s_dadda_pg_rca32_fa346_y0 ^ f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_11_21_y0;
  assign f_s_dadda_pg_rca32_fa346_y3 = f_s_dadda_pg_rca32_fa346_y0 & f_s_dadda_pg_rca32_fa346_f_s_dadda_pg_rca32_and_11_21_y0;
  assign f_s_dadda_pg_rca32_fa346_y4 = f_s_dadda_pg_rca32_fa346_y1 | f_s_dadda_pg_rca32_fa346_y3;
  assign f_s_dadda_pg_rca32_and_10_22_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_10_22_y0 = f_s_dadda_pg_rca32_and_10_22_a_10 & f_s_dadda_pg_rca32_and_10_22_b_22;
  assign f_s_dadda_pg_rca32_and_9_23_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_9_23_y0 = f_s_dadda_pg_rca32_and_9_23_a_9 & f_s_dadda_pg_rca32_and_9_23_b_23;
  assign f_s_dadda_pg_rca32_and_8_24_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_8_24_y0 = f_s_dadda_pg_rca32_and_8_24_a_8 & f_s_dadda_pg_rca32_and_8_24_b_24;
  assign f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_10_22_y0 = f_s_dadda_pg_rca32_and_10_22_y0;
  assign f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_9_23_y0 = f_s_dadda_pg_rca32_and_9_23_y0;
  assign f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_8_24_y0 = f_s_dadda_pg_rca32_and_8_24_y0;
  assign f_s_dadda_pg_rca32_fa347_y0 = f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_10_22_y0 ^ f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_9_23_y0;
  assign f_s_dadda_pg_rca32_fa347_y1 = f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_10_22_y0 & f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_9_23_y0;
  assign f_s_dadda_pg_rca32_fa347_y2 = f_s_dadda_pg_rca32_fa347_y0 ^ f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_8_24_y0;
  assign f_s_dadda_pg_rca32_fa347_y3 = f_s_dadda_pg_rca32_fa347_y0 & f_s_dadda_pg_rca32_fa347_f_s_dadda_pg_rca32_and_8_24_y0;
  assign f_s_dadda_pg_rca32_fa347_y4 = f_s_dadda_pg_rca32_fa347_y1 | f_s_dadda_pg_rca32_fa347_y3;
  assign f_s_dadda_pg_rca32_and_7_25_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_7_25_y0 = f_s_dadda_pg_rca32_and_7_25_a_7 & f_s_dadda_pg_rca32_and_7_25_b_25;
  assign f_s_dadda_pg_rca32_and_6_26_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_6_26_y0 = f_s_dadda_pg_rca32_and_6_26_a_6 & f_s_dadda_pg_rca32_and_6_26_b_26;
  assign f_s_dadda_pg_rca32_and_5_27_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_5_27_y0 = f_s_dadda_pg_rca32_and_5_27_a_5 & f_s_dadda_pg_rca32_and_5_27_b_27;
  assign f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_7_25_y0 = f_s_dadda_pg_rca32_and_7_25_y0;
  assign f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_6_26_y0 = f_s_dadda_pg_rca32_and_6_26_y0;
  assign f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_5_27_y0 = f_s_dadda_pg_rca32_and_5_27_y0;
  assign f_s_dadda_pg_rca32_fa348_y0 = f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_7_25_y0 ^ f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_6_26_y0;
  assign f_s_dadda_pg_rca32_fa348_y1 = f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_7_25_y0 & f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_6_26_y0;
  assign f_s_dadda_pg_rca32_fa348_y2 = f_s_dadda_pg_rca32_fa348_y0 ^ f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_5_27_y0;
  assign f_s_dadda_pg_rca32_fa348_y3 = f_s_dadda_pg_rca32_fa348_y0 & f_s_dadda_pg_rca32_fa348_f_s_dadda_pg_rca32_and_5_27_y0;
  assign f_s_dadda_pg_rca32_fa348_y4 = f_s_dadda_pg_rca32_fa348_y1 | f_s_dadda_pg_rca32_fa348_y3;
  assign f_s_dadda_pg_rca32_and_4_28_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_4_28_y0 = f_s_dadda_pg_rca32_and_4_28_a_4 & f_s_dadda_pg_rca32_and_4_28_b_28;
  assign f_s_dadda_pg_rca32_and_3_29_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_3_29_y0 = f_s_dadda_pg_rca32_and_3_29_a_3 & f_s_dadda_pg_rca32_and_3_29_b_29;
  assign f_s_dadda_pg_rca32_and_2_30_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_2_30_y0 = f_s_dadda_pg_rca32_and_2_30_a_2 & f_s_dadda_pg_rca32_and_2_30_b_30;
  assign f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_4_28_y0 = f_s_dadda_pg_rca32_and_4_28_y0;
  assign f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_3_29_y0 = f_s_dadda_pg_rca32_and_3_29_y0;
  assign f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_2_30_y0 = f_s_dadda_pg_rca32_and_2_30_y0;
  assign f_s_dadda_pg_rca32_fa349_y0 = f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_4_28_y0 ^ f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_3_29_y0;
  assign f_s_dadda_pg_rca32_fa349_y1 = f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_4_28_y0 & f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_3_29_y0;
  assign f_s_dadda_pg_rca32_fa349_y2 = f_s_dadda_pg_rca32_fa349_y0 ^ f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_2_30_y0;
  assign f_s_dadda_pg_rca32_fa349_y3 = f_s_dadda_pg_rca32_fa349_y0 & f_s_dadda_pg_rca32_fa349_f_s_dadda_pg_rca32_and_2_30_y0;
  assign f_s_dadda_pg_rca32_fa349_y4 = f_s_dadda_pg_rca32_fa349_y1 | f_s_dadda_pg_rca32_fa349_y3;
  assign f_s_dadda_pg_rca32_nand_1_31_a_1 = a_1;
  assign f_s_dadda_pg_rca32_nand_1_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_1_31_y0 = ~(f_s_dadda_pg_rca32_nand_1_31_a_1 & f_s_dadda_pg_rca32_nand_1_31_b_31);
  assign f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_nand_1_31_y0 = f_s_dadda_pg_rca32_nand_1_31_y0;
  assign f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_fa6_y2 = f_s_dadda_pg_rca32_fa6_y2;
  assign f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_fa7_y2 = f_s_dadda_pg_rca32_fa7_y2;
  assign f_s_dadda_pg_rca32_fa350_y0 = f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_nand_1_31_y0 ^ f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_fa6_y2;
  assign f_s_dadda_pg_rca32_fa350_y1 = f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_nand_1_31_y0 & f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_fa6_y2;
  assign f_s_dadda_pg_rca32_fa350_y2 = f_s_dadda_pg_rca32_fa350_y0 ^ f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_fa7_y2;
  assign f_s_dadda_pg_rca32_fa350_y3 = f_s_dadda_pg_rca32_fa350_y0 & f_s_dadda_pg_rca32_fa350_f_s_dadda_pg_rca32_fa7_y2;
  assign f_s_dadda_pg_rca32_fa350_y4 = f_s_dadda_pg_rca32_fa350_y1 | f_s_dadda_pg_rca32_fa350_y3;
  assign f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa8_y2 = f_s_dadda_pg_rca32_fa8_y2;
  assign f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa9_y2 = f_s_dadda_pg_rca32_fa9_y2;
  assign f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa335_y2 = f_s_dadda_pg_rca32_fa335_y2;
  assign f_s_dadda_pg_rca32_fa351_y0 = f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa8_y2 ^ f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa9_y2;
  assign f_s_dadda_pg_rca32_fa351_y1 = f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa8_y2 & f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa9_y2;
  assign f_s_dadda_pg_rca32_fa351_y2 = f_s_dadda_pg_rca32_fa351_y0 ^ f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa335_y2;
  assign f_s_dadda_pg_rca32_fa351_y3 = f_s_dadda_pg_rca32_fa351_y0 & f_s_dadda_pg_rca32_fa351_f_s_dadda_pg_rca32_fa335_y2;
  assign f_s_dadda_pg_rca32_fa351_y4 = f_s_dadda_pg_rca32_fa351_y1 | f_s_dadda_pg_rca32_fa351_y3;
  assign f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa336_y2 = f_s_dadda_pg_rca32_fa336_y2;
  assign f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa337_y2 = f_s_dadda_pg_rca32_fa337_y2;
  assign f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa338_y2 = f_s_dadda_pg_rca32_fa338_y2;
  assign f_s_dadda_pg_rca32_fa352_y0 = f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa336_y2 ^ f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa337_y2;
  assign f_s_dadda_pg_rca32_fa352_y1 = f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa336_y2 & f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa337_y2;
  assign f_s_dadda_pg_rca32_fa352_y2 = f_s_dadda_pg_rca32_fa352_y0 ^ f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa338_y2;
  assign f_s_dadda_pg_rca32_fa352_y3 = f_s_dadda_pg_rca32_fa352_y0 & f_s_dadda_pg_rca32_fa352_f_s_dadda_pg_rca32_fa338_y2;
  assign f_s_dadda_pg_rca32_fa352_y4 = f_s_dadda_pg_rca32_fa352_y1 | f_s_dadda_pg_rca32_fa352_y3;
  assign f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa339_y2 = f_s_dadda_pg_rca32_fa339_y2;
  assign f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa340_y2 = f_s_dadda_pg_rca32_fa340_y2;
  assign f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa341_y2 = f_s_dadda_pg_rca32_fa341_y2;
  assign f_s_dadda_pg_rca32_fa353_y0 = f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa339_y2 ^ f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa340_y2;
  assign f_s_dadda_pg_rca32_fa353_y1 = f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa339_y2 & f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa340_y2;
  assign f_s_dadda_pg_rca32_fa353_y2 = f_s_dadda_pg_rca32_fa353_y0 ^ f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa341_y2;
  assign f_s_dadda_pg_rca32_fa353_y3 = f_s_dadda_pg_rca32_fa353_y0 & f_s_dadda_pg_rca32_fa353_f_s_dadda_pg_rca32_fa341_y2;
  assign f_s_dadda_pg_rca32_fa353_y4 = f_s_dadda_pg_rca32_fa353_y1 | f_s_dadda_pg_rca32_fa353_y3;
  assign f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa342_y2 = f_s_dadda_pg_rca32_fa342_y2;
  assign f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa343_y2 = f_s_dadda_pg_rca32_fa343_y2;
  assign f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa344_y2 = f_s_dadda_pg_rca32_fa344_y2;
  assign f_s_dadda_pg_rca32_fa354_y0 = f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa342_y2 ^ f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa343_y2;
  assign f_s_dadda_pg_rca32_fa354_y1 = f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa342_y2 & f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa343_y2;
  assign f_s_dadda_pg_rca32_fa354_y2 = f_s_dadda_pg_rca32_fa354_y0 ^ f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa344_y2;
  assign f_s_dadda_pg_rca32_fa354_y3 = f_s_dadda_pg_rca32_fa354_y0 & f_s_dadda_pg_rca32_fa354_f_s_dadda_pg_rca32_fa344_y2;
  assign f_s_dadda_pg_rca32_fa354_y4 = f_s_dadda_pg_rca32_fa354_y1 | f_s_dadda_pg_rca32_fa354_y3;
  assign f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa345_y2 = f_s_dadda_pg_rca32_fa345_y2;
  assign f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa346_y2 = f_s_dadda_pg_rca32_fa346_y2;
  assign f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa347_y2 = f_s_dadda_pg_rca32_fa347_y2;
  assign f_s_dadda_pg_rca32_fa355_y0 = f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa345_y2 ^ f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa346_y2;
  assign f_s_dadda_pg_rca32_fa355_y1 = f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa345_y2 & f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa346_y2;
  assign f_s_dadda_pg_rca32_fa355_y2 = f_s_dadda_pg_rca32_fa355_y0 ^ f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa347_y2;
  assign f_s_dadda_pg_rca32_fa355_y3 = f_s_dadda_pg_rca32_fa355_y0 & f_s_dadda_pg_rca32_fa355_f_s_dadda_pg_rca32_fa347_y2;
  assign f_s_dadda_pg_rca32_fa355_y4 = f_s_dadda_pg_rca32_fa355_y1 | f_s_dadda_pg_rca32_fa355_y3;
  assign f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa348_y2 = f_s_dadda_pg_rca32_fa348_y2;
  assign f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa349_y2 = f_s_dadda_pg_rca32_fa349_y2;
  assign f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa350_y2 = f_s_dadda_pg_rca32_fa350_y2;
  assign f_s_dadda_pg_rca32_fa356_y0 = f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa348_y2 ^ f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa349_y2;
  assign f_s_dadda_pg_rca32_fa356_y1 = f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa348_y2 & f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa349_y2;
  assign f_s_dadda_pg_rca32_fa356_y2 = f_s_dadda_pg_rca32_fa356_y0 ^ f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa350_y2;
  assign f_s_dadda_pg_rca32_fa356_y3 = f_s_dadda_pg_rca32_fa356_y0 & f_s_dadda_pg_rca32_fa356_f_s_dadda_pg_rca32_fa350_y2;
  assign f_s_dadda_pg_rca32_fa356_y4 = f_s_dadda_pg_rca32_fa356_y1 | f_s_dadda_pg_rca32_fa356_y3;
  assign f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa356_y4 = f_s_dadda_pg_rca32_fa356_y4;
  assign f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa355_y4 = f_s_dadda_pg_rca32_fa355_y4;
  assign f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa354_y4 = f_s_dadda_pg_rca32_fa354_y4;
  assign f_s_dadda_pg_rca32_fa357_y0 = f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa356_y4 ^ f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa355_y4;
  assign f_s_dadda_pg_rca32_fa357_y1 = f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa356_y4 & f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa355_y4;
  assign f_s_dadda_pg_rca32_fa357_y2 = f_s_dadda_pg_rca32_fa357_y0 ^ f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa354_y4;
  assign f_s_dadda_pg_rca32_fa357_y3 = f_s_dadda_pg_rca32_fa357_y0 & f_s_dadda_pg_rca32_fa357_f_s_dadda_pg_rca32_fa354_y4;
  assign f_s_dadda_pg_rca32_fa357_y4 = f_s_dadda_pg_rca32_fa357_y1 | f_s_dadda_pg_rca32_fa357_y3;
  assign f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa353_y4 = f_s_dadda_pg_rca32_fa353_y4;
  assign f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa352_y4 = f_s_dadda_pg_rca32_fa352_y4;
  assign f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa351_y4 = f_s_dadda_pg_rca32_fa351_y4;
  assign f_s_dadda_pg_rca32_fa358_y0 = f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa353_y4 ^ f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa352_y4;
  assign f_s_dadda_pg_rca32_fa358_y1 = f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa353_y4 & f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa352_y4;
  assign f_s_dadda_pg_rca32_fa358_y2 = f_s_dadda_pg_rca32_fa358_y0 ^ f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa351_y4;
  assign f_s_dadda_pg_rca32_fa358_y3 = f_s_dadda_pg_rca32_fa358_y0 & f_s_dadda_pg_rca32_fa358_f_s_dadda_pg_rca32_fa351_y4;
  assign f_s_dadda_pg_rca32_fa358_y4 = f_s_dadda_pg_rca32_fa358_y1 | f_s_dadda_pg_rca32_fa358_y3;
  assign f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa350_y4 = f_s_dadda_pg_rca32_fa350_y4;
  assign f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa349_y4 = f_s_dadda_pg_rca32_fa349_y4;
  assign f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa348_y4 = f_s_dadda_pg_rca32_fa348_y4;
  assign f_s_dadda_pg_rca32_fa359_y0 = f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa350_y4 ^ f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa349_y4;
  assign f_s_dadda_pg_rca32_fa359_y1 = f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa350_y4 & f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa349_y4;
  assign f_s_dadda_pg_rca32_fa359_y2 = f_s_dadda_pg_rca32_fa359_y0 ^ f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa348_y4;
  assign f_s_dadda_pg_rca32_fa359_y3 = f_s_dadda_pg_rca32_fa359_y0 & f_s_dadda_pg_rca32_fa359_f_s_dadda_pg_rca32_fa348_y4;
  assign f_s_dadda_pg_rca32_fa359_y4 = f_s_dadda_pg_rca32_fa359_y1 | f_s_dadda_pg_rca32_fa359_y3;
  assign f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa347_y4 = f_s_dadda_pg_rca32_fa347_y4;
  assign f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa346_y4 = f_s_dadda_pg_rca32_fa346_y4;
  assign f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa345_y4 = f_s_dadda_pg_rca32_fa345_y4;
  assign f_s_dadda_pg_rca32_fa360_y0 = f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa347_y4 ^ f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa346_y4;
  assign f_s_dadda_pg_rca32_fa360_y1 = f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa347_y4 & f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa346_y4;
  assign f_s_dadda_pg_rca32_fa360_y2 = f_s_dadda_pg_rca32_fa360_y0 ^ f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa345_y4;
  assign f_s_dadda_pg_rca32_fa360_y3 = f_s_dadda_pg_rca32_fa360_y0 & f_s_dadda_pg_rca32_fa360_f_s_dadda_pg_rca32_fa345_y4;
  assign f_s_dadda_pg_rca32_fa360_y4 = f_s_dadda_pg_rca32_fa360_y1 | f_s_dadda_pg_rca32_fa360_y3;
  assign f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa344_y4 = f_s_dadda_pg_rca32_fa344_y4;
  assign f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa343_y4 = f_s_dadda_pg_rca32_fa343_y4;
  assign f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa342_y4 = f_s_dadda_pg_rca32_fa342_y4;
  assign f_s_dadda_pg_rca32_fa361_y0 = f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa344_y4 ^ f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa343_y4;
  assign f_s_dadda_pg_rca32_fa361_y1 = f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa344_y4 & f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa343_y4;
  assign f_s_dadda_pg_rca32_fa361_y2 = f_s_dadda_pg_rca32_fa361_y0 ^ f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa342_y4;
  assign f_s_dadda_pg_rca32_fa361_y3 = f_s_dadda_pg_rca32_fa361_y0 & f_s_dadda_pg_rca32_fa361_f_s_dadda_pg_rca32_fa342_y4;
  assign f_s_dadda_pg_rca32_fa361_y4 = f_s_dadda_pg_rca32_fa361_y1 | f_s_dadda_pg_rca32_fa361_y3;
  assign f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa341_y4 = f_s_dadda_pg_rca32_fa341_y4;
  assign f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa340_y4 = f_s_dadda_pg_rca32_fa340_y4;
  assign f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa339_y4 = f_s_dadda_pg_rca32_fa339_y4;
  assign f_s_dadda_pg_rca32_fa362_y0 = f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa341_y4 ^ f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa340_y4;
  assign f_s_dadda_pg_rca32_fa362_y1 = f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa341_y4 & f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa340_y4;
  assign f_s_dadda_pg_rca32_fa362_y2 = f_s_dadda_pg_rca32_fa362_y0 ^ f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa339_y4;
  assign f_s_dadda_pg_rca32_fa362_y3 = f_s_dadda_pg_rca32_fa362_y0 & f_s_dadda_pg_rca32_fa362_f_s_dadda_pg_rca32_fa339_y4;
  assign f_s_dadda_pg_rca32_fa362_y4 = f_s_dadda_pg_rca32_fa362_y1 | f_s_dadda_pg_rca32_fa362_y3;
  assign f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa338_y4 = f_s_dadda_pg_rca32_fa338_y4;
  assign f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa337_y4 = f_s_dadda_pg_rca32_fa337_y4;
  assign f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa336_y4 = f_s_dadda_pg_rca32_fa336_y4;
  assign f_s_dadda_pg_rca32_fa363_y0 = f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa338_y4 ^ f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa337_y4;
  assign f_s_dadda_pg_rca32_fa363_y1 = f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa338_y4 & f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa337_y4;
  assign f_s_dadda_pg_rca32_fa363_y2 = f_s_dadda_pg_rca32_fa363_y0 ^ f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa336_y4;
  assign f_s_dadda_pg_rca32_fa363_y3 = f_s_dadda_pg_rca32_fa363_y0 & f_s_dadda_pg_rca32_fa363_f_s_dadda_pg_rca32_fa336_y4;
  assign f_s_dadda_pg_rca32_fa363_y4 = f_s_dadda_pg_rca32_fa363_y1 | f_s_dadda_pg_rca32_fa363_y3;
  assign f_s_dadda_pg_rca32_and_26_7_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_26_7_y0 = f_s_dadda_pg_rca32_and_26_7_a_26 & f_s_dadda_pg_rca32_and_26_7_b_7;
  assign f_s_dadda_pg_rca32_and_25_8_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_25_8_y0 = f_s_dadda_pg_rca32_and_25_8_a_25 & f_s_dadda_pg_rca32_and_25_8_b_8;
  assign f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_fa335_y4 = f_s_dadda_pg_rca32_fa335_y4;
  assign f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_and_26_7_y0 = f_s_dadda_pg_rca32_and_26_7_y0;
  assign f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_and_25_8_y0 = f_s_dadda_pg_rca32_and_25_8_y0;
  assign f_s_dadda_pg_rca32_fa364_y0 = f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_fa335_y4 ^ f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_and_26_7_y0;
  assign f_s_dadda_pg_rca32_fa364_y1 = f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_fa335_y4 & f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_and_26_7_y0;
  assign f_s_dadda_pg_rca32_fa364_y2 = f_s_dadda_pg_rca32_fa364_y0 ^ f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_and_25_8_y0;
  assign f_s_dadda_pg_rca32_fa364_y3 = f_s_dadda_pg_rca32_fa364_y0 & f_s_dadda_pg_rca32_fa364_f_s_dadda_pg_rca32_and_25_8_y0;
  assign f_s_dadda_pg_rca32_fa364_y4 = f_s_dadda_pg_rca32_fa364_y1 | f_s_dadda_pg_rca32_fa364_y3;
  assign f_s_dadda_pg_rca32_and_24_9_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_24_9_y0 = f_s_dadda_pg_rca32_and_24_9_a_24 & f_s_dadda_pg_rca32_and_24_9_b_9;
  assign f_s_dadda_pg_rca32_and_23_10_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_23_10_y0 = f_s_dadda_pg_rca32_and_23_10_a_23 & f_s_dadda_pg_rca32_and_23_10_b_10;
  assign f_s_dadda_pg_rca32_and_22_11_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_22_11_y0 = f_s_dadda_pg_rca32_and_22_11_a_22 & f_s_dadda_pg_rca32_and_22_11_b_11;
  assign f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_24_9_y0 = f_s_dadda_pg_rca32_and_24_9_y0;
  assign f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_23_10_y0 = f_s_dadda_pg_rca32_and_23_10_y0;
  assign f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_22_11_y0 = f_s_dadda_pg_rca32_and_22_11_y0;
  assign f_s_dadda_pg_rca32_fa365_y0 = f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_24_9_y0 ^ f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_23_10_y0;
  assign f_s_dadda_pg_rca32_fa365_y1 = f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_24_9_y0 & f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_23_10_y0;
  assign f_s_dadda_pg_rca32_fa365_y2 = f_s_dadda_pg_rca32_fa365_y0 ^ f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_22_11_y0;
  assign f_s_dadda_pg_rca32_fa365_y3 = f_s_dadda_pg_rca32_fa365_y0 & f_s_dadda_pg_rca32_fa365_f_s_dadda_pg_rca32_and_22_11_y0;
  assign f_s_dadda_pg_rca32_fa365_y4 = f_s_dadda_pg_rca32_fa365_y1 | f_s_dadda_pg_rca32_fa365_y3;
  assign f_s_dadda_pg_rca32_and_21_12_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_21_12_y0 = f_s_dadda_pg_rca32_and_21_12_a_21 & f_s_dadda_pg_rca32_and_21_12_b_12;
  assign f_s_dadda_pg_rca32_and_20_13_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_20_13_y0 = f_s_dadda_pg_rca32_and_20_13_a_20 & f_s_dadda_pg_rca32_and_20_13_b_13;
  assign f_s_dadda_pg_rca32_and_19_14_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_19_14_y0 = f_s_dadda_pg_rca32_and_19_14_a_19 & f_s_dadda_pg_rca32_and_19_14_b_14;
  assign f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_21_12_y0 = f_s_dadda_pg_rca32_and_21_12_y0;
  assign f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_20_13_y0 = f_s_dadda_pg_rca32_and_20_13_y0;
  assign f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_19_14_y0 = f_s_dadda_pg_rca32_and_19_14_y0;
  assign f_s_dadda_pg_rca32_fa366_y0 = f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_21_12_y0 ^ f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_20_13_y0;
  assign f_s_dadda_pg_rca32_fa366_y1 = f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_21_12_y0 & f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_20_13_y0;
  assign f_s_dadda_pg_rca32_fa366_y2 = f_s_dadda_pg_rca32_fa366_y0 ^ f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_19_14_y0;
  assign f_s_dadda_pg_rca32_fa366_y3 = f_s_dadda_pg_rca32_fa366_y0 & f_s_dadda_pg_rca32_fa366_f_s_dadda_pg_rca32_and_19_14_y0;
  assign f_s_dadda_pg_rca32_fa366_y4 = f_s_dadda_pg_rca32_fa366_y1 | f_s_dadda_pg_rca32_fa366_y3;
  assign f_s_dadda_pg_rca32_and_18_15_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_18_15_y0 = f_s_dadda_pg_rca32_and_18_15_a_18 & f_s_dadda_pg_rca32_and_18_15_b_15;
  assign f_s_dadda_pg_rca32_and_17_16_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_17_16_y0 = f_s_dadda_pg_rca32_and_17_16_a_17 & f_s_dadda_pg_rca32_and_17_16_b_16;
  assign f_s_dadda_pg_rca32_and_16_17_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_16_17_y0 = f_s_dadda_pg_rca32_and_16_17_a_16 & f_s_dadda_pg_rca32_and_16_17_b_17;
  assign f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_18_15_y0 = f_s_dadda_pg_rca32_and_18_15_y0;
  assign f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_17_16_y0 = f_s_dadda_pg_rca32_and_17_16_y0;
  assign f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_16_17_y0 = f_s_dadda_pg_rca32_and_16_17_y0;
  assign f_s_dadda_pg_rca32_fa367_y0 = f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_18_15_y0 ^ f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_17_16_y0;
  assign f_s_dadda_pg_rca32_fa367_y1 = f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_18_15_y0 & f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_17_16_y0;
  assign f_s_dadda_pg_rca32_fa367_y2 = f_s_dadda_pg_rca32_fa367_y0 ^ f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_16_17_y0;
  assign f_s_dadda_pg_rca32_fa367_y3 = f_s_dadda_pg_rca32_fa367_y0 & f_s_dadda_pg_rca32_fa367_f_s_dadda_pg_rca32_and_16_17_y0;
  assign f_s_dadda_pg_rca32_fa367_y4 = f_s_dadda_pg_rca32_fa367_y1 | f_s_dadda_pg_rca32_fa367_y3;
  assign f_s_dadda_pg_rca32_and_15_18_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_15_18_y0 = f_s_dadda_pg_rca32_and_15_18_a_15 & f_s_dadda_pg_rca32_and_15_18_b_18;
  assign f_s_dadda_pg_rca32_and_14_19_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_14_19_y0 = f_s_dadda_pg_rca32_and_14_19_a_14 & f_s_dadda_pg_rca32_and_14_19_b_19;
  assign f_s_dadda_pg_rca32_and_13_20_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_13_20_y0 = f_s_dadda_pg_rca32_and_13_20_a_13 & f_s_dadda_pg_rca32_and_13_20_b_20;
  assign f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_15_18_y0 = f_s_dadda_pg_rca32_and_15_18_y0;
  assign f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_14_19_y0 = f_s_dadda_pg_rca32_and_14_19_y0;
  assign f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_13_20_y0 = f_s_dadda_pg_rca32_and_13_20_y0;
  assign f_s_dadda_pg_rca32_fa368_y0 = f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_15_18_y0 ^ f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_14_19_y0;
  assign f_s_dadda_pg_rca32_fa368_y1 = f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_15_18_y0 & f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_14_19_y0;
  assign f_s_dadda_pg_rca32_fa368_y2 = f_s_dadda_pg_rca32_fa368_y0 ^ f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_13_20_y0;
  assign f_s_dadda_pg_rca32_fa368_y3 = f_s_dadda_pg_rca32_fa368_y0 & f_s_dadda_pg_rca32_fa368_f_s_dadda_pg_rca32_and_13_20_y0;
  assign f_s_dadda_pg_rca32_fa368_y4 = f_s_dadda_pg_rca32_fa368_y1 | f_s_dadda_pg_rca32_fa368_y3;
  assign f_s_dadda_pg_rca32_and_12_21_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_12_21_y0 = f_s_dadda_pg_rca32_and_12_21_a_12 & f_s_dadda_pg_rca32_and_12_21_b_21;
  assign f_s_dadda_pg_rca32_and_11_22_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_11_22_y0 = f_s_dadda_pg_rca32_and_11_22_a_11 & f_s_dadda_pg_rca32_and_11_22_b_22;
  assign f_s_dadda_pg_rca32_and_10_23_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_10_23_y0 = f_s_dadda_pg_rca32_and_10_23_a_10 & f_s_dadda_pg_rca32_and_10_23_b_23;
  assign f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_12_21_y0 = f_s_dadda_pg_rca32_and_12_21_y0;
  assign f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_11_22_y0 = f_s_dadda_pg_rca32_and_11_22_y0;
  assign f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_10_23_y0 = f_s_dadda_pg_rca32_and_10_23_y0;
  assign f_s_dadda_pg_rca32_fa369_y0 = f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_12_21_y0 ^ f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_11_22_y0;
  assign f_s_dadda_pg_rca32_fa369_y1 = f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_12_21_y0 & f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_11_22_y0;
  assign f_s_dadda_pg_rca32_fa369_y2 = f_s_dadda_pg_rca32_fa369_y0 ^ f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_10_23_y0;
  assign f_s_dadda_pg_rca32_fa369_y3 = f_s_dadda_pg_rca32_fa369_y0 & f_s_dadda_pg_rca32_fa369_f_s_dadda_pg_rca32_and_10_23_y0;
  assign f_s_dadda_pg_rca32_fa369_y4 = f_s_dadda_pg_rca32_fa369_y1 | f_s_dadda_pg_rca32_fa369_y3;
  assign f_s_dadda_pg_rca32_and_9_24_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_9_24_y0 = f_s_dadda_pg_rca32_and_9_24_a_9 & f_s_dadda_pg_rca32_and_9_24_b_24;
  assign f_s_dadda_pg_rca32_and_8_25_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_8_25_y0 = f_s_dadda_pg_rca32_and_8_25_a_8 & f_s_dadda_pg_rca32_and_8_25_b_25;
  assign f_s_dadda_pg_rca32_and_7_26_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_7_26_y0 = f_s_dadda_pg_rca32_and_7_26_a_7 & f_s_dadda_pg_rca32_and_7_26_b_26;
  assign f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_9_24_y0 = f_s_dadda_pg_rca32_and_9_24_y0;
  assign f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_8_25_y0 = f_s_dadda_pg_rca32_and_8_25_y0;
  assign f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_7_26_y0 = f_s_dadda_pg_rca32_and_7_26_y0;
  assign f_s_dadda_pg_rca32_fa370_y0 = f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_9_24_y0 ^ f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_8_25_y0;
  assign f_s_dadda_pg_rca32_fa370_y1 = f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_9_24_y0 & f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_8_25_y0;
  assign f_s_dadda_pg_rca32_fa370_y2 = f_s_dadda_pg_rca32_fa370_y0 ^ f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_7_26_y0;
  assign f_s_dadda_pg_rca32_fa370_y3 = f_s_dadda_pg_rca32_fa370_y0 & f_s_dadda_pg_rca32_fa370_f_s_dadda_pg_rca32_and_7_26_y0;
  assign f_s_dadda_pg_rca32_fa370_y4 = f_s_dadda_pg_rca32_fa370_y1 | f_s_dadda_pg_rca32_fa370_y3;
  assign f_s_dadda_pg_rca32_and_6_27_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_6_27_y0 = f_s_dadda_pg_rca32_and_6_27_a_6 & f_s_dadda_pg_rca32_and_6_27_b_27;
  assign f_s_dadda_pg_rca32_and_5_28_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_5_28_y0 = f_s_dadda_pg_rca32_and_5_28_a_5 & f_s_dadda_pg_rca32_and_5_28_b_28;
  assign f_s_dadda_pg_rca32_and_4_29_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_4_29_y0 = f_s_dadda_pg_rca32_and_4_29_a_4 & f_s_dadda_pg_rca32_and_4_29_b_29;
  assign f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_6_27_y0 = f_s_dadda_pg_rca32_and_6_27_y0;
  assign f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_5_28_y0 = f_s_dadda_pg_rca32_and_5_28_y0;
  assign f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_4_29_y0 = f_s_dadda_pg_rca32_and_4_29_y0;
  assign f_s_dadda_pg_rca32_fa371_y0 = f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_6_27_y0 ^ f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_5_28_y0;
  assign f_s_dadda_pg_rca32_fa371_y1 = f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_6_27_y0 & f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_5_28_y0;
  assign f_s_dadda_pg_rca32_fa371_y2 = f_s_dadda_pg_rca32_fa371_y0 ^ f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_4_29_y0;
  assign f_s_dadda_pg_rca32_fa371_y3 = f_s_dadda_pg_rca32_fa371_y0 & f_s_dadda_pg_rca32_fa371_f_s_dadda_pg_rca32_and_4_29_y0;
  assign f_s_dadda_pg_rca32_fa371_y4 = f_s_dadda_pg_rca32_fa371_y1 | f_s_dadda_pg_rca32_fa371_y3;
  assign f_s_dadda_pg_rca32_and_3_30_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_3_30_y0 = f_s_dadda_pg_rca32_and_3_30_a_3 & f_s_dadda_pg_rca32_and_3_30_b_30;
  assign f_s_dadda_pg_rca32_nand_2_31_a_2 = a_2;
  assign f_s_dadda_pg_rca32_nand_2_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_2_31_y0 = ~(f_s_dadda_pg_rca32_nand_2_31_a_2 & f_s_dadda_pg_rca32_nand_2_31_b_31);
  assign f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_and_3_30_y0 = f_s_dadda_pg_rca32_and_3_30_y0;
  assign f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_nand_2_31_y0 = f_s_dadda_pg_rca32_nand_2_31_y0;
  assign f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_fa10_y2 = f_s_dadda_pg_rca32_fa10_y2;
  assign f_s_dadda_pg_rca32_fa372_y0 = f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_and_3_30_y0 ^ f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_nand_2_31_y0;
  assign f_s_dadda_pg_rca32_fa372_y1 = f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_and_3_30_y0 & f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_nand_2_31_y0;
  assign f_s_dadda_pg_rca32_fa372_y2 = f_s_dadda_pg_rca32_fa372_y0 ^ f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_fa10_y2;
  assign f_s_dadda_pg_rca32_fa372_y3 = f_s_dadda_pg_rca32_fa372_y0 & f_s_dadda_pg_rca32_fa372_f_s_dadda_pg_rca32_fa10_y2;
  assign f_s_dadda_pg_rca32_fa372_y4 = f_s_dadda_pg_rca32_fa372_y1 | f_s_dadda_pg_rca32_fa372_y3;
  assign f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa11_y2 = f_s_dadda_pg_rca32_fa11_y2;
  assign f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa12_y2 = f_s_dadda_pg_rca32_fa12_y2;
  assign f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa357_y2 = f_s_dadda_pg_rca32_fa357_y2;
  assign f_s_dadda_pg_rca32_fa373_y0 = f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa11_y2 ^ f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa12_y2;
  assign f_s_dadda_pg_rca32_fa373_y1 = f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa11_y2 & f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa12_y2;
  assign f_s_dadda_pg_rca32_fa373_y2 = f_s_dadda_pg_rca32_fa373_y0 ^ f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa357_y2;
  assign f_s_dadda_pg_rca32_fa373_y3 = f_s_dadda_pg_rca32_fa373_y0 & f_s_dadda_pg_rca32_fa373_f_s_dadda_pg_rca32_fa357_y2;
  assign f_s_dadda_pg_rca32_fa373_y4 = f_s_dadda_pg_rca32_fa373_y1 | f_s_dadda_pg_rca32_fa373_y3;
  assign f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa358_y2 = f_s_dadda_pg_rca32_fa358_y2;
  assign f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa359_y2 = f_s_dadda_pg_rca32_fa359_y2;
  assign f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa360_y2 = f_s_dadda_pg_rca32_fa360_y2;
  assign f_s_dadda_pg_rca32_fa374_y0 = f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa358_y2 ^ f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa359_y2;
  assign f_s_dadda_pg_rca32_fa374_y1 = f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa358_y2 & f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa359_y2;
  assign f_s_dadda_pg_rca32_fa374_y2 = f_s_dadda_pg_rca32_fa374_y0 ^ f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa360_y2;
  assign f_s_dadda_pg_rca32_fa374_y3 = f_s_dadda_pg_rca32_fa374_y0 & f_s_dadda_pg_rca32_fa374_f_s_dadda_pg_rca32_fa360_y2;
  assign f_s_dadda_pg_rca32_fa374_y4 = f_s_dadda_pg_rca32_fa374_y1 | f_s_dadda_pg_rca32_fa374_y3;
  assign f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa361_y2 = f_s_dadda_pg_rca32_fa361_y2;
  assign f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa362_y2 = f_s_dadda_pg_rca32_fa362_y2;
  assign f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa363_y2 = f_s_dadda_pg_rca32_fa363_y2;
  assign f_s_dadda_pg_rca32_fa375_y0 = f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa361_y2 ^ f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa362_y2;
  assign f_s_dadda_pg_rca32_fa375_y1 = f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa361_y2 & f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa362_y2;
  assign f_s_dadda_pg_rca32_fa375_y2 = f_s_dadda_pg_rca32_fa375_y0 ^ f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa363_y2;
  assign f_s_dadda_pg_rca32_fa375_y3 = f_s_dadda_pg_rca32_fa375_y0 & f_s_dadda_pg_rca32_fa375_f_s_dadda_pg_rca32_fa363_y2;
  assign f_s_dadda_pg_rca32_fa375_y4 = f_s_dadda_pg_rca32_fa375_y1 | f_s_dadda_pg_rca32_fa375_y3;
  assign f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa364_y2 = f_s_dadda_pg_rca32_fa364_y2;
  assign f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa365_y2 = f_s_dadda_pg_rca32_fa365_y2;
  assign f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa366_y2 = f_s_dadda_pg_rca32_fa366_y2;
  assign f_s_dadda_pg_rca32_fa376_y0 = f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa364_y2 ^ f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa365_y2;
  assign f_s_dadda_pg_rca32_fa376_y1 = f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa364_y2 & f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa365_y2;
  assign f_s_dadda_pg_rca32_fa376_y2 = f_s_dadda_pg_rca32_fa376_y0 ^ f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa366_y2;
  assign f_s_dadda_pg_rca32_fa376_y3 = f_s_dadda_pg_rca32_fa376_y0 & f_s_dadda_pg_rca32_fa376_f_s_dadda_pg_rca32_fa366_y2;
  assign f_s_dadda_pg_rca32_fa376_y4 = f_s_dadda_pg_rca32_fa376_y1 | f_s_dadda_pg_rca32_fa376_y3;
  assign f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa367_y2 = f_s_dadda_pg_rca32_fa367_y2;
  assign f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa368_y2 = f_s_dadda_pg_rca32_fa368_y2;
  assign f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa369_y2 = f_s_dadda_pg_rca32_fa369_y2;
  assign f_s_dadda_pg_rca32_fa377_y0 = f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa367_y2 ^ f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa368_y2;
  assign f_s_dadda_pg_rca32_fa377_y1 = f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa367_y2 & f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa368_y2;
  assign f_s_dadda_pg_rca32_fa377_y2 = f_s_dadda_pg_rca32_fa377_y0 ^ f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa369_y2;
  assign f_s_dadda_pg_rca32_fa377_y3 = f_s_dadda_pg_rca32_fa377_y0 & f_s_dadda_pg_rca32_fa377_f_s_dadda_pg_rca32_fa369_y2;
  assign f_s_dadda_pg_rca32_fa377_y4 = f_s_dadda_pg_rca32_fa377_y1 | f_s_dadda_pg_rca32_fa377_y3;
  assign f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa370_y2 = f_s_dadda_pg_rca32_fa370_y2;
  assign f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa371_y2 = f_s_dadda_pg_rca32_fa371_y2;
  assign f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa372_y2 = f_s_dadda_pg_rca32_fa372_y2;
  assign f_s_dadda_pg_rca32_fa378_y0 = f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa370_y2 ^ f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa371_y2;
  assign f_s_dadda_pg_rca32_fa378_y1 = f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa370_y2 & f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa371_y2;
  assign f_s_dadda_pg_rca32_fa378_y2 = f_s_dadda_pg_rca32_fa378_y0 ^ f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa372_y2;
  assign f_s_dadda_pg_rca32_fa378_y3 = f_s_dadda_pg_rca32_fa378_y0 & f_s_dadda_pg_rca32_fa378_f_s_dadda_pg_rca32_fa372_y2;
  assign f_s_dadda_pg_rca32_fa378_y4 = f_s_dadda_pg_rca32_fa378_y1 | f_s_dadda_pg_rca32_fa378_y3;
  assign f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa378_y4 = f_s_dadda_pg_rca32_fa378_y4;
  assign f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa377_y4 = f_s_dadda_pg_rca32_fa377_y4;
  assign f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa376_y4 = f_s_dadda_pg_rca32_fa376_y4;
  assign f_s_dadda_pg_rca32_fa379_y0 = f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa378_y4 ^ f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa377_y4;
  assign f_s_dadda_pg_rca32_fa379_y1 = f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa378_y4 & f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa377_y4;
  assign f_s_dadda_pg_rca32_fa379_y2 = f_s_dadda_pg_rca32_fa379_y0 ^ f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa376_y4;
  assign f_s_dadda_pg_rca32_fa379_y3 = f_s_dadda_pg_rca32_fa379_y0 & f_s_dadda_pg_rca32_fa379_f_s_dadda_pg_rca32_fa376_y4;
  assign f_s_dadda_pg_rca32_fa379_y4 = f_s_dadda_pg_rca32_fa379_y1 | f_s_dadda_pg_rca32_fa379_y3;
  assign f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa375_y4 = f_s_dadda_pg_rca32_fa375_y4;
  assign f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa374_y4 = f_s_dadda_pg_rca32_fa374_y4;
  assign f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa373_y4 = f_s_dadda_pg_rca32_fa373_y4;
  assign f_s_dadda_pg_rca32_fa380_y0 = f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa375_y4 ^ f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa374_y4;
  assign f_s_dadda_pg_rca32_fa380_y1 = f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa375_y4 & f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa374_y4;
  assign f_s_dadda_pg_rca32_fa380_y2 = f_s_dadda_pg_rca32_fa380_y0 ^ f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa373_y4;
  assign f_s_dadda_pg_rca32_fa380_y3 = f_s_dadda_pg_rca32_fa380_y0 & f_s_dadda_pg_rca32_fa380_f_s_dadda_pg_rca32_fa373_y4;
  assign f_s_dadda_pg_rca32_fa380_y4 = f_s_dadda_pg_rca32_fa380_y1 | f_s_dadda_pg_rca32_fa380_y3;
  assign f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa372_y4 = f_s_dadda_pg_rca32_fa372_y4;
  assign f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa371_y4 = f_s_dadda_pg_rca32_fa371_y4;
  assign f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa370_y4 = f_s_dadda_pg_rca32_fa370_y4;
  assign f_s_dadda_pg_rca32_fa381_y0 = f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa372_y4 ^ f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa371_y4;
  assign f_s_dadda_pg_rca32_fa381_y1 = f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa372_y4 & f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa371_y4;
  assign f_s_dadda_pg_rca32_fa381_y2 = f_s_dadda_pg_rca32_fa381_y0 ^ f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa370_y4;
  assign f_s_dadda_pg_rca32_fa381_y3 = f_s_dadda_pg_rca32_fa381_y0 & f_s_dadda_pg_rca32_fa381_f_s_dadda_pg_rca32_fa370_y4;
  assign f_s_dadda_pg_rca32_fa381_y4 = f_s_dadda_pg_rca32_fa381_y1 | f_s_dadda_pg_rca32_fa381_y3;
  assign f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa369_y4 = f_s_dadda_pg_rca32_fa369_y4;
  assign f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa368_y4 = f_s_dadda_pg_rca32_fa368_y4;
  assign f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa367_y4 = f_s_dadda_pg_rca32_fa367_y4;
  assign f_s_dadda_pg_rca32_fa382_y0 = f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa369_y4 ^ f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa368_y4;
  assign f_s_dadda_pg_rca32_fa382_y1 = f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa369_y4 & f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa368_y4;
  assign f_s_dadda_pg_rca32_fa382_y2 = f_s_dadda_pg_rca32_fa382_y0 ^ f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa367_y4;
  assign f_s_dadda_pg_rca32_fa382_y3 = f_s_dadda_pg_rca32_fa382_y0 & f_s_dadda_pg_rca32_fa382_f_s_dadda_pg_rca32_fa367_y4;
  assign f_s_dadda_pg_rca32_fa382_y4 = f_s_dadda_pg_rca32_fa382_y1 | f_s_dadda_pg_rca32_fa382_y3;
  assign f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa366_y4 = f_s_dadda_pg_rca32_fa366_y4;
  assign f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa365_y4 = f_s_dadda_pg_rca32_fa365_y4;
  assign f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa364_y4 = f_s_dadda_pg_rca32_fa364_y4;
  assign f_s_dadda_pg_rca32_fa383_y0 = f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa366_y4 ^ f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa365_y4;
  assign f_s_dadda_pg_rca32_fa383_y1 = f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa366_y4 & f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa365_y4;
  assign f_s_dadda_pg_rca32_fa383_y2 = f_s_dadda_pg_rca32_fa383_y0 ^ f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa364_y4;
  assign f_s_dadda_pg_rca32_fa383_y3 = f_s_dadda_pg_rca32_fa383_y0 & f_s_dadda_pg_rca32_fa383_f_s_dadda_pg_rca32_fa364_y4;
  assign f_s_dadda_pg_rca32_fa383_y4 = f_s_dadda_pg_rca32_fa383_y1 | f_s_dadda_pg_rca32_fa383_y3;
  assign f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa363_y4 = f_s_dadda_pg_rca32_fa363_y4;
  assign f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa362_y4 = f_s_dadda_pg_rca32_fa362_y4;
  assign f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa361_y4 = f_s_dadda_pg_rca32_fa361_y4;
  assign f_s_dadda_pg_rca32_fa384_y0 = f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa363_y4 ^ f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa362_y4;
  assign f_s_dadda_pg_rca32_fa384_y1 = f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa363_y4 & f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa362_y4;
  assign f_s_dadda_pg_rca32_fa384_y2 = f_s_dadda_pg_rca32_fa384_y0 ^ f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa361_y4;
  assign f_s_dadda_pg_rca32_fa384_y3 = f_s_dadda_pg_rca32_fa384_y0 & f_s_dadda_pg_rca32_fa384_f_s_dadda_pg_rca32_fa361_y4;
  assign f_s_dadda_pg_rca32_fa384_y4 = f_s_dadda_pg_rca32_fa384_y1 | f_s_dadda_pg_rca32_fa384_y3;
  assign f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa360_y4 = f_s_dadda_pg_rca32_fa360_y4;
  assign f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa359_y4 = f_s_dadda_pg_rca32_fa359_y4;
  assign f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa358_y4 = f_s_dadda_pg_rca32_fa358_y4;
  assign f_s_dadda_pg_rca32_fa385_y0 = f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa360_y4 ^ f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa359_y4;
  assign f_s_dadda_pg_rca32_fa385_y1 = f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa360_y4 & f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa359_y4;
  assign f_s_dadda_pg_rca32_fa385_y2 = f_s_dadda_pg_rca32_fa385_y0 ^ f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa358_y4;
  assign f_s_dadda_pg_rca32_fa385_y3 = f_s_dadda_pg_rca32_fa385_y0 & f_s_dadda_pg_rca32_fa385_f_s_dadda_pg_rca32_fa358_y4;
  assign f_s_dadda_pg_rca32_fa385_y4 = f_s_dadda_pg_rca32_fa385_y1 | f_s_dadda_pg_rca32_fa385_y3;
  assign f_s_dadda_pg_rca32_and_28_6_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_28_6_y0 = f_s_dadda_pg_rca32_and_28_6_a_28 & f_s_dadda_pg_rca32_and_28_6_b_6;
  assign f_s_dadda_pg_rca32_and_27_7_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_27_7_y0 = f_s_dadda_pg_rca32_and_27_7_a_27 & f_s_dadda_pg_rca32_and_27_7_b_7;
  assign f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_fa357_y4 = f_s_dadda_pg_rca32_fa357_y4;
  assign f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_and_28_6_y0 = f_s_dadda_pg_rca32_and_28_6_y0;
  assign f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_and_27_7_y0 = f_s_dadda_pg_rca32_and_27_7_y0;
  assign f_s_dadda_pg_rca32_fa386_y0 = f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_fa357_y4 ^ f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_and_28_6_y0;
  assign f_s_dadda_pg_rca32_fa386_y1 = f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_fa357_y4 & f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_and_28_6_y0;
  assign f_s_dadda_pg_rca32_fa386_y2 = f_s_dadda_pg_rca32_fa386_y0 ^ f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_and_27_7_y0;
  assign f_s_dadda_pg_rca32_fa386_y3 = f_s_dadda_pg_rca32_fa386_y0 & f_s_dadda_pg_rca32_fa386_f_s_dadda_pg_rca32_and_27_7_y0;
  assign f_s_dadda_pg_rca32_fa386_y4 = f_s_dadda_pg_rca32_fa386_y1 | f_s_dadda_pg_rca32_fa386_y3;
  assign f_s_dadda_pg_rca32_and_26_8_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_26_8_y0 = f_s_dadda_pg_rca32_and_26_8_a_26 & f_s_dadda_pg_rca32_and_26_8_b_8;
  assign f_s_dadda_pg_rca32_and_25_9_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_25_9_y0 = f_s_dadda_pg_rca32_and_25_9_a_25 & f_s_dadda_pg_rca32_and_25_9_b_9;
  assign f_s_dadda_pg_rca32_and_24_10_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_24_10_y0 = f_s_dadda_pg_rca32_and_24_10_a_24 & f_s_dadda_pg_rca32_and_24_10_b_10;
  assign f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_26_8_y0 = f_s_dadda_pg_rca32_and_26_8_y0;
  assign f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_25_9_y0 = f_s_dadda_pg_rca32_and_25_9_y0;
  assign f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_24_10_y0 = f_s_dadda_pg_rca32_and_24_10_y0;
  assign f_s_dadda_pg_rca32_fa387_y0 = f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_26_8_y0 ^ f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_25_9_y0;
  assign f_s_dadda_pg_rca32_fa387_y1 = f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_26_8_y0 & f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_25_9_y0;
  assign f_s_dadda_pg_rca32_fa387_y2 = f_s_dadda_pg_rca32_fa387_y0 ^ f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_24_10_y0;
  assign f_s_dadda_pg_rca32_fa387_y3 = f_s_dadda_pg_rca32_fa387_y0 & f_s_dadda_pg_rca32_fa387_f_s_dadda_pg_rca32_and_24_10_y0;
  assign f_s_dadda_pg_rca32_fa387_y4 = f_s_dadda_pg_rca32_fa387_y1 | f_s_dadda_pg_rca32_fa387_y3;
  assign f_s_dadda_pg_rca32_and_23_11_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_23_11_y0 = f_s_dadda_pg_rca32_and_23_11_a_23 & f_s_dadda_pg_rca32_and_23_11_b_11;
  assign f_s_dadda_pg_rca32_and_22_12_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_22_12_y0 = f_s_dadda_pg_rca32_and_22_12_a_22 & f_s_dadda_pg_rca32_and_22_12_b_12;
  assign f_s_dadda_pg_rca32_and_21_13_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_21_13_y0 = f_s_dadda_pg_rca32_and_21_13_a_21 & f_s_dadda_pg_rca32_and_21_13_b_13;
  assign f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_23_11_y0 = f_s_dadda_pg_rca32_and_23_11_y0;
  assign f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_22_12_y0 = f_s_dadda_pg_rca32_and_22_12_y0;
  assign f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_21_13_y0 = f_s_dadda_pg_rca32_and_21_13_y0;
  assign f_s_dadda_pg_rca32_fa388_y0 = f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_23_11_y0 ^ f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_22_12_y0;
  assign f_s_dadda_pg_rca32_fa388_y1 = f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_23_11_y0 & f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_22_12_y0;
  assign f_s_dadda_pg_rca32_fa388_y2 = f_s_dadda_pg_rca32_fa388_y0 ^ f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_21_13_y0;
  assign f_s_dadda_pg_rca32_fa388_y3 = f_s_dadda_pg_rca32_fa388_y0 & f_s_dadda_pg_rca32_fa388_f_s_dadda_pg_rca32_and_21_13_y0;
  assign f_s_dadda_pg_rca32_fa388_y4 = f_s_dadda_pg_rca32_fa388_y1 | f_s_dadda_pg_rca32_fa388_y3;
  assign f_s_dadda_pg_rca32_and_20_14_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_20_14_y0 = f_s_dadda_pg_rca32_and_20_14_a_20 & f_s_dadda_pg_rca32_and_20_14_b_14;
  assign f_s_dadda_pg_rca32_and_19_15_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_19_15_y0 = f_s_dadda_pg_rca32_and_19_15_a_19 & f_s_dadda_pg_rca32_and_19_15_b_15;
  assign f_s_dadda_pg_rca32_and_18_16_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_18_16_y0 = f_s_dadda_pg_rca32_and_18_16_a_18 & f_s_dadda_pg_rca32_and_18_16_b_16;
  assign f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_20_14_y0 = f_s_dadda_pg_rca32_and_20_14_y0;
  assign f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_19_15_y0 = f_s_dadda_pg_rca32_and_19_15_y0;
  assign f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_18_16_y0 = f_s_dadda_pg_rca32_and_18_16_y0;
  assign f_s_dadda_pg_rca32_fa389_y0 = f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_20_14_y0 ^ f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_19_15_y0;
  assign f_s_dadda_pg_rca32_fa389_y1 = f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_20_14_y0 & f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_19_15_y0;
  assign f_s_dadda_pg_rca32_fa389_y2 = f_s_dadda_pg_rca32_fa389_y0 ^ f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_18_16_y0;
  assign f_s_dadda_pg_rca32_fa389_y3 = f_s_dadda_pg_rca32_fa389_y0 & f_s_dadda_pg_rca32_fa389_f_s_dadda_pg_rca32_and_18_16_y0;
  assign f_s_dadda_pg_rca32_fa389_y4 = f_s_dadda_pg_rca32_fa389_y1 | f_s_dadda_pg_rca32_fa389_y3;
  assign f_s_dadda_pg_rca32_and_17_17_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_17_17_y0 = f_s_dadda_pg_rca32_and_17_17_a_17 & f_s_dadda_pg_rca32_and_17_17_b_17;
  assign f_s_dadda_pg_rca32_and_16_18_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_16_18_y0 = f_s_dadda_pg_rca32_and_16_18_a_16 & f_s_dadda_pg_rca32_and_16_18_b_18;
  assign f_s_dadda_pg_rca32_and_15_19_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_15_19_y0 = f_s_dadda_pg_rca32_and_15_19_a_15 & f_s_dadda_pg_rca32_and_15_19_b_19;
  assign f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_17_17_y0 = f_s_dadda_pg_rca32_and_17_17_y0;
  assign f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_16_18_y0 = f_s_dadda_pg_rca32_and_16_18_y0;
  assign f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_15_19_y0 = f_s_dadda_pg_rca32_and_15_19_y0;
  assign f_s_dadda_pg_rca32_fa390_y0 = f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_17_17_y0 ^ f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_16_18_y0;
  assign f_s_dadda_pg_rca32_fa390_y1 = f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_17_17_y0 & f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_16_18_y0;
  assign f_s_dadda_pg_rca32_fa390_y2 = f_s_dadda_pg_rca32_fa390_y0 ^ f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_15_19_y0;
  assign f_s_dadda_pg_rca32_fa390_y3 = f_s_dadda_pg_rca32_fa390_y0 & f_s_dadda_pg_rca32_fa390_f_s_dadda_pg_rca32_and_15_19_y0;
  assign f_s_dadda_pg_rca32_fa390_y4 = f_s_dadda_pg_rca32_fa390_y1 | f_s_dadda_pg_rca32_fa390_y3;
  assign f_s_dadda_pg_rca32_and_14_20_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_14_20_y0 = f_s_dadda_pg_rca32_and_14_20_a_14 & f_s_dadda_pg_rca32_and_14_20_b_20;
  assign f_s_dadda_pg_rca32_and_13_21_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_13_21_y0 = f_s_dadda_pg_rca32_and_13_21_a_13 & f_s_dadda_pg_rca32_and_13_21_b_21;
  assign f_s_dadda_pg_rca32_and_12_22_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_12_22_y0 = f_s_dadda_pg_rca32_and_12_22_a_12 & f_s_dadda_pg_rca32_and_12_22_b_22;
  assign f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_14_20_y0 = f_s_dadda_pg_rca32_and_14_20_y0;
  assign f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_13_21_y0 = f_s_dadda_pg_rca32_and_13_21_y0;
  assign f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_12_22_y0 = f_s_dadda_pg_rca32_and_12_22_y0;
  assign f_s_dadda_pg_rca32_fa391_y0 = f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_14_20_y0 ^ f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_13_21_y0;
  assign f_s_dadda_pg_rca32_fa391_y1 = f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_14_20_y0 & f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_13_21_y0;
  assign f_s_dadda_pg_rca32_fa391_y2 = f_s_dadda_pg_rca32_fa391_y0 ^ f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_12_22_y0;
  assign f_s_dadda_pg_rca32_fa391_y3 = f_s_dadda_pg_rca32_fa391_y0 & f_s_dadda_pg_rca32_fa391_f_s_dadda_pg_rca32_and_12_22_y0;
  assign f_s_dadda_pg_rca32_fa391_y4 = f_s_dadda_pg_rca32_fa391_y1 | f_s_dadda_pg_rca32_fa391_y3;
  assign f_s_dadda_pg_rca32_and_11_23_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_11_23_y0 = f_s_dadda_pg_rca32_and_11_23_a_11 & f_s_dadda_pg_rca32_and_11_23_b_23;
  assign f_s_dadda_pg_rca32_and_10_24_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_10_24_y0 = f_s_dadda_pg_rca32_and_10_24_a_10 & f_s_dadda_pg_rca32_and_10_24_b_24;
  assign f_s_dadda_pg_rca32_and_9_25_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_9_25_y0 = f_s_dadda_pg_rca32_and_9_25_a_9 & f_s_dadda_pg_rca32_and_9_25_b_25;
  assign f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_11_23_y0 = f_s_dadda_pg_rca32_and_11_23_y0;
  assign f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_10_24_y0 = f_s_dadda_pg_rca32_and_10_24_y0;
  assign f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_9_25_y0 = f_s_dadda_pg_rca32_and_9_25_y0;
  assign f_s_dadda_pg_rca32_fa392_y0 = f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_11_23_y0 ^ f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_10_24_y0;
  assign f_s_dadda_pg_rca32_fa392_y1 = f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_11_23_y0 & f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_10_24_y0;
  assign f_s_dadda_pg_rca32_fa392_y2 = f_s_dadda_pg_rca32_fa392_y0 ^ f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_9_25_y0;
  assign f_s_dadda_pg_rca32_fa392_y3 = f_s_dadda_pg_rca32_fa392_y0 & f_s_dadda_pg_rca32_fa392_f_s_dadda_pg_rca32_and_9_25_y0;
  assign f_s_dadda_pg_rca32_fa392_y4 = f_s_dadda_pg_rca32_fa392_y1 | f_s_dadda_pg_rca32_fa392_y3;
  assign f_s_dadda_pg_rca32_and_8_26_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_8_26_y0 = f_s_dadda_pg_rca32_and_8_26_a_8 & f_s_dadda_pg_rca32_and_8_26_b_26;
  assign f_s_dadda_pg_rca32_and_7_27_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_7_27_y0 = f_s_dadda_pg_rca32_and_7_27_a_7 & f_s_dadda_pg_rca32_and_7_27_b_27;
  assign f_s_dadda_pg_rca32_and_6_28_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_6_28_y0 = f_s_dadda_pg_rca32_and_6_28_a_6 & f_s_dadda_pg_rca32_and_6_28_b_28;
  assign f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_8_26_y0 = f_s_dadda_pg_rca32_and_8_26_y0;
  assign f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_7_27_y0 = f_s_dadda_pg_rca32_and_7_27_y0;
  assign f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_6_28_y0 = f_s_dadda_pg_rca32_and_6_28_y0;
  assign f_s_dadda_pg_rca32_fa393_y0 = f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_8_26_y0 ^ f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_7_27_y0;
  assign f_s_dadda_pg_rca32_fa393_y1 = f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_8_26_y0 & f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_7_27_y0;
  assign f_s_dadda_pg_rca32_fa393_y2 = f_s_dadda_pg_rca32_fa393_y0 ^ f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_6_28_y0;
  assign f_s_dadda_pg_rca32_fa393_y3 = f_s_dadda_pg_rca32_fa393_y0 & f_s_dadda_pg_rca32_fa393_f_s_dadda_pg_rca32_and_6_28_y0;
  assign f_s_dadda_pg_rca32_fa393_y4 = f_s_dadda_pg_rca32_fa393_y1 | f_s_dadda_pg_rca32_fa393_y3;
  assign f_s_dadda_pg_rca32_and_5_29_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_5_29_y0 = f_s_dadda_pg_rca32_and_5_29_a_5 & f_s_dadda_pg_rca32_and_5_29_b_29;
  assign f_s_dadda_pg_rca32_and_4_30_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_4_30_y0 = f_s_dadda_pg_rca32_and_4_30_a_4 & f_s_dadda_pg_rca32_and_4_30_b_30;
  assign f_s_dadda_pg_rca32_nand_3_31_a_3 = a_3;
  assign f_s_dadda_pg_rca32_nand_3_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_3_31_y0 = ~(f_s_dadda_pg_rca32_nand_3_31_a_3 & f_s_dadda_pg_rca32_nand_3_31_b_31);
  assign f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_and_5_29_y0 = f_s_dadda_pg_rca32_and_5_29_y0;
  assign f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_and_4_30_y0 = f_s_dadda_pg_rca32_and_4_30_y0;
  assign f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_nand_3_31_y0 = f_s_dadda_pg_rca32_nand_3_31_y0;
  assign f_s_dadda_pg_rca32_fa394_y0 = f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_and_5_29_y0 ^ f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_and_4_30_y0;
  assign f_s_dadda_pg_rca32_fa394_y1 = f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_and_5_29_y0 & f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_and_4_30_y0;
  assign f_s_dadda_pg_rca32_fa394_y2 = f_s_dadda_pg_rca32_fa394_y0 ^ f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_nand_3_31_y0;
  assign f_s_dadda_pg_rca32_fa394_y3 = f_s_dadda_pg_rca32_fa394_y0 & f_s_dadda_pg_rca32_fa394_f_s_dadda_pg_rca32_nand_3_31_y0;
  assign f_s_dadda_pg_rca32_fa394_y4 = f_s_dadda_pg_rca32_fa394_y1 | f_s_dadda_pg_rca32_fa394_y3;
  assign f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa13_y2 = f_s_dadda_pg_rca32_fa13_y2;
  assign f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa14_y2 = f_s_dadda_pg_rca32_fa14_y2;
  assign f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa379_y2 = f_s_dadda_pg_rca32_fa379_y2;
  assign f_s_dadda_pg_rca32_fa395_y0 = f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa13_y2 ^ f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa14_y2;
  assign f_s_dadda_pg_rca32_fa395_y1 = f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa13_y2 & f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa14_y2;
  assign f_s_dadda_pg_rca32_fa395_y2 = f_s_dadda_pg_rca32_fa395_y0 ^ f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa379_y2;
  assign f_s_dadda_pg_rca32_fa395_y3 = f_s_dadda_pg_rca32_fa395_y0 & f_s_dadda_pg_rca32_fa395_f_s_dadda_pg_rca32_fa379_y2;
  assign f_s_dadda_pg_rca32_fa395_y4 = f_s_dadda_pg_rca32_fa395_y1 | f_s_dadda_pg_rca32_fa395_y3;
  assign f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa380_y2 = f_s_dadda_pg_rca32_fa380_y2;
  assign f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa381_y2 = f_s_dadda_pg_rca32_fa381_y2;
  assign f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa382_y2 = f_s_dadda_pg_rca32_fa382_y2;
  assign f_s_dadda_pg_rca32_fa396_y0 = f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa380_y2 ^ f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa381_y2;
  assign f_s_dadda_pg_rca32_fa396_y1 = f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa380_y2 & f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa381_y2;
  assign f_s_dadda_pg_rca32_fa396_y2 = f_s_dadda_pg_rca32_fa396_y0 ^ f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa382_y2;
  assign f_s_dadda_pg_rca32_fa396_y3 = f_s_dadda_pg_rca32_fa396_y0 & f_s_dadda_pg_rca32_fa396_f_s_dadda_pg_rca32_fa382_y2;
  assign f_s_dadda_pg_rca32_fa396_y4 = f_s_dadda_pg_rca32_fa396_y1 | f_s_dadda_pg_rca32_fa396_y3;
  assign f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa383_y2 = f_s_dadda_pg_rca32_fa383_y2;
  assign f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa384_y2 = f_s_dadda_pg_rca32_fa384_y2;
  assign f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa385_y2 = f_s_dadda_pg_rca32_fa385_y2;
  assign f_s_dadda_pg_rca32_fa397_y0 = f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa383_y2 ^ f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa384_y2;
  assign f_s_dadda_pg_rca32_fa397_y1 = f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa383_y2 & f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa384_y2;
  assign f_s_dadda_pg_rca32_fa397_y2 = f_s_dadda_pg_rca32_fa397_y0 ^ f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa385_y2;
  assign f_s_dadda_pg_rca32_fa397_y3 = f_s_dadda_pg_rca32_fa397_y0 & f_s_dadda_pg_rca32_fa397_f_s_dadda_pg_rca32_fa385_y2;
  assign f_s_dadda_pg_rca32_fa397_y4 = f_s_dadda_pg_rca32_fa397_y1 | f_s_dadda_pg_rca32_fa397_y3;
  assign f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa386_y2 = f_s_dadda_pg_rca32_fa386_y2;
  assign f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa387_y2 = f_s_dadda_pg_rca32_fa387_y2;
  assign f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa388_y2 = f_s_dadda_pg_rca32_fa388_y2;
  assign f_s_dadda_pg_rca32_fa398_y0 = f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa386_y2 ^ f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa387_y2;
  assign f_s_dadda_pg_rca32_fa398_y1 = f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa386_y2 & f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa387_y2;
  assign f_s_dadda_pg_rca32_fa398_y2 = f_s_dadda_pg_rca32_fa398_y0 ^ f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa388_y2;
  assign f_s_dadda_pg_rca32_fa398_y3 = f_s_dadda_pg_rca32_fa398_y0 & f_s_dadda_pg_rca32_fa398_f_s_dadda_pg_rca32_fa388_y2;
  assign f_s_dadda_pg_rca32_fa398_y4 = f_s_dadda_pg_rca32_fa398_y1 | f_s_dadda_pg_rca32_fa398_y3;
  assign f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa389_y2 = f_s_dadda_pg_rca32_fa389_y2;
  assign f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa390_y2 = f_s_dadda_pg_rca32_fa390_y2;
  assign f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa391_y2 = f_s_dadda_pg_rca32_fa391_y2;
  assign f_s_dadda_pg_rca32_fa399_y0 = f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa389_y2 ^ f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa390_y2;
  assign f_s_dadda_pg_rca32_fa399_y1 = f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa389_y2 & f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa390_y2;
  assign f_s_dadda_pg_rca32_fa399_y2 = f_s_dadda_pg_rca32_fa399_y0 ^ f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa391_y2;
  assign f_s_dadda_pg_rca32_fa399_y3 = f_s_dadda_pg_rca32_fa399_y0 & f_s_dadda_pg_rca32_fa399_f_s_dadda_pg_rca32_fa391_y2;
  assign f_s_dadda_pg_rca32_fa399_y4 = f_s_dadda_pg_rca32_fa399_y1 | f_s_dadda_pg_rca32_fa399_y3;
  assign f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa392_y2 = f_s_dadda_pg_rca32_fa392_y2;
  assign f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa393_y2 = f_s_dadda_pg_rca32_fa393_y2;
  assign f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa394_y2 = f_s_dadda_pg_rca32_fa394_y2;
  assign f_s_dadda_pg_rca32_fa400_y0 = f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa392_y2 ^ f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa393_y2;
  assign f_s_dadda_pg_rca32_fa400_y1 = f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa392_y2 & f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa393_y2;
  assign f_s_dadda_pg_rca32_fa400_y2 = f_s_dadda_pg_rca32_fa400_y0 ^ f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa394_y2;
  assign f_s_dadda_pg_rca32_fa400_y3 = f_s_dadda_pg_rca32_fa400_y0 & f_s_dadda_pg_rca32_fa400_f_s_dadda_pg_rca32_fa394_y2;
  assign f_s_dadda_pg_rca32_fa400_y4 = f_s_dadda_pg_rca32_fa400_y1 | f_s_dadda_pg_rca32_fa400_y3;
  assign f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa400_y4 = f_s_dadda_pg_rca32_fa400_y4;
  assign f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa399_y4 = f_s_dadda_pg_rca32_fa399_y4;
  assign f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa398_y4 = f_s_dadda_pg_rca32_fa398_y4;
  assign f_s_dadda_pg_rca32_fa401_y0 = f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa400_y4 ^ f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa399_y4;
  assign f_s_dadda_pg_rca32_fa401_y1 = f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa400_y4 & f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa399_y4;
  assign f_s_dadda_pg_rca32_fa401_y2 = f_s_dadda_pg_rca32_fa401_y0 ^ f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa398_y4;
  assign f_s_dadda_pg_rca32_fa401_y3 = f_s_dadda_pg_rca32_fa401_y0 & f_s_dadda_pg_rca32_fa401_f_s_dadda_pg_rca32_fa398_y4;
  assign f_s_dadda_pg_rca32_fa401_y4 = f_s_dadda_pg_rca32_fa401_y1 | f_s_dadda_pg_rca32_fa401_y3;
  assign f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa397_y4 = f_s_dadda_pg_rca32_fa397_y4;
  assign f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa396_y4 = f_s_dadda_pg_rca32_fa396_y4;
  assign f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa395_y4 = f_s_dadda_pg_rca32_fa395_y4;
  assign f_s_dadda_pg_rca32_fa402_y0 = f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa397_y4 ^ f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa396_y4;
  assign f_s_dadda_pg_rca32_fa402_y1 = f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa397_y4 & f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa396_y4;
  assign f_s_dadda_pg_rca32_fa402_y2 = f_s_dadda_pg_rca32_fa402_y0 ^ f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa395_y4;
  assign f_s_dadda_pg_rca32_fa402_y3 = f_s_dadda_pg_rca32_fa402_y0 & f_s_dadda_pg_rca32_fa402_f_s_dadda_pg_rca32_fa395_y4;
  assign f_s_dadda_pg_rca32_fa402_y4 = f_s_dadda_pg_rca32_fa402_y1 | f_s_dadda_pg_rca32_fa402_y3;
  assign f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa394_y4 = f_s_dadda_pg_rca32_fa394_y4;
  assign f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa393_y4 = f_s_dadda_pg_rca32_fa393_y4;
  assign f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa392_y4 = f_s_dadda_pg_rca32_fa392_y4;
  assign f_s_dadda_pg_rca32_fa403_y0 = f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa394_y4 ^ f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa393_y4;
  assign f_s_dadda_pg_rca32_fa403_y1 = f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa394_y4 & f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa393_y4;
  assign f_s_dadda_pg_rca32_fa403_y2 = f_s_dadda_pg_rca32_fa403_y0 ^ f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa392_y4;
  assign f_s_dadda_pg_rca32_fa403_y3 = f_s_dadda_pg_rca32_fa403_y0 & f_s_dadda_pg_rca32_fa403_f_s_dadda_pg_rca32_fa392_y4;
  assign f_s_dadda_pg_rca32_fa403_y4 = f_s_dadda_pg_rca32_fa403_y1 | f_s_dadda_pg_rca32_fa403_y3;
  assign f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa391_y4 = f_s_dadda_pg_rca32_fa391_y4;
  assign f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa390_y4 = f_s_dadda_pg_rca32_fa390_y4;
  assign f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa389_y4 = f_s_dadda_pg_rca32_fa389_y4;
  assign f_s_dadda_pg_rca32_fa404_y0 = f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa391_y4 ^ f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa390_y4;
  assign f_s_dadda_pg_rca32_fa404_y1 = f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa391_y4 & f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa390_y4;
  assign f_s_dadda_pg_rca32_fa404_y2 = f_s_dadda_pg_rca32_fa404_y0 ^ f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa389_y4;
  assign f_s_dadda_pg_rca32_fa404_y3 = f_s_dadda_pg_rca32_fa404_y0 & f_s_dadda_pg_rca32_fa404_f_s_dadda_pg_rca32_fa389_y4;
  assign f_s_dadda_pg_rca32_fa404_y4 = f_s_dadda_pg_rca32_fa404_y1 | f_s_dadda_pg_rca32_fa404_y3;
  assign f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa388_y4 = f_s_dadda_pg_rca32_fa388_y4;
  assign f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa387_y4 = f_s_dadda_pg_rca32_fa387_y4;
  assign f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa386_y4 = f_s_dadda_pg_rca32_fa386_y4;
  assign f_s_dadda_pg_rca32_fa405_y0 = f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa388_y4 ^ f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa387_y4;
  assign f_s_dadda_pg_rca32_fa405_y1 = f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa388_y4 & f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa387_y4;
  assign f_s_dadda_pg_rca32_fa405_y2 = f_s_dadda_pg_rca32_fa405_y0 ^ f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa386_y4;
  assign f_s_dadda_pg_rca32_fa405_y3 = f_s_dadda_pg_rca32_fa405_y0 & f_s_dadda_pg_rca32_fa405_f_s_dadda_pg_rca32_fa386_y4;
  assign f_s_dadda_pg_rca32_fa405_y4 = f_s_dadda_pg_rca32_fa405_y1 | f_s_dadda_pg_rca32_fa405_y3;
  assign f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa385_y4 = f_s_dadda_pg_rca32_fa385_y4;
  assign f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa384_y4 = f_s_dadda_pg_rca32_fa384_y4;
  assign f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa383_y4 = f_s_dadda_pg_rca32_fa383_y4;
  assign f_s_dadda_pg_rca32_fa406_y0 = f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa385_y4 ^ f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa384_y4;
  assign f_s_dadda_pg_rca32_fa406_y1 = f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa385_y4 & f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa384_y4;
  assign f_s_dadda_pg_rca32_fa406_y2 = f_s_dadda_pg_rca32_fa406_y0 ^ f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa383_y4;
  assign f_s_dadda_pg_rca32_fa406_y3 = f_s_dadda_pg_rca32_fa406_y0 & f_s_dadda_pg_rca32_fa406_f_s_dadda_pg_rca32_fa383_y4;
  assign f_s_dadda_pg_rca32_fa406_y4 = f_s_dadda_pg_rca32_fa406_y1 | f_s_dadda_pg_rca32_fa406_y3;
  assign f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa382_y4 = f_s_dadda_pg_rca32_fa382_y4;
  assign f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa381_y4 = f_s_dadda_pg_rca32_fa381_y4;
  assign f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa380_y4 = f_s_dadda_pg_rca32_fa380_y4;
  assign f_s_dadda_pg_rca32_fa407_y0 = f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa382_y4 ^ f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa381_y4;
  assign f_s_dadda_pg_rca32_fa407_y1 = f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa382_y4 & f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa381_y4;
  assign f_s_dadda_pg_rca32_fa407_y2 = f_s_dadda_pg_rca32_fa407_y0 ^ f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa380_y4;
  assign f_s_dadda_pg_rca32_fa407_y3 = f_s_dadda_pg_rca32_fa407_y0 & f_s_dadda_pg_rca32_fa407_f_s_dadda_pg_rca32_fa380_y4;
  assign f_s_dadda_pg_rca32_fa407_y4 = f_s_dadda_pg_rca32_fa407_y1 | f_s_dadda_pg_rca32_fa407_y3;
  assign f_s_dadda_pg_rca32_and_30_5_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_30_5_y0 = f_s_dadda_pg_rca32_and_30_5_a_30 & f_s_dadda_pg_rca32_and_30_5_b_5;
  assign f_s_dadda_pg_rca32_and_29_6_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_29_6_y0 = f_s_dadda_pg_rca32_and_29_6_a_29 & f_s_dadda_pg_rca32_and_29_6_b_6;
  assign f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_fa379_y4 = f_s_dadda_pg_rca32_fa379_y4;
  assign f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_and_30_5_y0 = f_s_dadda_pg_rca32_and_30_5_y0;
  assign f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_and_29_6_y0 = f_s_dadda_pg_rca32_and_29_6_y0;
  assign f_s_dadda_pg_rca32_fa408_y0 = f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_fa379_y4 ^ f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_and_30_5_y0;
  assign f_s_dadda_pg_rca32_fa408_y1 = f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_fa379_y4 & f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_and_30_5_y0;
  assign f_s_dadda_pg_rca32_fa408_y2 = f_s_dadda_pg_rca32_fa408_y0 ^ f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_and_29_6_y0;
  assign f_s_dadda_pg_rca32_fa408_y3 = f_s_dadda_pg_rca32_fa408_y0 & f_s_dadda_pg_rca32_fa408_f_s_dadda_pg_rca32_and_29_6_y0;
  assign f_s_dadda_pg_rca32_fa408_y4 = f_s_dadda_pg_rca32_fa408_y1 | f_s_dadda_pg_rca32_fa408_y3;
  assign f_s_dadda_pg_rca32_and_28_7_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_28_7_y0 = f_s_dadda_pg_rca32_and_28_7_a_28 & f_s_dadda_pg_rca32_and_28_7_b_7;
  assign f_s_dadda_pg_rca32_and_27_8_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_27_8_y0 = f_s_dadda_pg_rca32_and_27_8_a_27 & f_s_dadda_pg_rca32_and_27_8_b_8;
  assign f_s_dadda_pg_rca32_and_26_9_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_26_9_y0 = f_s_dadda_pg_rca32_and_26_9_a_26 & f_s_dadda_pg_rca32_and_26_9_b_9;
  assign f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_28_7_y0 = f_s_dadda_pg_rca32_and_28_7_y0;
  assign f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_27_8_y0 = f_s_dadda_pg_rca32_and_27_8_y0;
  assign f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_26_9_y0 = f_s_dadda_pg_rca32_and_26_9_y0;
  assign f_s_dadda_pg_rca32_fa409_y0 = f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_28_7_y0 ^ f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_27_8_y0;
  assign f_s_dadda_pg_rca32_fa409_y1 = f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_28_7_y0 & f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_27_8_y0;
  assign f_s_dadda_pg_rca32_fa409_y2 = f_s_dadda_pg_rca32_fa409_y0 ^ f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_26_9_y0;
  assign f_s_dadda_pg_rca32_fa409_y3 = f_s_dadda_pg_rca32_fa409_y0 & f_s_dadda_pg_rca32_fa409_f_s_dadda_pg_rca32_and_26_9_y0;
  assign f_s_dadda_pg_rca32_fa409_y4 = f_s_dadda_pg_rca32_fa409_y1 | f_s_dadda_pg_rca32_fa409_y3;
  assign f_s_dadda_pg_rca32_and_25_10_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_25_10_y0 = f_s_dadda_pg_rca32_and_25_10_a_25 & f_s_dadda_pg_rca32_and_25_10_b_10;
  assign f_s_dadda_pg_rca32_and_24_11_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_24_11_y0 = f_s_dadda_pg_rca32_and_24_11_a_24 & f_s_dadda_pg_rca32_and_24_11_b_11;
  assign f_s_dadda_pg_rca32_and_23_12_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_23_12_y0 = f_s_dadda_pg_rca32_and_23_12_a_23 & f_s_dadda_pg_rca32_and_23_12_b_12;
  assign f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_25_10_y0 = f_s_dadda_pg_rca32_and_25_10_y0;
  assign f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_24_11_y0 = f_s_dadda_pg_rca32_and_24_11_y0;
  assign f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_23_12_y0 = f_s_dadda_pg_rca32_and_23_12_y0;
  assign f_s_dadda_pg_rca32_fa410_y0 = f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_25_10_y0 ^ f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_24_11_y0;
  assign f_s_dadda_pg_rca32_fa410_y1 = f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_25_10_y0 & f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_24_11_y0;
  assign f_s_dadda_pg_rca32_fa410_y2 = f_s_dadda_pg_rca32_fa410_y0 ^ f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_23_12_y0;
  assign f_s_dadda_pg_rca32_fa410_y3 = f_s_dadda_pg_rca32_fa410_y0 & f_s_dadda_pg_rca32_fa410_f_s_dadda_pg_rca32_and_23_12_y0;
  assign f_s_dadda_pg_rca32_fa410_y4 = f_s_dadda_pg_rca32_fa410_y1 | f_s_dadda_pg_rca32_fa410_y3;
  assign f_s_dadda_pg_rca32_and_22_13_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_22_13_y0 = f_s_dadda_pg_rca32_and_22_13_a_22 & f_s_dadda_pg_rca32_and_22_13_b_13;
  assign f_s_dadda_pg_rca32_and_21_14_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_21_14_y0 = f_s_dadda_pg_rca32_and_21_14_a_21 & f_s_dadda_pg_rca32_and_21_14_b_14;
  assign f_s_dadda_pg_rca32_and_20_15_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_20_15_y0 = f_s_dadda_pg_rca32_and_20_15_a_20 & f_s_dadda_pg_rca32_and_20_15_b_15;
  assign f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_22_13_y0 = f_s_dadda_pg_rca32_and_22_13_y0;
  assign f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_21_14_y0 = f_s_dadda_pg_rca32_and_21_14_y0;
  assign f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_20_15_y0 = f_s_dadda_pg_rca32_and_20_15_y0;
  assign f_s_dadda_pg_rca32_fa411_y0 = f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_22_13_y0 ^ f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_21_14_y0;
  assign f_s_dadda_pg_rca32_fa411_y1 = f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_22_13_y0 & f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_21_14_y0;
  assign f_s_dadda_pg_rca32_fa411_y2 = f_s_dadda_pg_rca32_fa411_y0 ^ f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_20_15_y0;
  assign f_s_dadda_pg_rca32_fa411_y3 = f_s_dadda_pg_rca32_fa411_y0 & f_s_dadda_pg_rca32_fa411_f_s_dadda_pg_rca32_and_20_15_y0;
  assign f_s_dadda_pg_rca32_fa411_y4 = f_s_dadda_pg_rca32_fa411_y1 | f_s_dadda_pg_rca32_fa411_y3;
  assign f_s_dadda_pg_rca32_and_19_16_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_19_16_y0 = f_s_dadda_pg_rca32_and_19_16_a_19 & f_s_dadda_pg_rca32_and_19_16_b_16;
  assign f_s_dadda_pg_rca32_and_18_17_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_18_17_y0 = f_s_dadda_pg_rca32_and_18_17_a_18 & f_s_dadda_pg_rca32_and_18_17_b_17;
  assign f_s_dadda_pg_rca32_and_17_18_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_17_18_y0 = f_s_dadda_pg_rca32_and_17_18_a_17 & f_s_dadda_pg_rca32_and_17_18_b_18;
  assign f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_19_16_y0 = f_s_dadda_pg_rca32_and_19_16_y0;
  assign f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_18_17_y0 = f_s_dadda_pg_rca32_and_18_17_y0;
  assign f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_17_18_y0 = f_s_dadda_pg_rca32_and_17_18_y0;
  assign f_s_dadda_pg_rca32_fa412_y0 = f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_19_16_y0 ^ f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_18_17_y0;
  assign f_s_dadda_pg_rca32_fa412_y1 = f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_19_16_y0 & f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_18_17_y0;
  assign f_s_dadda_pg_rca32_fa412_y2 = f_s_dadda_pg_rca32_fa412_y0 ^ f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_17_18_y0;
  assign f_s_dadda_pg_rca32_fa412_y3 = f_s_dadda_pg_rca32_fa412_y0 & f_s_dadda_pg_rca32_fa412_f_s_dadda_pg_rca32_and_17_18_y0;
  assign f_s_dadda_pg_rca32_fa412_y4 = f_s_dadda_pg_rca32_fa412_y1 | f_s_dadda_pg_rca32_fa412_y3;
  assign f_s_dadda_pg_rca32_and_16_19_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_16_19_y0 = f_s_dadda_pg_rca32_and_16_19_a_16 & f_s_dadda_pg_rca32_and_16_19_b_19;
  assign f_s_dadda_pg_rca32_and_15_20_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_15_20_y0 = f_s_dadda_pg_rca32_and_15_20_a_15 & f_s_dadda_pg_rca32_and_15_20_b_20;
  assign f_s_dadda_pg_rca32_and_14_21_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_14_21_y0 = f_s_dadda_pg_rca32_and_14_21_a_14 & f_s_dadda_pg_rca32_and_14_21_b_21;
  assign f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_16_19_y0 = f_s_dadda_pg_rca32_and_16_19_y0;
  assign f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_15_20_y0 = f_s_dadda_pg_rca32_and_15_20_y0;
  assign f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_14_21_y0 = f_s_dadda_pg_rca32_and_14_21_y0;
  assign f_s_dadda_pg_rca32_fa413_y0 = f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_16_19_y0 ^ f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_15_20_y0;
  assign f_s_dadda_pg_rca32_fa413_y1 = f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_16_19_y0 & f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_15_20_y0;
  assign f_s_dadda_pg_rca32_fa413_y2 = f_s_dadda_pg_rca32_fa413_y0 ^ f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_14_21_y0;
  assign f_s_dadda_pg_rca32_fa413_y3 = f_s_dadda_pg_rca32_fa413_y0 & f_s_dadda_pg_rca32_fa413_f_s_dadda_pg_rca32_and_14_21_y0;
  assign f_s_dadda_pg_rca32_fa413_y4 = f_s_dadda_pg_rca32_fa413_y1 | f_s_dadda_pg_rca32_fa413_y3;
  assign f_s_dadda_pg_rca32_and_13_22_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_13_22_y0 = f_s_dadda_pg_rca32_and_13_22_a_13 & f_s_dadda_pg_rca32_and_13_22_b_22;
  assign f_s_dadda_pg_rca32_and_12_23_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_12_23_y0 = f_s_dadda_pg_rca32_and_12_23_a_12 & f_s_dadda_pg_rca32_and_12_23_b_23;
  assign f_s_dadda_pg_rca32_and_11_24_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_11_24_y0 = f_s_dadda_pg_rca32_and_11_24_a_11 & f_s_dadda_pg_rca32_and_11_24_b_24;
  assign f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_13_22_y0 = f_s_dadda_pg_rca32_and_13_22_y0;
  assign f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_12_23_y0 = f_s_dadda_pg_rca32_and_12_23_y0;
  assign f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_11_24_y0 = f_s_dadda_pg_rca32_and_11_24_y0;
  assign f_s_dadda_pg_rca32_fa414_y0 = f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_13_22_y0 ^ f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_12_23_y0;
  assign f_s_dadda_pg_rca32_fa414_y1 = f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_13_22_y0 & f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_12_23_y0;
  assign f_s_dadda_pg_rca32_fa414_y2 = f_s_dadda_pg_rca32_fa414_y0 ^ f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_11_24_y0;
  assign f_s_dadda_pg_rca32_fa414_y3 = f_s_dadda_pg_rca32_fa414_y0 & f_s_dadda_pg_rca32_fa414_f_s_dadda_pg_rca32_and_11_24_y0;
  assign f_s_dadda_pg_rca32_fa414_y4 = f_s_dadda_pg_rca32_fa414_y1 | f_s_dadda_pg_rca32_fa414_y3;
  assign f_s_dadda_pg_rca32_and_10_25_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_10_25_y0 = f_s_dadda_pg_rca32_and_10_25_a_10 & f_s_dadda_pg_rca32_and_10_25_b_25;
  assign f_s_dadda_pg_rca32_and_9_26_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_9_26_y0 = f_s_dadda_pg_rca32_and_9_26_a_9 & f_s_dadda_pg_rca32_and_9_26_b_26;
  assign f_s_dadda_pg_rca32_and_8_27_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_8_27_y0 = f_s_dadda_pg_rca32_and_8_27_a_8 & f_s_dadda_pg_rca32_and_8_27_b_27;
  assign f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_10_25_y0 = f_s_dadda_pg_rca32_and_10_25_y0;
  assign f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_9_26_y0 = f_s_dadda_pg_rca32_and_9_26_y0;
  assign f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_8_27_y0 = f_s_dadda_pg_rca32_and_8_27_y0;
  assign f_s_dadda_pg_rca32_fa415_y0 = f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_10_25_y0 ^ f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_9_26_y0;
  assign f_s_dadda_pg_rca32_fa415_y1 = f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_10_25_y0 & f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_9_26_y0;
  assign f_s_dadda_pg_rca32_fa415_y2 = f_s_dadda_pg_rca32_fa415_y0 ^ f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_8_27_y0;
  assign f_s_dadda_pg_rca32_fa415_y3 = f_s_dadda_pg_rca32_fa415_y0 & f_s_dadda_pg_rca32_fa415_f_s_dadda_pg_rca32_and_8_27_y0;
  assign f_s_dadda_pg_rca32_fa415_y4 = f_s_dadda_pg_rca32_fa415_y1 | f_s_dadda_pg_rca32_fa415_y3;
  assign f_s_dadda_pg_rca32_and_7_28_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_7_28_y0 = f_s_dadda_pg_rca32_and_7_28_a_7 & f_s_dadda_pg_rca32_and_7_28_b_28;
  assign f_s_dadda_pg_rca32_and_6_29_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_6_29_y0 = f_s_dadda_pg_rca32_and_6_29_a_6 & f_s_dadda_pg_rca32_and_6_29_b_29;
  assign f_s_dadda_pg_rca32_and_5_30_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_5_30_y0 = f_s_dadda_pg_rca32_and_5_30_a_5 & f_s_dadda_pg_rca32_and_5_30_b_30;
  assign f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_7_28_y0 = f_s_dadda_pg_rca32_and_7_28_y0;
  assign f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_6_29_y0 = f_s_dadda_pg_rca32_and_6_29_y0;
  assign f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_5_30_y0 = f_s_dadda_pg_rca32_and_5_30_y0;
  assign f_s_dadda_pg_rca32_fa416_y0 = f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_7_28_y0 ^ f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_6_29_y0;
  assign f_s_dadda_pg_rca32_fa416_y1 = f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_7_28_y0 & f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_6_29_y0;
  assign f_s_dadda_pg_rca32_fa416_y2 = f_s_dadda_pg_rca32_fa416_y0 ^ f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_5_30_y0;
  assign f_s_dadda_pg_rca32_fa416_y3 = f_s_dadda_pg_rca32_fa416_y0 & f_s_dadda_pg_rca32_fa416_f_s_dadda_pg_rca32_and_5_30_y0;
  assign f_s_dadda_pg_rca32_fa416_y4 = f_s_dadda_pg_rca32_fa416_y1 | f_s_dadda_pg_rca32_fa416_y3;
  assign f_s_dadda_pg_rca32_nand_4_31_a_4 = a_4;
  assign f_s_dadda_pg_rca32_nand_4_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_4_31_y0 = ~(f_s_dadda_pg_rca32_nand_4_31_a_4 & f_s_dadda_pg_rca32_nand_4_31_b_31);
  assign f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_nand_4_31_y0 = f_s_dadda_pg_rca32_nand_4_31_y0;
  assign f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_fa15_y2 = f_s_dadda_pg_rca32_fa15_y2;
  assign f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_fa401_y2 = f_s_dadda_pg_rca32_fa401_y2;
  assign f_s_dadda_pg_rca32_fa417_y0 = f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_nand_4_31_y0 ^ f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_fa15_y2;
  assign f_s_dadda_pg_rca32_fa417_y1 = f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_nand_4_31_y0 & f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_fa15_y2;
  assign f_s_dadda_pg_rca32_fa417_y2 = f_s_dadda_pg_rca32_fa417_y0 ^ f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_fa401_y2;
  assign f_s_dadda_pg_rca32_fa417_y3 = f_s_dadda_pg_rca32_fa417_y0 & f_s_dadda_pg_rca32_fa417_f_s_dadda_pg_rca32_fa401_y2;
  assign f_s_dadda_pg_rca32_fa417_y4 = f_s_dadda_pg_rca32_fa417_y1 | f_s_dadda_pg_rca32_fa417_y3;
  assign f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa402_y2 = f_s_dadda_pg_rca32_fa402_y2;
  assign f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa403_y2 = f_s_dadda_pg_rca32_fa403_y2;
  assign f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa404_y2 = f_s_dadda_pg_rca32_fa404_y2;
  assign f_s_dadda_pg_rca32_fa418_y0 = f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa402_y2 ^ f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa403_y2;
  assign f_s_dadda_pg_rca32_fa418_y1 = f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa402_y2 & f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa403_y2;
  assign f_s_dadda_pg_rca32_fa418_y2 = f_s_dadda_pg_rca32_fa418_y0 ^ f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa404_y2;
  assign f_s_dadda_pg_rca32_fa418_y3 = f_s_dadda_pg_rca32_fa418_y0 & f_s_dadda_pg_rca32_fa418_f_s_dadda_pg_rca32_fa404_y2;
  assign f_s_dadda_pg_rca32_fa418_y4 = f_s_dadda_pg_rca32_fa418_y1 | f_s_dadda_pg_rca32_fa418_y3;
  assign f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa405_y2 = f_s_dadda_pg_rca32_fa405_y2;
  assign f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa406_y2 = f_s_dadda_pg_rca32_fa406_y2;
  assign f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa407_y2 = f_s_dadda_pg_rca32_fa407_y2;
  assign f_s_dadda_pg_rca32_fa419_y0 = f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa405_y2 ^ f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa406_y2;
  assign f_s_dadda_pg_rca32_fa419_y1 = f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa405_y2 & f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa406_y2;
  assign f_s_dadda_pg_rca32_fa419_y2 = f_s_dadda_pg_rca32_fa419_y0 ^ f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa407_y2;
  assign f_s_dadda_pg_rca32_fa419_y3 = f_s_dadda_pg_rca32_fa419_y0 & f_s_dadda_pg_rca32_fa419_f_s_dadda_pg_rca32_fa407_y2;
  assign f_s_dadda_pg_rca32_fa419_y4 = f_s_dadda_pg_rca32_fa419_y1 | f_s_dadda_pg_rca32_fa419_y3;
  assign f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa408_y2 = f_s_dadda_pg_rca32_fa408_y2;
  assign f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa409_y2 = f_s_dadda_pg_rca32_fa409_y2;
  assign f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa410_y2 = f_s_dadda_pg_rca32_fa410_y2;
  assign f_s_dadda_pg_rca32_fa420_y0 = f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa408_y2 ^ f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa409_y2;
  assign f_s_dadda_pg_rca32_fa420_y1 = f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa408_y2 & f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa409_y2;
  assign f_s_dadda_pg_rca32_fa420_y2 = f_s_dadda_pg_rca32_fa420_y0 ^ f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa410_y2;
  assign f_s_dadda_pg_rca32_fa420_y3 = f_s_dadda_pg_rca32_fa420_y0 & f_s_dadda_pg_rca32_fa420_f_s_dadda_pg_rca32_fa410_y2;
  assign f_s_dadda_pg_rca32_fa420_y4 = f_s_dadda_pg_rca32_fa420_y1 | f_s_dadda_pg_rca32_fa420_y3;
  assign f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa411_y2 = f_s_dadda_pg_rca32_fa411_y2;
  assign f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa412_y2 = f_s_dadda_pg_rca32_fa412_y2;
  assign f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa413_y2 = f_s_dadda_pg_rca32_fa413_y2;
  assign f_s_dadda_pg_rca32_fa421_y0 = f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa411_y2 ^ f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa412_y2;
  assign f_s_dadda_pg_rca32_fa421_y1 = f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa411_y2 & f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa412_y2;
  assign f_s_dadda_pg_rca32_fa421_y2 = f_s_dadda_pg_rca32_fa421_y0 ^ f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa413_y2;
  assign f_s_dadda_pg_rca32_fa421_y3 = f_s_dadda_pg_rca32_fa421_y0 & f_s_dadda_pg_rca32_fa421_f_s_dadda_pg_rca32_fa413_y2;
  assign f_s_dadda_pg_rca32_fa421_y4 = f_s_dadda_pg_rca32_fa421_y1 | f_s_dadda_pg_rca32_fa421_y3;
  assign f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa414_y2 = f_s_dadda_pg_rca32_fa414_y2;
  assign f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa415_y2 = f_s_dadda_pg_rca32_fa415_y2;
  assign f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa416_y2 = f_s_dadda_pg_rca32_fa416_y2;
  assign f_s_dadda_pg_rca32_fa422_y0 = f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa414_y2 ^ f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa415_y2;
  assign f_s_dadda_pg_rca32_fa422_y1 = f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa414_y2 & f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa415_y2;
  assign f_s_dadda_pg_rca32_fa422_y2 = f_s_dadda_pg_rca32_fa422_y0 ^ f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa416_y2;
  assign f_s_dadda_pg_rca32_fa422_y3 = f_s_dadda_pg_rca32_fa422_y0 & f_s_dadda_pg_rca32_fa422_f_s_dadda_pg_rca32_fa416_y2;
  assign f_s_dadda_pg_rca32_fa422_y4 = f_s_dadda_pg_rca32_fa422_y1 | f_s_dadda_pg_rca32_fa422_y3;
  assign f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa422_y4 = f_s_dadda_pg_rca32_fa422_y4;
  assign f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa421_y4 = f_s_dadda_pg_rca32_fa421_y4;
  assign f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa420_y4 = f_s_dadda_pg_rca32_fa420_y4;
  assign f_s_dadda_pg_rca32_fa423_y0 = f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa422_y4 ^ f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa421_y4;
  assign f_s_dadda_pg_rca32_fa423_y1 = f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa422_y4 & f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa421_y4;
  assign f_s_dadda_pg_rca32_fa423_y2 = f_s_dadda_pg_rca32_fa423_y0 ^ f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa420_y4;
  assign f_s_dadda_pg_rca32_fa423_y3 = f_s_dadda_pg_rca32_fa423_y0 & f_s_dadda_pg_rca32_fa423_f_s_dadda_pg_rca32_fa420_y4;
  assign f_s_dadda_pg_rca32_fa423_y4 = f_s_dadda_pg_rca32_fa423_y1 | f_s_dadda_pg_rca32_fa423_y3;
  assign f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa419_y4 = f_s_dadda_pg_rca32_fa419_y4;
  assign f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa418_y4 = f_s_dadda_pg_rca32_fa418_y4;
  assign f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa417_y4 = f_s_dadda_pg_rca32_fa417_y4;
  assign f_s_dadda_pg_rca32_fa424_y0 = f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa419_y4 ^ f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa418_y4;
  assign f_s_dadda_pg_rca32_fa424_y1 = f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa419_y4 & f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa418_y4;
  assign f_s_dadda_pg_rca32_fa424_y2 = f_s_dadda_pg_rca32_fa424_y0 ^ f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa417_y4;
  assign f_s_dadda_pg_rca32_fa424_y3 = f_s_dadda_pg_rca32_fa424_y0 & f_s_dadda_pg_rca32_fa424_f_s_dadda_pg_rca32_fa417_y4;
  assign f_s_dadda_pg_rca32_fa424_y4 = f_s_dadda_pg_rca32_fa424_y1 | f_s_dadda_pg_rca32_fa424_y3;
  assign f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa416_y4 = f_s_dadda_pg_rca32_fa416_y4;
  assign f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa415_y4 = f_s_dadda_pg_rca32_fa415_y4;
  assign f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa414_y4 = f_s_dadda_pg_rca32_fa414_y4;
  assign f_s_dadda_pg_rca32_fa425_y0 = f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa416_y4 ^ f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa415_y4;
  assign f_s_dadda_pg_rca32_fa425_y1 = f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa416_y4 & f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa415_y4;
  assign f_s_dadda_pg_rca32_fa425_y2 = f_s_dadda_pg_rca32_fa425_y0 ^ f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa414_y4;
  assign f_s_dadda_pg_rca32_fa425_y3 = f_s_dadda_pg_rca32_fa425_y0 & f_s_dadda_pg_rca32_fa425_f_s_dadda_pg_rca32_fa414_y4;
  assign f_s_dadda_pg_rca32_fa425_y4 = f_s_dadda_pg_rca32_fa425_y1 | f_s_dadda_pg_rca32_fa425_y3;
  assign f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa413_y4 = f_s_dadda_pg_rca32_fa413_y4;
  assign f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa412_y4 = f_s_dadda_pg_rca32_fa412_y4;
  assign f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa411_y4 = f_s_dadda_pg_rca32_fa411_y4;
  assign f_s_dadda_pg_rca32_fa426_y0 = f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa413_y4 ^ f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa412_y4;
  assign f_s_dadda_pg_rca32_fa426_y1 = f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa413_y4 & f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa412_y4;
  assign f_s_dadda_pg_rca32_fa426_y2 = f_s_dadda_pg_rca32_fa426_y0 ^ f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa411_y4;
  assign f_s_dadda_pg_rca32_fa426_y3 = f_s_dadda_pg_rca32_fa426_y0 & f_s_dadda_pg_rca32_fa426_f_s_dadda_pg_rca32_fa411_y4;
  assign f_s_dadda_pg_rca32_fa426_y4 = f_s_dadda_pg_rca32_fa426_y1 | f_s_dadda_pg_rca32_fa426_y3;
  assign f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa410_y4 = f_s_dadda_pg_rca32_fa410_y4;
  assign f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa409_y4 = f_s_dadda_pg_rca32_fa409_y4;
  assign f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa408_y4 = f_s_dadda_pg_rca32_fa408_y4;
  assign f_s_dadda_pg_rca32_fa427_y0 = f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa410_y4 ^ f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa409_y4;
  assign f_s_dadda_pg_rca32_fa427_y1 = f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa410_y4 & f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa409_y4;
  assign f_s_dadda_pg_rca32_fa427_y2 = f_s_dadda_pg_rca32_fa427_y0 ^ f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa408_y4;
  assign f_s_dadda_pg_rca32_fa427_y3 = f_s_dadda_pg_rca32_fa427_y0 & f_s_dadda_pg_rca32_fa427_f_s_dadda_pg_rca32_fa408_y4;
  assign f_s_dadda_pg_rca32_fa427_y4 = f_s_dadda_pg_rca32_fa427_y1 | f_s_dadda_pg_rca32_fa427_y3;
  assign f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa407_y4 = f_s_dadda_pg_rca32_fa407_y4;
  assign f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa406_y4 = f_s_dadda_pg_rca32_fa406_y4;
  assign f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa405_y4 = f_s_dadda_pg_rca32_fa405_y4;
  assign f_s_dadda_pg_rca32_fa428_y0 = f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa407_y4 ^ f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa406_y4;
  assign f_s_dadda_pg_rca32_fa428_y1 = f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa407_y4 & f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa406_y4;
  assign f_s_dadda_pg_rca32_fa428_y2 = f_s_dadda_pg_rca32_fa428_y0 ^ f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa405_y4;
  assign f_s_dadda_pg_rca32_fa428_y3 = f_s_dadda_pg_rca32_fa428_y0 & f_s_dadda_pg_rca32_fa428_f_s_dadda_pg_rca32_fa405_y4;
  assign f_s_dadda_pg_rca32_fa428_y4 = f_s_dadda_pg_rca32_fa428_y1 | f_s_dadda_pg_rca32_fa428_y3;
  assign f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa404_y4 = f_s_dadda_pg_rca32_fa404_y4;
  assign f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa403_y4 = f_s_dadda_pg_rca32_fa403_y4;
  assign f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa402_y4 = f_s_dadda_pg_rca32_fa402_y4;
  assign f_s_dadda_pg_rca32_fa429_y0 = f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa404_y4 ^ f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa403_y4;
  assign f_s_dadda_pg_rca32_fa429_y1 = f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa404_y4 & f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa403_y4;
  assign f_s_dadda_pg_rca32_fa429_y2 = f_s_dadda_pg_rca32_fa429_y0 ^ f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa402_y4;
  assign f_s_dadda_pg_rca32_fa429_y3 = f_s_dadda_pg_rca32_fa429_y0 & f_s_dadda_pg_rca32_fa429_f_s_dadda_pg_rca32_fa402_y4;
  assign f_s_dadda_pg_rca32_fa429_y4 = f_s_dadda_pg_rca32_fa429_y1 | f_s_dadda_pg_rca32_fa429_y3;
  assign f_s_dadda_pg_rca32_nand_31_5_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_nand_31_5_y0 = ~(f_s_dadda_pg_rca32_nand_31_5_a_31 & f_s_dadda_pg_rca32_nand_31_5_b_5);
  assign f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_fa401_y4 = f_s_dadda_pg_rca32_fa401_y4;
  assign f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_fa15_y4 = f_s_dadda_pg_rca32_fa15_y4;
  assign f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_nand_31_5_y0 = f_s_dadda_pg_rca32_nand_31_5_y0;
  assign f_s_dadda_pg_rca32_fa430_y0 = f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_fa401_y4 ^ f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_fa15_y4;
  assign f_s_dadda_pg_rca32_fa430_y1 = f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_fa401_y4 & f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_fa15_y4;
  assign f_s_dadda_pg_rca32_fa430_y2 = f_s_dadda_pg_rca32_fa430_y0 ^ f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_nand_31_5_y0;
  assign f_s_dadda_pg_rca32_fa430_y3 = f_s_dadda_pg_rca32_fa430_y0 & f_s_dadda_pg_rca32_fa430_f_s_dadda_pg_rca32_nand_31_5_y0;
  assign f_s_dadda_pg_rca32_fa430_y4 = f_s_dadda_pg_rca32_fa430_y1 | f_s_dadda_pg_rca32_fa430_y3;
  assign f_s_dadda_pg_rca32_and_30_6_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_30_6_y0 = f_s_dadda_pg_rca32_and_30_6_a_30 & f_s_dadda_pg_rca32_and_30_6_b_6;
  assign f_s_dadda_pg_rca32_and_29_7_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_29_7_y0 = f_s_dadda_pg_rca32_and_29_7_a_29 & f_s_dadda_pg_rca32_and_29_7_b_7;
  assign f_s_dadda_pg_rca32_and_28_8_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_28_8_y0 = f_s_dadda_pg_rca32_and_28_8_a_28 & f_s_dadda_pg_rca32_and_28_8_b_8;
  assign f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_30_6_y0 = f_s_dadda_pg_rca32_and_30_6_y0;
  assign f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_29_7_y0 = f_s_dadda_pg_rca32_and_29_7_y0;
  assign f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_28_8_y0 = f_s_dadda_pg_rca32_and_28_8_y0;
  assign f_s_dadda_pg_rca32_fa431_y0 = f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_30_6_y0 ^ f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_29_7_y0;
  assign f_s_dadda_pg_rca32_fa431_y1 = f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_30_6_y0 & f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_29_7_y0;
  assign f_s_dadda_pg_rca32_fa431_y2 = f_s_dadda_pg_rca32_fa431_y0 ^ f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_28_8_y0;
  assign f_s_dadda_pg_rca32_fa431_y3 = f_s_dadda_pg_rca32_fa431_y0 & f_s_dadda_pg_rca32_fa431_f_s_dadda_pg_rca32_and_28_8_y0;
  assign f_s_dadda_pg_rca32_fa431_y4 = f_s_dadda_pg_rca32_fa431_y1 | f_s_dadda_pg_rca32_fa431_y3;
  assign f_s_dadda_pg_rca32_and_27_9_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_27_9_y0 = f_s_dadda_pg_rca32_and_27_9_a_27 & f_s_dadda_pg_rca32_and_27_9_b_9;
  assign f_s_dadda_pg_rca32_and_26_10_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_26_10_y0 = f_s_dadda_pg_rca32_and_26_10_a_26 & f_s_dadda_pg_rca32_and_26_10_b_10;
  assign f_s_dadda_pg_rca32_and_25_11_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_25_11_y0 = f_s_dadda_pg_rca32_and_25_11_a_25 & f_s_dadda_pg_rca32_and_25_11_b_11;
  assign f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_27_9_y0 = f_s_dadda_pg_rca32_and_27_9_y0;
  assign f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_26_10_y0 = f_s_dadda_pg_rca32_and_26_10_y0;
  assign f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_25_11_y0 = f_s_dadda_pg_rca32_and_25_11_y0;
  assign f_s_dadda_pg_rca32_fa432_y0 = f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_27_9_y0 ^ f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_26_10_y0;
  assign f_s_dadda_pg_rca32_fa432_y1 = f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_27_9_y0 & f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_26_10_y0;
  assign f_s_dadda_pg_rca32_fa432_y2 = f_s_dadda_pg_rca32_fa432_y0 ^ f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_25_11_y0;
  assign f_s_dadda_pg_rca32_fa432_y3 = f_s_dadda_pg_rca32_fa432_y0 & f_s_dadda_pg_rca32_fa432_f_s_dadda_pg_rca32_and_25_11_y0;
  assign f_s_dadda_pg_rca32_fa432_y4 = f_s_dadda_pg_rca32_fa432_y1 | f_s_dadda_pg_rca32_fa432_y3;
  assign f_s_dadda_pg_rca32_and_24_12_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_24_12_y0 = f_s_dadda_pg_rca32_and_24_12_a_24 & f_s_dadda_pg_rca32_and_24_12_b_12;
  assign f_s_dadda_pg_rca32_and_23_13_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_23_13_y0 = f_s_dadda_pg_rca32_and_23_13_a_23 & f_s_dadda_pg_rca32_and_23_13_b_13;
  assign f_s_dadda_pg_rca32_and_22_14_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_22_14_y0 = f_s_dadda_pg_rca32_and_22_14_a_22 & f_s_dadda_pg_rca32_and_22_14_b_14;
  assign f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_24_12_y0 = f_s_dadda_pg_rca32_and_24_12_y0;
  assign f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_23_13_y0 = f_s_dadda_pg_rca32_and_23_13_y0;
  assign f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_22_14_y0 = f_s_dadda_pg_rca32_and_22_14_y0;
  assign f_s_dadda_pg_rca32_fa433_y0 = f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_24_12_y0 ^ f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_23_13_y0;
  assign f_s_dadda_pg_rca32_fa433_y1 = f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_24_12_y0 & f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_23_13_y0;
  assign f_s_dadda_pg_rca32_fa433_y2 = f_s_dadda_pg_rca32_fa433_y0 ^ f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_22_14_y0;
  assign f_s_dadda_pg_rca32_fa433_y3 = f_s_dadda_pg_rca32_fa433_y0 & f_s_dadda_pg_rca32_fa433_f_s_dadda_pg_rca32_and_22_14_y0;
  assign f_s_dadda_pg_rca32_fa433_y4 = f_s_dadda_pg_rca32_fa433_y1 | f_s_dadda_pg_rca32_fa433_y3;
  assign f_s_dadda_pg_rca32_and_21_15_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_21_15_y0 = f_s_dadda_pg_rca32_and_21_15_a_21 & f_s_dadda_pg_rca32_and_21_15_b_15;
  assign f_s_dadda_pg_rca32_and_20_16_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_20_16_y0 = f_s_dadda_pg_rca32_and_20_16_a_20 & f_s_dadda_pg_rca32_and_20_16_b_16;
  assign f_s_dadda_pg_rca32_and_19_17_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_19_17_y0 = f_s_dadda_pg_rca32_and_19_17_a_19 & f_s_dadda_pg_rca32_and_19_17_b_17;
  assign f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_21_15_y0 = f_s_dadda_pg_rca32_and_21_15_y0;
  assign f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_20_16_y0 = f_s_dadda_pg_rca32_and_20_16_y0;
  assign f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_19_17_y0 = f_s_dadda_pg_rca32_and_19_17_y0;
  assign f_s_dadda_pg_rca32_fa434_y0 = f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_21_15_y0 ^ f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_20_16_y0;
  assign f_s_dadda_pg_rca32_fa434_y1 = f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_21_15_y0 & f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_20_16_y0;
  assign f_s_dadda_pg_rca32_fa434_y2 = f_s_dadda_pg_rca32_fa434_y0 ^ f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_19_17_y0;
  assign f_s_dadda_pg_rca32_fa434_y3 = f_s_dadda_pg_rca32_fa434_y0 & f_s_dadda_pg_rca32_fa434_f_s_dadda_pg_rca32_and_19_17_y0;
  assign f_s_dadda_pg_rca32_fa434_y4 = f_s_dadda_pg_rca32_fa434_y1 | f_s_dadda_pg_rca32_fa434_y3;
  assign f_s_dadda_pg_rca32_and_18_18_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_18_18_y0 = f_s_dadda_pg_rca32_and_18_18_a_18 & f_s_dadda_pg_rca32_and_18_18_b_18;
  assign f_s_dadda_pg_rca32_and_17_19_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_17_19_y0 = f_s_dadda_pg_rca32_and_17_19_a_17 & f_s_dadda_pg_rca32_and_17_19_b_19;
  assign f_s_dadda_pg_rca32_and_16_20_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_16_20_y0 = f_s_dadda_pg_rca32_and_16_20_a_16 & f_s_dadda_pg_rca32_and_16_20_b_20;
  assign f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_18_18_y0 = f_s_dadda_pg_rca32_and_18_18_y0;
  assign f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_17_19_y0 = f_s_dadda_pg_rca32_and_17_19_y0;
  assign f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_16_20_y0 = f_s_dadda_pg_rca32_and_16_20_y0;
  assign f_s_dadda_pg_rca32_fa435_y0 = f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_18_18_y0 ^ f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_17_19_y0;
  assign f_s_dadda_pg_rca32_fa435_y1 = f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_18_18_y0 & f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_17_19_y0;
  assign f_s_dadda_pg_rca32_fa435_y2 = f_s_dadda_pg_rca32_fa435_y0 ^ f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_16_20_y0;
  assign f_s_dadda_pg_rca32_fa435_y3 = f_s_dadda_pg_rca32_fa435_y0 & f_s_dadda_pg_rca32_fa435_f_s_dadda_pg_rca32_and_16_20_y0;
  assign f_s_dadda_pg_rca32_fa435_y4 = f_s_dadda_pg_rca32_fa435_y1 | f_s_dadda_pg_rca32_fa435_y3;
  assign f_s_dadda_pg_rca32_and_15_21_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_15_21_y0 = f_s_dadda_pg_rca32_and_15_21_a_15 & f_s_dadda_pg_rca32_and_15_21_b_21;
  assign f_s_dadda_pg_rca32_and_14_22_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_14_22_y0 = f_s_dadda_pg_rca32_and_14_22_a_14 & f_s_dadda_pg_rca32_and_14_22_b_22;
  assign f_s_dadda_pg_rca32_and_13_23_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_13_23_y0 = f_s_dadda_pg_rca32_and_13_23_a_13 & f_s_dadda_pg_rca32_and_13_23_b_23;
  assign f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_15_21_y0 = f_s_dadda_pg_rca32_and_15_21_y0;
  assign f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_14_22_y0 = f_s_dadda_pg_rca32_and_14_22_y0;
  assign f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_13_23_y0 = f_s_dadda_pg_rca32_and_13_23_y0;
  assign f_s_dadda_pg_rca32_fa436_y0 = f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_15_21_y0 ^ f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_14_22_y0;
  assign f_s_dadda_pg_rca32_fa436_y1 = f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_15_21_y0 & f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_14_22_y0;
  assign f_s_dadda_pg_rca32_fa436_y2 = f_s_dadda_pg_rca32_fa436_y0 ^ f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_13_23_y0;
  assign f_s_dadda_pg_rca32_fa436_y3 = f_s_dadda_pg_rca32_fa436_y0 & f_s_dadda_pg_rca32_fa436_f_s_dadda_pg_rca32_and_13_23_y0;
  assign f_s_dadda_pg_rca32_fa436_y4 = f_s_dadda_pg_rca32_fa436_y1 | f_s_dadda_pg_rca32_fa436_y3;
  assign f_s_dadda_pg_rca32_and_12_24_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_12_24_y0 = f_s_dadda_pg_rca32_and_12_24_a_12 & f_s_dadda_pg_rca32_and_12_24_b_24;
  assign f_s_dadda_pg_rca32_and_11_25_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_11_25_y0 = f_s_dadda_pg_rca32_and_11_25_a_11 & f_s_dadda_pg_rca32_and_11_25_b_25;
  assign f_s_dadda_pg_rca32_and_10_26_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_10_26_y0 = f_s_dadda_pg_rca32_and_10_26_a_10 & f_s_dadda_pg_rca32_and_10_26_b_26;
  assign f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_12_24_y0 = f_s_dadda_pg_rca32_and_12_24_y0;
  assign f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_11_25_y0 = f_s_dadda_pg_rca32_and_11_25_y0;
  assign f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_10_26_y0 = f_s_dadda_pg_rca32_and_10_26_y0;
  assign f_s_dadda_pg_rca32_fa437_y0 = f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_12_24_y0 ^ f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_11_25_y0;
  assign f_s_dadda_pg_rca32_fa437_y1 = f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_12_24_y0 & f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_11_25_y0;
  assign f_s_dadda_pg_rca32_fa437_y2 = f_s_dadda_pg_rca32_fa437_y0 ^ f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_10_26_y0;
  assign f_s_dadda_pg_rca32_fa437_y3 = f_s_dadda_pg_rca32_fa437_y0 & f_s_dadda_pg_rca32_fa437_f_s_dadda_pg_rca32_and_10_26_y0;
  assign f_s_dadda_pg_rca32_fa437_y4 = f_s_dadda_pg_rca32_fa437_y1 | f_s_dadda_pg_rca32_fa437_y3;
  assign f_s_dadda_pg_rca32_and_9_27_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_9_27_y0 = f_s_dadda_pg_rca32_and_9_27_a_9 & f_s_dadda_pg_rca32_and_9_27_b_27;
  assign f_s_dadda_pg_rca32_and_8_28_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_8_28_y0 = f_s_dadda_pg_rca32_and_8_28_a_8 & f_s_dadda_pg_rca32_and_8_28_b_28;
  assign f_s_dadda_pg_rca32_and_7_29_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_7_29_y0 = f_s_dadda_pg_rca32_and_7_29_a_7 & f_s_dadda_pg_rca32_and_7_29_b_29;
  assign f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_9_27_y0 = f_s_dadda_pg_rca32_and_9_27_y0;
  assign f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_8_28_y0 = f_s_dadda_pg_rca32_and_8_28_y0;
  assign f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_7_29_y0 = f_s_dadda_pg_rca32_and_7_29_y0;
  assign f_s_dadda_pg_rca32_fa438_y0 = f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_9_27_y0 ^ f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_8_28_y0;
  assign f_s_dadda_pg_rca32_fa438_y1 = f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_9_27_y0 & f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_8_28_y0;
  assign f_s_dadda_pg_rca32_fa438_y2 = f_s_dadda_pg_rca32_fa438_y0 ^ f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_7_29_y0;
  assign f_s_dadda_pg_rca32_fa438_y3 = f_s_dadda_pg_rca32_fa438_y0 & f_s_dadda_pg_rca32_fa438_f_s_dadda_pg_rca32_and_7_29_y0;
  assign f_s_dadda_pg_rca32_fa438_y4 = f_s_dadda_pg_rca32_fa438_y1 | f_s_dadda_pg_rca32_fa438_y3;
  assign f_s_dadda_pg_rca32_and_6_30_a_6 = a_6;
  assign f_s_dadda_pg_rca32_and_6_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_6_30_y0 = f_s_dadda_pg_rca32_and_6_30_a_6 & f_s_dadda_pg_rca32_and_6_30_b_30;
  assign f_s_dadda_pg_rca32_nand_5_31_a_5 = a_5;
  assign f_s_dadda_pg_rca32_nand_5_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_5_31_y0 = ~(f_s_dadda_pg_rca32_nand_5_31_a_5 & f_s_dadda_pg_rca32_nand_5_31_b_31);
  assign f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_and_6_30_y0 = f_s_dadda_pg_rca32_and_6_30_y0;
  assign f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_nand_5_31_y0 = f_s_dadda_pg_rca32_nand_5_31_y0;
  assign f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_fa423_y2 = f_s_dadda_pg_rca32_fa423_y2;
  assign f_s_dadda_pg_rca32_fa439_y0 = f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_and_6_30_y0 ^ f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_nand_5_31_y0;
  assign f_s_dadda_pg_rca32_fa439_y1 = f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_and_6_30_y0 & f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_nand_5_31_y0;
  assign f_s_dadda_pg_rca32_fa439_y2 = f_s_dadda_pg_rca32_fa439_y0 ^ f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_fa423_y2;
  assign f_s_dadda_pg_rca32_fa439_y3 = f_s_dadda_pg_rca32_fa439_y0 & f_s_dadda_pg_rca32_fa439_f_s_dadda_pg_rca32_fa423_y2;
  assign f_s_dadda_pg_rca32_fa439_y4 = f_s_dadda_pg_rca32_fa439_y1 | f_s_dadda_pg_rca32_fa439_y3;
  assign f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa424_y2 = f_s_dadda_pg_rca32_fa424_y2;
  assign f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa425_y2 = f_s_dadda_pg_rca32_fa425_y2;
  assign f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa426_y2 = f_s_dadda_pg_rca32_fa426_y2;
  assign f_s_dadda_pg_rca32_fa440_y0 = f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa424_y2 ^ f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa425_y2;
  assign f_s_dadda_pg_rca32_fa440_y1 = f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa424_y2 & f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa425_y2;
  assign f_s_dadda_pg_rca32_fa440_y2 = f_s_dadda_pg_rca32_fa440_y0 ^ f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa426_y2;
  assign f_s_dadda_pg_rca32_fa440_y3 = f_s_dadda_pg_rca32_fa440_y0 & f_s_dadda_pg_rca32_fa440_f_s_dadda_pg_rca32_fa426_y2;
  assign f_s_dadda_pg_rca32_fa440_y4 = f_s_dadda_pg_rca32_fa440_y1 | f_s_dadda_pg_rca32_fa440_y3;
  assign f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa427_y2 = f_s_dadda_pg_rca32_fa427_y2;
  assign f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa428_y2 = f_s_dadda_pg_rca32_fa428_y2;
  assign f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa429_y2 = f_s_dadda_pg_rca32_fa429_y2;
  assign f_s_dadda_pg_rca32_fa441_y0 = f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa427_y2 ^ f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa428_y2;
  assign f_s_dadda_pg_rca32_fa441_y1 = f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa427_y2 & f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa428_y2;
  assign f_s_dadda_pg_rca32_fa441_y2 = f_s_dadda_pg_rca32_fa441_y0 ^ f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa429_y2;
  assign f_s_dadda_pg_rca32_fa441_y3 = f_s_dadda_pg_rca32_fa441_y0 & f_s_dadda_pg_rca32_fa441_f_s_dadda_pg_rca32_fa429_y2;
  assign f_s_dadda_pg_rca32_fa441_y4 = f_s_dadda_pg_rca32_fa441_y1 | f_s_dadda_pg_rca32_fa441_y3;
  assign f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa430_y2 = f_s_dadda_pg_rca32_fa430_y2;
  assign f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa431_y2 = f_s_dadda_pg_rca32_fa431_y2;
  assign f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa432_y2 = f_s_dadda_pg_rca32_fa432_y2;
  assign f_s_dadda_pg_rca32_fa442_y0 = f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa430_y2 ^ f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa431_y2;
  assign f_s_dadda_pg_rca32_fa442_y1 = f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa430_y2 & f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa431_y2;
  assign f_s_dadda_pg_rca32_fa442_y2 = f_s_dadda_pg_rca32_fa442_y0 ^ f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa432_y2;
  assign f_s_dadda_pg_rca32_fa442_y3 = f_s_dadda_pg_rca32_fa442_y0 & f_s_dadda_pg_rca32_fa442_f_s_dadda_pg_rca32_fa432_y2;
  assign f_s_dadda_pg_rca32_fa442_y4 = f_s_dadda_pg_rca32_fa442_y1 | f_s_dadda_pg_rca32_fa442_y3;
  assign f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa433_y2 = f_s_dadda_pg_rca32_fa433_y2;
  assign f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa434_y2 = f_s_dadda_pg_rca32_fa434_y2;
  assign f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa435_y2 = f_s_dadda_pg_rca32_fa435_y2;
  assign f_s_dadda_pg_rca32_fa443_y0 = f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa433_y2 ^ f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa434_y2;
  assign f_s_dadda_pg_rca32_fa443_y1 = f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa433_y2 & f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa434_y2;
  assign f_s_dadda_pg_rca32_fa443_y2 = f_s_dadda_pg_rca32_fa443_y0 ^ f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa435_y2;
  assign f_s_dadda_pg_rca32_fa443_y3 = f_s_dadda_pg_rca32_fa443_y0 & f_s_dadda_pg_rca32_fa443_f_s_dadda_pg_rca32_fa435_y2;
  assign f_s_dadda_pg_rca32_fa443_y4 = f_s_dadda_pg_rca32_fa443_y1 | f_s_dadda_pg_rca32_fa443_y3;
  assign f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa436_y2 = f_s_dadda_pg_rca32_fa436_y2;
  assign f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa437_y2 = f_s_dadda_pg_rca32_fa437_y2;
  assign f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa438_y2 = f_s_dadda_pg_rca32_fa438_y2;
  assign f_s_dadda_pg_rca32_fa444_y0 = f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa436_y2 ^ f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa437_y2;
  assign f_s_dadda_pg_rca32_fa444_y1 = f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa436_y2 & f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa437_y2;
  assign f_s_dadda_pg_rca32_fa444_y2 = f_s_dadda_pg_rca32_fa444_y0 ^ f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa438_y2;
  assign f_s_dadda_pg_rca32_fa444_y3 = f_s_dadda_pg_rca32_fa444_y0 & f_s_dadda_pg_rca32_fa444_f_s_dadda_pg_rca32_fa438_y2;
  assign f_s_dadda_pg_rca32_fa444_y4 = f_s_dadda_pg_rca32_fa444_y1 | f_s_dadda_pg_rca32_fa444_y3;
  assign f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa444_y4 = f_s_dadda_pg_rca32_fa444_y4;
  assign f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa443_y4 = f_s_dadda_pg_rca32_fa443_y4;
  assign f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa442_y4 = f_s_dadda_pg_rca32_fa442_y4;
  assign f_s_dadda_pg_rca32_fa445_y0 = f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa444_y4 ^ f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa443_y4;
  assign f_s_dadda_pg_rca32_fa445_y1 = f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa444_y4 & f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa443_y4;
  assign f_s_dadda_pg_rca32_fa445_y2 = f_s_dadda_pg_rca32_fa445_y0 ^ f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa442_y4;
  assign f_s_dadda_pg_rca32_fa445_y3 = f_s_dadda_pg_rca32_fa445_y0 & f_s_dadda_pg_rca32_fa445_f_s_dadda_pg_rca32_fa442_y4;
  assign f_s_dadda_pg_rca32_fa445_y4 = f_s_dadda_pg_rca32_fa445_y1 | f_s_dadda_pg_rca32_fa445_y3;
  assign f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa441_y4 = f_s_dadda_pg_rca32_fa441_y4;
  assign f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa440_y4 = f_s_dadda_pg_rca32_fa440_y4;
  assign f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa439_y4 = f_s_dadda_pg_rca32_fa439_y4;
  assign f_s_dadda_pg_rca32_fa446_y0 = f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa441_y4 ^ f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa440_y4;
  assign f_s_dadda_pg_rca32_fa446_y1 = f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa441_y4 & f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa440_y4;
  assign f_s_dadda_pg_rca32_fa446_y2 = f_s_dadda_pg_rca32_fa446_y0 ^ f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa439_y4;
  assign f_s_dadda_pg_rca32_fa446_y3 = f_s_dadda_pg_rca32_fa446_y0 & f_s_dadda_pg_rca32_fa446_f_s_dadda_pg_rca32_fa439_y4;
  assign f_s_dadda_pg_rca32_fa446_y4 = f_s_dadda_pg_rca32_fa446_y1 | f_s_dadda_pg_rca32_fa446_y3;
  assign f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa438_y4 = f_s_dadda_pg_rca32_fa438_y4;
  assign f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa437_y4 = f_s_dadda_pg_rca32_fa437_y4;
  assign f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa436_y4 = f_s_dadda_pg_rca32_fa436_y4;
  assign f_s_dadda_pg_rca32_fa447_y0 = f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa438_y4 ^ f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa437_y4;
  assign f_s_dadda_pg_rca32_fa447_y1 = f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa438_y4 & f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa437_y4;
  assign f_s_dadda_pg_rca32_fa447_y2 = f_s_dadda_pg_rca32_fa447_y0 ^ f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa436_y4;
  assign f_s_dadda_pg_rca32_fa447_y3 = f_s_dadda_pg_rca32_fa447_y0 & f_s_dadda_pg_rca32_fa447_f_s_dadda_pg_rca32_fa436_y4;
  assign f_s_dadda_pg_rca32_fa447_y4 = f_s_dadda_pg_rca32_fa447_y1 | f_s_dadda_pg_rca32_fa447_y3;
  assign f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa435_y4 = f_s_dadda_pg_rca32_fa435_y4;
  assign f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa434_y4 = f_s_dadda_pg_rca32_fa434_y4;
  assign f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa433_y4 = f_s_dadda_pg_rca32_fa433_y4;
  assign f_s_dadda_pg_rca32_fa448_y0 = f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa435_y4 ^ f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa434_y4;
  assign f_s_dadda_pg_rca32_fa448_y1 = f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa435_y4 & f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa434_y4;
  assign f_s_dadda_pg_rca32_fa448_y2 = f_s_dadda_pg_rca32_fa448_y0 ^ f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa433_y4;
  assign f_s_dadda_pg_rca32_fa448_y3 = f_s_dadda_pg_rca32_fa448_y0 & f_s_dadda_pg_rca32_fa448_f_s_dadda_pg_rca32_fa433_y4;
  assign f_s_dadda_pg_rca32_fa448_y4 = f_s_dadda_pg_rca32_fa448_y1 | f_s_dadda_pg_rca32_fa448_y3;
  assign f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa432_y4 = f_s_dadda_pg_rca32_fa432_y4;
  assign f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa431_y4 = f_s_dadda_pg_rca32_fa431_y4;
  assign f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa430_y4 = f_s_dadda_pg_rca32_fa430_y4;
  assign f_s_dadda_pg_rca32_fa449_y0 = f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa432_y4 ^ f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa431_y4;
  assign f_s_dadda_pg_rca32_fa449_y1 = f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa432_y4 & f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa431_y4;
  assign f_s_dadda_pg_rca32_fa449_y2 = f_s_dadda_pg_rca32_fa449_y0 ^ f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa430_y4;
  assign f_s_dadda_pg_rca32_fa449_y3 = f_s_dadda_pg_rca32_fa449_y0 & f_s_dadda_pg_rca32_fa449_f_s_dadda_pg_rca32_fa430_y4;
  assign f_s_dadda_pg_rca32_fa449_y4 = f_s_dadda_pg_rca32_fa449_y1 | f_s_dadda_pg_rca32_fa449_y3;
  assign f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa429_y4 = f_s_dadda_pg_rca32_fa429_y4;
  assign f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa428_y4 = f_s_dadda_pg_rca32_fa428_y4;
  assign f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa427_y4 = f_s_dadda_pg_rca32_fa427_y4;
  assign f_s_dadda_pg_rca32_fa450_y0 = f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa429_y4 ^ f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa428_y4;
  assign f_s_dadda_pg_rca32_fa450_y1 = f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa429_y4 & f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa428_y4;
  assign f_s_dadda_pg_rca32_fa450_y2 = f_s_dadda_pg_rca32_fa450_y0 ^ f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa427_y4;
  assign f_s_dadda_pg_rca32_fa450_y3 = f_s_dadda_pg_rca32_fa450_y0 & f_s_dadda_pg_rca32_fa450_f_s_dadda_pg_rca32_fa427_y4;
  assign f_s_dadda_pg_rca32_fa450_y4 = f_s_dadda_pg_rca32_fa450_y1 | f_s_dadda_pg_rca32_fa450_y3;
  assign f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa426_y4 = f_s_dadda_pg_rca32_fa426_y4;
  assign f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa425_y4 = f_s_dadda_pg_rca32_fa425_y4;
  assign f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa424_y4 = f_s_dadda_pg_rca32_fa424_y4;
  assign f_s_dadda_pg_rca32_fa451_y0 = f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa426_y4 ^ f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa425_y4;
  assign f_s_dadda_pg_rca32_fa451_y1 = f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa426_y4 & f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa425_y4;
  assign f_s_dadda_pg_rca32_fa451_y2 = f_s_dadda_pg_rca32_fa451_y0 ^ f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa424_y4;
  assign f_s_dadda_pg_rca32_fa451_y3 = f_s_dadda_pg_rca32_fa451_y0 & f_s_dadda_pg_rca32_fa451_f_s_dadda_pg_rca32_fa424_y4;
  assign f_s_dadda_pg_rca32_fa451_y4 = f_s_dadda_pg_rca32_fa451_y1 | f_s_dadda_pg_rca32_fa451_y3;
  assign f_s_dadda_pg_rca32_nand_31_6_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_nand_31_6_y0 = ~(f_s_dadda_pg_rca32_nand_31_6_a_31 & f_s_dadda_pg_rca32_nand_31_6_b_6);
  assign f_s_dadda_pg_rca32_and_30_7_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_30_7_y0 = f_s_dadda_pg_rca32_and_30_7_a_30 & f_s_dadda_pg_rca32_and_30_7_b_7;
  assign f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_fa423_y4 = f_s_dadda_pg_rca32_fa423_y4;
  assign f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_nand_31_6_y0 = f_s_dadda_pg_rca32_nand_31_6_y0;
  assign f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_and_30_7_y0 = f_s_dadda_pg_rca32_and_30_7_y0;
  assign f_s_dadda_pg_rca32_fa452_y0 = f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_fa423_y4 ^ f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_nand_31_6_y0;
  assign f_s_dadda_pg_rca32_fa452_y1 = f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_fa423_y4 & f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_nand_31_6_y0;
  assign f_s_dadda_pg_rca32_fa452_y2 = f_s_dadda_pg_rca32_fa452_y0 ^ f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_and_30_7_y0;
  assign f_s_dadda_pg_rca32_fa452_y3 = f_s_dadda_pg_rca32_fa452_y0 & f_s_dadda_pg_rca32_fa452_f_s_dadda_pg_rca32_and_30_7_y0;
  assign f_s_dadda_pg_rca32_fa452_y4 = f_s_dadda_pg_rca32_fa452_y1 | f_s_dadda_pg_rca32_fa452_y3;
  assign f_s_dadda_pg_rca32_and_29_8_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_29_8_y0 = f_s_dadda_pg_rca32_and_29_8_a_29 & f_s_dadda_pg_rca32_and_29_8_b_8;
  assign f_s_dadda_pg_rca32_and_28_9_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_28_9_y0 = f_s_dadda_pg_rca32_and_28_9_a_28 & f_s_dadda_pg_rca32_and_28_9_b_9;
  assign f_s_dadda_pg_rca32_and_27_10_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_27_10_y0 = f_s_dadda_pg_rca32_and_27_10_a_27 & f_s_dadda_pg_rca32_and_27_10_b_10;
  assign f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_29_8_y0 = f_s_dadda_pg_rca32_and_29_8_y0;
  assign f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_28_9_y0 = f_s_dadda_pg_rca32_and_28_9_y0;
  assign f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_27_10_y0 = f_s_dadda_pg_rca32_and_27_10_y0;
  assign f_s_dadda_pg_rca32_fa453_y0 = f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_29_8_y0 ^ f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_28_9_y0;
  assign f_s_dadda_pg_rca32_fa453_y1 = f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_29_8_y0 & f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_28_9_y0;
  assign f_s_dadda_pg_rca32_fa453_y2 = f_s_dadda_pg_rca32_fa453_y0 ^ f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_27_10_y0;
  assign f_s_dadda_pg_rca32_fa453_y3 = f_s_dadda_pg_rca32_fa453_y0 & f_s_dadda_pg_rca32_fa453_f_s_dadda_pg_rca32_and_27_10_y0;
  assign f_s_dadda_pg_rca32_fa453_y4 = f_s_dadda_pg_rca32_fa453_y1 | f_s_dadda_pg_rca32_fa453_y3;
  assign f_s_dadda_pg_rca32_and_26_11_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_26_11_y0 = f_s_dadda_pg_rca32_and_26_11_a_26 & f_s_dadda_pg_rca32_and_26_11_b_11;
  assign f_s_dadda_pg_rca32_and_25_12_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_25_12_y0 = f_s_dadda_pg_rca32_and_25_12_a_25 & f_s_dadda_pg_rca32_and_25_12_b_12;
  assign f_s_dadda_pg_rca32_and_24_13_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_24_13_y0 = f_s_dadda_pg_rca32_and_24_13_a_24 & f_s_dadda_pg_rca32_and_24_13_b_13;
  assign f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_26_11_y0 = f_s_dadda_pg_rca32_and_26_11_y0;
  assign f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_25_12_y0 = f_s_dadda_pg_rca32_and_25_12_y0;
  assign f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_24_13_y0 = f_s_dadda_pg_rca32_and_24_13_y0;
  assign f_s_dadda_pg_rca32_fa454_y0 = f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_26_11_y0 ^ f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_25_12_y0;
  assign f_s_dadda_pg_rca32_fa454_y1 = f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_26_11_y0 & f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_25_12_y0;
  assign f_s_dadda_pg_rca32_fa454_y2 = f_s_dadda_pg_rca32_fa454_y0 ^ f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_24_13_y0;
  assign f_s_dadda_pg_rca32_fa454_y3 = f_s_dadda_pg_rca32_fa454_y0 & f_s_dadda_pg_rca32_fa454_f_s_dadda_pg_rca32_and_24_13_y0;
  assign f_s_dadda_pg_rca32_fa454_y4 = f_s_dadda_pg_rca32_fa454_y1 | f_s_dadda_pg_rca32_fa454_y3;
  assign f_s_dadda_pg_rca32_and_23_14_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_23_14_y0 = f_s_dadda_pg_rca32_and_23_14_a_23 & f_s_dadda_pg_rca32_and_23_14_b_14;
  assign f_s_dadda_pg_rca32_and_22_15_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_22_15_y0 = f_s_dadda_pg_rca32_and_22_15_a_22 & f_s_dadda_pg_rca32_and_22_15_b_15;
  assign f_s_dadda_pg_rca32_and_21_16_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_21_16_y0 = f_s_dadda_pg_rca32_and_21_16_a_21 & f_s_dadda_pg_rca32_and_21_16_b_16;
  assign f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_23_14_y0 = f_s_dadda_pg_rca32_and_23_14_y0;
  assign f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_22_15_y0 = f_s_dadda_pg_rca32_and_22_15_y0;
  assign f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_21_16_y0 = f_s_dadda_pg_rca32_and_21_16_y0;
  assign f_s_dadda_pg_rca32_fa455_y0 = f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_23_14_y0 ^ f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_22_15_y0;
  assign f_s_dadda_pg_rca32_fa455_y1 = f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_23_14_y0 & f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_22_15_y0;
  assign f_s_dadda_pg_rca32_fa455_y2 = f_s_dadda_pg_rca32_fa455_y0 ^ f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_21_16_y0;
  assign f_s_dadda_pg_rca32_fa455_y3 = f_s_dadda_pg_rca32_fa455_y0 & f_s_dadda_pg_rca32_fa455_f_s_dadda_pg_rca32_and_21_16_y0;
  assign f_s_dadda_pg_rca32_fa455_y4 = f_s_dadda_pg_rca32_fa455_y1 | f_s_dadda_pg_rca32_fa455_y3;
  assign f_s_dadda_pg_rca32_and_20_17_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_20_17_y0 = f_s_dadda_pg_rca32_and_20_17_a_20 & f_s_dadda_pg_rca32_and_20_17_b_17;
  assign f_s_dadda_pg_rca32_and_19_18_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_19_18_y0 = f_s_dadda_pg_rca32_and_19_18_a_19 & f_s_dadda_pg_rca32_and_19_18_b_18;
  assign f_s_dadda_pg_rca32_and_18_19_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_18_19_y0 = f_s_dadda_pg_rca32_and_18_19_a_18 & f_s_dadda_pg_rca32_and_18_19_b_19;
  assign f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_20_17_y0 = f_s_dadda_pg_rca32_and_20_17_y0;
  assign f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_19_18_y0 = f_s_dadda_pg_rca32_and_19_18_y0;
  assign f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_18_19_y0 = f_s_dadda_pg_rca32_and_18_19_y0;
  assign f_s_dadda_pg_rca32_fa456_y0 = f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_20_17_y0 ^ f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_19_18_y0;
  assign f_s_dadda_pg_rca32_fa456_y1 = f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_20_17_y0 & f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_19_18_y0;
  assign f_s_dadda_pg_rca32_fa456_y2 = f_s_dadda_pg_rca32_fa456_y0 ^ f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_18_19_y0;
  assign f_s_dadda_pg_rca32_fa456_y3 = f_s_dadda_pg_rca32_fa456_y0 & f_s_dadda_pg_rca32_fa456_f_s_dadda_pg_rca32_and_18_19_y0;
  assign f_s_dadda_pg_rca32_fa456_y4 = f_s_dadda_pg_rca32_fa456_y1 | f_s_dadda_pg_rca32_fa456_y3;
  assign f_s_dadda_pg_rca32_and_17_20_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_17_20_y0 = f_s_dadda_pg_rca32_and_17_20_a_17 & f_s_dadda_pg_rca32_and_17_20_b_20;
  assign f_s_dadda_pg_rca32_and_16_21_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_16_21_y0 = f_s_dadda_pg_rca32_and_16_21_a_16 & f_s_dadda_pg_rca32_and_16_21_b_21;
  assign f_s_dadda_pg_rca32_and_15_22_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_15_22_y0 = f_s_dadda_pg_rca32_and_15_22_a_15 & f_s_dadda_pg_rca32_and_15_22_b_22;
  assign f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_17_20_y0 = f_s_dadda_pg_rca32_and_17_20_y0;
  assign f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_16_21_y0 = f_s_dadda_pg_rca32_and_16_21_y0;
  assign f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_15_22_y0 = f_s_dadda_pg_rca32_and_15_22_y0;
  assign f_s_dadda_pg_rca32_fa457_y0 = f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_17_20_y0 ^ f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_16_21_y0;
  assign f_s_dadda_pg_rca32_fa457_y1 = f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_17_20_y0 & f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_16_21_y0;
  assign f_s_dadda_pg_rca32_fa457_y2 = f_s_dadda_pg_rca32_fa457_y0 ^ f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_15_22_y0;
  assign f_s_dadda_pg_rca32_fa457_y3 = f_s_dadda_pg_rca32_fa457_y0 & f_s_dadda_pg_rca32_fa457_f_s_dadda_pg_rca32_and_15_22_y0;
  assign f_s_dadda_pg_rca32_fa457_y4 = f_s_dadda_pg_rca32_fa457_y1 | f_s_dadda_pg_rca32_fa457_y3;
  assign f_s_dadda_pg_rca32_and_14_23_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_14_23_y0 = f_s_dadda_pg_rca32_and_14_23_a_14 & f_s_dadda_pg_rca32_and_14_23_b_23;
  assign f_s_dadda_pg_rca32_and_13_24_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_13_24_y0 = f_s_dadda_pg_rca32_and_13_24_a_13 & f_s_dadda_pg_rca32_and_13_24_b_24;
  assign f_s_dadda_pg_rca32_and_12_25_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_12_25_y0 = f_s_dadda_pg_rca32_and_12_25_a_12 & f_s_dadda_pg_rca32_and_12_25_b_25;
  assign f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_14_23_y0 = f_s_dadda_pg_rca32_and_14_23_y0;
  assign f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_13_24_y0 = f_s_dadda_pg_rca32_and_13_24_y0;
  assign f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_12_25_y0 = f_s_dadda_pg_rca32_and_12_25_y0;
  assign f_s_dadda_pg_rca32_fa458_y0 = f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_14_23_y0 ^ f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_13_24_y0;
  assign f_s_dadda_pg_rca32_fa458_y1 = f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_14_23_y0 & f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_13_24_y0;
  assign f_s_dadda_pg_rca32_fa458_y2 = f_s_dadda_pg_rca32_fa458_y0 ^ f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_12_25_y0;
  assign f_s_dadda_pg_rca32_fa458_y3 = f_s_dadda_pg_rca32_fa458_y0 & f_s_dadda_pg_rca32_fa458_f_s_dadda_pg_rca32_and_12_25_y0;
  assign f_s_dadda_pg_rca32_fa458_y4 = f_s_dadda_pg_rca32_fa458_y1 | f_s_dadda_pg_rca32_fa458_y3;
  assign f_s_dadda_pg_rca32_and_11_26_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_11_26_y0 = f_s_dadda_pg_rca32_and_11_26_a_11 & f_s_dadda_pg_rca32_and_11_26_b_26;
  assign f_s_dadda_pg_rca32_and_10_27_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_10_27_y0 = f_s_dadda_pg_rca32_and_10_27_a_10 & f_s_dadda_pg_rca32_and_10_27_b_27;
  assign f_s_dadda_pg_rca32_and_9_28_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_9_28_y0 = f_s_dadda_pg_rca32_and_9_28_a_9 & f_s_dadda_pg_rca32_and_9_28_b_28;
  assign f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_11_26_y0 = f_s_dadda_pg_rca32_and_11_26_y0;
  assign f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_10_27_y0 = f_s_dadda_pg_rca32_and_10_27_y0;
  assign f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_9_28_y0 = f_s_dadda_pg_rca32_and_9_28_y0;
  assign f_s_dadda_pg_rca32_fa459_y0 = f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_11_26_y0 ^ f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_10_27_y0;
  assign f_s_dadda_pg_rca32_fa459_y1 = f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_11_26_y0 & f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_10_27_y0;
  assign f_s_dadda_pg_rca32_fa459_y2 = f_s_dadda_pg_rca32_fa459_y0 ^ f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_9_28_y0;
  assign f_s_dadda_pg_rca32_fa459_y3 = f_s_dadda_pg_rca32_fa459_y0 & f_s_dadda_pg_rca32_fa459_f_s_dadda_pg_rca32_and_9_28_y0;
  assign f_s_dadda_pg_rca32_fa459_y4 = f_s_dadda_pg_rca32_fa459_y1 | f_s_dadda_pg_rca32_fa459_y3;
  assign f_s_dadda_pg_rca32_and_8_29_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_8_29_y0 = f_s_dadda_pg_rca32_and_8_29_a_8 & f_s_dadda_pg_rca32_and_8_29_b_29;
  assign f_s_dadda_pg_rca32_and_7_30_a_7 = a_7;
  assign f_s_dadda_pg_rca32_and_7_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_7_30_y0 = f_s_dadda_pg_rca32_and_7_30_a_7 & f_s_dadda_pg_rca32_and_7_30_b_30;
  assign f_s_dadda_pg_rca32_nand_6_31_a_6 = a_6;
  assign f_s_dadda_pg_rca32_nand_6_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_6_31_y0 = ~(f_s_dadda_pg_rca32_nand_6_31_a_6 & f_s_dadda_pg_rca32_nand_6_31_b_31);
  assign f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_and_8_29_y0 = f_s_dadda_pg_rca32_and_8_29_y0;
  assign f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_and_7_30_y0 = f_s_dadda_pg_rca32_and_7_30_y0;
  assign f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_nand_6_31_y0 = f_s_dadda_pg_rca32_nand_6_31_y0;
  assign f_s_dadda_pg_rca32_fa460_y0 = f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_and_8_29_y0 ^ f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_and_7_30_y0;
  assign f_s_dadda_pg_rca32_fa460_y1 = f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_and_8_29_y0 & f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_and_7_30_y0;
  assign f_s_dadda_pg_rca32_fa460_y2 = f_s_dadda_pg_rca32_fa460_y0 ^ f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_nand_6_31_y0;
  assign f_s_dadda_pg_rca32_fa460_y3 = f_s_dadda_pg_rca32_fa460_y0 & f_s_dadda_pg_rca32_fa460_f_s_dadda_pg_rca32_nand_6_31_y0;
  assign f_s_dadda_pg_rca32_fa460_y4 = f_s_dadda_pg_rca32_fa460_y1 | f_s_dadda_pg_rca32_fa460_y3;
  assign f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa445_y2 = f_s_dadda_pg_rca32_fa445_y2;
  assign f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa446_y2 = f_s_dadda_pg_rca32_fa446_y2;
  assign f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa447_y2 = f_s_dadda_pg_rca32_fa447_y2;
  assign f_s_dadda_pg_rca32_fa461_y0 = f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa445_y2 ^ f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa446_y2;
  assign f_s_dadda_pg_rca32_fa461_y1 = f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa445_y2 & f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa446_y2;
  assign f_s_dadda_pg_rca32_fa461_y2 = f_s_dadda_pg_rca32_fa461_y0 ^ f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa447_y2;
  assign f_s_dadda_pg_rca32_fa461_y3 = f_s_dadda_pg_rca32_fa461_y0 & f_s_dadda_pg_rca32_fa461_f_s_dadda_pg_rca32_fa447_y2;
  assign f_s_dadda_pg_rca32_fa461_y4 = f_s_dadda_pg_rca32_fa461_y1 | f_s_dadda_pg_rca32_fa461_y3;
  assign f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa448_y2 = f_s_dadda_pg_rca32_fa448_y2;
  assign f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa449_y2 = f_s_dadda_pg_rca32_fa449_y2;
  assign f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa450_y2 = f_s_dadda_pg_rca32_fa450_y2;
  assign f_s_dadda_pg_rca32_fa462_y0 = f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa448_y2 ^ f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa449_y2;
  assign f_s_dadda_pg_rca32_fa462_y1 = f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa448_y2 & f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa449_y2;
  assign f_s_dadda_pg_rca32_fa462_y2 = f_s_dadda_pg_rca32_fa462_y0 ^ f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa450_y2;
  assign f_s_dadda_pg_rca32_fa462_y3 = f_s_dadda_pg_rca32_fa462_y0 & f_s_dadda_pg_rca32_fa462_f_s_dadda_pg_rca32_fa450_y2;
  assign f_s_dadda_pg_rca32_fa462_y4 = f_s_dadda_pg_rca32_fa462_y1 | f_s_dadda_pg_rca32_fa462_y3;
  assign f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa451_y2 = f_s_dadda_pg_rca32_fa451_y2;
  assign f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa452_y2 = f_s_dadda_pg_rca32_fa452_y2;
  assign f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa453_y2 = f_s_dadda_pg_rca32_fa453_y2;
  assign f_s_dadda_pg_rca32_fa463_y0 = f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa451_y2 ^ f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa452_y2;
  assign f_s_dadda_pg_rca32_fa463_y1 = f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa451_y2 & f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa452_y2;
  assign f_s_dadda_pg_rca32_fa463_y2 = f_s_dadda_pg_rca32_fa463_y0 ^ f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa453_y2;
  assign f_s_dadda_pg_rca32_fa463_y3 = f_s_dadda_pg_rca32_fa463_y0 & f_s_dadda_pg_rca32_fa463_f_s_dadda_pg_rca32_fa453_y2;
  assign f_s_dadda_pg_rca32_fa463_y4 = f_s_dadda_pg_rca32_fa463_y1 | f_s_dadda_pg_rca32_fa463_y3;
  assign f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa454_y2 = f_s_dadda_pg_rca32_fa454_y2;
  assign f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa455_y2 = f_s_dadda_pg_rca32_fa455_y2;
  assign f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa456_y2 = f_s_dadda_pg_rca32_fa456_y2;
  assign f_s_dadda_pg_rca32_fa464_y0 = f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa454_y2 ^ f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa455_y2;
  assign f_s_dadda_pg_rca32_fa464_y1 = f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa454_y2 & f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa455_y2;
  assign f_s_dadda_pg_rca32_fa464_y2 = f_s_dadda_pg_rca32_fa464_y0 ^ f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa456_y2;
  assign f_s_dadda_pg_rca32_fa464_y3 = f_s_dadda_pg_rca32_fa464_y0 & f_s_dadda_pg_rca32_fa464_f_s_dadda_pg_rca32_fa456_y2;
  assign f_s_dadda_pg_rca32_fa464_y4 = f_s_dadda_pg_rca32_fa464_y1 | f_s_dadda_pg_rca32_fa464_y3;
  assign f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa457_y2 = f_s_dadda_pg_rca32_fa457_y2;
  assign f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa458_y2 = f_s_dadda_pg_rca32_fa458_y2;
  assign f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa459_y2 = f_s_dadda_pg_rca32_fa459_y2;
  assign f_s_dadda_pg_rca32_fa465_y0 = f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa457_y2 ^ f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa458_y2;
  assign f_s_dadda_pg_rca32_fa465_y1 = f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa457_y2 & f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa458_y2;
  assign f_s_dadda_pg_rca32_fa465_y2 = f_s_dadda_pg_rca32_fa465_y0 ^ f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa459_y2;
  assign f_s_dadda_pg_rca32_fa465_y3 = f_s_dadda_pg_rca32_fa465_y0 & f_s_dadda_pg_rca32_fa465_f_s_dadda_pg_rca32_fa459_y2;
  assign f_s_dadda_pg_rca32_fa465_y4 = f_s_dadda_pg_rca32_fa465_y1 | f_s_dadda_pg_rca32_fa465_y3;
  assign f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa465_y4 = f_s_dadda_pg_rca32_fa465_y4;
  assign f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa464_y4 = f_s_dadda_pg_rca32_fa464_y4;
  assign f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa463_y4 = f_s_dadda_pg_rca32_fa463_y4;
  assign f_s_dadda_pg_rca32_fa466_y0 = f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa465_y4 ^ f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa464_y4;
  assign f_s_dadda_pg_rca32_fa466_y1 = f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa465_y4 & f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa464_y4;
  assign f_s_dadda_pg_rca32_fa466_y2 = f_s_dadda_pg_rca32_fa466_y0 ^ f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa463_y4;
  assign f_s_dadda_pg_rca32_fa466_y3 = f_s_dadda_pg_rca32_fa466_y0 & f_s_dadda_pg_rca32_fa466_f_s_dadda_pg_rca32_fa463_y4;
  assign f_s_dadda_pg_rca32_fa466_y4 = f_s_dadda_pg_rca32_fa466_y1 | f_s_dadda_pg_rca32_fa466_y3;
  assign f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa462_y4 = f_s_dadda_pg_rca32_fa462_y4;
  assign f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa461_y4 = f_s_dadda_pg_rca32_fa461_y4;
  assign f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa460_y4 = f_s_dadda_pg_rca32_fa460_y4;
  assign f_s_dadda_pg_rca32_fa467_y0 = f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa462_y4 ^ f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa461_y4;
  assign f_s_dadda_pg_rca32_fa467_y1 = f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa462_y4 & f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa461_y4;
  assign f_s_dadda_pg_rca32_fa467_y2 = f_s_dadda_pg_rca32_fa467_y0 ^ f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa460_y4;
  assign f_s_dadda_pg_rca32_fa467_y3 = f_s_dadda_pg_rca32_fa467_y0 & f_s_dadda_pg_rca32_fa467_f_s_dadda_pg_rca32_fa460_y4;
  assign f_s_dadda_pg_rca32_fa467_y4 = f_s_dadda_pg_rca32_fa467_y1 | f_s_dadda_pg_rca32_fa467_y3;
  assign f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa459_y4 = f_s_dadda_pg_rca32_fa459_y4;
  assign f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa458_y4 = f_s_dadda_pg_rca32_fa458_y4;
  assign f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa457_y4 = f_s_dadda_pg_rca32_fa457_y4;
  assign f_s_dadda_pg_rca32_fa468_y0 = f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa459_y4 ^ f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa458_y4;
  assign f_s_dadda_pg_rca32_fa468_y1 = f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa459_y4 & f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa458_y4;
  assign f_s_dadda_pg_rca32_fa468_y2 = f_s_dadda_pg_rca32_fa468_y0 ^ f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa457_y4;
  assign f_s_dadda_pg_rca32_fa468_y3 = f_s_dadda_pg_rca32_fa468_y0 & f_s_dadda_pg_rca32_fa468_f_s_dadda_pg_rca32_fa457_y4;
  assign f_s_dadda_pg_rca32_fa468_y4 = f_s_dadda_pg_rca32_fa468_y1 | f_s_dadda_pg_rca32_fa468_y3;
  assign f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa456_y4 = f_s_dadda_pg_rca32_fa456_y4;
  assign f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa455_y4 = f_s_dadda_pg_rca32_fa455_y4;
  assign f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa454_y4 = f_s_dadda_pg_rca32_fa454_y4;
  assign f_s_dadda_pg_rca32_fa469_y0 = f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa456_y4 ^ f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa455_y4;
  assign f_s_dadda_pg_rca32_fa469_y1 = f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa456_y4 & f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa455_y4;
  assign f_s_dadda_pg_rca32_fa469_y2 = f_s_dadda_pg_rca32_fa469_y0 ^ f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa454_y4;
  assign f_s_dadda_pg_rca32_fa469_y3 = f_s_dadda_pg_rca32_fa469_y0 & f_s_dadda_pg_rca32_fa469_f_s_dadda_pg_rca32_fa454_y4;
  assign f_s_dadda_pg_rca32_fa469_y4 = f_s_dadda_pg_rca32_fa469_y1 | f_s_dadda_pg_rca32_fa469_y3;
  assign f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa453_y4 = f_s_dadda_pg_rca32_fa453_y4;
  assign f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa452_y4 = f_s_dadda_pg_rca32_fa452_y4;
  assign f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa451_y4 = f_s_dadda_pg_rca32_fa451_y4;
  assign f_s_dadda_pg_rca32_fa470_y0 = f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa453_y4 ^ f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa452_y4;
  assign f_s_dadda_pg_rca32_fa470_y1 = f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa453_y4 & f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa452_y4;
  assign f_s_dadda_pg_rca32_fa470_y2 = f_s_dadda_pg_rca32_fa470_y0 ^ f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa451_y4;
  assign f_s_dadda_pg_rca32_fa470_y3 = f_s_dadda_pg_rca32_fa470_y0 & f_s_dadda_pg_rca32_fa470_f_s_dadda_pg_rca32_fa451_y4;
  assign f_s_dadda_pg_rca32_fa470_y4 = f_s_dadda_pg_rca32_fa470_y1 | f_s_dadda_pg_rca32_fa470_y3;
  assign f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa450_y4 = f_s_dadda_pg_rca32_fa450_y4;
  assign f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa449_y4 = f_s_dadda_pg_rca32_fa449_y4;
  assign f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa448_y4 = f_s_dadda_pg_rca32_fa448_y4;
  assign f_s_dadda_pg_rca32_fa471_y0 = f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa450_y4 ^ f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa449_y4;
  assign f_s_dadda_pg_rca32_fa471_y1 = f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa450_y4 & f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa449_y4;
  assign f_s_dadda_pg_rca32_fa471_y2 = f_s_dadda_pg_rca32_fa471_y0 ^ f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa448_y4;
  assign f_s_dadda_pg_rca32_fa471_y3 = f_s_dadda_pg_rca32_fa471_y0 & f_s_dadda_pg_rca32_fa471_f_s_dadda_pg_rca32_fa448_y4;
  assign f_s_dadda_pg_rca32_fa471_y4 = f_s_dadda_pg_rca32_fa471_y1 | f_s_dadda_pg_rca32_fa471_y3;
  assign f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa447_y4 = f_s_dadda_pg_rca32_fa447_y4;
  assign f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa446_y4 = f_s_dadda_pg_rca32_fa446_y4;
  assign f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa445_y4 = f_s_dadda_pg_rca32_fa445_y4;
  assign f_s_dadda_pg_rca32_fa472_y0 = f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa447_y4 ^ f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa446_y4;
  assign f_s_dadda_pg_rca32_fa472_y1 = f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa447_y4 & f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa446_y4;
  assign f_s_dadda_pg_rca32_fa472_y2 = f_s_dadda_pg_rca32_fa472_y0 ^ f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa445_y4;
  assign f_s_dadda_pg_rca32_fa472_y3 = f_s_dadda_pg_rca32_fa472_y0 & f_s_dadda_pg_rca32_fa472_f_s_dadda_pg_rca32_fa445_y4;
  assign f_s_dadda_pg_rca32_fa472_y4 = f_s_dadda_pg_rca32_fa472_y1 | f_s_dadda_pg_rca32_fa472_y3;
  assign f_s_dadda_pg_rca32_nand_31_7_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_nand_31_7_y0 = ~(f_s_dadda_pg_rca32_nand_31_7_a_31 & f_s_dadda_pg_rca32_nand_31_7_b_7);
  assign f_s_dadda_pg_rca32_and_30_8_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_30_8_y0 = f_s_dadda_pg_rca32_and_30_8_a_30 & f_s_dadda_pg_rca32_and_30_8_b_8;
  assign f_s_dadda_pg_rca32_and_29_9_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_29_9_y0 = f_s_dadda_pg_rca32_and_29_9_a_29 & f_s_dadda_pg_rca32_and_29_9_b_9;
  assign f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_nand_31_7_y0 = f_s_dadda_pg_rca32_nand_31_7_y0;
  assign f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_and_30_8_y0 = f_s_dadda_pg_rca32_and_30_8_y0;
  assign f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_and_29_9_y0 = f_s_dadda_pg_rca32_and_29_9_y0;
  assign f_s_dadda_pg_rca32_fa473_y0 = f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_nand_31_7_y0 ^ f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_and_30_8_y0;
  assign f_s_dadda_pg_rca32_fa473_y1 = f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_nand_31_7_y0 & f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_and_30_8_y0;
  assign f_s_dadda_pg_rca32_fa473_y2 = f_s_dadda_pg_rca32_fa473_y0 ^ f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_and_29_9_y0;
  assign f_s_dadda_pg_rca32_fa473_y3 = f_s_dadda_pg_rca32_fa473_y0 & f_s_dadda_pg_rca32_fa473_f_s_dadda_pg_rca32_and_29_9_y0;
  assign f_s_dadda_pg_rca32_fa473_y4 = f_s_dadda_pg_rca32_fa473_y1 | f_s_dadda_pg_rca32_fa473_y3;
  assign f_s_dadda_pg_rca32_and_28_10_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_28_10_y0 = f_s_dadda_pg_rca32_and_28_10_a_28 & f_s_dadda_pg_rca32_and_28_10_b_10;
  assign f_s_dadda_pg_rca32_and_27_11_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_27_11_y0 = f_s_dadda_pg_rca32_and_27_11_a_27 & f_s_dadda_pg_rca32_and_27_11_b_11;
  assign f_s_dadda_pg_rca32_and_26_12_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_26_12_y0 = f_s_dadda_pg_rca32_and_26_12_a_26 & f_s_dadda_pg_rca32_and_26_12_b_12;
  assign f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_28_10_y0 = f_s_dadda_pg_rca32_and_28_10_y0;
  assign f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_27_11_y0 = f_s_dadda_pg_rca32_and_27_11_y0;
  assign f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_26_12_y0 = f_s_dadda_pg_rca32_and_26_12_y0;
  assign f_s_dadda_pg_rca32_fa474_y0 = f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_28_10_y0 ^ f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_27_11_y0;
  assign f_s_dadda_pg_rca32_fa474_y1 = f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_28_10_y0 & f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_27_11_y0;
  assign f_s_dadda_pg_rca32_fa474_y2 = f_s_dadda_pg_rca32_fa474_y0 ^ f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_26_12_y0;
  assign f_s_dadda_pg_rca32_fa474_y3 = f_s_dadda_pg_rca32_fa474_y0 & f_s_dadda_pg_rca32_fa474_f_s_dadda_pg_rca32_and_26_12_y0;
  assign f_s_dadda_pg_rca32_fa474_y4 = f_s_dadda_pg_rca32_fa474_y1 | f_s_dadda_pg_rca32_fa474_y3;
  assign f_s_dadda_pg_rca32_and_25_13_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_25_13_y0 = f_s_dadda_pg_rca32_and_25_13_a_25 & f_s_dadda_pg_rca32_and_25_13_b_13;
  assign f_s_dadda_pg_rca32_and_24_14_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_24_14_y0 = f_s_dadda_pg_rca32_and_24_14_a_24 & f_s_dadda_pg_rca32_and_24_14_b_14;
  assign f_s_dadda_pg_rca32_and_23_15_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_23_15_y0 = f_s_dadda_pg_rca32_and_23_15_a_23 & f_s_dadda_pg_rca32_and_23_15_b_15;
  assign f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_25_13_y0 = f_s_dadda_pg_rca32_and_25_13_y0;
  assign f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_24_14_y0 = f_s_dadda_pg_rca32_and_24_14_y0;
  assign f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_23_15_y0 = f_s_dadda_pg_rca32_and_23_15_y0;
  assign f_s_dadda_pg_rca32_fa475_y0 = f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_25_13_y0 ^ f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_24_14_y0;
  assign f_s_dadda_pg_rca32_fa475_y1 = f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_25_13_y0 & f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_24_14_y0;
  assign f_s_dadda_pg_rca32_fa475_y2 = f_s_dadda_pg_rca32_fa475_y0 ^ f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_23_15_y0;
  assign f_s_dadda_pg_rca32_fa475_y3 = f_s_dadda_pg_rca32_fa475_y0 & f_s_dadda_pg_rca32_fa475_f_s_dadda_pg_rca32_and_23_15_y0;
  assign f_s_dadda_pg_rca32_fa475_y4 = f_s_dadda_pg_rca32_fa475_y1 | f_s_dadda_pg_rca32_fa475_y3;
  assign f_s_dadda_pg_rca32_and_22_16_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_22_16_y0 = f_s_dadda_pg_rca32_and_22_16_a_22 & f_s_dadda_pg_rca32_and_22_16_b_16;
  assign f_s_dadda_pg_rca32_and_21_17_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_21_17_y0 = f_s_dadda_pg_rca32_and_21_17_a_21 & f_s_dadda_pg_rca32_and_21_17_b_17;
  assign f_s_dadda_pg_rca32_and_20_18_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_20_18_y0 = f_s_dadda_pg_rca32_and_20_18_a_20 & f_s_dadda_pg_rca32_and_20_18_b_18;
  assign f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_22_16_y0 = f_s_dadda_pg_rca32_and_22_16_y0;
  assign f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_21_17_y0 = f_s_dadda_pg_rca32_and_21_17_y0;
  assign f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_20_18_y0 = f_s_dadda_pg_rca32_and_20_18_y0;
  assign f_s_dadda_pg_rca32_fa476_y0 = f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_22_16_y0 ^ f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_21_17_y0;
  assign f_s_dadda_pg_rca32_fa476_y1 = f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_22_16_y0 & f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_21_17_y0;
  assign f_s_dadda_pg_rca32_fa476_y2 = f_s_dadda_pg_rca32_fa476_y0 ^ f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_20_18_y0;
  assign f_s_dadda_pg_rca32_fa476_y3 = f_s_dadda_pg_rca32_fa476_y0 & f_s_dadda_pg_rca32_fa476_f_s_dadda_pg_rca32_and_20_18_y0;
  assign f_s_dadda_pg_rca32_fa476_y4 = f_s_dadda_pg_rca32_fa476_y1 | f_s_dadda_pg_rca32_fa476_y3;
  assign f_s_dadda_pg_rca32_and_19_19_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_19_19_y0 = f_s_dadda_pg_rca32_and_19_19_a_19 & f_s_dadda_pg_rca32_and_19_19_b_19;
  assign f_s_dadda_pg_rca32_and_18_20_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_18_20_y0 = f_s_dadda_pg_rca32_and_18_20_a_18 & f_s_dadda_pg_rca32_and_18_20_b_20;
  assign f_s_dadda_pg_rca32_and_17_21_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_17_21_y0 = f_s_dadda_pg_rca32_and_17_21_a_17 & f_s_dadda_pg_rca32_and_17_21_b_21;
  assign f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_19_19_y0 = f_s_dadda_pg_rca32_and_19_19_y0;
  assign f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_18_20_y0 = f_s_dadda_pg_rca32_and_18_20_y0;
  assign f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_17_21_y0 = f_s_dadda_pg_rca32_and_17_21_y0;
  assign f_s_dadda_pg_rca32_fa477_y0 = f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_19_19_y0 ^ f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_18_20_y0;
  assign f_s_dadda_pg_rca32_fa477_y1 = f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_19_19_y0 & f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_18_20_y0;
  assign f_s_dadda_pg_rca32_fa477_y2 = f_s_dadda_pg_rca32_fa477_y0 ^ f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_17_21_y0;
  assign f_s_dadda_pg_rca32_fa477_y3 = f_s_dadda_pg_rca32_fa477_y0 & f_s_dadda_pg_rca32_fa477_f_s_dadda_pg_rca32_and_17_21_y0;
  assign f_s_dadda_pg_rca32_fa477_y4 = f_s_dadda_pg_rca32_fa477_y1 | f_s_dadda_pg_rca32_fa477_y3;
  assign f_s_dadda_pg_rca32_and_16_22_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_16_22_y0 = f_s_dadda_pg_rca32_and_16_22_a_16 & f_s_dadda_pg_rca32_and_16_22_b_22;
  assign f_s_dadda_pg_rca32_and_15_23_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_15_23_y0 = f_s_dadda_pg_rca32_and_15_23_a_15 & f_s_dadda_pg_rca32_and_15_23_b_23;
  assign f_s_dadda_pg_rca32_and_14_24_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_14_24_y0 = f_s_dadda_pg_rca32_and_14_24_a_14 & f_s_dadda_pg_rca32_and_14_24_b_24;
  assign f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_16_22_y0 = f_s_dadda_pg_rca32_and_16_22_y0;
  assign f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_15_23_y0 = f_s_dadda_pg_rca32_and_15_23_y0;
  assign f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_14_24_y0 = f_s_dadda_pg_rca32_and_14_24_y0;
  assign f_s_dadda_pg_rca32_fa478_y0 = f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_16_22_y0 ^ f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_15_23_y0;
  assign f_s_dadda_pg_rca32_fa478_y1 = f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_16_22_y0 & f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_15_23_y0;
  assign f_s_dadda_pg_rca32_fa478_y2 = f_s_dadda_pg_rca32_fa478_y0 ^ f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_14_24_y0;
  assign f_s_dadda_pg_rca32_fa478_y3 = f_s_dadda_pg_rca32_fa478_y0 & f_s_dadda_pg_rca32_fa478_f_s_dadda_pg_rca32_and_14_24_y0;
  assign f_s_dadda_pg_rca32_fa478_y4 = f_s_dadda_pg_rca32_fa478_y1 | f_s_dadda_pg_rca32_fa478_y3;
  assign f_s_dadda_pg_rca32_and_13_25_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_13_25_y0 = f_s_dadda_pg_rca32_and_13_25_a_13 & f_s_dadda_pg_rca32_and_13_25_b_25;
  assign f_s_dadda_pg_rca32_and_12_26_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_12_26_y0 = f_s_dadda_pg_rca32_and_12_26_a_12 & f_s_dadda_pg_rca32_and_12_26_b_26;
  assign f_s_dadda_pg_rca32_and_11_27_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_11_27_y0 = f_s_dadda_pg_rca32_and_11_27_a_11 & f_s_dadda_pg_rca32_and_11_27_b_27;
  assign f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_13_25_y0 = f_s_dadda_pg_rca32_and_13_25_y0;
  assign f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_12_26_y0 = f_s_dadda_pg_rca32_and_12_26_y0;
  assign f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_11_27_y0 = f_s_dadda_pg_rca32_and_11_27_y0;
  assign f_s_dadda_pg_rca32_fa479_y0 = f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_13_25_y0 ^ f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_12_26_y0;
  assign f_s_dadda_pg_rca32_fa479_y1 = f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_13_25_y0 & f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_12_26_y0;
  assign f_s_dadda_pg_rca32_fa479_y2 = f_s_dadda_pg_rca32_fa479_y0 ^ f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_11_27_y0;
  assign f_s_dadda_pg_rca32_fa479_y3 = f_s_dadda_pg_rca32_fa479_y0 & f_s_dadda_pg_rca32_fa479_f_s_dadda_pg_rca32_and_11_27_y0;
  assign f_s_dadda_pg_rca32_fa479_y4 = f_s_dadda_pg_rca32_fa479_y1 | f_s_dadda_pg_rca32_fa479_y3;
  assign f_s_dadda_pg_rca32_and_10_28_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_10_28_y0 = f_s_dadda_pg_rca32_and_10_28_a_10 & f_s_dadda_pg_rca32_and_10_28_b_28;
  assign f_s_dadda_pg_rca32_and_9_29_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_9_29_y0 = f_s_dadda_pg_rca32_and_9_29_a_9 & f_s_dadda_pg_rca32_and_9_29_b_29;
  assign f_s_dadda_pg_rca32_and_8_30_a_8 = a_8;
  assign f_s_dadda_pg_rca32_and_8_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_8_30_y0 = f_s_dadda_pg_rca32_and_8_30_a_8 & f_s_dadda_pg_rca32_and_8_30_b_30;
  assign f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_10_28_y0 = f_s_dadda_pg_rca32_and_10_28_y0;
  assign f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_9_29_y0 = f_s_dadda_pg_rca32_and_9_29_y0;
  assign f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_8_30_y0 = f_s_dadda_pg_rca32_and_8_30_y0;
  assign f_s_dadda_pg_rca32_fa480_y0 = f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_10_28_y0 ^ f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_9_29_y0;
  assign f_s_dadda_pg_rca32_fa480_y1 = f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_10_28_y0 & f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_9_29_y0;
  assign f_s_dadda_pg_rca32_fa480_y2 = f_s_dadda_pg_rca32_fa480_y0 ^ f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_8_30_y0;
  assign f_s_dadda_pg_rca32_fa480_y3 = f_s_dadda_pg_rca32_fa480_y0 & f_s_dadda_pg_rca32_fa480_f_s_dadda_pg_rca32_and_8_30_y0;
  assign f_s_dadda_pg_rca32_fa480_y4 = f_s_dadda_pg_rca32_fa480_y1 | f_s_dadda_pg_rca32_fa480_y3;
  assign f_s_dadda_pg_rca32_nand_7_31_a_7 = a_7;
  assign f_s_dadda_pg_rca32_nand_7_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_7_31_y0 = ~(f_s_dadda_pg_rca32_nand_7_31_a_7 & f_s_dadda_pg_rca32_nand_7_31_b_31);
  assign f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_nand_7_31_y0 = f_s_dadda_pg_rca32_nand_7_31_y0;
  assign f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_fa466_y2 = f_s_dadda_pg_rca32_fa466_y2;
  assign f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_fa467_y2 = f_s_dadda_pg_rca32_fa467_y2;
  assign f_s_dadda_pg_rca32_fa481_y0 = f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_nand_7_31_y0 ^ f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_fa466_y2;
  assign f_s_dadda_pg_rca32_fa481_y1 = f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_nand_7_31_y0 & f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_fa466_y2;
  assign f_s_dadda_pg_rca32_fa481_y2 = f_s_dadda_pg_rca32_fa481_y0 ^ f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_fa467_y2;
  assign f_s_dadda_pg_rca32_fa481_y3 = f_s_dadda_pg_rca32_fa481_y0 & f_s_dadda_pg_rca32_fa481_f_s_dadda_pg_rca32_fa467_y2;
  assign f_s_dadda_pg_rca32_fa481_y4 = f_s_dadda_pg_rca32_fa481_y1 | f_s_dadda_pg_rca32_fa481_y3;
  assign f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa468_y2 = f_s_dadda_pg_rca32_fa468_y2;
  assign f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa469_y2 = f_s_dadda_pg_rca32_fa469_y2;
  assign f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa470_y2 = f_s_dadda_pg_rca32_fa470_y2;
  assign f_s_dadda_pg_rca32_fa482_y0 = f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa468_y2 ^ f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa469_y2;
  assign f_s_dadda_pg_rca32_fa482_y1 = f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa468_y2 & f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa469_y2;
  assign f_s_dadda_pg_rca32_fa482_y2 = f_s_dadda_pg_rca32_fa482_y0 ^ f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa470_y2;
  assign f_s_dadda_pg_rca32_fa482_y3 = f_s_dadda_pg_rca32_fa482_y0 & f_s_dadda_pg_rca32_fa482_f_s_dadda_pg_rca32_fa470_y2;
  assign f_s_dadda_pg_rca32_fa482_y4 = f_s_dadda_pg_rca32_fa482_y1 | f_s_dadda_pg_rca32_fa482_y3;
  assign f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa471_y2 = f_s_dadda_pg_rca32_fa471_y2;
  assign f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa472_y2 = f_s_dadda_pg_rca32_fa472_y2;
  assign f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa473_y2 = f_s_dadda_pg_rca32_fa473_y2;
  assign f_s_dadda_pg_rca32_fa483_y0 = f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa471_y2 ^ f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa472_y2;
  assign f_s_dadda_pg_rca32_fa483_y1 = f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa471_y2 & f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa472_y2;
  assign f_s_dadda_pg_rca32_fa483_y2 = f_s_dadda_pg_rca32_fa483_y0 ^ f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa473_y2;
  assign f_s_dadda_pg_rca32_fa483_y3 = f_s_dadda_pg_rca32_fa483_y0 & f_s_dadda_pg_rca32_fa483_f_s_dadda_pg_rca32_fa473_y2;
  assign f_s_dadda_pg_rca32_fa483_y4 = f_s_dadda_pg_rca32_fa483_y1 | f_s_dadda_pg_rca32_fa483_y3;
  assign f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa474_y2 = f_s_dadda_pg_rca32_fa474_y2;
  assign f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa475_y2 = f_s_dadda_pg_rca32_fa475_y2;
  assign f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa476_y2 = f_s_dadda_pg_rca32_fa476_y2;
  assign f_s_dadda_pg_rca32_fa484_y0 = f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa474_y2 ^ f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa475_y2;
  assign f_s_dadda_pg_rca32_fa484_y1 = f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa474_y2 & f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa475_y2;
  assign f_s_dadda_pg_rca32_fa484_y2 = f_s_dadda_pg_rca32_fa484_y0 ^ f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa476_y2;
  assign f_s_dadda_pg_rca32_fa484_y3 = f_s_dadda_pg_rca32_fa484_y0 & f_s_dadda_pg_rca32_fa484_f_s_dadda_pg_rca32_fa476_y2;
  assign f_s_dadda_pg_rca32_fa484_y4 = f_s_dadda_pg_rca32_fa484_y1 | f_s_dadda_pg_rca32_fa484_y3;
  assign f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa477_y2 = f_s_dadda_pg_rca32_fa477_y2;
  assign f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa478_y2 = f_s_dadda_pg_rca32_fa478_y2;
  assign f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa479_y2 = f_s_dadda_pg_rca32_fa479_y2;
  assign f_s_dadda_pg_rca32_fa485_y0 = f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa477_y2 ^ f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa478_y2;
  assign f_s_dadda_pg_rca32_fa485_y1 = f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa477_y2 & f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa478_y2;
  assign f_s_dadda_pg_rca32_fa485_y2 = f_s_dadda_pg_rca32_fa485_y0 ^ f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa479_y2;
  assign f_s_dadda_pg_rca32_fa485_y3 = f_s_dadda_pg_rca32_fa485_y0 & f_s_dadda_pg_rca32_fa485_f_s_dadda_pg_rca32_fa479_y2;
  assign f_s_dadda_pg_rca32_fa485_y4 = f_s_dadda_pg_rca32_fa485_y1 | f_s_dadda_pg_rca32_fa485_y3;
  assign f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa485_y4 = f_s_dadda_pg_rca32_fa485_y4;
  assign f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa484_y4 = f_s_dadda_pg_rca32_fa484_y4;
  assign f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa483_y4 = f_s_dadda_pg_rca32_fa483_y4;
  assign f_s_dadda_pg_rca32_fa486_y0 = f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa485_y4 ^ f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa484_y4;
  assign f_s_dadda_pg_rca32_fa486_y1 = f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa485_y4 & f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa484_y4;
  assign f_s_dadda_pg_rca32_fa486_y2 = f_s_dadda_pg_rca32_fa486_y0 ^ f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa483_y4;
  assign f_s_dadda_pg_rca32_fa486_y3 = f_s_dadda_pg_rca32_fa486_y0 & f_s_dadda_pg_rca32_fa486_f_s_dadda_pg_rca32_fa483_y4;
  assign f_s_dadda_pg_rca32_fa486_y4 = f_s_dadda_pg_rca32_fa486_y1 | f_s_dadda_pg_rca32_fa486_y3;
  assign f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa482_y4 = f_s_dadda_pg_rca32_fa482_y4;
  assign f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa481_y4 = f_s_dadda_pg_rca32_fa481_y4;
  assign f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa480_y4 = f_s_dadda_pg_rca32_fa480_y4;
  assign f_s_dadda_pg_rca32_fa487_y0 = f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa482_y4 ^ f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa481_y4;
  assign f_s_dadda_pg_rca32_fa487_y1 = f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa482_y4 & f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa481_y4;
  assign f_s_dadda_pg_rca32_fa487_y2 = f_s_dadda_pg_rca32_fa487_y0 ^ f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa480_y4;
  assign f_s_dadda_pg_rca32_fa487_y3 = f_s_dadda_pg_rca32_fa487_y0 & f_s_dadda_pg_rca32_fa487_f_s_dadda_pg_rca32_fa480_y4;
  assign f_s_dadda_pg_rca32_fa487_y4 = f_s_dadda_pg_rca32_fa487_y1 | f_s_dadda_pg_rca32_fa487_y3;
  assign f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa479_y4 = f_s_dadda_pg_rca32_fa479_y4;
  assign f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa478_y4 = f_s_dadda_pg_rca32_fa478_y4;
  assign f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa477_y4 = f_s_dadda_pg_rca32_fa477_y4;
  assign f_s_dadda_pg_rca32_fa488_y0 = f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa479_y4 ^ f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa478_y4;
  assign f_s_dadda_pg_rca32_fa488_y1 = f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa479_y4 & f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa478_y4;
  assign f_s_dadda_pg_rca32_fa488_y2 = f_s_dadda_pg_rca32_fa488_y0 ^ f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa477_y4;
  assign f_s_dadda_pg_rca32_fa488_y3 = f_s_dadda_pg_rca32_fa488_y0 & f_s_dadda_pg_rca32_fa488_f_s_dadda_pg_rca32_fa477_y4;
  assign f_s_dadda_pg_rca32_fa488_y4 = f_s_dadda_pg_rca32_fa488_y1 | f_s_dadda_pg_rca32_fa488_y3;
  assign f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa476_y4 = f_s_dadda_pg_rca32_fa476_y4;
  assign f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa475_y4 = f_s_dadda_pg_rca32_fa475_y4;
  assign f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa474_y4 = f_s_dadda_pg_rca32_fa474_y4;
  assign f_s_dadda_pg_rca32_fa489_y0 = f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa476_y4 ^ f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa475_y4;
  assign f_s_dadda_pg_rca32_fa489_y1 = f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa476_y4 & f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa475_y4;
  assign f_s_dadda_pg_rca32_fa489_y2 = f_s_dadda_pg_rca32_fa489_y0 ^ f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa474_y4;
  assign f_s_dadda_pg_rca32_fa489_y3 = f_s_dadda_pg_rca32_fa489_y0 & f_s_dadda_pg_rca32_fa489_f_s_dadda_pg_rca32_fa474_y4;
  assign f_s_dadda_pg_rca32_fa489_y4 = f_s_dadda_pg_rca32_fa489_y1 | f_s_dadda_pg_rca32_fa489_y3;
  assign f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa473_y4 = f_s_dadda_pg_rca32_fa473_y4;
  assign f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa472_y4 = f_s_dadda_pg_rca32_fa472_y4;
  assign f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa471_y4 = f_s_dadda_pg_rca32_fa471_y4;
  assign f_s_dadda_pg_rca32_fa490_y0 = f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa473_y4 ^ f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa472_y4;
  assign f_s_dadda_pg_rca32_fa490_y1 = f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa473_y4 & f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa472_y4;
  assign f_s_dadda_pg_rca32_fa490_y2 = f_s_dadda_pg_rca32_fa490_y0 ^ f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa471_y4;
  assign f_s_dadda_pg_rca32_fa490_y3 = f_s_dadda_pg_rca32_fa490_y0 & f_s_dadda_pg_rca32_fa490_f_s_dadda_pg_rca32_fa471_y4;
  assign f_s_dadda_pg_rca32_fa490_y4 = f_s_dadda_pg_rca32_fa490_y1 | f_s_dadda_pg_rca32_fa490_y3;
  assign f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa470_y4 = f_s_dadda_pg_rca32_fa470_y4;
  assign f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa469_y4 = f_s_dadda_pg_rca32_fa469_y4;
  assign f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa468_y4 = f_s_dadda_pg_rca32_fa468_y4;
  assign f_s_dadda_pg_rca32_fa491_y0 = f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa470_y4 ^ f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa469_y4;
  assign f_s_dadda_pg_rca32_fa491_y1 = f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa470_y4 & f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa469_y4;
  assign f_s_dadda_pg_rca32_fa491_y2 = f_s_dadda_pg_rca32_fa491_y0 ^ f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa468_y4;
  assign f_s_dadda_pg_rca32_fa491_y3 = f_s_dadda_pg_rca32_fa491_y0 & f_s_dadda_pg_rca32_fa491_f_s_dadda_pg_rca32_fa468_y4;
  assign f_s_dadda_pg_rca32_fa491_y4 = f_s_dadda_pg_rca32_fa491_y1 | f_s_dadda_pg_rca32_fa491_y3;
  assign f_s_dadda_pg_rca32_nand_31_8_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_nand_31_8_y0 = ~(f_s_dadda_pg_rca32_nand_31_8_a_31 & f_s_dadda_pg_rca32_nand_31_8_b_8);
  assign f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_fa467_y4 = f_s_dadda_pg_rca32_fa467_y4;
  assign f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_fa466_y4 = f_s_dadda_pg_rca32_fa466_y4;
  assign f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_nand_31_8_y0 = f_s_dadda_pg_rca32_nand_31_8_y0;
  assign f_s_dadda_pg_rca32_fa492_y0 = f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_fa467_y4 ^ f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_fa466_y4;
  assign f_s_dadda_pg_rca32_fa492_y1 = f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_fa467_y4 & f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_fa466_y4;
  assign f_s_dadda_pg_rca32_fa492_y2 = f_s_dadda_pg_rca32_fa492_y0 ^ f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_nand_31_8_y0;
  assign f_s_dadda_pg_rca32_fa492_y3 = f_s_dadda_pg_rca32_fa492_y0 & f_s_dadda_pg_rca32_fa492_f_s_dadda_pg_rca32_nand_31_8_y0;
  assign f_s_dadda_pg_rca32_fa492_y4 = f_s_dadda_pg_rca32_fa492_y1 | f_s_dadda_pg_rca32_fa492_y3;
  assign f_s_dadda_pg_rca32_and_30_9_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_30_9_y0 = f_s_dadda_pg_rca32_and_30_9_a_30 & f_s_dadda_pg_rca32_and_30_9_b_9;
  assign f_s_dadda_pg_rca32_and_29_10_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_29_10_y0 = f_s_dadda_pg_rca32_and_29_10_a_29 & f_s_dadda_pg_rca32_and_29_10_b_10;
  assign f_s_dadda_pg_rca32_and_28_11_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_28_11_y0 = f_s_dadda_pg_rca32_and_28_11_a_28 & f_s_dadda_pg_rca32_and_28_11_b_11;
  assign f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_30_9_y0 = f_s_dadda_pg_rca32_and_30_9_y0;
  assign f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_29_10_y0 = f_s_dadda_pg_rca32_and_29_10_y0;
  assign f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_28_11_y0 = f_s_dadda_pg_rca32_and_28_11_y0;
  assign f_s_dadda_pg_rca32_fa493_y0 = f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_30_9_y0 ^ f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_29_10_y0;
  assign f_s_dadda_pg_rca32_fa493_y1 = f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_30_9_y0 & f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_29_10_y0;
  assign f_s_dadda_pg_rca32_fa493_y2 = f_s_dadda_pg_rca32_fa493_y0 ^ f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_28_11_y0;
  assign f_s_dadda_pg_rca32_fa493_y3 = f_s_dadda_pg_rca32_fa493_y0 & f_s_dadda_pg_rca32_fa493_f_s_dadda_pg_rca32_and_28_11_y0;
  assign f_s_dadda_pg_rca32_fa493_y4 = f_s_dadda_pg_rca32_fa493_y1 | f_s_dadda_pg_rca32_fa493_y3;
  assign f_s_dadda_pg_rca32_and_27_12_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_27_12_y0 = f_s_dadda_pg_rca32_and_27_12_a_27 & f_s_dadda_pg_rca32_and_27_12_b_12;
  assign f_s_dadda_pg_rca32_and_26_13_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_26_13_y0 = f_s_dadda_pg_rca32_and_26_13_a_26 & f_s_dadda_pg_rca32_and_26_13_b_13;
  assign f_s_dadda_pg_rca32_and_25_14_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_25_14_y0 = f_s_dadda_pg_rca32_and_25_14_a_25 & f_s_dadda_pg_rca32_and_25_14_b_14;
  assign f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_27_12_y0 = f_s_dadda_pg_rca32_and_27_12_y0;
  assign f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_26_13_y0 = f_s_dadda_pg_rca32_and_26_13_y0;
  assign f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_25_14_y0 = f_s_dadda_pg_rca32_and_25_14_y0;
  assign f_s_dadda_pg_rca32_fa494_y0 = f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_27_12_y0 ^ f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_26_13_y0;
  assign f_s_dadda_pg_rca32_fa494_y1 = f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_27_12_y0 & f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_26_13_y0;
  assign f_s_dadda_pg_rca32_fa494_y2 = f_s_dadda_pg_rca32_fa494_y0 ^ f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_25_14_y0;
  assign f_s_dadda_pg_rca32_fa494_y3 = f_s_dadda_pg_rca32_fa494_y0 & f_s_dadda_pg_rca32_fa494_f_s_dadda_pg_rca32_and_25_14_y0;
  assign f_s_dadda_pg_rca32_fa494_y4 = f_s_dadda_pg_rca32_fa494_y1 | f_s_dadda_pg_rca32_fa494_y3;
  assign f_s_dadda_pg_rca32_and_24_15_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_24_15_y0 = f_s_dadda_pg_rca32_and_24_15_a_24 & f_s_dadda_pg_rca32_and_24_15_b_15;
  assign f_s_dadda_pg_rca32_and_23_16_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_23_16_y0 = f_s_dadda_pg_rca32_and_23_16_a_23 & f_s_dadda_pg_rca32_and_23_16_b_16;
  assign f_s_dadda_pg_rca32_and_22_17_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_22_17_y0 = f_s_dadda_pg_rca32_and_22_17_a_22 & f_s_dadda_pg_rca32_and_22_17_b_17;
  assign f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_24_15_y0 = f_s_dadda_pg_rca32_and_24_15_y0;
  assign f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_23_16_y0 = f_s_dadda_pg_rca32_and_23_16_y0;
  assign f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_22_17_y0 = f_s_dadda_pg_rca32_and_22_17_y0;
  assign f_s_dadda_pg_rca32_fa495_y0 = f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_24_15_y0 ^ f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_23_16_y0;
  assign f_s_dadda_pg_rca32_fa495_y1 = f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_24_15_y0 & f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_23_16_y0;
  assign f_s_dadda_pg_rca32_fa495_y2 = f_s_dadda_pg_rca32_fa495_y0 ^ f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_22_17_y0;
  assign f_s_dadda_pg_rca32_fa495_y3 = f_s_dadda_pg_rca32_fa495_y0 & f_s_dadda_pg_rca32_fa495_f_s_dadda_pg_rca32_and_22_17_y0;
  assign f_s_dadda_pg_rca32_fa495_y4 = f_s_dadda_pg_rca32_fa495_y1 | f_s_dadda_pg_rca32_fa495_y3;
  assign f_s_dadda_pg_rca32_and_21_18_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_21_18_y0 = f_s_dadda_pg_rca32_and_21_18_a_21 & f_s_dadda_pg_rca32_and_21_18_b_18;
  assign f_s_dadda_pg_rca32_and_20_19_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_20_19_y0 = f_s_dadda_pg_rca32_and_20_19_a_20 & f_s_dadda_pg_rca32_and_20_19_b_19;
  assign f_s_dadda_pg_rca32_and_19_20_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_19_20_y0 = f_s_dadda_pg_rca32_and_19_20_a_19 & f_s_dadda_pg_rca32_and_19_20_b_20;
  assign f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_21_18_y0 = f_s_dadda_pg_rca32_and_21_18_y0;
  assign f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_20_19_y0 = f_s_dadda_pg_rca32_and_20_19_y0;
  assign f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_19_20_y0 = f_s_dadda_pg_rca32_and_19_20_y0;
  assign f_s_dadda_pg_rca32_fa496_y0 = f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_21_18_y0 ^ f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_20_19_y0;
  assign f_s_dadda_pg_rca32_fa496_y1 = f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_21_18_y0 & f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_20_19_y0;
  assign f_s_dadda_pg_rca32_fa496_y2 = f_s_dadda_pg_rca32_fa496_y0 ^ f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_19_20_y0;
  assign f_s_dadda_pg_rca32_fa496_y3 = f_s_dadda_pg_rca32_fa496_y0 & f_s_dadda_pg_rca32_fa496_f_s_dadda_pg_rca32_and_19_20_y0;
  assign f_s_dadda_pg_rca32_fa496_y4 = f_s_dadda_pg_rca32_fa496_y1 | f_s_dadda_pg_rca32_fa496_y3;
  assign f_s_dadda_pg_rca32_and_18_21_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_18_21_y0 = f_s_dadda_pg_rca32_and_18_21_a_18 & f_s_dadda_pg_rca32_and_18_21_b_21;
  assign f_s_dadda_pg_rca32_and_17_22_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_17_22_y0 = f_s_dadda_pg_rca32_and_17_22_a_17 & f_s_dadda_pg_rca32_and_17_22_b_22;
  assign f_s_dadda_pg_rca32_and_16_23_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_16_23_y0 = f_s_dadda_pg_rca32_and_16_23_a_16 & f_s_dadda_pg_rca32_and_16_23_b_23;
  assign f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_18_21_y0 = f_s_dadda_pg_rca32_and_18_21_y0;
  assign f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_17_22_y0 = f_s_dadda_pg_rca32_and_17_22_y0;
  assign f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_16_23_y0 = f_s_dadda_pg_rca32_and_16_23_y0;
  assign f_s_dadda_pg_rca32_fa497_y0 = f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_18_21_y0 ^ f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_17_22_y0;
  assign f_s_dadda_pg_rca32_fa497_y1 = f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_18_21_y0 & f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_17_22_y0;
  assign f_s_dadda_pg_rca32_fa497_y2 = f_s_dadda_pg_rca32_fa497_y0 ^ f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_16_23_y0;
  assign f_s_dadda_pg_rca32_fa497_y3 = f_s_dadda_pg_rca32_fa497_y0 & f_s_dadda_pg_rca32_fa497_f_s_dadda_pg_rca32_and_16_23_y0;
  assign f_s_dadda_pg_rca32_fa497_y4 = f_s_dadda_pg_rca32_fa497_y1 | f_s_dadda_pg_rca32_fa497_y3;
  assign f_s_dadda_pg_rca32_and_15_24_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_15_24_y0 = f_s_dadda_pg_rca32_and_15_24_a_15 & f_s_dadda_pg_rca32_and_15_24_b_24;
  assign f_s_dadda_pg_rca32_and_14_25_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_14_25_y0 = f_s_dadda_pg_rca32_and_14_25_a_14 & f_s_dadda_pg_rca32_and_14_25_b_25;
  assign f_s_dadda_pg_rca32_and_13_26_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_13_26_y0 = f_s_dadda_pg_rca32_and_13_26_a_13 & f_s_dadda_pg_rca32_and_13_26_b_26;
  assign f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_15_24_y0 = f_s_dadda_pg_rca32_and_15_24_y0;
  assign f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_14_25_y0 = f_s_dadda_pg_rca32_and_14_25_y0;
  assign f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_13_26_y0 = f_s_dadda_pg_rca32_and_13_26_y0;
  assign f_s_dadda_pg_rca32_fa498_y0 = f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_15_24_y0 ^ f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_14_25_y0;
  assign f_s_dadda_pg_rca32_fa498_y1 = f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_15_24_y0 & f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_14_25_y0;
  assign f_s_dadda_pg_rca32_fa498_y2 = f_s_dadda_pg_rca32_fa498_y0 ^ f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_13_26_y0;
  assign f_s_dadda_pg_rca32_fa498_y3 = f_s_dadda_pg_rca32_fa498_y0 & f_s_dadda_pg_rca32_fa498_f_s_dadda_pg_rca32_and_13_26_y0;
  assign f_s_dadda_pg_rca32_fa498_y4 = f_s_dadda_pg_rca32_fa498_y1 | f_s_dadda_pg_rca32_fa498_y3;
  assign f_s_dadda_pg_rca32_and_12_27_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_12_27_y0 = f_s_dadda_pg_rca32_and_12_27_a_12 & f_s_dadda_pg_rca32_and_12_27_b_27;
  assign f_s_dadda_pg_rca32_and_11_28_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_11_28_y0 = f_s_dadda_pg_rca32_and_11_28_a_11 & f_s_dadda_pg_rca32_and_11_28_b_28;
  assign f_s_dadda_pg_rca32_and_10_29_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_10_29_y0 = f_s_dadda_pg_rca32_and_10_29_a_10 & f_s_dadda_pg_rca32_and_10_29_b_29;
  assign f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_12_27_y0 = f_s_dadda_pg_rca32_and_12_27_y0;
  assign f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_11_28_y0 = f_s_dadda_pg_rca32_and_11_28_y0;
  assign f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_10_29_y0 = f_s_dadda_pg_rca32_and_10_29_y0;
  assign f_s_dadda_pg_rca32_fa499_y0 = f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_12_27_y0 ^ f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_11_28_y0;
  assign f_s_dadda_pg_rca32_fa499_y1 = f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_12_27_y0 & f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_11_28_y0;
  assign f_s_dadda_pg_rca32_fa499_y2 = f_s_dadda_pg_rca32_fa499_y0 ^ f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_10_29_y0;
  assign f_s_dadda_pg_rca32_fa499_y3 = f_s_dadda_pg_rca32_fa499_y0 & f_s_dadda_pg_rca32_fa499_f_s_dadda_pg_rca32_and_10_29_y0;
  assign f_s_dadda_pg_rca32_fa499_y4 = f_s_dadda_pg_rca32_fa499_y1 | f_s_dadda_pg_rca32_fa499_y3;
  assign f_s_dadda_pg_rca32_and_9_30_a_9 = a_9;
  assign f_s_dadda_pg_rca32_and_9_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_9_30_y0 = f_s_dadda_pg_rca32_and_9_30_a_9 & f_s_dadda_pg_rca32_and_9_30_b_30;
  assign f_s_dadda_pg_rca32_nand_8_31_a_8 = a_8;
  assign f_s_dadda_pg_rca32_nand_8_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_8_31_y0 = ~(f_s_dadda_pg_rca32_nand_8_31_a_8 & f_s_dadda_pg_rca32_nand_8_31_b_31);
  assign f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_and_9_30_y0 = f_s_dadda_pg_rca32_and_9_30_y0;
  assign f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_nand_8_31_y0 = f_s_dadda_pg_rca32_nand_8_31_y0;
  assign f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_fa486_y2 = f_s_dadda_pg_rca32_fa486_y2;
  assign f_s_dadda_pg_rca32_fa500_y0 = f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_and_9_30_y0 ^ f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_nand_8_31_y0;
  assign f_s_dadda_pg_rca32_fa500_y1 = f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_and_9_30_y0 & f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_nand_8_31_y0;
  assign f_s_dadda_pg_rca32_fa500_y2 = f_s_dadda_pg_rca32_fa500_y0 ^ f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_fa486_y2;
  assign f_s_dadda_pg_rca32_fa500_y3 = f_s_dadda_pg_rca32_fa500_y0 & f_s_dadda_pg_rca32_fa500_f_s_dadda_pg_rca32_fa486_y2;
  assign f_s_dadda_pg_rca32_fa500_y4 = f_s_dadda_pg_rca32_fa500_y1 | f_s_dadda_pg_rca32_fa500_y3;
  assign f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa487_y2 = f_s_dadda_pg_rca32_fa487_y2;
  assign f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa488_y2 = f_s_dadda_pg_rca32_fa488_y2;
  assign f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa489_y2 = f_s_dadda_pg_rca32_fa489_y2;
  assign f_s_dadda_pg_rca32_fa501_y0 = f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa487_y2 ^ f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa488_y2;
  assign f_s_dadda_pg_rca32_fa501_y1 = f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa487_y2 & f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa488_y2;
  assign f_s_dadda_pg_rca32_fa501_y2 = f_s_dadda_pg_rca32_fa501_y0 ^ f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa489_y2;
  assign f_s_dadda_pg_rca32_fa501_y3 = f_s_dadda_pg_rca32_fa501_y0 & f_s_dadda_pg_rca32_fa501_f_s_dadda_pg_rca32_fa489_y2;
  assign f_s_dadda_pg_rca32_fa501_y4 = f_s_dadda_pg_rca32_fa501_y1 | f_s_dadda_pg_rca32_fa501_y3;
  assign f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa490_y2 = f_s_dadda_pg_rca32_fa490_y2;
  assign f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa491_y2 = f_s_dadda_pg_rca32_fa491_y2;
  assign f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa492_y2 = f_s_dadda_pg_rca32_fa492_y2;
  assign f_s_dadda_pg_rca32_fa502_y0 = f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa490_y2 ^ f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa491_y2;
  assign f_s_dadda_pg_rca32_fa502_y1 = f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa490_y2 & f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa491_y2;
  assign f_s_dadda_pg_rca32_fa502_y2 = f_s_dadda_pg_rca32_fa502_y0 ^ f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa492_y2;
  assign f_s_dadda_pg_rca32_fa502_y3 = f_s_dadda_pg_rca32_fa502_y0 & f_s_dadda_pg_rca32_fa502_f_s_dadda_pg_rca32_fa492_y2;
  assign f_s_dadda_pg_rca32_fa502_y4 = f_s_dadda_pg_rca32_fa502_y1 | f_s_dadda_pg_rca32_fa502_y3;
  assign f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa493_y2 = f_s_dadda_pg_rca32_fa493_y2;
  assign f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa494_y2 = f_s_dadda_pg_rca32_fa494_y2;
  assign f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa495_y2 = f_s_dadda_pg_rca32_fa495_y2;
  assign f_s_dadda_pg_rca32_fa503_y0 = f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa493_y2 ^ f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa494_y2;
  assign f_s_dadda_pg_rca32_fa503_y1 = f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa493_y2 & f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa494_y2;
  assign f_s_dadda_pg_rca32_fa503_y2 = f_s_dadda_pg_rca32_fa503_y0 ^ f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa495_y2;
  assign f_s_dadda_pg_rca32_fa503_y3 = f_s_dadda_pg_rca32_fa503_y0 & f_s_dadda_pg_rca32_fa503_f_s_dadda_pg_rca32_fa495_y2;
  assign f_s_dadda_pg_rca32_fa503_y4 = f_s_dadda_pg_rca32_fa503_y1 | f_s_dadda_pg_rca32_fa503_y3;
  assign f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa496_y2 = f_s_dadda_pg_rca32_fa496_y2;
  assign f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa497_y2 = f_s_dadda_pg_rca32_fa497_y2;
  assign f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa498_y2 = f_s_dadda_pg_rca32_fa498_y2;
  assign f_s_dadda_pg_rca32_fa504_y0 = f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa496_y2 ^ f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa497_y2;
  assign f_s_dadda_pg_rca32_fa504_y1 = f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa496_y2 & f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa497_y2;
  assign f_s_dadda_pg_rca32_fa504_y2 = f_s_dadda_pg_rca32_fa504_y0 ^ f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa498_y2;
  assign f_s_dadda_pg_rca32_fa504_y3 = f_s_dadda_pg_rca32_fa504_y0 & f_s_dadda_pg_rca32_fa504_f_s_dadda_pg_rca32_fa498_y2;
  assign f_s_dadda_pg_rca32_fa504_y4 = f_s_dadda_pg_rca32_fa504_y1 | f_s_dadda_pg_rca32_fa504_y3;
  assign f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa504_y4 = f_s_dadda_pg_rca32_fa504_y4;
  assign f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa503_y4 = f_s_dadda_pg_rca32_fa503_y4;
  assign f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa502_y4 = f_s_dadda_pg_rca32_fa502_y4;
  assign f_s_dadda_pg_rca32_fa505_y0 = f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa504_y4 ^ f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa503_y4;
  assign f_s_dadda_pg_rca32_fa505_y1 = f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa504_y4 & f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa503_y4;
  assign f_s_dadda_pg_rca32_fa505_y2 = f_s_dadda_pg_rca32_fa505_y0 ^ f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa502_y4;
  assign f_s_dadda_pg_rca32_fa505_y3 = f_s_dadda_pg_rca32_fa505_y0 & f_s_dadda_pg_rca32_fa505_f_s_dadda_pg_rca32_fa502_y4;
  assign f_s_dadda_pg_rca32_fa505_y4 = f_s_dadda_pg_rca32_fa505_y1 | f_s_dadda_pg_rca32_fa505_y3;
  assign f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa501_y4 = f_s_dadda_pg_rca32_fa501_y4;
  assign f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa500_y4 = f_s_dadda_pg_rca32_fa500_y4;
  assign f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa499_y4 = f_s_dadda_pg_rca32_fa499_y4;
  assign f_s_dadda_pg_rca32_fa506_y0 = f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa501_y4 ^ f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa500_y4;
  assign f_s_dadda_pg_rca32_fa506_y1 = f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa501_y4 & f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa500_y4;
  assign f_s_dadda_pg_rca32_fa506_y2 = f_s_dadda_pg_rca32_fa506_y0 ^ f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa499_y4;
  assign f_s_dadda_pg_rca32_fa506_y3 = f_s_dadda_pg_rca32_fa506_y0 & f_s_dadda_pg_rca32_fa506_f_s_dadda_pg_rca32_fa499_y4;
  assign f_s_dadda_pg_rca32_fa506_y4 = f_s_dadda_pg_rca32_fa506_y1 | f_s_dadda_pg_rca32_fa506_y3;
  assign f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa498_y4 = f_s_dadda_pg_rca32_fa498_y4;
  assign f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa497_y4 = f_s_dadda_pg_rca32_fa497_y4;
  assign f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa496_y4 = f_s_dadda_pg_rca32_fa496_y4;
  assign f_s_dadda_pg_rca32_fa507_y0 = f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa498_y4 ^ f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa497_y4;
  assign f_s_dadda_pg_rca32_fa507_y1 = f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa498_y4 & f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa497_y4;
  assign f_s_dadda_pg_rca32_fa507_y2 = f_s_dadda_pg_rca32_fa507_y0 ^ f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa496_y4;
  assign f_s_dadda_pg_rca32_fa507_y3 = f_s_dadda_pg_rca32_fa507_y0 & f_s_dadda_pg_rca32_fa507_f_s_dadda_pg_rca32_fa496_y4;
  assign f_s_dadda_pg_rca32_fa507_y4 = f_s_dadda_pg_rca32_fa507_y1 | f_s_dadda_pg_rca32_fa507_y3;
  assign f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa495_y4 = f_s_dadda_pg_rca32_fa495_y4;
  assign f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa494_y4 = f_s_dadda_pg_rca32_fa494_y4;
  assign f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa493_y4 = f_s_dadda_pg_rca32_fa493_y4;
  assign f_s_dadda_pg_rca32_fa508_y0 = f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa495_y4 ^ f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa494_y4;
  assign f_s_dadda_pg_rca32_fa508_y1 = f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa495_y4 & f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa494_y4;
  assign f_s_dadda_pg_rca32_fa508_y2 = f_s_dadda_pg_rca32_fa508_y0 ^ f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa493_y4;
  assign f_s_dadda_pg_rca32_fa508_y3 = f_s_dadda_pg_rca32_fa508_y0 & f_s_dadda_pg_rca32_fa508_f_s_dadda_pg_rca32_fa493_y4;
  assign f_s_dadda_pg_rca32_fa508_y4 = f_s_dadda_pg_rca32_fa508_y1 | f_s_dadda_pg_rca32_fa508_y3;
  assign f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa492_y4 = f_s_dadda_pg_rca32_fa492_y4;
  assign f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa491_y4 = f_s_dadda_pg_rca32_fa491_y4;
  assign f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa490_y4 = f_s_dadda_pg_rca32_fa490_y4;
  assign f_s_dadda_pg_rca32_fa509_y0 = f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa492_y4 ^ f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa491_y4;
  assign f_s_dadda_pg_rca32_fa509_y1 = f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa492_y4 & f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa491_y4;
  assign f_s_dadda_pg_rca32_fa509_y2 = f_s_dadda_pg_rca32_fa509_y0 ^ f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa490_y4;
  assign f_s_dadda_pg_rca32_fa509_y3 = f_s_dadda_pg_rca32_fa509_y0 & f_s_dadda_pg_rca32_fa509_f_s_dadda_pg_rca32_fa490_y4;
  assign f_s_dadda_pg_rca32_fa509_y4 = f_s_dadda_pg_rca32_fa509_y1 | f_s_dadda_pg_rca32_fa509_y3;
  assign f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa489_y4 = f_s_dadda_pg_rca32_fa489_y4;
  assign f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa488_y4 = f_s_dadda_pg_rca32_fa488_y4;
  assign f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa487_y4 = f_s_dadda_pg_rca32_fa487_y4;
  assign f_s_dadda_pg_rca32_fa510_y0 = f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa489_y4 ^ f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa488_y4;
  assign f_s_dadda_pg_rca32_fa510_y1 = f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa489_y4 & f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa488_y4;
  assign f_s_dadda_pg_rca32_fa510_y2 = f_s_dadda_pg_rca32_fa510_y0 ^ f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa487_y4;
  assign f_s_dadda_pg_rca32_fa510_y3 = f_s_dadda_pg_rca32_fa510_y0 & f_s_dadda_pg_rca32_fa510_f_s_dadda_pg_rca32_fa487_y4;
  assign f_s_dadda_pg_rca32_fa510_y4 = f_s_dadda_pg_rca32_fa510_y1 | f_s_dadda_pg_rca32_fa510_y3;
  assign f_s_dadda_pg_rca32_nand_31_9_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_nand_31_9_y0 = ~(f_s_dadda_pg_rca32_nand_31_9_a_31 & f_s_dadda_pg_rca32_nand_31_9_b_9);
  assign f_s_dadda_pg_rca32_and_30_10_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_30_10_y0 = f_s_dadda_pg_rca32_and_30_10_a_30 & f_s_dadda_pg_rca32_and_30_10_b_10;
  assign f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_fa486_y4 = f_s_dadda_pg_rca32_fa486_y4;
  assign f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_nand_31_9_y0 = f_s_dadda_pg_rca32_nand_31_9_y0;
  assign f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_and_30_10_y0 = f_s_dadda_pg_rca32_and_30_10_y0;
  assign f_s_dadda_pg_rca32_fa511_y0 = f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_fa486_y4 ^ f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_nand_31_9_y0;
  assign f_s_dadda_pg_rca32_fa511_y1 = f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_fa486_y4 & f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_nand_31_9_y0;
  assign f_s_dadda_pg_rca32_fa511_y2 = f_s_dadda_pg_rca32_fa511_y0 ^ f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_and_30_10_y0;
  assign f_s_dadda_pg_rca32_fa511_y3 = f_s_dadda_pg_rca32_fa511_y0 & f_s_dadda_pg_rca32_fa511_f_s_dadda_pg_rca32_and_30_10_y0;
  assign f_s_dadda_pg_rca32_fa511_y4 = f_s_dadda_pg_rca32_fa511_y1 | f_s_dadda_pg_rca32_fa511_y3;
  assign f_s_dadda_pg_rca32_and_29_11_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_29_11_y0 = f_s_dadda_pg_rca32_and_29_11_a_29 & f_s_dadda_pg_rca32_and_29_11_b_11;
  assign f_s_dadda_pg_rca32_and_28_12_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_28_12_y0 = f_s_dadda_pg_rca32_and_28_12_a_28 & f_s_dadda_pg_rca32_and_28_12_b_12;
  assign f_s_dadda_pg_rca32_and_27_13_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_27_13_y0 = f_s_dadda_pg_rca32_and_27_13_a_27 & f_s_dadda_pg_rca32_and_27_13_b_13;
  assign f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_29_11_y0 = f_s_dadda_pg_rca32_and_29_11_y0;
  assign f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_28_12_y0 = f_s_dadda_pg_rca32_and_28_12_y0;
  assign f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_27_13_y0 = f_s_dadda_pg_rca32_and_27_13_y0;
  assign f_s_dadda_pg_rca32_fa512_y0 = f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_29_11_y0 ^ f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_28_12_y0;
  assign f_s_dadda_pg_rca32_fa512_y1 = f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_29_11_y0 & f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_28_12_y0;
  assign f_s_dadda_pg_rca32_fa512_y2 = f_s_dadda_pg_rca32_fa512_y0 ^ f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_27_13_y0;
  assign f_s_dadda_pg_rca32_fa512_y3 = f_s_dadda_pg_rca32_fa512_y0 & f_s_dadda_pg_rca32_fa512_f_s_dadda_pg_rca32_and_27_13_y0;
  assign f_s_dadda_pg_rca32_fa512_y4 = f_s_dadda_pg_rca32_fa512_y1 | f_s_dadda_pg_rca32_fa512_y3;
  assign f_s_dadda_pg_rca32_and_26_14_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_26_14_y0 = f_s_dadda_pg_rca32_and_26_14_a_26 & f_s_dadda_pg_rca32_and_26_14_b_14;
  assign f_s_dadda_pg_rca32_and_25_15_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_25_15_y0 = f_s_dadda_pg_rca32_and_25_15_a_25 & f_s_dadda_pg_rca32_and_25_15_b_15;
  assign f_s_dadda_pg_rca32_and_24_16_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_24_16_y0 = f_s_dadda_pg_rca32_and_24_16_a_24 & f_s_dadda_pg_rca32_and_24_16_b_16;
  assign f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_26_14_y0 = f_s_dadda_pg_rca32_and_26_14_y0;
  assign f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_25_15_y0 = f_s_dadda_pg_rca32_and_25_15_y0;
  assign f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_24_16_y0 = f_s_dadda_pg_rca32_and_24_16_y0;
  assign f_s_dadda_pg_rca32_fa513_y0 = f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_26_14_y0 ^ f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_25_15_y0;
  assign f_s_dadda_pg_rca32_fa513_y1 = f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_26_14_y0 & f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_25_15_y0;
  assign f_s_dadda_pg_rca32_fa513_y2 = f_s_dadda_pg_rca32_fa513_y0 ^ f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_24_16_y0;
  assign f_s_dadda_pg_rca32_fa513_y3 = f_s_dadda_pg_rca32_fa513_y0 & f_s_dadda_pg_rca32_fa513_f_s_dadda_pg_rca32_and_24_16_y0;
  assign f_s_dadda_pg_rca32_fa513_y4 = f_s_dadda_pg_rca32_fa513_y1 | f_s_dadda_pg_rca32_fa513_y3;
  assign f_s_dadda_pg_rca32_and_23_17_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_23_17_y0 = f_s_dadda_pg_rca32_and_23_17_a_23 & f_s_dadda_pg_rca32_and_23_17_b_17;
  assign f_s_dadda_pg_rca32_and_22_18_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_22_18_y0 = f_s_dadda_pg_rca32_and_22_18_a_22 & f_s_dadda_pg_rca32_and_22_18_b_18;
  assign f_s_dadda_pg_rca32_and_21_19_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_21_19_y0 = f_s_dadda_pg_rca32_and_21_19_a_21 & f_s_dadda_pg_rca32_and_21_19_b_19;
  assign f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_23_17_y0 = f_s_dadda_pg_rca32_and_23_17_y0;
  assign f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_22_18_y0 = f_s_dadda_pg_rca32_and_22_18_y0;
  assign f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_21_19_y0 = f_s_dadda_pg_rca32_and_21_19_y0;
  assign f_s_dadda_pg_rca32_fa514_y0 = f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_23_17_y0 ^ f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_22_18_y0;
  assign f_s_dadda_pg_rca32_fa514_y1 = f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_23_17_y0 & f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_22_18_y0;
  assign f_s_dadda_pg_rca32_fa514_y2 = f_s_dadda_pg_rca32_fa514_y0 ^ f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_21_19_y0;
  assign f_s_dadda_pg_rca32_fa514_y3 = f_s_dadda_pg_rca32_fa514_y0 & f_s_dadda_pg_rca32_fa514_f_s_dadda_pg_rca32_and_21_19_y0;
  assign f_s_dadda_pg_rca32_fa514_y4 = f_s_dadda_pg_rca32_fa514_y1 | f_s_dadda_pg_rca32_fa514_y3;
  assign f_s_dadda_pg_rca32_and_20_20_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_20_20_y0 = f_s_dadda_pg_rca32_and_20_20_a_20 & f_s_dadda_pg_rca32_and_20_20_b_20;
  assign f_s_dadda_pg_rca32_and_19_21_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_19_21_y0 = f_s_dadda_pg_rca32_and_19_21_a_19 & f_s_dadda_pg_rca32_and_19_21_b_21;
  assign f_s_dadda_pg_rca32_and_18_22_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_18_22_y0 = f_s_dadda_pg_rca32_and_18_22_a_18 & f_s_dadda_pg_rca32_and_18_22_b_22;
  assign f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_20_20_y0 = f_s_dadda_pg_rca32_and_20_20_y0;
  assign f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_19_21_y0 = f_s_dadda_pg_rca32_and_19_21_y0;
  assign f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_18_22_y0 = f_s_dadda_pg_rca32_and_18_22_y0;
  assign f_s_dadda_pg_rca32_fa515_y0 = f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_20_20_y0 ^ f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_19_21_y0;
  assign f_s_dadda_pg_rca32_fa515_y1 = f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_20_20_y0 & f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_19_21_y0;
  assign f_s_dadda_pg_rca32_fa515_y2 = f_s_dadda_pg_rca32_fa515_y0 ^ f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_18_22_y0;
  assign f_s_dadda_pg_rca32_fa515_y3 = f_s_dadda_pg_rca32_fa515_y0 & f_s_dadda_pg_rca32_fa515_f_s_dadda_pg_rca32_and_18_22_y0;
  assign f_s_dadda_pg_rca32_fa515_y4 = f_s_dadda_pg_rca32_fa515_y1 | f_s_dadda_pg_rca32_fa515_y3;
  assign f_s_dadda_pg_rca32_and_17_23_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_17_23_y0 = f_s_dadda_pg_rca32_and_17_23_a_17 & f_s_dadda_pg_rca32_and_17_23_b_23;
  assign f_s_dadda_pg_rca32_and_16_24_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_16_24_y0 = f_s_dadda_pg_rca32_and_16_24_a_16 & f_s_dadda_pg_rca32_and_16_24_b_24;
  assign f_s_dadda_pg_rca32_and_15_25_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_15_25_y0 = f_s_dadda_pg_rca32_and_15_25_a_15 & f_s_dadda_pg_rca32_and_15_25_b_25;
  assign f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_17_23_y0 = f_s_dadda_pg_rca32_and_17_23_y0;
  assign f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_16_24_y0 = f_s_dadda_pg_rca32_and_16_24_y0;
  assign f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_15_25_y0 = f_s_dadda_pg_rca32_and_15_25_y0;
  assign f_s_dadda_pg_rca32_fa516_y0 = f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_17_23_y0 ^ f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_16_24_y0;
  assign f_s_dadda_pg_rca32_fa516_y1 = f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_17_23_y0 & f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_16_24_y0;
  assign f_s_dadda_pg_rca32_fa516_y2 = f_s_dadda_pg_rca32_fa516_y0 ^ f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_15_25_y0;
  assign f_s_dadda_pg_rca32_fa516_y3 = f_s_dadda_pg_rca32_fa516_y0 & f_s_dadda_pg_rca32_fa516_f_s_dadda_pg_rca32_and_15_25_y0;
  assign f_s_dadda_pg_rca32_fa516_y4 = f_s_dadda_pg_rca32_fa516_y1 | f_s_dadda_pg_rca32_fa516_y3;
  assign f_s_dadda_pg_rca32_and_14_26_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_14_26_y0 = f_s_dadda_pg_rca32_and_14_26_a_14 & f_s_dadda_pg_rca32_and_14_26_b_26;
  assign f_s_dadda_pg_rca32_and_13_27_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_13_27_y0 = f_s_dadda_pg_rca32_and_13_27_a_13 & f_s_dadda_pg_rca32_and_13_27_b_27;
  assign f_s_dadda_pg_rca32_and_12_28_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_12_28_y0 = f_s_dadda_pg_rca32_and_12_28_a_12 & f_s_dadda_pg_rca32_and_12_28_b_28;
  assign f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_14_26_y0 = f_s_dadda_pg_rca32_and_14_26_y0;
  assign f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_13_27_y0 = f_s_dadda_pg_rca32_and_13_27_y0;
  assign f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_12_28_y0 = f_s_dadda_pg_rca32_and_12_28_y0;
  assign f_s_dadda_pg_rca32_fa517_y0 = f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_14_26_y0 ^ f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_13_27_y0;
  assign f_s_dadda_pg_rca32_fa517_y1 = f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_14_26_y0 & f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_13_27_y0;
  assign f_s_dadda_pg_rca32_fa517_y2 = f_s_dadda_pg_rca32_fa517_y0 ^ f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_12_28_y0;
  assign f_s_dadda_pg_rca32_fa517_y3 = f_s_dadda_pg_rca32_fa517_y0 & f_s_dadda_pg_rca32_fa517_f_s_dadda_pg_rca32_and_12_28_y0;
  assign f_s_dadda_pg_rca32_fa517_y4 = f_s_dadda_pg_rca32_fa517_y1 | f_s_dadda_pg_rca32_fa517_y3;
  assign f_s_dadda_pg_rca32_and_11_29_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_11_29_y0 = f_s_dadda_pg_rca32_and_11_29_a_11 & f_s_dadda_pg_rca32_and_11_29_b_29;
  assign f_s_dadda_pg_rca32_and_10_30_a_10 = a_10;
  assign f_s_dadda_pg_rca32_and_10_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_10_30_y0 = f_s_dadda_pg_rca32_and_10_30_a_10 & f_s_dadda_pg_rca32_and_10_30_b_30;
  assign f_s_dadda_pg_rca32_nand_9_31_a_9 = a_9;
  assign f_s_dadda_pg_rca32_nand_9_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_9_31_y0 = ~(f_s_dadda_pg_rca32_nand_9_31_a_9 & f_s_dadda_pg_rca32_nand_9_31_b_31);
  assign f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_and_11_29_y0 = f_s_dadda_pg_rca32_and_11_29_y0;
  assign f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_and_10_30_y0 = f_s_dadda_pg_rca32_and_10_30_y0;
  assign f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_nand_9_31_y0 = f_s_dadda_pg_rca32_nand_9_31_y0;
  assign f_s_dadda_pg_rca32_fa518_y0 = f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_and_11_29_y0 ^ f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_and_10_30_y0;
  assign f_s_dadda_pg_rca32_fa518_y1 = f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_and_11_29_y0 & f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_and_10_30_y0;
  assign f_s_dadda_pg_rca32_fa518_y2 = f_s_dadda_pg_rca32_fa518_y0 ^ f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_nand_9_31_y0;
  assign f_s_dadda_pg_rca32_fa518_y3 = f_s_dadda_pg_rca32_fa518_y0 & f_s_dadda_pg_rca32_fa518_f_s_dadda_pg_rca32_nand_9_31_y0;
  assign f_s_dadda_pg_rca32_fa518_y4 = f_s_dadda_pg_rca32_fa518_y1 | f_s_dadda_pg_rca32_fa518_y3;
  assign f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa505_y2 = f_s_dadda_pg_rca32_fa505_y2;
  assign f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa506_y2 = f_s_dadda_pg_rca32_fa506_y2;
  assign f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa507_y2 = f_s_dadda_pg_rca32_fa507_y2;
  assign f_s_dadda_pg_rca32_fa519_y0 = f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa505_y2 ^ f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa506_y2;
  assign f_s_dadda_pg_rca32_fa519_y1 = f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa505_y2 & f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa506_y2;
  assign f_s_dadda_pg_rca32_fa519_y2 = f_s_dadda_pg_rca32_fa519_y0 ^ f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa507_y2;
  assign f_s_dadda_pg_rca32_fa519_y3 = f_s_dadda_pg_rca32_fa519_y0 & f_s_dadda_pg_rca32_fa519_f_s_dadda_pg_rca32_fa507_y2;
  assign f_s_dadda_pg_rca32_fa519_y4 = f_s_dadda_pg_rca32_fa519_y1 | f_s_dadda_pg_rca32_fa519_y3;
  assign f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa508_y2 = f_s_dadda_pg_rca32_fa508_y2;
  assign f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa509_y2 = f_s_dadda_pg_rca32_fa509_y2;
  assign f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa510_y2 = f_s_dadda_pg_rca32_fa510_y2;
  assign f_s_dadda_pg_rca32_fa520_y0 = f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa508_y2 ^ f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa509_y2;
  assign f_s_dadda_pg_rca32_fa520_y1 = f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa508_y2 & f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa509_y2;
  assign f_s_dadda_pg_rca32_fa520_y2 = f_s_dadda_pg_rca32_fa520_y0 ^ f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa510_y2;
  assign f_s_dadda_pg_rca32_fa520_y3 = f_s_dadda_pg_rca32_fa520_y0 & f_s_dadda_pg_rca32_fa520_f_s_dadda_pg_rca32_fa510_y2;
  assign f_s_dadda_pg_rca32_fa520_y4 = f_s_dadda_pg_rca32_fa520_y1 | f_s_dadda_pg_rca32_fa520_y3;
  assign f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa511_y2 = f_s_dadda_pg_rca32_fa511_y2;
  assign f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa512_y2 = f_s_dadda_pg_rca32_fa512_y2;
  assign f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa513_y2 = f_s_dadda_pg_rca32_fa513_y2;
  assign f_s_dadda_pg_rca32_fa521_y0 = f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa511_y2 ^ f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa512_y2;
  assign f_s_dadda_pg_rca32_fa521_y1 = f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa511_y2 & f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa512_y2;
  assign f_s_dadda_pg_rca32_fa521_y2 = f_s_dadda_pg_rca32_fa521_y0 ^ f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa513_y2;
  assign f_s_dadda_pg_rca32_fa521_y3 = f_s_dadda_pg_rca32_fa521_y0 & f_s_dadda_pg_rca32_fa521_f_s_dadda_pg_rca32_fa513_y2;
  assign f_s_dadda_pg_rca32_fa521_y4 = f_s_dadda_pg_rca32_fa521_y1 | f_s_dadda_pg_rca32_fa521_y3;
  assign f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa514_y2 = f_s_dadda_pg_rca32_fa514_y2;
  assign f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa515_y2 = f_s_dadda_pg_rca32_fa515_y2;
  assign f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa516_y2 = f_s_dadda_pg_rca32_fa516_y2;
  assign f_s_dadda_pg_rca32_fa522_y0 = f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa514_y2 ^ f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa515_y2;
  assign f_s_dadda_pg_rca32_fa522_y1 = f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa514_y2 & f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa515_y2;
  assign f_s_dadda_pg_rca32_fa522_y2 = f_s_dadda_pg_rca32_fa522_y0 ^ f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa516_y2;
  assign f_s_dadda_pg_rca32_fa522_y3 = f_s_dadda_pg_rca32_fa522_y0 & f_s_dadda_pg_rca32_fa522_f_s_dadda_pg_rca32_fa516_y2;
  assign f_s_dadda_pg_rca32_fa522_y4 = f_s_dadda_pg_rca32_fa522_y1 | f_s_dadda_pg_rca32_fa522_y3;
  assign f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa522_y4 = f_s_dadda_pg_rca32_fa522_y4;
  assign f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa521_y4 = f_s_dadda_pg_rca32_fa521_y4;
  assign f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa520_y4 = f_s_dadda_pg_rca32_fa520_y4;
  assign f_s_dadda_pg_rca32_fa523_y0 = f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa522_y4 ^ f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa521_y4;
  assign f_s_dadda_pg_rca32_fa523_y1 = f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa522_y4 & f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa521_y4;
  assign f_s_dadda_pg_rca32_fa523_y2 = f_s_dadda_pg_rca32_fa523_y0 ^ f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa520_y4;
  assign f_s_dadda_pg_rca32_fa523_y3 = f_s_dadda_pg_rca32_fa523_y0 & f_s_dadda_pg_rca32_fa523_f_s_dadda_pg_rca32_fa520_y4;
  assign f_s_dadda_pg_rca32_fa523_y4 = f_s_dadda_pg_rca32_fa523_y1 | f_s_dadda_pg_rca32_fa523_y3;
  assign f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa519_y4 = f_s_dadda_pg_rca32_fa519_y4;
  assign f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa518_y4 = f_s_dadda_pg_rca32_fa518_y4;
  assign f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa517_y4 = f_s_dadda_pg_rca32_fa517_y4;
  assign f_s_dadda_pg_rca32_fa524_y0 = f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa519_y4 ^ f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa518_y4;
  assign f_s_dadda_pg_rca32_fa524_y1 = f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa519_y4 & f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa518_y4;
  assign f_s_dadda_pg_rca32_fa524_y2 = f_s_dadda_pg_rca32_fa524_y0 ^ f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa517_y4;
  assign f_s_dadda_pg_rca32_fa524_y3 = f_s_dadda_pg_rca32_fa524_y0 & f_s_dadda_pg_rca32_fa524_f_s_dadda_pg_rca32_fa517_y4;
  assign f_s_dadda_pg_rca32_fa524_y4 = f_s_dadda_pg_rca32_fa524_y1 | f_s_dadda_pg_rca32_fa524_y3;
  assign f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa516_y4 = f_s_dadda_pg_rca32_fa516_y4;
  assign f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa515_y4 = f_s_dadda_pg_rca32_fa515_y4;
  assign f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa514_y4 = f_s_dadda_pg_rca32_fa514_y4;
  assign f_s_dadda_pg_rca32_fa525_y0 = f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa516_y4 ^ f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa515_y4;
  assign f_s_dadda_pg_rca32_fa525_y1 = f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa516_y4 & f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa515_y4;
  assign f_s_dadda_pg_rca32_fa525_y2 = f_s_dadda_pg_rca32_fa525_y0 ^ f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa514_y4;
  assign f_s_dadda_pg_rca32_fa525_y3 = f_s_dadda_pg_rca32_fa525_y0 & f_s_dadda_pg_rca32_fa525_f_s_dadda_pg_rca32_fa514_y4;
  assign f_s_dadda_pg_rca32_fa525_y4 = f_s_dadda_pg_rca32_fa525_y1 | f_s_dadda_pg_rca32_fa525_y3;
  assign f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa513_y4 = f_s_dadda_pg_rca32_fa513_y4;
  assign f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa512_y4 = f_s_dadda_pg_rca32_fa512_y4;
  assign f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa511_y4 = f_s_dadda_pg_rca32_fa511_y4;
  assign f_s_dadda_pg_rca32_fa526_y0 = f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa513_y4 ^ f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa512_y4;
  assign f_s_dadda_pg_rca32_fa526_y1 = f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa513_y4 & f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa512_y4;
  assign f_s_dadda_pg_rca32_fa526_y2 = f_s_dadda_pg_rca32_fa526_y0 ^ f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa511_y4;
  assign f_s_dadda_pg_rca32_fa526_y3 = f_s_dadda_pg_rca32_fa526_y0 & f_s_dadda_pg_rca32_fa526_f_s_dadda_pg_rca32_fa511_y4;
  assign f_s_dadda_pg_rca32_fa526_y4 = f_s_dadda_pg_rca32_fa526_y1 | f_s_dadda_pg_rca32_fa526_y3;
  assign f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa510_y4 = f_s_dadda_pg_rca32_fa510_y4;
  assign f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa509_y4 = f_s_dadda_pg_rca32_fa509_y4;
  assign f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa508_y4 = f_s_dadda_pg_rca32_fa508_y4;
  assign f_s_dadda_pg_rca32_fa527_y0 = f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa510_y4 ^ f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa509_y4;
  assign f_s_dadda_pg_rca32_fa527_y1 = f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa510_y4 & f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa509_y4;
  assign f_s_dadda_pg_rca32_fa527_y2 = f_s_dadda_pg_rca32_fa527_y0 ^ f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa508_y4;
  assign f_s_dadda_pg_rca32_fa527_y3 = f_s_dadda_pg_rca32_fa527_y0 & f_s_dadda_pg_rca32_fa527_f_s_dadda_pg_rca32_fa508_y4;
  assign f_s_dadda_pg_rca32_fa527_y4 = f_s_dadda_pg_rca32_fa527_y1 | f_s_dadda_pg_rca32_fa527_y3;
  assign f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa507_y4 = f_s_dadda_pg_rca32_fa507_y4;
  assign f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa506_y4 = f_s_dadda_pg_rca32_fa506_y4;
  assign f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa505_y4 = f_s_dadda_pg_rca32_fa505_y4;
  assign f_s_dadda_pg_rca32_fa528_y0 = f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa507_y4 ^ f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa506_y4;
  assign f_s_dadda_pg_rca32_fa528_y1 = f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa507_y4 & f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa506_y4;
  assign f_s_dadda_pg_rca32_fa528_y2 = f_s_dadda_pg_rca32_fa528_y0 ^ f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa505_y4;
  assign f_s_dadda_pg_rca32_fa528_y3 = f_s_dadda_pg_rca32_fa528_y0 & f_s_dadda_pg_rca32_fa528_f_s_dadda_pg_rca32_fa505_y4;
  assign f_s_dadda_pg_rca32_fa528_y4 = f_s_dadda_pg_rca32_fa528_y1 | f_s_dadda_pg_rca32_fa528_y3;
  assign f_s_dadda_pg_rca32_nand_31_10_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_nand_31_10_y0 = ~(f_s_dadda_pg_rca32_nand_31_10_a_31 & f_s_dadda_pg_rca32_nand_31_10_b_10);
  assign f_s_dadda_pg_rca32_and_30_11_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_and_30_11_y0 = f_s_dadda_pg_rca32_and_30_11_a_30 & f_s_dadda_pg_rca32_and_30_11_b_11;
  assign f_s_dadda_pg_rca32_and_29_12_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_29_12_y0 = f_s_dadda_pg_rca32_and_29_12_a_29 & f_s_dadda_pg_rca32_and_29_12_b_12;
  assign f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_nand_31_10_y0 = f_s_dadda_pg_rca32_nand_31_10_y0;
  assign f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_and_30_11_y0 = f_s_dadda_pg_rca32_and_30_11_y0;
  assign f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_and_29_12_y0 = f_s_dadda_pg_rca32_and_29_12_y0;
  assign f_s_dadda_pg_rca32_fa529_y0 = f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_nand_31_10_y0 ^ f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_and_30_11_y0;
  assign f_s_dadda_pg_rca32_fa529_y1 = f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_nand_31_10_y0 & f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_and_30_11_y0;
  assign f_s_dadda_pg_rca32_fa529_y2 = f_s_dadda_pg_rca32_fa529_y0 ^ f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_and_29_12_y0;
  assign f_s_dadda_pg_rca32_fa529_y3 = f_s_dadda_pg_rca32_fa529_y0 & f_s_dadda_pg_rca32_fa529_f_s_dadda_pg_rca32_and_29_12_y0;
  assign f_s_dadda_pg_rca32_fa529_y4 = f_s_dadda_pg_rca32_fa529_y1 | f_s_dadda_pg_rca32_fa529_y3;
  assign f_s_dadda_pg_rca32_and_28_13_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_28_13_y0 = f_s_dadda_pg_rca32_and_28_13_a_28 & f_s_dadda_pg_rca32_and_28_13_b_13;
  assign f_s_dadda_pg_rca32_and_27_14_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_27_14_y0 = f_s_dadda_pg_rca32_and_27_14_a_27 & f_s_dadda_pg_rca32_and_27_14_b_14;
  assign f_s_dadda_pg_rca32_and_26_15_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_26_15_y0 = f_s_dadda_pg_rca32_and_26_15_a_26 & f_s_dadda_pg_rca32_and_26_15_b_15;
  assign f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_28_13_y0 = f_s_dadda_pg_rca32_and_28_13_y0;
  assign f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_27_14_y0 = f_s_dadda_pg_rca32_and_27_14_y0;
  assign f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_26_15_y0 = f_s_dadda_pg_rca32_and_26_15_y0;
  assign f_s_dadda_pg_rca32_fa530_y0 = f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_28_13_y0 ^ f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_27_14_y0;
  assign f_s_dadda_pg_rca32_fa530_y1 = f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_28_13_y0 & f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_27_14_y0;
  assign f_s_dadda_pg_rca32_fa530_y2 = f_s_dadda_pg_rca32_fa530_y0 ^ f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_26_15_y0;
  assign f_s_dadda_pg_rca32_fa530_y3 = f_s_dadda_pg_rca32_fa530_y0 & f_s_dadda_pg_rca32_fa530_f_s_dadda_pg_rca32_and_26_15_y0;
  assign f_s_dadda_pg_rca32_fa530_y4 = f_s_dadda_pg_rca32_fa530_y1 | f_s_dadda_pg_rca32_fa530_y3;
  assign f_s_dadda_pg_rca32_and_25_16_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_25_16_y0 = f_s_dadda_pg_rca32_and_25_16_a_25 & f_s_dadda_pg_rca32_and_25_16_b_16;
  assign f_s_dadda_pg_rca32_and_24_17_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_24_17_y0 = f_s_dadda_pg_rca32_and_24_17_a_24 & f_s_dadda_pg_rca32_and_24_17_b_17;
  assign f_s_dadda_pg_rca32_and_23_18_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_23_18_y0 = f_s_dadda_pg_rca32_and_23_18_a_23 & f_s_dadda_pg_rca32_and_23_18_b_18;
  assign f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_25_16_y0 = f_s_dadda_pg_rca32_and_25_16_y0;
  assign f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_24_17_y0 = f_s_dadda_pg_rca32_and_24_17_y0;
  assign f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_23_18_y0 = f_s_dadda_pg_rca32_and_23_18_y0;
  assign f_s_dadda_pg_rca32_fa531_y0 = f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_25_16_y0 ^ f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_24_17_y0;
  assign f_s_dadda_pg_rca32_fa531_y1 = f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_25_16_y0 & f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_24_17_y0;
  assign f_s_dadda_pg_rca32_fa531_y2 = f_s_dadda_pg_rca32_fa531_y0 ^ f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_23_18_y0;
  assign f_s_dadda_pg_rca32_fa531_y3 = f_s_dadda_pg_rca32_fa531_y0 & f_s_dadda_pg_rca32_fa531_f_s_dadda_pg_rca32_and_23_18_y0;
  assign f_s_dadda_pg_rca32_fa531_y4 = f_s_dadda_pg_rca32_fa531_y1 | f_s_dadda_pg_rca32_fa531_y3;
  assign f_s_dadda_pg_rca32_and_22_19_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_22_19_y0 = f_s_dadda_pg_rca32_and_22_19_a_22 & f_s_dadda_pg_rca32_and_22_19_b_19;
  assign f_s_dadda_pg_rca32_and_21_20_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_21_20_y0 = f_s_dadda_pg_rca32_and_21_20_a_21 & f_s_dadda_pg_rca32_and_21_20_b_20;
  assign f_s_dadda_pg_rca32_and_20_21_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_20_21_y0 = f_s_dadda_pg_rca32_and_20_21_a_20 & f_s_dadda_pg_rca32_and_20_21_b_21;
  assign f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_22_19_y0 = f_s_dadda_pg_rca32_and_22_19_y0;
  assign f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_21_20_y0 = f_s_dadda_pg_rca32_and_21_20_y0;
  assign f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_20_21_y0 = f_s_dadda_pg_rca32_and_20_21_y0;
  assign f_s_dadda_pg_rca32_fa532_y0 = f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_22_19_y0 ^ f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_21_20_y0;
  assign f_s_dadda_pg_rca32_fa532_y1 = f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_22_19_y0 & f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_21_20_y0;
  assign f_s_dadda_pg_rca32_fa532_y2 = f_s_dadda_pg_rca32_fa532_y0 ^ f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_20_21_y0;
  assign f_s_dadda_pg_rca32_fa532_y3 = f_s_dadda_pg_rca32_fa532_y0 & f_s_dadda_pg_rca32_fa532_f_s_dadda_pg_rca32_and_20_21_y0;
  assign f_s_dadda_pg_rca32_fa532_y4 = f_s_dadda_pg_rca32_fa532_y1 | f_s_dadda_pg_rca32_fa532_y3;
  assign f_s_dadda_pg_rca32_and_19_22_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_19_22_y0 = f_s_dadda_pg_rca32_and_19_22_a_19 & f_s_dadda_pg_rca32_and_19_22_b_22;
  assign f_s_dadda_pg_rca32_and_18_23_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_18_23_y0 = f_s_dadda_pg_rca32_and_18_23_a_18 & f_s_dadda_pg_rca32_and_18_23_b_23;
  assign f_s_dadda_pg_rca32_and_17_24_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_17_24_y0 = f_s_dadda_pg_rca32_and_17_24_a_17 & f_s_dadda_pg_rca32_and_17_24_b_24;
  assign f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_19_22_y0 = f_s_dadda_pg_rca32_and_19_22_y0;
  assign f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_18_23_y0 = f_s_dadda_pg_rca32_and_18_23_y0;
  assign f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_17_24_y0 = f_s_dadda_pg_rca32_and_17_24_y0;
  assign f_s_dadda_pg_rca32_fa533_y0 = f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_19_22_y0 ^ f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_18_23_y0;
  assign f_s_dadda_pg_rca32_fa533_y1 = f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_19_22_y0 & f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_18_23_y0;
  assign f_s_dadda_pg_rca32_fa533_y2 = f_s_dadda_pg_rca32_fa533_y0 ^ f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_17_24_y0;
  assign f_s_dadda_pg_rca32_fa533_y3 = f_s_dadda_pg_rca32_fa533_y0 & f_s_dadda_pg_rca32_fa533_f_s_dadda_pg_rca32_and_17_24_y0;
  assign f_s_dadda_pg_rca32_fa533_y4 = f_s_dadda_pg_rca32_fa533_y1 | f_s_dadda_pg_rca32_fa533_y3;
  assign f_s_dadda_pg_rca32_and_16_25_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_16_25_y0 = f_s_dadda_pg_rca32_and_16_25_a_16 & f_s_dadda_pg_rca32_and_16_25_b_25;
  assign f_s_dadda_pg_rca32_and_15_26_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_15_26_y0 = f_s_dadda_pg_rca32_and_15_26_a_15 & f_s_dadda_pg_rca32_and_15_26_b_26;
  assign f_s_dadda_pg_rca32_and_14_27_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_14_27_y0 = f_s_dadda_pg_rca32_and_14_27_a_14 & f_s_dadda_pg_rca32_and_14_27_b_27;
  assign f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_16_25_y0 = f_s_dadda_pg_rca32_and_16_25_y0;
  assign f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_15_26_y0 = f_s_dadda_pg_rca32_and_15_26_y0;
  assign f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_14_27_y0 = f_s_dadda_pg_rca32_and_14_27_y0;
  assign f_s_dadda_pg_rca32_fa534_y0 = f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_16_25_y0 ^ f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_15_26_y0;
  assign f_s_dadda_pg_rca32_fa534_y1 = f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_16_25_y0 & f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_15_26_y0;
  assign f_s_dadda_pg_rca32_fa534_y2 = f_s_dadda_pg_rca32_fa534_y0 ^ f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_14_27_y0;
  assign f_s_dadda_pg_rca32_fa534_y3 = f_s_dadda_pg_rca32_fa534_y0 & f_s_dadda_pg_rca32_fa534_f_s_dadda_pg_rca32_and_14_27_y0;
  assign f_s_dadda_pg_rca32_fa534_y4 = f_s_dadda_pg_rca32_fa534_y1 | f_s_dadda_pg_rca32_fa534_y3;
  assign f_s_dadda_pg_rca32_and_13_28_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_13_28_y0 = f_s_dadda_pg_rca32_and_13_28_a_13 & f_s_dadda_pg_rca32_and_13_28_b_28;
  assign f_s_dadda_pg_rca32_and_12_29_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_12_29_y0 = f_s_dadda_pg_rca32_and_12_29_a_12 & f_s_dadda_pg_rca32_and_12_29_b_29;
  assign f_s_dadda_pg_rca32_and_11_30_a_11 = a_11;
  assign f_s_dadda_pg_rca32_and_11_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_11_30_y0 = f_s_dadda_pg_rca32_and_11_30_a_11 & f_s_dadda_pg_rca32_and_11_30_b_30;
  assign f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_13_28_y0 = f_s_dadda_pg_rca32_and_13_28_y0;
  assign f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_12_29_y0 = f_s_dadda_pg_rca32_and_12_29_y0;
  assign f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_11_30_y0 = f_s_dadda_pg_rca32_and_11_30_y0;
  assign f_s_dadda_pg_rca32_fa535_y0 = f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_13_28_y0 ^ f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_12_29_y0;
  assign f_s_dadda_pg_rca32_fa535_y1 = f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_13_28_y0 & f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_12_29_y0;
  assign f_s_dadda_pg_rca32_fa535_y2 = f_s_dadda_pg_rca32_fa535_y0 ^ f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_11_30_y0;
  assign f_s_dadda_pg_rca32_fa535_y3 = f_s_dadda_pg_rca32_fa535_y0 & f_s_dadda_pg_rca32_fa535_f_s_dadda_pg_rca32_and_11_30_y0;
  assign f_s_dadda_pg_rca32_fa535_y4 = f_s_dadda_pg_rca32_fa535_y1 | f_s_dadda_pg_rca32_fa535_y3;
  assign f_s_dadda_pg_rca32_nand_10_31_a_10 = a_10;
  assign f_s_dadda_pg_rca32_nand_10_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_10_31_y0 = ~(f_s_dadda_pg_rca32_nand_10_31_a_10 & f_s_dadda_pg_rca32_nand_10_31_b_31);
  assign f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_nand_10_31_y0 = f_s_dadda_pg_rca32_nand_10_31_y0;
  assign f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_fa523_y2 = f_s_dadda_pg_rca32_fa523_y2;
  assign f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_fa524_y2 = f_s_dadda_pg_rca32_fa524_y2;
  assign f_s_dadda_pg_rca32_fa536_y0 = f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_nand_10_31_y0 ^ f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_fa523_y2;
  assign f_s_dadda_pg_rca32_fa536_y1 = f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_nand_10_31_y0 & f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_fa523_y2;
  assign f_s_dadda_pg_rca32_fa536_y2 = f_s_dadda_pg_rca32_fa536_y0 ^ f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_fa524_y2;
  assign f_s_dadda_pg_rca32_fa536_y3 = f_s_dadda_pg_rca32_fa536_y0 & f_s_dadda_pg_rca32_fa536_f_s_dadda_pg_rca32_fa524_y2;
  assign f_s_dadda_pg_rca32_fa536_y4 = f_s_dadda_pg_rca32_fa536_y1 | f_s_dadda_pg_rca32_fa536_y3;
  assign f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa525_y2 = f_s_dadda_pg_rca32_fa525_y2;
  assign f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa526_y2 = f_s_dadda_pg_rca32_fa526_y2;
  assign f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa527_y2 = f_s_dadda_pg_rca32_fa527_y2;
  assign f_s_dadda_pg_rca32_fa537_y0 = f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa525_y2 ^ f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa526_y2;
  assign f_s_dadda_pg_rca32_fa537_y1 = f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa525_y2 & f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa526_y2;
  assign f_s_dadda_pg_rca32_fa537_y2 = f_s_dadda_pg_rca32_fa537_y0 ^ f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa527_y2;
  assign f_s_dadda_pg_rca32_fa537_y3 = f_s_dadda_pg_rca32_fa537_y0 & f_s_dadda_pg_rca32_fa537_f_s_dadda_pg_rca32_fa527_y2;
  assign f_s_dadda_pg_rca32_fa537_y4 = f_s_dadda_pg_rca32_fa537_y1 | f_s_dadda_pg_rca32_fa537_y3;
  assign f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa528_y2 = f_s_dadda_pg_rca32_fa528_y2;
  assign f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa529_y2 = f_s_dadda_pg_rca32_fa529_y2;
  assign f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa530_y2 = f_s_dadda_pg_rca32_fa530_y2;
  assign f_s_dadda_pg_rca32_fa538_y0 = f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa528_y2 ^ f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa529_y2;
  assign f_s_dadda_pg_rca32_fa538_y1 = f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa528_y2 & f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa529_y2;
  assign f_s_dadda_pg_rca32_fa538_y2 = f_s_dadda_pg_rca32_fa538_y0 ^ f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa530_y2;
  assign f_s_dadda_pg_rca32_fa538_y3 = f_s_dadda_pg_rca32_fa538_y0 & f_s_dadda_pg_rca32_fa538_f_s_dadda_pg_rca32_fa530_y2;
  assign f_s_dadda_pg_rca32_fa538_y4 = f_s_dadda_pg_rca32_fa538_y1 | f_s_dadda_pg_rca32_fa538_y3;
  assign f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa531_y2 = f_s_dadda_pg_rca32_fa531_y2;
  assign f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa532_y2 = f_s_dadda_pg_rca32_fa532_y2;
  assign f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa533_y2 = f_s_dadda_pg_rca32_fa533_y2;
  assign f_s_dadda_pg_rca32_fa539_y0 = f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa531_y2 ^ f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa532_y2;
  assign f_s_dadda_pg_rca32_fa539_y1 = f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa531_y2 & f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa532_y2;
  assign f_s_dadda_pg_rca32_fa539_y2 = f_s_dadda_pg_rca32_fa539_y0 ^ f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa533_y2;
  assign f_s_dadda_pg_rca32_fa539_y3 = f_s_dadda_pg_rca32_fa539_y0 & f_s_dadda_pg_rca32_fa539_f_s_dadda_pg_rca32_fa533_y2;
  assign f_s_dadda_pg_rca32_fa539_y4 = f_s_dadda_pg_rca32_fa539_y1 | f_s_dadda_pg_rca32_fa539_y3;
  assign f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa539_y4 = f_s_dadda_pg_rca32_fa539_y4;
  assign f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa538_y4 = f_s_dadda_pg_rca32_fa538_y4;
  assign f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa537_y4 = f_s_dadda_pg_rca32_fa537_y4;
  assign f_s_dadda_pg_rca32_fa540_y0 = f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa539_y4 ^ f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa538_y4;
  assign f_s_dadda_pg_rca32_fa540_y1 = f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa539_y4 & f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa538_y4;
  assign f_s_dadda_pg_rca32_fa540_y2 = f_s_dadda_pg_rca32_fa540_y0 ^ f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa537_y4;
  assign f_s_dadda_pg_rca32_fa540_y3 = f_s_dadda_pg_rca32_fa540_y0 & f_s_dadda_pg_rca32_fa540_f_s_dadda_pg_rca32_fa537_y4;
  assign f_s_dadda_pg_rca32_fa540_y4 = f_s_dadda_pg_rca32_fa540_y1 | f_s_dadda_pg_rca32_fa540_y3;
  assign f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa536_y4 = f_s_dadda_pg_rca32_fa536_y4;
  assign f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa535_y4 = f_s_dadda_pg_rca32_fa535_y4;
  assign f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa534_y4 = f_s_dadda_pg_rca32_fa534_y4;
  assign f_s_dadda_pg_rca32_fa541_y0 = f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa536_y4 ^ f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa535_y4;
  assign f_s_dadda_pg_rca32_fa541_y1 = f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa536_y4 & f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa535_y4;
  assign f_s_dadda_pg_rca32_fa541_y2 = f_s_dadda_pg_rca32_fa541_y0 ^ f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa534_y4;
  assign f_s_dadda_pg_rca32_fa541_y3 = f_s_dadda_pg_rca32_fa541_y0 & f_s_dadda_pg_rca32_fa541_f_s_dadda_pg_rca32_fa534_y4;
  assign f_s_dadda_pg_rca32_fa541_y4 = f_s_dadda_pg_rca32_fa541_y1 | f_s_dadda_pg_rca32_fa541_y3;
  assign f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa533_y4 = f_s_dadda_pg_rca32_fa533_y4;
  assign f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa532_y4 = f_s_dadda_pg_rca32_fa532_y4;
  assign f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa531_y4 = f_s_dadda_pg_rca32_fa531_y4;
  assign f_s_dadda_pg_rca32_fa542_y0 = f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa533_y4 ^ f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa532_y4;
  assign f_s_dadda_pg_rca32_fa542_y1 = f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa533_y4 & f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa532_y4;
  assign f_s_dadda_pg_rca32_fa542_y2 = f_s_dadda_pg_rca32_fa542_y0 ^ f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa531_y4;
  assign f_s_dadda_pg_rca32_fa542_y3 = f_s_dadda_pg_rca32_fa542_y0 & f_s_dadda_pg_rca32_fa542_f_s_dadda_pg_rca32_fa531_y4;
  assign f_s_dadda_pg_rca32_fa542_y4 = f_s_dadda_pg_rca32_fa542_y1 | f_s_dadda_pg_rca32_fa542_y3;
  assign f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa530_y4 = f_s_dadda_pg_rca32_fa530_y4;
  assign f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa529_y4 = f_s_dadda_pg_rca32_fa529_y4;
  assign f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa528_y4 = f_s_dadda_pg_rca32_fa528_y4;
  assign f_s_dadda_pg_rca32_fa543_y0 = f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa530_y4 ^ f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa529_y4;
  assign f_s_dadda_pg_rca32_fa543_y1 = f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa530_y4 & f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa529_y4;
  assign f_s_dadda_pg_rca32_fa543_y2 = f_s_dadda_pg_rca32_fa543_y0 ^ f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa528_y4;
  assign f_s_dadda_pg_rca32_fa543_y3 = f_s_dadda_pg_rca32_fa543_y0 & f_s_dadda_pg_rca32_fa543_f_s_dadda_pg_rca32_fa528_y4;
  assign f_s_dadda_pg_rca32_fa543_y4 = f_s_dadda_pg_rca32_fa543_y1 | f_s_dadda_pg_rca32_fa543_y3;
  assign f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa527_y4 = f_s_dadda_pg_rca32_fa527_y4;
  assign f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa526_y4 = f_s_dadda_pg_rca32_fa526_y4;
  assign f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa525_y4 = f_s_dadda_pg_rca32_fa525_y4;
  assign f_s_dadda_pg_rca32_fa544_y0 = f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa527_y4 ^ f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa526_y4;
  assign f_s_dadda_pg_rca32_fa544_y1 = f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa527_y4 & f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa526_y4;
  assign f_s_dadda_pg_rca32_fa544_y2 = f_s_dadda_pg_rca32_fa544_y0 ^ f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa525_y4;
  assign f_s_dadda_pg_rca32_fa544_y3 = f_s_dadda_pg_rca32_fa544_y0 & f_s_dadda_pg_rca32_fa544_f_s_dadda_pg_rca32_fa525_y4;
  assign f_s_dadda_pg_rca32_fa544_y4 = f_s_dadda_pg_rca32_fa544_y1 | f_s_dadda_pg_rca32_fa544_y3;
  assign f_s_dadda_pg_rca32_nand_31_11_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_11_b_11 = b_11;
  assign f_s_dadda_pg_rca32_nand_31_11_y0 = ~(f_s_dadda_pg_rca32_nand_31_11_a_31 & f_s_dadda_pg_rca32_nand_31_11_b_11);
  assign f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_fa524_y4 = f_s_dadda_pg_rca32_fa524_y4;
  assign f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_fa523_y4 = f_s_dadda_pg_rca32_fa523_y4;
  assign f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_nand_31_11_y0 = f_s_dadda_pg_rca32_nand_31_11_y0;
  assign f_s_dadda_pg_rca32_fa545_y0 = f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_fa524_y4 ^ f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_fa523_y4;
  assign f_s_dadda_pg_rca32_fa545_y1 = f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_fa524_y4 & f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_fa523_y4;
  assign f_s_dadda_pg_rca32_fa545_y2 = f_s_dadda_pg_rca32_fa545_y0 ^ f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_nand_31_11_y0;
  assign f_s_dadda_pg_rca32_fa545_y3 = f_s_dadda_pg_rca32_fa545_y0 & f_s_dadda_pg_rca32_fa545_f_s_dadda_pg_rca32_nand_31_11_y0;
  assign f_s_dadda_pg_rca32_fa545_y4 = f_s_dadda_pg_rca32_fa545_y1 | f_s_dadda_pg_rca32_fa545_y3;
  assign f_s_dadda_pg_rca32_and_30_12_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_and_30_12_y0 = f_s_dadda_pg_rca32_and_30_12_a_30 & f_s_dadda_pg_rca32_and_30_12_b_12;
  assign f_s_dadda_pg_rca32_and_29_13_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_29_13_y0 = f_s_dadda_pg_rca32_and_29_13_a_29 & f_s_dadda_pg_rca32_and_29_13_b_13;
  assign f_s_dadda_pg_rca32_and_28_14_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_28_14_y0 = f_s_dadda_pg_rca32_and_28_14_a_28 & f_s_dadda_pg_rca32_and_28_14_b_14;
  assign f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_30_12_y0 = f_s_dadda_pg_rca32_and_30_12_y0;
  assign f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_29_13_y0 = f_s_dadda_pg_rca32_and_29_13_y0;
  assign f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_28_14_y0 = f_s_dadda_pg_rca32_and_28_14_y0;
  assign f_s_dadda_pg_rca32_fa546_y0 = f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_30_12_y0 ^ f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_29_13_y0;
  assign f_s_dadda_pg_rca32_fa546_y1 = f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_30_12_y0 & f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_29_13_y0;
  assign f_s_dadda_pg_rca32_fa546_y2 = f_s_dadda_pg_rca32_fa546_y0 ^ f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_28_14_y0;
  assign f_s_dadda_pg_rca32_fa546_y3 = f_s_dadda_pg_rca32_fa546_y0 & f_s_dadda_pg_rca32_fa546_f_s_dadda_pg_rca32_and_28_14_y0;
  assign f_s_dadda_pg_rca32_fa546_y4 = f_s_dadda_pg_rca32_fa546_y1 | f_s_dadda_pg_rca32_fa546_y3;
  assign f_s_dadda_pg_rca32_and_27_15_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_27_15_y0 = f_s_dadda_pg_rca32_and_27_15_a_27 & f_s_dadda_pg_rca32_and_27_15_b_15;
  assign f_s_dadda_pg_rca32_and_26_16_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_26_16_y0 = f_s_dadda_pg_rca32_and_26_16_a_26 & f_s_dadda_pg_rca32_and_26_16_b_16;
  assign f_s_dadda_pg_rca32_and_25_17_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_25_17_y0 = f_s_dadda_pg_rca32_and_25_17_a_25 & f_s_dadda_pg_rca32_and_25_17_b_17;
  assign f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_27_15_y0 = f_s_dadda_pg_rca32_and_27_15_y0;
  assign f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_26_16_y0 = f_s_dadda_pg_rca32_and_26_16_y0;
  assign f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_25_17_y0 = f_s_dadda_pg_rca32_and_25_17_y0;
  assign f_s_dadda_pg_rca32_fa547_y0 = f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_27_15_y0 ^ f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_26_16_y0;
  assign f_s_dadda_pg_rca32_fa547_y1 = f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_27_15_y0 & f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_26_16_y0;
  assign f_s_dadda_pg_rca32_fa547_y2 = f_s_dadda_pg_rca32_fa547_y0 ^ f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_25_17_y0;
  assign f_s_dadda_pg_rca32_fa547_y3 = f_s_dadda_pg_rca32_fa547_y0 & f_s_dadda_pg_rca32_fa547_f_s_dadda_pg_rca32_and_25_17_y0;
  assign f_s_dadda_pg_rca32_fa547_y4 = f_s_dadda_pg_rca32_fa547_y1 | f_s_dadda_pg_rca32_fa547_y3;
  assign f_s_dadda_pg_rca32_and_24_18_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_24_18_y0 = f_s_dadda_pg_rca32_and_24_18_a_24 & f_s_dadda_pg_rca32_and_24_18_b_18;
  assign f_s_dadda_pg_rca32_and_23_19_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_23_19_y0 = f_s_dadda_pg_rca32_and_23_19_a_23 & f_s_dadda_pg_rca32_and_23_19_b_19;
  assign f_s_dadda_pg_rca32_and_22_20_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_22_20_y0 = f_s_dadda_pg_rca32_and_22_20_a_22 & f_s_dadda_pg_rca32_and_22_20_b_20;
  assign f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_24_18_y0 = f_s_dadda_pg_rca32_and_24_18_y0;
  assign f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_23_19_y0 = f_s_dadda_pg_rca32_and_23_19_y0;
  assign f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_22_20_y0 = f_s_dadda_pg_rca32_and_22_20_y0;
  assign f_s_dadda_pg_rca32_fa548_y0 = f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_24_18_y0 ^ f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_23_19_y0;
  assign f_s_dadda_pg_rca32_fa548_y1 = f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_24_18_y0 & f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_23_19_y0;
  assign f_s_dadda_pg_rca32_fa548_y2 = f_s_dadda_pg_rca32_fa548_y0 ^ f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_22_20_y0;
  assign f_s_dadda_pg_rca32_fa548_y3 = f_s_dadda_pg_rca32_fa548_y0 & f_s_dadda_pg_rca32_fa548_f_s_dadda_pg_rca32_and_22_20_y0;
  assign f_s_dadda_pg_rca32_fa548_y4 = f_s_dadda_pg_rca32_fa548_y1 | f_s_dadda_pg_rca32_fa548_y3;
  assign f_s_dadda_pg_rca32_and_21_21_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_21_21_y0 = f_s_dadda_pg_rca32_and_21_21_a_21 & f_s_dadda_pg_rca32_and_21_21_b_21;
  assign f_s_dadda_pg_rca32_and_20_22_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_20_22_y0 = f_s_dadda_pg_rca32_and_20_22_a_20 & f_s_dadda_pg_rca32_and_20_22_b_22;
  assign f_s_dadda_pg_rca32_and_19_23_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_19_23_y0 = f_s_dadda_pg_rca32_and_19_23_a_19 & f_s_dadda_pg_rca32_and_19_23_b_23;
  assign f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_21_21_y0 = f_s_dadda_pg_rca32_and_21_21_y0;
  assign f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_20_22_y0 = f_s_dadda_pg_rca32_and_20_22_y0;
  assign f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_19_23_y0 = f_s_dadda_pg_rca32_and_19_23_y0;
  assign f_s_dadda_pg_rca32_fa549_y0 = f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_21_21_y0 ^ f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_20_22_y0;
  assign f_s_dadda_pg_rca32_fa549_y1 = f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_21_21_y0 & f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_20_22_y0;
  assign f_s_dadda_pg_rca32_fa549_y2 = f_s_dadda_pg_rca32_fa549_y0 ^ f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_19_23_y0;
  assign f_s_dadda_pg_rca32_fa549_y3 = f_s_dadda_pg_rca32_fa549_y0 & f_s_dadda_pg_rca32_fa549_f_s_dadda_pg_rca32_and_19_23_y0;
  assign f_s_dadda_pg_rca32_fa549_y4 = f_s_dadda_pg_rca32_fa549_y1 | f_s_dadda_pg_rca32_fa549_y3;
  assign f_s_dadda_pg_rca32_and_18_24_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_18_24_y0 = f_s_dadda_pg_rca32_and_18_24_a_18 & f_s_dadda_pg_rca32_and_18_24_b_24;
  assign f_s_dadda_pg_rca32_and_17_25_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_17_25_y0 = f_s_dadda_pg_rca32_and_17_25_a_17 & f_s_dadda_pg_rca32_and_17_25_b_25;
  assign f_s_dadda_pg_rca32_and_16_26_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_16_26_y0 = f_s_dadda_pg_rca32_and_16_26_a_16 & f_s_dadda_pg_rca32_and_16_26_b_26;
  assign f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_18_24_y0 = f_s_dadda_pg_rca32_and_18_24_y0;
  assign f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_17_25_y0 = f_s_dadda_pg_rca32_and_17_25_y0;
  assign f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_16_26_y0 = f_s_dadda_pg_rca32_and_16_26_y0;
  assign f_s_dadda_pg_rca32_fa550_y0 = f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_18_24_y0 ^ f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_17_25_y0;
  assign f_s_dadda_pg_rca32_fa550_y1 = f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_18_24_y0 & f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_17_25_y0;
  assign f_s_dadda_pg_rca32_fa550_y2 = f_s_dadda_pg_rca32_fa550_y0 ^ f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_16_26_y0;
  assign f_s_dadda_pg_rca32_fa550_y3 = f_s_dadda_pg_rca32_fa550_y0 & f_s_dadda_pg_rca32_fa550_f_s_dadda_pg_rca32_and_16_26_y0;
  assign f_s_dadda_pg_rca32_fa550_y4 = f_s_dadda_pg_rca32_fa550_y1 | f_s_dadda_pg_rca32_fa550_y3;
  assign f_s_dadda_pg_rca32_and_15_27_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_15_27_y0 = f_s_dadda_pg_rca32_and_15_27_a_15 & f_s_dadda_pg_rca32_and_15_27_b_27;
  assign f_s_dadda_pg_rca32_and_14_28_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_14_28_y0 = f_s_dadda_pg_rca32_and_14_28_a_14 & f_s_dadda_pg_rca32_and_14_28_b_28;
  assign f_s_dadda_pg_rca32_and_13_29_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_13_29_y0 = f_s_dadda_pg_rca32_and_13_29_a_13 & f_s_dadda_pg_rca32_and_13_29_b_29;
  assign f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_15_27_y0 = f_s_dadda_pg_rca32_and_15_27_y0;
  assign f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_14_28_y0 = f_s_dadda_pg_rca32_and_14_28_y0;
  assign f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_13_29_y0 = f_s_dadda_pg_rca32_and_13_29_y0;
  assign f_s_dadda_pg_rca32_fa551_y0 = f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_15_27_y0 ^ f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_14_28_y0;
  assign f_s_dadda_pg_rca32_fa551_y1 = f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_15_27_y0 & f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_14_28_y0;
  assign f_s_dadda_pg_rca32_fa551_y2 = f_s_dadda_pg_rca32_fa551_y0 ^ f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_13_29_y0;
  assign f_s_dadda_pg_rca32_fa551_y3 = f_s_dadda_pg_rca32_fa551_y0 & f_s_dadda_pg_rca32_fa551_f_s_dadda_pg_rca32_and_13_29_y0;
  assign f_s_dadda_pg_rca32_fa551_y4 = f_s_dadda_pg_rca32_fa551_y1 | f_s_dadda_pg_rca32_fa551_y3;
  assign f_s_dadda_pg_rca32_and_12_30_a_12 = a_12;
  assign f_s_dadda_pg_rca32_and_12_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_12_30_y0 = f_s_dadda_pg_rca32_and_12_30_a_12 & f_s_dadda_pg_rca32_and_12_30_b_30;
  assign f_s_dadda_pg_rca32_nand_11_31_a_11 = a_11;
  assign f_s_dadda_pg_rca32_nand_11_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_11_31_y0 = ~(f_s_dadda_pg_rca32_nand_11_31_a_11 & f_s_dadda_pg_rca32_nand_11_31_b_31);
  assign f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_and_12_30_y0 = f_s_dadda_pg_rca32_and_12_30_y0;
  assign f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_nand_11_31_y0 = f_s_dadda_pg_rca32_nand_11_31_y0;
  assign f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_fa540_y2 = f_s_dadda_pg_rca32_fa540_y2;
  assign f_s_dadda_pg_rca32_fa552_y0 = f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_and_12_30_y0 ^ f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_nand_11_31_y0;
  assign f_s_dadda_pg_rca32_fa552_y1 = f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_and_12_30_y0 & f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_nand_11_31_y0;
  assign f_s_dadda_pg_rca32_fa552_y2 = f_s_dadda_pg_rca32_fa552_y0 ^ f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_fa540_y2;
  assign f_s_dadda_pg_rca32_fa552_y3 = f_s_dadda_pg_rca32_fa552_y0 & f_s_dadda_pg_rca32_fa552_f_s_dadda_pg_rca32_fa540_y2;
  assign f_s_dadda_pg_rca32_fa552_y4 = f_s_dadda_pg_rca32_fa552_y1 | f_s_dadda_pg_rca32_fa552_y3;
  assign f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa541_y2 = f_s_dadda_pg_rca32_fa541_y2;
  assign f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa542_y2 = f_s_dadda_pg_rca32_fa542_y2;
  assign f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa543_y2 = f_s_dadda_pg_rca32_fa543_y2;
  assign f_s_dadda_pg_rca32_fa553_y0 = f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa541_y2 ^ f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa542_y2;
  assign f_s_dadda_pg_rca32_fa553_y1 = f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa541_y2 & f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa542_y2;
  assign f_s_dadda_pg_rca32_fa553_y2 = f_s_dadda_pg_rca32_fa553_y0 ^ f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa543_y2;
  assign f_s_dadda_pg_rca32_fa553_y3 = f_s_dadda_pg_rca32_fa553_y0 & f_s_dadda_pg_rca32_fa553_f_s_dadda_pg_rca32_fa543_y2;
  assign f_s_dadda_pg_rca32_fa553_y4 = f_s_dadda_pg_rca32_fa553_y1 | f_s_dadda_pg_rca32_fa553_y3;
  assign f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa544_y2 = f_s_dadda_pg_rca32_fa544_y2;
  assign f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa545_y2 = f_s_dadda_pg_rca32_fa545_y2;
  assign f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa546_y2 = f_s_dadda_pg_rca32_fa546_y2;
  assign f_s_dadda_pg_rca32_fa554_y0 = f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa544_y2 ^ f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa545_y2;
  assign f_s_dadda_pg_rca32_fa554_y1 = f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa544_y2 & f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa545_y2;
  assign f_s_dadda_pg_rca32_fa554_y2 = f_s_dadda_pg_rca32_fa554_y0 ^ f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa546_y2;
  assign f_s_dadda_pg_rca32_fa554_y3 = f_s_dadda_pg_rca32_fa554_y0 & f_s_dadda_pg_rca32_fa554_f_s_dadda_pg_rca32_fa546_y2;
  assign f_s_dadda_pg_rca32_fa554_y4 = f_s_dadda_pg_rca32_fa554_y1 | f_s_dadda_pg_rca32_fa554_y3;
  assign f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa547_y2 = f_s_dadda_pg_rca32_fa547_y2;
  assign f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa548_y2 = f_s_dadda_pg_rca32_fa548_y2;
  assign f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa549_y2 = f_s_dadda_pg_rca32_fa549_y2;
  assign f_s_dadda_pg_rca32_fa555_y0 = f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa547_y2 ^ f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa548_y2;
  assign f_s_dadda_pg_rca32_fa555_y1 = f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa547_y2 & f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa548_y2;
  assign f_s_dadda_pg_rca32_fa555_y2 = f_s_dadda_pg_rca32_fa555_y0 ^ f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa549_y2;
  assign f_s_dadda_pg_rca32_fa555_y3 = f_s_dadda_pg_rca32_fa555_y0 & f_s_dadda_pg_rca32_fa555_f_s_dadda_pg_rca32_fa549_y2;
  assign f_s_dadda_pg_rca32_fa555_y4 = f_s_dadda_pg_rca32_fa555_y1 | f_s_dadda_pg_rca32_fa555_y3;
  assign f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa555_y4 = f_s_dadda_pg_rca32_fa555_y4;
  assign f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa554_y4 = f_s_dadda_pg_rca32_fa554_y4;
  assign f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa553_y4 = f_s_dadda_pg_rca32_fa553_y4;
  assign f_s_dadda_pg_rca32_fa556_y0 = f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa555_y4 ^ f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa554_y4;
  assign f_s_dadda_pg_rca32_fa556_y1 = f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa555_y4 & f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa554_y4;
  assign f_s_dadda_pg_rca32_fa556_y2 = f_s_dadda_pg_rca32_fa556_y0 ^ f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa553_y4;
  assign f_s_dadda_pg_rca32_fa556_y3 = f_s_dadda_pg_rca32_fa556_y0 & f_s_dadda_pg_rca32_fa556_f_s_dadda_pg_rca32_fa553_y4;
  assign f_s_dadda_pg_rca32_fa556_y4 = f_s_dadda_pg_rca32_fa556_y1 | f_s_dadda_pg_rca32_fa556_y3;
  assign f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa552_y4 = f_s_dadda_pg_rca32_fa552_y4;
  assign f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa551_y4 = f_s_dadda_pg_rca32_fa551_y4;
  assign f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa550_y4 = f_s_dadda_pg_rca32_fa550_y4;
  assign f_s_dadda_pg_rca32_fa557_y0 = f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa552_y4 ^ f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa551_y4;
  assign f_s_dadda_pg_rca32_fa557_y1 = f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa552_y4 & f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa551_y4;
  assign f_s_dadda_pg_rca32_fa557_y2 = f_s_dadda_pg_rca32_fa557_y0 ^ f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa550_y4;
  assign f_s_dadda_pg_rca32_fa557_y3 = f_s_dadda_pg_rca32_fa557_y0 & f_s_dadda_pg_rca32_fa557_f_s_dadda_pg_rca32_fa550_y4;
  assign f_s_dadda_pg_rca32_fa557_y4 = f_s_dadda_pg_rca32_fa557_y1 | f_s_dadda_pg_rca32_fa557_y3;
  assign f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa549_y4 = f_s_dadda_pg_rca32_fa549_y4;
  assign f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa548_y4 = f_s_dadda_pg_rca32_fa548_y4;
  assign f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa547_y4 = f_s_dadda_pg_rca32_fa547_y4;
  assign f_s_dadda_pg_rca32_fa558_y0 = f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa549_y4 ^ f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa548_y4;
  assign f_s_dadda_pg_rca32_fa558_y1 = f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa549_y4 & f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa548_y4;
  assign f_s_dadda_pg_rca32_fa558_y2 = f_s_dadda_pg_rca32_fa558_y0 ^ f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa547_y4;
  assign f_s_dadda_pg_rca32_fa558_y3 = f_s_dadda_pg_rca32_fa558_y0 & f_s_dadda_pg_rca32_fa558_f_s_dadda_pg_rca32_fa547_y4;
  assign f_s_dadda_pg_rca32_fa558_y4 = f_s_dadda_pg_rca32_fa558_y1 | f_s_dadda_pg_rca32_fa558_y3;
  assign f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa546_y4 = f_s_dadda_pg_rca32_fa546_y4;
  assign f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa545_y4 = f_s_dadda_pg_rca32_fa545_y4;
  assign f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa544_y4 = f_s_dadda_pg_rca32_fa544_y4;
  assign f_s_dadda_pg_rca32_fa559_y0 = f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa546_y4 ^ f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa545_y4;
  assign f_s_dadda_pg_rca32_fa559_y1 = f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa546_y4 & f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa545_y4;
  assign f_s_dadda_pg_rca32_fa559_y2 = f_s_dadda_pg_rca32_fa559_y0 ^ f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa544_y4;
  assign f_s_dadda_pg_rca32_fa559_y3 = f_s_dadda_pg_rca32_fa559_y0 & f_s_dadda_pg_rca32_fa559_f_s_dadda_pg_rca32_fa544_y4;
  assign f_s_dadda_pg_rca32_fa559_y4 = f_s_dadda_pg_rca32_fa559_y1 | f_s_dadda_pg_rca32_fa559_y3;
  assign f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa543_y4 = f_s_dadda_pg_rca32_fa543_y4;
  assign f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa542_y4 = f_s_dadda_pg_rca32_fa542_y4;
  assign f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa541_y4 = f_s_dadda_pg_rca32_fa541_y4;
  assign f_s_dadda_pg_rca32_fa560_y0 = f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa543_y4 ^ f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa542_y4;
  assign f_s_dadda_pg_rca32_fa560_y1 = f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa543_y4 & f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa542_y4;
  assign f_s_dadda_pg_rca32_fa560_y2 = f_s_dadda_pg_rca32_fa560_y0 ^ f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa541_y4;
  assign f_s_dadda_pg_rca32_fa560_y3 = f_s_dadda_pg_rca32_fa560_y0 & f_s_dadda_pg_rca32_fa560_f_s_dadda_pg_rca32_fa541_y4;
  assign f_s_dadda_pg_rca32_fa560_y4 = f_s_dadda_pg_rca32_fa560_y1 | f_s_dadda_pg_rca32_fa560_y3;
  assign f_s_dadda_pg_rca32_nand_31_12_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_12_b_12 = b_12;
  assign f_s_dadda_pg_rca32_nand_31_12_y0 = ~(f_s_dadda_pg_rca32_nand_31_12_a_31 & f_s_dadda_pg_rca32_nand_31_12_b_12);
  assign f_s_dadda_pg_rca32_and_30_13_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_and_30_13_y0 = f_s_dadda_pg_rca32_and_30_13_a_30 & f_s_dadda_pg_rca32_and_30_13_b_13;
  assign f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_fa540_y4 = f_s_dadda_pg_rca32_fa540_y4;
  assign f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_nand_31_12_y0 = f_s_dadda_pg_rca32_nand_31_12_y0;
  assign f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_and_30_13_y0 = f_s_dadda_pg_rca32_and_30_13_y0;
  assign f_s_dadda_pg_rca32_fa561_y0 = f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_fa540_y4 ^ f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_nand_31_12_y0;
  assign f_s_dadda_pg_rca32_fa561_y1 = f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_fa540_y4 & f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_nand_31_12_y0;
  assign f_s_dadda_pg_rca32_fa561_y2 = f_s_dadda_pg_rca32_fa561_y0 ^ f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_and_30_13_y0;
  assign f_s_dadda_pg_rca32_fa561_y3 = f_s_dadda_pg_rca32_fa561_y0 & f_s_dadda_pg_rca32_fa561_f_s_dadda_pg_rca32_and_30_13_y0;
  assign f_s_dadda_pg_rca32_fa561_y4 = f_s_dadda_pg_rca32_fa561_y1 | f_s_dadda_pg_rca32_fa561_y3;
  assign f_s_dadda_pg_rca32_and_29_14_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_29_14_y0 = f_s_dadda_pg_rca32_and_29_14_a_29 & f_s_dadda_pg_rca32_and_29_14_b_14;
  assign f_s_dadda_pg_rca32_and_28_15_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_28_15_y0 = f_s_dadda_pg_rca32_and_28_15_a_28 & f_s_dadda_pg_rca32_and_28_15_b_15;
  assign f_s_dadda_pg_rca32_and_27_16_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_27_16_y0 = f_s_dadda_pg_rca32_and_27_16_a_27 & f_s_dadda_pg_rca32_and_27_16_b_16;
  assign f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_29_14_y0 = f_s_dadda_pg_rca32_and_29_14_y0;
  assign f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_28_15_y0 = f_s_dadda_pg_rca32_and_28_15_y0;
  assign f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_27_16_y0 = f_s_dadda_pg_rca32_and_27_16_y0;
  assign f_s_dadda_pg_rca32_fa562_y0 = f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_29_14_y0 ^ f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_28_15_y0;
  assign f_s_dadda_pg_rca32_fa562_y1 = f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_29_14_y0 & f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_28_15_y0;
  assign f_s_dadda_pg_rca32_fa562_y2 = f_s_dadda_pg_rca32_fa562_y0 ^ f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_27_16_y0;
  assign f_s_dadda_pg_rca32_fa562_y3 = f_s_dadda_pg_rca32_fa562_y0 & f_s_dadda_pg_rca32_fa562_f_s_dadda_pg_rca32_and_27_16_y0;
  assign f_s_dadda_pg_rca32_fa562_y4 = f_s_dadda_pg_rca32_fa562_y1 | f_s_dadda_pg_rca32_fa562_y3;
  assign f_s_dadda_pg_rca32_and_26_17_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_26_17_y0 = f_s_dadda_pg_rca32_and_26_17_a_26 & f_s_dadda_pg_rca32_and_26_17_b_17;
  assign f_s_dadda_pg_rca32_and_25_18_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_25_18_y0 = f_s_dadda_pg_rca32_and_25_18_a_25 & f_s_dadda_pg_rca32_and_25_18_b_18;
  assign f_s_dadda_pg_rca32_and_24_19_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_24_19_y0 = f_s_dadda_pg_rca32_and_24_19_a_24 & f_s_dadda_pg_rca32_and_24_19_b_19;
  assign f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_26_17_y0 = f_s_dadda_pg_rca32_and_26_17_y0;
  assign f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_25_18_y0 = f_s_dadda_pg_rca32_and_25_18_y0;
  assign f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_24_19_y0 = f_s_dadda_pg_rca32_and_24_19_y0;
  assign f_s_dadda_pg_rca32_fa563_y0 = f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_26_17_y0 ^ f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_25_18_y0;
  assign f_s_dadda_pg_rca32_fa563_y1 = f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_26_17_y0 & f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_25_18_y0;
  assign f_s_dadda_pg_rca32_fa563_y2 = f_s_dadda_pg_rca32_fa563_y0 ^ f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_24_19_y0;
  assign f_s_dadda_pg_rca32_fa563_y3 = f_s_dadda_pg_rca32_fa563_y0 & f_s_dadda_pg_rca32_fa563_f_s_dadda_pg_rca32_and_24_19_y0;
  assign f_s_dadda_pg_rca32_fa563_y4 = f_s_dadda_pg_rca32_fa563_y1 | f_s_dadda_pg_rca32_fa563_y3;
  assign f_s_dadda_pg_rca32_and_23_20_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_23_20_y0 = f_s_dadda_pg_rca32_and_23_20_a_23 & f_s_dadda_pg_rca32_and_23_20_b_20;
  assign f_s_dadda_pg_rca32_and_22_21_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_22_21_y0 = f_s_dadda_pg_rca32_and_22_21_a_22 & f_s_dadda_pg_rca32_and_22_21_b_21;
  assign f_s_dadda_pg_rca32_and_21_22_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_21_22_y0 = f_s_dadda_pg_rca32_and_21_22_a_21 & f_s_dadda_pg_rca32_and_21_22_b_22;
  assign f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_23_20_y0 = f_s_dadda_pg_rca32_and_23_20_y0;
  assign f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_22_21_y0 = f_s_dadda_pg_rca32_and_22_21_y0;
  assign f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_21_22_y0 = f_s_dadda_pg_rca32_and_21_22_y0;
  assign f_s_dadda_pg_rca32_fa564_y0 = f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_23_20_y0 ^ f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_22_21_y0;
  assign f_s_dadda_pg_rca32_fa564_y1 = f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_23_20_y0 & f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_22_21_y0;
  assign f_s_dadda_pg_rca32_fa564_y2 = f_s_dadda_pg_rca32_fa564_y0 ^ f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_21_22_y0;
  assign f_s_dadda_pg_rca32_fa564_y3 = f_s_dadda_pg_rca32_fa564_y0 & f_s_dadda_pg_rca32_fa564_f_s_dadda_pg_rca32_and_21_22_y0;
  assign f_s_dadda_pg_rca32_fa564_y4 = f_s_dadda_pg_rca32_fa564_y1 | f_s_dadda_pg_rca32_fa564_y3;
  assign f_s_dadda_pg_rca32_and_20_23_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_20_23_y0 = f_s_dadda_pg_rca32_and_20_23_a_20 & f_s_dadda_pg_rca32_and_20_23_b_23;
  assign f_s_dadda_pg_rca32_and_19_24_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_19_24_y0 = f_s_dadda_pg_rca32_and_19_24_a_19 & f_s_dadda_pg_rca32_and_19_24_b_24;
  assign f_s_dadda_pg_rca32_and_18_25_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_18_25_y0 = f_s_dadda_pg_rca32_and_18_25_a_18 & f_s_dadda_pg_rca32_and_18_25_b_25;
  assign f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_20_23_y0 = f_s_dadda_pg_rca32_and_20_23_y0;
  assign f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_19_24_y0 = f_s_dadda_pg_rca32_and_19_24_y0;
  assign f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_18_25_y0 = f_s_dadda_pg_rca32_and_18_25_y0;
  assign f_s_dadda_pg_rca32_fa565_y0 = f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_20_23_y0 ^ f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_19_24_y0;
  assign f_s_dadda_pg_rca32_fa565_y1 = f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_20_23_y0 & f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_19_24_y0;
  assign f_s_dadda_pg_rca32_fa565_y2 = f_s_dadda_pg_rca32_fa565_y0 ^ f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_18_25_y0;
  assign f_s_dadda_pg_rca32_fa565_y3 = f_s_dadda_pg_rca32_fa565_y0 & f_s_dadda_pg_rca32_fa565_f_s_dadda_pg_rca32_and_18_25_y0;
  assign f_s_dadda_pg_rca32_fa565_y4 = f_s_dadda_pg_rca32_fa565_y1 | f_s_dadda_pg_rca32_fa565_y3;
  assign f_s_dadda_pg_rca32_and_17_26_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_17_26_y0 = f_s_dadda_pg_rca32_and_17_26_a_17 & f_s_dadda_pg_rca32_and_17_26_b_26;
  assign f_s_dadda_pg_rca32_and_16_27_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_16_27_y0 = f_s_dadda_pg_rca32_and_16_27_a_16 & f_s_dadda_pg_rca32_and_16_27_b_27;
  assign f_s_dadda_pg_rca32_and_15_28_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_15_28_y0 = f_s_dadda_pg_rca32_and_15_28_a_15 & f_s_dadda_pg_rca32_and_15_28_b_28;
  assign f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_17_26_y0 = f_s_dadda_pg_rca32_and_17_26_y0;
  assign f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_16_27_y0 = f_s_dadda_pg_rca32_and_16_27_y0;
  assign f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_15_28_y0 = f_s_dadda_pg_rca32_and_15_28_y0;
  assign f_s_dadda_pg_rca32_fa566_y0 = f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_17_26_y0 ^ f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_16_27_y0;
  assign f_s_dadda_pg_rca32_fa566_y1 = f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_17_26_y0 & f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_16_27_y0;
  assign f_s_dadda_pg_rca32_fa566_y2 = f_s_dadda_pg_rca32_fa566_y0 ^ f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_15_28_y0;
  assign f_s_dadda_pg_rca32_fa566_y3 = f_s_dadda_pg_rca32_fa566_y0 & f_s_dadda_pg_rca32_fa566_f_s_dadda_pg_rca32_and_15_28_y0;
  assign f_s_dadda_pg_rca32_fa566_y4 = f_s_dadda_pg_rca32_fa566_y1 | f_s_dadda_pg_rca32_fa566_y3;
  assign f_s_dadda_pg_rca32_and_14_29_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_14_29_y0 = f_s_dadda_pg_rca32_and_14_29_a_14 & f_s_dadda_pg_rca32_and_14_29_b_29;
  assign f_s_dadda_pg_rca32_and_13_30_a_13 = a_13;
  assign f_s_dadda_pg_rca32_and_13_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_13_30_y0 = f_s_dadda_pg_rca32_and_13_30_a_13 & f_s_dadda_pg_rca32_and_13_30_b_30;
  assign f_s_dadda_pg_rca32_nand_12_31_a_12 = a_12;
  assign f_s_dadda_pg_rca32_nand_12_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_12_31_y0 = ~(f_s_dadda_pg_rca32_nand_12_31_a_12 & f_s_dadda_pg_rca32_nand_12_31_b_31);
  assign f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_and_14_29_y0 = f_s_dadda_pg_rca32_and_14_29_y0;
  assign f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_and_13_30_y0 = f_s_dadda_pg_rca32_and_13_30_y0;
  assign f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_nand_12_31_y0 = f_s_dadda_pg_rca32_nand_12_31_y0;
  assign f_s_dadda_pg_rca32_fa567_y0 = f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_and_14_29_y0 ^ f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_and_13_30_y0;
  assign f_s_dadda_pg_rca32_fa567_y1 = f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_and_14_29_y0 & f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_and_13_30_y0;
  assign f_s_dadda_pg_rca32_fa567_y2 = f_s_dadda_pg_rca32_fa567_y0 ^ f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_nand_12_31_y0;
  assign f_s_dadda_pg_rca32_fa567_y3 = f_s_dadda_pg_rca32_fa567_y0 & f_s_dadda_pg_rca32_fa567_f_s_dadda_pg_rca32_nand_12_31_y0;
  assign f_s_dadda_pg_rca32_fa567_y4 = f_s_dadda_pg_rca32_fa567_y1 | f_s_dadda_pg_rca32_fa567_y3;
  assign f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa556_y2 = f_s_dadda_pg_rca32_fa556_y2;
  assign f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa557_y2 = f_s_dadda_pg_rca32_fa557_y2;
  assign f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa558_y2 = f_s_dadda_pg_rca32_fa558_y2;
  assign f_s_dadda_pg_rca32_fa568_y0 = f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa556_y2 ^ f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa557_y2;
  assign f_s_dadda_pg_rca32_fa568_y1 = f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa556_y2 & f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa557_y2;
  assign f_s_dadda_pg_rca32_fa568_y2 = f_s_dadda_pg_rca32_fa568_y0 ^ f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa558_y2;
  assign f_s_dadda_pg_rca32_fa568_y3 = f_s_dadda_pg_rca32_fa568_y0 & f_s_dadda_pg_rca32_fa568_f_s_dadda_pg_rca32_fa558_y2;
  assign f_s_dadda_pg_rca32_fa568_y4 = f_s_dadda_pg_rca32_fa568_y1 | f_s_dadda_pg_rca32_fa568_y3;
  assign f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa559_y2 = f_s_dadda_pg_rca32_fa559_y2;
  assign f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa560_y2 = f_s_dadda_pg_rca32_fa560_y2;
  assign f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa561_y2 = f_s_dadda_pg_rca32_fa561_y2;
  assign f_s_dadda_pg_rca32_fa569_y0 = f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa559_y2 ^ f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa560_y2;
  assign f_s_dadda_pg_rca32_fa569_y1 = f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa559_y2 & f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa560_y2;
  assign f_s_dadda_pg_rca32_fa569_y2 = f_s_dadda_pg_rca32_fa569_y0 ^ f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa561_y2;
  assign f_s_dadda_pg_rca32_fa569_y3 = f_s_dadda_pg_rca32_fa569_y0 & f_s_dadda_pg_rca32_fa569_f_s_dadda_pg_rca32_fa561_y2;
  assign f_s_dadda_pg_rca32_fa569_y4 = f_s_dadda_pg_rca32_fa569_y1 | f_s_dadda_pg_rca32_fa569_y3;
  assign f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa562_y2 = f_s_dadda_pg_rca32_fa562_y2;
  assign f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa563_y2 = f_s_dadda_pg_rca32_fa563_y2;
  assign f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa564_y2 = f_s_dadda_pg_rca32_fa564_y2;
  assign f_s_dadda_pg_rca32_fa570_y0 = f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa562_y2 ^ f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa563_y2;
  assign f_s_dadda_pg_rca32_fa570_y1 = f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa562_y2 & f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa563_y2;
  assign f_s_dadda_pg_rca32_fa570_y2 = f_s_dadda_pg_rca32_fa570_y0 ^ f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa564_y2;
  assign f_s_dadda_pg_rca32_fa570_y3 = f_s_dadda_pg_rca32_fa570_y0 & f_s_dadda_pg_rca32_fa570_f_s_dadda_pg_rca32_fa564_y2;
  assign f_s_dadda_pg_rca32_fa570_y4 = f_s_dadda_pg_rca32_fa570_y1 | f_s_dadda_pg_rca32_fa570_y3;
  assign f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa570_y4 = f_s_dadda_pg_rca32_fa570_y4;
  assign f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa569_y4 = f_s_dadda_pg_rca32_fa569_y4;
  assign f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa568_y4 = f_s_dadda_pg_rca32_fa568_y4;
  assign f_s_dadda_pg_rca32_fa571_y0 = f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa570_y4 ^ f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa569_y4;
  assign f_s_dadda_pg_rca32_fa571_y1 = f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa570_y4 & f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa569_y4;
  assign f_s_dadda_pg_rca32_fa571_y2 = f_s_dadda_pg_rca32_fa571_y0 ^ f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa568_y4;
  assign f_s_dadda_pg_rca32_fa571_y3 = f_s_dadda_pg_rca32_fa571_y0 & f_s_dadda_pg_rca32_fa571_f_s_dadda_pg_rca32_fa568_y4;
  assign f_s_dadda_pg_rca32_fa571_y4 = f_s_dadda_pg_rca32_fa571_y1 | f_s_dadda_pg_rca32_fa571_y3;
  assign f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa567_y4 = f_s_dadda_pg_rca32_fa567_y4;
  assign f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa566_y4 = f_s_dadda_pg_rca32_fa566_y4;
  assign f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa565_y4 = f_s_dadda_pg_rca32_fa565_y4;
  assign f_s_dadda_pg_rca32_fa572_y0 = f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa567_y4 ^ f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa566_y4;
  assign f_s_dadda_pg_rca32_fa572_y1 = f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa567_y4 & f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa566_y4;
  assign f_s_dadda_pg_rca32_fa572_y2 = f_s_dadda_pg_rca32_fa572_y0 ^ f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa565_y4;
  assign f_s_dadda_pg_rca32_fa572_y3 = f_s_dadda_pg_rca32_fa572_y0 & f_s_dadda_pg_rca32_fa572_f_s_dadda_pg_rca32_fa565_y4;
  assign f_s_dadda_pg_rca32_fa572_y4 = f_s_dadda_pg_rca32_fa572_y1 | f_s_dadda_pg_rca32_fa572_y3;
  assign f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa564_y4 = f_s_dadda_pg_rca32_fa564_y4;
  assign f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa563_y4 = f_s_dadda_pg_rca32_fa563_y4;
  assign f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa562_y4 = f_s_dadda_pg_rca32_fa562_y4;
  assign f_s_dadda_pg_rca32_fa573_y0 = f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa564_y4 ^ f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa563_y4;
  assign f_s_dadda_pg_rca32_fa573_y1 = f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa564_y4 & f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa563_y4;
  assign f_s_dadda_pg_rca32_fa573_y2 = f_s_dadda_pg_rca32_fa573_y0 ^ f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa562_y4;
  assign f_s_dadda_pg_rca32_fa573_y3 = f_s_dadda_pg_rca32_fa573_y0 & f_s_dadda_pg_rca32_fa573_f_s_dadda_pg_rca32_fa562_y4;
  assign f_s_dadda_pg_rca32_fa573_y4 = f_s_dadda_pg_rca32_fa573_y1 | f_s_dadda_pg_rca32_fa573_y3;
  assign f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa561_y4 = f_s_dadda_pg_rca32_fa561_y4;
  assign f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa560_y4 = f_s_dadda_pg_rca32_fa560_y4;
  assign f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa559_y4 = f_s_dadda_pg_rca32_fa559_y4;
  assign f_s_dadda_pg_rca32_fa574_y0 = f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa561_y4 ^ f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa560_y4;
  assign f_s_dadda_pg_rca32_fa574_y1 = f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa561_y4 & f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa560_y4;
  assign f_s_dadda_pg_rca32_fa574_y2 = f_s_dadda_pg_rca32_fa574_y0 ^ f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa559_y4;
  assign f_s_dadda_pg_rca32_fa574_y3 = f_s_dadda_pg_rca32_fa574_y0 & f_s_dadda_pg_rca32_fa574_f_s_dadda_pg_rca32_fa559_y4;
  assign f_s_dadda_pg_rca32_fa574_y4 = f_s_dadda_pg_rca32_fa574_y1 | f_s_dadda_pg_rca32_fa574_y3;
  assign f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa558_y4 = f_s_dadda_pg_rca32_fa558_y4;
  assign f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa557_y4 = f_s_dadda_pg_rca32_fa557_y4;
  assign f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa556_y4 = f_s_dadda_pg_rca32_fa556_y4;
  assign f_s_dadda_pg_rca32_fa575_y0 = f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa558_y4 ^ f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa557_y4;
  assign f_s_dadda_pg_rca32_fa575_y1 = f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa558_y4 & f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa557_y4;
  assign f_s_dadda_pg_rca32_fa575_y2 = f_s_dadda_pg_rca32_fa575_y0 ^ f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa556_y4;
  assign f_s_dadda_pg_rca32_fa575_y3 = f_s_dadda_pg_rca32_fa575_y0 & f_s_dadda_pg_rca32_fa575_f_s_dadda_pg_rca32_fa556_y4;
  assign f_s_dadda_pg_rca32_fa575_y4 = f_s_dadda_pg_rca32_fa575_y1 | f_s_dadda_pg_rca32_fa575_y3;
  assign f_s_dadda_pg_rca32_nand_31_13_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_13_b_13 = b_13;
  assign f_s_dadda_pg_rca32_nand_31_13_y0 = ~(f_s_dadda_pg_rca32_nand_31_13_a_31 & f_s_dadda_pg_rca32_nand_31_13_b_13);
  assign f_s_dadda_pg_rca32_and_30_14_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_and_30_14_y0 = f_s_dadda_pg_rca32_and_30_14_a_30 & f_s_dadda_pg_rca32_and_30_14_b_14;
  assign f_s_dadda_pg_rca32_and_29_15_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_29_15_y0 = f_s_dadda_pg_rca32_and_29_15_a_29 & f_s_dadda_pg_rca32_and_29_15_b_15;
  assign f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_nand_31_13_y0 = f_s_dadda_pg_rca32_nand_31_13_y0;
  assign f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_and_30_14_y0 = f_s_dadda_pg_rca32_and_30_14_y0;
  assign f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_and_29_15_y0 = f_s_dadda_pg_rca32_and_29_15_y0;
  assign f_s_dadda_pg_rca32_fa576_y0 = f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_nand_31_13_y0 ^ f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_and_30_14_y0;
  assign f_s_dadda_pg_rca32_fa576_y1 = f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_nand_31_13_y0 & f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_and_30_14_y0;
  assign f_s_dadda_pg_rca32_fa576_y2 = f_s_dadda_pg_rca32_fa576_y0 ^ f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_and_29_15_y0;
  assign f_s_dadda_pg_rca32_fa576_y3 = f_s_dadda_pg_rca32_fa576_y0 & f_s_dadda_pg_rca32_fa576_f_s_dadda_pg_rca32_and_29_15_y0;
  assign f_s_dadda_pg_rca32_fa576_y4 = f_s_dadda_pg_rca32_fa576_y1 | f_s_dadda_pg_rca32_fa576_y3;
  assign f_s_dadda_pg_rca32_and_28_16_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_28_16_y0 = f_s_dadda_pg_rca32_and_28_16_a_28 & f_s_dadda_pg_rca32_and_28_16_b_16;
  assign f_s_dadda_pg_rca32_and_27_17_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_27_17_y0 = f_s_dadda_pg_rca32_and_27_17_a_27 & f_s_dadda_pg_rca32_and_27_17_b_17;
  assign f_s_dadda_pg_rca32_and_26_18_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_26_18_y0 = f_s_dadda_pg_rca32_and_26_18_a_26 & f_s_dadda_pg_rca32_and_26_18_b_18;
  assign f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_28_16_y0 = f_s_dadda_pg_rca32_and_28_16_y0;
  assign f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_27_17_y0 = f_s_dadda_pg_rca32_and_27_17_y0;
  assign f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_26_18_y0 = f_s_dadda_pg_rca32_and_26_18_y0;
  assign f_s_dadda_pg_rca32_fa577_y0 = f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_28_16_y0 ^ f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_27_17_y0;
  assign f_s_dadda_pg_rca32_fa577_y1 = f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_28_16_y0 & f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_27_17_y0;
  assign f_s_dadda_pg_rca32_fa577_y2 = f_s_dadda_pg_rca32_fa577_y0 ^ f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_26_18_y0;
  assign f_s_dadda_pg_rca32_fa577_y3 = f_s_dadda_pg_rca32_fa577_y0 & f_s_dadda_pg_rca32_fa577_f_s_dadda_pg_rca32_and_26_18_y0;
  assign f_s_dadda_pg_rca32_fa577_y4 = f_s_dadda_pg_rca32_fa577_y1 | f_s_dadda_pg_rca32_fa577_y3;
  assign f_s_dadda_pg_rca32_and_25_19_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_25_19_y0 = f_s_dadda_pg_rca32_and_25_19_a_25 & f_s_dadda_pg_rca32_and_25_19_b_19;
  assign f_s_dadda_pg_rca32_and_24_20_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_24_20_y0 = f_s_dadda_pg_rca32_and_24_20_a_24 & f_s_dadda_pg_rca32_and_24_20_b_20;
  assign f_s_dadda_pg_rca32_and_23_21_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_23_21_y0 = f_s_dadda_pg_rca32_and_23_21_a_23 & f_s_dadda_pg_rca32_and_23_21_b_21;
  assign f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_25_19_y0 = f_s_dadda_pg_rca32_and_25_19_y0;
  assign f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_24_20_y0 = f_s_dadda_pg_rca32_and_24_20_y0;
  assign f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_23_21_y0 = f_s_dadda_pg_rca32_and_23_21_y0;
  assign f_s_dadda_pg_rca32_fa578_y0 = f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_25_19_y0 ^ f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_24_20_y0;
  assign f_s_dadda_pg_rca32_fa578_y1 = f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_25_19_y0 & f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_24_20_y0;
  assign f_s_dadda_pg_rca32_fa578_y2 = f_s_dadda_pg_rca32_fa578_y0 ^ f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_23_21_y0;
  assign f_s_dadda_pg_rca32_fa578_y3 = f_s_dadda_pg_rca32_fa578_y0 & f_s_dadda_pg_rca32_fa578_f_s_dadda_pg_rca32_and_23_21_y0;
  assign f_s_dadda_pg_rca32_fa578_y4 = f_s_dadda_pg_rca32_fa578_y1 | f_s_dadda_pg_rca32_fa578_y3;
  assign f_s_dadda_pg_rca32_and_22_22_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_22_22_y0 = f_s_dadda_pg_rca32_and_22_22_a_22 & f_s_dadda_pg_rca32_and_22_22_b_22;
  assign f_s_dadda_pg_rca32_and_21_23_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_21_23_y0 = f_s_dadda_pg_rca32_and_21_23_a_21 & f_s_dadda_pg_rca32_and_21_23_b_23;
  assign f_s_dadda_pg_rca32_and_20_24_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_20_24_y0 = f_s_dadda_pg_rca32_and_20_24_a_20 & f_s_dadda_pg_rca32_and_20_24_b_24;
  assign f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_22_22_y0 = f_s_dadda_pg_rca32_and_22_22_y0;
  assign f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_21_23_y0 = f_s_dadda_pg_rca32_and_21_23_y0;
  assign f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_20_24_y0 = f_s_dadda_pg_rca32_and_20_24_y0;
  assign f_s_dadda_pg_rca32_fa579_y0 = f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_22_22_y0 ^ f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_21_23_y0;
  assign f_s_dadda_pg_rca32_fa579_y1 = f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_22_22_y0 & f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_21_23_y0;
  assign f_s_dadda_pg_rca32_fa579_y2 = f_s_dadda_pg_rca32_fa579_y0 ^ f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_20_24_y0;
  assign f_s_dadda_pg_rca32_fa579_y3 = f_s_dadda_pg_rca32_fa579_y0 & f_s_dadda_pg_rca32_fa579_f_s_dadda_pg_rca32_and_20_24_y0;
  assign f_s_dadda_pg_rca32_fa579_y4 = f_s_dadda_pg_rca32_fa579_y1 | f_s_dadda_pg_rca32_fa579_y3;
  assign f_s_dadda_pg_rca32_and_19_25_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_19_25_y0 = f_s_dadda_pg_rca32_and_19_25_a_19 & f_s_dadda_pg_rca32_and_19_25_b_25;
  assign f_s_dadda_pg_rca32_and_18_26_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_18_26_y0 = f_s_dadda_pg_rca32_and_18_26_a_18 & f_s_dadda_pg_rca32_and_18_26_b_26;
  assign f_s_dadda_pg_rca32_and_17_27_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_17_27_y0 = f_s_dadda_pg_rca32_and_17_27_a_17 & f_s_dadda_pg_rca32_and_17_27_b_27;
  assign f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_19_25_y0 = f_s_dadda_pg_rca32_and_19_25_y0;
  assign f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_18_26_y0 = f_s_dadda_pg_rca32_and_18_26_y0;
  assign f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_17_27_y0 = f_s_dadda_pg_rca32_and_17_27_y0;
  assign f_s_dadda_pg_rca32_fa580_y0 = f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_19_25_y0 ^ f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_18_26_y0;
  assign f_s_dadda_pg_rca32_fa580_y1 = f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_19_25_y0 & f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_18_26_y0;
  assign f_s_dadda_pg_rca32_fa580_y2 = f_s_dadda_pg_rca32_fa580_y0 ^ f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_17_27_y0;
  assign f_s_dadda_pg_rca32_fa580_y3 = f_s_dadda_pg_rca32_fa580_y0 & f_s_dadda_pg_rca32_fa580_f_s_dadda_pg_rca32_and_17_27_y0;
  assign f_s_dadda_pg_rca32_fa580_y4 = f_s_dadda_pg_rca32_fa580_y1 | f_s_dadda_pg_rca32_fa580_y3;
  assign f_s_dadda_pg_rca32_and_16_28_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_16_28_y0 = f_s_dadda_pg_rca32_and_16_28_a_16 & f_s_dadda_pg_rca32_and_16_28_b_28;
  assign f_s_dadda_pg_rca32_and_15_29_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_15_29_y0 = f_s_dadda_pg_rca32_and_15_29_a_15 & f_s_dadda_pg_rca32_and_15_29_b_29;
  assign f_s_dadda_pg_rca32_and_14_30_a_14 = a_14;
  assign f_s_dadda_pg_rca32_and_14_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_14_30_y0 = f_s_dadda_pg_rca32_and_14_30_a_14 & f_s_dadda_pg_rca32_and_14_30_b_30;
  assign f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_16_28_y0 = f_s_dadda_pg_rca32_and_16_28_y0;
  assign f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_15_29_y0 = f_s_dadda_pg_rca32_and_15_29_y0;
  assign f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_14_30_y0 = f_s_dadda_pg_rca32_and_14_30_y0;
  assign f_s_dadda_pg_rca32_fa581_y0 = f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_16_28_y0 ^ f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_15_29_y0;
  assign f_s_dadda_pg_rca32_fa581_y1 = f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_16_28_y0 & f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_15_29_y0;
  assign f_s_dadda_pg_rca32_fa581_y2 = f_s_dadda_pg_rca32_fa581_y0 ^ f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_14_30_y0;
  assign f_s_dadda_pg_rca32_fa581_y3 = f_s_dadda_pg_rca32_fa581_y0 & f_s_dadda_pg_rca32_fa581_f_s_dadda_pg_rca32_and_14_30_y0;
  assign f_s_dadda_pg_rca32_fa581_y4 = f_s_dadda_pg_rca32_fa581_y1 | f_s_dadda_pg_rca32_fa581_y3;
  assign f_s_dadda_pg_rca32_nand_13_31_a_13 = a_13;
  assign f_s_dadda_pg_rca32_nand_13_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_13_31_y0 = ~(f_s_dadda_pg_rca32_nand_13_31_a_13 & f_s_dadda_pg_rca32_nand_13_31_b_31);
  assign f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_nand_13_31_y0 = f_s_dadda_pg_rca32_nand_13_31_y0;
  assign f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_fa571_y2 = f_s_dadda_pg_rca32_fa571_y2;
  assign f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_fa572_y2 = f_s_dadda_pg_rca32_fa572_y2;
  assign f_s_dadda_pg_rca32_fa582_y0 = f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_nand_13_31_y0 ^ f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_fa571_y2;
  assign f_s_dadda_pg_rca32_fa582_y1 = f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_nand_13_31_y0 & f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_fa571_y2;
  assign f_s_dadda_pg_rca32_fa582_y2 = f_s_dadda_pg_rca32_fa582_y0 ^ f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_fa572_y2;
  assign f_s_dadda_pg_rca32_fa582_y3 = f_s_dadda_pg_rca32_fa582_y0 & f_s_dadda_pg_rca32_fa582_f_s_dadda_pg_rca32_fa572_y2;
  assign f_s_dadda_pg_rca32_fa582_y4 = f_s_dadda_pg_rca32_fa582_y1 | f_s_dadda_pg_rca32_fa582_y3;
  assign f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa573_y2 = f_s_dadda_pg_rca32_fa573_y2;
  assign f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa574_y2 = f_s_dadda_pg_rca32_fa574_y2;
  assign f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa575_y2 = f_s_dadda_pg_rca32_fa575_y2;
  assign f_s_dadda_pg_rca32_fa583_y0 = f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa573_y2 ^ f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa574_y2;
  assign f_s_dadda_pg_rca32_fa583_y1 = f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa573_y2 & f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa574_y2;
  assign f_s_dadda_pg_rca32_fa583_y2 = f_s_dadda_pg_rca32_fa583_y0 ^ f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa575_y2;
  assign f_s_dadda_pg_rca32_fa583_y3 = f_s_dadda_pg_rca32_fa583_y0 & f_s_dadda_pg_rca32_fa583_f_s_dadda_pg_rca32_fa575_y2;
  assign f_s_dadda_pg_rca32_fa583_y4 = f_s_dadda_pg_rca32_fa583_y1 | f_s_dadda_pg_rca32_fa583_y3;
  assign f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa576_y2 = f_s_dadda_pg_rca32_fa576_y2;
  assign f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa577_y2 = f_s_dadda_pg_rca32_fa577_y2;
  assign f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa578_y2 = f_s_dadda_pg_rca32_fa578_y2;
  assign f_s_dadda_pg_rca32_fa584_y0 = f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa576_y2 ^ f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa577_y2;
  assign f_s_dadda_pg_rca32_fa584_y1 = f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa576_y2 & f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa577_y2;
  assign f_s_dadda_pg_rca32_fa584_y2 = f_s_dadda_pg_rca32_fa584_y0 ^ f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa578_y2;
  assign f_s_dadda_pg_rca32_fa584_y3 = f_s_dadda_pg_rca32_fa584_y0 & f_s_dadda_pg_rca32_fa584_f_s_dadda_pg_rca32_fa578_y2;
  assign f_s_dadda_pg_rca32_fa584_y4 = f_s_dadda_pg_rca32_fa584_y1 | f_s_dadda_pg_rca32_fa584_y3;
  assign f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa584_y4 = f_s_dadda_pg_rca32_fa584_y4;
  assign f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa583_y4 = f_s_dadda_pg_rca32_fa583_y4;
  assign f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa582_y4 = f_s_dadda_pg_rca32_fa582_y4;
  assign f_s_dadda_pg_rca32_fa585_y0 = f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa584_y4 ^ f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa583_y4;
  assign f_s_dadda_pg_rca32_fa585_y1 = f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa584_y4 & f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa583_y4;
  assign f_s_dadda_pg_rca32_fa585_y2 = f_s_dadda_pg_rca32_fa585_y0 ^ f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa582_y4;
  assign f_s_dadda_pg_rca32_fa585_y3 = f_s_dadda_pg_rca32_fa585_y0 & f_s_dadda_pg_rca32_fa585_f_s_dadda_pg_rca32_fa582_y4;
  assign f_s_dadda_pg_rca32_fa585_y4 = f_s_dadda_pg_rca32_fa585_y1 | f_s_dadda_pg_rca32_fa585_y3;
  assign f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa581_y4 = f_s_dadda_pg_rca32_fa581_y4;
  assign f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa580_y4 = f_s_dadda_pg_rca32_fa580_y4;
  assign f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa579_y4 = f_s_dadda_pg_rca32_fa579_y4;
  assign f_s_dadda_pg_rca32_fa586_y0 = f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa581_y4 ^ f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa580_y4;
  assign f_s_dadda_pg_rca32_fa586_y1 = f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa581_y4 & f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa580_y4;
  assign f_s_dadda_pg_rca32_fa586_y2 = f_s_dadda_pg_rca32_fa586_y0 ^ f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa579_y4;
  assign f_s_dadda_pg_rca32_fa586_y3 = f_s_dadda_pg_rca32_fa586_y0 & f_s_dadda_pg_rca32_fa586_f_s_dadda_pg_rca32_fa579_y4;
  assign f_s_dadda_pg_rca32_fa586_y4 = f_s_dadda_pg_rca32_fa586_y1 | f_s_dadda_pg_rca32_fa586_y3;
  assign f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa578_y4 = f_s_dadda_pg_rca32_fa578_y4;
  assign f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa577_y4 = f_s_dadda_pg_rca32_fa577_y4;
  assign f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa576_y4 = f_s_dadda_pg_rca32_fa576_y4;
  assign f_s_dadda_pg_rca32_fa587_y0 = f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa578_y4 ^ f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa577_y4;
  assign f_s_dadda_pg_rca32_fa587_y1 = f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa578_y4 & f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa577_y4;
  assign f_s_dadda_pg_rca32_fa587_y2 = f_s_dadda_pg_rca32_fa587_y0 ^ f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa576_y4;
  assign f_s_dadda_pg_rca32_fa587_y3 = f_s_dadda_pg_rca32_fa587_y0 & f_s_dadda_pg_rca32_fa587_f_s_dadda_pg_rca32_fa576_y4;
  assign f_s_dadda_pg_rca32_fa587_y4 = f_s_dadda_pg_rca32_fa587_y1 | f_s_dadda_pg_rca32_fa587_y3;
  assign f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa575_y4 = f_s_dadda_pg_rca32_fa575_y4;
  assign f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa574_y4 = f_s_dadda_pg_rca32_fa574_y4;
  assign f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa573_y4 = f_s_dadda_pg_rca32_fa573_y4;
  assign f_s_dadda_pg_rca32_fa588_y0 = f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa575_y4 ^ f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa574_y4;
  assign f_s_dadda_pg_rca32_fa588_y1 = f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa575_y4 & f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa574_y4;
  assign f_s_dadda_pg_rca32_fa588_y2 = f_s_dadda_pg_rca32_fa588_y0 ^ f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa573_y4;
  assign f_s_dadda_pg_rca32_fa588_y3 = f_s_dadda_pg_rca32_fa588_y0 & f_s_dadda_pg_rca32_fa588_f_s_dadda_pg_rca32_fa573_y4;
  assign f_s_dadda_pg_rca32_fa588_y4 = f_s_dadda_pg_rca32_fa588_y1 | f_s_dadda_pg_rca32_fa588_y3;
  assign f_s_dadda_pg_rca32_nand_31_14_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_14_b_14 = b_14;
  assign f_s_dadda_pg_rca32_nand_31_14_y0 = ~(f_s_dadda_pg_rca32_nand_31_14_a_31 & f_s_dadda_pg_rca32_nand_31_14_b_14);
  assign f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_fa572_y4 = f_s_dadda_pg_rca32_fa572_y4;
  assign f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_fa571_y4 = f_s_dadda_pg_rca32_fa571_y4;
  assign f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_nand_31_14_y0 = f_s_dadda_pg_rca32_nand_31_14_y0;
  assign f_s_dadda_pg_rca32_fa589_y0 = f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_fa572_y4 ^ f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_fa571_y4;
  assign f_s_dadda_pg_rca32_fa589_y1 = f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_fa572_y4 & f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_fa571_y4;
  assign f_s_dadda_pg_rca32_fa589_y2 = f_s_dadda_pg_rca32_fa589_y0 ^ f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_nand_31_14_y0;
  assign f_s_dadda_pg_rca32_fa589_y3 = f_s_dadda_pg_rca32_fa589_y0 & f_s_dadda_pg_rca32_fa589_f_s_dadda_pg_rca32_nand_31_14_y0;
  assign f_s_dadda_pg_rca32_fa589_y4 = f_s_dadda_pg_rca32_fa589_y1 | f_s_dadda_pg_rca32_fa589_y3;
  assign f_s_dadda_pg_rca32_and_30_15_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_and_30_15_y0 = f_s_dadda_pg_rca32_and_30_15_a_30 & f_s_dadda_pg_rca32_and_30_15_b_15;
  assign f_s_dadda_pg_rca32_and_29_16_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_29_16_y0 = f_s_dadda_pg_rca32_and_29_16_a_29 & f_s_dadda_pg_rca32_and_29_16_b_16;
  assign f_s_dadda_pg_rca32_and_28_17_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_28_17_y0 = f_s_dadda_pg_rca32_and_28_17_a_28 & f_s_dadda_pg_rca32_and_28_17_b_17;
  assign f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_30_15_y0 = f_s_dadda_pg_rca32_and_30_15_y0;
  assign f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_29_16_y0 = f_s_dadda_pg_rca32_and_29_16_y0;
  assign f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_28_17_y0 = f_s_dadda_pg_rca32_and_28_17_y0;
  assign f_s_dadda_pg_rca32_fa590_y0 = f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_30_15_y0 ^ f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_29_16_y0;
  assign f_s_dadda_pg_rca32_fa590_y1 = f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_30_15_y0 & f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_29_16_y0;
  assign f_s_dadda_pg_rca32_fa590_y2 = f_s_dadda_pg_rca32_fa590_y0 ^ f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_28_17_y0;
  assign f_s_dadda_pg_rca32_fa590_y3 = f_s_dadda_pg_rca32_fa590_y0 & f_s_dadda_pg_rca32_fa590_f_s_dadda_pg_rca32_and_28_17_y0;
  assign f_s_dadda_pg_rca32_fa590_y4 = f_s_dadda_pg_rca32_fa590_y1 | f_s_dadda_pg_rca32_fa590_y3;
  assign f_s_dadda_pg_rca32_and_27_18_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_27_18_y0 = f_s_dadda_pg_rca32_and_27_18_a_27 & f_s_dadda_pg_rca32_and_27_18_b_18;
  assign f_s_dadda_pg_rca32_and_26_19_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_26_19_y0 = f_s_dadda_pg_rca32_and_26_19_a_26 & f_s_dadda_pg_rca32_and_26_19_b_19;
  assign f_s_dadda_pg_rca32_and_25_20_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_25_20_y0 = f_s_dadda_pg_rca32_and_25_20_a_25 & f_s_dadda_pg_rca32_and_25_20_b_20;
  assign f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_27_18_y0 = f_s_dadda_pg_rca32_and_27_18_y0;
  assign f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_26_19_y0 = f_s_dadda_pg_rca32_and_26_19_y0;
  assign f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_25_20_y0 = f_s_dadda_pg_rca32_and_25_20_y0;
  assign f_s_dadda_pg_rca32_fa591_y0 = f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_27_18_y0 ^ f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_26_19_y0;
  assign f_s_dadda_pg_rca32_fa591_y1 = f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_27_18_y0 & f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_26_19_y0;
  assign f_s_dadda_pg_rca32_fa591_y2 = f_s_dadda_pg_rca32_fa591_y0 ^ f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_25_20_y0;
  assign f_s_dadda_pg_rca32_fa591_y3 = f_s_dadda_pg_rca32_fa591_y0 & f_s_dadda_pg_rca32_fa591_f_s_dadda_pg_rca32_and_25_20_y0;
  assign f_s_dadda_pg_rca32_fa591_y4 = f_s_dadda_pg_rca32_fa591_y1 | f_s_dadda_pg_rca32_fa591_y3;
  assign f_s_dadda_pg_rca32_and_24_21_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_24_21_y0 = f_s_dadda_pg_rca32_and_24_21_a_24 & f_s_dadda_pg_rca32_and_24_21_b_21;
  assign f_s_dadda_pg_rca32_and_23_22_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_23_22_y0 = f_s_dadda_pg_rca32_and_23_22_a_23 & f_s_dadda_pg_rca32_and_23_22_b_22;
  assign f_s_dadda_pg_rca32_and_22_23_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_22_23_y0 = f_s_dadda_pg_rca32_and_22_23_a_22 & f_s_dadda_pg_rca32_and_22_23_b_23;
  assign f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_24_21_y0 = f_s_dadda_pg_rca32_and_24_21_y0;
  assign f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_23_22_y0 = f_s_dadda_pg_rca32_and_23_22_y0;
  assign f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_22_23_y0 = f_s_dadda_pg_rca32_and_22_23_y0;
  assign f_s_dadda_pg_rca32_fa592_y0 = f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_24_21_y0 ^ f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_23_22_y0;
  assign f_s_dadda_pg_rca32_fa592_y1 = f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_24_21_y0 & f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_23_22_y0;
  assign f_s_dadda_pg_rca32_fa592_y2 = f_s_dadda_pg_rca32_fa592_y0 ^ f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_22_23_y0;
  assign f_s_dadda_pg_rca32_fa592_y3 = f_s_dadda_pg_rca32_fa592_y0 & f_s_dadda_pg_rca32_fa592_f_s_dadda_pg_rca32_and_22_23_y0;
  assign f_s_dadda_pg_rca32_fa592_y4 = f_s_dadda_pg_rca32_fa592_y1 | f_s_dadda_pg_rca32_fa592_y3;
  assign f_s_dadda_pg_rca32_and_21_24_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_21_24_y0 = f_s_dadda_pg_rca32_and_21_24_a_21 & f_s_dadda_pg_rca32_and_21_24_b_24;
  assign f_s_dadda_pg_rca32_and_20_25_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_20_25_y0 = f_s_dadda_pg_rca32_and_20_25_a_20 & f_s_dadda_pg_rca32_and_20_25_b_25;
  assign f_s_dadda_pg_rca32_and_19_26_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_19_26_y0 = f_s_dadda_pg_rca32_and_19_26_a_19 & f_s_dadda_pg_rca32_and_19_26_b_26;
  assign f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_21_24_y0 = f_s_dadda_pg_rca32_and_21_24_y0;
  assign f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_20_25_y0 = f_s_dadda_pg_rca32_and_20_25_y0;
  assign f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_19_26_y0 = f_s_dadda_pg_rca32_and_19_26_y0;
  assign f_s_dadda_pg_rca32_fa593_y0 = f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_21_24_y0 ^ f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_20_25_y0;
  assign f_s_dadda_pg_rca32_fa593_y1 = f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_21_24_y0 & f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_20_25_y0;
  assign f_s_dadda_pg_rca32_fa593_y2 = f_s_dadda_pg_rca32_fa593_y0 ^ f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_19_26_y0;
  assign f_s_dadda_pg_rca32_fa593_y3 = f_s_dadda_pg_rca32_fa593_y0 & f_s_dadda_pg_rca32_fa593_f_s_dadda_pg_rca32_and_19_26_y0;
  assign f_s_dadda_pg_rca32_fa593_y4 = f_s_dadda_pg_rca32_fa593_y1 | f_s_dadda_pg_rca32_fa593_y3;
  assign f_s_dadda_pg_rca32_and_18_27_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_18_27_y0 = f_s_dadda_pg_rca32_and_18_27_a_18 & f_s_dadda_pg_rca32_and_18_27_b_27;
  assign f_s_dadda_pg_rca32_and_17_28_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_17_28_y0 = f_s_dadda_pg_rca32_and_17_28_a_17 & f_s_dadda_pg_rca32_and_17_28_b_28;
  assign f_s_dadda_pg_rca32_and_16_29_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_16_29_y0 = f_s_dadda_pg_rca32_and_16_29_a_16 & f_s_dadda_pg_rca32_and_16_29_b_29;
  assign f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_18_27_y0 = f_s_dadda_pg_rca32_and_18_27_y0;
  assign f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_17_28_y0 = f_s_dadda_pg_rca32_and_17_28_y0;
  assign f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_16_29_y0 = f_s_dadda_pg_rca32_and_16_29_y0;
  assign f_s_dadda_pg_rca32_fa594_y0 = f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_18_27_y0 ^ f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_17_28_y0;
  assign f_s_dadda_pg_rca32_fa594_y1 = f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_18_27_y0 & f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_17_28_y0;
  assign f_s_dadda_pg_rca32_fa594_y2 = f_s_dadda_pg_rca32_fa594_y0 ^ f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_16_29_y0;
  assign f_s_dadda_pg_rca32_fa594_y3 = f_s_dadda_pg_rca32_fa594_y0 & f_s_dadda_pg_rca32_fa594_f_s_dadda_pg_rca32_and_16_29_y0;
  assign f_s_dadda_pg_rca32_fa594_y4 = f_s_dadda_pg_rca32_fa594_y1 | f_s_dadda_pg_rca32_fa594_y3;
  assign f_s_dadda_pg_rca32_and_15_30_a_15 = a_15;
  assign f_s_dadda_pg_rca32_and_15_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_15_30_y0 = f_s_dadda_pg_rca32_and_15_30_a_15 & f_s_dadda_pg_rca32_and_15_30_b_30;
  assign f_s_dadda_pg_rca32_nand_14_31_a_14 = a_14;
  assign f_s_dadda_pg_rca32_nand_14_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_14_31_y0 = ~(f_s_dadda_pg_rca32_nand_14_31_a_14 & f_s_dadda_pg_rca32_nand_14_31_b_31);
  assign f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_and_15_30_y0 = f_s_dadda_pg_rca32_and_15_30_y0;
  assign f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_nand_14_31_y0 = f_s_dadda_pg_rca32_nand_14_31_y0;
  assign f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_fa585_y2 = f_s_dadda_pg_rca32_fa585_y2;
  assign f_s_dadda_pg_rca32_fa595_y0 = f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_and_15_30_y0 ^ f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_nand_14_31_y0;
  assign f_s_dadda_pg_rca32_fa595_y1 = f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_and_15_30_y0 & f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_nand_14_31_y0;
  assign f_s_dadda_pg_rca32_fa595_y2 = f_s_dadda_pg_rca32_fa595_y0 ^ f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_fa585_y2;
  assign f_s_dadda_pg_rca32_fa595_y3 = f_s_dadda_pg_rca32_fa595_y0 & f_s_dadda_pg_rca32_fa595_f_s_dadda_pg_rca32_fa585_y2;
  assign f_s_dadda_pg_rca32_fa595_y4 = f_s_dadda_pg_rca32_fa595_y1 | f_s_dadda_pg_rca32_fa595_y3;
  assign f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa586_y2 = f_s_dadda_pg_rca32_fa586_y2;
  assign f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa587_y2 = f_s_dadda_pg_rca32_fa587_y2;
  assign f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa588_y2 = f_s_dadda_pg_rca32_fa588_y2;
  assign f_s_dadda_pg_rca32_fa596_y0 = f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa586_y2 ^ f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa587_y2;
  assign f_s_dadda_pg_rca32_fa596_y1 = f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa586_y2 & f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa587_y2;
  assign f_s_dadda_pg_rca32_fa596_y2 = f_s_dadda_pg_rca32_fa596_y0 ^ f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa588_y2;
  assign f_s_dadda_pg_rca32_fa596_y3 = f_s_dadda_pg_rca32_fa596_y0 & f_s_dadda_pg_rca32_fa596_f_s_dadda_pg_rca32_fa588_y2;
  assign f_s_dadda_pg_rca32_fa596_y4 = f_s_dadda_pg_rca32_fa596_y1 | f_s_dadda_pg_rca32_fa596_y3;
  assign f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa589_y2 = f_s_dadda_pg_rca32_fa589_y2;
  assign f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa590_y2 = f_s_dadda_pg_rca32_fa590_y2;
  assign f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa591_y2 = f_s_dadda_pg_rca32_fa591_y2;
  assign f_s_dadda_pg_rca32_fa597_y0 = f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa589_y2 ^ f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa590_y2;
  assign f_s_dadda_pg_rca32_fa597_y1 = f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa589_y2 & f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa590_y2;
  assign f_s_dadda_pg_rca32_fa597_y2 = f_s_dadda_pg_rca32_fa597_y0 ^ f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa591_y2;
  assign f_s_dadda_pg_rca32_fa597_y3 = f_s_dadda_pg_rca32_fa597_y0 & f_s_dadda_pg_rca32_fa597_f_s_dadda_pg_rca32_fa591_y2;
  assign f_s_dadda_pg_rca32_fa597_y4 = f_s_dadda_pg_rca32_fa597_y1 | f_s_dadda_pg_rca32_fa597_y3;
  assign f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa597_y4 = f_s_dadda_pg_rca32_fa597_y4;
  assign f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa596_y4 = f_s_dadda_pg_rca32_fa596_y4;
  assign f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa595_y4 = f_s_dadda_pg_rca32_fa595_y4;
  assign f_s_dadda_pg_rca32_fa598_y0 = f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa597_y4 ^ f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa596_y4;
  assign f_s_dadda_pg_rca32_fa598_y1 = f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa597_y4 & f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa596_y4;
  assign f_s_dadda_pg_rca32_fa598_y2 = f_s_dadda_pg_rca32_fa598_y0 ^ f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa595_y4;
  assign f_s_dadda_pg_rca32_fa598_y3 = f_s_dadda_pg_rca32_fa598_y0 & f_s_dadda_pg_rca32_fa598_f_s_dadda_pg_rca32_fa595_y4;
  assign f_s_dadda_pg_rca32_fa598_y4 = f_s_dadda_pg_rca32_fa598_y1 | f_s_dadda_pg_rca32_fa598_y3;
  assign f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa594_y4 = f_s_dadda_pg_rca32_fa594_y4;
  assign f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa593_y4 = f_s_dadda_pg_rca32_fa593_y4;
  assign f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa592_y4 = f_s_dadda_pg_rca32_fa592_y4;
  assign f_s_dadda_pg_rca32_fa599_y0 = f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa594_y4 ^ f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa593_y4;
  assign f_s_dadda_pg_rca32_fa599_y1 = f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa594_y4 & f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa593_y4;
  assign f_s_dadda_pg_rca32_fa599_y2 = f_s_dadda_pg_rca32_fa599_y0 ^ f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa592_y4;
  assign f_s_dadda_pg_rca32_fa599_y3 = f_s_dadda_pg_rca32_fa599_y0 & f_s_dadda_pg_rca32_fa599_f_s_dadda_pg_rca32_fa592_y4;
  assign f_s_dadda_pg_rca32_fa599_y4 = f_s_dadda_pg_rca32_fa599_y1 | f_s_dadda_pg_rca32_fa599_y3;
  assign f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa591_y4 = f_s_dadda_pg_rca32_fa591_y4;
  assign f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa590_y4 = f_s_dadda_pg_rca32_fa590_y4;
  assign f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa589_y4 = f_s_dadda_pg_rca32_fa589_y4;
  assign f_s_dadda_pg_rca32_fa600_y0 = f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa591_y4 ^ f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa590_y4;
  assign f_s_dadda_pg_rca32_fa600_y1 = f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa591_y4 & f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa590_y4;
  assign f_s_dadda_pg_rca32_fa600_y2 = f_s_dadda_pg_rca32_fa600_y0 ^ f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa589_y4;
  assign f_s_dadda_pg_rca32_fa600_y3 = f_s_dadda_pg_rca32_fa600_y0 & f_s_dadda_pg_rca32_fa600_f_s_dadda_pg_rca32_fa589_y4;
  assign f_s_dadda_pg_rca32_fa600_y4 = f_s_dadda_pg_rca32_fa600_y1 | f_s_dadda_pg_rca32_fa600_y3;
  assign f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa588_y4 = f_s_dadda_pg_rca32_fa588_y4;
  assign f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa587_y4 = f_s_dadda_pg_rca32_fa587_y4;
  assign f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa586_y4 = f_s_dadda_pg_rca32_fa586_y4;
  assign f_s_dadda_pg_rca32_fa601_y0 = f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa588_y4 ^ f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa587_y4;
  assign f_s_dadda_pg_rca32_fa601_y1 = f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa588_y4 & f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa587_y4;
  assign f_s_dadda_pg_rca32_fa601_y2 = f_s_dadda_pg_rca32_fa601_y0 ^ f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa586_y4;
  assign f_s_dadda_pg_rca32_fa601_y3 = f_s_dadda_pg_rca32_fa601_y0 & f_s_dadda_pg_rca32_fa601_f_s_dadda_pg_rca32_fa586_y4;
  assign f_s_dadda_pg_rca32_fa601_y4 = f_s_dadda_pg_rca32_fa601_y1 | f_s_dadda_pg_rca32_fa601_y3;
  assign f_s_dadda_pg_rca32_nand_31_15_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_15_b_15 = b_15;
  assign f_s_dadda_pg_rca32_nand_31_15_y0 = ~(f_s_dadda_pg_rca32_nand_31_15_a_31 & f_s_dadda_pg_rca32_nand_31_15_b_15);
  assign f_s_dadda_pg_rca32_and_30_16_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_and_30_16_y0 = f_s_dadda_pg_rca32_and_30_16_a_30 & f_s_dadda_pg_rca32_and_30_16_b_16;
  assign f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_fa585_y4 = f_s_dadda_pg_rca32_fa585_y4;
  assign f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_nand_31_15_y0 = f_s_dadda_pg_rca32_nand_31_15_y0;
  assign f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_and_30_16_y0 = f_s_dadda_pg_rca32_and_30_16_y0;
  assign f_s_dadda_pg_rca32_fa602_y0 = f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_fa585_y4 ^ f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_nand_31_15_y0;
  assign f_s_dadda_pg_rca32_fa602_y1 = f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_fa585_y4 & f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_nand_31_15_y0;
  assign f_s_dadda_pg_rca32_fa602_y2 = f_s_dadda_pg_rca32_fa602_y0 ^ f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_and_30_16_y0;
  assign f_s_dadda_pg_rca32_fa602_y3 = f_s_dadda_pg_rca32_fa602_y0 & f_s_dadda_pg_rca32_fa602_f_s_dadda_pg_rca32_and_30_16_y0;
  assign f_s_dadda_pg_rca32_fa602_y4 = f_s_dadda_pg_rca32_fa602_y1 | f_s_dadda_pg_rca32_fa602_y3;
  assign f_s_dadda_pg_rca32_and_29_17_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_29_17_y0 = f_s_dadda_pg_rca32_and_29_17_a_29 & f_s_dadda_pg_rca32_and_29_17_b_17;
  assign f_s_dadda_pg_rca32_and_28_18_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_28_18_y0 = f_s_dadda_pg_rca32_and_28_18_a_28 & f_s_dadda_pg_rca32_and_28_18_b_18;
  assign f_s_dadda_pg_rca32_and_27_19_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_27_19_y0 = f_s_dadda_pg_rca32_and_27_19_a_27 & f_s_dadda_pg_rca32_and_27_19_b_19;
  assign f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_29_17_y0 = f_s_dadda_pg_rca32_and_29_17_y0;
  assign f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_28_18_y0 = f_s_dadda_pg_rca32_and_28_18_y0;
  assign f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_27_19_y0 = f_s_dadda_pg_rca32_and_27_19_y0;
  assign f_s_dadda_pg_rca32_fa603_y0 = f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_29_17_y0 ^ f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_28_18_y0;
  assign f_s_dadda_pg_rca32_fa603_y1 = f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_29_17_y0 & f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_28_18_y0;
  assign f_s_dadda_pg_rca32_fa603_y2 = f_s_dadda_pg_rca32_fa603_y0 ^ f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_27_19_y0;
  assign f_s_dadda_pg_rca32_fa603_y3 = f_s_dadda_pg_rca32_fa603_y0 & f_s_dadda_pg_rca32_fa603_f_s_dadda_pg_rca32_and_27_19_y0;
  assign f_s_dadda_pg_rca32_fa603_y4 = f_s_dadda_pg_rca32_fa603_y1 | f_s_dadda_pg_rca32_fa603_y3;
  assign f_s_dadda_pg_rca32_and_26_20_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_26_20_y0 = f_s_dadda_pg_rca32_and_26_20_a_26 & f_s_dadda_pg_rca32_and_26_20_b_20;
  assign f_s_dadda_pg_rca32_and_25_21_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_25_21_y0 = f_s_dadda_pg_rca32_and_25_21_a_25 & f_s_dadda_pg_rca32_and_25_21_b_21;
  assign f_s_dadda_pg_rca32_and_24_22_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_24_22_y0 = f_s_dadda_pg_rca32_and_24_22_a_24 & f_s_dadda_pg_rca32_and_24_22_b_22;
  assign f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_26_20_y0 = f_s_dadda_pg_rca32_and_26_20_y0;
  assign f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_25_21_y0 = f_s_dadda_pg_rca32_and_25_21_y0;
  assign f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_24_22_y0 = f_s_dadda_pg_rca32_and_24_22_y0;
  assign f_s_dadda_pg_rca32_fa604_y0 = f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_26_20_y0 ^ f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_25_21_y0;
  assign f_s_dadda_pg_rca32_fa604_y1 = f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_26_20_y0 & f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_25_21_y0;
  assign f_s_dadda_pg_rca32_fa604_y2 = f_s_dadda_pg_rca32_fa604_y0 ^ f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_24_22_y0;
  assign f_s_dadda_pg_rca32_fa604_y3 = f_s_dadda_pg_rca32_fa604_y0 & f_s_dadda_pg_rca32_fa604_f_s_dadda_pg_rca32_and_24_22_y0;
  assign f_s_dadda_pg_rca32_fa604_y4 = f_s_dadda_pg_rca32_fa604_y1 | f_s_dadda_pg_rca32_fa604_y3;
  assign f_s_dadda_pg_rca32_and_23_23_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_23_23_y0 = f_s_dadda_pg_rca32_and_23_23_a_23 & f_s_dadda_pg_rca32_and_23_23_b_23;
  assign f_s_dadda_pg_rca32_and_22_24_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_22_24_y0 = f_s_dadda_pg_rca32_and_22_24_a_22 & f_s_dadda_pg_rca32_and_22_24_b_24;
  assign f_s_dadda_pg_rca32_and_21_25_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_21_25_y0 = f_s_dadda_pg_rca32_and_21_25_a_21 & f_s_dadda_pg_rca32_and_21_25_b_25;
  assign f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_23_23_y0 = f_s_dadda_pg_rca32_and_23_23_y0;
  assign f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_22_24_y0 = f_s_dadda_pg_rca32_and_22_24_y0;
  assign f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_21_25_y0 = f_s_dadda_pg_rca32_and_21_25_y0;
  assign f_s_dadda_pg_rca32_fa605_y0 = f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_23_23_y0 ^ f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_22_24_y0;
  assign f_s_dadda_pg_rca32_fa605_y1 = f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_23_23_y0 & f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_22_24_y0;
  assign f_s_dadda_pg_rca32_fa605_y2 = f_s_dadda_pg_rca32_fa605_y0 ^ f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_21_25_y0;
  assign f_s_dadda_pg_rca32_fa605_y3 = f_s_dadda_pg_rca32_fa605_y0 & f_s_dadda_pg_rca32_fa605_f_s_dadda_pg_rca32_and_21_25_y0;
  assign f_s_dadda_pg_rca32_fa605_y4 = f_s_dadda_pg_rca32_fa605_y1 | f_s_dadda_pg_rca32_fa605_y3;
  assign f_s_dadda_pg_rca32_and_20_26_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_20_26_y0 = f_s_dadda_pg_rca32_and_20_26_a_20 & f_s_dadda_pg_rca32_and_20_26_b_26;
  assign f_s_dadda_pg_rca32_and_19_27_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_19_27_y0 = f_s_dadda_pg_rca32_and_19_27_a_19 & f_s_dadda_pg_rca32_and_19_27_b_27;
  assign f_s_dadda_pg_rca32_and_18_28_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_18_28_y0 = f_s_dadda_pg_rca32_and_18_28_a_18 & f_s_dadda_pg_rca32_and_18_28_b_28;
  assign f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_20_26_y0 = f_s_dadda_pg_rca32_and_20_26_y0;
  assign f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_19_27_y0 = f_s_dadda_pg_rca32_and_19_27_y0;
  assign f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_18_28_y0 = f_s_dadda_pg_rca32_and_18_28_y0;
  assign f_s_dadda_pg_rca32_fa606_y0 = f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_20_26_y0 ^ f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_19_27_y0;
  assign f_s_dadda_pg_rca32_fa606_y1 = f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_20_26_y0 & f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_19_27_y0;
  assign f_s_dadda_pg_rca32_fa606_y2 = f_s_dadda_pg_rca32_fa606_y0 ^ f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_18_28_y0;
  assign f_s_dadda_pg_rca32_fa606_y3 = f_s_dadda_pg_rca32_fa606_y0 & f_s_dadda_pg_rca32_fa606_f_s_dadda_pg_rca32_and_18_28_y0;
  assign f_s_dadda_pg_rca32_fa606_y4 = f_s_dadda_pg_rca32_fa606_y1 | f_s_dadda_pg_rca32_fa606_y3;
  assign f_s_dadda_pg_rca32_and_17_29_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_17_29_y0 = f_s_dadda_pg_rca32_and_17_29_a_17 & f_s_dadda_pg_rca32_and_17_29_b_29;
  assign f_s_dadda_pg_rca32_and_16_30_a_16 = a_16;
  assign f_s_dadda_pg_rca32_and_16_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_16_30_y0 = f_s_dadda_pg_rca32_and_16_30_a_16 & f_s_dadda_pg_rca32_and_16_30_b_30;
  assign f_s_dadda_pg_rca32_nand_15_31_a_15 = a_15;
  assign f_s_dadda_pg_rca32_nand_15_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_15_31_y0 = ~(f_s_dadda_pg_rca32_nand_15_31_a_15 & f_s_dadda_pg_rca32_nand_15_31_b_31);
  assign f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_and_17_29_y0 = f_s_dadda_pg_rca32_and_17_29_y0;
  assign f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_and_16_30_y0 = f_s_dadda_pg_rca32_and_16_30_y0;
  assign f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_nand_15_31_y0 = f_s_dadda_pg_rca32_nand_15_31_y0;
  assign f_s_dadda_pg_rca32_fa607_y0 = f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_and_17_29_y0 ^ f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_and_16_30_y0;
  assign f_s_dadda_pg_rca32_fa607_y1 = f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_and_17_29_y0 & f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_and_16_30_y0;
  assign f_s_dadda_pg_rca32_fa607_y2 = f_s_dadda_pg_rca32_fa607_y0 ^ f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_nand_15_31_y0;
  assign f_s_dadda_pg_rca32_fa607_y3 = f_s_dadda_pg_rca32_fa607_y0 & f_s_dadda_pg_rca32_fa607_f_s_dadda_pg_rca32_nand_15_31_y0;
  assign f_s_dadda_pg_rca32_fa607_y4 = f_s_dadda_pg_rca32_fa607_y1 | f_s_dadda_pg_rca32_fa607_y3;
  assign f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa598_y2 = f_s_dadda_pg_rca32_fa598_y2;
  assign f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa599_y2 = f_s_dadda_pg_rca32_fa599_y2;
  assign f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa600_y2 = f_s_dadda_pg_rca32_fa600_y2;
  assign f_s_dadda_pg_rca32_fa608_y0 = f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa598_y2 ^ f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa599_y2;
  assign f_s_dadda_pg_rca32_fa608_y1 = f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa598_y2 & f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa599_y2;
  assign f_s_dadda_pg_rca32_fa608_y2 = f_s_dadda_pg_rca32_fa608_y0 ^ f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa600_y2;
  assign f_s_dadda_pg_rca32_fa608_y3 = f_s_dadda_pg_rca32_fa608_y0 & f_s_dadda_pg_rca32_fa608_f_s_dadda_pg_rca32_fa600_y2;
  assign f_s_dadda_pg_rca32_fa608_y4 = f_s_dadda_pg_rca32_fa608_y1 | f_s_dadda_pg_rca32_fa608_y3;
  assign f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa601_y2 = f_s_dadda_pg_rca32_fa601_y2;
  assign f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa602_y2 = f_s_dadda_pg_rca32_fa602_y2;
  assign f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa603_y2 = f_s_dadda_pg_rca32_fa603_y2;
  assign f_s_dadda_pg_rca32_fa609_y0 = f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa601_y2 ^ f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa602_y2;
  assign f_s_dadda_pg_rca32_fa609_y1 = f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa601_y2 & f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa602_y2;
  assign f_s_dadda_pg_rca32_fa609_y2 = f_s_dadda_pg_rca32_fa609_y0 ^ f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa603_y2;
  assign f_s_dadda_pg_rca32_fa609_y3 = f_s_dadda_pg_rca32_fa609_y0 & f_s_dadda_pg_rca32_fa609_f_s_dadda_pg_rca32_fa603_y2;
  assign f_s_dadda_pg_rca32_fa609_y4 = f_s_dadda_pg_rca32_fa609_y1 | f_s_dadda_pg_rca32_fa609_y3;
  assign f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa609_y4 = f_s_dadda_pg_rca32_fa609_y4;
  assign f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa608_y4 = f_s_dadda_pg_rca32_fa608_y4;
  assign f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa607_y4 = f_s_dadda_pg_rca32_fa607_y4;
  assign f_s_dadda_pg_rca32_fa610_y0 = f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa609_y4 ^ f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa608_y4;
  assign f_s_dadda_pg_rca32_fa610_y1 = f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa609_y4 & f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa608_y4;
  assign f_s_dadda_pg_rca32_fa610_y2 = f_s_dadda_pg_rca32_fa610_y0 ^ f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa607_y4;
  assign f_s_dadda_pg_rca32_fa610_y3 = f_s_dadda_pg_rca32_fa610_y0 & f_s_dadda_pg_rca32_fa610_f_s_dadda_pg_rca32_fa607_y4;
  assign f_s_dadda_pg_rca32_fa610_y4 = f_s_dadda_pg_rca32_fa610_y1 | f_s_dadda_pg_rca32_fa610_y3;
  assign f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa606_y4 = f_s_dadda_pg_rca32_fa606_y4;
  assign f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa605_y4 = f_s_dadda_pg_rca32_fa605_y4;
  assign f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa604_y4 = f_s_dadda_pg_rca32_fa604_y4;
  assign f_s_dadda_pg_rca32_fa611_y0 = f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa606_y4 ^ f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa605_y4;
  assign f_s_dadda_pg_rca32_fa611_y1 = f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa606_y4 & f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa605_y4;
  assign f_s_dadda_pg_rca32_fa611_y2 = f_s_dadda_pg_rca32_fa611_y0 ^ f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa604_y4;
  assign f_s_dadda_pg_rca32_fa611_y3 = f_s_dadda_pg_rca32_fa611_y0 & f_s_dadda_pg_rca32_fa611_f_s_dadda_pg_rca32_fa604_y4;
  assign f_s_dadda_pg_rca32_fa611_y4 = f_s_dadda_pg_rca32_fa611_y1 | f_s_dadda_pg_rca32_fa611_y3;
  assign f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa603_y4 = f_s_dadda_pg_rca32_fa603_y4;
  assign f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa602_y4 = f_s_dadda_pg_rca32_fa602_y4;
  assign f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa601_y4 = f_s_dadda_pg_rca32_fa601_y4;
  assign f_s_dadda_pg_rca32_fa612_y0 = f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa603_y4 ^ f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa602_y4;
  assign f_s_dadda_pg_rca32_fa612_y1 = f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa603_y4 & f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa602_y4;
  assign f_s_dadda_pg_rca32_fa612_y2 = f_s_dadda_pg_rca32_fa612_y0 ^ f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa601_y4;
  assign f_s_dadda_pg_rca32_fa612_y3 = f_s_dadda_pg_rca32_fa612_y0 & f_s_dadda_pg_rca32_fa612_f_s_dadda_pg_rca32_fa601_y4;
  assign f_s_dadda_pg_rca32_fa612_y4 = f_s_dadda_pg_rca32_fa612_y1 | f_s_dadda_pg_rca32_fa612_y3;
  assign f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa600_y4 = f_s_dadda_pg_rca32_fa600_y4;
  assign f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa599_y4 = f_s_dadda_pg_rca32_fa599_y4;
  assign f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa598_y4 = f_s_dadda_pg_rca32_fa598_y4;
  assign f_s_dadda_pg_rca32_fa613_y0 = f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa600_y4 ^ f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa599_y4;
  assign f_s_dadda_pg_rca32_fa613_y1 = f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa600_y4 & f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa599_y4;
  assign f_s_dadda_pg_rca32_fa613_y2 = f_s_dadda_pg_rca32_fa613_y0 ^ f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa598_y4;
  assign f_s_dadda_pg_rca32_fa613_y3 = f_s_dadda_pg_rca32_fa613_y0 & f_s_dadda_pg_rca32_fa613_f_s_dadda_pg_rca32_fa598_y4;
  assign f_s_dadda_pg_rca32_fa613_y4 = f_s_dadda_pg_rca32_fa613_y1 | f_s_dadda_pg_rca32_fa613_y3;
  assign f_s_dadda_pg_rca32_nand_31_16_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_16_b_16 = b_16;
  assign f_s_dadda_pg_rca32_nand_31_16_y0 = ~(f_s_dadda_pg_rca32_nand_31_16_a_31 & f_s_dadda_pg_rca32_nand_31_16_b_16);
  assign f_s_dadda_pg_rca32_and_30_17_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_and_30_17_y0 = f_s_dadda_pg_rca32_and_30_17_a_30 & f_s_dadda_pg_rca32_and_30_17_b_17;
  assign f_s_dadda_pg_rca32_and_29_18_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_29_18_y0 = f_s_dadda_pg_rca32_and_29_18_a_29 & f_s_dadda_pg_rca32_and_29_18_b_18;
  assign f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_nand_31_16_y0 = f_s_dadda_pg_rca32_nand_31_16_y0;
  assign f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_and_30_17_y0 = f_s_dadda_pg_rca32_and_30_17_y0;
  assign f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_and_29_18_y0 = f_s_dadda_pg_rca32_and_29_18_y0;
  assign f_s_dadda_pg_rca32_fa614_y0 = f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_nand_31_16_y0 ^ f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_and_30_17_y0;
  assign f_s_dadda_pg_rca32_fa614_y1 = f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_nand_31_16_y0 & f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_and_30_17_y0;
  assign f_s_dadda_pg_rca32_fa614_y2 = f_s_dadda_pg_rca32_fa614_y0 ^ f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_and_29_18_y0;
  assign f_s_dadda_pg_rca32_fa614_y3 = f_s_dadda_pg_rca32_fa614_y0 & f_s_dadda_pg_rca32_fa614_f_s_dadda_pg_rca32_and_29_18_y0;
  assign f_s_dadda_pg_rca32_fa614_y4 = f_s_dadda_pg_rca32_fa614_y1 | f_s_dadda_pg_rca32_fa614_y3;
  assign f_s_dadda_pg_rca32_and_28_19_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_28_19_y0 = f_s_dadda_pg_rca32_and_28_19_a_28 & f_s_dadda_pg_rca32_and_28_19_b_19;
  assign f_s_dadda_pg_rca32_and_27_20_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_27_20_y0 = f_s_dadda_pg_rca32_and_27_20_a_27 & f_s_dadda_pg_rca32_and_27_20_b_20;
  assign f_s_dadda_pg_rca32_and_26_21_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_26_21_y0 = f_s_dadda_pg_rca32_and_26_21_a_26 & f_s_dadda_pg_rca32_and_26_21_b_21;
  assign f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_28_19_y0 = f_s_dadda_pg_rca32_and_28_19_y0;
  assign f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_27_20_y0 = f_s_dadda_pg_rca32_and_27_20_y0;
  assign f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_26_21_y0 = f_s_dadda_pg_rca32_and_26_21_y0;
  assign f_s_dadda_pg_rca32_fa615_y0 = f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_28_19_y0 ^ f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_27_20_y0;
  assign f_s_dadda_pg_rca32_fa615_y1 = f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_28_19_y0 & f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_27_20_y0;
  assign f_s_dadda_pg_rca32_fa615_y2 = f_s_dadda_pg_rca32_fa615_y0 ^ f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_26_21_y0;
  assign f_s_dadda_pg_rca32_fa615_y3 = f_s_dadda_pg_rca32_fa615_y0 & f_s_dadda_pg_rca32_fa615_f_s_dadda_pg_rca32_and_26_21_y0;
  assign f_s_dadda_pg_rca32_fa615_y4 = f_s_dadda_pg_rca32_fa615_y1 | f_s_dadda_pg_rca32_fa615_y3;
  assign f_s_dadda_pg_rca32_and_25_22_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_25_22_y0 = f_s_dadda_pg_rca32_and_25_22_a_25 & f_s_dadda_pg_rca32_and_25_22_b_22;
  assign f_s_dadda_pg_rca32_and_24_23_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_24_23_y0 = f_s_dadda_pg_rca32_and_24_23_a_24 & f_s_dadda_pg_rca32_and_24_23_b_23;
  assign f_s_dadda_pg_rca32_and_23_24_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_23_24_y0 = f_s_dadda_pg_rca32_and_23_24_a_23 & f_s_dadda_pg_rca32_and_23_24_b_24;
  assign f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_25_22_y0 = f_s_dadda_pg_rca32_and_25_22_y0;
  assign f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_24_23_y0 = f_s_dadda_pg_rca32_and_24_23_y0;
  assign f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_23_24_y0 = f_s_dadda_pg_rca32_and_23_24_y0;
  assign f_s_dadda_pg_rca32_fa616_y0 = f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_25_22_y0 ^ f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_24_23_y0;
  assign f_s_dadda_pg_rca32_fa616_y1 = f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_25_22_y0 & f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_24_23_y0;
  assign f_s_dadda_pg_rca32_fa616_y2 = f_s_dadda_pg_rca32_fa616_y0 ^ f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_23_24_y0;
  assign f_s_dadda_pg_rca32_fa616_y3 = f_s_dadda_pg_rca32_fa616_y0 & f_s_dadda_pg_rca32_fa616_f_s_dadda_pg_rca32_and_23_24_y0;
  assign f_s_dadda_pg_rca32_fa616_y4 = f_s_dadda_pg_rca32_fa616_y1 | f_s_dadda_pg_rca32_fa616_y3;
  assign f_s_dadda_pg_rca32_and_22_25_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_22_25_y0 = f_s_dadda_pg_rca32_and_22_25_a_22 & f_s_dadda_pg_rca32_and_22_25_b_25;
  assign f_s_dadda_pg_rca32_and_21_26_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_21_26_y0 = f_s_dadda_pg_rca32_and_21_26_a_21 & f_s_dadda_pg_rca32_and_21_26_b_26;
  assign f_s_dadda_pg_rca32_and_20_27_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_20_27_y0 = f_s_dadda_pg_rca32_and_20_27_a_20 & f_s_dadda_pg_rca32_and_20_27_b_27;
  assign f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_22_25_y0 = f_s_dadda_pg_rca32_and_22_25_y0;
  assign f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_21_26_y0 = f_s_dadda_pg_rca32_and_21_26_y0;
  assign f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_20_27_y0 = f_s_dadda_pg_rca32_and_20_27_y0;
  assign f_s_dadda_pg_rca32_fa617_y0 = f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_22_25_y0 ^ f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_21_26_y0;
  assign f_s_dadda_pg_rca32_fa617_y1 = f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_22_25_y0 & f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_21_26_y0;
  assign f_s_dadda_pg_rca32_fa617_y2 = f_s_dadda_pg_rca32_fa617_y0 ^ f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_20_27_y0;
  assign f_s_dadda_pg_rca32_fa617_y3 = f_s_dadda_pg_rca32_fa617_y0 & f_s_dadda_pg_rca32_fa617_f_s_dadda_pg_rca32_and_20_27_y0;
  assign f_s_dadda_pg_rca32_fa617_y4 = f_s_dadda_pg_rca32_fa617_y1 | f_s_dadda_pg_rca32_fa617_y3;
  assign f_s_dadda_pg_rca32_and_19_28_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_19_28_y0 = f_s_dadda_pg_rca32_and_19_28_a_19 & f_s_dadda_pg_rca32_and_19_28_b_28;
  assign f_s_dadda_pg_rca32_and_18_29_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_18_29_y0 = f_s_dadda_pg_rca32_and_18_29_a_18 & f_s_dadda_pg_rca32_and_18_29_b_29;
  assign f_s_dadda_pg_rca32_and_17_30_a_17 = a_17;
  assign f_s_dadda_pg_rca32_and_17_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_17_30_y0 = f_s_dadda_pg_rca32_and_17_30_a_17 & f_s_dadda_pg_rca32_and_17_30_b_30;
  assign f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_19_28_y0 = f_s_dadda_pg_rca32_and_19_28_y0;
  assign f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_18_29_y0 = f_s_dadda_pg_rca32_and_18_29_y0;
  assign f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_17_30_y0 = f_s_dadda_pg_rca32_and_17_30_y0;
  assign f_s_dadda_pg_rca32_fa618_y0 = f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_19_28_y0 ^ f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_18_29_y0;
  assign f_s_dadda_pg_rca32_fa618_y1 = f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_19_28_y0 & f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_18_29_y0;
  assign f_s_dadda_pg_rca32_fa618_y2 = f_s_dadda_pg_rca32_fa618_y0 ^ f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_17_30_y0;
  assign f_s_dadda_pg_rca32_fa618_y3 = f_s_dadda_pg_rca32_fa618_y0 & f_s_dadda_pg_rca32_fa618_f_s_dadda_pg_rca32_and_17_30_y0;
  assign f_s_dadda_pg_rca32_fa618_y4 = f_s_dadda_pg_rca32_fa618_y1 | f_s_dadda_pg_rca32_fa618_y3;
  assign f_s_dadda_pg_rca32_nand_16_31_a_16 = a_16;
  assign f_s_dadda_pg_rca32_nand_16_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_16_31_y0 = ~(f_s_dadda_pg_rca32_nand_16_31_a_16 & f_s_dadda_pg_rca32_nand_16_31_b_31);
  assign f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_nand_16_31_y0 = f_s_dadda_pg_rca32_nand_16_31_y0;
  assign f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_fa610_y2 = f_s_dadda_pg_rca32_fa610_y2;
  assign f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_fa611_y2 = f_s_dadda_pg_rca32_fa611_y2;
  assign f_s_dadda_pg_rca32_fa619_y0 = f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_nand_16_31_y0 ^ f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_fa610_y2;
  assign f_s_dadda_pg_rca32_fa619_y1 = f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_nand_16_31_y0 & f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_fa610_y2;
  assign f_s_dadda_pg_rca32_fa619_y2 = f_s_dadda_pg_rca32_fa619_y0 ^ f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_fa611_y2;
  assign f_s_dadda_pg_rca32_fa619_y3 = f_s_dadda_pg_rca32_fa619_y0 & f_s_dadda_pg_rca32_fa619_f_s_dadda_pg_rca32_fa611_y2;
  assign f_s_dadda_pg_rca32_fa619_y4 = f_s_dadda_pg_rca32_fa619_y1 | f_s_dadda_pg_rca32_fa619_y3;
  assign f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa612_y2 = f_s_dadda_pg_rca32_fa612_y2;
  assign f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa613_y2 = f_s_dadda_pg_rca32_fa613_y2;
  assign f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa614_y2 = f_s_dadda_pg_rca32_fa614_y2;
  assign f_s_dadda_pg_rca32_fa620_y0 = f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa612_y2 ^ f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa613_y2;
  assign f_s_dadda_pg_rca32_fa620_y1 = f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa612_y2 & f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa613_y2;
  assign f_s_dadda_pg_rca32_fa620_y2 = f_s_dadda_pg_rca32_fa620_y0 ^ f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa614_y2;
  assign f_s_dadda_pg_rca32_fa620_y3 = f_s_dadda_pg_rca32_fa620_y0 & f_s_dadda_pg_rca32_fa620_f_s_dadda_pg_rca32_fa614_y2;
  assign f_s_dadda_pg_rca32_fa620_y4 = f_s_dadda_pg_rca32_fa620_y1 | f_s_dadda_pg_rca32_fa620_y3;
  assign f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa620_y4 = f_s_dadda_pg_rca32_fa620_y4;
  assign f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa619_y4 = f_s_dadda_pg_rca32_fa619_y4;
  assign f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa618_y4 = f_s_dadda_pg_rca32_fa618_y4;
  assign f_s_dadda_pg_rca32_fa621_y0 = f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa620_y4 ^ f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa619_y4;
  assign f_s_dadda_pg_rca32_fa621_y1 = f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa620_y4 & f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa619_y4;
  assign f_s_dadda_pg_rca32_fa621_y2 = f_s_dadda_pg_rca32_fa621_y0 ^ f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa618_y4;
  assign f_s_dadda_pg_rca32_fa621_y3 = f_s_dadda_pg_rca32_fa621_y0 & f_s_dadda_pg_rca32_fa621_f_s_dadda_pg_rca32_fa618_y4;
  assign f_s_dadda_pg_rca32_fa621_y4 = f_s_dadda_pg_rca32_fa621_y1 | f_s_dadda_pg_rca32_fa621_y3;
  assign f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa617_y4 = f_s_dadda_pg_rca32_fa617_y4;
  assign f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa616_y4 = f_s_dadda_pg_rca32_fa616_y4;
  assign f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa615_y4 = f_s_dadda_pg_rca32_fa615_y4;
  assign f_s_dadda_pg_rca32_fa622_y0 = f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa617_y4 ^ f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa616_y4;
  assign f_s_dadda_pg_rca32_fa622_y1 = f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa617_y4 & f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa616_y4;
  assign f_s_dadda_pg_rca32_fa622_y2 = f_s_dadda_pg_rca32_fa622_y0 ^ f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa615_y4;
  assign f_s_dadda_pg_rca32_fa622_y3 = f_s_dadda_pg_rca32_fa622_y0 & f_s_dadda_pg_rca32_fa622_f_s_dadda_pg_rca32_fa615_y4;
  assign f_s_dadda_pg_rca32_fa622_y4 = f_s_dadda_pg_rca32_fa622_y1 | f_s_dadda_pg_rca32_fa622_y3;
  assign f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa614_y4 = f_s_dadda_pg_rca32_fa614_y4;
  assign f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa613_y4 = f_s_dadda_pg_rca32_fa613_y4;
  assign f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa612_y4 = f_s_dadda_pg_rca32_fa612_y4;
  assign f_s_dadda_pg_rca32_fa623_y0 = f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa614_y4 ^ f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa613_y4;
  assign f_s_dadda_pg_rca32_fa623_y1 = f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa614_y4 & f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa613_y4;
  assign f_s_dadda_pg_rca32_fa623_y2 = f_s_dadda_pg_rca32_fa623_y0 ^ f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa612_y4;
  assign f_s_dadda_pg_rca32_fa623_y3 = f_s_dadda_pg_rca32_fa623_y0 & f_s_dadda_pg_rca32_fa623_f_s_dadda_pg_rca32_fa612_y4;
  assign f_s_dadda_pg_rca32_fa623_y4 = f_s_dadda_pg_rca32_fa623_y1 | f_s_dadda_pg_rca32_fa623_y3;
  assign f_s_dadda_pg_rca32_nand_31_17_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_17_b_17 = b_17;
  assign f_s_dadda_pg_rca32_nand_31_17_y0 = ~(f_s_dadda_pg_rca32_nand_31_17_a_31 & f_s_dadda_pg_rca32_nand_31_17_b_17);
  assign f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_fa611_y4 = f_s_dadda_pg_rca32_fa611_y4;
  assign f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_fa610_y4 = f_s_dadda_pg_rca32_fa610_y4;
  assign f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_nand_31_17_y0 = f_s_dadda_pg_rca32_nand_31_17_y0;
  assign f_s_dadda_pg_rca32_fa624_y0 = f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_fa611_y4 ^ f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_fa610_y4;
  assign f_s_dadda_pg_rca32_fa624_y1 = f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_fa611_y4 & f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_fa610_y4;
  assign f_s_dadda_pg_rca32_fa624_y2 = f_s_dadda_pg_rca32_fa624_y0 ^ f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_nand_31_17_y0;
  assign f_s_dadda_pg_rca32_fa624_y3 = f_s_dadda_pg_rca32_fa624_y0 & f_s_dadda_pg_rca32_fa624_f_s_dadda_pg_rca32_nand_31_17_y0;
  assign f_s_dadda_pg_rca32_fa624_y4 = f_s_dadda_pg_rca32_fa624_y1 | f_s_dadda_pg_rca32_fa624_y3;
  assign f_s_dadda_pg_rca32_and_30_18_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_and_30_18_y0 = f_s_dadda_pg_rca32_and_30_18_a_30 & f_s_dadda_pg_rca32_and_30_18_b_18;
  assign f_s_dadda_pg_rca32_and_29_19_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_29_19_y0 = f_s_dadda_pg_rca32_and_29_19_a_29 & f_s_dadda_pg_rca32_and_29_19_b_19;
  assign f_s_dadda_pg_rca32_and_28_20_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_28_20_y0 = f_s_dadda_pg_rca32_and_28_20_a_28 & f_s_dadda_pg_rca32_and_28_20_b_20;
  assign f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_30_18_y0 = f_s_dadda_pg_rca32_and_30_18_y0;
  assign f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_29_19_y0 = f_s_dadda_pg_rca32_and_29_19_y0;
  assign f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_28_20_y0 = f_s_dadda_pg_rca32_and_28_20_y0;
  assign f_s_dadda_pg_rca32_fa625_y0 = f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_30_18_y0 ^ f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_29_19_y0;
  assign f_s_dadda_pg_rca32_fa625_y1 = f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_30_18_y0 & f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_29_19_y0;
  assign f_s_dadda_pg_rca32_fa625_y2 = f_s_dadda_pg_rca32_fa625_y0 ^ f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_28_20_y0;
  assign f_s_dadda_pg_rca32_fa625_y3 = f_s_dadda_pg_rca32_fa625_y0 & f_s_dadda_pg_rca32_fa625_f_s_dadda_pg_rca32_and_28_20_y0;
  assign f_s_dadda_pg_rca32_fa625_y4 = f_s_dadda_pg_rca32_fa625_y1 | f_s_dadda_pg_rca32_fa625_y3;
  assign f_s_dadda_pg_rca32_and_27_21_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_27_21_y0 = f_s_dadda_pg_rca32_and_27_21_a_27 & f_s_dadda_pg_rca32_and_27_21_b_21;
  assign f_s_dadda_pg_rca32_and_26_22_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_26_22_y0 = f_s_dadda_pg_rca32_and_26_22_a_26 & f_s_dadda_pg_rca32_and_26_22_b_22;
  assign f_s_dadda_pg_rca32_and_25_23_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_25_23_y0 = f_s_dadda_pg_rca32_and_25_23_a_25 & f_s_dadda_pg_rca32_and_25_23_b_23;
  assign f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_27_21_y0 = f_s_dadda_pg_rca32_and_27_21_y0;
  assign f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_26_22_y0 = f_s_dadda_pg_rca32_and_26_22_y0;
  assign f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_25_23_y0 = f_s_dadda_pg_rca32_and_25_23_y0;
  assign f_s_dadda_pg_rca32_fa626_y0 = f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_27_21_y0 ^ f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_26_22_y0;
  assign f_s_dadda_pg_rca32_fa626_y1 = f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_27_21_y0 & f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_26_22_y0;
  assign f_s_dadda_pg_rca32_fa626_y2 = f_s_dadda_pg_rca32_fa626_y0 ^ f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_25_23_y0;
  assign f_s_dadda_pg_rca32_fa626_y3 = f_s_dadda_pg_rca32_fa626_y0 & f_s_dadda_pg_rca32_fa626_f_s_dadda_pg_rca32_and_25_23_y0;
  assign f_s_dadda_pg_rca32_fa626_y4 = f_s_dadda_pg_rca32_fa626_y1 | f_s_dadda_pg_rca32_fa626_y3;
  assign f_s_dadda_pg_rca32_and_24_24_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_24_24_y0 = f_s_dadda_pg_rca32_and_24_24_a_24 & f_s_dadda_pg_rca32_and_24_24_b_24;
  assign f_s_dadda_pg_rca32_and_23_25_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_23_25_y0 = f_s_dadda_pg_rca32_and_23_25_a_23 & f_s_dadda_pg_rca32_and_23_25_b_25;
  assign f_s_dadda_pg_rca32_and_22_26_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_22_26_y0 = f_s_dadda_pg_rca32_and_22_26_a_22 & f_s_dadda_pg_rca32_and_22_26_b_26;
  assign f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_24_24_y0 = f_s_dadda_pg_rca32_and_24_24_y0;
  assign f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_23_25_y0 = f_s_dadda_pg_rca32_and_23_25_y0;
  assign f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_22_26_y0 = f_s_dadda_pg_rca32_and_22_26_y0;
  assign f_s_dadda_pg_rca32_fa627_y0 = f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_24_24_y0 ^ f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_23_25_y0;
  assign f_s_dadda_pg_rca32_fa627_y1 = f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_24_24_y0 & f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_23_25_y0;
  assign f_s_dadda_pg_rca32_fa627_y2 = f_s_dadda_pg_rca32_fa627_y0 ^ f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_22_26_y0;
  assign f_s_dadda_pg_rca32_fa627_y3 = f_s_dadda_pg_rca32_fa627_y0 & f_s_dadda_pg_rca32_fa627_f_s_dadda_pg_rca32_and_22_26_y0;
  assign f_s_dadda_pg_rca32_fa627_y4 = f_s_dadda_pg_rca32_fa627_y1 | f_s_dadda_pg_rca32_fa627_y3;
  assign f_s_dadda_pg_rca32_and_21_27_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_21_27_y0 = f_s_dadda_pg_rca32_and_21_27_a_21 & f_s_dadda_pg_rca32_and_21_27_b_27;
  assign f_s_dadda_pg_rca32_and_20_28_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_20_28_y0 = f_s_dadda_pg_rca32_and_20_28_a_20 & f_s_dadda_pg_rca32_and_20_28_b_28;
  assign f_s_dadda_pg_rca32_and_19_29_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_19_29_y0 = f_s_dadda_pg_rca32_and_19_29_a_19 & f_s_dadda_pg_rca32_and_19_29_b_29;
  assign f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_21_27_y0 = f_s_dadda_pg_rca32_and_21_27_y0;
  assign f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_20_28_y0 = f_s_dadda_pg_rca32_and_20_28_y0;
  assign f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_19_29_y0 = f_s_dadda_pg_rca32_and_19_29_y0;
  assign f_s_dadda_pg_rca32_fa628_y0 = f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_21_27_y0 ^ f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_20_28_y0;
  assign f_s_dadda_pg_rca32_fa628_y1 = f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_21_27_y0 & f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_20_28_y0;
  assign f_s_dadda_pg_rca32_fa628_y2 = f_s_dadda_pg_rca32_fa628_y0 ^ f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_19_29_y0;
  assign f_s_dadda_pg_rca32_fa628_y3 = f_s_dadda_pg_rca32_fa628_y0 & f_s_dadda_pg_rca32_fa628_f_s_dadda_pg_rca32_and_19_29_y0;
  assign f_s_dadda_pg_rca32_fa628_y4 = f_s_dadda_pg_rca32_fa628_y1 | f_s_dadda_pg_rca32_fa628_y3;
  assign f_s_dadda_pg_rca32_and_18_30_a_18 = a_18;
  assign f_s_dadda_pg_rca32_and_18_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_18_30_y0 = f_s_dadda_pg_rca32_and_18_30_a_18 & f_s_dadda_pg_rca32_and_18_30_b_30;
  assign f_s_dadda_pg_rca32_nand_17_31_a_17 = a_17;
  assign f_s_dadda_pg_rca32_nand_17_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_17_31_y0 = ~(f_s_dadda_pg_rca32_nand_17_31_a_17 & f_s_dadda_pg_rca32_nand_17_31_b_31);
  assign f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_and_18_30_y0 = f_s_dadda_pg_rca32_and_18_30_y0;
  assign f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_nand_17_31_y0 = f_s_dadda_pg_rca32_nand_17_31_y0;
  assign f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_fa621_y2 = f_s_dadda_pg_rca32_fa621_y2;
  assign f_s_dadda_pg_rca32_fa629_y0 = f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_and_18_30_y0 ^ f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_nand_17_31_y0;
  assign f_s_dadda_pg_rca32_fa629_y1 = f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_and_18_30_y0 & f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_nand_17_31_y0;
  assign f_s_dadda_pg_rca32_fa629_y2 = f_s_dadda_pg_rca32_fa629_y0 ^ f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_fa621_y2;
  assign f_s_dadda_pg_rca32_fa629_y3 = f_s_dadda_pg_rca32_fa629_y0 & f_s_dadda_pg_rca32_fa629_f_s_dadda_pg_rca32_fa621_y2;
  assign f_s_dadda_pg_rca32_fa629_y4 = f_s_dadda_pg_rca32_fa629_y1 | f_s_dadda_pg_rca32_fa629_y3;
  assign f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa622_y2 = f_s_dadda_pg_rca32_fa622_y2;
  assign f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa623_y2 = f_s_dadda_pg_rca32_fa623_y2;
  assign f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa624_y2 = f_s_dadda_pg_rca32_fa624_y2;
  assign f_s_dadda_pg_rca32_fa630_y0 = f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa622_y2 ^ f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa623_y2;
  assign f_s_dadda_pg_rca32_fa630_y1 = f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa622_y2 & f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa623_y2;
  assign f_s_dadda_pg_rca32_fa630_y2 = f_s_dadda_pg_rca32_fa630_y0 ^ f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa624_y2;
  assign f_s_dadda_pg_rca32_fa630_y3 = f_s_dadda_pg_rca32_fa630_y0 & f_s_dadda_pg_rca32_fa630_f_s_dadda_pg_rca32_fa624_y2;
  assign f_s_dadda_pg_rca32_fa630_y4 = f_s_dadda_pg_rca32_fa630_y1 | f_s_dadda_pg_rca32_fa630_y3;
  assign f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa630_y4 = f_s_dadda_pg_rca32_fa630_y4;
  assign f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa629_y4 = f_s_dadda_pg_rca32_fa629_y4;
  assign f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa628_y4 = f_s_dadda_pg_rca32_fa628_y4;
  assign f_s_dadda_pg_rca32_fa631_y0 = f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa630_y4 ^ f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa629_y4;
  assign f_s_dadda_pg_rca32_fa631_y1 = f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa630_y4 & f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa629_y4;
  assign f_s_dadda_pg_rca32_fa631_y2 = f_s_dadda_pg_rca32_fa631_y0 ^ f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa628_y4;
  assign f_s_dadda_pg_rca32_fa631_y3 = f_s_dadda_pg_rca32_fa631_y0 & f_s_dadda_pg_rca32_fa631_f_s_dadda_pg_rca32_fa628_y4;
  assign f_s_dadda_pg_rca32_fa631_y4 = f_s_dadda_pg_rca32_fa631_y1 | f_s_dadda_pg_rca32_fa631_y3;
  assign f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa627_y4 = f_s_dadda_pg_rca32_fa627_y4;
  assign f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa626_y4 = f_s_dadda_pg_rca32_fa626_y4;
  assign f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa625_y4 = f_s_dadda_pg_rca32_fa625_y4;
  assign f_s_dadda_pg_rca32_fa632_y0 = f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa627_y4 ^ f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa626_y4;
  assign f_s_dadda_pg_rca32_fa632_y1 = f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa627_y4 & f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa626_y4;
  assign f_s_dadda_pg_rca32_fa632_y2 = f_s_dadda_pg_rca32_fa632_y0 ^ f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa625_y4;
  assign f_s_dadda_pg_rca32_fa632_y3 = f_s_dadda_pg_rca32_fa632_y0 & f_s_dadda_pg_rca32_fa632_f_s_dadda_pg_rca32_fa625_y4;
  assign f_s_dadda_pg_rca32_fa632_y4 = f_s_dadda_pg_rca32_fa632_y1 | f_s_dadda_pg_rca32_fa632_y3;
  assign f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa624_y4 = f_s_dadda_pg_rca32_fa624_y4;
  assign f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa623_y4 = f_s_dadda_pg_rca32_fa623_y4;
  assign f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa622_y4 = f_s_dadda_pg_rca32_fa622_y4;
  assign f_s_dadda_pg_rca32_fa633_y0 = f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa624_y4 ^ f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa623_y4;
  assign f_s_dadda_pg_rca32_fa633_y1 = f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa624_y4 & f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa623_y4;
  assign f_s_dadda_pg_rca32_fa633_y2 = f_s_dadda_pg_rca32_fa633_y0 ^ f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa622_y4;
  assign f_s_dadda_pg_rca32_fa633_y3 = f_s_dadda_pg_rca32_fa633_y0 & f_s_dadda_pg_rca32_fa633_f_s_dadda_pg_rca32_fa622_y4;
  assign f_s_dadda_pg_rca32_fa633_y4 = f_s_dadda_pg_rca32_fa633_y1 | f_s_dadda_pg_rca32_fa633_y3;
  assign f_s_dadda_pg_rca32_nand_31_18_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_18_b_18 = b_18;
  assign f_s_dadda_pg_rca32_nand_31_18_y0 = ~(f_s_dadda_pg_rca32_nand_31_18_a_31 & f_s_dadda_pg_rca32_nand_31_18_b_18);
  assign f_s_dadda_pg_rca32_and_30_19_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_and_30_19_y0 = f_s_dadda_pg_rca32_and_30_19_a_30 & f_s_dadda_pg_rca32_and_30_19_b_19;
  assign f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_fa621_y4 = f_s_dadda_pg_rca32_fa621_y4;
  assign f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_nand_31_18_y0 = f_s_dadda_pg_rca32_nand_31_18_y0;
  assign f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_and_30_19_y0 = f_s_dadda_pg_rca32_and_30_19_y0;
  assign f_s_dadda_pg_rca32_fa634_y0 = f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_fa621_y4 ^ f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_nand_31_18_y0;
  assign f_s_dadda_pg_rca32_fa634_y1 = f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_fa621_y4 & f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_nand_31_18_y0;
  assign f_s_dadda_pg_rca32_fa634_y2 = f_s_dadda_pg_rca32_fa634_y0 ^ f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_and_30_19_y0;
  assign f_s_dadda_pg_rca32_fa634_y3 = f_s_dadda_pg_rca32_fa634_y0 & f_s_dadda_pg_rca32_fa634_f_s_dadda_pg_rca32_and_30_19_y0;
  assign f_s_dadda_pg_rca32_fa634_y4 = f_s_dadda_pg_rca32_fa634_y1 | f_s_dadda_pg_rca32_fa634_y3;
  assign f_s_dadda_pg_rca32_and_29_20_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_29_20_y0 = f_s_dadda_pg_rca32_and_29_20_a_29 & f_s_dadda_pg_rca32_and_29_20_b_20;
  assign f_s_dadda_pg_rca32_and_28_21_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_28_21_y0 = f_s_dadda_pg_rca32_and_28_21_a_28 & f_s_dadda_pg_rca32_and_28_21_b_21;
  assign f_s_dadda_pg_rca32_and_27_22_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_27_22_y0 = f_s_dadda_pg_rca32_and_27_22_a_27 & f_s_dadda_pg_rca32_and_27_22_b_22;
  assign f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_29_20_y0 = f_s_dadda_pg_rca32_and_29_20_y0;
  assign f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_28_21_y0 = f_s_dadda_pg_rca32_and_28_21_y0;
  assign f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_27_22_y0 = f_s_dadda_pg_rca32_and_27_22_y0;
  assign f_s_dadda_pg_rca32_fa635_y0 = f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_29_20_y0 ^ f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_28_21_y0;
  assign f_s_dadda_pg_rca32_fa635_y1 = f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_29_20_y0 & f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_28_21_y0;
  assign f_s_dadda_pg_rca32_fa635_y2 = f_s_dadda_pg_rca32_fa635_y0 ^ f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_27_22_y0;
  assign f_s_dadda_pg_rca32_fa635_y3 = f_s_dadda_pg_rca32_fa635_y0 & f_s_dadda_pg_rca32_fa635_f_s_dadda_pg_rca32_and_27_22_y0;
  assign f_s_dadda_pg_rca32_fa635_y4 = f_s_dadda_pg_rca32_fa635_y1 | f_s_dadda_pg_rca32_fa635_y3;
  assign f_s_dadda_pg_rca32_and_26_23_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_26_23_y0 = f_s_dadda_pg_rca32_and_26_23_a_26 & f_s_dadda_pg_rca32_and_26_23_b_23;
  assign f_s_dadda_pg_rca32_and_25_24_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_25_24_y0 = f_s_dadda_pg_rca32_and_25_24_a_25 & f_s_dadda_pg_rca32_and_25_24_b_24;
  assign f_s_dadda_pg_rca32_and_24_25_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_24_25_y0 = f_s_dadda_pg_rca32_and_24_25_a_24 & f_s_dadda_pg_rca32_and_24_25_b_25;
  assign f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_26_23_y0 = f_s_dadda_pg_rca32_and_26_23_y0;
  assign f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_25_24_y0 = f_s_dadda_pg_rca32_and_25_24_y0;
  assign f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_24_25_y0 = f_s_dadda_pg_rca32_and_24_25_y0;
  assign f_s_dadda_pg_rca32_fa636_y0 = f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_26_23_y0 ^ f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_25_24_y0;
  assign f_s_dadda_pg_rca32_fa636_y1 = f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_26_23_y0 & f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_25_24_y0;
  assign f_s_dadda_pg_rca32_fa636_y2 = f_s_dadda_pg_rca32_fa636_y0 ^ f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_24_25_y0;
  assign f_s_dadda_pg_rca32_fa636_y3 = f_s_dadda_pg_rca32_fa636_y0 & f_s_dadda_pg_rca32_fa636_f_s_dadda_pg_rca32_and_24_25_y0;
  assign f_s_dadda_pg_rca32_fa636_y4 = f_s_dadda_pg_rca32_fa636_y1 | f_s_dadda_pg_rca32_fa636_y3;
  assign f_s_dadda_pg_rca32_and_23_26_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_23_26_y0 = f_s_dadda_pg_rca32_and_23_26_a_23 & f_s_dadda_pg_rca32_and_23_26_b_26;
  assign f_s_dadda_pg_rca32_and_22_27_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_22_27_y0 = f_s_dadda_pg_rca32_and_22_27_a_22 & f_s_dadda_pg_rca32_and_22_27_b_27;
  assign f_s_dadda_pg_rca32_and_21_28_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_21_28_y0 = f_s_dadda_pg_rca32_and_21_28_a_21 & f_s_dadda_pg_rca32_and_21_28_b_28;
  assign f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_23_26_y0 = f_s_dadda_pg_rca32_and_23_26_y0;
  assign f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_22_27_y0 = f_s_dadda_pg_rca32_and_22_27_y0;
  assign f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_21_28_y0 = f_s_dadda_pg_rca32_and_21_28_y0;
  assign f_s_dadda_pg_rca32_fa637_y0 = f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_23_26_y0 ^ f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_22_27_y0;
  assign f_s_dadda_pg_rca32_fa637_y1 = f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_23_26_y0 & f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_22_27_y0;
  assign f_s_dadda_pg_rca32_fa637_y2 = f_s_dadda_pg_rca32_fa637_y0 ^ f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_21_28_y0;
  assign f_s_dadda_pg_rca32_fa637_y3 = f_s_dadda_pg_rca32_fa637_y0 & f_s_dadda_pg_rca32_fa637_f_s_dadda_pg_rca32_and_21_28_y0;
  assign f_s_dadda_pg_rca32_fa637_y4 = f_s_dadda_pg_rca32_fa637_y1 | f_s_dadda_pg_rca32_fa637_y3;
  assign f_s_dadda_pg_rca32_and_20_29_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_20_29_y0 = f_s_dadda_pg_rca32_and_20_29_a_20 & f_s_dadda_pg_rca32_and_20_29_b_29;
  assign f_s_dadda_pg_rca32_and_19_30_a_19 = a_19;
  assign f_s_dadda_pg_rca32_and_19_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_19_30_y0 = f_s_dadda_pg_rca32_and_19_30_a_19 & f_s_dadda_pg_rca32_and_19_30_b_30;
  assign f_s_dadda_pg_rca32_nand_18_31_a_18 = a_18;
  assign f_s_dadda_pg_rca32_nand_18_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_18_31_y0 = ~(f_s_dadda_pg_rca32_nand_18_31_a_18 & f_s_dadda_pg_rca32_nand_18_31_b_31);
  assign f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_and_20_29_y0 = f_s_dadda_pg_rca32_and_20_29_y0;
  assign f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_and_19_30_y0 = f_s_dadda_pg_rca32_and_19_30_y0;
  assign f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_nand_18_31_y0 = f_s_dadda_pg_rca32_nand_18_31_y0;
  assign f_s_dadda_pg_rca32_fa638_y0 = f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_and_20_29_y0 ^ f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_and_19_30_y0;
  assign f_s_dadda_pg_rca32_fa638_y1 = f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_and_20_29_y0 & f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_and_19_30_y0;
  assign f_s_dadda_pg_rca32_fa638_y2 = f_s_dadda_pg_rca32_fa638_y0 ^ f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_nand_18_31_y0;
  assign f_s_dadda_pg_rca32_fa638_y3 = f_s_dadda_pg_rca32_fa638_y0 & f_s_dadda_pg_rca32_fa638_f_s_dadda_pg_rca32_nand_18_31_y0;
  assign f_s_dadda_pg_rca32_fa638_y4 = f_s_dadda_pg_rca32_fa638_y1 | f_s_dadda_pg_rca32_fa638_y3;
  assign f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa631_y2 = f_s_dadda_pg_rca32_fa631_y2;
  assign f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa632_y2 = f_s_dadda_pg_rca32_fa632_y2;
  assign f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa633_y2 = f_s_dadda_pg_rca32_fa633_y2;
  assign f_s_dadda_pg_rca32_fa639_y0 = f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa631_y2 ^ f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa632_y2;
  assign f_s_dadda_pg_rca32_fa639_y1 = f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa631_y2 & f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa632_y2;
  assign f_s_dadda_pg_rca32_fa639_y2 = f_s_dadda_pg_rca32_fa639_y0 ^ f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa633_y2;
  assign f_s_dadda_pg_rca32_fa639_y3 = f_s_dadda_pg_rca32_fa639_y0 & f_s_dadda_pg_rca32_fa639_f_s_dadda_pg_rca32_fa633_y2;
  assign f_s_dadda_pg_rca32_fa639_y4 = f_s_dadda_pg_rca32_fa639_y1 | f_s_dadda_pg_rca32_fa639_y3;
  assign f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa639_y4 = f_s_dadda_pg_rca32_fa639_y4;
  assign f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa638_y4 = f_s_dadda_pg_rca32_fa638_y4;
  assign f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa637_y4 = f_s_dadda_pg_rca32_fa637_y4;
  assign f_s_dadda_pg_rca32_fa640_y0 = f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa639_y4 ^ f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa638_y4;
  assign f_s_dadda_pg_rca32_fa640_y1 = f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa639_y4 & f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa638_y4;
  assign f_s_dadda_pg_rca32_fa640_y2 = f_s_dadda_pg_rca32_fa640_y0 ^ f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa637_y4;
  assign f_s_dadda_pg_rca32_fa640_y3 = f_s_dadda_pg_rca32_fa640_y0 & f_s_dadda_pg_rca32_fa640_f_s_dadda_pg_rca32_fa637_y4;
  assign f_s_dadda_pg_rca32_fa640_y4 = f_s_dadda_pg_rca32_fa640_y1 | f_s_dadda_pg_rca32_fa640_y3;
  assign f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa636_y4 = f_s_dadda_pg_rca32_fa636_y4;
  assign f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa635_y4 = f_s_dadda_pg_rca32_fa635_y4;
  assign f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa634_y4 = f_s_dadda_pg_rca32_fa634_y4;
  assign f_s_dadda_pg_rca32_fa641_y0 = f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa636_y4 ^ f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa635_y4;
  assign f_s_dadda_pg_rca32_fa641_y1 = f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa636_y4 & f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa635_y4;
  assign f_s_dadda_pg_rca32_fa641_y2 = f_s_dadda_pg_rca32_fa641_y0 ^ f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa634_y4;
  assign f_s_dadda_pg_rca32_fa641_y3 = f_s_dadda_pg_rca32_fa641_y0 & f_s_dadda_pg_rca32_fa641_f_s_dadda_pg_rca32_fa634_y4;
  assign f_s_dadda_pg_rca32_fa641_y4 = f_s_dadda_pg_rca32_fa641_y1 | f_s_dadda_pg_rca32_fa641_y3;
  assign f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa633_y4 = f_s_dadda_pg_rca32_fa633_y4;
  assign f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa632_y4 = f_s_dadda_pg_rca32_fa632_y4;
  assign f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa631_y4 = f_s_dadda_pg_rca32_fa631_y4;
  assign f_s_dadda_pg_rca32_fa642_y0 = f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa633_y4 ^ f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa632_y4;
  assign f_s_dadda_pg_rca32_fa642_y1 = f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa633_y4 & f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa632_y4;
  assign f_s_dadda_pg_rca32_fa642_y2 = f_s_dadda_pg_rca32_fa642_y0 ^ f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa631_y4;
  assign f_s_dadda_pg_rca32_fa642_y3 = f_s_dadda_pg_rca32_fa642_y0 & f_s_dadda_pg_rca32_fa642_f_s_dadda_pg_rca32_fa631_y4;
  assign f_s_dadda_pg_rca32_fa642_y4 = f_s_dadda_pg_rca32_fa642_y1 | f_s_dadda_pg_rca32_fa642_y3;
  assign f_s_dadda_pg_rca32_nand_31_19_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_19_b_19 = b_19;
  assign f_s_dadda_pg_rca32_nand_31_19_y0 = ~(f_s_dadda_pg_rca32_nand_31_19_a_31 & f_s_dadda_pg_rca32_nand_31_19_b_19);
  assign f_s_dadda_pg_rca32_and_30_20_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_and_30_20_y0 = f_s_dadda_pg_rca32_and_30_20_a_30 & f_s_dadda_pg_rca32_and_30_20_b_20;
  assign f_s_dadda_pg_rca32_and_29_21_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_29_21_y0 = f_s_dadda_pg_rca32_and_29_21_a_29 & f_s_dadda_pg_rca32_and_29_21_b_21;
  assign f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_nand_31_19_y0 = f_s_dadda_pg_rca32_nand_31_19_y0;
  assign f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_and_30_20_y0 = f_s_dadda_pg_rca32_and_30_20_y0;
  assign f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_and_29_21_y0 = f_s_dadda_pg_rca32_and_29_21_y0;
  assign f_s_dadda_pg_rca32_fa643_y0 = f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_nand_31_19_y0 ^ f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_and_30_20_y0;
  assign f_s_dadda_pg_rca32_fa643_y1 = f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_nand_31_19_y0 & f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_and_30_20_y0;
  assign f_s_dadda_pg_rca32_fa643_y2 = f_s_dadda_pg_rca32_fa643_y0 ^ f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_and_29_21_y0;
  assign f_s_dadda_pg_rca32_fa643_y3 = f_s_dadda_pg_rca32_fa643_y0 & f_s_dadda_pg_rca32_fa643_f_s_dadda_pg_rca32_and_29_21_y0;
  assign f_s_dadda_pg_rca32_fa643_y4 = f_s_dadda_pg_rca32_fa643_y1 | f_s_dadda_pg_rca32_fa643_y3;
  assign f_s_dadda_pg_rca32_and_28_22_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_28_22_y0 = f_s_dadda_pg_rca32_and_28_22_a_28 & f_s_dadda_pg_rca32_and_28_22_b_22;
  assign f_s_dadda_pg_rca32_and_27_23_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_27_23_y0 = f_s_dadda_pg_rca32_and_27_23_a_27 & f_s_dadda_pg_rca32_and_27_23_b_23;
  assign f_s_dadda_pg_rca32_and_26_24_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_26_24_y0 = f_s_dadda_pg_rca32_and_26_24_a_26 & f_s_dadda_pg_rca32_and_26_24_b_24;
  assign f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_28_22_y0 = f_s_dadda_pg_rca32_and_28_22_y0;
  assign f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_27_23_y0 = f_s_dadda_pg_rca32_and_27_23_y0;
  assign f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_26_24_y0 = f_s_dadda_pg_rca32_and_26_24_y0;
  assign f_s_dadda_pg_rca32_fa644_y0 = f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_28_22_y0 ^ f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_27_23_y0;
  assign f_s_dadda_pg_rca32_fa644_y1 = f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_28_22_y0 & f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_27_23_y0;
  assign f_s_dadda_pg_rca32_fa644_y2 = f_s_dadda_pg_rca32_fa644_y0 ^ f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_26_24_y0;
  assign f_s_dadda_pg_rca32_fa644_y3 = f_s_dadda_pg_rca32_fa644_y0 & f_s_dadda_pg_rca32_fa644_f_s_dadda_pg_rca32_and_26_24_y0;
  assign f_s_dadda_pg_rca32_fa644_y4 = f_s_dadda_pg_rca32_fa644_y1 | f_s_dadda_pg_rca32_fa644_y3;
  assign f_s_dadda_pg_rca32_and_25_25_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_25_25_y0 = f_s_dadda_pg_rca32_and_25_25_a_25 & f_s_dadda_pg_rca32_and_25_25_b_25;
  assign f_s_dadda_pg_rca32_and_24_26_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_24_26_y0 = f_s_dadda_pg_rca32_and_24_26_a_24 & f_s_dadda_pg_rca32_and_24_26_b_26;
  assign f_s_dadda_pg_rca32_and_23_27_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_23_27_y0 = f_s_dadda_pg_rca32_and_23_27_a_23 & f_s_dadda_pg_rca32_and_23_27_b_27;
  assign f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_25_25_y0 = f_s_dadda_pg_rca32_and_25_25_y0;
  assign f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_24_26_y0 = f_s_dadda_pg_rca32_and_24_26_y0;
  assign f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_23_27_y0 = f_s_dadda_pg_rca32_and_23_27_y0;
  assign f_s_dadda_pg_rca32_fa645_y0 = f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_25_25_y0 ^ f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_24_26_y0;
  assign f_s_dadda_pg_rca32_fa645_y1 = f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_25_25_y0 & f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_24_26_y0;
  assign f_s_dadda_pg_rca32_fa645_y2 = f_s_dadda_pg_rca32_fa645_y0 ^ f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_23_27_y0;
  assign f_s_dadda_pg_rca32_fa645_y3 = f_s_dadda_pg_rca32_fa645_y0 & f_s_dadda_pg_rca32_fa645_f_s_dadda_pg_rca32_and_23_27_y0;
  assign f_s_dadda_pg_rca32_fa645_y4 = f_s_dadda_pg_rca32_fa645_y1 | f_s_dadda_pg_rca32_fa645_y3;
  assign f_s_dadda_pg_rca32_and_22_28_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_22_28_y0 = f_s_dadda_pg_rca32_and_22_28_a_22 & f_s_dadda_pg_rca32_and_22_28_b_28;
  assign f_s_dadda_pg_rca32_and_21_29_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_21_29_y0 = f_s_dadda_pg_rca32_and_21_29_a_21 & f_s_dadda_pg_rca32_and_21_29_b_29;
  assign f_s_dadda_pg_rca32_and_20_30_a_20 = a_20;
  assign f_s_dadda_pg_rca32_and_20_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_20_30_y0 = f_s_dadda_pg_rca32_and_20_30_a_20 & f_s_dadda_pg_rca32_and_20_30_b_30;
  assign f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_22_28_y0 = f_s_dadda_pg_rca32_and_22_28_y0;
  assign f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_21_29_y0 = f_s_dadda_pg_rca32_and_21_29_y0;
  assign f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_20_30_y0 = f_s_dadda_pg_rca32_and_20_30_y0;
  assign f_s_dadda_pg_rca32_fa646_y0 = f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_22_28_y0 ^ f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_21_29_y0;
  assign f_s_dadda_pg_rca32_fa646_y1 = f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_22_28_y0 & f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_21_29_y0;
  assign f_s_dadda_pg_rca32_fa646_y2 = f_s_dadda_pg_rca32_fa646_y0 ^ f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_20_30_y0;
  assign f_s_dadda_pg_rca32_fa646_y3 = f_s_dadda_pg_rca32_fa646_y0 & f_s_dadda_pg_rca32_fa646_f_s_dadda_pg_rca32_and_20_30_y0;
  assign f_s_dadda_pg_rca32_fa646_y4 = f_s_dadda_pg_rca32_fa646_y1 | f_s_dadda_pg_rca32_fa646_y3;
  assign f_s_dadda_pg_rca32_nand_19_31_a_19 = a_19;
  assign f_s_dadda_pg_rca32_nand_19_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_19_31_y0 = ~(f_s_dadda_pg_rca32_nand_19_31_a_19 & f_s_dadda_pg_rca32_nand_19_31_b_31);
  assign f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_nand_19_31_y0 = f_s_dadda_pg_rca32_nand_19_31_y0;
  assign f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_fa640_y2 = f_s_dadda_pg_rca32_fa640_y2;
  assign f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_fa641_y2 = f_s_dadda_pg_rca32_fa641_y2;
  assign f_s_dadda_pg_rca32_fa647_y0 = f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_nand_19_31_y0 ^ f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_fa640_y2;
  assign f_s_dadda_pg_rca32_fa647_y1 = f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_nand_19_31_y0 & f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_fa640_y2;
  assign f_s_dadda_pg_rca32_fa647_y2 = f_s_dadda_pg_rca32_fa647_y0 ^ f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_fa641_y2;
  assign f_s_dadda_pg_rca32_fa647_y3 = f_s_dadda_pg_rca32_fa647_y0 & f_s_dadda_pg_rca32_fa647_f_s_dadda_pg_rca32_fa641_y2;
  assign f_s_dadda_pg_rca32_fa647_y4 = f_s_dadda_pg_rca32_fa647_y1 | f_s_dadda_pg_rca32_fa647_y3;
  assign f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa647_y4 = f_s_dadda_pg_rca32_fa647_y4;
  assign f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa646_y4 = f_s_dadda_pg_rca32_fa646_y4;
  assign f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa645_y4 = f_s_dadda_pg_rca32_fa645_y4;
  assign f_s_dadda_pg_rca32_fa648_y0 = f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa647_y4 ^ f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa646_y4;
  assign f_s_dadda_pg_rca32_fa648_y1 = f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa647_y4 & f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa646_y4;
  assign f_s_dadda_pg_rca32_fa648_y2 = f_s_dadda_pg_rca32_fa648_y0 ^ f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa645_y4;
  assign f_s_dadda_pg_rca32_fa648_y3 = f_s_dadda_pg_rca32_fa648_y0 & f_s_dadda_pg_rca32_fa648_f_s_dadda_pg_rca32_fa645_y4;
  assign f_s_dadda_pg_rca32_fa648_y4 = f_s_dadda_pg_rca32_fa648_y1 | f_s_dadda_pg_rca32_fa648_y3;
  assign f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa644_y4 = f_s_dadda_pg_rca32_fa644_y4;
  assign f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa643_y4 = f_s_dadda_pg_rca32_fa643_y4;
  assign f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa642_y4 = f_s_dadda_pg_rca32_fa642_y4;
  assign f_s_dadda_pg_rca32_fa649_y0 = f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa644_y4 ^ f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa643_y4;
  assign f_s_dadda_pg_rca32_fa649_y1 = f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa644_y4 & f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa643_y4;
  assign f_s_dadda_pg_rca32_fa649_y2 = f_s_dadda_pg_rca32_fa649_y0 ^ f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa642_y4;
  assign f_s_dadda_pg_rca32_fa649_y3 = f_s_dadda_pg_rca32_fa649_y0 & f_s_dadda_pg_rca32_fa649_f_s_dadda_pg_rca32_fa642_y4;
  assign f_s_dadda_pg_rca32_fa649_y4 = f_s_dadda_pg_rca32_fa649_y1 | f_s_dadda_pg_rca32_fa649_y3;
  assign f_s_dadda_pg_rca32_nand_31_20_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_20_b_20 = b_20;
  assign f_s_dadda_pg_rca32_nand_31_20_y0 = ~(f_s_dadda_pg_rca32_nand_31_20_a_31 & f_s_dadda_pg_rca32_nand_31_20_b_20);
  assign f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_fa641_y4 = f_s_dadda_pg_rca32_fa641_y4;
  assign f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_fa640_y4 = f_s_dadda_pg_rca32_fa640_y4;
  assign f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_nand_31_20_y0 = f_s_dadda_pg_rca32_nand_31_20_y0;
  assign f_s_dadda_pg_rca32_fa650_y0 = f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_fa641_y4 ^ f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_fa640_y4;
  assign f_s_dadda_pg_rca32_fa650_y1 = f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_fa641_y4 & f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_fa640_y4;
  assign f_s_dadda_pg_rca32_fa650_y2 = f_s_dadda_pg_rca32_fa650_y0 ^ f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_nand_31_20_y0;
  assign f_s_dadda_pg_rca32_fa650_y3 = f_s_dadda_pg_rca32_fa650_y0 & f_s_dadda_pg_rca32_fa650_f_s_dadda_pg_rca32_nand_31_20_y0;
  assign f_s_dadda_pg_rca32_fa650_y4 = f_s_dadda_pg_rca32_fa650_y1 | f_s_dadda_pg_rca32_fa650_y3;
  assign f_s_dadda_pg_rca32_and_30_21_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_and_30_21_y0 = f_s_dadda_pg_rca32_and_30_21_a_30 & f_s_dadda_pg_rca32_and_30_21_b_21;
  assign f_s_dadda_pg_rca32_and_29_22_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_29_22_y0 = f_s_dadda_pg_rca32_and_29_22_a_29 & f_s_dadda_pg_rca32_and_29_22_b_22;
  assign f_s_dadda_pg_rca32_and_28_23_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_28_23_y0 = f_s_dadda_pg_rca32_and_28_23_a_28 & f_s_dadda_pg_rca32_and_28_23_b_23;
  assign f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_30_21_y0 = f_s_dadda_pg_rca32_and_30_21_y0;
  assign f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_29_22_y0 = f_s_dadda_pg_rca32_and_29_22_y0;
  assign f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_28_23_y0 = f_s_dadda_pg_rca32_and_28_23_y0;
  assign f_s_dadda_pg_rca32_fa651_y0 = f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_30_21_y0 ^ f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_29_22_y0;
  assign f_s_dadda_pg_rca32_fa651_y1 = f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_30_21_y0 & f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_29_22_y0;
  assign f_s_dadda_pg_rca32_fa651_y2 = f_s_dadda_pg_rca32_fa651_y0 ^ f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_28_23_y0;
  assign f_s_dadda_pg_rca32_fa651_y3 = f_s_dadda_pg_rca32_fa651_y0 & f_s_dadda_pg_rca32_fa651_f_s_dadda_pg_rca32_and_28_23_y0;
  assign f_s_dadda_pg_rca32_fa651_y4 = f_s_dadda_pg_rca32_fa651_y1 | f_s_dadda_pg_rca32_fa651_y3;
  assign f_s_dadda_pg_rca32_and_27_24_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_27_24_y0 = f_s_dadda_pg_rca32_and_27_24_a_27 & f_s_dadda_pg_rca32_and_27_24_b_24;
  assign f_s_dadda_pg_rca32_and_26_25_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_26_25_y0 = f_s_dadda_pg_rca32_and_26_25_a_26 & f_s_dadda_pg_rca32_and_26_25_b_25;
  assign f_s_dadda_pg_rca32_and_25_26_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_25_26_y0 = f_s_dadda_pg_rca32_and_25_26_a_25 & f_s_dadda_pg_rca32_and_25_26_b_26;
  assign f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_27_24_y0 = f_s_dadda_pg_rca32_and_27_24_y0;
  assign f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_26_25_y0 = f_s_dadda_pg_rca32_and_26_25_y0;
  assign f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_25_26_y0 = f_s_dadda_pg_rca32_and_25_26_y0;
  assign f_s_dadda_pg_rca32_fa652_y0 = f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_27_24_y0 ^ f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_26_25_y0;
  assign f_s_dadda_pg_rca32_fa652_y1 = f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_27_24_y0 & f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_26_25_y0;
  assign f_s_dadda_pg_rca32_fa652_y2 = f_s_dadda_pg_rca32_fa652_y0 ^ f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_25_26_y0;
  assign f_s_dadda_pg_rca32_fa652_y3 = f_s_dadda_pg_rca32_fa652_y0 & f_s_dadda_pg_rca32_fa652_f_s_dadda_pg_rca32_and_25_26_y0;
  assign f_s_dadda_pg_rca32_fa652_y4 = f_s_dadda_pg_rca32_fa652_y1 | f_s_dadda_pg_rca32_fa652_y3;
  assign f_s_dadda_pg_rca32_and_24_27_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_24_27_y0 = f_s_dadda_pg_rca32_and_24_27_a_24 & f_s_dadda_pg_rca32_and_24_27_b_27;
  assign f_s_dadda_pg_rca32_and_23_28_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_23_28_y0 = f_s_dadda_pg_rca32_and_23_28_a_23 & f_s_dadda_pg_rca32_and_23_28_b_28;
  assign f_s_dadda_pg_rca32_and_22_29_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_22_29_y0 = f_s_dadda_pg_rca32_and_22_29_a_22 & f_s_dadda_pg_rca32_and_22_29_b_29;
  assign f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_24_27_y0 = f_s_dadda_pg_rca32_and_24_27_y0;
  assign f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_23_28_y0 = f_s_dadda_pg_rca32_and_23_28_y0;
  assign f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_22_29_y0 = f_s_dadda_pg_rca32_and_22_29_y0;
  assign f_s_dadda_pg_rca32_fa653_y0 = f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_24_27_y0 ^ f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_23_28_y0;
  assign f_s_dadda_pg_rca32_fa653_y1 = f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_24_27_y0 & f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_23_28_y0;
  assign f_s_dadda_pg_rca32_fa653_y2 = f_s_dadda_pg_rca32_fa653_y0 ^ f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_22_29_y0;
  assign f_s_dadda_pg_rca32_fa653_y3 = f_s_dadda_pg_rca32_fa653_y0 & f_s_dadda_pg_rca32_fa653_f_s_dadda_pg_rca32_and_22_29_y0;
  assign f_s_dadda_pg_rca32_fa653_y4 = f_s_dadda_pg_rca32_fa653_y1 | f_s_dadda_pg_rca32_fa653_y3;
  assign f_s_dadda_pg_rca32_and_21_30_a_21 = a_21;
  assign f_s_dadda_pg_rca32_and_21_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_21_30_y0 = f_s_dadda_pg_rca32_and_21_30_a_21 & f_s_dadda_pg_rca32_and_21_30_b_30;
  assign f_s_dadda_pg_rca32_nand_20_31_a_20 = a_20;
  assign f_s_dadda_pg_rca32_nand_20_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_20_31_y0 = ~(f_s_dadda_pg_rca32_nand_20_31_a_20 & f_s_dadda_pg_rca32_nand_20_31_b_31);
  assign f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_and_21_30_y0 = f_s_dadda_pg_rca32_and_21_30_y0;
  assign f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_nand_20_31_y0 = f_s_dadda_pg_rca32_nand_20_31_y0;
  assign f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_fa648_y2 = f_s_dadda_pg_rca32_fa648_y2;
  assign f_s_dadda_pg_rca32_fa654_y0 = f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_and_21_30_y0 ^ f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_nand_20_31_y0;
  assign f_s_dadda_pg_rca32_fa654_y1 = f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_and_21_30_y0 & f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_nand_20_31_y0;
  assign f_s_dadda_pg_rca32_fa654_y2 = f_s_dadda_pg_rca32_fa654_y0 ^ f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_fa648_y2;
  assign f_s_dadda_pg_rca32_fa654_y3 = f_s_dadda_pg_rca32_fa654_y0 & f_s_dadda_pg_rca32_fa654_f_s_dadda_pg_rca32_fa648_y2;
  assign f_s_dadda_pg_rca32_fa654_y4 = f_s_dadda_pg_rca32_fa654_y1 | f_s_dadda_pg_rca32_fa654_y3;
  assign f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa654_y4 = f_s_dadda_pg_rca32_fa654_y4;
  assign f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa653_y4 = f_s_dadda_pg_rca32_fa653_y4;
  assign f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa652_y4 = f_s_dadda_pg_rca32_fa652_y4;
  assign f_s_dadda_pg_rca32_fa655_y0 = f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa654_y4 ^ f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa653_y4;
  assign f_s_dadda_pg_rca32_fa655_y1 = f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa654_y4 & f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa653_y4;
  assign f_s_dadda_pg_rca32_fa655_y2 = f_s_dadda_pg_rca32_fa655_y0 ^ f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa652_y4;
  assign f_s_dadda_pg_rca32_fa655_y3 = f_s_dadda_pg_rca32_fa655_y0 & f_s_dadda_pg_rca32_fa655_f_s_dadda_pg_rca32_fa652_y4;
  assign f_s_dadda_pg_rca32_fa655_y4 = f_s_dadda_pg_rca32_fa655_y1 | f_s_dadda_pg_rca32_fa655_y3;
  assign f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa651_y4 = f_s_dadda_pg_rca32_fa651_y4;
  assign f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa650_y4 = f_s_dadda_pg_rca32_fa650_y4;
  assign f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa649_y4 = f_s_dadda_pg_rca32_fa649_y4;
  assign f_s_dadda_pg_rca32_fa656_y0 = f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa651_y4 ^ f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa650_y4;
  assign f_s_dadda_pg_rca32_fa656_y1 = f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa651_y4 & f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa650_y4;
  assign f_s_dadda_pg_rca32_fa656_y2 = f_s_dadda_pg_rca32_fa656_y0 ^ f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa649_y4;
  assign f_s_dadda_pg_rca32_fa656_y3 = f_s_dadda_pg_rca32_fa656_y0 & f_s_dadda_pg_rca32_fa656_f_s_dadda_pg_rca32_fa649_y4;
  assign f_s_dadda_pg_rca32_fa656_y4 = f_s_dadda_pg_rca32_fa656_y1 | f_s_dadda_pg_rca32_fa656_y3;
  assign f_s_dadda_pg_rca32_nand_31_21_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_21_b_21 = b_21;
  assign f_s_dadda_pg_rca32_nand_31_21_y0 = ~(f_s_dadda_pg_rca32_nand_31_21_a_31 & f_s_dadda_pg_rca32_nand_31_21_b_21);
  assign f_s_dadda_pg_rca32_and_30_22_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_and_30_22_y0 = f_s_dadda_pg_rca32_and_30_22_a_30 & f_s_dadda_pg_rca32_and_30_22_b_22;
  assign f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_fa648_y4 = f_s_dadda_pg_rca32_fa648_y4;
  assign f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_nand_31_21_y0 = f_s_dadda_pg_rca32_nand_31_21_y0;
  assign f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_and_30_22_y0 = f_s_dadda_pg_rca32_and_30_22_y0;
  assign f_s_dadda_pg_rca32_fa657_y0 = f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_fa648_y4 ^ f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_nand_31_21_y0;
  assign f_s_dadda_pg_rca32_fa657_y1 = f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_fa648_y4 & f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_nand_31_21_y0;
  assign f_s_dadda_pg_rca32_fa657_y2 = f_s_dadda_pg_rca32_fa657_y0 ^ f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_and_30_22_y0;
  assign f_s_dadda_pg_rca32_fa657_y3 = f_s_dadda_pg_rca32_fa657_y0 & f_s_dadda_pg_rca32_fa657_f_s_dadda_pg_rca32_and_30_22_y0;
  assign f_s_dadda_pg_rca32_fa657_y4 = f_s_dadda_pg_rca32_fa657_y1 | f_s_dadda_pg_rca32_fa657_y3;
  assign f_s_dadda_pg_rca32_and_29_23_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_29_23_y0 = f_s_dadda_pg_rca32_and_29_23_a_29 & f_s_dadda_pg_rca32_and_29_23_b_23;
  assign f_s_dadda_pg_rca32_and_28_24_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_28_24_y0 = f_s_dadda_pg_rca32_and_28_24_a_28 & f_s_dadda_pg_rca32_and_28_24_b_24;
  assign f_s_dadda_pg_rca32_and_27_25_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_27_25_y0 = f_s_dadda_pg_rca32_and_27_25_a_27 & f_s_dadda_pg_rca32_and_27_25_b_25;
  assign f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_29_23_y0 = f_s_dadda_pg_rca32_and_29_23_y0;
  assign f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_28_24_y0 = f_s_dadda_pg_rca32_and_28_24_y0;
  assign f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_27_25_y0 = f_s_dadda_pg_rca32_and_27_25_y0;
  assign f_s_dadda_pg_rca32_fa658_y0 = f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_29_23_y0 ^ f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_28_24_y0;
  assign f_s_dadda_pg_rca32_fa658_y1 = f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_29_23_y0 & f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_28_24_y0;
  assign f_s_dadda_pg_rca32_fa658_y2 = f_s_dadda_pg_rca32_fa658_y0 ^ f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_27_25_y0;
  assign f_s_dadda_pg_rca32_fa658_y3 = f_s_dadda_pg_rca32_fa658_y0 & f_s_dadda_pg_rca32_fa658_f_s_dadda_pg_rca32_and_27_25_y0;
  assign f_s_dadda_pg_rca32_fa658_y4 = f_s_dadda_pg_rca32_fa658_y1 | f_s_dadda_pg_rca32_fa658_y3;
  assign f_s_dadda_pg_rca32_and_26_26_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_26_26_y0 = f_s_dadda_pg_rca32_and_26_26_a_26 & f_s_dadda_pg_rca32_and_26_26_b_26;
  assign f_s_dadda_pg_rca32_and_25_27_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_25_27_y0 = f_s_dadda_pg_rca32_and_25_27_a_25 & f_s_dadda_pg_rca32_and_25_27_b_27;
  assign f_s_dadda_pg_rca32_and_24_28_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_24_28_y0 = f_s_dadda_pg_rca32_and_24_28_a_24 & f_s_dadda_pg_rca32_and_24_28_b_28;
  assign f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_26_26_y0 = f_s_dadda_pg_rca32_and_26_26_y0;
  assign f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_25_27_y0 = f_s_dadda_pg_rca32_and_25_27_y0;
  assign f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_24_28_y0 = f_s_dadda_pg_rca32_and_24_28_y0;
  assign f_s_dadda_pg_rca32_fa659_y0 = f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_26_26_y0 ^ f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_25_27_y0;
  assign f_s_dadda_pg_rca32_fa659_y1 = f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_26_26_y0 & f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_25_27_y0;
  assign f_s_dadda_pg_rca32_fa659_y2 = f_s_dadda_pg_rca32_fa659_y0 ^ f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_24_28_y0;
  assign f_s_dadda_pg_rca32_fa659_y3 = f_s_dadda_pg_rca32_fa659_y0 & f_s_dadda_pg_rca32_fa659_f_s_dadda_pg_rca32_and_24_28_y0;
  assign f_s_dadda_pg_rca32_fa659_y4 = f_s_dadda_pg_rca32_fa659_y1 | f_s_dadda_pg_rca32_fa659_y3;
  assign f_s_dadda_pg_rca32_and_23_29_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_23_29_y0 = f_s_dadda_pg_rca32_and_23_29_a_23 & f_s_dadda_pg_rca32_and_23_29_b_29;
  assign f_s_dadda_pg_rca32_and_22_30_a_22 = a_22;
  assign f_s_dadda_pg_rca32_and_22_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_22_30_y0 = f_s_dadda_pg_rca32_and_22_30_a_22 & f_s_dadda_pg_rca32_and_22_30_b_30;
  assign f_s_dadda_pg_rca32_nand_21_31_a_21 = a_21;
  assign f_s_dadda_pg_rca32_nand_21_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_21_31_y0 = ~(f_s_dadda_pg_rca32_nand_21_31_a_21 & f_s_dadda_pg_rca32_nand_21_31_b_31);
  assign f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_and_23_29_y0 = f_s_dadda_pg_rca32_and_23_29_y0;
  assign f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_and_22_30_y0 = f_s_dadda_pg_rca32_and_22_30_y0;
  assign f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_nand_21_31_y0 = f_s_dadda_pg_rca32_nand_21_31_y0;
  assign f_s_dadda_pg_rca32_fa660_y0 = f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_and_23_29_y0 ^ f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_and_22_30_y0;
  assign f_s_dadda_pg_rca32_fa660_y1 = f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_and_23_29_y0 & f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_and_22_30_y0;
  assign f_s_dadda_pg_rca32_fa660_y2 = f_s_dadda_pg_rca32_fa660_y0 ^ f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_nand_21_31_y0;
  assign f_s_dadda_pg_rca32_fa660_y3 = f_s_dadda_pg_rca32_fa660_y0 & f_s_dadda_pg_rca32_fa660_f_s_dadda_pg_rca32_nand_21_31_y0;
  assign f_s_dadda_pg_rca32_fa660_y4 = f_s_dadda_pg_rca32_fa660_y1 | f_s_dadda_pg_rca32_fa660_y3;
  assign f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa660_y4 = f_s_dadda_pg_rca32_fa660_y4;
  assign f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa659_y4 = f_s_dadda_pg_rca32_fa659_y4;
  assign f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa658_y4 = f_s_dadda_pg_rca32_fa658_y4;
  assign f_s_dadda_pg_rca32_fa661_y0 = f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa660_y4 ^ f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa659_y4;
  assign f_s_dadda_pg_rca32_fa661_y1 = f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa660_y4 & f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa659_y4;
  assign f_s_dadda_pg_rca32_fa661_y2 = f_s_dadda_pg_rca32_fa661_y0 ^ f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa658_y4;
  assign f_s_dadda_pg_rca32_fa661_y3 = f_s_dadda_pg_rca32_fa661_y0 & f_s_dadda_pg_rca32_fa661_f_s_dadda_pg_rca32_fa658_y4;
  assign f_s_dadda_pg_rca32_fa661_y4 = f_s_dadda_pg_rca32_fa661_y1 | f_s_dadda_pg_rca32_fa661_y3;
  assign f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa657_y4 = f_s_dadda_pg_rca32_fa657_y4;
  assign f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa656_y4 = f_s_dadda_pg_rca32_fa656_y4;
  assign f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa655_y4 = f_s_dadda_pg_rca32_fa655_y4;
  assign f_s_dadda_pg_rca32_fa662_y0 = f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa657_y4 ^ f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa656_y4;
  assign f_s_dadda_pg_rca32_fa662_y1 = f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa657_y4 & f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa656_y4;
  assign f_s_dadda_pg_rca32_fa662_y2 = f_s_dadda_pg_rca32_fa662_y0 ^ f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa655_y4;
  assign f_s_dadda_pg_rca32_fa662_y3 = f_s_dadda_pg_rca32_fa662_y0 & f_s_dadda_pg_rca32_fa662_f_s_dadda_pg_rca32_fa655_y4;
  assign f_s_dadda_pg_rca32_fa662_y4 = f_s_dadda_pg_rca32_fa662_y1 | f_s_dadda_pg_rca32_fa662_y3;
  assign f_s_dadda_pg_rca32_nand_31_22_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_22_b_22 = b_22;
  assign f_s_dadda_pg_rca32_nand_31_22_y0 = ~(f_s_dadda_pg_rca32_nand_31_22_a_31 & f_s_dadda_pg_rca32_nand_31_22_b_22);
  assign f_s_dadda_pg_rca32_and_30_23_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_and_30_23_y0 = f_s_dadda_pg_rca32_and_30_23_a_30 & f_s_dadda_pg_rca32_and_30_23_b_23;
  assign f_s_dadda_pg_rca32_and_29_24_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_29_24_y0 = f_s_dadda_pg_rca32_and_29_24_a_29 & f_s_dadda_pg_rca32_and_29_24_b_24;
  assign f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_nand_31_22_y0 = f_s_dadda_pg_rca32_nand_31_22_y0;
  assign f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_and_30_23_y0 = f_s_dadda_pg_rca32_and_30_23_y0;
  assign f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_and_29_24_y0 = f_s_dadda_pg_rca32_and_29_24_y0;
  assign f_s_dadda_pg_rca32_fa663_y0 = f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_nand_31_22_y0 ^ f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_and_30_23_y0;
  assign f_s_dadda_pg_rca32_fa663_y1 = f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_nand_31_22_y0 & f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_and_30_23_y0;
  assign f_s_dadda_pg_rca32_fa663_y2 = f_s_dadda_pg_rca32_fa663_y0 ^ f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_and_29_24_y0;
  assign f_s_dadda_pg_rca32_fa663_y3 = f_s_dadda_pg_rca32_fa663_y0 & f_s_dadda_pg_rca32_fa663_f_s_dadda_pg_rca32_and_29_24_y0;
  assign f_s_dadda_pg_rca32_fa663_y4 = f_s_dadda_pg_rca32_fa663_y1 | f_s_dadda_pg_rca32_fa663_y3;
  assign f_s_dadda_pg_rca32_and_28_25_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_28_25_y0 = f_s_dadda_pg_rca32_and_28_25_a_28 & f_s_dadda_pg_rca32_and_28_25_b_25;
  assign f_s_dadda_pg_rca32_and_27_26_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_27_26_y0 = f_s_dadda_pg_rca32_and_27_26_a_27 & f_s_dadda_pg_rca32_and_27_26_b_26;
  assign f_s_dadda_pg_rca32_and_26_27_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_26_27_y0 = f_s_dadda_pg_rca32_and_26_27_a_26 & f_s_dadda_pg_rca32_and_26_27_b_27;
  assign f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_28_25_y0 = f_s_dadda_pg_rca32_and_28_25_y0;
  assign f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_27_26_y0 = f_s_dadda_pg_rca32_and_27_26_y0;
  assign f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_26_27_y0 = f_s_dadda_pg_rca32_and_26_27_y0;
  assign f_s_dadda_pg_rca32_fa664_y0 = f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_28_25_y0 ^ f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_27_26_y0;
  assign f_s_dadda_pg_rca32_fa664_y1 = f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_28_25_y0 & f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_27_26_y0;
  assign f_s_dadda_pg_rca32_fa664_y2 = f_s_dadda_pg_rca32_fa664_y0 ^ f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_26_27_y0;
  assign f_s_dadda_pg_rca32_fa664_y3 = f_s_dadda_pg_rca32_fa664_y0 & f_s_dadda_pg_rca32_fa664_f_s_dadda_pg_rca32_and_26_27_y0;
  assign f_s_dadda_pg_rca32_fa664_y4 = f_s_dadda_pg_rca32_fa664_y1 | f_s_dadda_pg_rca32_fa664_y3;
  assign f_s_dadda_pg_rca32_and_25_28_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_25_28_y0 = f_s_dadda_pg_rca32_and_25_28_a_25 & f_s_dadda_pg_rca32_and_25_28_b_28;
  assign f_s_dadda_pg_rca32_and_24_29_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_24_29_y0 = f_s_dadda_pg_rca32_and_24_29_a_24 & f_s_dadda_pg_rca32_and_24_29_b_29;
  assign f_s_dadda_pg_rca32_and_23_30_a_23 = a_23;
  assign f_s_dadda_pg_rca32_and_23_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_23_30_y0 = f_s_dadda_pg_rca32_and_23_30_a_23 & f_s_dadda_pg_rca32_and_23_30_b_30;
  assign f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_25_28_y0 = f_s_dadda_pg_rca32_and_25_28_y0;
  assign f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_24_29_y0 = f_s_dadda_pg_rca32_and_24_29_y0;
  assign f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_23_30_y0 = f_s_dadda_pg_rca32_and_23_30_y0;
  assign f_s_dadda_pg_rca32_fa665_y0 = f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_25_28_y0 ^ f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_24_29_y0;
  assign f_s_dadda_pg_rca32_fa665_y1 = f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_25_28_y0 & f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_24_29_y0;
  assign f_s_dadda_pg_rca32_fa665_y2 = f_s_dadda_pg_rca32_fa665_y0 ^ f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_23_30_y0;
  assign f_s_dadda_pg_rca32_fa665_y3 = f_s_dadda_pg_rca32_fa665_y0 & f_s_dadda_pg_rca32_fa665_f_s_dadda_pg_rca32_and_23_30_y0;
  assign f_s_dadda_pg_rca32_fa665_y4 = f_s_dadda_pg_rca32_fa665_y1 | f_s_dadda_pg_rca32_fa665_y3;
  assign f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa665_y4 = f_s_dadda_pg_rca32_fa665_y4;
  assign f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa664_y4 = f_s_dadda_pg_rca32_fa664_y4;
  assign f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa663_y4 = f_s_dadda_pg_rca32_fa663_y4;
  assign f_s_dadda_pg_rca32_fa666_y0 = f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa665_y4 ^ f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa664_y4;
  assign f_s_dadda_pg_rca32_fa666_y1 = f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa665_y4 & f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa664_y4;
  assign f_s_dadda_pg_rca32_fa666_y2 = f_s_dadda_pg_rca32_fa666_y0 ^ f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa663_y4;
  assign f_s_dadda_pg_rca32_fa666_y3 = f_s_dadda_pg_rca32_fa666_y0 & f_s_dadda_pg_rca32_fa666_f_s_dadda_pg_rca32_fa663_y4;
  assign f_s_dadda_pg_rca32_fa666_y4 = f_s_dadda_pg_rca32_fa666_y1 | f_s_dadda_pg_rca32_fa666_y3;
  assign f_s_dadda_pg_rca32_nand_31_23_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_23_b_23 = b_23;
  assign f_s_dadda_pg_rca32_nand_31_23_y0 = ~(f_s_dadda_pg_rca32_nand_31_23_a_31 & f_s_dadda_pg_rca32_nand_31_23_b_23);
  assign f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_fa662_y4 = f_s_dadda_pg_rca32_fa662_y4;
  assign f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_fa661_y4 = f_s_dadda_pg_rca32_fa661_y4;
  assign f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_nand_31_23_y0 = f_s_dadda_pg_rca32_nand_31_23_y0;
  assign f_s_dadda_pg_rca32_fa667_y0 = f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_fa662_y4 ^ f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_fa661_y4;
  assign f_s_dadda_pg_rca32_fa667_y1 = f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_fa662_y4 & f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_fa661_y4;
  assign f_s_dadda_pg_rca32_fa667_y2 = f_s_dadda_pg_rca32_fa667_y0 ^ f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_nand_31_23_y0;
  assign f_s_dadda_pg_rca32_fa667_y3 = f_s_dadda_pg_rca32_fa667_y0 & f_s_dadda_pg_rca32_fa667_f_s_dadda_pg_rca32_nand_31_23_y0;
  assign f_s_dadda_pg_rca32_fa667_y4 = f_s_dadda_pg_rca32_fa667_y1 | f_s_dadda_pg_rca32_fa667_y3;
  assign f_s_dadda_pg_rca32_and_30_24_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_and_30_24_y0 = f_s_dadda_pg_rca32_and_30_24_a_30 & f_s_dadda_pg_rca32_and_30_24_b_24;
  assign f_s_dadda_pg_rca32_and_29_25_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_29_25_y0 = f_s_dadda_pg_rca32_and_29_25_a_29 & f_s_dadda_pg_rca32_and_29_25_b_25;
  assign f_s_dadda_pg_rca32_and_28_26_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_28_26_y0 = f_s_dadda_pg_rca32_and_28_26_a_28 & f_s_dadda_pg_rca32_and_28_26_b_26;
  assign f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_30_24_y0 = f_s_dadda_pg_rca32_and_30_24_y0;
  assign f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_29_25_y0 = f_s_dadda_pg_rca32_and_29_25_y0;
  assign f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_28_26_y0 = f_s_dadda_pg_rca32_and_28_26_y0;
  assign f_s_dadda_pg_rca32_fa668_y0 = f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_30_24_y0 ^ f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_29_25_y0;
  assign f_s_dadda_pg_rca32_fa668_y1 = f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_30_24_y0 & f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_29_25_y0;
  assign f_s_dadda_pg_rca32_fa668_y2 = f_s_dadda_pg_rca32_fa668_y0 ^ f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_28_26_y0;
  assign f_s_dadda_pg_rca32_fa668_y3 = f_s_dadda_pg_rca32_fa668_y0 & f_s_dadda_pg_rca32_fa668_f_s_dadda_pg_rca32_and_28_26_y0;
  assign f_s_dadda_pg_rca32_fa668_y4 = f_s_dadda_pg_rca32_fa668_y1 | f_s_dadda_pg_rca32_fa668_y3;
  assign f_s_dadda_pg_rca32_and_27_27_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_27_27_y0 = f_s_dadda_pg_rca32_and_27_27_a_27 & f_s_dadda_pg_rca32_and_27_27_b_27;
  assign f_s_dadda_pg_rca32_and_26_28_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_26_28_y0 = f_s_dadda_pg_rca32_and_26_28_a_26 & f_s_dadda_pg_rca32_and_26_28_b_28;
  assign f_s_dadda_pg_rca32_and_25_29_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_25_29_y0 = f_s_dadda_pg_rca32_and_25_29_a_25 & f_s_dadda_pg_rca32_and_25_29_b_29;
  assign f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_27_27_y0 = f_s_dadda_pg_rca32_and_27_27_y0;
  assign f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_26_28_y0 = f_s_dadda_pg_rca32_and_26_28_y0;
  assign f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_25_29_y0 = f_s_dadda_pg_rca32_and_25_29_y0;
  assign f_s_dadda_pg_rca32_fa669_y0 = f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_27_27_y0 ^ f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_26_28_y0;
  assign f_s_dadda_pg_rca32_fa669_y1 = f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_27_27_y0 & f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_26_28_y0;
  assign f_s_dadda_pg_rca32_fa669_y2 = f_s_dadda_pg_rca32_fa669_y0 ^ f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_25_29_y0;
  assign f_s_dadda_pg_rca32_fa669_y3 = f_s_dadda_pg_rca32_fa669_y0 & f_s_dadda_pg_rca32_fa669_f_s_dadda_pg_rca32_and_25_29_y0;
  assign f_s_dadda_pg_rca32_fa669_y4 = f_s_dadda_pg_rca32_fa669_y1 | f_s_dadda_pg_rca32_fa669_y3;
  assign f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa669_y4 = f_s_dadda_pg_rca32_fa669_y4;
  assign f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa668_y4 = f_s_dadda_pg_rca32_fa668_y4;
  assign f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa667_y4 = f_s_dadda_pg_rca32_fa667_y4;
  assign f_s_dadda_pg_rca32_fa670_y0 = f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa669_y4 ^ f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa668_y4;
  assign f_s_dadda_pg_rca32_fa670_y1 = f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa669_y4 & f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa668_y4;
  assign f_s_dadda_pg_rca32_fa670_y2 = f_s_dadda_pg_rca32_fa670_y0 ^ f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa667_y4;
  assign f_s_dadda_pg_rca32_fa670_y3 = f_s_dadda_pg_rca32_fa670_y0 & f_s_dadda_pg_rca32_fa670_f_s_dadda_pg_rca32_fa667_y4;
  assign f_s_dadda_pg_rca32_fa670_y4 = f_s_dadda_pg_rca32_fa670_y1 | f_s_dadda_pg_rca32_fa670_y3;
  assign f_s_dadda_pg_rca32_nand_31_24_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_24_b_24 = b_24;
  assign f_s_dadda_pg_rca32_nand_31_24_y0 = ~(f_s_dadda_pg_rca32_nand_31_24_a_31 & f_s_dadda_pg_rca32_nand_31_24_b_24);
  assign f_s_dadda_pg_rca32_and_30_25_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_and_30_25_y0 = f_s_dadda_pg_rca32_and_30_25_a_30 & f_s_dadda_pg_rca32_and_30_25_b_25;
  assign f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_fa666_y4 = f_s_dadda_pg_rca32_fa666_y4;
  assign f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_nand_31_24_y0 = f_s_dadda_pg_rca32_nand_31_24_y0;
  assign f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_and_30_25_y0 = f_s_dadda_pg_rca32_and_30_25_y0;
  assign f_s_dadda_pg_rca32_fa671_y0 = f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_fa666_y4 ^ f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_nand_31_24_y0;
  assign f_s_dadda_pg_rca32_fa671_y1 = f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_fa666_y4 & f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_nand_31_24_y0;
  assign f_s_dadda_pg_rca32_fa671_y2 = f_s_dadda_pg_rca32_fa671_y0 ^ f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_and_30_25_y0;
  assign f_s_dadda_pg_rca32_fa671_y3 = f_s_dadda_pg_rca32_fa671_y0 & f_s_dadda_pg_rca32_fa671_f_s_dadda_pg_rca32_and_30_25_y0;
  assign f_s_dadda_pg_rca32_fa671_y4 = f_s_dadda_pg_rca32_fa671_y1 | f_s_dadda_pg_rca32_fa671_y3;
  assign f_s_dadda_pg_rca32_and_29_26_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_29_26_y0 = f_s_dadda_pg_rca32_and_29_26_a_29 & f_s_dadda_pg_rca32_and_29_26_b_26;
  assign f_s_dadda_pg_rca32_and_28_27_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_28_27_y0 = f_s_dadda_pg_rca32_and_28_27_a_28 & f_s_dadda_pg_rca32_and_28_27_b_27;
  assign f_s_dadda_pg_rca32_and_27_28_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_27_28_y0 = f_s_dadda_pg_rca32_and_27_28_a_27 & f_s_dadda_pg_rca32_and_27_28_b_28;
  assign f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_29_26_y0 = f_s_dadda_pg_rca32_and_29_26_y0;
  assign f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_28_27_y0 = f_s_dadda_pg_rca32_and_28_27_y0;
  assign f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_27_28_y0 = f_s_dadda_pg_rca32_and_27_28_y0;
  assign f_s_dadda_pg_rca32_fa672_y0 = f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_29_26_y0 ^ f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_28_27_y0;
  assign f_s_dadda_pg_rca32_fa672_y1 = f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_29_26_y0 & f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_28_27_y0;
  assign f_s_dadda_pg_rca32_fa672_y2 = f_s_dadda_pg_rca32_fa672_y0 ^ f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_27_28_y0;
  assign f_s_dadda_pg_rca32_fa672_y3 = f_s_dadda_pg_rca32_fa672_y0 & f_s_dadda_pg_rca32_fa672_f_s_dadda_pg_rca32_and_27_28_y0;
  assign f_s_dadda_pg_rca32_fa672_y4 = f_s_dadda_pg_rca32_fa672_y1 | f_s_dadda_pg_rca32_fa672_y3;
  assign f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa672_y4 = f_s_dadda_pg_rca32_fa672_y4;
  assign f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa671_y4 = f_s_dadda_pg_rca32_fa671_y4;
  assign f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa670_y4 = f_s_dadda_pg_rca32_fa670_y4;
  assign f_s_dadda_pg_rca32_fa673_y0 = f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa672_y4 ^ f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa671_y4;
  assign f_s_dadda_pg_rca32_fa673_y1 = f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa672_y4 & f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa671_y4;
  assign f_s_dadda_pg_rca32_fa673_y2 = f_s_dadda_pg_rca32_fa673_y0 ^ f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa670_y4;
  assign f_s_dadda_pg_rca32_fa673_y3 = f_s_dadda_pg_rca32_fa673_y0 & f_s_dadda_pg_rca32_fa673_f_s_dadda_pg_rca32_fa670_y4;
  assign f_s_dadda_pg_rca32_fa673_y4 = f_s_dadda_pg_rca32_fa673_y1 | f_s_dadda_pg_rca32_fa673_y3;
  assign f_s_dadda_pg_rca32_nand_31_25_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_25_b_25 = b_25;
  assign f_s_dadda_pg_rca32_nand_31_25_y0 = ~(f_s_dadda_pg_rca32_nand_31_25_a_31 & f_s_dadda_pg_rca32_nand_31_25_b_25);
  assign f_s_dadda_pg_rca32_and_30_26_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_and_30_26_y0 = f_s_dadda_pg_rca32_and_30_26_a_30 & f_s_dadda_pg_rca32_and_30_26_b_26;
  assign f_s_dadda_pg_rca32_and_29_27_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_29_27_y0 = f_s_dadda_pg_rca32_and_29_27_a_29 & f_s_dadda_pg_rca32_and_29_27_b_27;
  assign f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_nand_31_25_y0 = f_s_dadda_pg_rca32_nand_31_25_y0;
  assign f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_and_30_26_y0 = f_s_dadda_pg_rca32_and_30_26_y0;
  assign f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_and_29_27_y0 = f_s_dadda_pg_rca32_and_29_27_y0;
  assign f_s_dadda_pg_rca32_fa674_y0 = f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_nand_31_25_y0 ^ f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_and_30_26_y0;
  assign f_s_dadda_pg_rca32_fa674_y1 = f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_nand_31_25_y0 & f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_and_30_26_y0;
  assign f_s_dadda_pg_rca32_fa674_y2 = f_s_dadda_pg_rca32_fa674_y0 ^ f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_and_29_27_y0;
  assign f_s_dadda_pg_rca32_fa674_y3 = f_s_dadda_pg_rca32_fa674_y0 & f_s_dadda_pg_rca32_fa674_f_s_dadda_pg_rca32_and_29_27_y0;
  assign f_s_dadda_pg_rca32_fa674_y4 = f_s_dadda_pg_rca32_fa674_y1 | f_s_dadda_pg_rca32_fa674_y3;
  assign f_s_dadda_pg_rca32_nand_31_26_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_26_b_26 = b_26;
  assign f_s_dadda_pg_rca32_nand_31_26_y0 = ~(f_s_dadda_pg_rca32_nand_31_26_a_31 & f_s_dadda_pg_rca32_nand_31_26_b_26);
  assign f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_fa674_y4 = f_s_dadda_pg_rca32_fa674_y4;
  assign f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_fa673_y4 = f_s_dadda_pg_rca32_fa673_y4;
  assign f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_nand_31_26_y0 = f_s_dadda_pg_rca32_nand_31_26_y0;
  assign f_s_dadda_pg_rca32_fa675_y0 = f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_fa674_y4 ^ f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_fa673_y4;
  assign f_s_dadda_pg_rca32_fa675_y1 = f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_fa674_y4 & f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_fa673_y4;
  assign f_s_dadda_pg_rca32_fa675_y2 = f_s_dadda_pg_rca32_fa675_y0 ^ f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_nand_31_26_y0;
  assign f_s_dadda_pg_rca32_fa675_y3 = f_s_dadda_pg_rca32_fa675_y0 & f_s_dadda_pg_rca32_fa675_f_s_dadda_pg_rca32_nand_31_26_y0;
  assign f_s_dadda_pg_rca32_fa675_y4 = f_s_dadda_pg_rca32_fa675_y1 | f_s_dadda_pg_rca32_fa675_y3;
  assign f_s_dadda_pg_rca32_and_4_0_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_4_0_y0 = f_s_dadda_pg_rca32_and_4_0_a_4 & f_s_dadda_pg_rca32_and_4_0_b_0;
  assign f_s_dadda_pg_rca32_and_3_1_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_3_1_y0 = f_s_dadda_pg_rca32_and_3_1_a_3 & f_s_dadda_pg_rca32_and_3_1_b_1;
  assign f_s_dadda_pg_rca32_ha26_f_s_dadda_pg_rca32_and_4_0_y0 = f_s_dadda_pg_rca32_and_4_0_y0;
  assign f_s_dadda_pg_rca32_ha26_f_s_dadda_pg_rca32_and_3_1_y0 = f_s_dadda_pg_rca32_and_3_1_y0;
  assign f_s_dadda_pg_rca32_ha26_y0 = f_s_dadda_pg_rca32_ha26_f_s_dadda_pg_rca32_and_4_0_y0 ^ f_s_dadda_pg_rca32_ha26_f_s_dadda_pg_rca32_and_3_1_y0;
  assign f_s_dadda_pg_rca32_ha26_y1 = f_s_dadda_pg_rca32_ha26_f_s_dadda_pg_rca32_and_4_0_y0 & f_s_dadda_pg_rca32_ha26_f_s_dadda_pg_rca32_and_3_1_y0;
  assign f_s_dadda_pg_rca32_and_5_0_a_5 = a_5;
  assign f_s_dadda_pg_rca32_and_5_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_5_0_y0 = f_s_dadda_pg_rca32_and_5_0_a_5 & f_s_dadda_pg_rca32_and_5_0_b_0;
  assign f_s_dadda_pg_rca32_and_4_1_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_4_1_y0 = f_s_dadda_pg_rca32_and_4_1_a_4 & f_s_dadda_pg_rca32_and_4_1_b_1;
  assign f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_ha26_y1 = f_s_dadda_pg_rca32_ha26_y1;
  assign f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_and_5_0_y0 = f_s_dadda_pg_rca32_and_5_0_y0;
  assign f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_and_4_1_y0 = f_s_dadda_pg_rca32_and_4_1_y0;
  assign f_s_dadda_pg_rca32_fa676_y0 = f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_ha26_y1 ^ f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_and_5_0_y0;
  assign f_s_dadda_pg_rca32_fa676_y1 = f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_ha26_y1 & f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_and_5_0_y0;
  assign f_s_dadda_pg_rca32_fa676_y2 = f_s_dadda_pg_rca32_fa676_y0 ^ f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_and_4_1_y0;
  assign f_s_dadda_pg_rca32_fa676_y3 = f_s_dadda_pg_rca32_fa676_y0 & f_s_dadda_pg_rca32_fa676_f_s_dadda_pg_rca32_and_4_1_y0;
  assign f_s_dadda_pg_rca32_fa676_y4 = f_s_dadda_pg_rca32_fa676_y1 | f_s_dadda_pg_rca32_fa676_y3;
  assign f_s_dadda_pg_rca32_and_3_2_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_3_2_y0 = f_s_dadda_pg_rca32_and_3_2_a_3 & f_s_dadda_pg_rca32_and_3_2_b_2;
  assign f_s_dadda_pg_rca32_and_2_3_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_2_3_y0 = f_s_dadda_pg_rca32_and_2_3_a_2 & f_s_dadda_pg_rca32_and_2_3_b_3;
  assign f_s_dadda_pg_rca32_ha27_f_s_dadda_pg_rca32_and_3_2_y0 = f_s_dadda_pg_rca32_and_3_2_y0;
  assign f_s_dadda_pg_rca32_ha27_f_s_dadda_pg_rca32_and_2_3_y0 = f_s_dadda_pg_rca32_and_2_3_y0;
  assign f_s_dadda_pg_rca32_ha27_y0 = f_s_dadda_pg_rca32_ha27_f_s_dadda_pg_rca32_and_3_2_y0 ^ f_s_dadda_pg_rca32_ha27_f_s_dadda_pg_rca32_and_2_3_y0;
  assign f_s_dadda_pg_rca32_ha27_y1 = f_s_dadda_pg_rca32_ha27_f_s_dadda_pg_rca32_and_3_2_y0 & f_s_dadda_pg_rca32_ha27_f_s_dadda_pg_rca32_and_2_3_y0;
  assign f_s_dadda_pg_rca32_and_4_2_a_4 = a_4;
  assign f_s_dadda_pg_rca32_and_4_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_4_2_y0 = f_s_dadda_pg_rca32_and_4_2_a_4 & f_s_dadda_pg_rca32_and_4_2_b_2;
  assign f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_ha27_y1 = f_s_dadda_pg_rca32_ha27_y1;
  assign f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_fa676_y4 = f_s_dadda_pg_rca32_fa676_y4;
  assign f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_and_4_2_y0 = f_s_dadda_pg_rca32_and_4_2_y0;
  assign f_s_dadda_pg_rca32_fa677_y0 = f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_ha27_y1 ^ f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_fa676_y4;
  assign f_s_dadda_pg_rca32_fa677_y1 = f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_ha27_y1 & f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_fa676_y4;
  assign f_s_dadda_pg_rca32_fa677_y2 = f_s_dadda_pg_rca32_fa677_y0 ^ f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_and_4_2_y0;
  assign f_s_dadda_pg_rca32_fa677_y3 = f_s_dadda_pg_rca32_fa677_y0 & f_s_dadda_pg_rca32_fa677_f_s_dadda_pg_rca32_and_4_2_y0;
  assign f_s_dadda_pg_rca32_fa677_y4 = f_s_dadda_pg_rca32_fa677_y1 | f_s_dadda_pg_rca32_fa677_y3;
  assign f_s_dadda_pg_rca32_and_3_3_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_3_3_y0 = f_s_dadda_pg_rca32_and_3_3_a_3 & f_s_dadda_pg_rca32_and_3_3_b_3;
  assign f_s_dadda_pg_rca32_and_2_4_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_2_4_y0 = f_s_dadda_pg_rca32_and_2_4_a_2 & f_s_dadda_pg_rca32_and_2_4_b_4;
  assign f_s_dadda_pg_rca32_and_1_5_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_1_5_y0 = f_s_dadda_pg_rca32_and_1_5_a_1 & f_s_dadda_pg_rca32_and_1_5_b_5;
  assign f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_3_3_y0 = f_s_dadda_pg_rca32_and_3_3_y0;
  assign f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_2_4_y0 = f_s_dadda_pg_rca32_and_2_4_y0;
  assign f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_1_5_y0 = f_s_dadda_pg_rca32_and_1_5_y0;
  assign f_s_dadda_pg_rca32_fa678_y0 = f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_3_3_y0 ^ f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_2_4_y0;
  assign f_s_dadda_pg_rca32_fa678_y1 = f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_3_3_y0 & f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_2_4_y0;
  assign f_s_dadda_pg_rca32_fa678_y2 = f_s_dadda_pg_rca32_fa678_y0 ^ f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_1_5_y0;
  assign f_s_dadda_pg_rca32_fa678_y3 = f_s_dadda_pg_rca32_fa678_y0 & f_s_dadda_pg_rca32_fa678_f_s_dadda_pg_rca32_and_1_5_y0;
  assign f_s_dadda_pg_rca32_fa678_y4 = f_s_dadda_pg_rca32_fa678_y1 | f_s_dadda_pg_rca32_fa678_y3;
  assign f_s_dadda_pg_rca32_and_3_4_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_3_4_y0 = f_s_dadda_pg_rca32_and_3_4_a_3 & f_s_dadda_pg_rca32_and_3_4_b_4;
  assign f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_fa678_y4 = f_s_dadda_pg_rca32_fa678_y4;
  assign f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_fa677_y4 = f_s_dadda_pg_rca32_fa677_y4;
  assign f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_and_3_4_y0 = f_s_dadda_pg_rca32_and_3_4_y0;
  assign f_s_dadda_pg_rca32_fa679_y0 = f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_fa678_y4 ^ f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_fa677_y4;
  assign f_s_dadda_pg_rca32_fa679_y1 = f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_fa678_y4 & f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_fa677_y4;
  assign f_s_dadda_pg_rca32_fa679_y2 = f_s_dadda_pg_rca32_fa679_y0 ^ f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_and_3_4_y0;
  assign f_s_dadda_pg_rca32_fa679_y3 = f_s_dadda_pg_rca32_fa679_y0 & f_s_dadda_pg_rca32_fa679_f_s_dadda_pg_rca32_and_3_4_y0;
  assign f_s_dadda_pg_rca32_fa679_y4 = f_s_dadda_pg_rca32_fa679_y1 | f_s_dadda_pg_rca32_fa679_y3;
  assign f_s_dadda_pg_rca32_and_2_5_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_2_5_y0 = f_s_dadda_pg_rca32_and_2_5_a_2 & f_s_dadda_pg_rca32_and_2_5_b_5;
  assign f_s_dadda_pg_rca32_and_1_6_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_1_6_y0 = f_s_dadda_pg_rca32_and_1_6_a_1 & f_s_dadda_pg_rca32_and_1_6_b_6;
  assign f_s_dadda_pg_rca32_and_0_7_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_0_7_y0 = f_s_dadda_pg_rca32_and_0_7_a_0 & f_s_dadda_pg_rca32_and_0_7_b_7;
  assign f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_2_5_y0 = f_s_dadda_pg_rca32_and_2_5_y0;
  assign f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_1_6_y0 = f_s_dadda_pg_rca32_and_1_6_y0;
  assign f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_0_7_y0 = f_s_dadda_pg_rca32_and_0_7_y0;
  assign f_s_dadda_pg_rca32_fa680_y0 = f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_2_5_y0 ^ f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_1_6_y0;
  assign f_s_dadda_pg_rca32_fa680_y1 = f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_2_5_y0 & f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_1_6_y0;
  assign f_s_dadda_pg_rca32_fa680_y2 = f_s_dadda_pg_rca32_fa680_y0 ^ f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_0_7_y0;
  assign f_s_dadda_pg_rca32_fa680_y3 = f_s_dadda_pg_rca32_fa680_y0 & f_s_dadda_pg_rca32_fa680_f_s_dadda_pg_rca32_and_0_7_y0;
  assign f_s_dadda_pg_rca32_fa680_y4 = f_s_dadda_pg_rca32_fa680_y1 | f_s_dadda_pg_rca32_fa680_y3;
  assign f_s_dadda_pg_rca32_and_2_6_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_2_6_y0 = f_s_dadda_pg_rca32_and_2_6_a_2 & f_s_dadda_pg_rca32_and_2_6_b_6;
  assign f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_fa680_y4 = f_s_dadda_pg_rca32_fa680_y4;
  assign f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_fa679_y4 = f_s_dadda_pg_rca32_fa679_y4;
  assign f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_and_2_6_y0 = f_s_dadda_pg_rca32_and_2_6_y0;
  assign f_s_dadda_pg_rca32_fa681_y0 = f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_fa680_y4 ^ f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_fa679_y4;
  assign f_s_dadda_pg_rca32_fa681_y1 = f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_fa680_y4 & f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_fa679_y4;
  assign f_s_dadda_pg_rca32_fa681_y2 = f_s_dadda_pg_rca32_fa681_y0 ^ f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_and_2_6_y0;
  assign f_s_dadda_pg_rca32_fa681_y3 = f_s_dadda_pg_rca32_fa681_y0 & f_s_dadda_pg_rca32_fa681_f_s_dadda_pg_rca32_and_2_6_y0;
  assign f_s_dadda_pg_rca32_fa681_y4 = f_s_dadda_pg_rca32_fa681_y1 | f_s_dadda_pg_rca32_fa681_y3;
  assign f_s_dadda_pg_rca32_and_1_7_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_7_b_7 = b_7;
  assign f_s_dadda_pg_rca32_and_1_7_y0 = f_s_dadda_pg_rca32_and_1_7_a_1 & f_s_dadda_pg_rca32_and_1_7_b_7;
  assign f_s_dadda_pg_rca32_and_0_8_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_0_8_y0 = f_s_dadda_pg_rca32_and_0_8_a_0 & f_s_dadda_pg_rca32_and_0_8_b_8;
  assign f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_and_1_7_y0 = f_s_dadda_pg_rca32_and_1_7_y0;
  assign f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_and_0_8_y0 = f_s_dadda_pg_rca32_and_0_8_y0;
  assign f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_fa17_y2 = f_s_dadda_pg_rca32_fa17_y2;
  assign f_s_dadda_pg_rca32_fa682_y0 = f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_and_1_7_y0 ^ f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_and_0_8_y0;
  assign f_s_dadda_pg_rca32_fa682_y1 = f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_and_1_7_y0 & f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_and_0_8_y0;
  assign f_s_dadda_pg_rca32_fa682_y2 = f_s_dadda_pg_rca32_fa682_y0 ^ f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_fa17_y2;
  assign f_s_dadda_pg_rca32_fa682_y3 = f_s_dadda_pg_rca32_fa682_y0 & f_s_dadda_pg_rca32_fa682_f_s_dadda_pg_rca32_fa17_y2;
  assign f_s_dadda_pg_rca32_fa682_y4 = f_s_dadda_pg_rca32_fa682_y1 | f_s_dadda_pg_rca32_fa682_y3;
  assign f_s_dadda_pg_rca32_and_1_8_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_8_b_8 = b_8;
  assign f_s_dadda_pg_rca32_and_1_8_y0 = f_s_dadda_pg_rca32_and_1_8_a_1 & f_s_dadda_pg_rca32_and_1_8_b_8;
  assign f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_fa682_y4 = f_s_dadda_pg_rca32_fa682_y4;
  assign f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_fa681_y4 = f_s_dadda_pg_rca32_fa681_y4;
  assign f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_and_1_8_y0 = f_s_dadda_pg_rca32_and_1_8_y0;
  assign f_s_dadda_pg_rca32_fa683_y0 = f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_fa682_y4 ^ f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_fa681_y4;
  assign f_s_dadda_pg_rca32_fa683_y1 = f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_fa682_y4 & f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_fa681_y4;
  assign f_s_dadda_pg_rca32_fa683_y2 = f_s_dadda_pg_rca32_fa683_y0 ^ f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_and_1_8_y0;
  assign f_s_dadda_pg_rca32_fa683_y3 = f_s_dadda_pg_rca32_fa683_y0 & f_s_dadda_pg_rca32_fa683_f_s_dadda_pg_rca32_and_1_8_y0;
  assign f_s_dadda_pg_rca32_fa683_y4 = f_s_dadda_pg_rca32_fa683_y1 | f_s_dadda_pg_rca32_fa683_y3;
  assign f_s_dadda_pg_rca32_and_0_9_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_9_b_9 = b_9;
  assign f_s_dadda_pg_rca32_and_0_9_y0 = f_s_dadda_pg_rca32_and_0_9_a_0 & f_s_dadda_pg_rca32_and_0_9_b_9;
  assign f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_and_0_9_y0 = f_s_dadda_pg_rca32_and_0_9_y0;
  assign f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_fa19_y2 = f_s_dadda_pg_rca32_fa19_y2;
  assign f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_fa20_y2 = f_s_dadda_pg_rca32_fa20_y2;
  assign f_s_dadda_pg_rca32_fa684_y0 = f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_and_0_9_y0 ^ f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_fa19_y2;
  assign f_s_dadda_pg_rca32_fa684_y1 = f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_and_0_9_y0 & f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_fa19_y2;
  assign f_s_dadda_pg_rca32_fa684_y2 = f_s_dadda_pg_rca32_fa684_y0 ^ f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_fa20_y2;
  assign f_s_dadda_pg_rca32_fa684_y3 = f_s_dadda_pg_rca32_fa684_y0 & f_s_dadda_pg_rca32_fa684_f_s_dadda_pg_rca32_fa20_y2;
  assign f_s_dadda_pg_rca32_fa684_y4 = f_s_dadda_pg_rca32_fa684_y1 | f_s_dadda_pg_rca32_fa684_y3;
  assign f_s_dadda_pg_rca32_and_0_10_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_10_b_10 = b_10;
  assign f_s_dadda_pg_rca32_and_0_10_y0 = f_s_dadda_pg_rca32_and_0_10_a_0 & f_s_dadda_pg_rca32_and_0_10_b_10;
  assign f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_fa684_y4 = f_s_dadda_pg_rca32_fa684_y4;
  assign f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_fa683_y4 = f_s_dadda_pg_rca32_fa683_y4;
  assign f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_and_0_10_y0 = f_s_dadda_pg_rca32_and_0_10_y0;
  assign f_s_dadda_pg_rca32_fa685_y0 = f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_fa684_y4 ^ f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_fa683_y4;
  assign f_s_dadda_pg_rca32_fa685_y1 = f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_fa684_y4 & f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_fa683_y4;
  assign f_s_dadda_pg_rca32_fa685_y2 = f_s_dadda_pg_rca32_fa685_y0 ^ f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_and_0_10_y0;
  assign f_s_dadda_pg_rca32_fa685_y3 = f_s_dadda_pg_rca32_fa685_y0 & f_s_dadda_pg_rca32_fa685_f_s_dadda_pg_rca32_and_0_10_y0;
  assign f_s_dadda_pg_rca32_fa685_y4 = f_s_dadda_pg_rca32_fa685_y1 | f_s_dadda_pg_rca32_fa685_y3;
  assign f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa22_y2 = f_s_dadda_pg_rca32_fa22_y2;
  assign f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa23_y2 = f_s_dadda_pg_rca32_fa23_y2;
  assign f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa24_y2 = f_s_dadda_pg_rca32_fa24_y2;
  assign f_s_dadda_pg_rca32_fa686_y0 = f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa22_y2 ^ f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa23_y2;
  assign f_s_dadda_pg_rca32_fa686_y1 = f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa22_y2 & f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa23_y2;
  assign f_s_dadda_pg_rca32_fa686_y2 = f_s_dadda_pg_rca32_fa686_y0 ^ f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa24_y2;
  assign f_s_dadda_pg_rca32_fa686_y3 = f_s_dadda_pg_rca32_fa686_y0 & f_s_dadda_pg_rca32_fa686_f_s_dadda_pg_rca32_fa24_y2;
  assign f_s_dadda_pg_rca32_fa686_y4 = f_s_dadda_pg_rca32_fa686_y1 | f_s_dadda_pg_rca32_fa686_y3;
  assign f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa686_y4 = f_s_dadda_pg_rca32_fa686_y4;
  assign f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa685_y4 = f_s_dadda_pg_rca32_fa685_y4;
  assign f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa26_y2 = f_s_dadda_pg_rca32_fa26_y2;
  assign f_s_dadda_pg_rca32_fa687_y0 = f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa686_y4 ^ f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa685_y4;
  assign f_s_dadda_pg_rca32_fa687_y1 = f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa686_y4 & f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa685_y4;
  assign f_s_dadda_pg_rca32_fa687_y2 = f_s_dadda_pg_rca32_fa687_y0 ^ f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa26_y2;
  assign f_s_dadda_pg_rca32_fa687_y3 = f_s_dadda_pg_rca32_fa687_y0 & f_s_dadda_pg_rca32_fa687_f_s_dadda_pg_rca32_fa26_y2;
  assign f_s_dadda_pg_rca32_fa687_y4 = f_s_dadda_pg_rca32_fa687_y1 | f_s_dadda_pg_rca32_fa687_y3;
  assign f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa27_y2 = f_s_dadda_pg_rca32_fa27_y2;
  assign f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa28_y2 = f_s_dadda_pg_rca32_fa28_y2;
  assign f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa29_y2 = f_s_dadda_pg_rca32_fa29_y2;
  assign f_s_dadda_pg_rca32_fa688_y0 = f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa27_y2 ^ f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa28_y2;
  assign f_s_dadda_pg_rca32_fa688_y1 = f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa27_y2 & f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa28_y2;
  assign f_s_dadda_pg_rca32_fa688_y2 = f_s_dadda_pg_rca32_fa688_y0 ^ f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa29_y2;
  assign f_s_dadda_pg_rca32_fa688_y3 = f_s_dadda_pg_rca32_fa688_y0 & f_s_dadda_pg_rca32_fa688_f_s_dadda_pg_rca32_fa29_y2;
  assign f_s_dadda_pg_rca32_fa688_y4 = f_s_dadda_pg_rca32_fa688_y1 | f_s_dadda_pg_rca32_fa688_y3;
  assign f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa688_y4 = f_s_dadda_pg_rca32_fa688_y4;
  assign f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa687_y4 = f_s_dadda_pg_rca32_fa687_y4;
  assign f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa32_y2 = f_s_dadda_pg_rca32_fa32_y2;
  assign f_s_dadda_pg_rca32_fa689_y0 = f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa688_y4 ^ f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa687_y4;
  assign f_s_dadda_pg_rca32_fa689_y1 = f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa688_y4 & f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa687_y4;
  assign f_s_dadda_pg_rca32_fa689_y2 = f_s_dadda_pg_rca32_fa689_y0 ^ f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa32_y2;
  assign f_s_dadda_pg_rca32_fa689_y3 = f_s_dadda_pg_rca32_fa689_y0 & f_s_dadda_pg_rca32_fa689_f_s_dadda_pg_rca32_fa32_y2;
  assign f_s_dadda_pg_rca32_fa689_y4 = f_s_dadda_pg_rca32_fa689_y1 | f_s_dadda_pg_rca32_fa689_y3;
  assign f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa33_y2 = f_s_dadda_pg_rca32_fa33_y2;
  assign f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa34_y2 = f_s_dadda_pg_rca32_fa34_y2;
  assign f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa35_y2 = f_s_dadda_pg_rca32_fa35_y2;
  assign f_s_dadda_pg_rca32_fa690_y0 = f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa33_y2 ^ f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa34_y2;
  assign f_s_dadda_pg_rca32_fa690_y1 = f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa33_y2 & f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa34_y2;
  assign f_s_dadda_pg_rca32_fa690_y2 = f_s_dadda_pg_rca32_fa690_y0 ^ f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa35_y2;
  assign f_s_dadda_pg_rca32_fa690_y3 = f_s_dadda_pg_rca32_fa690_y0 & f_s_dadda_pg_rca32_fa690_f_s_dadda_pg_rca32_fa35_y2;
  assign f_s_dadda_pg_rca32_fa690_y4 = f_s_dadda_pg_rca32_fa690_y1 | f_s_dadda_pg_rca32_fa690_y3;
  assign f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa690_y4 = f_s_dadda_pg_rca32_fa690_y4;
  assign f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa689_y4 = f_s_dadda_pg_rca32_fa689_y4;
  assign f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa39_y2 = f_s_dadda_pg_rca32_fa39_y2;
  assign f_s_dadda_pg_rca32_fa691_y0 = f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa690_y4 ^ f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa689_y4;
  assign f_s_dadda_pg_rca32_fa691_y1 = f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa690_y4 & f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa689_y4;
  assign f_s_dadda_pg_rca32_fa691_y2 = f_s_dadda_pg_rca32_fa691_y0 ^ f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa39_y2;
  assign f_s_dadda_pg_rca32_fa691_y3 = f_s_dadda_pg_rca32_fa691_y0 & f_s_dadda_pg_rca32_fa691_f_s_dadda_pg_rca32_fa39_y2;
  assign f_s_dadda_pg_rca32_fa691_y4 = f_s_dadda_pg_rca32_fa691_y1 | f_s_dadda_pg_rca32_fa691_y3;
  assign f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa40_y2 = f_s_dadda_pg_rca32_fa40_y2;
  assign f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa41_y2 = f_s_dadda_pg_rca32_fa41_y2;
  assign f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa42_y2 = f_s_dadda_pg_rca32_fa42_y2;
  assign f_s_dadda_pg_rca32_fa692_y0 = f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa40_y2 ^ f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa41_y2;
  assign f_s_dadda_pg_rca32_fa692_y1 = f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa40_y2 & f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa41_y2;
  assign f_s_dadda_pg_rca32_fa692_y2 = f_s_dadda_pg_rca32_fa692_y0 ^ f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa42_y2;
  assign f_s_dadda_pg_rca32_fa692_y3 = f_s_dadda_pg_rca32_fa692_y0 & f_s_dadda_pg_rca32_fa692_f_s_dadda_pg_rca32_fa42_y2;
  assign f_s_dadda_pg_rca32_fa692_y4 = f_s_dadda_pg_rca32_fa692_y1 | f_s_dadda_pg_rca32_fa692_y3;
  assign f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa692_y4 = f_s_dadda_pg_rca32_fa692_y4;
  assign f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa691_y4 = f_s_dadda_pg_rca32_fa691_y4;
  assign f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa47_y2 = f_s_dadda_pg_rca32_fa47_y2;
  assign f_s_dadda_pg_rca32_fa693_y0 = f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa692_y4 ^ f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa691_y4;
  assign f_s_dadda_pg_rca32_fa693_y1 = f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa692_y4 & f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa691_y4;
  assign f_s_dadda_pg_rca32_fa693_y2 = f_s_dadda_pg_rca32_fa693_y0 ^ f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa47_y2;
  assign f_s_dadda_pg_rca32_fa693_y3 = f_s_dadda_pg_rca32_fa693_y0 & f_s_dadda_pg_rca32_fa693_f_s_dadda_pg_rca32_fa47_y2;
  assign f_s_dadda_pg_rca32_fa693_y4 = f_s_dadda_pg_rca32_fa693_y1 | f_s_dadda_pg_rca32_fa693_y3;
  assign f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa48_y2 = f_s_dadda_pg_rca32_fa48_y2;
  assign f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa49_y2 = f_s_dadda_pg_rca32_fa49_y2;
  assign f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa50_y2 = f_s_dadda_pg_rca32_fa50_y2;
  assign f_s_dadda_pg_rca32_fa694_y0 = f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa48_y2 ^ f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa49_y2;
  assign f_s_dadda_pg_rca32_fa694_y1 = f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa48_y2 & f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa49_y2;
  assign f_s_dadda_pg_rca32_fa694_y2 = f_s_dadda_pg_rca32_fa694_y0 ^ f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa50_y2;
  assign f_s_dadda_pg_rca32_fa694_y3 = f_s_dadda_pg_rca32_fa694_y0 & f_s_dadda_pg_rca32_fa694_f_s_dadda_pg_rca32_fa50_y2;
  assign f_s_dadda_pg_rca32_fa694_y4 = f_s_dadda_pg_rca32_fa694_y1 | f_s_dadda_pg_rca32_fa694_y3;
  assign f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa694_y4 = f_s_dadda_pg_rca32_fa694_y4;
  assign f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa693_y4 = f_s_dadda_pg_rca32_fa693_y4;
  assign f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa56_y2 = f_s_dadda_pg_rca32_fa56_y2;
  assign f_s_dadda_pg_rca32_fa695_y0 = f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa694_y4 ^ f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa693_y4;
  assign f_s_dadda_pg_rca32_fa695_y1 = f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa694_y4 & f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa693_y4;
  assign f_s_dadda_pg_rca32_fa695_y2 = f_s_dadda_pg_rca32_fa695_y0 ^ f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa56_y2;
  assign f_s_dadda_pg_rca32_fa695_y3 = f_s_dadda_pg_rca32_fa695_y0 & f_s_dadda_pg_rca32_fa695_f_s_dadda_pg_rca32_fa56_y2;
  assign f_s_dadda_pg_rca32_fa695_y4 = f_s_dadda_pg_rca32_fa695_y1 | f_s_dadda_pg_rca32_fa695_y3;
  assign f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa57_y2 = f_s_dadda_pg_rca32_fa57_y2;
  assign f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa58_y2 = f_s_dadda_pg_rca32_fa58_y2;
  assign f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa59_y2 = f_s_dadda_pg_rca32_fa59_y2;
  assign f_s_dadda_pg_rca32_fa696_y0 = f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa57_y2 ^ f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa58_y2;
  assign f_s_dadda_pg_rca32_fa696_y1 = f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa57_y2 & f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa58_y2;
  assign f_s_dadda_pg_rca32_fa696_y2 = f_s_dadda_pg_rca32_fa696_y0 ^ f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa59_y2;
  assign f_s_dadda_pg_rca32_fa696_y3 = f_s_dadda_pg_rca32_fa696_y0 & f_s_dadda_pg_rca32_fa696_f_s_dadda_pg_rca32_fa59_y2;
  assign f_s_dadda_pg_rca32_fa696_y4 = f_s_dadda_pg_rca32_fa696_y1 | f_s_dadda_pg_rca32_fa696_y3;
  assign f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa696_y4 = f_s_dadda_pg_rca32_fa696_y4;
  assign f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa695_y4 = f_s_dadda_pg_rca32_fa695_y4;
  assign f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa66_y2 = f_s_dadda_pg_rca32_fa66_y2;
  assign f_s_dadda_pg_rca32_fa697_y0 = f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa696_y4 ^ f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa695_y4;
  assign f_s_dadda_pg_rca32_fa697_y1 = f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa696_y4 & f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa695_y4;
  assign f_s_dadda_pg_rca32_fa697_y2 = f_s_dadda_pg_rca32_fa697_y0 ^ f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa66_y2;
  assign f_s_dadda_pg_rca32_fa697_y3 = f_s_dadda_pg_rca32_fa697_y0 & f_s_dadda_pg_rca32_fa697_f_s_dadda_pg_rca32_fa66_y2;
  assign f_s_dadda_pg_rca32_fa697_y4 = f_s_dadda_pg_rca32_fa697_y1 | f_s_dadda_pg_rca32_fa697_y3;
  assign f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa67_y2 = f_s_dadda_pg_rca32_fa67_y2;
  assign f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa68_y2 = f_s_dadda_pg_rca32_fa68_y2;
  assign f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa69_y2 = f_s_dadda_pg_rca32_fa69_y2;
  assign f_s_dadda_pg_rca32_fa698_y0 = f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa67_y2 ^ f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa68_y2;
  assign f_s_dadda_pg_rca32_fa698_y1 = f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa67_y2 & f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa68_y2;
  assign f_s_dadda_pg_rca32_fa698_y2 = f_s_dadda_pg_rca32_fa698_y0 ^ f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa69_y2;
  assign f_s_dadda_pg_rca32_fa698_y3 = f_s_dadda_pg_rca32_fa698_y0 & f_s_dadda_pg_rca32_fa698_f_s_dadda_pg_rca32_fa69_y2;
  assign f_s_dadda_pg_rca32_fa698_y4 = f_s_dadda_pg_rca32_fa698_y1 | f_s_dadda_pg_rca32_fa698_y3;
  assign f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa698_y4 = f_s_dadda_pg_rca32_fa698_y4;
  assign f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa697_y4 = f_s_dadda_pg_rca32_fa697_y4;
  assign f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa77_y2 = f_s_dadda_pg_rca32_fa77_y2;
  assign f_s_dadda_pg_rca32_fa699_y0 = f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa698_y4 ^ f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa697_y4;
  assign f_s_dadda_pg_rca32_fa699_y1 = f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa698_y4 & f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa697_y4;
  assign f_s_dadda_pg_rca32_fa699_y2 = f_s_dadda_pg_rca32_fa699_y0 ^ f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa77_y2;
  assign f_s_dadda_pg_rca32_fa699_y3 = f_s_dadda_pg_rca32_fa699_y0 & f_s_dadda_pg_rca32_fa699_f_s_dadda_pg_rca32_fa77_y2;
  assign f_s_dadda_pg_rca32_fa699_y4 = f_s_dadda_pg_rca32_fa699_y1 | f_s_dadda_pg_rca32_fa699_y3;
  assign f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa78_y2 = f_s_dadda_pg_rca32_fa78_y2;
  assign f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa79_y2 = f_s_dadda_pg_rca32_fa79_y2;
  assign f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa80_y2 = f_s_dadda_pg_rca32_fa80_y2;
  assign f_s_dadda_pg_rca32_fa700_y0 = f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa78_y2 ^ f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa79_y2;
  assign f_s_dadda_pg_rca32_fa700_y1 = f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa78_y2 & f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa79_y2;
  assign f_s_dadda_pg_rca32_fa700_y2 = f_s_dadda_pg_rca32_fa700_y0 ^ f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa80_y2;
  assign f_s_dadda_pg_rca32_fa700_y3 = f_s_dadda_pg_rca32_fa700_y0 & f_s_dadda_pg_rca32_fa700_f_s_dadda_pg_rca32_fa80_y2;
  assign f_s_dadda_pg_rca32_fa700_y4 = f_s_dadda_pg_rca32_fa700_y1 | f_s_dadda_pg_rca32_fa700_y3;
  assign f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa700_y4 = f_s_dadda_pg_rca32_fa700_y4;
  assign f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa699_y4 = f_s_dadda_pg_rca32_fa699_y4;
  assign f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa89_y2 = f_s_dadda_pg_rca32_fa89_y2;
  assign f_s_dadda_pg_rca32_fa701_y0 = f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa700_y4 ^ f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa699_y4;
  assign f_s_dadda_pg_rca32_fa701_y1 = f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa700_y4 & f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa699_y4;
  assign f_s_dadda_pg_rca32_fa701_y2 = f_s_dadda_pg_rca32_fa701_y0 ^ f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa89_y2;
  assign f_s_dadda_pg_rca32_fa701_y3 = f_s_dadda_pg_rca32_fa701_y0 & f_s_dadda_pg_rca32_fa701_f_s_dadda_pg_rca32_fa89_y2;
  assign f_s_dadda_pg_rca32_fa701_y4 = f_s_dadda_pg_rca32_fa701_y1 | f_s_dadda_pg_rca32_fa701_y3;
  assign f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa90_y2 = f_s_dadda_pg_rca32_fa90_y2;
  assign f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa91_y2 = f_s_dadda_pg_rca32_fa91_y2;
  assign f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa92_y2 = f_s_dadda_pg_rca32_fa92_y2;
  assign f_s_dadda_pg_rca32_fa702_y0 = f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa90_y2 ^ f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa91_y2;
  assign f_s_dadda_pg_rca32_fa702_y1 = f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa90_y2 & f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa91_y2;
  assign f_s_dadda_pg_rca32_fa702_y2 = f_s_dadda_pg_rca32_fa702_y0 ^ f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa92_y2;
  assign f_s_dadda_pg_rca32_fa702_y3 = f_s_dadda_pg_rca32_fa702_y0 & f_s_dadda_pg_rca32_fa702_f_s_dadda_pg_rca32_fa92_y2;
  assign f_s_dadda_pg_rca32_fa702_y4 = f_s_dadda_pg_rca32_fa702_y1 | f_s_dadda_pg_rca32_fa702_y3;
  assign f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa702_y4 = f_s_dadda_pg_rca32_fa702_y4;
  assign f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa701_y4 = f_s_dadda_pg_rca32_fa701_y4;
  assign f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa102_y2 = f_s_dadda_pg_rca32_fa102_y2;
  assign f_s_dadda_pg_rca32_fa703_y0 = f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa702_y4 ^ f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa701_y4;
  assign f_s_dadda_pg_rca32_fa703_y1 = f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa702_y4 & f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa701_y4;
  assign f_s_dadda_pg_rca32_fa703_y2 = f_s_dadda_pg_rca32_fa703_y0 ^ f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa102_y2;
  assign f_s_dadda_pg_rca32_fa703_y3 = f_s_dadda_pg_rca32_fa703_y0 & f_s_dadda_pg_rca32_fa703_f_s_dadda_pg_rca32_fa102_y2;
  assign f_s_dadda_pg_rca32_fa703_y4 = f_s_dadda_pg_rca32_fa703_y1 | f_s_dadda_pg_rca32_fa703_y3;
  assign f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa103_y2 = f_s_dadda_pg_rca32_fa103_y2;
  assign f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa104_y2 = f_s_dadda_pg_rca32_fa104_y2;
  assign f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa105_y2 = f_s_dadda_pg_rca32_fa105_y2;
  assign f_s_dadda_pg_rca32_fa704_y0 = f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa103_y2 ^ f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa104_y2;
  assign f_s_dadda_pg_rca32_fa704_y1 = f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa103_y2 & f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa104_y2;
  assign f_s_dadda_pg_rca32_fa704_y2 = f_s_dadda_pg_rca32_fa704_y0 ^ f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa105_y2;
  assign f_s_dadda_pg_rca32_fa704_y3 = f_s_dadda_pg_rca32_fa704_y0 & f_s_dadda_pg_rca32_fa704_f_s_dadda_pg_rca32_fa105_y2;
  assign f_s_dadda_pg_rca32_fa704_y4 = f_s_dadda_pg_rca32_fa704_y1 | f_s_dadda_pg_rca32_fa704_y3;
  assign f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa704_y4 = f_s_dadda_pg_rca32_fa704_y4;
  assign f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa703_y4 = f_s_dadda_pg_rca32_fa703_y4;
  assign f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa116_y2 = f_s_dadda_pg_rca32_fa116_y2;
  assign f_s_dadda_pg_rca32_fa705_y0 = f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa704_y4 ^ f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa703_y4;
  assign f_s_dadda_pg_rca32_fa705_y1 = f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa704_y4 & f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa703_y4;
  assign f_s_dadda_pg_rca32_fa705_y2 = f_s_dadda_pg_rca32_fa705_y0 ^ f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa116_y2;
  assign f_s_dadda_pg_rca32_fa705_y3 = f_s_dadda_pg_rca32_fa705_y0 & f_s_dadda_pg_rca32_fa705_f_s_dadda_pg_rca32_fa116_y2;
  assign f_s_dadda_pg_rca32_fa705_y4 = f_s_dadda_pg_rca32_fa705_y1 | f_s_dadda_pg_rca32_fa705_y3;
  assign f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa117_y2 = f_s_dadda_pg_rca32_fa117_y2;
  assign f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa118_y2 = f_s_dadda_pg_rca32_fa118_y2;
  assign f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa119_y2 = f_s_dadda_pg_rca32_fa119_y2;
  assign f_s_dadda_pg_rca32_fa706_y0 = f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa117_y2 ^ f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa118_y2;
  assign f_s_dadda_pg_rca32_fa706_y1 = f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa117_y2 & f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa118_y2;
  assign f_s_dadda_pg_rca32_fa706_y2 = f_s_dadda_pg_rca32_fa706_y0 ^ f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa119_y2;
  assign f_s_dadda_pg_rca32_fa706_y3 = f_s_dadda_pg_rca32_fa706_y0 & f_s_dadda_pg_rca32_fa706_f_s_dadda_pg_rca32_fa119_y2;
  assign f_s_dadda_pg_rca32_fa706_y4 = f_s_dadda_pg_rca32_fa706_y1 | f_s_dadda_pg_rca32_fa706_y3;
  assign f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa706_y4 = f_s_dadda_pg_rca32_fa706_y4;
  assign f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa705_y4 = f_s_dadda_pg_rca32_fa705_y4;
  assign f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa131_y2 = f_s_dadda_pg_rca32_fa131_y2;
  assign f_s_dadda_pg_rca32_fa707_y0 = f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa706_y4 ^ f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa705_y4;
  assign f_s_dadda_pg_rca32_fa707_y1 = f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa706_y4 & f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa705_y4;
  assign f_s_dadda_pg_rca32_fa707_y2 = f_s_dadda_pg_rca32_fa707_y0 ^ f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa131_y2;
  assign f_s_dadda_pg_rca32_fa707_y3 = f_s_dadda_pg_rca32_fa707_y0 & f_s_dadda_pg_rca32_fa707_f_s_dadda_pg_rca32_fa131_y2;
  assign f_s_dadda_pg_rca32_fa707_y4 = f_s_dadda_pg_rca32_fa707_y1 | f_s_dadda_pg_rca32_fa707_y3;
  assign f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa132_y2 = f_s_dadda_pg_rca32_fa132_y2;
  assign f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa133_y2 = f_s_dadda_pg_rca32_fa133_y2;
  assign f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa134_y2 = f_s_dadda_pg_rca32_fa134_y2;
  assign f_s_dadda_pg_rca32_fa708_y0 = f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa132_y2 ^ f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa133_y2;
  assign f_s_dadda_pg_rca32_fa708_y1 = f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa132_y2 & f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa133_y2;
  assign f_s_dadda_pg_rca32_fa708_y2 = f_s_dadda_pg_rca32_fa708_y0 ^ f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa134_y2;
  assign f_s_dadda_pg_rca32_fa708_y3 = f_s_dadda_pg_rca32_fa708_y0 & f_s_dadda_pg_rca32_fa708_f_s_dadda_pg_rca32_fa134_y2;
  assign f_s_dadda_pg_rca32_fa708_y4 = f_s_dadda_pg_rca32_fa708_y1 | f_s_dadda_pg_rca32_fa708_y3;
  assign f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa708_y4 = f_s_dadda_pg_rca32_fa708_y4;
  assign f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa707_y4 = f_s_dadda_pg_rca32_fa707_y4;
  assign f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa147_y2 = f_s_dadda_pg_rca32_fa147_y2;
  assign f_s_dadda_pg_rca32_fa709_y0 = f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa708_y4 ^ f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa707_y4;
  assign f_s_dadda_pg_rca32_fa709_y1 = f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa708_y4 & f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa707_y4;
  assign f_s_dadda_pg_rca32_fa709_y2 = f_s_dadda_pg_rca32_fa709_y0 ^ f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa147_y2;
  assign f_s_dadda_pg_rca32_fa709_y3 = f_s_dadda_pg_rca32_fa709_y0 & f_s_dadda_pg_rca32_fa709_f_s_dadda_pg_rca32_fa147_y2;
  assign f_s_dadda_pg_rca32_fa709_y4 = f_s_dadda_pg_rca32_fa709_y1 | f_s_dadda_pg_rca32_fa709_y3;
  assign f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa148_y2 = f_s_dadda_pg_rca32_fa148_y2;
  assign f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa149_y2 = f_s_dadda_pg_rca32_fa149_y2;
  assign f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa150_y2 = f_s_dadda_pg_rca32_fa150_y2;
  assign f_s_dadda_pg_rca32_fa710_y0 = f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa148_y2 ^ f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa149_y2;
  assign f_s_dadda_pg_rca32_fa710_y1 = f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa148_y2 & f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa149_y2;
  assign f_s_dadda_pg_rca32_fa710_y2 = f_s_dadda_pg_rca32_fa710_y0 ^ f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa150_y2;
  assign f_s_dadda_pg_rca32_fa710_y3 = f_s_dadda_pg_rca32_fa710_y0 & f_s_dadda_pg_rca32_fa710_f_s_dadda_pg_rca32_fa150_y2;
  assign f_s_dadda_pg_rca32_fa710_y4 = f_s_dadda_pg_rca32_fa710_y1 | f_s_dadda_pg_rca32_fa710_y3;
  assign f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa710_y4 = f_s_dadda_pg_rca32_fa710_y4;
  assign f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa709_y4 = f_s_dadda_pg_rca32_fa709_y4;
  assign f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa164_y2 = f_s_dadda_pg_rca32_fa164_y2;
  assign f_s_dadda_pg_rca32_fa711_y0 = f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa710_y4 ^ f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa709_y4;
  assign f_s_dadda_pg_rca32_fa711_y1 = f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa710_y4 & f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa709_y4;
  assign f_s_dadda_pg_rca32_fa711_y2 = f_s_dadda_pg_rca32_fa711_y0 ^ f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa164_y2;
  assign f_s_dadda_pg_rca32_fa711_y3 = f_s_dadda_pg_rca32_fa711_y0 & f_s_dadda_pg_rca32_fa711_f_s_dadda_pg_rca32_fa164_y2;
  assign f_s_dadda_pg_rca32_fa711_y4 = f_s_dadda_pg_rca32_fa711_y1 | f_s_dadda_pg_rca32_fa711_y3;
  assign f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa165_y2 = f_s_dadda_pg_rca32_fa165_y2;
  assign f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa166_y2 = f_s_dadda_pg_rca32_fa166_y2;
  assign f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa167_y2 = f_s_dadda_pg_rca32_fa167_y2;
  assign f_s_dadda_pg_rca32_fa712_y0 = f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa165_y2 ^ f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa166_y2;
  assign f_s_dadda_pg_rca32_fa712_y1 = f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa165_y2 & f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa166_y2;
  assign f_s_dadda_pg_rca32_fa712_y2 = f_s_dadda_pg_rca32_fa712_y0 ^ f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa167_y2;
  assign f_s_dadda_pg_rca32_fa712_y3 = f_s_dadda_pg_rca32_fa712_y0 & f_s_dadda_pg_rca32_fa712_f_s_dadda_pg_rca32_fa167_y2;
  assign f_s_dadda_pg_rca32_fa712_y4 = f_s_dadda_pg_rca32_fa712_y1 | f_s_dadda_pg_rca32_fa712_y3;
  assign f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa712_y4 = f_s_dadda_pg_rca32_fa712_y4;
  assign f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa711_y4 = f_s_dadda_pg_rca32_fa711_y4;
  assign f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa182_y2 = f_s_dadda_pg_rca32_fa182_y2;
  assign f_s_dadda_pg_rca32_fa713_y0 = f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa712_y4 ^ f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa711_y4;
  assign f_s_dadda_pg_rca32_fa713_y1 = f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa712_y4 & f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa711_y4;
  assign f_s_dadda_pg_rca32_fa713_y2 = f_s_dadda_pg_rca32_fa713_y0 ^ f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa182_y2;
  assign f_s_dadda_pg_rca32_fa713_y3 = f_s_dadda_pg_rca32_fa713_y0 & f_s_dadda_pg_rca32_fa713_f_s_dadda_pg_rca32_fa182_y2;
  assign f_s_dadda_pg_rca32_fa713_y4 = f_s_dadda_pg_rca32_fa713_y1 | f_s_dadda_pg_rca32_fa713_y3;
  assign f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa183_y2 = f_s_dadda_pg_rca32_fa183_y2;
  assign f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa184_y2 = f_s_dadda_pg_rca32_fa184_y2;
  assign f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa185_y2 = f_s_dadda_pg_rca32_fa185_y2;
  assign f_s_dadda_pg_rca32_fa714_y0 = f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa183_y2 ^ f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa184_y2;
  assign f_s_dadda_pg_rca32_fa714_y1 = f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa183_y2 & f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa184_y2;
  assign f_s_dadda_pg_rca32_fa714_y2 = f_s_dadda_pg_rca32_fa714_y0 ^ f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa185_y2;
  assign f_s_dadda_pg_rca32_fa714_y3 = f_s_dadda_pg_rca32_fa714_y0 & f_s_dadda_pg_rca32_fa714_f_s_dadda_pg_rca32_fa185_y2;
  assign f_s_dadda_pg_rca32_fa714_y4 = f_s_dadda_pg_rca32_fa714_y1 | f_s_dadda_pg_rca32_fa714_y3;
  assign f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa714_y4 = f_s_dadda_pg_rca32_fa714_y4;
  assign f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa713_y4 = f_s_dadda_pg_rca32_fa713_y4;
  assign f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa201_y2 = f_s_dadda_pg_rca32_fa201_y2;
  assign f_s_dadda_pg_rca32_fa715_y0 = f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa714_y4 ^ f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa713_y4;
  assign f_s_dadda_pg_rca32_fa715_y1 = f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa714_y4 & f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa713_y4;
  assign f_s_dadda_pg_rca32_fa715_y2 = f_s_dadda_pg_rca32_fa715_y0 ^ f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa201_y2;
  assign f_s_dadda_pg_rca32_fa715_y3 = f_s_dadda_pg_rca32_fa715_y0 & f_s_dadda_pg_rca32_fa715_f_s_dadda_pg_rca32_fa201_y2;
  assign f_s_dadda_pg_rca32_fa715_y4 = f_s_dadda_pg_rca32_fa715_y1 | f_s_dadda_pg_rca32_fa715_y3;
  assign f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa202_y2 = f_s_dadda_pg_rca32_fa202_y2;
  assign f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa203_y2 = f_s_dadda_pg_rca32_fa203_y2;
  assign f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa204_y2 = f_s_dadda_pg_rca32_fa204_y2;
  assign f_s_dadda_pg_rca32_fa716_y0 = f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa202_y2 ^ f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa203_y2;
  assign f_s_dadda_pg_rca32_fa716_y1 = f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa202_y2 & f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa203_y2;
  assign f_s_dadda_pg_rca32_fa716_y2 = f_s_dadda_pg_rca32_fa716_y0 ^ f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa204_y2;
  assign f_s_dadda_pg_rca32_fa716_y3 = f_s_dadda_pg_rca32_fa716_y0 & f_s_dadda_pg_rca32_fa716_f_s_dadda_pg_rca32_fa204_y2;
  assign f_s_dadda_pg_rca32_fa716_y4 = f_s_dadda_pg_rca32_fa716_y1 | f_s_dadda_pg_rca32_fa716_y3;
  assign f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa716_y4 = f_s_dadda_pg_rca32_fa716_y4;
  assign f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa715_y4 = f_s_dadda_pg_rca32_fa715_y4;
  assign f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa221_y2 = f_s_dadda_pg_rca32_fa221_y2;
  assign f_s_dadda_pg_rca32_fa717_y0 = f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa716_y4 ^ f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa715_y4;
  assign f_s_dadda_pg_rca32_fa717_y1 = f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa716_y4 & f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa715_y4;
  assign f_s_dadda_pg_rca32_fa717_y2 = f_s_dadda_pg_rca32_fa717_y0 ^ f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa221_y2;
  assign f_s_dadda_pg_rca32_fa717_y3 = f_s_dadda_pg_rca32_fa717_y0 & f_s_dadda_pg_rca32_fa717_f_s_dadda_pg_rca32_fa221_y2;
  assign f_s_dadda_pg_rca32_fa717_y4 = f_s_dadda_pg_rca32_fa717_y1 | f_s_dadda_pg_rca32_fa717_y3;
  assign f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa222_y2 = f_s_dadda_pg_rca32_fa222_y2;
  assign f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa223_y2 = f_s_dadda_pg_rca32_fa223_y2;
  assign f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa224_y2 = f_s_dadda_pg_rca32_fa224_y2;
  assign f_s_dadda_pg_rca32_fa718_y0 = f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa222_y2 ^ f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa223_y2;
  assign f_s_dadda_pg_rca32_fa718_y1 = f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa222_y2 & f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa223_y2;
  assign f_s_dadda_pg_rca32_fa718_y2 = f_s_dadda_pg_rca32_fa718_y0 ^ f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa224_y2;
  assign f_s_dadda_pg_rca32_fa718_y3 = f_s_dadda_pg_rca32_fa718_y0 & f_s_dadda_pg_rca32_fa718_f_s_dadda_pg_rca32_fa224_y2;
  assign f_s_dadda_pg_rca32_fa718_y4 = f_s_dadda_pg_rca32_fa718_y1 | f_s_dadda_pg_rca32_fa718_y3;
  assign f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa718_y4 = f_s_dadda_pg_rca32_fa718_y4;
  assign f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa717_y4 = f_s_dadda_pg_rca32_fa717_y4;
  assign f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa242_y2 = f_s_dadda_pg_rca32_fa242_y2;
  assign f_s_dadda_pg_rca32_fa719_y0 = f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa718_y4 ^ f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa717_y4;
  assign f_s_dadda_pg_rca32_fa719_y1 = f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa718_y4 & f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa717_y4;
  assign f_s_dadda_pg_rca32_fa719_y2 = f_s_dadda_pg_rca32_fa719_y0 ^ f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa242_y2;
  assign f_s_dadda_pg_rca32_fa719_y3 = f_s_dadda_pg_rca32_fa719_y0 & f_s_dadda_pg_rca32_fa719_f_s_dadda_pg_rca32_fa242_y2;
  assign f_s_dadda_pg_rca32_fa719_y4 = f_s_dadda_pg_rca32_fa719_y1 | f_s_dadda_pg_rca32_fa719_y3;
  assign f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa243_y2 = f_s_dadda_pg_rca32_fa243_y2;
  assign f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa244_y2 = f_s_dadda_pg_rca32_fa244_y2;
  assign f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa245_y2 = f_s_dadda_pg_rca32_fa245_y2;
  assign f_s_dadda_pg_rca32_fa720_y0 = f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa243_y2 ^ f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa244_y2;
  assign f_s_dadda_pg_rca32_fa720_y1 = f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa243_y2 & f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa244_y2;
  assign f_s_dadda_pg_rca32_fa720_y2 = f_s_dadda_pg_rca32_fa720_y0 ^ f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa245_y2;
  assign f_s_dadda_pg_rca32_fa720_y3 = f_s_dadda_pg_rca32_fa720_y0 & f_s_dadda_pg_rca32_fa720_f_s_dadda_pg_rca32_fa245_y2;
  assign f_s_dadda_pg_rca32_fa720_y4 = f_s_dadda_pg_rca32_fa720_y1 | f_s_dadda_pg_rca32_fa720_y3;
  assign f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa720_y4 = f_s_dadda_pg_rca32_fa720_y4;
  assign f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa719_y4 = f_s_dadda_pg_rca32_fa719_y4;
  assign f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa263_y2 = f_s_dadda_pg_rca32_fa263_y2;
  assign f_s_dadda_pg_rca32_fa721_y0 = f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa720_y4 ^ f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa719_y4;
  assign f_s_dadda_pg_rca32_fa721_y1 = f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa720_y4 & f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa719_y4;
  assign f_s_dadda_pg_rca32_fa721_y2 = f_s_dadda_pg_rca32_fa721_y0 ^ f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa263_y2;
  assign f_s_dadda_pg_rca32_fa721_y3 = f_s_dadda_pg_rca32_fa721_y0 & f_s_dadda_pg_rca32_fa721_f_s_dadda_pg_rca32_fa263_y2;
  assign f_s_dadda_pg_rca32_fa721_y4 = f_s_dadda_pg_rca32_fa721_y1 | f_s_dadda_pg_rca32_fa721_y3;
  assign f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa264_y2 = f_s_dadda_pg_rca32_fa264_y2;
  assign f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa265_y2 = f_s_dadda_pg_rca32_fa265_y2;
  assign f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa266_y2 = f_s_dadda_pg_rca32_fa266_y2;
  assign f_s_dadda_pg_rca32_fa722_y0 = f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa264_y2 ^ f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa265_y2;
  assign f_s_dadda_pg_rca32_fa722_y1 = f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa264_y2 & f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa265_y2;
  assign f_s_dadda_pg_rca32_fa722_y2 = f_s_dadda_pg_rca32_fa722_y0 ^ f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa266_y2;
  assign f_s_dadda_pg_rca32_fa722_y3 = f_s_dadda_pg_rca32_fa722_y0 & f_s_dadda_pg_rca32_fa722_f_s_dadda_pg_rca32_fa266_y2;
  assign f_s_dadda_pg_rca32_fa722_y4 = f_s_dadda_pg_rca32_fa722_y1 | f_s_dadda_pg_rca32_fa722_y3;
  assign f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa722_y4 = f_s_dadda_pg_rca32_fa722_y4;
  assign f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa721_y4 = f_s_dadda_pg_rca32_fa721_y4;
  assign f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa285_y2 = f_s_dadda_pg_rca32_fa285_y2;
  assign f_s_dadda_pg_rca32_fa723_y0 = f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa722_y4 ^ f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa721_y4;
  assign f_s_dadda_pg_rca32_fa723_y1 = f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa722_y4 & f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa721_y4;
  assign f_s_dadda_pg_rca32_fa723_y2 = f_s_dadda_pg_rca32_fa723_y0 ^ f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa285_y2;
  assign f_s_dadda_pg_rca32_fa723_y3 = f_s_dadda_pg_rca32_fa723_y0 & f_s_dadda_pg_rca32_fa723_f_s_dadda_pg_rca32_fa285_y2;
  assign f_s_dadda_pg_rca32_fa723_y4 = f_s_dadda_pg_rca32_fa723_y1 | f_s_dadda_pg_rca32_fa723_y3;
  assign f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa286_y2 = f_s_dadda_pg_rca32_fa286_y2;
  assign f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa287_y2 = f_s_dadda_pg_rca32_fa287_y2;
  assign f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa288_y2 = f_s_dadda_pg_rca32_fa288_y2;
  assign f_s_dadda_pg_rca32_fa724_y0 = f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa286_y2 ^ f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa287_y2;
  assign f_s_dadda_pg_rca32_fa724_y1 = f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa286_y2 & f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa287_y2;
  assign f_s_dadda_pg_rca32_fa724_y2 = f_s_dadda_pg_rca32_fa724_y0 ^ f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa288_y2;
  assign f_s_dadda_pg_rca32_fa724_y3 = f_s_dadda_pg_rca32_fa724_y0 & f_s_dadda_pg_rca32_fa724_f_s_dadda_pg_rca32_fa288_y2;
  assign f_s_dadda_pg_rca32_fa724_y4 = f_s_dadda_pg_rca32_fa724_y1 | f_s_dadda_pg_rca32_fa724_y3;
  assign f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa724_y4 = f_s_dadda_pg_rca32_fa724_y4;
  assign f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa723_y4 = f_s_dadda_pg_rca32_fa723_y4;
  assign f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa307_y2 = f_s_dadda_pg_rca32_fa307_y2;
  assign f_s_dadda_pg_rca32_fa725_y0 = f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa724_y4 ^ f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa723_y4;
  assign f_s_dadda_pg_rca32_fa725_y1 = f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa724_y4 & f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa723_y4;
  assign f_s_dadda_pg_rca32_fa725_y2 = f_s_dadda_pg_rca32_fa725_y0 ^ f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa307_y2;
  assign f_s_dadda_pg_rca32_fa725_y3 = f_s_dadda_pg_rca32_fa725_y0 & f_s_dadda_pg_rca32_fa725_f_s_dadda_pg_rca32_fa307_y2;
  assign f_s_dadda_pg_rca32_fa725_y4 = f_s_dadda_pg_rca32_fa725_y1 | f_s_dadda_pg_rca32_fa725_y3;
  assign f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa308_y2 = f_s_dadda_pg_rca32_fa308_y2;
  assign f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa309_y2 = f_s_dadda_pg_rca32_fa309_y2;
  assign f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa310_y2 = f_s_dadda_pg_rca32_fa310_y2;
  assign f_s_dadda_pg_rca32_fa726_y0 = f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa308_y2 ^ f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa309_y2;
  assign f_s_dadda_pg_rca32_fa726_y1 = f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa308_y2 & f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa309_y2;
  assign f_s_dadda_pg_rca32_fa726_y2 = f_s_dadda_pg_rca32_fa726_y0 ^ f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa310_y2;
  assign f_s_dadda_pg_rca32_fa726_y3 = f_s_dadda_pg_rca32_fa726_y0 & f_s_dadda_pg_rca32_fa726_f_s_dadda_pg_rca32_fa310_y2;
  assign f_s_dadda_pg_rca32_fa726_y4 = f_s_dadda_pg_rca32_fa726_y1 | f_s_dadda_pg_rca32_fa726_y3;
  assign f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa726_y4 = f_s_dadda_pg_rca32_fa726_y4;
  assign f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa725_y4 = f_s_dadda_pg_rca32_fa725_y4;
  assign f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa329_y2 = f_s_dadda_pg_rca32_fa329_y2;
  assign f_s_dadda_pg_rca32_fa727_y0 = f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa726_y4 ^ f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa725_y4;
  assign f_s_dadda_pg_rca32_fa727_y1 = f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa726_y4 & f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa725_y4;
  assign f_s_dadda_pg_rca32_fa727_y2 = f_s_dadda_pg_rca32_fa727_y0 ^ f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa329_y2;
  assign f_s_dadda_pg_rca32_fa727_y3 = f_s_dadda_pg_rca32_fa727_y0 & f_s_dadda_pg_rca32_fa727_f_s_dadda_pg_rca32_fa329_y2;
  assign f_s_dadda_pg_rca32_fa727_y4 = f_s_dadda_pg_rca32_fa727_y1 | f_s_dadda_pg_rca32_fa727_y3;
  assign f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa330_y2 = f_s_dadda_pg_rca32_fa330_y2;
  assign f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa331_y2 = f_s_dadda_pg_rca32_fa331_y2;
  assign f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa332_y2 = f_s_dadda_pg_rca32_fa332_y2;
  assign f_s_dadda_pg_rca32_fa728_y0 = f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa330_y2 ^ f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa331_y2;
  assign f_s_dadda_pg_rca32_fa728_y1 = f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa330_y2 & f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa331_y2;
  assign f_s_dadda_pg_rca32_fa728_y2 = f_s_dadda_pg_rca32_fa728_y0 ^ f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa332_y2;
  assign f_s_dadda_pg_rca32_fa728_y3 = f_s_dadda_pg_rca32_fa728_y0 & f_s_dadda_pg_rca32_fa728_f_s_dadda_pg_rca32_fa332_y2;
  assign f_s_dadda_pg_rca32_fa728_y4 = f_s_dadda_pg_rca32_fa728_y1 | f_s_dadda_pg_rca32_fa728_y3;
  assign f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa728_y4 = f_s_dadda_pg_rca32_fa728_y4;
  assign f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa727_y4 = f_s_dadda_pg_rca32_fa727_y4;
  assign f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa351_y2 = f_s_dadda_pg_rca32_fa351_y2;
  assign f_s_dadda_pg_rca32_fa729_y0 = f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa728_y4 ^ f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa727_y4;
  assign f_s_dadda_pg_rca32_fa729_y1 = f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa728_y4 & f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa727_y4;
  assign f_s_dadda_pg_rca32_fa729_y2 = f_s_dadda_pg_rca32_fa729_y0 ^ f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa351_y2;
  assign f_s_dadda_pg_rca32_fa729_y3 = f_s_dadda_pg_rca32_fa729_y0 & f_s_dadda_pg_rca32_fa729_f_s_dadda_pg_rca32_fa351_y2;
  assign f_s_dadda_pg_rca32_fa729_y4 = f_s_dadda_pg_rca32_fa729_y1 | f_s_dadda_pg_rca32_fa729_y3;
  assign f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa352_y2 = f_s_dadda_pg_rca32_fa352_y2;
  assign f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa353_y2 = f_s_dadda_pg_rca32_fa353_y2;
  assign f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa354_y2 = f_s_dadda_pg_rca32_fa354_y2;
  assign f_s_dadda_pg_rca32_fa730_y0 = f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa352_y2 ^ f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa353_y2;
  assign f_s_dadda_pg_rca32_fa730_y1 = f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa352_y2 & f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa353_y2;
  assign f_s_dadda_pg_rca32_fa730_y2 = f_s_dadda_pg_rca32_fa730_y0 ^ f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa354_y2;
  assign f_s_dadda_pg_rca32_fa730_y3 = f_s_dadda_pg_rca32_fa730_y0 & f_s_dadda_pg_rca32_fa730_f_s_dadda_pg_rca32_fa354_y2;
  assign f_s_dadda_pg_rca32_fa730_y4 = f_s_dadda_pg_rca32_fa730_y1 | f_s_dadda_pg_rca32_fa730_y3;
  assign f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa730_y4 = f_s_dadda_pg_rca32_fa730_y4;
  assign f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa729_y4 = f_s_dadda_pg_rca32_fa729_y4;
  assign f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa373_y2 = f_s_dadda_pg_rca32_fa373_y2;
  assign f_s_dadda_pg_rca32_fa731_y0 = f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa730_y4 ^ f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa729_y4;
  assign f_s_dadda_pg_rca32_fa731_y1 = f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa730_y4 & f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa729_y4;
  assign f_s_dadda_pg_rca32_fa731_y2 = f_s_dadda_pg_rca32_fa731_y0 ^ f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa373_y2;
  assign f_s_dadda_pg_rca32_fa731_y3 = f_s_dadda_pg_rca32_fa731_y0 & f_s_dadda_pg_rca32_fa731_f_s_dadda_pg_rca32_fa373_y2;
  assign f_s_dadda_pg_rca32_fa731_y4 = f_s_dadda_pg_rca32_fa731_y1 | f_s_dadda_pg_rca32_fa731_y3;
  assign f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa374_y2 = f_s_dadda_pg_rca32_fa374_y2;
  assign f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa375_y2 = f_s_dadda_pg_rca32_fa375_y2;
  assign f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa376_y2 = f_s_dadda_pg_rca32_fa376_y2;
  assign f_s_dadda_pg_rca32_fa732_y0 = f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa374_y2 ^ f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa375_y2;
  assign f_s_dadda_pg_rca32_fa732_y1 = f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa374_y2 & f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa375_y2;
  assign f_s_dadda_pg_rca32_fa732_y2 = f_s_dadda_pg_rca32_fa732_y0 ^ f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa376_y2;
  assign f_s_dadda_pg_rca32_fa732_y3 = f_s_dadda_pg_rca32_fa732_y0 & f_s_dadda_pg_rca32_fa732_f_s_dadda_pg_rca32_fa376_y2;
  assign f_s_dadda_pg_rca32_fa732_y4 = f_s_dadda_pg_rca32_fa732_y1 | f_s_dadda_pg_rca32_fa732_y3;
  assign f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa732_y4 = f_s_dadda_pg_rca32_fa732_y4;
  assign f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa731_y4 = f_s_dadda_pg_rca32_fa731_y4;
  assign f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa395_y2 = f_s_dadda_pg_rca32_fa395_y2;
  assign f_s_dadda_pg_rca32_fa733_y0 = f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa732_y4 ^ f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa731_y4;
  assign f_s_dadda_pg_rca32_fa733_y1 = f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa732_y4 & f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa731_y4;
  assign f_s_dadda_pg_rca32_fa733_y2 = f_s_dadda_pg_rca32_fa733_y0 ^ f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa395_y2;
  assign f_s_dadda_pg_rca32_fa733_y3 = f_s_dadda_pg_rca32_fa733_y0 & f_s_dadda_pg_rca32_fa733_f_s_dadda_pg_rca32_fa395_y2;
  assign f_s_dadda_pg_rca32_fa733_y4 = f_s_dadda_pg_rca32_fa733_y1 | f_s_dadda_pg_rca32_fa733_y3;
  assign f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa396_y2 = f_s_dadda_pg_rca32_fa396_y2;
  assign f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa397_y2 = f_s_dadda_pg_rca32_fa397_y2;
  assign f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa398_y2 = f_s_dadda_pg_rca32_fa398_y2;
  assign f_s_dadda_pg_rca32_fa734_y0 = f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa396_y2 ^ f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa397_y2;
  assign f_s_dadda_pg_rca32_fa734_y1 = f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa396_y2 & f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa397_y2;
  assign f_s_dadda_pg_rca32_fa734_y2 = f_s_dadda_pg_rca32_fa734_y0 ^ f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa398_y2;
  assign f_s_dadda_pg_rca32_fa734_y3 = f_s_dadda_pg_rca32_fa734_y0 & f_s_dadda_pg_rca32_fa734_f_s_dadda_pg_rca32_fa398_y2;
  assign f_s_dadda_pg_rca32_fa734_y4 = f_s_dadda_pg_rca32_fa734_y1 | f_s_dadda_pg_rca32_fa734_y3;
  assign f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa734_y4 = f_s_dadda_pg_rca32_fa734_y4;
  assign f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa733_y4 = f_s_dadda_pg_rca32_fa733_y4;
  assign f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa417_y2 = f_s_dadda_pg_rca32_fa417_y2;
  assign f_s_dadda_pg_rca32_fa735_y0 = f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa734_y4 ^ f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa733_y4;
  assign f_s_dadda_pg_rca32_fa735_y1 = f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa734_y4 & f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa733_y4;
  assign f_s_dadda_pg_rca32_fa735_y2 = f_s_dadda_pg_rca32_fa735_y0 ^ f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa417_y2;
  assign f_s_dadda_pg_rca32_fa735_y3 = f_s_dadda_pg_rca32_fa735_y0 & f_s_dadda_pg_rca32_fa735_f_s_dadda_pg_rca32_fa417_y2;
  assign f_s_dadda_pg_rca32_fa735_y4 = f_s_dadda_pg_rca32_fa735_y1 | f_s_dadda_pg_rca32_fa735_y3;
  assign f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa418_y2 = f_s_dadda_pg_rca32_fa418_y2;
  assign f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa419_y2 = f_s_dadda_pg_rca32_fa419_y2;
  assign f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa420_y2 = f_s_dadda_pg_rca32_fa420_y2;
  assign f_s_dadda_pg_rca32_fa736_y0 = f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa418_y2 ^ f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa419_y2;
  assign f_s_dadda_pg_rca32_fa736_y1 = f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa418_y2 & f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa419_y2;
  assign f_s_dadda_pg_rca32_fa736_y2 = f_s_dadda_pg_rca32_fa736_y0 ^ f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa420_y2;
  assign f_s_dadda_pg_rca32_fa736_y3 = f_s_dadda_pg_rca32_fa736_y0 & f_s_dadda_pg_rca32_fa736_f_s_dadda_pg_rca32_fa420_y2;
  assign f_s_dadda_pg_rca32_fa736_y4 = f_s_dadda_pg_rca32_fa736_y1 | f_s_dadda_pg_rca32_fa736_y3;
  assign f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa736_y4 = f_s_dadda_pg_rca32_fa736_y4;
  assign f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa735_y4 = f_s_dadda_pg_rca32_fa735_y4;
  assign f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa439_y2 = f_s_dadda_pg_rca32_fa439_y2;
  assign f_s_dadda_pg_rca32_fa737_y0 = f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa736_y4 ^ f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa735_y4;
  assign f_s_dadda_pg_rca32_fa737_y1 = f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa736_y4 & f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa735_y4;
  assign f_s_dadda_pg_rca32_fa737_y2 = f_s_dadda_pg_rca32_fa737_y0 ^ f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa439_y2;
  assign f_s_dadda_pg_rca32_fa737_y3 = f_s_dadda_pg_rca32_fa737_y0 & f_s_dadda_pg_rca32_fa737_f_s_dadda_pg_rca32_fa439_y2;
  assign f_s_dadda_pg_rca32_fa737_y4 = f_s_dadda_pg_rca32_fa737_y1 | f_s_dadda_pg_rca32_fa737_y3;
  assign f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa440_y2 = f_s_dadda_pg_rca32_fa440_y2;
  assign f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa441_y2 = f_s_dadda_pg_rca32_fa441_y2;
  assign f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa442_y2 = f_s_dadda_pg_rca32_fa442_y2;
  assign f_s_dadda_pg_rca32_fa738_y0 = f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa440_y2 ^ f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa441_y2;
  assign f_s_dadda_pg_rca32_fa738_y1 = f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa440_y2 & f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa441_y2;
  assign f_s_dadda_pg_rca32_fa738_y2 = f_s_dadda_pg_rca32_fa738_y0 ^ f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa442_y2;
  assign f_s_dadda_pg_rca32_fa738_y3 = f_s_dadda_pg_rca32_fa738_y0 & f_s_dadda_pg_rca32_fa738_f_s_dadda_pg_rca32_fa442_y2;
  assign f_s_dadda_pg_rca32_fa738_y4 = f_s_dadda_pg_rca32_fa738_y1 | f_s_dadda_pg_rca32_fa738_y3;
  assign f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa738_y4 = f_s_dadda_pg_rca32_fa738_y4;
  assign f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa737_y4 = f_s_dadda_pg_rca32_fa737_y4;
  assign f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa460_y2 = f_s_dadda_pg_rca32_fa460_y2;
  assign f_s_dadda_pg_rca32_fa739_y0 = f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa738_y4 ^ f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa737_y4;
  assign f_s_dadda_pg_rca32_fa739_y1 = f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa738_y4 & f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa737_y4;
  assign f_s_dadda_pg_rca32_fa739_y2 = f_s_dadda_pg_rca32_fa739_y0 ^ f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa460_y2;
  assign f_s_dadda_pg_rca32_fa739_y3 = f_s_dadda_pg_rca32_fa739_y0 & f_s_dadda_pg_rca32_fa739_f_s_dadda_pg_rca32_fa460_y2;
  assign f_s_dadda_pg_rca32_fa739_y4 = f_s_dadda_pg_rca32_fa739_y1 | f_s_dadda_pg_rca32_fa739_y3;
  assign f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa461_y2 = f_s_dadda_pg_rca32_fa461_y2;
  assign f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa462_y2 = f_s_dadda_pg_rca32_fa462_y2;
  assign f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa463_y2 = f_s_dadda_pg_rca32_fa463_y2;
  assign f_s_dadda_pg_rca32_fa740_y0 = f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa461_y2 ^ f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa462_y2;
  assign f_s_dadda_pg_rca32_fa740_y1 = f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa461_y2 & f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa462_y2;
  assign f_s_dadda_pg_rca32_fa740_y2 = f_s_dadda_pg_rca32_fa740_y0 ^ f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa463_y2;
  assign f_s_dadda_pg_rca32_fa740_y3 = f_s_dadda_pg_rca32_fa740_y0 & f_s_dadda_pg_rca32_fa740_f_s_dadda_pg_rca32_fa463_y2;
  assign f_s_dadda_pg_rca32_fa740_y4 = f_s_dadda_pg_rca32_fa740_y1 | f_s_dadda_pg_rca32_fa740_y3;
  assign f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa740_y4 = f_s_dadda_pg_rca32_fa740_y4;
  assign f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa739_y4 = f_s_dadda_pg_rca32_fa739_y4;
  assign f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa480_y2 = f_s_dadda_pg_rca32_fa480_y2;
  assign f_s_dadda_pg_rca32_fa741_y0 = f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa740_y4 ^ f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa739_y4;
  assign f_s_dadda_pg_rca32_fa741_y1 = f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa740_y4 & f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa739_y4;
  assign f_s_dadda_pg_rca32_fa741_y2 = f_s_dadda_pg_rca32_fa741_y0 ^ f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa480_y2;
  assign f_s_dadda_pg_rca32_fa741_y3 = f_s_dadda_pg_rca32_fa741_y0 & f_s_dadda_pg_rca32_fa741_f_s_dadda_pg_rca32_fa480_y2;
  assign f_s_dadda_pg_rca32_fa741_y4 = f_s_dadda_pg_rca32_fa741_y1 | f_s_dadda_pg_rca32_fa741_y3;
  assign f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa481_y2 = f_s_dadda_pg_rca32_fa481_y2;
  assign f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa482_y2 = f_s_dadda_pg_rca32_fa482_y2;
  assign f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa483_y2 = f_s_dadda_pg_rca32_fa483_y2;
  assign f_s_dadda_pg_rca32_fa742_y0 = f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa481_y2 ^ f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa482_y2;
  assign f_s_dadda_pg_rca32_fa742_y1 = f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa481_y2 & f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa482_y2;
  assign f_s_dadda_pg_rca32_fa742_y2 = f_s_dadda_pg_rca32_fa742_y0 ^ f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa483_y2;
  assign f_s_dadda_pg_rca32_fa742_y3 = f_s_dadda_pg_rca32_fa742_y0 & f_s_dadda_pg_rca32_fa742_f_s_dadda_pg_rca32_fa483_y2;
  assign f_s_dadda_pg_rca32_fa742_y4 = f_s_dadda_pg_rca32_fa742_y1 | f_s_dadda_pg_rca32_fa742_y3;
  assign f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa742_y4 = f_s_dadda_pg_rca32_fa742_y4;
  assign f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa741_y4 = f_s_dadda_pg_rca32_fa741_y4;
  assign f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa499_y2 = f_s_dadda_pg_rca32_fa499_y2;
  assign f_s_dadda_pg_rca32_fa743_y0 = f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa742_y4 ^ f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa741_y4;
  assign f_s_dadda_pg_rca32_fa743_y1 = f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa742_y4 & f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa741_y4;
  assign f_s_dadda_pg_rca32_fa743_y2 = f_s_dadda_pg_rca32_fa743_y0 ^ f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa499_y2;
  assign f_s_dadda_pg_rca32_fa743_y3 = f_s_dadda_pg_rca32_fa743_y0 & f_s_dadda_pg_rca32_fa743_f_s_dadda_pg_rca32_fa499_y2;
  assign f_s_dadda_pg_rca32_fa743_y4 = f_s_dadda_pg_rca32_fa743_y1 | f_s_dadda_pg_rca32_fa743_y3;
  assign f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa500_y2 = f_s_dadda_pg_rca32_fa500_y2;
  assign f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa501_y2 = f_s_dadda_pg_rca32_fa501_y2;
  assign f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa502_y2 = f_s_dadda_pg_rca32_fa502_y2;
  assign f_s_dadda_pg_rca32_fa744_y0 = f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa500_y2 ^ f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa501_y2;
  assign f_s_dadda_pg_rca32_fa744_y1 = f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa500_y2 & f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa501_y2;
  assign f_s_dadda_pg_rca32_fa744_y2 = f_s_dadda_pg_rca32_fa744_y0 ^ f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa502_y2;
  assign f_s_dadda_pg_rca32_fa744_y3 = f_s_dadda_pg_rca32_fa744_y0 & f_s_dadda_pg_rca32_fa744_f_s_dadda_pg_rca32_fa502_y2;
  assign f_s_dadda_pg_rca32_fa744_y4 = f_s_dadda_pg_rca32_fa744_y1 | f_s_dadda_pg_rca32_fa744_y3;
  assign f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa744_y4 = f_s_dadda_pg_rca32_fa744_y4;
  assign f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa743_y4 = f_s_dadda_pg_rca32_fa743_y4;
  assign f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa517_y2 = f_s_dadda_pg_rca32_fa517_y2;
  assign f_s_dadda_pg_rca32_fa745_y0 = f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa744_y4 ^ f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa743_y4;
  assign f_s_dadda_pg_rca32_fa745_y1 = f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa744_y4 & f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa743_y4;
  assign f_s_dadda_pg_rca32_fa745_y2 = f_s_dadda_pg_rca32_fa745_y0 ^ f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa517_y2;
  assign f_s_dadda_pg_rca32_fa745_y3 = f_s_dadda_pg_rca32_fa745_y0 & f_s_dadda_pg_rca32_fa745_f_s_dadda_pg_rca32_fa517_y2;
  assign f_s_dadda_pg_rca32_fa745_y4 = f_s_dadda_pg_rca32_fa745_y1 | f_s_dadda_pg_rca32_fa745_y3;
  assign f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa518_y2 = f_s_dadda_pg_rca32_fa518_y2;
  assign f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa519_y2 = f_s_dadda_pg_rca32_fa519_y2;
  assign f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa520_y2 = f_s_dadda_pg_rca32_fa520_y2;
  assign f_s_dadda_pg_rca32_fa746_y0 = f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa518_y2 ^ f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa519_y2;
  assign f_s_dadda_pg_rca32_fa746_y1 = f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa518_y2 & f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa519_y2;
  assign f_s_dadda_pg_rca32_fa746_y2 = f_s_dadda_pg_rca32_fa746_y0 ^ f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa520_y2;
  assign f_s_dadda_pg_rca32_fa746_y3 = f_s_dadda_pg_rca32_fa746_y0 & f_s_dadda_pg_rca32_fa746_f_s_dadda_pg_rca32_fa520_y2;
  assign f_s_dadda_pg_rca32_fa746_y4 = f_s_dadda_pg_rca32_fa746_y1 | f_s_dadda_pg_rca32_fa746_y3;
  assign f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa746_y4 = f_s_dadda_pg_rca32_fa746_y4;
  assign f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa745_y4 = f_s_dadda_pg_rca32_fa745_y4;
  assign f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa534_y2 = f_s_dadda_pg_rca32_fa534_y2;
  assign f_s_dadda_pg_rca32_fa747_y0 = f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa746_y4 ^ f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa745_y4;
  assign f_s_dadda_pg_rca32_fa747_y1 = f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa746_y4 & f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa745_y4;
  assign f_s_dadda_pg_rca32_fa747_y2 = f_s_dadda_pg_rca32_fa747_y0 ^ f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa534_y2;
  assign f_s_dadda_pg_rca32_fa747_y3 = f_s_dadda_pg_rca32_fa747_y0 & f_s_dadda_pg_rca32_fa747_f_s_dadda_pg_rca32_fa534_y2;
  assign f_s_dadda_pg_rca32_fa747_y4 = f_s_dadda_pg_rca32_fa747_y1 | f_s_dadda_pg_rca32_fa747_y3;
  assign f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa535_y2 = f_s_dadda_pg_rca32_fa535_y2;
  assign f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa536_y2 = f_s_dadda_pg_rca32_fa536_y2;
  assign f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa537_y2 = f_s_dadda_pg_rca32_fa537_y2;
  assign f_s_dadda_pg_rca32_fa748_y0 = f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa535_y2 ^ f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa536_y2;
  assign f_s_dadda_pg_rca32_fa748_y1 = f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa535_y2 & f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa536_y2;
  assign f_s_dadda_pg_rca32_fa748_y2 = f_s_dadda_pg_rca32_fa748_y0 ^ f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa537_y2;
  assign f_s_dadda_pg_rca32_fa748_y3 = f_s_dadda_pg_rca32_fa748_y0 & f_s_dadda_pg_rca32_fa748_f_s_dadda_pg_rca32_fa537_y2;
  assign f_s_dadda_pg_rca32_fa748_y4 = f_s_dadda_pg_rca32_fa748_y1 | f_s_dadda_pg_rca32_fa748_y3;
  assign f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa748_y4 = f_s_dadda_pg_rca32_fa748_y4;
  assign f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa747_y4 = f_s_dadda_pg_rca32_fa747_y4;
  assign f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa550_y2 = f_s_dadda_pg_rca32_fa550_y2;
  assign f_s_dadda_pg_rca32_fa749_y0 = f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa748_y4 ^ f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa747_y4;
  assign f_s_dadda_pg_rca32_fa749_y1 = f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa748_y4 & f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa747_y4;
  assign f_s_dadda_pg_rca32_fa749_y2 = f_s_dadda_pg_rca32_fa749_y0 ^ f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa550_y2;
  assign f_s_dadda_pg_rca32_fa749_y3 = f_s_dadda_pg_rca32_fa749_y0 & f_s_dadda_pg_rca32_fa749_f_s_dadda_pg_rca32_fa550_y2;
  assign f_s_dadda_pg_rca32_fa749_y4 = f_s_dadda_pg_rca32_fa749_y1 | f_s_dadda_pg_rca32_fa749_y3;
  assign f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa551_y2 = f_s_dadda_pg_rca32_fa551_y2;
  assign f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa552_y2 = f_s_dadda_pg_rca32_fa552_y2;
  assign f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa553_y2 = f_s_dadda_pg_rca32_fa553_y2;
  assign f_s_dadda_pg_rca32_fa750_y0 = f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa551_y2 ^ f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa552_y2;
  assign f_s_dadda_pg_rca32_fa750_y1 = f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa551_y2 & f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa552_y2;
  assign f_s_dadda_pg_rca32_fa750_y2 = f_s_dadda_pg_rca32_fa750_y0 ^ f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa553_y2;
  assign f_s_dadda_pg_rca32_fa750_y3 = f_s_dadda_pg_rca32_fa750_y0 & f_s_dadda_pg_rca32_fa750_f_s_dadda_pg_rca32_fa553_y2;
  assign f_s_dadda_pg_rca32_fa750_y4 = f_s_dadda_pg_rca32_fa750_y1 | f_s_dadda_pg_rca32_fa750_y3;
  assign f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa750_y4 = f_s_dadda_pg_rca32_fa750_y4;
  assign f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa749_y4 = f_s_dadda_pg_rca32_fa749_y4;
  assign f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa565_y2 = f_s_dadda_pg_rca32_fa565_y2;
  assign f_s_dadda_pg_rca32_fa751_y0 = f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa750_y4 ^ f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa749_y4;
  assign f_s_dadda_pg_rca32_fa751_y1 = f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa750_y4 & f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa749_y4;
  assign f_s_dadda_pg_rca32_fa751_y2 = f_s_dadda_pg_rca32_fa751_y0 ^ f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa565_y2;
  assign f_s_dadda_pg_rca32_fa751_y3 = f_s_dadda_pg_rca32_fa751_y0 & f_s_dadda_pg_rca32_fa751_f_s_dadda_pg_rca32_fa565_y2;
  assign f_s_dadda_pg_rca32_fa751_y4 = f_s_dadda_pg_rca32_fa751_y1 | f_s_dadda_pg_rca32_fa751_y3;
  assign f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa566_y2 = f_s_dadda_pg_rca32_fa566_y2;
  assign f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa567_y2 = f_s_dadda_pg_rca32_fa567_y2;
  assign f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa568_y2 = f_s_dadda_pg_rca32_fa568_y2;
  assign f_s_dadda_pg_rca32_fa752_y0 = f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa566_y2 ^ f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa567_y2;
  assign f_s_dadda_pg_rca32_fa752_y1 = f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa566_y2 & f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa567_y2;
  assign f_s_dadda_pg_rca32_fa752_y2 = f_s_dadda_pg_rca32_fa752_y0 ^ f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa568_y2;
  assign f_s_dadda_pg_rca32_fa752_y3 = f_s_dadda_pg_rca32_fa752_y0 & f_s_dadda_pg_rca32_fa752_f_s_dadda_pg_rca32_fa568_y2;
  assign f_s_dadda_pg_rca32_fa752_y4 = f_s_dadda_pg_rca32_fa752_y1 | f_s_dadda_pg_rca32_fa752_y3;
  assign f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa752_y4 = f_s_dadda_pg_rca32_fa752_y4;
  assign f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa751_y4 = f_s_dadda_pg_rca32_fa751_y4;
  assign f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa579_y2 = f_s_dadda_pg_rca32_fa579_y2;
  assign f_s_dadda_pg_rca32_fa753_y0 = f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa752_y4 ^ f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa751_y4;
  assign f_s_dadda_pg_rca32_fa753_y1 = f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa752_y4 & f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa751_y4;
  assign f_s_dadda_pg_rca32_fa753_y2 = f_s_dadda_pg_rca32_fa753_y0 ^ f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa579_y2;
  assign f_s_dadda_pg_rca32_fa753_y3 = f_s_dadda_pg_rca32_fa753_y0 & f_s_dadda_pg_rca32_fa753_f_s_dadda_pg_rca32_fa579_y2;
  assign f_s_dadda_pg_rca32_fa753_y4 = f_s_dadda_pg_rca32_fa753_y1 | f_s_dadda_pg_rca32_fa753_y3;
  assign f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa580_y2 = f_s_dadda_pg_rca32_fa580_y2;
  assign f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa581_y2 = f_s_dadda_pg_rca32_fa581_y2;
  assign f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa582_y2 = f_s_dadda_pg_rca32_fa582_y2;
  assign f_s_dadda_pg_rca32_fa754_y0 = f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa580_y2 ^ f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa581_y2;
  assign f_s_dadda_pg_rca32_fa754_y1 = f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa580_y2 & f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa581_y2;
  assign f_s_dadda_pg_rca32_fa754_y2 = f_s_dadda_pg_rca32_fa754_y0 ^ f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa582_y2;
  assign f_s_dadda_pg_rca32_fa754_y3 = f_s_dadda_pg_rca32_fa754_y0 & f_s_dadda_pg_rca32_fa754_f_s_dadda_pg_rca32_fa582_y2;
  assign f_s_dadda_pg_rca32_fa754_y4 = f_s_dadda_pg_rca32_fa754_y1 | f_s_dadda_pg_rca32_fa754_y3;
  assign f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa754_y4 = f_s_dadda_pg_rca32_fa754_y4;
  assign f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa753_y4 = f_s_dadda_pg_rca32_fa753_y4;
  assign f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa592_y2 = f_s_dadda_pg_rca32_fa592_y2;
  assign f_s_dadda_pg_rca32_fa755_y0 = f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa754_y4 ^ f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa753_y4;
  assign f_s_dadda_pg_rca32_fa755_y1 = f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa754_y4 & f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa753_y4;
  assign f_s_dadda_pg_rca32_fa755_y2 = f_s_dadda_pg_rca32_fa755_y0 ^ f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa592_y2;
  assign f_s_dadda_pg_rca32_fa755_y3 = f_s_dadda_pg_rca32_fa755_y0 & f_s_dadda_pg_rca32_fa755_f_s_dadda_pg_rca32_fa592_y2;
  assign f_s_dadda_pg_rca32_fa755_y4 = f_s_dadda_pg_rca32_fa755_y1 | f_s_dadda_pg_rca32_fa755_y3;
  assign f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa593_y2 = f_s_dadda_pg_rca32_fa593_y2;
  assign f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa594_y2 = f_s_dadda_pg_rca32_fa594_y2;
  assign f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa595_y2 = f_s_dadda_pg_rca32_fa595_y2;
  assign f_s_dadda_pg_rca32_fa756_y0 = f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa593_y2 ^ f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa594_y2;
  assign f_s_dadda_pg_rca32_fa756_y1 = f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa593_y2 & f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa594_y2;
  assign f_s_dadda_pg_rca32_fa756_y2 = f_s_dadda_pg_rca32_fa756_y0 ^ f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa595_y2;
  assign f_s_dadda_pg_rca32_fa756_y3 = f_s_dadda_pg_rca32_fa756_y0 & f_s_dadda_pg_rca32_fa756_f_s_dadda_pg_rca32_fa595_y2;
  assign f_s_dadda_pg_rca32_fa756_y4 = f_s_dadda_pg_rca32_fa756_y1 | f_s_dadda_pg_rca32_fa756_y3;
  assign f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa756_y4 = f_s_dadda_pg_rca32_fa756_y4;
  assign f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa755_y4 = f_s_dadda_pg_rca32_fa755_y4;
  assign f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa604_y2 = f_s_dadda_pg_rca32_fa604_y2;
  assign f_s_dadda_pg_rca32_fa757_y0 = f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa756_y4 ^ f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa755_y4;
  assign f_s_dadda_pg_rca32_fa757_y1 = f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa756_y4 & f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa755_y4;
  assign f_s_dadda_pg_rca32_fa757_y2 = f_s_dadda_pg_rca32_fa757_y0 ^ f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa604_y2;
  assign f_s_dadda_pg_rca32_fa757_y3 = f_s_dadda_pg_rca32_fa757_y0 & f_s_dadda_pg_rca32_fa757_f_s_dadda_pg_rca32_fa604_y2;
  assign f_s_dadda_pg_rca32_fa757_y4 = f_s_dadda_pg_rca32_fa757_y1 | f_s_dadda_pg_rca32_fa757_y3;
  assign f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa605_y2 = f_s_dadda_pg_rca32_fa605_y2;
  assign f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa606_y2 = f_s_dadda_pg_rca32_fa606_y2;
  assign f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa607_y2 = f_s_dadda_pg_rca32_fa607_y2;
  assign f_s_dadda_pg_rca32_fa758_y0 = f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa605_y2 ^ f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa606_y2;
  assign f_s_dadda_pg_rca32_fa758_y1 = f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa605_y2 & f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa606_y2;
  assign f_s_dadda_pg_rca32_fa758_y2 = f_s_dadda_pg_rca32_fa758_y0 ^ f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa607_y2;
  assign f_s_dadda_pg_rca32_fa758_y3 = f_s_dadda_pg_rca32_fa758_y0 & f_s_dadda_pg_rca32_fa758_f_s_dadda_pg_rca32_fa607_y2;
  assign f_s_dadda_pg_rca32_fa758_y4 = f_s_dadda_pg_rca32_fa758_y1 | f_s_dadda_pg_rca32_fa758_y3;
  assign f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa758_y4 = f_s_dadda_pg_rca32_fa758_y4;
  assign f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa757_y4 = f_s_dadda_pg_rca32_fa757_y4;
  assign f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa615_y2 = f_s_dadda_pg_rca32_fa615_y2;
  assign f_s_dadda_pg_rca32_fa759_y0 = f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa758_y4 ^ f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa757_y4;
  assign f_s_dadda_pg_rca32_fa759_y1 = f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa758_y4 & f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa757_y4;
  assign f_s_dadda_pg_rca32_fa759_y2 = f_s_dadda_pg_rca32_fa759_y0 ^ f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa615_y2;
  assign f_s_dadda_pg_rca32_fa759_y3 = f_s_dadda_pg_rca32_fa759_y0 & f_s_dadda_pg_rca32_fa759_f_s_dadda_pg_rca32_fa615_y2;
  assign f_s_dadda_pg_rca32_fa759_y4 = f_s_dadda_pg_rca32_fa759_y1 | f_s_dadda_pg_rca32_fa759_y3;
  assign f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa616_y2 = f_s_dadda_pg_rca32_fa616_y2;
  assign f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa617_y2 = f_s_dadda_pg_rca32_fa617_y2;
  assign f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa618_y2 = f_s_dadda_pg_rca32_fa618_y2;
  assign f_s_dadda_pg_rca32_fa760_y0 = f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa616_y2 ^ f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa617_y2;
  assign f_s_dadda_pg_rca32_fa760_y1 = f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa616_y2 & f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa617_y2;
  assign f_s_dadda_pg_rca32_fa760_y2 = f_s_dadda_pg_rca32_fa760_y0 ^ f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa618_y2;
  assign f_s_dadda_pg_rca32_fa760_y3 = f_s_dadda_pg_rca32_fa760_y0 & f_s_dadda_pg_rca32_fa760_f_s_dadda_pg_rca32_fa618_y2;
  assign f_s_dadda_pg_rca32_fa760_y4 = f_s_dadda_pg_rca32_fa760_y1 | f_s_dadda_pg_rca32_fa760_y3;
  assign f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa760_y4 = f_s_dadda_pg_rca32_fa760_y4;
  assign f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa759_y4 = f_s_dadda_pg_rca32_fa759_y4;
  assign f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa625_y2 = f_s_dadda_pg_rca32_fa625_y2;
  assign f_s_dadda_pg_rca32_fa761_y0 = f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa760_y4 ^ f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa759_y4;
  assign f_s_dadda_pg_rca32_fa761_y1 = f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa760_y4 & f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa759_y4;
  assign f_s_dadda_pg_rca32_fa761_y2 = f_s_dadda_pg_rca32_fa761_y0 ^ f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa625_y2;
  assign f_s_dadda_pg_rca32_fa761_y3 = f_s_dadda_pg_rca32_fa761_y0 & f_s_dadda_pg_rca32_fa761_f_s_dadda_pg_rca32_fa625_y2;
  assign f_s_dadda_pg_rca32_fa761_y4 = f_s_dadda_pg_rca32_fa761_y1 | f_s_dadda_pg_rca32_fa761_y3;
  assign f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa626_y2 = f_s_dadda_pg_rca32_fa626_y2;
  assign f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa627_y2 = f_s_dadda_pg_rca32_fa627_y2;
  assign f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa628_y2 = f_s_dadda_pg_rca32_fa628_y2;
  assign f_s_dadda_pg_rca32_fa762_y0 = f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa626_y2 ^ f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa627_y2;
  assign f_s_dadda_pg_rca32_fa762_y1 = f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa626_y2 & f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa627_y2;
  assign f_s_dadda_pg_rca32_fa762_y2 = f_s_dadda_pg_rca32_fa762_y0 ^ f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa628_y2;
  assign f_s_dadda_pg_rca32_fa762_y3 = f_s_dadda_pg_rca32_fa762_y0 & f_s_dadda_pg_rca32_fa762_f_s_dadda_pg_rca32_fa628_y2;
  assign f_s_dadda_pg_rca32_fa762_y4 = f_s_dadda_pg_rca32_fa762_y1 | f_s_dadda_pg_rca32_fa762_y3;
  assign f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa762_y4 = f_s_dadda_pg_rca32_fa762_y4;
  assign f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa761_y4 = f_s_dadda_pg_rca32_fa761_y4;
  assign f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa634_y2 = f_s_dadda_pg_rca32_fa634_y2;
  assign f_s_dadda_pg_rca32_fa763_y0 = f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa762_y4 ^ f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa761_y4;
  assign f_s_dadda_pg_rca32_fa763_y1 = f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa762_y4 & f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa761_y4;
  assign f_s_dadda_pg_rca32_fa763_y2 = f_s_dadda_pg_rca32_fa763_y0 ^ f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa634_y2;
  assign f_s_dadda_pg_rca32_fa763_y3 = f_s_dadda_pg_rca32_fa763_y0 & f_s_dadda_pg_rca32_fa763_f_s_dadda_pg_rca32_fa634_y2;
  assign f_s_dadda_pg_rca32_fa763_y4 = f_s_dadda_pg_rca32_fa763_y1 | f_s_dadda_pg_rca32_fa763_y3;
  assign f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa635_y2 = f_s_dadda_pg_rca32_fa635_y2;
  assign f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa636_y2 = f_s_dadda_pg_rca32_fa636_y2;
  assign f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa637_y2 = f_s_dadda_pg_rca32_fa637_y2;
  assign f_s_dadda_pg_rca32_fa764_y0 = f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa635_y2 ^ f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa636_y2;
  assign f_s_dadda_pg_rca32_fa764_y1 = f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa635_y2 & f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa636_y2;
  assign f_s_dadda_pg_rca32_fa764_y2 = f_s_dadda_pg_rca32_fa764_y0 ^ f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa637_y2;
  assign f_s_dadda_pg_rca32_fa764_y3 = f_s_dadda_pg_rca32_fa764_y0 & f_s_dadda_pg_rca32_fa764_f_s_dadda_pg_rca32_fa637_y2;
  assign f_s_dadda_pg_rca32_fa764_y4 = f_s_dadda_pg_rca32_fa764_y1 | f_s_dadda_pg_rca32_fa764_y3;
  assign f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa764_y4 = f_s_dadda_pg_rca32_fa764_y4;
  assign f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa763_y4 = f_s_dadda_pg_rca32_fa763_y4;
  assign f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa642_y2 = f_s_dadda_pg_rca32_fa642_y2;
  assign f_s_dadda_pg_rca32_fa765_y0 = f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa764_y4 ^ f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa763_y4;
  assign f_s_dadda_pg_rca32_fa765_y1 = f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa764_y4 & f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa763_y4;
  assign f_s_dadda_pg_rca32_fa765_y2 = f_s_dadda_pg_rca32_fa765_y0 ^ f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa642_y2;
  assign f_s_dadda_pg_rca32_fa765_y3 = f_s_dadda_pg_rca32_fa765_y0 & f_s_dadda_pg_rca32_fa765_f_s_dadda_pg_rca32_fa642_y2;
  assign f_s_dadda_pg_rca32_fa765_y4 = f_s_dadda_pg_rca32_fa765_y1 | f_s_dadda_pg_rca32_fa765_y3;
  assign f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa643_y2 = f_s_dadda_pg_rca32_fa643_y2;
  assign f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa644_y2 = f_s_dadda_pg_rca32_fa644_y2;
  assign f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa645_y2 = f_s_dadda_pg_rca32_fa645_y2;
  assign f_s_dadda_pg_rca32_fa766_y0 = f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa643_y2 ^ f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa644_y2;
  assign f_s_dadda_pg_rca32_fa766_y1 = f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa643_y2 & f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa644_y2;
  assign f_s_dadda_pg_rca32_fa766_y2 = f_s_dadda_pg_rca32_fa766_y0 ^ f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa645_y2;
  assign f_s_dadda_pg_rca32_fa766_y3 = f_s_dadda_pg_rca32_fa766_y0 & f_s_dadda_pg_rca32_fa766_f_s_dadda_pg_rca32_fa645_y2;
  assign f_s_dadda_pg_rca32_fa766_y4 = f_s_dadda_pg_rca32_fa766_y1 | f_s_dadda_pg_rca32_fa766_y3;
  assign f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa766_y4 = f_s_dadda_pg_rca32_fa766_y4;
  assign f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa765_y4 = f_s_dadda_pg_rca32_fa765_y4;
  assign f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa649_y2 = f_s_dadda_pg_rca32_fa649_y2;
  assign f_s_dadda_pg_rca32_fa767_y0 = f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa766_y4 ^ f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa765_y4;
  assign f_s_dadda_pg_rca32_fa767_y1 = f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa766_y4 & f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa765_y4;
  assign f_s_dadda_pg_rca32_fa767_y2 = f_s_dadda_pg_rca32_fa767_y0 ^ f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa649_y2;
  assign f_s_dadda_pg_rca32_fa767_y3 = f_s_dadda_pg_rca32_fa767_y0 & f_s_dadda_pg_rca32_fa767_f_s_dadda_pg_rca32_fa649_y2;
  assign f_s_dadda_pg_rca32_fa767_y4 = f_s_dadda_pg_rca32_fa767_y1 | f_s_dadda_pg_rca32_fa767_y3;
  assign f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa650_y2 = f_s_dadda_pg_rca32_fa650_y2;
  assign f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa651_y2 = f_s_dadda_pg_rca32_fa651_y2;
  assign f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa652_y2 = f_s_dadda_pg_rca32_fa652_y2;
  assign f_s_dadda_pg_rca32_fa768_y0 = f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa650_y2 ^ f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa651_y2;
  assign f_s_dadda_pg_rca32_fa768_y1 = f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa650_y2 & f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa651_y2;
  assign f_s_dadda_pg_rca32_fa768_y2 = f_s_dadda_pg_rca32_fa768_y0 ^ f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa652_y2;
  assign f_s_dadda_pg_rca32_fa768_y3 = f_s_dadda_pg_rca32_fa768_y0 & f_s_dadda_pg_rca32_fa768_f_s_dadda_pg_rca32_fa652_y2;
  assign f_s_dadda_pg_rca32_fa768_y4 = f_s_dadda_pg_rca32_fa768_y1 | f_s_dadda_pg_rca32_fa768_y3;
  assign f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa768_y4 = f_s_dadda_pg_rca32_fa768_y4;
  assign f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa767_y4 = f_s_dadda_pg_rca32_fa767_y4;
  assign f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa655_y2 = f_s_dadda_pg_rca32_fa655_y2;
  assign f_s_dadda_pg_rca32_fa769_y0 = f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa768_y4 ^ f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa767_y4;
  assign f_s_dadda_pg_rca32_fa769_y1 = f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa768_y4 & f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa767_y4;
  assign f_s_dadda_pg_rca32_fa769_y2 = f_s_dadda_pg_rca32_fa769_y0 ^ f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa655_y2;
  assign f_s_dadda_pg_rca32_fa769_y3 = f_s_dadda_pg_rca32_fa769_y0 & f_s_dadda_pg_rca32_fa769_f_s_dadda_pg_rca32_fa655_y2;
  assign f_s_dadda_pg_rca32_fa769_y4 = f_s_dadda_pg_rca32_fa769_y1 | f_s_dadda_pg_rca32_fa769_y3;
  assign f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa656_y2 = f_s_dadda_pg_rca32_fa656_y2;
  assign f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa657_y2 = f_s_dadda_pg_rca32_fa657_y2;
  assign f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa658_y2 = f_s_dadda_pg_rca32_fa658_y2;
  assign f_s_dadda_pg_rca32_fa770_y0 = f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa656_y2 ^ f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa657_y2;
  assign f_s_dadda_pg_rca32_fa770_y1 = f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa656_y2 & f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa657_y2;
  assign f_s_dadda_pg_rca32_fa770_y2 = f_s_dadda_pg_rca32_fa770_y0 ^ f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa658_y2;
  assign f_s_dadda_pg_rca32_fa770_y3 = f_s_dadda_pg_rca32_fa770_y0 & f_s_dadda_pg_rca32_fa770_f_s_dadda_pg_rca32_fa658_y2;
  assign f_s_dadda_pg_rca32_fa770_y4 = f_s_dadda_pg_rca32_fa770_y1 | f_s_dadda_pg_rca32_fa770_y3;
  assign f_s_dadda_pg_rca32_nand_22_31_a_22 = a_22;
  assign f_s_dadda_pg_rca32_nand_22_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_22_31_y0 = ~(f_s_dadda_pg_rca32_nand_22_31_a_22 & f_s_dadda_pg_rca32_nand_22_31_b_31);
  assign f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_fa770_y4 = f_s_dadda_pg_rca32_fa770_y4;
  assign f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_fa769_y4 = f_s_dadda_pg_rca32_fa769_y4;
  assign f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_nand_22_31_y0 = f_s_dadda_pg_rca32_nand_22_31_y0;
  assign f_s_dadda_pg_rca32_fa771_y0 = f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_fa770_y4 ^ f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_fa769_y4;
  assign f_s_dadda_pg_rca32_fa771_y1 = f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_fa770_y4 & f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_fa769_y4;
  assign f_s_dadda_pg_rca32_fa771_y2 = f_s_dadda_pg_rca32_fa771_y0 ^ f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_nand_22_31_y0;
  assign f_s_dadda_pg_rca32_fa771_y3 = f_s_dadda_pg_rca32_fa771_y0 & f_s_dadda_pg_rca32_fa771_f_s_dadda_pg_rca32_nand_22_31_y0;
  assign f_s_dadda_pg_rca32_fa771_y4 = f_s_dadda_pg_rca32_fa771_y1 | f_s_dadda_pg_rca32_fa771_y3;
  assign f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa661_y2 = f_s_dadda_pg_rca32_fa661_y2;
  assign f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa662_y2 = f_s_dadda_pg_rca32_fa662_y2;
  assign f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa663_y2 = f_s_dadda_pg_rca32_fa663_y2;
  assign f_s_dadda_pg_rca32_fa772_y0 = f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa661_y2 ^ f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa662_y2;
  assign f_s_dadda_pg_rca32_fa772_y1 = f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa661_y2 & f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa662_y2;
  assign f_s_dadda_pg_rca32_fa772_y2 = f_s_dadda_pg_rca32_fa772_y0 ^ f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa663_y2;
  assign f_s_dadda_pg_rca32_fa772_y3 = f_s_dadda_pg_rca32_fa772_y0 & f_s_dadda_pg_rca32_fa772_f_s_dadda_pg_rca32_fa663_y2;
  assign f_s_dadda_pg_rca32_fa772_y4 = f_s_dadda_pg_rca32_fa772_y1 | f_s_dadda_pg_rca32_fa772_y3;
  assign f_s_dadda_pg_rca32_and_24_30_a_24 = a_24;
  assign f_s_dadda_pg_rca32_and_24_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_24_30_y0 = f_s_dadda_pg_rca32_and_24_30_a_24 & f_s_dadda_pg_rca32_and_24_30_b_30;
  assign f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_fa772_y4 = f_s_dadda_pg_rca32_fa772_y4;
  assign f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_fa771_y4 = f_s_dadda_pg_rca32_fa771_y4;
  assign f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_and_24_30_y0 = f_s_dadda_pg_rca32_and_24_30_y0;
  assign f_s_dadda_pg_rca32_fa773_y0 = f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_fa772_y4 ^ f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_fa771_y4;
  assign f_s_dadda_pg_rca32_fa773_y1 = f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_fa772_y4 & f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_fa771_y4;
  assign f_s_dadda_pg_rca32_fa773_y2 = f_s_dadda_pg_rca32_fa773_y0 ^ f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_and_24_30_y0;
  assign f_s_dadda_pg_rca32_fa773_y3 = f_s_dadda_pg_rca32_fa773_y0 & f_s_dadda_pg_rca32_fa773_f_s_dadda_pg_rca32_and_24_30_y0;
  assign f_s_dadda_pg_rca32_fa773_y4 = f_s_dadda_pg_rca32_fa773_y1 | f_s_dadda_pg_rca32_fa773_y3;
  assign f_s_dadda_pg_rca32_nand_23_31_a_23 = a_23;
  assign f_s_dadda_pg_rca32_nand_23_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_23_31_y0 = ~(f_s_dadda_pg_rca32_nand_23_31_a_23 & f_s_dadda_pg_rca32_nand_23_31_b_31);
  assign f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_nand_23_31_y0 = f_s_dadda_pg_rca32_nand_23_31_y0;
  assign f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_fa666_y2 = f_s_dadda_pg_rca32_fa666_y2;
  assign f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_fa667_y2 = f_s_dadda_pg_rca32_fa667_y2;
  assign f_s_dadda_pg_rca32_fa774_y0 = f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_nand_23_31_y0 ^ f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_fa666_y2;
  assign f_s_dadda_pg_rca32_fa774_y1 = f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_nand_23_31_y0 & f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_fa666_y2;
  assign f_s_dadda_pg_rca32_fa774_y2 = f_s_dadda_pg_rca32_fa774_y0 ^ f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_fa667_y2;
  assign f_s_dadda_pg_rca32_fa774_y3 = f_s_dadda_pg_rca32_fa774_y0 & f_s_dadda_pg_rca32_fa774_f_s_dadda_pg_rca32_fa667_y2;
  assign f_s_dadda_pg_rca32_fa774_y4 = f_s_dadda_pg_rca32_fa774_y1 | f_s_dadda_pg_rca32_fa774_y3;
  assign f_s_dadda_pg_rca32_and_26_29_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_26_29_y0 = f_s_dadda_pg_rca32_and_26_29_a_26 & f_s_dadda_pg_rca32_and_26_29_b_29;
  assign f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_fa774_y4 = f_s_dadda_pg_rca32_fa774_y4;
  assign f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_fa773_y4 = f_s_dadda_pg_rca32_fa773_y4;
  assign f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_and_26_29_y0 = f_s_dadda_pg_rca32_and_26_29_y0;
  assign f_s_dadda_pg_rca32_fa775_y0 = f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_fa774_y4 ^ f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_fa773_y4;
  assign f_s_dadda_pg_rca32_fa775_y1 = f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_fa774_y4 & f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_fa773_y4;
  assign f_s_dadda_pg_rca32_fa775_y2 = f_s_dadda_pg_rca32_fa775_y0 ^ f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_and_26_29_y0;
  assign f_s_dadda_pg_rca32_fa775_y3 = f_s_dadda_pg_rca32_fa775_y0 & f_s_dadda_pg_rca32_fa775_f_s_dadda_pg_rca32_and_26_29_y0;
  assign f_s_dadda_pg_rca32_fa775_y4 = f_s_dadda_pg_rca32_fa775_y1 | f_s_dadda_pg_rca32_fa775_y3;
  assign f_s_dadda_pg_rca32_and_25_30_a_25 = a_25;
  assign f_s_dadda_pg_rca32_and_25_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_25_30_y0 = f_s_dadda_pg_rca32_and_25_30_a_25 & f_s_dadda_pg_rca32_and_25_30_b_30;
  assign f_s_dadda_pg_rca32_nand_24_31_a_24 = a_24;
  assign f_s_dadda_pg_rca32_nand_24_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_24_31_y0 = ~(f_s_dadda_pg_rca32_nand_24_31_a_24 & f_s_dadda_pg_rca32_nand_24_31_b_31);
  assign f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_and_25_30_y0 = f_s_dadda_pg_rca32_and_25_30_y0;
  assign f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_nand_24_31_y0 = f_s_dadda_pg_rca32_nand_24_31_y0;
  assign f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_fa670_y2 = f_s_dadda_pg_rca32_fa670_y2;
  assign f_s_dadda_pg_rca32_fa776_y0 = f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_and_25_30_y0 ^ f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_nand_24_31_y0;
  assign f_s_dadda_pg_rca32_fa776_y1 = f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_and_25_30_y0 & f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_nand_24_31_y0;
  assign f_s_dadda_pg_rca32_fa776_y2 = f_s_dadda_pg_rca32_fa776_y0 ^ f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_fa670_y2;
  assign f_s_dadda_pg_rca32_fa776_y3 = f_s_dadda_pg_rca32_fa776_y0 & f_s_dadda_pg_rca32_fa776_f_s_dadda_pg_rca32_fa670_y2;
  assign f_s_dadda_pg_rca32_fa776_y4 = f_s_dadda_pg_rca32_fa776_y1 | f_s_dadda_pg_rca32_fa776_y3;
  assign f_s_dadda_pg_rca32_and_28_28_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_28_28_y0 = f_s_dadda_pg_rca32_and_28_28_a_28 & f_s_dadda_pg_rca32_and_28_28_b_28;
  assign f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_fa776_y4 = f_s_dadda_pg_rca32_fa776_y4;
  assign f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_fa775_y4 = f_s_dadda_pg_rca32_fa775_y4;
  assign f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_and_28_28_y0 = f_s_dadda_pg_rca32_and_28_28_y0;
  assign f_s_dadda_pg_rca32_fa777_y0 = f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_fa776_y4 ^ f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_fa775_y4;
  assign f_s_dadda_pg_rca32_fa777_y1 = f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_fa776_y4 & f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_fa775_y4;
  assign f_s_dadda_pg_rca32_fa777_y2 = f_s_dadda_pg_rca32_fa777_y0 ^ f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_and_28_28_y0;
  assign f_s_dadda_pg_rca32_fa777_y3 = f_s_dadda_pg_rca32_fa777_y0 & f_s_dadda_pg_rca32_fa777_f_s_dadda_pg_rca32_and_28_28_y0;
  assign f_s_dadda_pg_rca32_fa777_y4 = f_s_dadda_pg_rca32_fa777_y1 | f_s_dadda_pg_rca32_fa777_y3;
  assign f_s_dadda_pg_rca32_and_27_29_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_27_29_y0 = f_s_dadda_pg_rca32_and_27_29_a_27 & f_s_dadda_pg_rca32_and_27_29_b_29;
  assign f_s_dadda_pg_rca32_and_26_30_a_26 = a_26;
  assign f_s_dadda_pg_rca32_and_26_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_26_30_y0 = f_s_dadda_pg_rca32_and_26_30_a_26 & f_s_dadda_pg_rca32_and_26_30_b_30;
  assign f_s_dadda_pg_rca32_nand_25_31_a_25 = a_25;
  assign f_s_dadda_pg_rca32_nand_25_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_25_31_y0 = ~(f_s_dadda_pg_rca32_nand_25_31_a_25 & f_s_dadda_pg_rca32_nand_25_31_b_31);
  assign f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_and_27_29_y0 = f_s_dadda_pg_rca32_and_27_29_y0;
  assign f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_and_26_30_y0 = f_s_dadda_pg_rca32_and_26_30_y0;
  assign f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_nand_25_31_y0 = f_s_dadda_pg_rca32_nand_25_31_y0;
  assign f_s_dadda_pg_rca32_fa778_y0 = f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_and_27_29_y0 ^ f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_and_26_30_y0;
  assign f_s_dadda_pg_rca32_fa778_y1 = f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_and_27_29_y0 & f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_and_26_30_y0;
  assign f_s_dadda_pg_rca32_fa778_y2 = f_s_dadda_pg_rca32_fa778_y0 ^ f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_nand_25_31_y0;
  assign f_s_dadda_pg_rca32_fa778_y3 = f_s_dadda_pg_rca32_fa778_y0 & f_s_dadda_pg_rca32_fa778_f_s_dadda_pg_rca32_nand_25_31_y0;
  assign f_s_dadda_pg_rca32_fa778_y4 = f_s_dadda_pg_rca32_fa778_y1 | f_s_dadda_pg_rca32_fa778_y3;
  assign f_s_dadda_pg_rca32_and_30_27_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_and_30_27_y0 = f_s_dadda_pg_rca32_and_30_27_a_30 & f_s_dadda_pg_rca32_and_30_27_b_27;
  assign f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_fa778_y4 = f_s_dadda_pg_rca32_fa778_y4;
  assign f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_fa777_y4 = f_s_dadda_pg_rca32_fa777_y4;
  assign f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_and_30_27_y0 = f_s_dadda_pg_rca32_and_30_27_y0;
  assign f_s_dadda_pg_rca32_fa779_y0 = f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_fa778_y4 ^ f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_fa777_y4;
  assign f_s_dadda_pg_rca32_fa779_y1 = f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_fa778_y4 & f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_fa777_y4;
  assign f_s_dadda_pg_rca32_fa779_y2 = f_s_dadda_pg_rca32_fa779_y0 ^ f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_and_30_27_y0;
  assign f_s_dadda_pg_rca32_fa779_y3 = f_s_dadda_pg_rca32_fa779_y0 & f_s_dadda_pg_rca32_fa779_f_s_dadda_pg_rca32_and_30_27_y0;
  assign f_s_dadda_pg_rca32_fa779_y4 = f_s_dadda_pg_rca32_fa779_y1 | f_s_dadda_pg_rca32_fa779_y3;
  assign f_s_dadda_pg_rca32_and_29_28_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_29_28_y0 = f_s_dadda_pg_rca32_and_29_28_a_29 & f_s_dadda_pg_rca32_and_29_28_b_28;
  assign f_s_dadda_pg_rca32_and_28_29_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_28_29_y0 = f_s_dadda_pg_rca32_and_28_29_a_28 & f_s_dadda_pg_rca32_and_28_29_b_29;
  assign f_s_dadda_pg_rca32_and_27_30_a_27 = a_27;
  assign f_s_dadda_pg_rca32_and_27_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_27_30_y0 = f_s_dadda_pg_rca32_and_27_30_a_27 & f_s_dadda_pg_rca32_and_27_30_b_30;
  assign f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_29_28_y0 = f_s_dadda_pg_rca32_and_29_28_y0;
  assign f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_28_29_y0 = f_s_dadda_pg_rca32_and_28_29_y0;
  assign f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_27_30_y0 = f_s_dadda_pg_rca32_and_27_30_y0;
  assign f_s_dadda_pg_rca32_fa780_y0 = f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_29_28_y0 ^ f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_28_29_y0;
  assign f_s_dadda_pg_rca32_fa780_y1 = f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_29_28_y0 & f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_28_29_y0;
  assign f_s_dadda_pg_rca32_fa780_y2 = f_s_dadda_pg_rca32_fa780_y0 ^ f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_27_30_y0;
  assign f_s_dadda_pg_rca32_fa780_y3 = f_s_dadda_pg_rca32_fa780_y0 & f_s_dadda_pg_rca32_fa780_f_s_dadda_pg_rca32_and_27_30_y0;
  assign f_s_dadda_pg_rca32_fa780_y4 = f_s_dadda_pg_rca32_fa780_y1 | f_s_dadda_pg_rca32_fa780_y3;
  assign f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa780_y4 = f_s_dadda_pg_rca32_fa780_y4;
  assign f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa779_y4 = f_s_dadda_pg_rca32_fa779_y4;
  assign f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa675_y4 = f_s_dadda_pg_rca32_fa675_y4;
  assign f_s_dadda_pg_rca32_fa781_y0 = f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa780_y4 ^ f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa779_y4;
  assign f_s_dadda_pg_rca32_fa781_y1 = f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa780_y4 & f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa779_y4;
  assign f_s_dadda_pg_rca32_fa781_y2 = f_s_dadda_pg_rca32_fa781_y0 ^ f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa675_y4;
  assign f_s_dadda_pg_rca32_fa781_y3 = f_s_dadda_pg_rca32_fa781_y0 & f_s_dadda_pg_rca32_fa781_f_s_dadda_pg_rca32_fa675_y4;
  assign f_s_dadda_pg_rca32_fa781_y4 = f_s_dadda_pg_rca32_fa781_y1 | f_s_dadda_pg_rca32_fa781_y3;
  assign f_s_dadda_pg_rca32_nand_31_27_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_27_b_27 = b_27;
  assign f_s_dadda_pg_rca32_nand_31_27_y0 = ~(f_s_dadda_pg_rca32_nand_31_27_a_31 & f_s_dadda_pg_rca32_nand_31_27_b_27);
  assign f_s_dadda_pg_rca32_and_30_28_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_and_30_28_y0 = f_s_dadda_pg_rca32_and_30_28_a_30 & f_s_dadda_pg_rca32_and_30_28_b_28;
  assign f_s_dadda_pg_rca32_and_29_29_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_29_29_y0 = f_s_dadda_pg_rca32_and_29_29_a_29 & f_s_dadda_pg_rca32_and_29_29_b_29;
  assign f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_nand_31_27_y0 = f_s_dadda_pg_rca32_nand_31_27_y0;
  assign f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_and_30_28_y0 = f_s_dadda_pg_rca32_and_30_28_y0;
  assign f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_and_29_29_y0 = f_s_dadda_pg_rca32_and_29_29_y0;
  assign f_s_dadda_pg_rca32_fa782_y0 = f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_nand_31_27_y0 ^ f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_and_30_28_y0;
  assign f_s_dadda_pg_rca32_fa782_y1 = f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_nand_31_27_y0 & f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_and_30_28_y0;
  assign f_s_dadda_pg_rca32_fa782_y2 = f_s_dadda_pg_rca32_fa782_y0 ^ f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_and_29_29_y0;
  assign f_s_dadda_pg_rca32_fa782_y3 = f_s_dadda_pg_rca32_fa782_y0 & f_s_dadda_pg_rca32_fa782_f_s_dadda_pg_rca32_and_29_29_y0;
  assign f_s_dadda_pg_rca32_fa782_y4 = f_s_dadda_pg_rca32_fa782_y1 | f_s_dadda_pg_rca32_fa782_y3;
  assign f_s_dadda_pg_rca32_nand_31_28_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_28_b_28 = b_28;
  assign f_s_dadda_pg_rca32_nand_31_28_y0 = ~(f_s_dadda_pg_rca32_nand_31_28_a_31 & f_s_dadda_pg_rca32_nand_31_28_b_28);
  assign f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_fa782_y4 = f_s_dadda_pg_rca32_fa782_y4;
  assign f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_fa781_y4 = f_s_dadda_pg_rca32_fa781_y4;
  assign f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_nand_31_28_y0 = f_s_dadda_pg_rca32_nand_31_28_y0;
  assign f_s_dadda_pg_rca32_fa783_y0 = f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_fa782_y4 ^ f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_fa781_y4;
  assign f_s_dadda_pg_rca32_fa783_y1 = f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_fa782_y4 & f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_fa781_y4;
  assign f_s_dadda_pg_rca32_fa783_y2 = f_s_dadda_pg_rca32_fa783_y0 ^ f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_nand_31_28_y0;
  assign f_s_dadda_pg_rca32_fa783_y3 = f_s_dadda_pg_rca32_fa783_y0 & f_s_dadda_pg_rca32_fa783_f_s_dadda_pg_rca32_nand_31_28_y0;
  assign f_s_dadda_pg_rca32_fa783_y4 = f_s_dadda_pg_rca32_fa783_y1 | f_s_dadda_pg_rca32_fa783_y3;
  assign f_s_dadda_pg_rca32_and_3_0_a_3 = a_3;
  assign f_s_dadda_pg_rca32_and_3_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_3_0_y0 = f_s_dadda_pg_rca32_and_3_0_a_3 & f_s_dadda_pg_rca32_and_3_0_b_0;
  assign f_s_dadda_pg_rca32_and_2_1_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_2_1_y0 = f_s_dadda_pg_rca32_and_2_1_a_2 & f_s_dadda_pg_rca32_and_2_1_b_1;
  assign f_s_dadda_pg_rca32_ha28_f_s_dadda_pg_rca32_and_3_0_y0 = f_s_dadda_pg_rca32_and_3_0_y0;
  assign f_s_dadda_pg_rca32_ha28_f_s_dadda_pg_rca32_and_2_1_y0 = f_s_dadda_pg_rca32_and_2_1_y0;
  assign f_s_dadda_pg_rca32_ha28_y0 = f_s_dadda_pg_rca32_ha28_f_s_dadda_pg_rca32_and_3_0_y0 ^ f_s_dadda_pg_rca32_ha28_f_s_dadda_pg_rca32_and_2_1_y0;
  assign f_s_dadda_pg_rca32_ha28_y1 = f_s_dadda_pg_rca32_ha28_f_s_dadda_pg_rca32_and_3_0_y0 & f_s_dadda_pg_rca32_ha28_f_s_dadda_pg_rca32_and_2_1_y0;
  assign f_s_dadda_pg_rca32_and_2_2_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_2_2_y0 = f_s_dadda_pg_rca32_and_2_2_a_2 & f_s_dadda_pg_rca32_and_2_2_b_2;
  assign f_s_dadda_pg_rca32_and_1_3_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_1_3_y0 = f_s_dadda_pg_rca32_and_1_3_a_1 & f_s_dadda_pg_rca32_and_1_3_b_3;
  assign f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_ha28_y1 = f_s_dadda_pg_rca32_ha28_y1;
  assign f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_and_2_2_y0 = f_s_dadda_pg_rca32_and_2_2_y0;
  assign f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_and_1_3_y0 = f_s_dadda_pg_rca32_and_1_3_y0;
  assign f_s_dadda_pg_rca32_fa784_y0 = f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_ha28_y1 ^ f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_and_2_2_y0;
  assign f_s_dadda_pg_rca32_fa784_y1 = f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_ha28_y1 & f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_and_2_2_y0;
  assign f_s_dadda_pg_rca32_fa784_y2 = f_s_dadda_pg_rca32_fa784_y0 ^ f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_and_1_3_y0;
  assign f_s_dadda_pg_rca32_fa784_y3 = f_s_dadda_pg_rca32_fa784_y0 & f_s_dadda_pg_rca32_fa784_f_s_dadda_pg_rca32_and_1_3_y0;
  assign f_s_dadda_pg_rca32_fa784_y4 = f_s_dadda_pg_rca32_fa784_y1 | f_s_dadda_pg_rca32_fa784_y3;
  assign f_s_dadda_pg_rca32_and_1_4_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_1_4_y0 = f_s_dadda_pg_rca32_and_1_4_a_1 & f_s_dadda_pg_rca32_and_1_4_b_4;
  assign f_s_dadda_pg_rca32_and_0_5_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_5_b_5 = b_5;
  assign f_s_dadda_pg_rca32_and_0_5_y0 = f_s_dadda_pg_rca32_and_0_5_a_0 & f_s_dadda_pg_rca32_and_0_5_b_5;
  assign f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_fa784_y4 = f_s_dadda_pg_rca32_fa784_y4;
  assign f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_and_1_4_y0 = f_s_dadda_pg_rca32_and_1_4_y0;
  assign f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_and_0_5_y0 = f_s_dadda_pg_rca32_and_0_5_y0;
  assign f_s_dadda_pg_rca32_fa785_y0 = f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_fa784_y4 ^ f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_and_1_4_y0;
  assign f_s_dadda_pg_rca32_fa785_y1 = f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_fa784_y4 & f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_and_1_4_y0;
  assign f_s_dadda_pg_rca32_fa785_y2 = f_s_dadda_pg_rca32_fa785_y0 ^ f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_and_0_5_y0;
  assign f_s_dadda_pg_rca32_fa785_y3 = f_s_dadda_pg_rca32_fa785_y0 & f_s_dadda_pg_rca32_fa785_f_s_dadda_pg_rca32_and_0_5_y0;
  assign f_s_dadda_pg_rca32_fa785_y4 = f_s_dadda_pg_rca32_fa785_y1 | f_s_dadda_pg_rca32_fa785_y3;
  assign f_s_dadda_pg_rca32_and_0_6_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_6_b_6 = b_6;
  assign f_s_dadda_pg_rca32_and_0_6_y0 = f_s_dadda_pg_rca32_and_0_6_a_0 & f_s_dadda_pg_rca32_and_0_6_b_6;
  assign f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_fa785_y4 = f_s_dadda_pg_rca32_fa785_y4;
  assign f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_and_0_6_y0 = f_s_dadda_pg_rca32_and_0_6_y0;
  assign f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_ha4_y0 = f_s_dadda_pg_rca32_ha4_y0;
  assign f_s_dadda_pg_rca32_fa786_y0 = f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_fa785_y4 ^ f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_and_0_6_y0;
  assign f_s_dadda_pg_rca32_fa786_y1 = f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_fa785_y4 & f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_and_0_6_y0;
  assign f_s_dadda_pg_rca32_fa786_y2 = f_s_dadda_pg_rca32_fa786_y0 ^ f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_ha4_y0;
  assign f_s_dadda_pg_rca32_fa786_y3 = f_s_dadda_pg_rca32_fa786_y0 & f_s_dadda_pg_rca32_fa786_f_s_dadda_pg_rca32_ha4_y0;
  assign f_s_dadda_pg_rca32_fa786_y4 = f_s_dadda_pg_rca32_fa786_y1 | f_s_dadda_pg_rca32_fa786_y3;
  assign f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_fa786_y4 = f_s_dadda_pg_rca32_fa786_y4;
  assign f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_fa16_y2 = f_s_dadda_pg_rca32_fa16_y2;
  assign f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_ha5_y0 = f_s_dadda_pg_rca32_ha5_y0;
  assign f_s_dadda_pg_rca32_fa787_y0 = f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_fa786_y4 ^ f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_fa16_y2;
  assign f_s_dadda_pg_rca32_fa787_y1 = f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_fa786_y4 & f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_fa16_y2;
  assign f_s_dadda_pg_rca32_fa787_y2 = f_s_dadda_pg_rca32_fa787_y0 ^ f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_ha5_y0;
  assign f_s_dadda_pg_rca32_fa787_y3 = f_s_dadda_pg_rca32_fa787_y0 & f_s_dadda_pg_rca32_fa787_f_s_dadda_pg_rca32_ha5_y0;
  assign f_s_dadda_pg_rca32_fa787_y4 = f_s_dadda_pg_rca32_fa787_y1 | f_s_dadda_pg_rca32_fa787_y3;
  assign f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_fa787_y4 = f_s_dadda_pg_rca32_fa787_y4;
  assign f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_fa18_y2 = f_s_dadda_pg_rca32_fa18_y2;
  assign f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_ha6_y0 = f_s_dadda_pg_rca32_ha6_y0;
  assign f_s_dadda_pg_rca32_fa788_y0 = f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_fa787_y4 ^ f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_fa18_y2;
  assign f_s_dadda_pg_rca32_fa788_y1 = f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_fa787_y4 & f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_fa18_y2;
  assign f_s_dadda_pg_rca32_fa788_y2 = f_s_dadda_pg_rca32_fa788_y0 ^ f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_ha6_y0;
  assign f_s_dadda_pg_rca32_fa788_y3 = f_s_dadda_pg_rca32_fa788_y0 & f_s_dadda_pg_rca32_fa788_f_s_dadda_pg_rca32_ha6_y0;
  assign f_s_dadda_pg_rca32_fa788_y4 = f_s_dadda_pg_rca32_fa788_y1 | f_s_dadda_pg_rca32_fa788_y3;
  assign f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_fa788_y4 = f_s_dadda_pg_rca32_fa788_y4;
  assign f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_fa21_y2 = f_s_dadda_pg_rca32_fa21_y2;
  assign f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_ha7_y0 = f_s_dadda_pg_rca32_ha7_y0;
  assign f_s_dadda_pg_rca32_fa789_y0 = f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_fa788_y4 ^ f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_fa21_y2;
  assign f_s_dadda_pg_rca32_fa789_y1 = f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_fa788_y4 & f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_fa21_y2;
  assign f_s_dadda_pg_rca32_fa789_y2 = f_s_dadda_pg_rca32_fa789_y0 ^ f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_ha7_y0;
  assign f_s_dadda_pg_rca32_fa789_y3 = f_s_dadda_pg_rca32_fa789_y0 & f_s_dadda_pg_rca32_fa789_f_s_dadda_pg_rca32_ha7_y0;
  assign f_s_dadda_pg_rca32_fa789_y4 = f_s_dadda_pg_rca32_fa789_y1 | f_s_dadda_pg_rca32_fa789_y3;
  assign f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_fa789_y4 = f_s_dadda_pg_rca32_fa789_y4;
  assign f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_fa25_y2 = f_s_dadda_pg_rca32_fa25_y2;
  assign f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_ha8_y0 = f_s_dadda_pg_rca32_ha8_y0;
  assign f_s_dadda_pg_rca32_fa790_y0 = f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_fa789_y4 ^ f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_fa25_y2;
  assign f_s_dadda_pg_rca32_fa790_y1 = f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_fa789_y4 & f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_fa25_y2;
  assign f_s_dadda_pg_rca32_fa790_y2 = f_s_dadda_pg_rca32_fa790_y0 ^ f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_ha8_y0;
  assign f_s_dadda_pg_rca32_fa790_y3 = f_s_dadda_pg_rca32_fa790_y0 & f_s_dadda_pg_rca32_fa790_f_s_dadda_pg_rca32_ha8_y0;
  assign f_s_dadda_pg_rca32_fa790_y4 = f_s_dadda_pg_rca32_fa790_y1 | f_s_dadda_pg_rca32_fa790_y3;
  assign f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_fa790_y4 = f_s_dadda_pg_rca32_fa790_y4;
  assign f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_fa30_y2 = f_s_dadda_pg_rca32_fa30_y2;
  assign f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_ha9_y0 = f_s_dadda_pg_rca32_ha9_y0;
  assign f_s_dadda_pg_rca32_fa791_y0 = f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_fa790_y4 ^ f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_fa30_y2;
  assign f_s_dadda_pg_rca32_fa791_y1 = f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_fa790_y4 & f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_fa30_y2;
  assign f_s_dadda_pg_rca32_fa791_y2 = f_s_dadda_pg_rca32_fa791_y0 ^ f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_ha9_y0;
  assign f_s_dadda_pg_rca32_fa791_y3 = f_s_dadda_pg_rca32_fa791_y0 & f_s_dadda_pg_rca32_fa791_f_s_dadda_pg_rca32_ha9_y0;
  assign f_s_dadda_pg_rca32_fa791_y4 = f_s_dadda_pg_rca32_fa791_y1 | f_s_dadda_pg_rca32_fa791_y3;
  assign f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_fa791_y4 = f_s_dadda_pg_rca32_fa791_y4;
  assign f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_fa36_y2 = f_s_dadda_pg_rca32_fa36_y2;
  assign f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_ha10_y0 = f_s_dadda_pg_rca32_ha10_y0;
  assign f_s_dadda_pg_rca32_fa792_y0 = f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_fa791_y4 ^ f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_fa36_y2;
  assign f_s_dadda_pg_rca32_fa792_y1 = f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_fa791_y4 & f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_fa36_y2;
  assign f_s_dadda_pg_rca32_fa792_y2 = f_s_dadda_pg_rca32_fa792_y0 ^ f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_ha10_y0;
  assign f_s_dadda_pg_rca32_fa792_y3 = f_s_dadda_pg_rca32_fa792_y0 & f_s_dadda_pg_rca32_fa792_f_s_dadda_pg_rca32_ha10_y0;
  assign f_s_dadda_pg_rca32_fa792_y4 = f_s_dadda_pg_rca32_fa792_y1 | f_s_dadda_pg_rca32_fa792_y3;
  assign f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_fa792_y4 = f_s_dadda_pg_rca32_fa792_y4;
  assign f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_fa43_y2 = f_s_dadda_pg_rca32_fa43_y2;
  assign f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_ha11_y0 = f_s_dadda_pg_rca32_ha11_y0;
  assign f_s_dadda_pg_rca32_fa793_y0 = f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_fa792_y4 ^ f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_fa43_y2;
  assign f_s_dadda_pg_rca32_fa793_y1 = f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_fa792_y4 & f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_fa43_y2;
  assign f_s_dadda_pg_rca32_fa793_y2 = f_s_dadda_pg_rca32_fa793_y0 ^ f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_ha11_y0;
  assign f_s_dadda_pg_rca32_fa793_y3 = f_s_dadda_pg_rca32_fa793_y0 & f_s_dadda_pg_rca32_fa793_f_s_dadda_pg_rca32_ha11_y0;
  assign f_s_dadda_pg_rca32_fa793_y4 = f_s_dadda_pg_rca32_fa793_y1 | f_s_dadda_pg_rca32_fa793_y3;
  assign f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_fa793_y4 = f_s_dadda_pg_rca32_fa793_y4;
  assign f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_fa51_y2 = f_s_dadda_pg_rca32_fa51_y2;
  assign f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_ha12_y0 = f_s_dadda_pg_rca32_ha12_y0;
  assign f_s_dadda_pg_rca32_fa794_y0 = f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_fa793_y4 ^ f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_fa51_y2;
  assign f_s_dadda_pg_rca32_fa794_y1 = f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_fa793_y4 & f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_fa51_y2;
  assign f_s_dadda_pg_rca32_fa794_y2 = f_s_dadda_pg_rca32_fa794_y0 ^ f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_ha12_y0;
  assign f_s_dadda_pg_rca32_fa794_y3 = f_s_dadda_pg_rca32_fa794_y0 & f_s_dadda_pg_rca32_fa794_f_s_dadda_pg_rca32_ha12_y0;
  assign f_s_dadda_pg_rca32_fa794_y4 = f_s_dadda_pg_rca32_fa794_y1 | f_s_dadda_pg_rca32_fa794_y3;
  assign f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_fa794_y4 = f_s_dadda_pg_rca32_fa794_y4;
  assign f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_fa60_y2 = f_s_dadda_pg_rca32_fa60_y2;
  assign f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_ha13_y0 = f_s_dadda_pg_rca32_ha13_y0;
  assign f_s_dadda_pg_rca32_fa795_y0 = f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_fa794_y4 ^ f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_fa60_y2;
  assign f_s_dadda_pg_rca32_fa795_y1 = f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_fa794_y4 & f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_fa60_y2;
  assign f_s_dadda_pg_rca32_fa795_y2 = f_s_dadda_pg_rca32_fa795_y0 ^ f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_ha13_y0;
  assign f_s_dadda_pg_rca32_fa795_y3 = f_s_dadda_pg_rca32_fa795_y0 & f_s_dadda_pg_rca32_fa795_f_s_dadda_pg_rca32_ha13_y0;
  assign f_s_dadda_pg_rca32_fa795_y4 = f_s_dadda_pg_rca32_fa795_y1 | f_s_dadda_pg_rca32_fa795_y3;
  assign f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_fa795_y4 = f_s_dadda_pg_rca32_fa795_y4;
  assign f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_fa70_y2 = f_s_dadda_pg_rca32_fa70_y2;
  assign f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_ha14_y0 = f_s_dadda_pg_rca32_ha14_y0;
  assign f_s_dadda_pg_rca32_fa796_y0 = f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_fa795_y4 ^ f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_fa70_y2;
  assign f_s_dadda_pg_rca32_fa796_y1 = f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_fa795_y4 & f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_fa70_y2;
  assign f_s_dadda_pg_rca32_fa796_y2 = f_s_dadda_pg_rca32_fa796_y0 ^ f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_ha14_y0;
  assign f_s_dadda_pg_rca32_fa796_y3 = f_s_dadda_pg_rca32_fa796_y0 & f_s_dadda_pg_rca32_fa796_f_s_dadda_pg_rca32_ha14_y0;
  assign f_s_dadda_pg_rca32_fa796_y4 = f_s_dadda_pg_rca32_fa796_y1 | f_s_dadda_pg_rca32_fa796_y3;
  assign f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_fa796_y4 = f_s_dadda_pg_rca32_fa796_y4;
  assign f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_fa81_y2 = f_s_dadda_pg_rca32_fa81_y2;
  assign f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_ha15_y0 = f_s_dadda_pg_rca32_ha15_y0;
  assign f_s_dadda_pg_rca32_fa797_y0 = f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_fa796_y4 ^ f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_fa81_y2;
  assign f_s_dadda_pg_rca32_fa797_y1 = f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_fa796_y4 & f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_fa81_y2;
  assign f_s_dadda_pg_rca32_fa797_y2 = f_s_dadda_pg_rca32_fa797_y0 ^ f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_ha15_y0;
  assign f_s_dadda_pg_rca32_fa797_y3 = f_s_dadda_pg_rca32_fa797_y0 & f_s_dadda_pg_rca32_fa797_f_s_dadda_pg_rca32_ha15_y0;
  assign f_s_dadda_pg_rca32_fa797_y4 = f_s_dadda_pg_rca32_fa797_y1 | f_s_dadda_pg_rca32_fa797_y3;
  assign f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_fa797_y4 = f_s_dadda_pg_rca32_fa797_y4;
  assign f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_fa93_y2 = f_s_dadda_pg_rca32_fa93_y2;
  assign f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_ha16_y0 = f_s_dadda_pg_rca32_ha16_y0;
  assign f_s_dadda_pg_rca32_fa798_y0 = f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_fa797_y4 ^ f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_fa93_y2;
  assign f_s_dadda_pg_rca32_fa798_y1 = f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_fa797_y4 & f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_fa93_y2;
  assign f_s_dadda_pg_rca32_fa798_y2 = f_s_dadda_pg_rca32_fa798_y0 ^ f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_ha16_y0;
  assign f_s_dadda_pg_rca32_fa798_y3 = f_s_dadda_pg_rca32_fa798_y0 & f_s_dadda_pg_rca32_fa798_f_s_dadda_pg_rca32_ha16_y0;
  assign f_s_dadda_pg_rca32_fa798_y4 = f_s_dadda_pg_rca32_fa798_y1 | f_s_dadda_pg_rca32_fa798_y3;
  assign f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_fa798_y4 = f_s_dadda_pg_rca32_fa798_y4;
  assign f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_fa106_y2 = f_s_dadda_pg_rca32_fa106_y2;
  assign f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_ha17_y0 = f_s_dadda_pg_rca32_ha17_y0;
  assign f_s_dadda_pg_rca32_fa799_y0 = f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_fa798_y4 ^ f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_fa106_y2;
  assign f_s_dadda_pg_rca32_fa799_y1 = f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_fa798_y4 & f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_fa106_y2;
  assign f_s_dadda_pg_rca32_fa799_y2 = f_s_dadda_pg_rca32_fa799_y0 ^ f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_ha17_y0;
  assign f_s_dadda_pg_rca32_fa799_y3 = f_s_dadda_pg_rca32_fa799_y0 & f_s_dadda_pg_rca32_fa799_f_s_dadda_pg_rca32_ha17_y0;
  assign f_s_dadda_pg_rca32_fa799_y4 = f_s_dadda_pg_rca32_fa799_y1 | f_s_dadda_pg_rca32_fa799_y3;
  assign f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_fa799_y4 = f_s_dadda_pg_rca32_fa799_y4;
  assign f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_fa120_y2 = f_s_dadda_pg_rca32_fa120_y2;
  assign f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_ha18_y0 = f_s_dadda_pg_rca32_ha18_y0;
  assign f_s_dadda_pg_rca32_fa800_y0 = f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_fa799_y4 ^ f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_fa120_y2;
  assign f_s_dadda_pg_rca32_fa800_y1 = f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_fa799_y4 & f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_fa120_y2;
  assign f_s_dadda_pg_rca32_fa800_y2 = f_s_dadda_pg_rca32_fa800_y0 ^ f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_ha18_y0;
  assign f_s_dadda_pg_rca32_fa800_y3 = f_s_dadda_pg_rca32_fa800_y0 & f_s_dadda_pg_rca32_fa800_f_s_dadda_pg_rca32_ha18_y0;
  assign f_s_dadda_pg_rca32_fa800_y4 = f_s_dadda_pg_rca32_fa800_y1 | f_s_dadda_pg_rca32_fa800_y3;
  assign f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_fa800_y4 = f_s_dadda_pg_rca32_fa800_y4;
  assign f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_fa135_y2 = f_s_dadda_pg_rca32_fa135_y2;
  assign f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_ha19_y0 = f_s_dadda_pg_rca32_ha19_y0;
  assign f_s_dadda_pg_rca32_fa801_y0 = f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_fa800_y4 ^ f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_fa135_y2;
  assign f_s_dadda_pg_rca32_fa801_y1 = f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_fa800_y4 & f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_fa135_y2;
  assign f_s_dadda_pg_rca32_fa801_y2 = f_s_dadda_pg_rca32_fa801_y0 ^ f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_ha19_y0;
  assign f_s_dadda_pg_rca32_fa801_y3 = f_s_dadda_pg_rca32_fa801_y0 & f_s_dadda_pg_rca32_fa801_f_s_dadda_pg_rca32_ha19_y0;
  assign f_s_dadda_pg_rca32_fa801_y4 = f_s_dadda_pg_rca32_fa801_y1 | f_s_dadda_pg_rca32_fa801_y3;
  assign f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_fa801_y4 = f_s_dadda_pg_rca32_fa801_y4;
  assign f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_fa151_y2 = f_s_dadda_pg_rca32_fa151_y2;
  assign f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_ha20_y0 = f_s_dadda_pg_rca32_ha20_y0;
  assign f_s_dadda_pg_rca32_fa802_y0 = f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_fa801_y4 ^ f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_fa151_y2;
  assign f_s_dadda_pg_rca32_fa802_y1 = f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_fa801_y4 & f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_fa151_y2;
  assign f_s_dadda_pg_rca32_fa802_y2 = f_s_dadda_pg_rca32_fa802_y0 ^ f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_ha20_y0;
  assign f_s_dadda_pg_rca32_fa802_y3 = f_s_dadda_pg_rca32_fa802_y0 & f_s_dadda_pg_rca32_fa802_f_s_dadda_pg_rca32_ha20_y0;
  assign f_s_dadda_pg_rca32_fa802_y4 = f_s_dadda_pg_rca32_fa802_y1 | f_s_dadda_pg_rca32_fa802_y3;
  assign f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_fa802_y4 = f_s_dadda_pg_rca32_fa802_y4;
  assign f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_fa168_y2 = f_s_dadda_pg_rca32_fa168_y2;
  assign f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_ha21_y0 = f_s_dadda_pg_rca32_ha21_y0;
  assign f_s_dadda_pg_rca32_fa803_y0 = f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_fa802_y4 ^ f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_fa168_y2;
  assign f_s_dadda_pg_rca32_fa803_y1 = f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_fa802_y4 & f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_fa168_y2;
  assign f_s_dadda_pg_rca32_fa803_y2 = f_s_dadda_pg_rca32_fa803_y0 ^ f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_ha21_y0;
  assign f_s_dadda_pg_rca32_fa803_y3 = f_s_dadda_pg_rca32_fa803_y0 & f_s_dadda_pg_rca32_fa803_f_s_dadda_pg_rca32_ha21_y0;
  assign f_s_dadda_pg_rca32_fa803_y4 = f_s_dadda_pg_rca32_fa803_y1 | f_s_dadda_pg_rca32_fa803_y3;
  assign f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_fa803_y4 = f_s_dadda_pg_rca32_fa803_y4;
  assign f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_fa186_y2 = f_s_dadda_pg_rca32_fa186_y2;
  assign f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_ha22_y0 = f_s_dadda_pg_rca32_ha22_y0;
  assign f_s_dadda_pg_rca32_fa804_y0 = f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_fa803_y4 ^ f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_fa186_y2;
  assign f_s_dadda_pg_rca32_fa804_y1 = f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_fa803_y4 & f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_fa186_y2;
  assign f_s_dadda_pg_rca32_fa804_y2 = f_s_dadda_pg_rca32_fa804_y0 ^ f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_ha22_y0;
  assign f_s_dadda_pg_rca32_fa804_y3 = f_s_dadda_pg_rca32_fa804_y0 & f_s_dadda_pg_rca32_fa804_f_s_dadda_pg_rca32_ha22_y0;
  assign f_s_dadda_pg_rca32_fa804_y4 = f_s_dadda_pg_rca32_fa804_y1 | f_s_dadda_pg_rca32_fa804_y3;
  assign f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_fa804_y4 = f_s_dadda_pg_rca32_fa804_y4;
  assign f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_fa205_y2 = f_s_dadda_pg_rca32_fa205_y2;
  assign f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_ha23_y0 = f_s_dadda_pg_rca32_ha23_y0;
  assign f_s_dadda_pg_rca32_fa805_y0 = f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_fa804_y4 ^ f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_fa205_y2;
  assign f_s_dadda_pg_rca32_fa805_y1 = f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_fa804_y4 & f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_fa205_y2;
  assign f_s_dadda_pg_rca32_fa805_y2 = f_s_dadda_pg_rca32_fa805_y0 ^ f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_ha23_y0;
  assign f_s_dadda_pg_rca32_fa805_y3 = f_s_dadda_pg_rca32_fa805_y0 & f_s_dadda_pg_rca32_fa805_f_s_dadda_pg_rca32_ha23_y0;
  assign f_s_dadda_pg_rca32_fa805_y4 = f_s_dadda_pg_rca32_fa805_y1 | f_s_dadda_pg_rca32_fa805_y3;
  assign f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_fa805_y4 = f_s_dadda_pg_rca32_fa805_y4;
  assign f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_fa225_y2 = f_s_dadda_pg_rca32_fa225_y2;
  assign f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_ha24_y0 = f_s_dadda_pg_rca32_ha24_y0;
  assign f_s_dadda_pg_rca32_fa806_y0 = f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_fa805_y4 ^ f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_fa225_y2;
  assign f_s_dadda_pg_rca32_fa806_y1 = f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_fa805_y4 & f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_fa225_y2;
  assign f_s_dadda_pg_rca32_fa806_y2 = f_s_dadda_pg_rca32_fa806_y0 ^ f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_ha24_y0;
  assign f_s_dadda_pg_rca32_fa806_y3 = f_s_dadda_pg_rca32_fa806_y0 & f_s_dadda_pg_rca32_fa806_f_s_dadda_pg_rca32_ha24_y0;
  assign f_s_dadda_pg_rca32_fa806_y4 = f_s_dadda_pg_rca32_fa806_y1 | f_s_dadda_pg_rca32_fa806_y3;
  assign f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_fa806_y4 = f_s_dadda_pg_rca32_fa806_y4;
  assign f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_fa246_y2 = f_s_dadda_pg_rca32_fa246_y2;
  assign f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_ha25_y0 = f_s_dadda_pg_rca32_ha25_y0;
  assign f_s_dadda_pg_rca32_fa807_y0 = f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_fa806_y4 ^ f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_fa246_y2;
  assign f_s_dadda_pg_rca32_fa807_y1 = f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_fa806_y4 & f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_fa246_y2;
  assign f_s_dadda_pg_rca32_fa807_y2 = f_s_dadda_pg_rca32_fa807_y0 ^ f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_ha25_y0;
  assign f_s_dadda_pg_rca32_fa807_y3 = f_s_dadda_pg_rca32_fa807_y0 & f_s_dadda_pg_rca32_fa807_f_s_dadda_pg_rca32_ha25_y0;
  assign f_s_dadda_pg_rca32_fa807_y4 = f_s_dadda_pg_rca32_fa807_y1 | f_s_dadda_pg_rca32_fa807_y3;
  assign f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa807_y4 = f_s_dadda_pg_rca32_fa807_y4;
  assign f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa267_y2 = f_s_dadda_pg_rca32_fa267_y2;
  assign f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa268_y2 = f_s_dadda_pg_rca32_fa268_y2;
  assign f_s_dadda_pg_rca32_fa808_y0 = f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa807_y4 ^ f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa267_y2;
  assign f_s_dadda_pg_rca32_fa808_y1 = f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa807_y4 & f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa267_y2;
  assign f_s_dadda_pg_rca32_fa808_y2 = f_s_dadda_pg_rca32_fa808_y0 ^ f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa268_y2;
  assign f_s_dadda_pg_rca32_fa808_y3 = f_s_dadda_pg_rca32_fa808_y0 & f_s_dadda_pg_rca32_fa808_f_s_dadda_pg_rca32_fa268_y2;
  assign f_s_dadda_pg_rca32_fa808_y4 = f_s_dadda_pg_rca32_fa808_y1 | f_s_dadda_pg_rca32_fa808_y3;
  assign f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa808_y4 = f_s_dadda_pg_rca32_fa808_y4;
  assign f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa289_y2 = f_s_dadda_pg_rca32_fa289_y2;
  assign f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa290_y2 = f_s_dadda_pg_rca32_fa290_y2;
  assign f_s_dadda_pg_rca32_fa809_y0 = f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa808_y4 ^ f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa289_y2;
  assign f_s_dadda_pg_rca32_fa809_y1 = f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa808_y4 & f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa289_y2;
  assign f_s_dadda_pg_rca32_fa809_y2 = f_s_dadda_pg_rca32_fa809_y0 ^ f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa290_y2;
  assign f_s_dadda_pg_rca32_fa809_y3 = f_s_dadda_pg_rca32_fa809_y0 & f_s_dadda_pg_rca32_fa809_f_s_dadda_pg_rca32_fa290_y2;
  assign f_s_dadda_pg_rca32_fa809_y4 = f_s_dadda_pg_rca32_fa809_y1 | f_s_dadda_pg_rca32_fa809_y3;
  assign f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa809_y4 = f_s_dadda_pg_rca32_fa809_y4;
  assign f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa311_y2 = f_s_dadda_pg_rca32_fa311_y2;
  assign f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa312_y2 = f_s_dadda_pg_rca32_fa312_y2;
  assign f_s_dadda_pg_rca32_fa810_y0 = f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa809_y4 ^ f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa311_y2;
  assign f_s_dadda_pg_rca32_fa810_y1 = f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa809_y4 & f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa311_y2;
  assign f_s_dadda_pg_rca32_fa810_y2 = f_s_dadda_pg_rca32_fa810_y0 ^ f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa312_y2;
  assign f_s_dadda_pg_rca32_fa810_y3 = f_s_dadda_pg_rca32_fa810_y0 & f_s_dadda_pg_rca32_fa810_f_s_dadda_pg_rca32_fa312_y2;
  assign f_s_dadda_pg_rca32_fa810_y4 = f_s_dadda_pg_rca32_fa810_y1 | f_s_dadda_pg_rca32_fa810_y3;
  assign f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa810_y4 = f_s_dadda_pg_rca32_fa810_y4;
  assign f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa333_y2 = f_s_dadda_pg_rca32_fa333_y2;
  assign f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa334_y2 = f_s_dadda_pg_rca32_fa334_y2;
  assign f_s_dadda_pg_rca32_fa811_y0 = f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa810_y4 ^ f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa333_y2;
  assign f_s_dadda_pg_rca32_fa811_y1 = f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa810_y4 & f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa333_y2;
  assign f_s_dadda_pg_rca32_fa811_y2 = f_s_dadda_pg_rca32_fa811_y0 ^ f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa334_y2;
  assign f_s_dadda_pg_rca32_fa811_y3 = f_s_dadda_pg_rca32_fa811_y0 & f_s_dadda_pg_rca32_fa811_f_s_dadda_pg_rca32_fa334_y2;
  assign f_s_dadda_pg_rca32_fa811_y4 = f_s_dadda_pg_rca32_fa811_y1 | f_s_dadda_pg_rca32_fa811_y3;
  assign f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa811_y4 = f_s_dadda_pg_rca32_fa811_y4;
  assign f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa355_y2 = f_s_dadda_pg_rca32_fa355_y2;
  assign f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa356_y2 = f_s_dadda_pg_rca32_fa356_y2;
  assign f_s_dadda_pg_rca32_fa812_y0 = f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa811_y4 ^ f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa355_y2;
  assign f_s_dadda_pg_rca32_fa812_y1 = f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa811_y4 & f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa355_y2;
  assign f_s_dadda_pg_rca32_fa812_y2 = f_s_dadda_pg_rca32_fa812_y0 ^ f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa356_y2;
  assign f_s_dadda_pg_rca32_fa812_y3 = f_s_dadda_pg_rca32_fa812_y0 & f_s_dadda_pg_rca32_fa812_f_s_dadda_pg_rca32_fa356_y2;
  assign f_s_dadda_pg_rca32_fa812_y4 = f_s_dadda_pg_rca32_fa812_y1 | f_s_dadda_pg_rca32_fa812_y3;
  assign f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa812_y4 = f_s_dadda_pg_rca32_fa812_y4;
  assign f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa377_y2 = f_s_dadda_pg_rca32_fa377_y2;
  assign f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa378_y2 = f_s_dadda_pg_rca32_fa378_y2;
  assign f_s_dadda_pg_rca32_fa813_y0 = f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa812_y4 ^ f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa377_y2;
  assign f_s_dadda_pg_rca32_fa813_y1 = f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa812_y4 & f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa377_y2;
  assign f_s_dadda_pg_rca32_fa813_y2 = f_s_dadda_pg_rca32_fa813_y0 ^ f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa378_y2;
  assign f_s_dadda_pg_rca32_fa813_y3 = f_s_dadda_pg_rca32_fa813_y0 & f_s_dadda_pg_rca32_fa813_f_s_dadda_pg_rca32_fa378_y2;
  assign f_s_dadda_pg_rca32_fa813_y4 = f_s_dadda_pg_rca32_fa813_y1 | f_s_dadda_pg_rca32_fa813_y3;
  assign f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa813_y4 = f_s_dadda_pg_rca32_fa813_y4;
  assign f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa399_y2 = f_s_dadda_pg_rca32_fa399_y2;
  assign f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa400_y2 = f_s_dadda_pg_rca32_fa400_y2;
  assign f_s_dadda_pg_rca32_fa814_y0 = f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa813_y4 ^ f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa399_y2;
  assign f_s_dadda_pg_rca32_fa814_y1 = f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa813_y4 & f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa399_y2;
  assign f_s_dadda_pg_rca32_fa814_y2 = f_s_dadda_pg_rca32_fa814_y0 ^ f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa400_y2;
  assign f_s_dadda_pg_rca32_fa814_y3 = f_s_dadda_pg_rca32_fa814_y0 & f_s_dadda_pg_rca32_fa814_f_s_dadda_pg_rca32_fa400_y2;
  assign f_s_dadda_pg_rca32_fa814_y4 = f_s_dadda_pg_rca32_fa814_y1 | f_s_dadda_pg_rca32_fa814_y3;
  assign f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa814_y4 = f_s_dadda_pg_rca32_fa814_y4;
  assign f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa421_y2 = f_s_dadda_pg_rca32_fa421_y2;
  assign f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa422_y2 = f_s_dadda_pg_rca32_fa422_y2;
  assign f_s_dadda_pg_rca32_fa815_y0 = f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa814_y4 ^ f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa421_y2;
  assign f_s_dadda_pg_rca32_fa815_y1 = f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa814_y4 & f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa421_y2;
  assign f_s_dadda_pg_rca32_fa815_y2 = f_s_dadda_pg_rca32_fa815_y0 ^ f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa422_y2;
  assign f_s_dadda_pg_rca32_fa815_y3 = f_s_dadda_pg_rca32_fa815_y0 & f_s_dadda_pg_rca32_fa815_f_s_dadda_pg_rca32_fa422_y2;
  assign f_s_dadda_pg_rca32_fa815_y4 = f_s_dadda_pg_rca32_fa815_y1 | f_s_dadda_pg_rca32_fa815_y3;
  assign f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa815_y4 = f_s_dadda_pg_rca32_fa815_y4;
  assign f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa443_y2 = f_s_dadda_pg_rca32_fa443_y2;
  assign f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa444_y2 = f_s_dadda_pg_rca32_fa444_y2;
  assign f_s_dadda_pg_rca32_fa816_y0 = f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa815_y4 ^ f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa443_y2;
  assign f_s_dadda_pg_rca32_fa816_y1 = f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa815_y4 & f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa443_y2;
  assign f_s_dadda_pg_rca32_fa816_y2 = f_s_dadda_pg_rca32_fa816_y0 ^ f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa444_y2;
  assign f_s_dadda_pg_rca32_fa816_y3 = f_s_dadda_pg_rca32_fa816_y0 & f_s_dadda_pg_rca32_fa816_f_s_dadda_pg_rca32_fa444_y2;
  assign f_s_dadda_pg_rca32_fa816_y4 = f_s_dadda_pg_rca32_fa816_y1 | f_s_dadda_pg_rca32_fa816_y3;
  assign f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa816_y4 = f_s_dadda_pg_rca32_fa816_y4;
  assign f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa464_y2 = f_s_dadda_pg_rca32_fa464_y2;
  assign f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa465_y2 = f_s_dadda_pg_rca32_fa465_y2;
  assign f_s_dadda_pg_rca32_fa817_y0 = f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa816_y4 ^ f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa464_y2;
  assign f_s_dadda_pg_rca32_fa817_y1 = f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa816_y4 & f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa464_y2;
  assign f_s_dadda_pg_rca32_fa817_y2 = f_s_dadda_pg_rca32_fa817_y0 ^ f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa465_y2;
  assign f_s_dadda_pg_rca32_fa817_y3 = f_s_dadda_pg_rca32_fa817_y0 & f_s_dadda_pg_rca32_fa817_f_s_dadda_pg_rca32_fa465_y2;
  assign f_s_dadda_pg_rca32_fa817_y4 = f_s_dadda_pg_rca32_fa817_y1 | f_s_dadda_pg_rca32_fa817_y3;
  assign f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa817_y4 = f_s_dadda_pg_rca32_fa817_y4;
  assign f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa484_y2 = f_s_dadda_pg_rca32_fa484_y2;
  assign f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa485_y2 = f_s_dadda_pg_rca32_fa485_y2;
  assign f_s_dadda_pg_rca32_fa818_y0 = f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa817_y4 ^ f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa484_y2;
  assign f_s_dadda_pg_rca32_fa818_y1 = f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa817_y4 & f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa484_y2;
  assign f_s_dadda_pg_rca32_fa818_y2 = f_s_dadda_pg_rca32_fa818_y0 ^ f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa485_y2;
  assign f_s_dadda_pg_rca32_fa818_y3 = f_s_dadda_pg_rca32_fa818_y0 & f_s_dadda_pg_rca32_fa818_f_s_dadda_pg_rca32_fa485_y2;
  assign f_s_dadda_pg_rca32_fa818_y4 = f_s_dadda_pg_rca32_fa818_y1 | f_s_dadda_pg_rca32_fa818_y3;
  assign f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa818_y4 = f_s_dadda_pg_rca32_fa818_y4;
  assign f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa503_y2 = f_s_dadda_pg_rca32_fa503_y2;
  assign f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa504_y2 = f_s_dadda_pg_rca32_fa504_y2;
  assign f_s_dadda_pg_rca32_fa819_y0 = f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa818_y4 ^ f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa503_y2;
  assign f_s_dadda_pg_rca32_fa819_y1 = f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa818_y4 & f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa503_y2;
  assign f_s_dadda_pg_rca32_fa819_y2 = f_s_dadda_pg_rca32_fa819_y0 ^ f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa504_y2;
  assign f_s_dadda_pg_rca32_fa819_y3 = f_s_dadda_pg_rca32_fa819_y0 & f_s_dadda_pg_rca32_fa819_f_s_dadda_pg_rca32_fa504_y2;
  assign f_s_dadda_pg_rca32_fa819_y4 = f_s_dadda_pg_rca32_fa819_y1 | f_s_dadda_pg_rca32_fa819_y3;
  assign f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa819_y4 = f_s_dadda_pg_rca32_fa819_y4;
  assign f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa521_y2 = f_s_dadda_pg_rca32_fa521_y2;
  assign f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa522_y2 = f_s_dadda_pg_rca32_fa522_y2;
  assign f_s_dadda_pg_rca32_fa820_y0 = f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa819_y4 ^ f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa521_y2;
  assign f_s_dadda_pg_rca32_fa820_y1 = f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa819_y4 & f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa521_y2;
  assign f_s_dadda_pg_rca32_fa820_y2 = f_s_dadda_pg_rca32_fa820_y0 ^ f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa522_y2;
  assign f_s_dadda_pg_rca32_fa820_y3 = f_s_dadda_pg_rca32_fa820_y0 & f_s_dadda_pg_rca32_fa820_f_s_dadda_pg_rca32_fa522_y2;
  assign f_s_dadda_pg_rca32_fa820_y4 = f_s_dadda_pg_rca32_fa820_y1 | f_s_dadda_pg_rca32_fa820_y3;
  assign f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa820_y4 = f_s_dadda_pg_rca32_fa820_y4;
  assign f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa538_y2 = f_s_dadda_pg_rca32_fa538_y2;
  assign f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa539_y2 = f_s_dadda_pg_rca32_fa539_y2;
  assign f_s_dadda_pg_rca32_fa821_y0 = f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa820_y4 ^ f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa538_y2;
  assign f_s_dadda_pg_rca32_fa821_y1 = f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa820_y4 & f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa538_y2;
  assign f_s_dadda_pg_rca32_fa821_y2 = f_s_dadda_pg_rca32_fa821_y0 ^ f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa539_y2;
  assign f_s_dadda_pg_rca32_fa821_y3 = f_s_dadda_pg_rca32_fa821_y0 & f_s_dadda_pg_rca32_fa821_f_s_dadda_pg_rca32_fa539_y2;
  assign f_s_dadda_pg_rca32_fa821_y4 = f_s_dadda_pg_rca32_fa821_y1 | f_s_dadda_pg_rca32_fa821_y3;
  assign f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa821_y4 = f_s_dadda_pg_rca32_fa821_y4;
  assign f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa554_y2 = f_s_dadda_pg_rca32_fa554_y2;
  assign f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa555_y2 = f_s_dadda_pg_rca32_fa555_y2;
  assign f_s_dadda_pg_rca32_fa822_y0 = f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa821_y4 ^ f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa554_y2;
  assign f_s_dadda_pg_rca32_fa822_y1 = f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa821_y4 & f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa554_y2;
  assign f_s_dadda_pg_rca32_fa822_y2 = f_s_dadda_pg_rca32_fa822_y0 ^ f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa555_y2;
  assign f_s_dadda_pg_rca32_fa822_y3 = f_s_dadda_pg_rca32_fa822_y0 & f_s_dadda_pg_rca32_fa822_f_s_dadda_pg_rca32_fa555_y2;
  assign f_s_dadda_pg_rca32_fa822_y4 = f_s_dadda_pg_rca32_fa822_y1 | f_s_dadda_pg_rca32_fa822_y3;
  assign f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa822_y4 = f_s_dadda_pg_rca32_fa822_y4;
  assign f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa569_y2 = f_s_dadda_pg_rca32_fa569_y2;
  assign f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa570_y2 = f_s_dadda_pg_rca32_fa570_y2;
  assign f_s_dadda_pg_rca32_fa823_y0 = f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa822_y4 ^ f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa569_y2;
  assign f_s_dadda_pg_rca32_fa823_y1 = f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa822_y4 & f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa569_y2;
  assign f_s_dadda_pg_rca32_fa823_y2 = f_s_dadda_pg_rca32_fa823_y0 ^ f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa570_y2;
  assign f_s_dadda_pg_rca32_fa823_y3 = f_s_dadda_pg_rca32_fa823_y0 & f_s_dadda_pg_rca32_fa823_f_s_dadda_pg_rca32_fa570_y2;
  assign f_s_dadda_pg_rca32_fa823_y4 = f_s_dadda_pg_rca32_fa823_y1 | f_s_dadda_pg_rca32_fa823_y3;
  assign f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa823_y4 = f_s_dadda_pg_rca32_fa823_y4;
  assign f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa583_y2 = f_s_dadda_pg_rca32_fa583_y2;
  assign f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa584_y2 = f_s_dadda_pg_rca32_fa584_y2;
  assign f_s_dadda_pg_rca32_fa824_y0 = f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa823_y4 ^ f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa583_y2;
  assign f_s_dadda_pg_rca32_fa824_y1 = f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa823_y4 & f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa583_y2;
  assign f_s_dadda_pg_rca32_fa824_y2 = f_s_dadda_pg_rca32_fa824_y0 ^ f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa584_y2;
  assign f_s_dadda_pg_rca32_fa824_y3 = f_s_dadda_pg_rca32_fa824_y0 & f_s_dadda_pg_rca32_fa824_f_s_dadda_pg_rca32_fa584_y2;
  assign f_s_dadda_pg_rca32_fa824_y4 = f_s_dadda_pg_rca32_fa824_y1 | f_s_dadda_pg_rca32_fa824_y3;
  assign f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa824_y4 = f_s_dadda_pg_rca32_fa824_y4;
  assign f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa596_y2 = f_s_dadda_pg_rca32_fa596_y2;
  assign f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa597_y2 = f_s_dadda_pg_rca32_fa597_y2;
  assign f_s_dadda_pg_rca32_fa825_y0 = f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa824_y4 ^ f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa596_y2;
  assign f_s_dadda_pg_rca32_fa825_y1 = f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa824_y4 & f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa596_y2;
  assign f_s_dadda_pg_rca32_fa825_y2 = f_s_dadda_pg_rca32_fa825_y0 ^ f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa597_y2;
  assign f_s_dadda_pg_rca32_fa825_y3 = f_s_dadda_pg_rca32_fa825_y0 & f_s_dadda_pg_rca32_fa825_f_s_dadda_pg_rca32_fa597_y2;
  assign f_s_dadda_pg_rca32_fa825_y4 = f_s_dadda_pg_rca32_fa825_y1 | f_s_dadda_pg_rca32_fa825_y3;
  assign f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa825_y4 = f_s_dadda_pg_rca32_fa825_y4;
  assign f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa608_y2 = f_s_dadda_pg_rca32_fa608_y2;
  assign f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa609_y2 = f_s_dadda_pg_rca32_fa609_y2;
  assign f_s_dadda_pg_rca32_fa826_y0 = f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa825_y4 ^ f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa608_y2;
  assign f_s_dadda_pg_rca32_fa826_y1 = f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa825_y4 & f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa608_y2;
  assign f_s_dadda_pg_rca32_fa826_y2 = f_s_dadda_pg_rca32_fa826_y0 ^ f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa609_y2;
  assign f_s_dadda_pg_rca32_fa826_y3 = f_s_dadda_pg_rca32_fa826_y0 & f_s_dadda_pg_rca32_fa826_f_s_dadda_pg_rca32_fa609_y2;
  assign f_s_dadda_pg_rca32_fa826_y4 = f_s_dadda_pg_rca32_fa826_y1 | f_s_dadda_pg_rca32_fa826_y3;
  assign f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa826_y4 = f_s_dadda_pg_rca32_fa826_y4;
  assign f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa619_y2 = f_s_dadda_pg_rca32_fa619_y2;
  assign f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa620_y2 = f_s_dadda_pg_rca32_fa620_y2;
  assign f_s_dadda_pg_rca32_fa827_y0 = f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa826_y4 ^ f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa619_y2;
  assign f_s_dadda_pg_rca32_fa827_y1 = f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa826_y4 & f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa619_y2;
  assign f_s_dadda_pg_rca32_fa827_y2 = f_s_dadda_pg_rca32_fa827_y0 ^ f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa620_y2;
  assign f_s_dadda_pg_rca32_fa827_y3 = f_s_dadda_pg_rca32_fa827_y0 & f_s_dadda_pg_rca32_fa827_f_s_dadda_pg_rca32_fa620_y2;
  assign f_s_dadda_pg_rca32_fa827_y4 = f_s_dadda_pg_rca32_fa827_y1 | f_s_dadda_pg_rca32_fa827_y3;
  assign f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa827_y4 = f_s_dadda_pg_rca32_fa827_y4;
  assign f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa629_y2 = f_s_dadda_pg_rca32_fa629_y2;
  assign f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa630_y2 = f_s_dadda_pg_rca32_fa630_y2;
  assign f_s_dadda_pg_rca32_fa828_y0 = f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa827_y4 ^ f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa629_y2;
  assign f_s_dadda_pg_rca32_fa828_y1 = f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa827_y4 & f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa629_y2;
  assign f_s_dadda_pg_rca32_fa828_y2 = f_s_dadda_pg_rca32_fa828_y0 ^ f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa630_y2;
  assign f_s_dadda_pg_rca32_fa828_y3 = f_s_dadda_pg_rca32_fa828_y0 & f_s_dadda_pg_rca32_fa828_f_s_dadda_pg_rca32_fa630_y2;
  assign f_s_dadda_pg_rca32_fa828_y4 = f_s_dadda_pg_rca32_fa828_y1 | f_s_dadda_pg_rca32_fa828_y3;
  assign f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa828_y4 = f_s_dadda_pg_rca32_fa828_y4;
  assign f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa638_y2 = f_s_dadda_pg_rca32_fa638_y2;
  assign f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa639_y2 = f_s_dadda_pg_rca32_fa639_y2;
  assign f_s_dadda_pg_rca32_fa829_y0 = f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa828_y4 ^ f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa638_y2;
  assign f_s_dadda_pg_rca32_fa829_y1 = f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa828_y4 & f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa638_y2;
  assign f_s_dadda_pg_rca32_fa829_y2 = f_s_dadda_pg_rca32_fa829_y0 ^ f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa639_y2;
  assign f_s_dadda_pg_rca32_fa829_y3 = f_s_dadda_pg_rca32_fa829_y0 & f_s_dadda_pg_rca32_fa829_f_s_dadda_pg_rca32_fa639_y2;
  assign f_s_dadda_pg_rca32_fa829_y4 = f_s_dadda_pg_rca32_fa829_y1 | f_s_dadda_pg_rca32_fa829_y3;
  assign f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa829_y4 = f_s_dadda_pg_rca32_fa829_y4;
  assign f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa646_y2 = f_s_dadda_pg_rca32_fa646_y2;
  assign f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa647_y2 = f_s_dadda_pg_rca32_fa647_y2;
  assign f_s_dadda_pg_rca32_fa830_y0 = f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa829_y4 ^ f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa646_y2;
  assign f_s_dadda_pg_rca32_fa830_y1 = f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa829_y4 & f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa646_y2;
  assign f_s_dadda_pg_rca32_fa830_y2 = f_s_dadda_pg_rca32_fa830_y0 ^ f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa647_y2;
  assign f_s_dadda_pg_rca32_fa830_y3 = f_s_dadda_pg_rca32_fa830_y0 & f_s_dadda_pg_rca32_fa830_f_s_dadda_pg_rca32_fa647_y2;
  assign f_s_dadda_pg_rca32_fa830_y4 = f_s_dadda_pg_rca32_fa830_y1 | f_s_dadda_pg_rca32_fa830_y3;
  assign f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa830_y4 = f_s_dadda_pg_rca32_fa830_y4;
  assign f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa653_y2 = f_s_dadda_pg_rca32_fa653_y2;
  assign f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa654_y2 = f_s_dadda_pg_rca32_fa654_y2;
  assign f_s_dadda_pg_rca32_fa831_y0 = f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa830_y4 ^ f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa653_y2;
  assign f_s_dadda_pg_rca32_fa831_y1 = f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa830_y4 & f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa653_y2;
  assign f_s_dadda_pg_rca32_fa831_y2 = f_s_dadda_pg_rca32_fa831_y0 ^ f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa654_y2;
  assign f_s_dadda_pg_rca32_fa831_y3 = f_s_dadda_pg_rca32_fa831_y0 & f_s_dadda_pg_rca32_fa831_f_s_dadda_pg_rca32_fa654_y2;
  assign f_s_dadda_pg_rca32_fa831_y4 = f_s_dadda_pg_rca32_fa831_y1 | f_s_dadda_pg_rca32_fa831_y3;
  assign f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa831_y4 = f_s_dadda_pg_rca32_fa831_y4;
  assign f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa659_y2 = f_s_dadda_pg_rca32_fa659_y2;
  assign f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa660_y2 = f_s_dadda_pg_rca32_fa660_y2;
  assign f_s_dadda_pg_rca32_fa832_y0 = f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa831_y4 ^ f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa659_y2;
  assign f_s_dadda_pg_rca32_fa832_y1 = f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa831_y4 & f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa659_y2;
  assign f_s_dadda_pg_rca32_fa832_y2 = f_s_dadda_pg_rca32_fa832_y0 ^ f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa660_y2;
  assign f_s_dadda_pg_rca32_fa832_y3 = f_s_dadda_pg_rca32_fa832_y0 & f_s_dadda_pg_rca32_fa832_f_s_dadda_pg_rca32_fa660_y2;
  assign f_s_dadda_pg_rca32_fa832_y4 = f_s_dadda_pg_rca32_fa832_y1 | f_s_dadda_pg_rca32_fa832_y3;
  assign f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa832_y4 = f_s_dadda_pg_rca32_fa832_y4;
  assign f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa664_y2 = f_s_dadda_pg_rca32_fa664_y2;
  assign f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa665_y2 = f_s_dadda_pg_rca32_fa665_y2;
  assign f_s_dadda_pg_rca32_fa833_y0 = f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa832_y4 ^ f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa664_y2;
  assign f_s_dadda_pg_rca32_fa833_y1 = f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa832_y4 & f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa664_y2;
  assign f_s_dadda_pg_rca32_fa833_y2 = f_s_dadda_pg_rca32_fa833_y0 ^ f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa665_y2;
  assign f_s_dadda_pg_rca32_fa833_y3 = f_s_dadda_pg_rca32_fa833_y0 & f_s_dadda_pg_rca32_fa833_f_s_dadda_pg_rca32_fa665_y2;
  assign f_s_dadda_pg_rca32_fa833_y4 = f_s_dadda_pg_rca32_fa833_y1 | f_s_dadda_pg_rca32_fa833_y3;
  assign f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa833_y4 = f_s_dadda_pg_rca32_fa833_y4;
  assign f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa668_y2 = f_s_dadda_pg_rca32_fa668_y2;
  assign f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa669_y2 = f_s_dadda_pg_rca32_fa669_y2;
  assign f_s_dadda_pg_rca32_fa834_y0 = f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa833_y4 ^ f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa668_y2;
  assign f_s_dadda_pg_rca32_fa834_y1 = f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa833_y4 & f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa668_y2;
  assign f_s_dadda_pg_rca32_fa834_y2 = f_s_dadda_pg_rca32_fa834_y0 ^ f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa669_y2;
  assign f_s_dadda_pg_rca32_fa834_y3 = f_s_dadda_pg_rca32_fa834_y0 & f_s_dadda_pg_rca32_fa834_f_s_dadda_pg_rca32_fa669_y2;
  assign f_s_dadda_pg_rca32_fa834_y4 = f_s_dadda_pg_rca32_fa834_y1 | f_s_dadda_pg_rca32_fa834_y3;
  assign f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa834_y4 = f_s_dadda_pg_rca32_fa834_y4;
  assign f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa671_y2 = f_s_dadda_pg_rca32_fa671_y2;
  assign f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa672_y2 = f_s_dadda_pg_rca32_fa672_y2;
  assign f_s_dadda_pg_rca32_fa835_y0 = f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa834_y4 ^ f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa671_y2;
  assign f_s_dadda_pg_rca32_fa835_y1 = f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa834_y4 & f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa671_y2;
  assign f_s_dadda_pg_rca32_fa835_y2 = f_s_dadda_pg_rca32_fa835_y0 ^ f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa672_y2;
  assign f_s_dadda_pg_rca32_fa835_y3 = f_s_dadda_pg_rca32_fa835_y0 & f_s_dadda_pg_rca32_fa835_f_s_dadda_pg_rca32_fa672_y2;
  assign f_s_dadda_pg_rca32_fa835_y4 = f_s_dadda_pg_rca32_fa835_y1 | f_s_dadda_pg_rca32_fa835_y3;
  assign f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa835_y4 = f_s_dadda_pg_rca32_fa835_y4;
  assign f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa673_y2 = f_s_dadda_pg_rca32_fa673_y2;
  assign f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa674_y2 = f_s_dadda_pg_rca32_fa674_y2;
  assign f_s_dadda_pg_rca32_fa836_y0 = f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa835_y4 ^ f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa673_y2;
  assign f_s_dadda_pg_rca32_fa836_y1 = f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa835_y4 & f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa673_y2;
  assign f_s_dadda_pg_rca32_fa836_y2 = f_s_dadda_pg_rca32_fa836_y0 ^ f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa674_y2;
  assign f_s_dadda_pg_rca32_fa836_y3 = f_s_dadda_pg_rca32_fa836_y0 & f_s_dadda_pg_rca32_fa836_f_s_dadda_pg_rca32_fa674_y2;
  assign f_s_dadda_pg_rca32_fa836_y4 = f_s_dadda_pg_rca32_fa836_y1 | f_s_dadda_pg_rca32_fa836_y3;
  assign f_s_dadda_pg_rca32_nand_26_31_a_26 = a_26;
  assign f_s_dadda_pg_rca32_nand_26_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_26_31_y0 = ~(f_s_dadda_pg_rca32_nand_26_31_a_26 & f_s_dadda_pg_rca32_nand_26_31_b_31);
  assign f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_fa836_y4 = f_s_dadda_pg_rca32_fa836_y4;
  assign f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_nand_26_31_y0 = f_s_dadda_pg_rca32_nand_26_31_y0;
  assign f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_fa675_y2 = f_s_dadda_pg_rca32_fa675_y2;
  assign f_s_dadda_pg_rca32_fa837_y0 = f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_fa836_y4 ^ f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_nand_26_31_y0;
  assign f_s_dadda_pg_rca32_fa837_y1 = f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_fa836_y4 & f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_nand_26_31_y0;
  assign f_s_dadda_pg_rca32_fa837_y2 = f_s_dadda_pg_rca32_fa837_y0 ^ f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_fa675_y2;
  assign f_s_dadda_pg_rca32_fa837_y3 = f_s_dadda_pg_rca32_fa837_y0 & f_s_dadda_pg_rca32_fa837_f_s_dadda_pg_rca32_fa675_y2;
  assign f_s_dadda_pg_rca32_fa837_y4 = f_s_dadda_pg_rca32_fa837_y1 | f_s_dadda_pg_rca32_fa837_y3;
  assign f_s_dadda_pg_rca32_and_28_30_a_28 = a_28;
  assign f_s_dadda_pg_rca32_and_28_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_28_30_y0 = f_s_dadda_pg_rca32_and_28_30_a_28 & f_s_dadda_pg_rca32_and_28_30_b_30;
  assign f_s_dadda_pg_rca32_nand_27_31_a_27 = a_27;
  assign f_s_dadda_pg_rca32_nand_27_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_27_31_y0 = ~(f_s_dadda_pg_rca32_nand_27_31_a_27 & f_s_dadda_pg_rca32_nand_27_31_b_31);
  assign f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_fa837_y4 = f_s_dadda_pg_rca32_fa837_y4;
  assign f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_and_28_30_y0 = f_s_dadda_pg_rca32_and_28_30_y0;
  assign f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_nand_27_31_y0 = f_s_dadda_pg_rca32_nand_27_31_y0;
  assign f_s_dadda_pg_rca32_fa838_y0 = f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_fa837_y4 ^ f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_and_28_30_y0;
  assign f_s_dadda_pg_rca32_fa838_y1 = f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_fa837_y4 & f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_and_28_30_y0;
  assign f_s_dadda_pg_rca32_fa838_y2 = f_s_dadda_pg_rca32_fa838_y0 ^ f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_nand_27_31_y0;
  assign f_s_dadda_pg_rca32_fa838_y3 = f_s_dadda_pg_rca32_fa838_y0 & f_s_dadda_pg_rca32_fa838_f_s_dadda_pg_rca32_nand_27_31_y0;
  assign f_s_dadda_pg_rca32_fa838_y4 = f_s_dadda_pg_rca32_fa838_y1 | f_s_dadda_pg_rca32_fa838_y3;
  assign f_s_dadda_pg_rca32_and_30_29_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_and_30_29_y0 = f_s_dadda_pg_rca32_and_30_29_a_30 & f_s_dadda_pg_rca32_and_30_29_b_29;
  assign f_s_dadda_pg_rca32_and_29_30_a_29 = a_29;
  assign f_s_dadda_pg_rca32_and_29_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_29_30_y0 = f_s_dadda_pg_rca32_and_29_30_a_29 & f_s_dadda_pg_rca32_and_29_30_b_30;
  assign f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_fa838_y4 = f_s_dadda_pg_rca32_fa838_y4;
  assign f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_and_30_29_y0 = f_s_dadda_pg_rca32_and_30_29_y0;
  assign f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_and_29_30_y0 = f_s_dadda_pg_rca32_and_29_30_y0;
  assign f_s_dadda_pg_rca32_fa839_y0 = f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_fa838_y4 ^ f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_and_30_29_y0;
  assign f_s_dadda_pg_rca32_fa839_y1 = f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_fa838_y4 & f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_and_30_29_y0;
  assign f_s_dadda_pg_rca32_fa839_y2 = f_s_dadda_pg_rca32_fa839_y0 ^ f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_and_29_30_y0;
  assign f_s_dadda_pg_rca32_fa839_y3 = f_s_dadda_pg_rca32_fa839_y0 & f_s_dadda_pg_rca32_fa839_f_s_dadda_pg_rca32_and_29_30_y0;
  assign f_s_dadda_pg_rca32_fa839_y4 = f_s_dadda_pg_rca32_fa839_y1 | f_s_dadda_pg_rca32_fa839_y3;
  assign f_s_dadda_pg_rca32_nand_31_29_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_29_b_29 = b_29;
  assign f_s_dadda_pg_rca32_nand_31_29_y0 = ~(f_s_dadda_pg_rca32_nand_31_29_a_31 & f_s_dadda_pg_rca32_nand_31_29_b_29);
  assign f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_fa839_y4 = f_s_dadda_pg_rca32_fa839_y4;
  assign f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_fa783_y4 = f_s_dadda_pg_rca32_fa783_y4;
  assign f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_nand_31_29_y0 = f_s_dadda_pg_rca32_nand_31_29_y0;
  assign f_s_dadda_pg_rca32_fa840_y0 = f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_fa839_y4 ^ f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_fa783_y4;
  assign f_s_dadda_pg_rca32_fa840_y1 = f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_fa839_y4 & f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_fa783_y4;
  assign f_s_dadda_pg_rca32_fa840_y2 = f_s_dadda_pg_rca32_fa840_y0 ^ f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_nand_31_29_y0;
  assign f_s_dadda_pg_rca32_fa840_y3 = f_s_dadda_pg_rca32_fa840_y0 & f_s_dadda_pg_rca32_fa840_f_s_dadda_pg_rca32_nand_31_29_y0;
  assign f_s_dadda_pg_rca32_fa840_y4 = f_s_dadda_pg_rca32_fa840_y1 | f_s_dadda_pg_rca32_fa840_y3;
  assign f_s_dadda_pg_rca32_and_2_0_a_2 = a_2;
  assign f_s_dadda_pg_rca32_and_2_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_2_0_y0 = f_s_dadda_pg_rca32_and_2_0_a_2 & f_s_dadda_pg_rca32_and_2_0_b_0;
  assign f_s_dadda_pg_rca32_and_1_1_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_1_1_y0 = f_s_dadda_pg_rca32_and_1_1_a_1 & f_s_dadda_pg_rca32_and_1_1_b_1;
  assign f_s_dadda_pg_rca32_ha29_f_s_dadda_pg_rca32_and_2_0_y0 = f_s_dadda_pg_rca32_and_2_0_y0;
  assign f_s_dadda_pg_rca32_ha29_f_s_dadda_pg_rca32_and_1_1_y0 = f_s_dadda_pg_rca32_and_1_1_y0;
  assign f_s_dadda_pg_rca32_ha29_y0 = f_s_dadda_pg_rca32_ha29_f_s_dadda_pg_rca32_and_2_0_y0 ^ f_s_dadda_pg_rca32_ha29_f_s_dadda_pg_rca32_and_1_1_y0;
  assign f_s_dadda_pg_rca32_ha29_y1 = f_s_dadda_pg_rca32_ha29_f_s_dadda_pg_rca32_and_2_0_y0 & f_s_dadda_pg_rca32_ha29_f_s_dadda_pg_rca32_and_1_1_y0;
  assign f_s_dadda_pg_rca32_and_1_2_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_1_2_y0 = f_s_dadda_pg_rca32_and_1_2_a_1 & f_s_dadda_pg_rca32_and_1_2_b_2;
  assign f_s_dadda_pg_rca32_and_0_3_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_3_b_3 = b_3;
  assign f_s_dadda_pg_rca32_and_0_3_y0 = f_s_dadda_pg_rca32_and_0_3_a_0 & f_s_dadda_pg_rca32_and_0_3_b_3;
  assign f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_ha29_y1 = f_s_dadda_pg_rca32_ha29_y1;
  assign f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_and_1_2_y0 = f_s_dadda_pg_rca32_and_1_2_y0;
  assign f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_and_0_3_y0 = f_s_dadda_pg_rca32_and_0_3_y0;
  assign f_s_dadda_pg_rca32_fa841_y0 = f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_ha29_y1 ^ f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_and_1_2_y0;
  assign f_s_dadda_pg_rca32_fa841_y1 = f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_ha29_y1 & f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_and_1_2_y0;
  assign f_s_dadda_pg_rca32_fa841_y2 = f_s_dadda_pg_rca32_fa841_y0 ^ f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_and_0_3_y0;
  assign f_s_dadda_pg_rca32_fa841_y3 = f_s_dadda_pg_rca32_fa841_y0 & f_s_dadda_pg_rca32_fa841_f_s_dadda_pg_rca32_and_0_3_y0;
  assign f_s_dadda_pg_rca32_fa841_y4 = f_s_dadda_pg_rca32_fa841_y1 | f_s_dadda_pg_rca32_fa841_y3;
  assign f_s_dadda_pg_rca32_and_0_4_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_4_b_4 = b_4;
  assign f_s_dadda_pg_rca32_and_0_4_y0 = f_s_dadda_pg_rca32_and_0_4_a_0 & f_s_dadda_pg_rca32_and_0_4_b_4;
  assign f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_fa841_y4 = f_s_dadda_pg_rca32_fa841_y4;
  assign f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_and_0_4_y0 = f_s_dadda_pg_rca32_and_0_4_y0;
  assign f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_ha26_y0 = f_s_dadda_pg_rca32_ha26_y0;
  assign f_s_dadda_pg_rca32_fa842_y0 = f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_fa841_y4 ^ f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_and_0_4_y0;
  assign f_s_dadda_pg_rca32_fa842_y1 = f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_fa841_y4 & f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_and_0_4_y0;
  assign f_s_dadda_pg_rca32_fa842_y2 = f_s_dadda_pg_rca32_fa842_y0 ^ f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_ha26_y0;
  assign f_s_dadda_pg_rca32_fa842_y3 = f_s_dadda_pg_rca32_fa842_y0 & f_s_dadda_pg_rca32_fa842_f_s_dadda_pg_rca32_ha26_y0;
  assign f_s_dadda_pg_rca32_fa842_y4 = f_s_dadda_pg_rca32_fa842_y1 | f_s_dadda_pg_rca32_fa842_y3;
  assign f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_fa842_y4 = f_s_dadda_pg_rca32_fa842_y4;
  assign f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_fa676_y2 = f_s_dadda_pg_rca32_fa676_y2;
  assign f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_ha27_y0 = f_s_dadda_pg_rca32_ha27_y0;
  assign f_s_dadda_pg_rca32_fa843_y0 = f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_fa842_y4 ^ f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_fa676_y2;
  assign f_s_dadda_pg_rca32_fa843_y1 = f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_fa842_y4 & f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_fa676_y2;
  assign f_s_dadda_pg_rca32_fa843_y2 = f_s_dadda_pg_rca32_fa843_y0 ^ f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_ha27_y0;
  assign f_s_dadda_pg_rca32_fa843_y3 = f_s_dadda_pg_rca32_fa843_y0 & f_s_dadda_pg_rca32_fa843_f_s_dadda_pg_rca32_ha27_y0;
  assign f_s_dadda_pg_rca32_fa843_y4 = f_s_dadda_pg_rca32_fa843_y1 | f_s_dadda_pg_rca32_fa843_y3;
  assign f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa843_y4 = f_s_dadda_pg_rca32_fa843_y4;
  assign f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa677_y2 = f_s_dadda_pg_rca32_fa677_y2;
  assign f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa678_y2 = f_s_dadda_pg_rca32_fa678_y2;
  assign f_s_dadda_pg_rca32_fa844_y0 = f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa843_y4 ^ f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa677_y2;
  assign f_s_dadda_pg_rca32_fa844_y1 = f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa843_y4 & f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa677_y2;
  assign f_s_dadda_pg_rca32_fa844_y2 = f_s_dadda_pg_rca32_fa844_y0 ^ f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa678_y2;
  assign f_s_dadda_pg_rca32_fa844_y3 = f_s_dadda_pg_rca32_fa844_y0 & f_s_dadda_pg_rca32_fa844_f_s_dadda_pg_rca32_fa678_y2;
  assign f_s_dadda_pg_rca32_fa844_y4 = f_s_dadda_pg_rca32_fa844_y1 | f_s_dadda_pg_rca32_fa844_y3;
  assign f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa844_y4 = f_s_dadda_pg_rca32_fa844_y4;
  assign f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa679_y2 = f_s_dadda_pg_rca32_fa679_y2;
  assign f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa680_y2 = f_s_dadda_pg_rca32_fa680_y2;
  assign f_s_dadda_pg_rca32_fa845_y0 = f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa844_y4 ^ f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa679_y2;
  assign f_s_dadda_pg_rca32_fa845_y1 = f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa844_y4 & f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa679_y2;
  assign f_s_dadda_pg_rca32_fa845_y2 = f_s_dadda_pg_rca32_fa845_y0 ^ f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa680_y2;
  assign f_s_dadda_pg_rca32_fa845_y3 = f_s_dadda_pg_rca32_fa845_y0 & f_s_dadda_pg_rca32_fa845_f_s_dadda_pg_rca32_fa680_y2;
  assign f_s_dadda_pg_rca32_fa845_y4 = f_s_dadda_pg_rca32_fa845_y1 | f_s_dadda_pg_rca32_fa845_y3;
  assign f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa845_y4 = f_s_dadda_pg_rca32_fa845_y4;
  assign f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa681_y2 = f_s_dadda_pg_rca32_fa681_y2;
  assign f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa682_y2 = f_s_dadda_pg_rca32_fa682_y2;
  assign f_s_dadda_pg_rca32_fa846_y0 = f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa845_y4 ^ f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa681_y2;
  assign f_s_dadda_pg_rca32_fa846_y1 = f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa845_y4 & f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa681_y2;
  assign f_s_dadda_pg_rca32_fa846_y2 = f_s_dadda_pg_rca32_fa846_y0 ^ f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa682_y2;
  assign f_s_dadda_pg_rca32_fa846_y3 = f_s_dadda_pg_rca32_fa846_y0 & f_s_dadda_pg_rca32_fa846_f_s_dadda_pg_rca32_fa682_y2;
  assign f_s_dadda_pg_rca32_fa846_y4 = f_s_dadda_pg_rca32_fa846_y1 | f_s_dadda_pg_rca32_fa846_y3;
  assign f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa846_y4 = f_s_dadda_pg_rca32_fa846_y4;
  assign f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa683_y2 = f_s_dadda_pg_rca32_fa683_y2;
  assign f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa684_y2 = f_s_dadda_pg_rca32_fa684_y2;
  assign f_s_dadda_pg_rca32_fa847_y0 = f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa846_y4 ^ f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa683_y2;
  assign f_s_dadda_pg_rca32_fa847_y1 = f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa846_y4 & f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa683_y2;
  assign f_s_dadda_pg_rca32_fa847_y2 = f_s_dadda_pg_rca32_fa847_y0 ^ f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa684_y2;
  assign f_s_dadda_pg_rca32_fa847_y3 = f_s_dadda_pg_rca32_fa847_y0 & f_s_dadda_pg_rca32_fa847_f_s_dadda_pg_rca32_fa684_y2;
  assign f_s_dadda_pg_rca32_fa847_y4 = f_s_dadda_pg_rca32_fa847_y1 | f_s_dadda_pg_rca32_fa847_y3;
  assign f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa847_y4 = f_s_dadda_pg_rca32_fa847_y4;
  assign f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa685_y2 = f_s_dadda_pg_rca32_fa685_y2;
  assign f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa686_y2 = f_s_dadda_pg_rca32_fa686_y2;
  assign f_s_dadda_pg_rca32_fa848_y0 = f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa847_y4 ^ f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa685_y2;
  assign f_s_dadda_pg_rca32_fa848_y1 = f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa847_y4 & f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa685_y2;
  assign f_s_dadda_pg_rca32_fa848_y2 = f_s_dadda_pg_rca32_fa848_y0 ^ f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa686_y2;
  assign f_s_dadda_pg_rca32_fa848_y3 = f_s_dadda_pg_rca32_fa848_y0 & f_s_dadda_pg_rca32_fa848_f_s_dadda_pg_rca32_fa686_y2;
  assign f_s_dadda_pg_rca32_fa848_y4 = f_s_dadda_pg_rca32_fa848_y1 | f_s_dadda_pg_rca32_fa848_y3;
  assign f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa848_y4 = f_s_dadda_pg_rca32_fa848_y4;
  assign f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa687_y2 = f_s_dadda_pg_rca32_fa687_y2;
  assign f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa688_y2 = f_s_dadda_pg_rca32_fa688_y2;
  assign f_s_dadda_pg_rca32_fa849_y0 = f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa848_y4 ^ f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa687_y2;
  assign f_s_dadda_pg_rca32_fa849_y1 = f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa848_y4 & f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa687_y2;
  assign f_s_dadda_pg_rca32_fa849_y2 = f_s_dadda_pg_rca32_fa849_y0 ^ f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa688_y2;
  assign f_s_dadda_pg_rca32_fa849_y3 = f_s_dadda_pg_rca32_fa849_y0 & f_s_dadda_pg_rca32_fa849_f_s_dadda_pg_rca32_fa688_y2;
  assign f_s_dadda_pg_rca32_fa849_y4 = f_s_dadda_pg_rca32_fa849_y1 | f_s_dadda_pg_rca32_fa849_y3;
  assign f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa849_y4 = f_s_dadda_pg_rca32_fa849_y4;
  assign f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa689_y2 = f_s_dadda_pg_rca32_fa689_y2;
  assign f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa690_y2 = f_s_dadda_pg_rca32_fa690_y2;
  assign f_s_dadda_pg_rca32_fa850_y0 = f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa849_y4 ^ f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa689_y2;
  assign f_s_dadda_pg_rca32_fa850_y1 = f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa849_y4 & f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa689_y2;
  assign f_s_dadda_pg_rca32_fa850_y2 = f_s_dadda_pg_rca32_fa850_y0 ^ f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa690_y2;
  assign f_s_dadda_pg_rca32_fa850_y3 = f_s_dadda_pg_rca32_fa850_y0 & f_s_dadda_pg_rca32_fa850_f_s_dadda_pg_rca32_fa690_y2;
  assign f_s_dadda_pg_rca32_fa850_y4 = f_s_dadda_pg_rca32_fa850_y1 | f_s_dadda_pg_rca32_fa850_y3;
  assign f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa850_y4 = f_s_dadda_pg_rca32_fa850_y4;
  assign f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa691_y2 = f_s_dadda_pg_rca32_fa691_y2;
  assign f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa692_y2 = f_s_dadda_pg_rca32_fa692_y2;
  assign f_s_dadda_pg_rca32_fa851_y0 = f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa850_y4 ^ f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa691_y2;
  assign f_s_dadda_pg_rca32_fa851_y1 = f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa850_y4 & f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa691_y2;
  assign f_s_dadda_pg_rca32_fa851_y2 = f_s_dadda_pg_rca32_fa851_y0 ^ f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa692_y2;
  assign f_s_dadda_pg_rca32_fa851_y3 = f_s_dadda_pg_rca32_fa851_y0 & f_s_dadda_pg_rca32_fa851_f_s_dadda_pg_rca32_fa692_y2;
  assign f_s_dadda_pg_rca32_fa851_y4 = f_s_dadda_pg_rca32_fa851_y1 | f_s_dadda_pg_rca32_fa851_y3;
  assign f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa851_y4 = f_s_dadda_pg_rca32_fa851_y4;
  assign f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa693_y2 = f_s_dadda_pg_rca32_fa693_y2;
  assign f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa694_y2 = f_s_dadda_pg_rca32_fa694_y2;
  assign f_s_dadda_pg_rca32_fa852_y0 = f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa851_y4 ^ f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa693_y2;
  assign f_s_dadda_pg_rca32_fa852_y1 = f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa851_y4 & f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa693_y2;
  assign f_s_dadda_pg_rca32_fa852_y2 = f_s_dadda_pg_rca32_fa852_y0 ^ f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa694_y2;
  assign f_s_dadda_pg_rca32_fa852_y3 = f_s_dadda_pg_rca32_fa852_y0 & f_s_dadda_pg_rca32_fa852_f_s_dadda_pg_rca32_fa694_y2;
  assign f_s_dadda_pg_rca32_fa852_y4 = f_s_dadda_pg_rca32_fa852_y1 | f_s_dadda_pg_rca32_fa852_y3;
  assign f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa852_y4 = f_s_dadda_pg_rca32_fa852_y4;
  assign f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa695_y2 = f_s_dadda_pg_rca32_fa695_y2;
  assign f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa696_y2 = f_s_dadda_pg_rca32_fa696_y2;
  assign f_s_dadda_pg_rca32_fa853_y0 = f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa852_y4 ^ f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa695_y2;
  assign f_s_dadda_pg_rca32_fa853_y1 = f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa852_y4 & f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa695_y2;
  assign f_s_dadda_pg_rca32_fa853_y2 = f_s_dadda_pg_rca32_fa853_y0 ^ f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa696_y2;
  assign f_s_dadda_pg_rca32_fa853_y3 = f_s_dadda_pg_rca32_fa853_y0 & f_s_dadda_pg_rca32_fa853_f_s_dadda_pg_rca32_fa696_y2;
  assign f_s_dadda_pg_rca32_fa853_y4 = f_s_dadda_pg_rca32_fa853_y1 | f_s_dadda_pg_rca32_fa853_y3;
  assign f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa853_y4 = f_s_dadda_pg_rca32_fa853_y4;
  assign f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa697_y2 = f_s_dadda_pg_rca32_fa697_y2;
  assign f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa698_y2 = f_s_dadda_pg_rca32_fa698_y2;
  assign f_s_dadda_pg_rca32_fa854_y0 = f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa853_y4 ^ f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa697_y2;
  assign f_s_dadda_pg_rca32_fa854_y1 = f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa853_y4 & f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa697_y2;
  assign f_s_dadda_pg_rca32_fa854_y2 = f_s_dadda_pg_rca32_fa854_y0 ^ f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa698_y2;
  assign f_s_dadda_pg_rca32_fa854_y3 = f_s_dadda_pg_rca32_fa854_y0 & f_s_dadda_pg_rca32_fa854_f_s_dadda_pg_rca32_fa698_y2;
  assign f_s_dadda_pg_rca32_fa854_y4 = f_s_dadda_pg_rca32_fa854_y1 | f_s_dadda_pg_rca32_fa854_y3;
  assign f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa854_y4 = f_s_dadda_pg_rca32_fa854_y4;
  assign f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa699_y2 = f_s_dadda_pg_rca32_fa699_y2;
  assign f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa700_y2 = f_s_dadda_pg_rca32_fa700_y2;
  assign f_s_dadda_pg_rca32_fa855_y0 = f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa854_y4 ^ f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa699_y2;
  assign f_s_dadda_pg_rca32_fa855_y1 = f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa854_y4 & f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa699_y2;
  assign f_s_dadda_pg_rca32_fa855_y2 = f_s_dadda_pg_rca32_fa855_y0 ^ f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa700_y2;
  assign f_s_dadda_pg_rca32_fa855_y3 = f_s_dadda_pg_rca32_fa855_y0 & f_s_dadda_pg_rca32_fa855_f_s_dadda_pg_rca32_fa700_y2;
  assign f_s_dadda_pg_rca32_fa855_y4 = f_s_dadda_pg_rca32_fa855_y1 | f_s_dadda_pg_rca32_fa855_y3;
  assign f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa855_y4 = f_s_dadda_pg_rca32_fa855_y4;
  assign f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa701_y2 = f_s_dadda_pg_rca32_fa701_y2;
  assign f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa702_y2 = f_s_dadda_pg_rca32_fa702_y2;
  assign f_s_dadda_pg_rca32_fa856_y0 = f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa855_y4 ^ f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa701_y2;
  assign f_s_dadda_pg_rca32_fa856_y1 = f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa855_y4 & f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa701_y2;
  assign f_s_dadda_pg_rca32_fa856_y2 = f_s_dadda_pg_rca32_fa856_y0 ^ f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa702_y2;
  assign f_s_dadda_pg_rca32_fa856_y3 = f_s_dadda_pg_rca32_fa856_y0 & f_s_dadda_pg_rca32_fa856_f_s_dadda_pg_rca32_fa702_y2;
  assign f_s_dadda_pg_rca32_fa856_y4 = f_s_dadda_pg_rca32_fa856_y1 | f_s_dadda_pg_rca32_fa856_y3;
  assign f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa856_y4 = f_s_dadda_pg_rca32_fa856_y4;
  assign f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa703_y2 = f_s_dadda_pg_rca32_fa703_y2;
  assign f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa704_y2 = f_s_dadda_pg_rca32_fa704_y2;
  assign f_s_dadda_pg_rca32_fa857_y0 = f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa856_y4 ^ f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa703_y2;
  assign f_s_dadda_pg_rca32_fa857_y1 = f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa856_y4 & f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa703_y2;
  assign f_s_dadda_pg_rca32_fa857_y2 = f_s_dadda_pg_rca32_fa857_y0 ^ f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa704_y2;
  assign f_s_dadda_pg_rca32_fa857_y3 = f_s_dadda_pg_rca32_fa857_y0 & f_s_dadda_pg_rca32_fa857_f_s_dadda_pg_rca32_fa704_y2;
  assign f_s_dadda_pg_rca32_fa857_y4 = f_s_dadda_pg_rca32_fa857_y1 | f_s_dadda_pg_rca32_fa857_y3;
  assign f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa857_y4 = f_s_dadda_pg_rca32_fa857_y4;
  assign f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa705_y2 = f_s_dadda_pg_rca32_fa705_y2;
  assign f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa706_y2 = f_s_dadda_pg_rca32_fa706_y2;
  assign f_s_dadda_pg_rca32_fa858_y0 = f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa857_y4 ^ f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa705_y2;
  assign f_s_dadda_pg_rca32_fa858_y1 = f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa857_y4 & f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa705_y2;
  assign f_s_dadda_pg_rca32_fa858_y2 = f_s_dadda_pg_rca32_fa858_y0 ^ f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa706_y2;
  assign f_s_dadda_pg_rca32_fa858_y3 = f_s_dadda_pg_rca32_fa858_y0 & f_s_dadda_pg_rca32_fa858_f_s_dadda_pg_rca32_fa706_y2;
  assign f_s_dadda_pg_rca32_fa858_y4 = f_s_dadda_pg_rca32_fa858_y1 | f_s_dadda_pg_rca32_fa858_y3;
  assign f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa858_y4 = f_s_dadda_pg_rca32_fa858_y4;
  assign f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa707_y2 = f_s_dadda_pg_rca32_fa707_y2;
  assign f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa708_y2 = f_s_dadda_pg_rca32_fa708_y2;
  assign f_s_dadda_pg_rca32_fa859_y0 = f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa858_y4 ^ f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa707_y2;
  assign f_s_dadda_pg_rca32_fa859_y1 = f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa858_y4 & f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa707_y2;
  assign f_s_dadda_pg_rca32_fa859_y2 = f_s_dadda_pg_rca32_fa859_y0 ^ f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa708_y2;
  assign f_s_dadda_pg_rca32_fa859_y3 = f_s_dadda_pg_rca32_fa859_y0 & f_s_dadda_pg_rca32_fa859_f_s_dadda_pg_rca32_fa708_y2;
  assign f_s_dadda_pg_rca32_fa859_y4 = f_s_dadda_pg_rca32_fa859_y1 | f_s_dadda_pg_rca32_fa859_y3;
  assign f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa859_y4 = f_s_dadda_pg_rca32_fa859_y4;
  assign f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa709_y2 = f_s_dadda_pg_rca32_fa709_y2;
  assign f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa710_y2 = f_s_dadda_pg_rca32_fa710_y2;
  assign f_s_dadda_pg_rca32_fa860_y0 = f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa859_y4 ^ f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa709_y2;
  assign f_s_dadda_pg_rca32_fa860_y1 = f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa859_y4 & f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa709_y2;
  assign f_s_dadda_pg_rca32_fa860_y2 = f_s_dadda_pg_rca32_fa860_y0 ^ f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa710_y2;
  assign f_s_dadda_pg_rca32_fa860_y3 = f_s_dadda_pg_rca32_fa860_y0 & f_s_dadda_pg_rca32_fa860_f_s_dadda_pg_rca32_fa710_y2;
  assign f_s_dadda_pg_rca32_fa860_y4 = f_s_dadda_pg_rca32_fa860_y1 | f_s_dadda_pg_rca32_fa860_y3;
  assign f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa860_y4 = f_s_dadda_pg_rca32_fa860_y4;
  assign f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa711_y2 = f_s_dadda_pg_rca32_fa711_y2;
  assign f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa712_y2 = f_s_dadda_pg_rca32_fa712_y2;
  assign f_s_dadda_pg_rca32_fa861_y0 = f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa860_y4 ^ f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa711_y2;
  assign f_s_dadda_pg_rca32_fa861_y1 = f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa860_y4 & f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa711_y2;
  assign f_s_dadda_pg_rca32_fa861_y2 = f_s_dadda_pg_rca32_fa861_y0 ^ f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa712_y2;
  assign f_s_dadda_pg_rca32_fa861_y3 = f_s_dadda_pg_rca32_fa861_y0 & f_s_dadda_pg_rca32_fa861_f_s_dadda_pg_rca32_fa712_y2;
  assign f_s_dadda_pg_rca32_fa861_y4 = f_s_dadda_pg_rca32_fa861_y1 | f_s_dadda_pg_rca32_fa861_y3;
  assign f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa861_y4 = f_s_dadda_pg_rca32_fa861_y4;
  assign f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa713_y2 = f_s_dadda_pg_rca32_fa713_y2;
  assign f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa714_y2 = f_s_dadda_pg_rca32_fa714_y2;
  assign f_s_dadda_pg_rca32_fa862_y0 = f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa861_y4 ^ f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa713_y2;
  assign f_s_dadda_pg_rca32_fa862_y1 = f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa861_y4 & f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa713_y2;
  assign f_s_dadda_pg_rca32_fa862_y2 = f_s_dadda_pg_rca32_fa862_y0 ^ f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa714_y2;
  assign f_s_dadda_pg_rca32_fa862_y3 = f_s_dadda_pg_rca32_fa862_y0 & f_s_dadda_pg_rca32_fa862_f_s_dadda_pg_rca32_fa714_y2;
  assign f_s_dadda_pg_rca32_fa862_y4 = f_s_dadda_pg_rca32_fa862_y1 | f_s_dadda_pg_rca32_fa862_y3;
  assign f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa862_y4 = f_s_dadda_pg_rca32_fa862_y4;
  assign f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa715_y2 = f_s_dadda_pg_rca32_fa715_y2;
  assign f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa716_y2 = f_s_dadda_pg_rca32_fa716_y2;
  assign f_s_dadda_pg_rca32_fa863_y0 = f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa862_y4 ^ f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa715_y2;
  assign f_s_dadda_pg_rca32_fa863_y1 = f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa862_y4 & f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa715_y2;
  assign f_s_dadda_pg_rca32_fa863_y2 = f_s_dadda_pg_rca32_fa863_y0 ^ f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa716_y2;
  assign f_s_dadda_pg_rca32_fa863_y3 = f_s_dadda_pg_rca32_fa863_y0 & f_s_dadda_pg_rca32_fa863_f_s_dadda_pg_rca32_fa716_y2;
  assign f_s_dadda_pg_rca32_fa863_y4 = f_s_dadda_pg_rca32_fa863_y1 | f_s_dadda_pg_rca32_fa863_y3;
  assign f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa863_y4 = f_s_dadda_pg_rca32_fa863_y4;
  assign f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa717_y2 = f_s_dadda_pg_rca32_fa717_y2;
  assign f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa718_y2 = f_s_dadda_pg_rca32_fa718_y2;
  assign f_s_dadda_pg_rca32_fa864_y0 = f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa863_y4 ^ f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa717_y2;
  assign f_s_dadda_pg_rca32_fa864_y1 = f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa863_y4 & f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa717_y2;
  assign f_s_dadda_pg_rca32_fa864_y2 = f_s_dadda_pg_rca32_fa864_y0 ^ f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa718_y2;
  assign f_s_dadda_pg_rca32_fa864_y3 = f_s_dadda_pg_rca32_fa864_y0 & f_s_dadda_pg_rca32_fa864_f_s_dadda_pg_rca32_fa718_y2;
  assign f_s_dadda_pg_rca32_fa864_y4 = f_s_dadda_pg_rca32_fa864_y1 | f_s_dadda_pg_rca32_fa864_y3;
  assign f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa864_y4 = f_s_dadda_pg_rca32_fa864_y4;
  assign f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa719_y2 = f_s_dadda_pg_rca32_fa719_y2;
  assign f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa720_y2 = f_s_dadda_pg_rca32_fa720_y2;
  assign f_s_dadda_pg_rca32_fa865_y0 = f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa864_y4 ^ f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa719_y2;
  assign f_s_dadda_pg_rca32_fa865_y1 = f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa864_y4 & f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa719_y2;
  assign f_s_dadda_pg_rca32_fa865_y2 = f_s_dadda_pg_rca32_fa865_y0 ^ f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa720_y2;
  assign f_s_dadda_pg_rca32_fa865_y3 = f_s_dadda_pg_rca32_fa865_y0 & f_s_dadda_pg_rca32_fa865_f_s_dadda_pg_rca32_fa720_y2;
  assign f_s_dadda_pg_rca32_fa865_y4 = f_s_dadda_pg_rca32_fa865_y1 | f_s_dadda_pg_rca32_fa865_y3;
  assign f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa865_y4 = f_s_dadda_pg_rca32_fa865_y4;
  assign f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa721_y2 = f_s_dadda_pg_rca32_fa721_y2;
  assign f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa722_y2 = f_s_dadda_pg_rca32_fa722_y2;
  assign f_s_dadda_pg_rca32_fa866_y0 = f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa865_y4 ^ f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa721_y2;
  assign f_s_dadda_pg_rca32_fa866_y1 = f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa865_y4 & f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa721_y2;
  assign f_s_dadda_pg_rca32_fa866_y2 = f_s_dadda_pg_rca32_fa866_y0 ^ f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa722_y2;
  assign f_s_dadda_pg_rca32_fa866_y3 = f_s_dadda_pg_rca32_fa866_y0 & f_s_dadda_pg_rca32_fa866_f_s_dadda_pg_rca32_fa722_y2;
  assign f_s_dadda_pg_rca32_fa866_y4 = f_s_dadda_pg_rca32_fa866_y1 | f_s_dadda_pg_rca32_fa866_y3;
  assign f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa866_y4 = f_s_dadda_pg_rca32_fa866_y4;
  assign f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa723_y2 = f_s_dadda_pg_rca32_fa723_y2;
  assign f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa724_y2 = f_s_dadda_pg_rca32_fa724_y2;
  assign f_s_dadda_pg_rca32_fa867_y0 = f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa866_y4 ^ f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa723_y2;
  assign f_s_dadda_pg_rca32_fa867_y1 = f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa866_y4 & f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa723_y2;
  assign f_s_dadda_pg_rca32_fa867_y2 = f_s_dadda_pg_rca32_fa867_y0 ^ f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa724_y2;
  assign f_s_dadda_pg_rca32_fa867_y3 = f_s_dadda_pg_rca32_fa867_y0 & f_s_dadda_pg_rca32_fa867_f_s_dadda_pg_rca32_fa724_y2;
  assign f_s_dadda_pg_rca32_fa867_y4 = f_s_dadda_pg_rca32_fa867_y1 | f_s_dadda_pg_rca32_fa867_y3;
  assign f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa867_y4 = f_s_dadda_pg_rca32_fa867_y4;
  assign f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa725_y2 = f_s_dadda_pg_rca32_fa725_y2;
  assign f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa726_y2 = f_s_dadda_pg_rca32_fa726_y2;
  assign f_s_dadda_pg_rca32_fa868_y0 = f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa867_y4 ^ f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa725_y2;
  assign f_s_dadda_pg_rca32_fa868_y1 = f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa867_y4 & f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa725_y2;
  assign f_s_dadda_pg_rca32_fa868_y2 = f_s_dadda_pg_rca32_fa868_y0 ^ f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa726_y2;
  assign f_s_dadda_pg_rca32_fa868_y3 = f_s_dadda_pg_rca32_fa868_y0 & f_s_dadda_pg_rca32_fa868_f_s_dadda_pg_rca32_fa726_y2;
  assign f_s_dadda_pg_rca32_fa868_y4 = f_s_dadda_pg_rca32_fa868_y1 | f_s_dadda_pg_rca32_fa868_y3;
  assign f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa868_y4 = f_s_dadda_pg_rca32_fa868_y4;
  assign f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa727_y2 = f_s_dadda_pg_rca32_fa727_y2;
  assign f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa728_y2 = f_s_dadda_pg_rca32_fa728_y2;
  assign f_s_dadda_pg_rca32_fa869_y0 = f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa868_y4 ^ f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa727_y2;
  assign f_s_dadda_pg_rca32_fa869_y1 = f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa868_y4 & f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa727_y2;
  assign f_s_dadda_pg_rca32_fa869_y2 = f_s_dadda_pg_rca32_fa869_y0 ^ f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa728_y2;
  assign f_s_dadda_pg_rca32_fa869_y3 = f_s_dadda_pg_rca32_fa869_y0 & f_s_dadda_pg_rca32_fa869_f_s_dadda_pg_rca32_fa728_y2;
  assign f_s_dadda_pg_rca32_fa869_y4 = f_s_dadda_pg_rca32_fa869_y1 | f_s_dadda_pg_rca32_fa869_y3;
  assign f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa869_y4 = f_s_dadda_pg_rca32_fa869_y4;
  assign f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa729_y2 = f_s_dadda_pg_rca32_fa729_y2;
  assign f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa730_y2 = f_s_dadda_pg_rca32_fa730_y2;
  assign f_s_dadda_pg_rca32_fa870_y0 = f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa869_y4 ^ f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa729_y2;
  assign f_s_dadda_pg_rca32_fa870_y1 = f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa869_y4 & f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa729_y2;
  assign f_s_dadda_pg_rca32_fa870_y2 = f_s_dadda_pg_rca32_fa870_y0 ^ f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa730_y2;
  assign f_s_dadda_pg_rca32_fa870_y3 = f_s_dadda_pg_rca32_fa870_y0 & f_s_dadda_pg_rca32_fa870_f_s_dadda_pg_rca32_fa730_y2;
  assign f_s_dadda_pg_rca32_fa870_y4 = f_s_dadda_pg_rca32_fa870_y1 | f_s_dadda_pg_rca32_fa870_y3;
  assign f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa870_y4 = f_s_dadda_pg_rca32_fa870_y4;
  assign f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa731_y2 = f_s_dadda_pg_rca32_fa731_y2;
  assign f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa732_y2 = f_s_dadda_pg_rca32_fa732_y2;
  assign f_s_dadda_pg_rca32_fa871_y0 = f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa870_y4 ^ f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa731_y2;
  assign f_s_dadda_pg_rca32_fa871_y1 = f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa870_y4 & f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa731_y2;
  assign f_s_dadda_pg_rca32_fa871_y2 = f_s_dadda_pg_rca32_fa871_y0 ^ f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa732_y2;
  assign f_s_dadda_pg_rca32_fa871_y3 = f_s_dadda_pg_rca32_fa871_y0 & f_s_dadda_pg_rca32_fa871_f_s_dadda_pg_rca32_fa732_y2;
  assign f_s_dadda_pg_rca32_fa871_y4 = f_s_dadda_pg_rca32_fa871_y1 | f_s_dadda_pg_rca32_fa871_y3;
  assign f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa871_y4 = f_s_dadda_pg_rca32_fa871_y4;
  assign f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa733_y2 = f_s_dadda_pg_rca32_fa733_y2;
  assign f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa734_y2 = f_s_dadda_pg_rca32_fa734_y2;
  assign f_s_dadda_pg_rca32_fa872_y0 = f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa871_y4 ^ f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa733_y2;
  assign f_s_dadda_pg_rca32_fa872_y1 = f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa871_y4 & f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa733_y2;
  assign f_s_dadda_pg_rca32_fa872_y2 = f_s_dadda_pg_rca32_fa872_y0 ^ f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa734_y2;
  assign f_s_dadda_pg_rca32_fa872_y3 = f_s_dadda_pg_rca32_fa872_y0 & f_s_dadda_pg_rca32_fa872_f_s_dadda_pg_rca32_fa734_y2;
  assign f_s_dadda_pg_rca32_fa872_y4 = f_s_dadda_pg_rca32_fa872_y1 | f_s_dadda_pg_rca32_fa872_y3;
  assign f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa872_y4 = f_s_dadda_pg_rca32_fa872_y4;
  assign f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa735_y2 = f_s_dadda_pg_rca32_fa735_y2;
  assign f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa736_y2 = f_s_dadda_pg_rca32_fa736_y2;
  assign f_s_dadda_pg_rca32_fa873_y0 = f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa872_y4 ^ f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa735_y2;
  assign f_s_dadda_pg_rca32_fa873_y1 = f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa872_y4 & f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa735_y2;
  assign f_s_dadda_pg_rca32_fa873_y2 = f_s_dadda_pg_rca32_fa873_y0 ^ f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa736_y2;
  assign f_s_dadda_pg_rca32_fa873_y3 = f_s_dadda_pg_rca32_fa873_y0 & f_s_dadda_pg_rca32_fa873_f_s_dadda_pg_rca32_fa736_y2;
  assign f_s_dadda_pg_rca32_fa873_y4 = f_s_dadda_pg_rca32_fa873_y1 | f_s_dadda_pg_rca32_fa873_y3;
  assign f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa873_y4 = f_s_dadda_pg_rca32_fa873_y4;
  assign f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa737_y2 = f_s_dadda_pg_rca32_fa737_y2;
  assign f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa738_y2 = f_s_dadda_pg_rca32_fa738_y2;
  assign f_s_dadda_pg_rca32_fa874_y0 = f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa873_y4 ^ f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa737_y2;
  assign f_s_dadda_pg_rca32_fa874_y1 = f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa873_y4 & f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa737_y2;
  assign f_s_dadda_pg_rca32_fa874_y2 = f_s_dadda_pg_rca32_fa874_y0 ^ f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa738_y2;
  assign f_s_dadda_pg_rca32_fa874_y3 = f_s_dadda_pg_rca32_fa874_y0 & f_s_dadda_pg_rca32_fa874_f_s_dadda_pg_rca32_fa738_y2;
  assign f_s_dadda_pg_rca32_fa874_y4 = f_s_dadda_pg_rca32_fa874_y1 | f_s_dadda_pg_rca32_fa874_y3;
  assign f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa874_y4 = f_s_dadda_pg_rca32_fa874_y4;
  assign f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa739_y2 = f_s_dadda_pg_rca32_fa739_y2;
  assign f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa740_y2 = f_s_dadda_pg_rca32_fa740_y2;
  assign f_s_dadda_pg_rca32_fa875_y0 = f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa874_y4 ^ f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa739_y2;
  assign f_s_dadda_pg_rca32_fa875_y1 = f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa874_y4 & f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa739_y2;
  assign f_s_dadda_pg_rca32_fa875_y2 = f_s_dadda_pg_rca32_fa875_y0 ^ f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa740_y2;
  assign f_s_dadda_pg_rca32_fa875_y3 = f_s_dadda_pg_rca32_fa875_y0 & f_s_dadda_pg_rca32_fa875_f_s_dadda_pg_rca32_fa740_y2;
  assign f_s_dadda_pg_rca32_fa875_y4 = f_s_dadda_pg_rca32_fa875_y1 | f_s_dadda_pg_rca32_fa875_y3;
  assign f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa875_y4 = f_s_dadda_pg_rca32_fa875_y4;
  assign f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa741_y2 = f_s_dadda_pg_rca32_fa741_y2;
  assign f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa742_y2 = f_s_dadda_pg_rca32_fa742_y2;
  assign f_s_dadda_pg_rca32_fa876_y0 = f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa875_y4 ^ f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa741_y2;
  assign f_s_dadda_pg_rca32_fa876_y1 = f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa875_y4 & f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa741_y2;
  assign f_s_dadda_pg_rca32_fa876_y2 = f_s_dadda_pg_rca32_fa876_y0 ^ f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa742_y2;
  assign f_s_dadda_pg_rca32_fa876_y3 = f_s_dadda_pg_rca32_fa876_y0 & f_s_dadda_pg_rca32_fa876_f_s_dadda_pg_rca32_fa742_y2;
  assign f_s_dadda_pg_rca32_fa876_y4 = f_s_dadda_pg_rca32_fa876_y1 | f_s_dadda_pg_rca32_fa876_y3;
  assign f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa876_y4 = f_s_dadda_pg_rca32_fa876_y4;
  assign f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa743_y2 = f_s_dadda_pg_rca32_fa743_y2;
  assign f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa744_y2 = f_s_dadda_pg_rca32_fa744_y2;
  assign f_s_dadda_pg_rca32_fa877_y0 = f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa876_y4 ^ f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa743_y2;
  assign f_s_dadda_pg_rca32_fa877_y1 = f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa876_y4 & f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa743_y2;
  assign f_s_dadda_pg_rca32_fa877_y2 = f_s_dadda_pg_rca32_fa877_y0 ^ f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa744_y2;
  assign f_s_dadda_pg_rca32_fa877_y3 = f_s_dadda_pg_rca32_fa877_y0 & f_s_dadda_pg_rca32_fa877_f_s_dadda_pg_rca32_fa744_y2;
  assign f_s_dadda_pg_rca32_fa877_y4 = f_s_dadda_pg_rca32_fa877_y1 | f_s_dadda_pg_rca32_fa877_y3;
  assign f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa877_y4 = f_s_dadda_pg_rca32_fa877_y4;
  assign f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa745_y2 = f_s_dadda_pg_rca32_fa745_y2;
  assign f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa746_y2 = f_s_dadda_pg_rca32_fa746_y2;
  assign f_s_dadda_pg_rca32_fa878_y0 = f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa877_y4 ^ f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa745_y2;
  assign f_s_dadda_pg_rca32_fa878_y1 = f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa877_y4 & f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa745_y2;
  assign f_s_dadda_pg_rca32_fa878_y2 = f_s_dadda_pg_rca32_fa878_y0 ^ f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa746_y2;
  assign f_s_dadda_pg_rca32_fa878_y3 = f_s_dadda_pg_rca32_fa878_y0 & f_s_dadda_pg_rca32_fa878_f_s_dadda_pg_rca32_fa746_y2;
  assign f_s_dadda_pg_rca32_fa878_y4 = f_s_dadda_pg_rca32_fa878_y1 | f_s_dadda_pg_rca32_fa878_y3;
  assign f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa878_y4 = f_s_dadda_pg_rca32_fa878_y4;
  assign f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa747_y2 = f_s_dadda_pg_rca32_fa747_y2;
  assign f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa748_y2 = f_s_dadda_pg_rca32_fa748_y2;
  assign f_s_dadda_pg_rca32_fa879_y0 = f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa878_y4 ^ f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa747_y2;
  assign f_s_dadda_pg_rca32_fa879_y1 = f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa878_y4 & f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa747_y2;
  assign f_s_dadda_pg_rca32_fa879_y2 = f_s_dadda_pg_rca32_fa879_y0 ^ f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa748_y2;
  assign f_s_dadda_pg_rca32_fa879_y3 = f_s_dadda_pg_rca32_fa879_y0 & f_s_dadda_pg_rca32_fa879_f_s_dadda_pg_rca32_fa748_y2;
  assign f_s_dadda_pg_rca32_fa879_y4 = f_s_dadda_pg_rca32_fa879_y1 | f_s_dadda_pg_rca32_fa879_y3;
  assign f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa879_y4 = f_s_dadda_pg_rca32_fa879_y4;
  assign f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa749_y2 = f_s_dadda_pg_rca32_fa749_y2;
  assign f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa750_y2 = f_s_dadda_pg_rca32_fa750_y2;
  assign f_s_dadda_pg_rca32_fa880_y0 = f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa879_y4 ^ f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa749_y2;
  assign f_s_dadda_pg_rca32_fa880_y1 = f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa879_y4 & f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa749_y2;
  assign f_s_dadda_pg_rca32_fa880_y2 = f_s_dadda_pg_rca32_fa880_y0 ^ f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa750_y2;
  assign f_s_dadda_pg_rca32_fa880_y3 = f_s_dadda_pg_rca32_fa880_y0 & f_s_dadda_pg_rca32_fa880_f_s_dadda_pg_rca32_fa750_y2;
  assign f_s_dadda_pg_rca32_fa880_y4 = f_s_dadda_pg_rca32_fa880_y1 | f_s_dadda_pg_rca32_fa880_y3;
  assign f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa880_y4 = f_s_dadda_pg_rca32_fa880_y4;
  assign f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa751_y2 = f_s_dadda_pg_rca32_fa751_y2;
  assign f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa752_y2 = f_s_dadda_pg_rca32_fa752_y2;
  assign f_s_dadda_pg_rca32_fa881_y0 = f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa880_y4 ^ f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa751_y2;
  assign f_s_dadda_pg_rca32_fa881_y1 = f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa880_y4 & f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa751_y2;
  assign f_s_dadda_pg_rca32_fa881_y2 = f_s_dadda_pg_rca32_fa881_y0 ^ f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa752_y2;
  assign f_s_dadda_pg_rca32_fa881_y3 = f_s_dadda_pg_rca32_fa881_y0 & f_s_dadda_pg_rca32_fa881_f_s_dadda_pg_rca32_fa752_y2;
  assign f_s_dadda_pg_rca32_fa881_y4 = f_s_dadda_pg_rca32_fa881_y1 | f_s_dadda_pg_rca32_fa881_y3;
  assign f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa881_y4 = f_s_dadda_pg_rca32_fa881_y4;
  assign f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa753_y2 = f_s_dadda_pg_rca32_fa753_y2;
  assign f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa754_y2 = f_s_dadda_pg_rca32_fa754_y2;
  assign f_s_dadda_pg_rca32_fa882_y0 = f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa881_y4 ^ f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa753_y2;
  assign f_s_dadda_pg_rca32_fa882_y1 = f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa881_y4 & f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa753_y2;
  assign f_s_dadda_pg_rca32_fa882_y2 = f_s_dadda_pg_rca32_fa882_y0 ^ f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa754_y2;
  assign f_s_dadda_pg_rca32_fa882_y3 = f_s_dadda_pg_rca32_fa882_y0 & f_s_dadda_pg_rca32_fa882_f_s_dadda_pg_rca32_fa754_y2;
  assign f_s_dadda_pg_rca32_fa882_y4 = f_s_dadda_pg_rca32_fa882_y1 | f_s_dadda_pg_rca32_fa882_y3;
  assign f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa882_y4 = f_s_dadda_pg_rca32_fa882_y4;
  assign f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa755_y2 = f_s_dadda_pg_rca32_fa755_y2;
  assign f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa756_y2 = f_s_dadda_pg_rca32_fa756_y2;
  assign f_s_dadda_pg_rca32_fa883_y0 = f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa882_y4 ^ f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa755_y2;
  assign f_s_dadda_pg_rca32_fa883_y1 = f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa882_y4 & f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa755_y2;
  assign f_s_dadda_pg_rca32_fa883_y2 = f_s_dadda_pg_rca32_fa883_y0 ^ f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa756_y2;
  assign f_s_dadda_pg_rca32_fa883_y3 = f_s_dadda_pg_rca32_fa883_y0 & f_s_dadda_pg_rca32_fa883_f_s_dadda_pg_rca32_fa756_y2;
  assign f_s_dadda_pg_rca32_fa883_y4 = f_s_dadda_pg_rca32_fa883_y1 | f_s_dadda_pg_rca32_fa883_y3;
  assign f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa883_y4 = f_s_dadda_pg_rca32_fa883_y4;
  assign f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa757_y2 = f_s_dadda_pg_rca32_fa757_y2;
  assign f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa758_y2 = f_s_dadda_pg_rca32_fa758_y2;
  assign f_s_dadda_pg_rca32_fa884_y0 = f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa883_y4 ^ f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa757_y2;
  assign f_s_dadda_pg_rca32_fa884_y1 = f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa883_y4 & f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa757_y2;
  assign f_s_dadda_pg_rca32_fa884_y2 = f_s_dadda_pg_rca32_fa884_y0 ^ f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa758_y2;
  assign f_s_dadda_pg_rca32_fa884_y3 = f_s_dadda_pg_rca32_fa884_y0 & f_s_dadda_pg_rca32_fa884_f_s_dadda_pg_rca32_fa758_y2;
  assign f_s_dadda_pg_rca32_fa884_y4 = f_s_dadda_pg_rca32_fa884_y1 | f_s_dadda_pg_rca32_fa884_y3;
  assign f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa884_y4 = f_s_dadda_pg_rca32_fa884_y4;
  assign f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa759_y2 = f_s_dadda_pg_rca32_fa759_y2;
  assign f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa760_y2 = f_s_dadda_pg_rca32_fa760_y2;
  assign f_s_dadda_pg_rca32_fa885_y0 = f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa884_y4 ^ f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa759_y2;
  assign f_s_dadda_pg_rca32_fa885_y1 = f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa884_y4 & f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa759_y2;
  assign f_s_dadda_pg_rca32_fa885_y2 = f_s_dadda_pg_rca32_fa885_y0 ^ f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa760_y2;
  assign f_s_dadda_pg_rca32_fa885_y3 = f_s_dadda_pg_rca32_fa885_y0 & f_s_dadda_pg_rca32_fa885_f_s_dadda_pg_rca32_fa760_y2;
  assign f_s_dadda_pg_rca32_fa885_y4 = f_s_dadda_pg_rca32_fa885_y1 | f_s_dadda_pg_rca32_fa885_y3;
  assign f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa885_y4 = f_s_dadda_pg_rca32_fa885_y4;
  assign f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa761_y2 = f_s_dadda_pg_rca32_fa761_y2;
  assign f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa762_y2 = f_s_dadda_pg_rca32_fa762_y2;
  assign f_s_dadda_pg_rca32_fa886_y0 = f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa885_y4 ^ f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa761_y2;
  assign f_s_dadda_pg_rca32_fa886_y1 = f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa885_y4 & f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa761_y2;
  assign f_s_dadda_pg_rca32_fa886_y2 = f_s_dadda_pg_rca32_fa886_y0 ^ f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa762_y2;
  assign f_s_dadda_pg_rca32_fa886_y3 = f_s_dadda_pg_rca32_fa886_y0 & f_s_dadda_pg_rca32_fa886_f_s_dadda_pg_rca32_fa762_y2;
  assign f_s_dadda_pg_rca32_fa886_y4 = f_s_dadda_pg_rca32_fa886_y1 | f_s_dadda_pg_rca32_fa886_y3;
  assign f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa886_y4 = f_s_dadda_pg_rca32_fa886_y4;
  assign f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa763_y2 = f_s_dadda_pg_rca32_fa763_y2;
  assign f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa764_y2 = f_s_dadda_pg_rca32_fa764_y2;
  assign f_s_dadda_pg_rca32_fa887_y0 = f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa886_y4 ^ f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa763_y2;
  assign f_s_dadda_pg_rca32_fa887_y1 = f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa886_y4 & f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa763_y2;
  assign f_s_dadda_pg_rca32_fa887_y2 = f_s_dadda_pg_rca32_fa887_y0 ^ f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa764_y2;
  assign f_s_dadda_pg_rca32_fa887_y3 = f_s_dadda_pg_rca32_fa887_y0 & f_s_dadda_pg_rca32_fa887_f_s_dadda_pg_rca32_fa764_y2;
  assign f_s_dadda_pg_rca32_fa887_y4 = f_s_dadda_pg_rca32_fa887_y1 | f_s_dadda_pg_rca32_fa887_y3;
  assign f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa887_y4 = f_s_dadda_pg_rca32_fa887_y4;
  assign f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa765_y2 = f_s_dadda_pg_rca32_fa765_y2;
  assign f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa766_y2 = f_s_dadda_pg_rca32_fa766_y2;
  assign f_s_dadda_pg_rca32_fa888_y0 = f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa887_y4 ^ f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa765_y2;
  assign f_s_dadda_pg_rca32_fa888_y1 = f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa887_y4 & f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa765_y2;
  assign f_s_dadda_pg_rca32_fa888_y2 = f_s_dadda_pg_rca32_fa888_y0 ^ f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa766_y2;
  assign f_s_dadda_pg_rca32_fa888_y3 = f_s_dadda_pg_rca32_fa888_y0 & f_s_dadda_pg_rca32_fa888_f_s_dadda_pg_rca32_fa766_y2;
  assign f_s_dadda_pg_rca32_fa888_y4 = f_s_dadda_pg_rca32_fa888_y1 | f_s_dadda_pg_rca32_fa888_y3;
  assign f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa888_y4 = f_s_dadda_pg_rca32_fa888_y4;
  assign f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa767_y2 = f_s_dadda_pg_rca32_fa767_y2;
  assign f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa768_y2 = f_s_dadda_pg_rca32_fa768_y2;
  assign f_s_dadda_pg_rca32_fa889_y0 = f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa888_y4 ^ f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa767_y2;
  assign f_s_dadda_pg_rca32_fa889_y1 = f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa888_y4 & f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa767_y2;
  assign f_s_dadda_pg_rca32_fa889_y2 = f_s_dadda_pg_rca32_fa889_y0 ^ f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa768_y2;
  assign f_s_dadda_pg_rca32_fa889_y3 = f_s_dadda_pg_rca32_fa889_y0 & f_s_dadda_pg_rca32_fa889_f_s_dadda_pg_rca32_fa768_y2;
  assign f_s_dadda_pg_rca32_fa889_y4 = f_s_dadda_pg_rca32_fa889_y1 | f_s_dadda_pg_rca32_fa889_y3;
  assign f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa889_y4 = f_s_dadda_pg_rca32_fa889_y4;
  assign f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa769_y2 = f_s_dadda_pg_rca32_fa769_y2;
  assign f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa770_y2 = f_s_dadda_pg_rca32_fa770_y2;
  assign f_s_dadda_pg_rca32_fa890_y0 = f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa889_y4 ^ f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa769_y2;
  assign f_s_dadda_pg_rca32_fa890_y1 = f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa889_y4 & f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa769_y2;
  assign f_s_dadda_pg_rca32_fa890_y2 = f_s_dadda_pg_rca32_fa890_y0 ^ f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa770_y2;
  assign f_s_dadda_pg_rca32_fa890_y3 = f_s_dadda_pg_rca32_fa890_y0 & f_s_dadda_pg_rca32_fa890_f_s_dadda_pg_rca32_fa770_y2;
  assign f_s_dadda_pg_rca32_fa890_y4 = f_s_dadda_pg_rca32_fa890_y1 | f_s_dadda_pg_rca32_fa890_y3;
  assign f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa890_y4 = f_s_dadda_pg_rca32_fa890_y4;
  assign f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa771_y2 = f_s_dadda_pg_rca32_fa771_y2;
  assign f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa772_y2 = f_s_dadda_pg_rca32_fa772_y2;
  assign f_s_dadda_pg_rca32_fa891_y0 = f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa890_y4 ^ f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa771_y2;
  assign f_s_dadda_pg_rca32_fa891_y1 = f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa890_y4 & f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa771_y2;
  assign f_s_dadda_pg_rca32_fa891_y2 = f_s_dadda_pg_rca32_fa891_y0 ^ f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa772_y2;
  assign f_s_dadda_pg_rca32_fa891_y3 = f_s_dadda_pg_rca32_fa891_y0 & f_s_dadda_pg_rca32_fa891_f_s_dadda_pg_rca32_fa772_y2;
  assign f_s_dadda_pg_rca32_fa891_y4 = f_s_dadda_pg_rca32_fa891_y1 | f_s_dadda_pg_rca32_fa891_y3;
  assign f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa891_y4 = f_s_dadda_pg_rca32_fa891_y4;
  assign f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa773_y2 = f_s_dadda_pg_rca32_fa773_y2;
  assign f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa774_y2 = f_s_dadda_pg_rca32_fa774_y2;
  assign f_s_dadda_pg_rca32_fa892_y0 = f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa891_y4 ^ f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa773_y2;
  assign f_s_dadda_pg_rca32_fa892_y1 = f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa891_y4 & f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa773_y2;
  assign f_s_dadda_pg_rca32_fa892_y2 = f_s_dadda_pg_rca32_fa892_y0 ^ f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa774_y2;
  assign f_s_dadda_pg_rca32_fa892_y3 = f_s_dadda_pg_rca32_fa892_y0 & f_s_dadda_pg_rca32_fa892_f_s_dadda_pg_rca32_fa774_y2;
  assign f_s_dadda_pg_rca32_fa892_y4 = f_s_dadda_pg_rca32_fa892_y1 | f_s_dadda_pg_rca32_fa892_y3;
  assign f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa892_y4 = f_s_dadda_pg_rca32_fa892_y4;
  assign f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa775_y2 = f_s_dadda_pg_rca32_fa775_y2;
  assign f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa776_y2 = f_s_dadda_pg_rca32_fa776_y2;
  assign f_s_dadda_pg_rca32_fa893_y0 = f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa892_y4 ^ f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa775_y2;
  assign f_s_dadda_pg_rca32_fa893_y1 = f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa892_y4 & f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa775_y2;
  assign f_s_dadda_pg_rca32_fa893_y2 = f_s_dadda_pg_rca32_fa893_y0 ^ f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa776_y2;
  assign f_s_dadda_pg_rca32_fa893_y3 = f_s_dadda_pg_rca32_fa893_y0 & f_s_dadda_pg_rca32_fa893_f_s_dadda_pg_rca32_fa776_y2;
  assign f_s_dadda_pg_rca32_fa893_y4 = f_s_dadda_pg_rca32_fa893_y1 | f_s_dadda_pg_rca32_fa893_y3;
  assign f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa893_y4 = f_s_dadda_pg_rca32_fa893_y4;
  assign f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa777_y2 = f_s_dadda_pg_rca32_fa777_y2;
  assign f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa778_y2 = f_s_dadda_pg_rca32_fa778_y2;
  assign f_s_dadda_pg_rca32_fa894_y0 = f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa893_y4 ^ f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa777_y2;
  assign f_s_dadda_pg_rca32_fa894_y1 = f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa893_y4 & f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa777_y2;
  assign f_s_dadda_pg_rca32_fa894_y2 = f_s_dadda_pg_rca32_fa894_y0 ^ f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa778_y2;
  assign f_s_dadda_pg_rca32_fa894_y3 = f_s_dadda_pg_rca32_fa894_y0 & f_s_dadda_pg_rca32_fa894_f_s_dadda_pg_rca32_fa778_y2;
  assign f_s_dadda_pg_rca32_fa894_y4 = f_s_dadda_pg_rca32_fa894_y1 | f_s_dadda_pg_rca32_fa894_y3;
  assign f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa894_y4 = f_s_dadda_pg_rca32_fa894_y4;
  assign f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa779_y2 = f_s_dadda_pg_rca32_fa779_y2;
  assign f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa780_y2 = f_s_dadda_pg_rca32_fa780_y2;
  assign f_s_dadda_pg_rca32_fa895_y0 = f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa894_y4 ^ f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa779_y2;
  assign f_s_dadda_pg_rca32_fa895_y1 = f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa894_y4 & f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa779_y2;
  assign f_s_dadda_pg_rca32_fa895_y2 = f_s_dadda_pg_rca32_fa895_y0 ^ f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa780_y2;
  assign f_s_dadda_pg_rca32_fa895_y3 = f_s_dadda_pg_rca32_fa895_y0 & f_s_dadda_pg_rca32_fa895_f_s_dadda_pg_rca32_fa780_y2;
  assign f_s_dadda_pg_rca32_fa895_y4 = f_s_dadda_pg_rca32_fa895_y1 | f_s_dadda_pg_rca32_fa895_y3;
  assign f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa895_y4 = f_s_dadda_pg_rca32_fa895_y4;
  assign f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa781_y2 = f_s_dadda_pg_rca32_fa781_y2;
  assign f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa782_y2 = f_s_dadda_pg_rca32_fa782_y2;
  assign f_s_dadda_pg_rca32_fa896_y0 = f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa895_y4 ^ f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa781_y2;
  assign f_s_dadda_pg_rca32_fa896_y1 = f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa895_y4 & f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa781_y2;
  assign f_s_dadda_pg_rca32_fa896_y2 = f_s_dadda_pg_rca32_fa896_y0 ^ f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa782_y2;
  assign f_s_dadda_pg_rca32_fa896_y3 = f_s_dadda_pg_rca32_fa896_y0 & f_s_dadda_pg_rca32_fa896_f_s_dadda_pg_rca32_fa782_y2;
  assign f_s_dadda_pg_rca32_fa896_y4 = f_s_dadda_pg_rca32_fa896_y1 | f_s_dadda_pg_rca32_fa896_y3;
  assign f_s_dadda_pg_rca32_nand_28_31_a_28 = a_28;
  assign f_s_dadda_pg_rca32_nand_28_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_28_31_y0 = ~(f_s_dadda_pg_rca32_nand_28_31_a_28 & f_s_dadda_pg_rca32_nand_28_31_b_31);
  assign f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_fa896_y4 = f_s_dadda_pg_rca32_fa896_y4;
  assign f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_nand_28_31_y0 = f_s_dadda_pg_rca32_nand_28_31_y0;
  assign f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_fa783_y2 = f_s_dadda_pg_rca32_fa783_y2;
  assign f_s_dadda_pg_rca32_fa897_y0 = f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_fa896_y4 ^ f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_nand_28_31_y0;
  assign f_s_dadda_pg_rca32_fa897_y1 = f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_fa896_y4 & f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_nand_28_31_y0;
  assign f_s_dadda_pg_rca32_fa897_y2 = f_s_dadda_pg_rca32_fa897_y0 ^ f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_fa783_y2;
  assign f_s_dadda_pg_rca32_fa897_y3 = f_s_dadda_pg_rca32_fa897_y0 & f_s_dadda_pg_rca32_fa897_f_s_dadda_pg_rca32_fa783_y2;
  assign f_s_dadda_pg_rca32_fa897_y4 = f_s_dadda_pg_rca32_fa897_y1 | f_s_dadda_pg_rca32_fa897_y3;
  assign f_s_dadda_pg_rca32_and_30_30_a_30 = a_30;
  assign f_s_dadda_pg_rca32_and_30_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_and_30_30_y0 = f_s_dadda_pg_rca32_and_30_30_a_30 & f_s_dadda_pg_rca32_and_30_30_b_30;
  assign f_s_dadda_pg_rca32_nand_29_31_a_29 = a_29;
  assign f_s_dadda_pg_rca32_nand_29_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_29_31_y0 = ~(f_s_dadda_pg_rca32_nand_29_31_a_29 & f_s_dadda_pg_rca32_nand_29_31_b_31);
  assign f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_fa897_y4 = f_s_dadda_pg_rca32_fa897_y4;
  assign f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_and_30_30_y0 = f_s_dadda_pg_rca32_and_30_30_y0;
  assign f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_nand_29_31_y0 = f_s_dadda_pg_rca32_nand_29_31_y0;
  assign f_s_dadda_pg_rca32_fa898_y0 = f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_fa897_y4 ^ f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_and_30_30_y0;
  assign f_s_dadda_pg_rca32_fa898_y1 = f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_fa897_y4 & f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_and_30_30_y0;
  assign f_s_dadda_pg_rca32_fa898_y2 = f_s_dadda_pg_rca32_fa898_y0 ^ f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_nand_29_31_y0;
  assign f_s_dadda_pg_rca32_fa898_y3 = f_s_dadda_pg_rca32_fa898_y0 & f_s_dadda_pg_rca32_fa898_f_s_dadda_pg_rca32_nand_29_31_y0;
  assign f_s_dadda_pg_rca32_fa898_y4 = f_s_dadda_pg_rca32_fa898_y1 | f_s_dadda_pg_rca32_fa898_y3;
  assign f_s_dadda_pg_rca32_nand_31_30_a_31 = a_31;
  assign f_s_dadda_pg_rca32_nand_31_30_b_30 = b_30;
  assign f_s_dadda_pg_rca32_nand_31_30_y0 = ~(f_s_dadda_pg_rca32_nand_31_30_a_31 & f_s_dadda_pg_rca32_nand_31_30_b_30);
  assign f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_fa898_y4 = f_s_dadda_pg_rca32_fa898_y4;
  assign f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_fa840_y4 = f_s_dadda_pg_rca32_fa840_y4;
  assign f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_nand_31_30_y0 = f_s_dadda_pg_rca32_nand_31_30_y0;
  assign f_s_dadda_pg_rca32_fa899_y0 = f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_fa898_y4 ^ f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_fa840_y4;
  assign f_s_dadda_pg_rca32_fa899_y1 = f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_fa898_y4 & f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_fa840_y4;
  assign f_s_dadda_pg_rca32_fa899_y2 = f_s_dadda_pg_rca32_fa899_y0 ^ f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_nand_31_30_y0;
  assign f_s_dadda_pg_rca32_fa899_y3 = f_s_dadda_pg_rca32_fa899_y0 & f_s_dadda_pg_rca32_fa899_f_s_dadda_pg_rca32_nand_31_30_y0;
  assign f_s_dadda_pg_rca32_fa899_y4 = f_s_dadda_pg_rca32_fa899_y1 | f_s_dadda_pg_rca32_fa899_y3;
  assign f_s_dadda_pg_rca32_and_0_0_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_0_0_y0 = f_s_dadda_pg_rca32_and_0_0_a_0 & f_s_dadda_pg_rca32_and_0_0_b_0;
  assign f_s_dadda_pg_rca32_and_1_0_a_1 = a_1;
  assign f_s_dadda_pg_rca32_and_1_0_b_0 = b_0;
  assign f_s_dadda_pg_rca32_and_1_0_y0 = f_s_dadda_pg_rca32_and_1_0_a_1 & f_s_dadda_pg_rca32_and_1_0_b_0;
  assign f_s_dadda_pg_rca32_and_0_2_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_2_b_2 = b_2;
  assign f_s_dadda_pg_rca32_and_0_2_y0 = f_s_dadda_pg_rca32_and_0_2_a_0 & f_s_dadda_pg_rca32_and_0_2_b_2;
  assign f_s_dadda_pg_rca32_nand_30_31_a_30 = a_30;
  assign f_s_dadda_pg_rca32_nand_30_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_nand_30_31_y0 = ~(f_s_dadda_pg_rca32_nand_30_31_a_30 & f_s_dadda_pg_rca32_nand_30_31_b_31);
  assign f_s_dadda_pg_rca32_and_0_1_a_0 = a_0;
  assign f_s_dadda_pg_rca32_and_0_1_b_1 = b_1;
  assign f_s_dadda_pg_rca32_and_0_1_y0 = f_s_dadda_pg_rca32_and_0_1_a_0 & f_s_dadda_pg_rca32_and_0_1_b_1;
  assign f_s_dadda_pg_rca32_and_31_31_a_31 = a_31;
  assign f_s_dadda_pg_rca32_and_31_31_b_31 = b_31;
  assign f_s_dadda_pg_rca32_and_31_31_y0 = f_s_dadda_pg_rca32_and_31_31_a_31 & f_s_dadda_pg_rca32_and_31_31_b_31;
  assign constant_wire_value_0_f_s_dadda_pg_rca32_and_1_0_y0 = f_s_dadda_pg_rca32_and_1_0_y0;
  assign constant_wire_value_0_f_s_dadda_pg_rca32_and_0_1_y0 = f_s_dadda_pg_rca32_and_0_1_y0;
  assign constant_wire_value_0_y0 = constant_wire_value_0_f_s_dadda_pg_rca32_and_1_0_y0 ^ constant_wire_value_0_f_s_dadda_pg_rca32_and_0_1_y0;
  assign constant_wire_value_0_y1 = ~(constant_wire_value_0_f_s_dadda_pg_rca32_and_1_0_y0 ^ constant_wire_value_0_f_s_dadda_pg_rca32_and_0_1_y0);
  assign constant_wire_0 = ~(constant_wire_value_0_y0 | constant_wire_value_0_y1);
  assign f_s_dadda_pg_rca32_u_pg_rca_fa0_f_s_dadda_pg_rca32_and_1_0_y0 = f_s_dadda_pg_rca32_and_1_0_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa0_f_s_dadda_pg_rca32_and_0_1_y0 = f_s_dadda_pg_rca32_and_0_1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa0_constant_wire_0 = constant_wire_0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa0_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa0_f_s_dadda_pg_rca32_and_1_0_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa0_f_s_dadda_pg_rca32_and_0_1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa0_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa0_f_s_dadda_pg_rca32_and_1_0_y0 & f_s_dadda_pg_rca32_u_pg_rca_fa0_f_s_dadda_pg_rca32_and_0_1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa0_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa0_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa0_constant_wire_0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and0_constant_wire_0 = constant_wire_0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and0_f_s_dadda_pg_rca32_u_pg_rca_fa0_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa0_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and0_y0 = f_s_dadda_pg_rca32_u_pg_rca_and0_constant_wire_0 & f_s_dadda_pg_rca32_u_pg_rca_and0_f_s_dadda_pg_rca32_u_pg_rca_fa0_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or0_f_s_dadda_pg_rca32_u_pg_rca_and0_y0 = f_s_dadda_pg_rca32_u_pg_rca_and0_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or0_f_s_dadda_pg_rca32_u_pg_rca_fa0_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa0_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or0_y0 = f_s_dadda_pg_rca32_u_pg_rca_or0_f_s_dadda_pg_rca32_u_pg_rca_and0_y0 | f_s_dadda_pg_rca32_u_pg_rca_or0_f_s_dadda_pg_rca32_u_pg_rca_fa0_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_and_0_2_y0 = f_s_dadda_pg_rca32_and_0_2_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_ha29_y0 = f_s_dadda_pg_rca32_ha29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_u_pg_rca_or0_y0 = f_s_dadda_pg_rca32_u_pg_rca_or0_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa1_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_and_0_2_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_ha29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa1_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_and_0_2_y0 & f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_ha29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa1_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa1_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa1_f_s_dadda_pg_rca32_u_pg_rca_or0_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and1_f_s_dadda_pg_rca32_u_pg_rca_or0_y0 = f_s_dadda_pg_rca32_u_pg_rca_or0_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and1_f_s_dadda_pg_rca32_u_pg_rca_fa1_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and1_y0 = f_s_dadda_pg_rca32_u_pg_rca_and1_f_s_dadda_pg_rca32_u_pg_rca_or0_y0 & f_s_dadda_pg_rca32_u_pg_rca_and1_f_s_dadda_pg_rca32_u_pg_rca_fa1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or1_f_s_dadda_pg_rca32_u_pg_rca_and1_y0 = f_s_dadda_pg_rca32_u_pg_rca_and1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or1_f_s_dadda_pg_rca32_u_pg_rca_fa1_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa1_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or1_y0 = f_s_dadda_pg_rca32_u_pg_rca_or1_f_s_dadda_pg_rca32_u_pg_rca_and1_y0 | f_s_dadda_pg_rca32_u_pg_rca_or1_f_s_dadda_pg_rca32_u_pg_rca_fa1_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_ha28_y0 = f_s_dadda_pg_rca32_ha28_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_fa841_y2 = f_s_dadda_pg_rca32_fa841_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_u_pg_rca_or1_y0 = f_s_dadda_pg_rca32_u_pg_rca_or1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa2_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_ha28_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_fa841_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa2_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_ha28_y0 & f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_fa841_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa2_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa2_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa2_f_s_dadda_pg_rca32_u_pg_rca_or1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and2_f_s_dadda_pg_rca32_u_pg_rca_or1_y0 = f_s_dadda_pg_rca32_u_pg_rca_or1_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and2_f_s_dadda_pg_rca32_u_pg_rca_fa2_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa2_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and2_y0 = f_s_dadda_pg_rca32_u_pg_rca_and2_f_s_dadda_pg_rca32_u_pg_rca_or1_y0 & f_s_dadda_pg_rca32_u_pg_rca_and2_f_s_dadda_pg_rca32_u_pg_rca_fa2_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or2_f_s_dadda_pg_rca32_u_pg_rca_and2_y0 = f_s_dadda_pg_rca32_u_pg_rca_and2_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or2_f_s_dadda_pg_rca32_u_pg_rca_fa2_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa2_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or2_y0 = f_s_dadda_pg_rca32_u_pg_rca_or2_f_s_dadda_pg_rca32_u_pg_rca_and2_y0 | f_s_dadda_pg_rca32_u_pg_rca_or2_f_s_dadda_pg_rca32_u_pg_rca_fa2_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_fa784_y2 = f_s_dadda_pg_rca32_fa784_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_fa842_y2 = f_s_dadda_pg_rca32_fa842_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_u_pg_rca_or2_y0 = f_s_dadda_pg_rca32_u_pg_rca_or2_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa3_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_fa784_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_fa842_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa3_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_fa784_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_fa842_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa3_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa3_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa3_f_s_dadda_pg_rca32_u_pg_rca_or2_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and3_f_s_dadda_pg_rca32_u_pg_rca_or2_y0 = f_s_dadda_pg_rca32_u_pg_rca_or2_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and3_f_s_dadda_pg_rca32_u_pg_rca_fa3_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa3_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and3_y0 = f_s_dadda_pg_rca32_u_pg_rca_and3_f_s_dadda_pg_rca32_u_pg_rca_or2_y0 & f_s_dadda_pg_rca32_u_pg_rca_and3_f_s_dadda_pg_rca32_u_pg_rca_fa3_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or3_f_s_dadda_pg_rca32_u_pg_rca_and3_y0 = f_s_dadda_pg_rca32_u_pg_rca_and3_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or3_f_s_dadda_pg_rca32_u_pg_rca_fa3_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa3_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or3_y0 = f_s_dadda_pg_rca32_u_pg_rca_or3_f_s_dadda_pg_rca32_u_pg_rca_and3_y0 | f_s_dadda_pg_rca32_u_pg_rca_or3_f_s_dadda_pg_rca32_u_pg_rca_fa3_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_fa785_y2 = f_s_dadda_pg_rca32_fa785_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_fa843_y2 = f_s_dadda_pg_rca32_fa843_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_u_pg_rca_or3_y0 = f_s_dadda_pg_rca32_u_pg_rca_or3_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa4_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_fa785_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_fa843_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa4_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_fa785_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_fa843_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa4_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa4_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa4_f_s_dadda_pg_rca32_u_pg_rca_or3_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and4_f_s_dadda_pg_rca32_u_pg_rca_or3_y0 = f_s_dadda_pg_rca32_u_pg_rca_or3_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and4_f_s_dadda_pg_rca32_u_pg_rca_fa4_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa4_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and4_y0 = f_s_dadda_pg_rca32_u_pg_rca_and4_f_s_dadda_pg_rca32_u_pg_rca_or3_y0 & f_s_dadda_pg_rca32_u_pg_rca_and4_f_s_dadda_pg_rca32_u_pg_rca_fa4_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or4_f_s_dadda_pg_rca32_u_pg_rca_and4_y0 = f_s_dadda_pg_rca32_u_pg_rca_and4_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or4_f_s_dadda_pg_rca32_u_pg_rca_fa4_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa4_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or4_y0 = f_s_dadda_pg_rca32_u_pg_rca_or4_f_s_dadda_pg_rca32_u_pg_rca_and4_y0 | f_s_dadda_pg_rca32_u_pg_rca_or4_f_s_dadda_pg_rca32_u_pg_rca_fa4_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_fa786_y2 = f_s_dadda_pg_rca32_fa786_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_fa844_y2 = f_s_dadda_pg_rca32_fa844_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_u_pg_rca_or4_y0 = f_s_dadda_pg_rca32_u_pg_rca_or4_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa5_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_fa786_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_fa844_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa5_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_fa786_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_fa844_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa5_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa5_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa5_f_s_dadda_pg_rca32_u_pg_rca_or4_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and5_f_s_dadda_pg_rca32_u_pg_rca_or4_y0 = f_s_dadda_pg_rca32_u_pg_rca_or4_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and5_f_s_dadda_pg_rca32_u_pg_rca_fa5_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa5_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and5_y0 = f_s_dadda_pg_rca32_u_pg_rca_and5_f_s_dadda_pg_rca32_u_pg_rca_or4_y0 & f_s_dadda_pg_rca32_u_pg_rca_and5_f_s_dadda_pg_rca32_u_pg_rca_fa5_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or5_f_s_dadda_pg_rca32_u_pg_rca_and5_y0 = f_s_dadda_pg_rca32_u_pg_rca_and5_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or5_f_s_dadda_pg_rca32_u_pg_rca_fa5_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa5_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or5_y0 = f_s_dadda_pg_rca32_u_pg_rca_or5_f_s_dadda_pg_rca32_u_pg_rca_and5_y0 | f_s_dadda_pg_rca32_u_pg_rca_or5_f_s_dadda_pg_rca32_u_pg_rca_fa5_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_fa787_y2 = f_s_dadda_pg_rca32_fa787_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_fa845_y2 = f_s_dadda_pg_rca32_fa845_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_u_pg_rca_or5_y0 = f_s_dadda_pg_rca32_u_pg_rca_or5_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa6_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_fa787_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_fa845_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa6_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_fa787_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_fa845_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa6_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa6_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa6_f_s_dadda_pg_rca32_u_pg_rca_or5_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and6_f_s_dadda_pg_rca32_u_pg_rca_or5_y0 = f_s_dadda_pg_rca32_u_pg_rca_or5_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and6_f_s_dadda_pg_rca32_u_pg_rca_fa6_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa6_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and6_y0 = f_s_dadda_pg_rca32_u_pg_rca_and6_f_s_dadda_pg_rca32_u_pg_rca_or5_y0 & f_s_dadda_pg_rca32_u_pg_rca_and6_f_s_dadda_pg_rca32_u_pg_rca_fa6_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or6_f_s_dadda_pg_rca32_u_pg_rca_and6_y0 = f_s_dadda_pg_rca32_u_pg_rca_and6_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or6_f_s_dadda_pg_rca32_u_pg_rca_fa6_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa6_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or6_y0 = f_s_dadda_pg_rca32_u_pg_rca_or6_f_s_dadda_pg_rca32_u_pg_rca_and6_y0 | f_s_dadda_pg_rca32_u_pg_rca_or6_f_s_dadda_pg_rca32_u_pg_rca_fa6_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_fa788_y2 = f_s_dadda_pg_rca32_fa788_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_fa846_y2 = f_s_dadda_pg_rca32_fa846_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_u_pg_rca_or6_y0 = f_s_dadda_pg_rca32_u_pg_rca_or6_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa7_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_fa788_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_fa846_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa7_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_fa788_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_fa846_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa7_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa7_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa7_f_s_dadda_pg_rca32_u_pg_rca_or6_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and7_f_s_dadda_pg_rca32_u_pg_rca_or6_y0 = f_s_dadda_pg_rca32_u_pg_rca_or6_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and7_f_s_dadda_pg_rca32_u_pg_rca_fa7_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa7_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and7_y0 = f_s_dadda_pg_rca32_u_pg_rca_and7_f_s_dadda_pg_rca32_u_pg_rca_or6_y0 & f_s_dadda_pg_rca32_u_pg_rca_and7_f_s_dadda_pg_rca32_u_pg_rca_fa7_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or7_f_s_dadda_pg_rca32_u_pg_rca_and7_y0 = f_s_dadda_pg_rca32_u_pg_rca_and7_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or7_f_s_dadda_pg_rca32_u_pg_rca_fa7_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa7_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or7_y0 = f_s_dadda_pg_rca32_u_pg_rca_or7_f_s_dadda_pg_rca32_u_pg_rca_and7_y0 | f_s_dadda_pg_rca32_u_pg_rca_or7_f_s_dadda_pg_rca32_u_pg_rca_fa7_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_fa789_y2 = f_s_dadda_pg_rca32_fa789_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_fa847_y2 = f_s_dadda_pg_rca32_fa847_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_u_pg_rca_or7_y0 = f_s_dadda_pg_rca32_u_pg_rca_or7_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa8_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_fa789_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_fa847_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa8_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_fa789_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_fa847_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa8_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa8_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa8_f_s_dadda_pg_rca32_u_pg_rca_or7_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and8_f_s_dadda_pg_rca32_u_pg_rca_or7_y0 = f_s_dadda_pg_rca32_u_pg_rca_or7_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and8_f_s_dadda_pg_rca32_u_pg_rca_fa8_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa8_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and8_y0 = f_s_dadda_pg_rca32_u_pg_rca_and8_f_s_dadda_pg_rca32_u_pg_rca_or7_y0 & f_s_dadda_pg_rca32_u_pg_rca_and8_f_s_dadda_pg_rca32_u_pg_rca_fa8_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or8_f_s_dadda_pg_rca32_u_pg_rca_and8_y0 = f_s_dadda_pg_rca32_u_pg_rca_and8_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or8_f_s_dadda_pg_rca32_u_pg_rca_fa8_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa8_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or8_y0 = f_s_dadda_pg_rca32_u_pg_rca_or8_f_s_dadda_pg_rca32_u_pg_rca_and8_y0 | f_s_dadda_pg_rca32_u_pg_rca_or8_f_s_dadda_pg_rca32_u_pg_rca_fa8_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_fa790_y2 = f_s_dadda_pg_rca32_fa790_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_fa848_y2 = f_s_dadda_pg_rca32_fa848_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_u_pg_rca_or8_y0 = f_s_dadda_pg_rca32_u_pg_rca_or8_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa9_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_fa790_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_fa848_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa9_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_fa790_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_fa848_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa9_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa9_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa9_f_s_dadda_pg_rca32_u_pg_rca_or8_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and9_f_s_dadda_pg_rca32_u_pg_rca_or8_y0 = f_s_dadda_pg_rca32_u_pg_rca_or8_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and9_f_s_dadda_pg_rca32_u_pg_rca_fa9_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa9_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and9_y0 = f_s_dadda_pg_rca32_u_pg_rca_and9_f_s_dadda_pg_rca32_u_pg_rca_or8_y0 & f_s_dadda_pg_rca32_u_pg_rca_and9_f_s_dadda_pg_rca32_u_pg_rca_fa9_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or9_f_s_dadda_pg_rca32_u_pg_rca_and9_y0 = f_s_dadda_pg_rca32_u_pg_rca_and9_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or9_f_s_dadda_pg_rca32_u_pg_rca_fa9_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa9_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or9_y0 = f_s_dadda_pg_rca32_u_pg_rca_or9_f_s_dadda_pg_rca32_u_pg_rca_and9_y0 | f_s_dadda_pg_rca32_u_pg_rca_or9_f_s_dadda_pg_rca32_u_pg_rca_fa9_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_fa791_y2 = f_s_dadda_pg_rca32_fa791_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_fa849_y2 = f_s_dadda_pg_rca32_fa849_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_u_pg_rca_or9_y0 = f_s_dadda_pg_rca32_u_pg_rca_or9_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa10_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_fa791_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_fa849_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa10_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_fa791_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_fa849_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa10_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa10_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa10_f_s_dadda_pg_rca32_u_pg_rca_or9_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and10_f_s_dadda_pg_rca32_u_pg_rca_or9_y0 = f_s_dadda_pg_rca32_u_pg_rca_or9_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and10_f_s_dadda_pg_rca32_u_pg_rca_fa10_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa10_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and10_y0 = f_s_dadda_pg_rca32_u_pg_rca_and10_f_s_dadda_pg_rca32_u_pg_rca_or9_y0 & f_s_dadda_pg_rca32_u_pg_rca_and10_f_s_dadda_pg_rca32_u_pg_rca_fa10_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or10_f_s_dadda_pg_rca32_u_pg_rca_and10_y0 = f_s_dadda_pg_rca32_u_pg_rca_and10_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or10_f_s_dadda_pg_rca32_u_pg_rca_fa10_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa10_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or10_y0 = f_s_dadda_pg_rca32_u_pg_rca_or10_f_s_dadda_pg_rca32_u_pg_rca_and10_y0 | f_s_dadda_pg_rca32_u_pg_rca_or10_f_s_dadda_pg_rca32_u_pg_rca_fa10_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_fa792_y2 = f_s_dadda_pg_rca32_fa792_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_fa850_y2 = f_s_dadda_pg_rca32_fa850_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_u_pg_rca_or10_y0 = f_s_dadda_pg_rca32_u_pg_rca_or10_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa11_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_fa792_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_fa850_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa11_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_fa792_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_fa850_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa11_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa11_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa11_f_s_dadda_pg_rca32_u_pg_rca_or10_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and11_f_s_dadda_pg_rca32_u_pg_rca_or10_y0 = f_s_dadda_pg_rca32_u_pg_rca_or10_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and11_f_s_dadda_pg_rca32_u_pg_rca_fa11_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa11_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and11_y0 = f_s_dadda_pg_rca32_u_pg_rca_and11_f_s_dadda_pg_rca32_u_pg_rca_or10_y0 & f_s_dadda_pg_rca32_u_pg_rca_and11_f_s_dadda_pg_rca32_u_pg_rca_fa11_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or11_f_s_dadda_pg_rca32_u_pg_rca_and11_y0 = f_s_dadda_pg_rca32_u_pg_rca_and11_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or11_f_s_dadda_pg_rca32_u_pg_rca_fa11_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa11_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or11_y0 = f_s_dadda_pg_rca32_u_pg_rca_or11_f_s_dadda_pg_rca32_u_pg_rca_and11_y0 | f_s_dadda_pg_rca32_u_pg_rca_or11_f_s_dadda_pg_rca32_u_pg_rca_fa11_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_fa793_y2 = f_s_dadda_pg_rca32_fa793_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_fa851_y2 = f_s_dadda_pg_rca32_fa851_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_u_pg_rca_or11_y0 = f_s_dadda_pg_rca32_u_pg_rca_or11_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa12_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_fa793_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_fa851_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa12_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_fa793_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_fa851_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa12_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa12_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa12_f_s_dadda_pg_rca32_u_pg_rca_or11_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and12_f_s_dadda_pg_rca32_u_pg_rca_or11_y0 = f_s_dadda_pg_rca32_u_pg_rca_or11_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and12_f_s_dadda_pg_rca32_u_pg_rca_fa12_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa12_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and12_y0 = f_s_dadda_pg_rca32_u_pg_rca_and12_f_s_dadda_pg_rca32_u_pg_rca_or11_y0 & f_s_dadda_pg_rca32_u_pg_rca_and12_f_s_dadda_pg_rca32_u_pg_rca_fa12_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or12_f_s_dadda_pg_rca32_u_pg_rca_and12_y0 = f_s_dadda_pg_rca32_u_pg_rca_and12_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or12_f_s_dadda_pg_rca32_u_pg_rca_fa12_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa12_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or12_y0 = f_s_dadda_pg_rca32_u_pg_rca_or12_f_s_dadda_pg_rca32_u_pg_rca_and12_y0 | f_s_dadda_pg_rca32_u_pg_rca_or12_f_s_dadda_pg_rca32_u_pg_rca_fa12_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_fa794_y2 = f_s_dadda_pg_rca32_fa794_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_fa852_y2 = f_s_dadda_pg_rca32_fa852_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_u_pg_rca_or12_y0 = f_s_dadda_pg_rca32_u_pg_rca_or12_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa13_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_fa794_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_fa852_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa13_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_fa794_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_fa852_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa13_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa13_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa13_f_s_dadda_pg_rca32_u_pg_rca_or12_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and13_f_s_dadda_pg_rca32_u_pg_rca_or12_y0 = f_s_dadda_pg_rca32_u_pg_rca_or12_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and13_f_s_dadda_pg_rca32_u_pg_rca_fa13_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa13_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and13_y0 = f_s_dadda_pg_rca32_u_pg_rca_and13_f_s_dadda_pg_rca32_u_pg_rca_or12_y0 & f_s_dadda_pg_rca32_u_pg_rca_and13_f_s_dadda_pg_rca32_u_pg_rca_fa13_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or13_f_s_dadda_pg_rca32_u_pg_rca_and13_y0 = f_s_dadda_pg_rca32_u_pg_rca_and13_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or13_f_s_dadda_pg_rca32_u_pg_rca_fa13_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa13_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or13_y0 = f_s_dadda_pg_rca32_u_pg_rca_or13_f_s_dadda_pg_rca32_u_pg_rca_and13_y0 | f_s_dadda_pg_rca32_u_pg_rca_or13_f_s_dadda_pg_rca32_u_pg_rca_fa13_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_fa795_y2 = f_s_dadda_pg_rca32_fa795_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_fa853_y2 = f_s_dadda_pg_rca32_fa853_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_u_pg_rca_or13_y0 = f_s_dadda_pg_rca32_u_pg_rca_or13_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa14_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_fa795_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_fa853_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa14_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_fa795_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_fa853_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa14_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa14_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa14_f_s_dadda_pg_rca32_u_pg_rca_or13_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and14_f_s_dadda_pg_rca32_u_pg_rca_or13_y0 = f_s_dadda_pg_rca32_u_pg_rca_or13_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and14_f_s_dadda_pg_rca32_u_pg_rca_fa14_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa14_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and14_y0 = f_s_dadda_pg_rca32_u_pg_rca_and14_f_s_dadda_pg_rca32_u_pg_rca_or13_y0 & f_s_dadda_pg_rca32_u_pg_rca_and14_f_s_dadda_pg_rca32_u_pg_rca_fa14_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or14_f_s_dadda_pg_rca32_u_pg_rca_and14_y0 = f_s_dadda_pg_rca32_u_pg_rca_and14_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or14_f_s_dadda_pg_rca32_u_pg_rca_fa14_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa14_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or14_y0 = f_s_dadda_pg_rca32_u_pg_rca_or14_f_s_dadda_pg_rca32_u_pg_rca_and14_y0 | f_s_dadda_pg_rca32_u_pg_rca_or14_f_s_dadda_pg_rca32_u_pg_rca_fa14_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_fa796_y2 = f_s_dadda_pg_rca32_fa796_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_fa854_y2 = f_s_dadda_pg_rca32_fa854_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_u_pg_rca_or14_y0 = f_s_dadda_pg_rca32_u_pg_rca_or14_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa15_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_fa796_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_fa854_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa15_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_fa796_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_fa854_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa15_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa15_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa15_f_s_dadda_pg_rca32_u_pg_rca_or14_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and15_f_s_dadda_pg_rca32_u_pg_rca_or14_y0 = f_s_dadda_pg_rca32_u_pg_rca_or14_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and15_f_s_dadda_pg_rca32_u_pg_rca_fa15_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa15_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and15_y0 = f_s_dadda_pg_rca32_u_pg_rca_and15_f_s_dadda_pg_rca32_u_pg_rca_or14_y0 & f_s_dadda_pg_rca32_u_pg_rca_and15_f_s_dadda_pg_rca32_u_pg_rca_fa15_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or15_f_s_dadda_pg_rca32_u_pg_rca_and15_y0 = f_s_dadda_pg_rca32_u_pg_rca_and15_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or15_f_s_dadda_pg_rca32_u_pg_rca_fa15_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa15_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or15_y0 = f_s_dadda_pg_rca32_u_pg_rca_or15_f_s_dadda_pg_rca32_u_pg_rca_and15_y0 | f_s_dadda_pg_rca32_u_pg_rca_or15_f_s_dadda_pg_rca32_u_pg_rca_fa15_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_fa797_y2 = f_s_dadda_pg_rca32_fa797_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_fa855_y2 = f_s_dadda_pg_rca32_fa855_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_u_pg_rca_or15_y0 = f_s_dadda_pg_rca32_u_pg_rca_or15_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa16_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_fa797_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_fa855_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa16_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_fa797_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_fa855_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa16_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa16_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa16_f_s_dadda_pg_rca32_u_pg_rca_or15_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and16_f_s_dadda_pg_rca32_u_pg_rca_or15_y0 = f_s_dadda_pg_rca32_u_pg_rca_or15_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and16_f_s_dadda_pg_rca32_u_pg_rca_fa16_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa16_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and16_y0 = f_s_dadda_pg_rca32_u_pg_rca_and16_f_s_dadda_pg_rca32_u_pg_rca_or15_y0 & f_s_dadda_pg_rca32_u_pg_rca_and16_f_s_dadda_pg_rca32_u_pg_rca_fa16_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or16_f_s_dadda_pg_rca32_u_pg_rca_and16_y0 = f_s_dadda_pg_rca32_u_pg_rca_and16_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or16_f_s_dadda_pg_rca32_u_pg_rca_fa16_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa16_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or16_y0 = f_s_dadda_pg_rca32_u_pg_rca_or16_f_s_dadda_pg_rca32_u_pg_rca_and16_y0 | f_s_dadda_pg_rca32_u_pg_rca_or16_f_s_dadda_pg_rca32_u_pg_rca_fa16_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_fa798_y2 = f_s_dadda_pg_rca32_fa798_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_fa856_y2 = f_s_dadda_pg_rca32_fa856_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_u_pg_rca_or16_y0 = f_s_dadda_pg_rca32_u_pg_rca_or16_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa17_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_fa798_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_fa856_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa17_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_fa798_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_fa856_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa17_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa17_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa17_f_s_dadda_pg_rca32_u_pg_rca_or16_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and17_f_s_dadda_pg_rca32_u_pg_rca_or16_y0 = f_s_dadda_pg_rca32_u_pg_rca_or16_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and17_f_s_dadda_pg_rca32_u_pg_rca_fa17_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa17_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and17_y0 = f_s_dadda_pg_rca32_u_pg_rca_and17_f_s_dadda_pg_rca32_u_pg_rca_or16_y0 & f_s_dadda_pg_rca32_u_pg_rca_and17_f_s_dadda_pg_rca32_u_pg_rca_fa17_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or17_f_s_dadda_pg_rca32_u_pg_rca_and17_y0 = f_s_dadda_pg_rca32_u_pg_rca_and17_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or17_f_s_dadda_pg_rca32_u_pg_rca_fa17_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa17_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or17_y0 = f_s_dadda_pg_rca32_u_pg_rca_or17_f_s_dadda_pg_rca32_u_pg_rca_and17_y0 | f_s_dadda_pg_rca32_u_pg_rca_or17_f_s_dadda_pg_rca32_u_pg_rca_fa17_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_fa799_y2 = f_s_dadda_pg_rca32_fa799_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_fa857_y2 = f_s_dadda_pg_rca32_fa857_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_u_pg_rca_or17_y0 = f_s_dadda_pg_rca32_u_pg_rca_or17_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa18_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_fa799_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_fa857_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa18_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_fa799_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_fa857_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa18_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa18_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa18_f_s_dadda_pg_rca32_u_pg_rca_or17_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and18_f_s_dadda_pg_rca32_u_pg_rca_or17_y0 = f_s_dadda_pg_rca32_u_pg_rca_or17_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and18_f_s_dadda_pg_rca32_u_pg_rca_fa18_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa18_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and18_y0 = f_s_dadda_pg_rca32_u_pg_rca_and18_f_s_dadda_pg_rca32_u_pg_rca_or17_y0 & f_s_dadda_pg_rca32_u_pg_rca_and18_f_s_dadda_pg_rca32_u_pg_rca_fa18_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or18_f_s_dadda_pg_rca32_u_pg_rca_and18_y0 = f_s_dadda_pg_rca32_u_pg_rca_and18_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or18_f_s_dadda_pg_rca32_u_pg_rca_fa18_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa18_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or18_y0 = f_s_dadda_pg_rca32_u_pg_rca_or18_f_s_dadda_pg_rca32_u_pg_rca_and18_y0 | f_s_dadda_pg_rca32_u_pg_rca_or18_f_s_dadda_pg_rca32_u_pg_rca_fa18_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_fa800_y2 = f_s_dadda_pg_rca32_fa800_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_fa858_y2 = f_s_dadda_pg_rca32_fa858_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_u_pg_rca_or18_y0 = f_s_dadda_pg_rca32_u_pg_rca_or18_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa19_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_fa800_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_fa858_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa19_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_fa800_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_fa858_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa19_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa19_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa19_f_s_dadda_pg_rca32_u_pg_rca_or18_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and19_f_s_dadda_pg_rca32_u_pg_rca_or18_y0 = f_s_dadda_pg_rca32_u_pg_rca_or18_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and19_f_s_dadda_pg_rca32_u_pg_rca_fa19_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa19_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and19_y0 = f_s_dadda_pg_rca32_u_pg_rca_and19_f_s_dadda_pg_rca32_u_pg_rca_or18_y0 & f_s_dadda_pg_rca32_u_pg_rca_and19_f_s_dadda_pg_rca32_u_pg_rca_fa19_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or19_f_s_dadda_pg_rca32_u_pg_rca_and19_y0 = f_s_dadda_pg_rca32_u_pg_rca_and19_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or19_f_s_dadda_pg_rca32_u_pg_rca_fa19_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa19_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or19_y0 = f_s_dadda_pg_rca32_u_pg_rca_or19_f_s_dadda_pg_rca32_u_pg_rca_and19_y0 | f_s_dadda_pg_rca32_u_pg_rca_or19_f_s_dadda_pg_rca32_u_pg_rca_fa19_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_fa801_y2 = f_s_dadda_pg_rca32_fa801_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_fa859_y2 = f_s_dadda_pg_rca32_fa859_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_u_pg_rca_or19_y0 = f_s_dadda_pg_rca32_u_pg_rca_or19_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa20_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_fa801_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_fa859_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa20_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_fa801_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_fa859_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa20_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa20_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa20_f_s_dadda_pg_rca32_u_pg_rca_or19_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and20_f_s_dadda_pg_rca32_u_pg_rca_or19_y0 = f_s_dadda_pg_rca32_u_pg_rca_or19_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and20_f_s_dadda_pg_rca32_u_pg_rca_fa20_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa20_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and20_y0 = f_s_dadda_pg_rca32_u_pg_rca_and20_f_s_dadda_pg_rca32_u_pg_rca_or19_y0 & f_s_dadda_pg_rca32_u_pg_rca_and20_f_s_dadda_pg_rca32_u_pg_rca_fa20_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or20_f_s_dadda_pg_rca32_u_pg_rca_and20_y0 = f_s_dadda_pg_rca32_u_pg_rca_and20_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or20_f_s_dadda_pg_rca32_u_pg_rca_fa20_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa20_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or20_y0 = f_s_dadda_pg_rca32_u_pg_rca_or20_f_s_dadda_pg_rca32_u_pg_rca_and20_y0 | f_s_dadda_pg_rca32_u_pg_rca_or20_f_s_dadda_pg_rca32_u_pg_rca_fa20_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_fa802_y2 = f_s_dadda_pg_rca32_fa802_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_fa860_y2 = f_s_dadda_pg_rca32_fa860_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_u_pg_rca_or20_y0 = f_s_dadda_pg_rca32_u_pg_rca_or20_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa21_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_fa802_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_fa860_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa21_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_fa802_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_fa860_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa21_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa21_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa21_f_s_dadda_pg_rca32_u_pg_rca_or20_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and21_f_s_dadda_pg_rca32_u_pg_rca_or20_y0 = f_s_dadda_pg_rca32_u_pg_rca_or20_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and21_f_s_dadda_pg_rca32_u_pg_rca_fa21_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa21_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and21_y0 = f_s_dadda_pg_rca32_u_pg_rca_and21_f_s_dadda_pg_rca32_u_pg_rca_or20_y0 & f_s_dadda_pg_rca32_u_pg_rca_and21_f_s_dadda_pg_rca32_u_pg_rca_fa21_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or21_f_s_dadda_pg_rca32_u_pg_rca_and21_y0 = f_s_dadda_pg_rca32_u_pg_rca_and21_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or21_f_s_dadda_pg_rca32_u_pg_rca_fa21_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa21_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or21_y0 = f_s_dadda_pg_rca32_u_pg_rca_or21_f_s_dadda_pg_rca32_u_pg_rca_and21_y0 | f_s_dadda_pg_rca32_u_pg_rca_or21_f_s_dadda_pg_rca32_u_pg_rca_fa21_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_fa803_y2 = f_s_dadda_pg_rca32_fa803_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_fa861_y2 = f_s_dadda_pg_rca32_fa861_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_u_pg_rca_or21_y0 = f_s_dadda_pg_rca32_u_pg_rca_or21_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa22_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_fa803_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_fa861_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa22_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_fa803_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_fa861_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa22_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa22_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa22_f_s_dadda_pg_rca32_u_pg_rca_or21_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and22_f_s_dadda_pg_rca32_u_pg_rca_or21_y0 = f_s_dadda_pg_rca32_u_pg_rca_or21_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and22_f_s_dadda_pg_rca32_u_pg_rca_fa22_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa22_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and22_y0 = f_s_dadda_pg_rca32_u_pg_rca_and22_f_s_dadda_pg_rca32_u_pg_rca_or21_y0 & f_s_dadda_pg_rca32_u_pg_rca_and22_f_s_dadda_pg_rca32_u_pg_rca_fa22_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or22_f_s_dadda_pg_rca32_u_pg_rca_and22_y0 = f_s_dadda_pg_rca32_u_pg_rca_and22_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or22_f_s_dadda_pg_rca32_u_pg_rca_fa22_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa22_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or22_y0 = f_s_dadda_pg_rca32_u_pg_rca_or22_f_s_dadda_pg_rca32_u_pg_rca_and22_y0 | f_s_dadda_pg_rca32_u_pg_rca_or22_f_s_dadda_pg_rca32_u_pg_rca_fa22_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_fa804_y2 = f_s_dadda_pg_rca32_fa804_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_fa862_y2 = f_s_dadda_pg_rca32_fa862_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_u_pg_rca_or22_y0 = f_s_dadda_pg_rca32_u_pg_rca_or22_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa23_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_fa804_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_fa862_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa23_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_fa804_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_fa862_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa23_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa23_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa23_f_s_dadda_pg_rca32_u_pg_rca_or22_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and23_f_s_dadda_pg_rca32_u_pg_rca_or22_y0 = f_s_dadda_pg_rca32_u_pg_rca_or22_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and23_f_s_dadda_pg_rca32_u_pg_rca_fa23_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa23_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and23_y0 = f_s_dadda_pg_rca32_u_pg_rca_and23_f_s_dadda_pg_rca32_u_pg_rca_or22_y0 & f_s_dadda_pg_rca32_u_pg_rca_and23_f_s_dadda_pg_rca32_u_pg_rca_fa23_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or23_f_s_dadda_pg_rca32_u_pg_rca_and23_y0 = f_s_dadda_pg_rca32_u_pg_rca_and23_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or23_f_s_dadda_pg_rca32_u_pg_rca_fa23_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa23_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or23_y0 = f_s_dadda_pg_rca32_u_pg_rca_or23_f_s_dadda_pg_rca32_u_pg_rca_and23_y0 | f_s_dadda_pg_rca32_u_pg_rca_or23_f_s_dadda_pg_rca32_u_pg_rca_fa23_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_fa805_y2 = f_s_dadda_pg_rca32_fa805_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_fa863_y2 = f_s_dadda_pg_rca32_fa863_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_u_pg_rca_or23_y0 = f_s_dadda_pg_rca32_u_pg_rca_or23_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa24_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_fa805_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_fa863_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa24_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_fa805_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_fa863_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa24_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa24_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa24_f_s_dadda_pg_rca32_u_pg_rca_or23_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and24_f_s_dadda_pg_rca32_u_pg_rca_or23_y0 = f_s_dadda_pg_rca32_u_pg_rca_or23_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and24_f_s_dadda_pg_rca32_u_pg_rca_fa24_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa24_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and24_y0 = f_s_dadda_pg_rca32_u_pg_rca_and24_f_s_dadda_pg_rca32_u_pg_rca_or23_y0 & f_s_dadda_pg_rca32_u_pg_rca_and24_f_s_dadda_pg_rca32_u_pg_rca_fa24_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or24_f_s_dadda_pg_rca32_u_pg_rca_and24_y0 = f_s_dadda_pg_rca32_u_pg_rca_and24_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or24_f_s_dadda_pg_rca32_u_pg_rca_fa24_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa24_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or24_y0 = f_s_dadda_pg_rca32_u_pg_rca_or24_f_s_dadda_pg_rca32_u_pg_rca_and24_y0 | f_s_dadda_pg_rca32_u_pg_rca_or24_f_s_dadda_pg_rca32_u_pg_rca_fa24_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_fa806_y2 = f_s_dadda_pg_rca32_fa806_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_fa864_y2 = f_s_dadda_pg_rca32_fa864_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_u_pg_rca_or24_y0 = f_s_dadda_pg_rca32_u_pg_rca_or24_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa25_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_fa806_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_fa864_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa25_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_fa806_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_fa864_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa25_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa25_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa25_f_s_dadda_pg_rca32_u_pg_rca_or24_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and25_f_s_dadda_pg_rca32_u_pg_rca_or24_y0 = f_s_dadda_pg_rca32_u_pg_rca_or24_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and25_f_s_dadda_pg_rca32_u_pg_rca_fa25_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa25_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and25_y0 = f_s_dadda_pg_rca32_u_pg_rca_and25_f_s_dadda_pg_rca32_u_pg_rca_or24_y0 & f_s_dadda_pg_rca32_u_pg_rca_and25_f_s_dadda_pg_rca32_u_pg_rca_fa25_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or25_f_s_dadda_pg_rca32_u_pg_rca_and25_y0 = f_s_dadda_pg_rca32_u_pg_rca_and25_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or25_f_s_dadda_pg_rca32_u_pg_rca_fa25_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa25_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or25_y0 = f_s_dadda_pg_rca32_u_pg_rca_or25_f_s_dadda_pg_rca32_u_pg_rca_and25_y0 | f_s_dadda_pg_rca32_u_pg_rca_or25_f_s_dadda_pg_rca32_u_pg_rca_fa25_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_fa807_y2 = f_s_dadda_pg_rca32_fa807_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_fa865_y2 = f_s_dadda_pg_rca32_fa865_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_u_pg_rca_or25_y0 = f_s_dadda_pg_rca32_u_pg_rca_or25_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa26_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_fa807_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_fa865_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa26_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_fa807_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_fa865_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa26_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa26_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa26_f_s_dadda_pg_rca32_u_pg_rca_or25_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and26_f_s_dadda_pg_rca32_u_pg_rca_or25_y0 = f_s_dadda_pg_rca32_u_pg_rca_or25_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and26_f_s_dadda_pg_rca32_u_pg_rca_fa26_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa26_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and26_y0 = f_s_dadda_pg_rca32_u_pg_rca_and26_f_s_dadda_pg_rca32_u_pg_rca_or25_y0 & f_s_dadda_pg_rca32_u_pg_rca_and26_f_s_dadda_pg_rca32_u_pg_rca_fa26_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or26_f_s_dadda_pg_rca32_u_pg_rca_and26_y0 = f_s_dadda_pg_rca32_u_pg_rca_and26_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or26_f_s_dadda_pg_rca32_u_pg_rca_fa26_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa26_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or26_y0 = f_s_dadda_pg_rca32_u_pg_rca_or26_f_s_dadda_pg_rca32_u_pg_rca_and26_y0 | f_s_dadda_pg_rca32_u_pg_rca_or26_f_s_dadda_pg_rca32_u_pg_rca_fa26_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_fa808_y2 = f_s_dadda_pg_rca32_fa808_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_fa866_y2 = f_s_dadda_pg_rca32_fa866_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_u_pg_rca_or26_y0 = f_s_dadda_pg_rca32_u_pg_rca_or26_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa27_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_fa808_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_fa866_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa27_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_fa808_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_fa866_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa27_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa27_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa27_f_s_dadda_pg_rca32_u_pg_rca_or26_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and27_f_s_dadda_pg_rca32_u_pg_rca_or26_y0 = f_s_dadda_pg_rca32_u_pg_rca_or26_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and27_f_s_dadda_pg_rca32_u_pg_rca_fa27_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa27_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and27_y0 = f_s_dadda_pg_rca32_u_pg_rca_and27_f_s_dadda_pg_rca32_u_pg_rca_or26_y0 & f_s_dadda_pg_rca32_u_pg_rca_and27_f_s_dadda_pg_rca32_u_pg_rca_fa27_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or27_f_s_dadda_pg_rca32_u_pg_rca_and27_y0 = f_s_dadda_pg_rca32_u_pg_rca_and27_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or27_f_s_dadda_pg_rca32_u_pg_rca_fa27_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa27_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or27_y0 = f_s_dadda_pg_rca32_u_pg_rca_or27_f_s_dadda_pg_rca32_u_pg_rca_and27_y0 | f_s_dadda_pg_rca32_u_pg_rca_or27_f_s_dadda_pg_rca32_u_pg_rca_fa27_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_fa809_y2 = f_s_dadda_pg_rca32_fa809_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_fa867_y2 = f_s_dadda_pg_rca32_fa867_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_u_pg_rca_or27_y0 = f_s_dadda_pg_rca32_u_pg_rca_or27_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa28_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_fa809_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_fa867_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa28_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_fa809_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_fa867_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa28_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa28_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa28_f_s_dadda_pg_rca32_u_pg_rca_or27_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and28_f_s_dadda_pg_rca32_u_pg_rca_or27_y0 = f_s_dadda_pg_rca32_u_pg_rca_or27_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and28_f_s_dadda_pg_rca32_u_pg_rca_fa28_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa28_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and28_y0 = f_s_dadda_pg_rca32_u_pg_rca_and28_f_s_dadda_pg_rca32_u_pg_rca_or27_y0 & f_s_dadda_pg_rca32_u_pg_rca_and28_f_s_dadda_pg_rca32_u_pg_rca_fa28_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or28_f_s_dadda_pg_rca32_u_pg_rca_and28_y0 = f_s_dadda_pg_rca32_u_pg_rca_and28_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or28_f_s_dadda_pg_rca32_u_pg_rca_fa28_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa28_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or28_y0 = f_s_dadda_pg_rca32_u_pg_rca_or28_f_s_dadda_pg_rca32_u_pg_rca_and28_y0 | f_s_dadda_pg_rca32_u_pg_rca_or28_f_s_dadda_pg_rca32_u_pg_rca_fa28_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_fa810_y2 = f_s_dadda_pg_rca32_fa810_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_fa868_y2 = f_s_dadda_pg_rca32_fa868_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_u_pg_rca_or28_y0 = f_s_dadda_pg_rca32_u_pg_rca_or28_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa29_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_fa810_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_fa868_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa29_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_fa810_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_fa868_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa29_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa29_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa29_f_s_dadda_pg_rca32_u_pg_rca_or28_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and29_f_s_dadda_pg_rca32_u_pg_rca_or28_y0 = f_s_dadda_pg_rca32_u_pg_rca_or28_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and29_f_s_dadda_pg_rca32_u_pg_rca_fa29_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and29_y0 = f_s_dadda_pg_rca32_u_pg_rca_and29_f_s_dadda_pg_rca32_u_pg_rca_or28_y0 & f_s_dadda_pg_rca32_u_pg_rca_and29_f_s_dadda_pg_rca32_u_pg_rca_fa29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or29_f_s_dadda_pg_rca32_u_pg_rca_and29_y0 = f_s_dadda_pg_rca32_u_pg_rca_and29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or29_f_s_dadda_pg_rca32_u_pg_rca_fa29_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa29_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or29_y0 = f_s_dadda_pg_rca32_u_pg_rca_or29_f_s_dadda_pg_rca32_u_pg_rca_and29_y0 | f_s_dadda_pg_rca32_u_pg_rca_or29_f_s_dadda_pg_rca32_u_pg_rca_fa29_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_fa811_y2 = f_s_dadda_pg_rca32_fa811_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_fa869_y2 = f_s_dadda_pg_rca32_fa869_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_u_pg_rca_or29_y0 = f_s_dadda_pg_rca32_u_pg_rca_or29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa30_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_fa811_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_fa869_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa30_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_fa811_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_fa869_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa30_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa30_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa30_f_s_dadda_pg_rca32_u_pg_rca_or29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and30_f_s_dadda_pg_rca32_u_pg_rca_or29_y0 = f_s_dadda_pg_rca32_u_pg_rca_or29_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and30_f_s_dadda_pg_rca32_u_pg_rca_fa30_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa30_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and30_y0 = f_s_dadda_pg_rca32_u_pg_rca_and30_f_s_dadda_pg_rca32_u_pg_rca_or29_y0 & f_s_dadda_pg_rca32_u_pg_rca_and30_f_s_dadda_pg_rca32_u_pg_rca_fa30_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or30_f_s_dadda_pg_rca32_u_pg_rca_and30_y0 = f_s_dadda_pg_rca32_u_pg_rca_and30_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or30_f_s_dadda_pg_rca32_u_pg_rca_fa30_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa30_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or30_y0 = f_s_dadda_pg_rca32_u_pg_rca_or30_f_s_dadda_pg_rca32_u_pg_rca_and30_y0 | f_s_dadda_pg_rca32_u_pg_rca_or30_f_s_dadda_pg_rca32_u_pg_rca_fa30_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_fa812_y2 = f_s_dadda_pg_rca32_fa812_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_fa870_y2 = f_s_dadda_pg_rca32_fa870_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_u_pg_rca_or30_y0 = f_s_dadda_pg_rca32_u_pg_rca_or30_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa31_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_fa812_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_fa870_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa31_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_fa812_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_fa870_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa31_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa31_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa31_f_s_dadda_pg_rca32_u_pg_rca_or30_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and31_f_s_dadda_pg_rca32_u_pg_rca_or30_y0 = f_s_dadda_pg_rca32_u_pg_rca_or30_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and31_f_s_dadda_pg_rca32_u_pg_rca_fa31_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and31_y0 = f_s_dadda_pg_rca32_u_pg_rca_and31_f_s_dadda_pg_rca32_u_pg_rca_or30_y0 & f_s_dadda_pg_rca32_u_pg_rca_and31_f_s_dadda_pg_rca32_u_pg_rca_fa31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or31_f_s_dadda_pg_rca32_u_pg_rca_and31_y0 = f_s_dadda_pg_rca32_u_pg_rca_and31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or31_f_s_dadda_pg_rca32_u_pg_rca_fa31_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa31_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or31_y0 = f_s_dadda_pg_rca32_u_pg_rca_or31_f_s_dadda_pg_rca32_u_pg_rca_and31_y0 | f_s_dadda_pg_rca32_u_pg_rca_or31_f_s_dadda_pg_rca32_u_pg_rca_fa31_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_fa813_y2 = f_s_dadda_pg_rca32_fa813_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_fa871_y2 = f_s_dadda_pg_rca32_fa871_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_u_pg_rca_or31_y0 = f_s_dadda_pg_rca32_u_pg_rca_or31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa32_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_fa813_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_fa871_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa32_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_fa813_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_fa871_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa32_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa32_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa32_f_s_dadda_pg_rca32_u_pg_rca_or31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and32_f_s_dadda_pg_rca32_u_pg_rca_or31_y0 = f_s_dadda_pg_rca32_u_pg_rca_or31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and32_f_s_dadda_pg_rca32_u_pg_rca_fa32_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa32_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and32_y0 = f_s_dadda_pg_rca32_u_pg_rca_and32_f_s_dadda_pg_rca32_u_pg_rca_or31_y0 & f_s_dadda_pg_rca32_u_pg_rca_and32_f_s_dadda_pg_rca32_u_pg_rca_fa32_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or32_f_s_dadda_pg_rca32_u_pg_rca_and32_y0 = f_s_dadda_pg_rca32_u_pg_rca_and32_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or32_f_s_dadda_pg_rca32_u_pg_rca_fa32_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa32_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or32_y0 = f_s_dadda_pg_rca32_u_pg_rca_or32_f_s_dadda_pg_rca32_u_pg_rca_and32_y0 | f_s_dadda_pg_rca32_u_pg_rca_or32_f_s_dadda_pg_rca32_u_pg_rca_fa32_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_fa814_y2 = f_s_dadda_pg_rca32_fa814_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_fa872_y2 = f_s_dadda_pg_rca32_fa872_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_u_pg_rca_or32_y0 = f_s_dadda_pg_rca32_u_pg_rca_or32_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa33_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_fa814_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_fa872_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa33_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_fa814_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_fa872_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa33_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa33_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa33_f_s_dadda_pg_rca32_u_pg_rca_or32_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and33_f_s_dadda_pg_rca32_u_pg_rca_or32_y0 = f_s_dadda_pg_rca32_u_pg_rca_or32_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and33_f_s_dadda_pg_rca32_u_pg_rca_fa33_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa33_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and33_y0 = f_s_dadda_pg_rca32_u_pg_rca_and33_f_s_dadda_pg_rca32_u_pg_rca_or32_y0 & f_s_dadda_pg_rca32_u_pg_rca_and33_f_s_dadda_pg_rca32_u_pg_rca_fa33_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or33_f_s_dadda_pg_rca32_u_pg_rca_and33_y0 = f_s_dadda_pg_rca32_u_pg_rca_and33_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or33_f_s_dadda_pg_rca32_u_pg_rca_fa33_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa33_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or33_y0 = f_s_dadda_pg_rca32_u_pg_rca_or33_f_s_dadda_pg_rca32_u_pg_rca_and33_y0 | f_s_dadda_pg_rca32_u_pg_rca_or33_f_s_dadda_pg_rca32_u_pg_rca_fa33_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_fa815_y2 = f_s_dadda_pg_rca32_fa815_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_fa873_y2 = f_s_dadda_pg_rca32_fa873_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_u_pg_rca_or33_y0 = f_s_dadda_pg_rca32_u_pg_rca_or33_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa34_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_fa815_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_fa873_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa34_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_fa815_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_fa873_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa34_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa34_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa34_f_s_dadda_pg_rca32_u_pg_rca_or33_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and34_f_s_dadda_pg_rca32_u_pg_rca_or33_y0 = f_s_dadda_pg_rca32_u_pg_rca_or33_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and34_f_s_dadda_pg_rca32_u_pg_rca_fa34_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa34_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and34_y0 = f_s_dadda_pg_rca32_u_pg_rca_and34_f_s_dadda_pg_rca32_u_pg_rca_or33_y0 & f_s_dadda_pg_rca32_u_pg_rca_and34_f_s_dadda_pg_rca32_u_pg_rca_fa34_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or34_f_s_dadda_pg_rca32_u_pg_rca_and34_y0 = f_s_dadda_pg_rca32_u_pg_rca_and34_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or34_f_s_dadda_pg_rca32_u_pg_rca_fa34_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa34_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or34_y0 = f_s_dadda_pg_rca32_u_pg_rca_or34_f_s_dadda_pg_rca32_u_pg_rca_and34_y0 | f_s_dadda_pg_rca32_u_pg_rca_or34_f_s_dadda_pg_rca32_u_pg_rca_fa34_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_fa816_y2 = f_s_dadda_pg_rca32_fa816_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_fa874_y2 = f_s_dadda_pg_rca32_fa874_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_u_pg_rca_or34_y0 = f_s_dadda_pg_rca32_u_pg_rca_or34_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa35_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_fa816_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_fa874_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa35_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_fa816_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_fa874_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa35_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa35_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa35_f_s_dadda_pg_rca32_u_pg_rca_or34_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and35_f_s_dadda_pg_rca32_u_pg_rca_or34_y0 = f_s_dadda_pg_rca32_u_pg_rca_or34_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and35_f_s_dadda_pg_rca32_u_pg_rca_fa35_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa35_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and35_y0 = f_s_dadda_pg_rca32_u_pg_rca_and35_f_s_dadda_pg_rca32_u_pg_rca_or34_y0 & f_s_dadda_pg_rca32_u_pg_rca_and35_f_s_dadda_pg_rca32_u_pg_rca_fa35_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or35_f_s_dadda_pg_rca32_u_pg_rca_and35_y0 = f_s_dadda_pg_rca32_u_pg_rca_and35_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or35_f_s_dadda_pg_rca32_u_pg_rca_fa35_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa35_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or35_y0 = f_s_dadda_pg_rca32_u_pg_rca_or35_f_s_dadda_pg_rca32_u_pg_rca_and35_y0 | f_s_dadda_pg_rca32_u_pg_rca_or35_f_s_dadda_pg_rca32_u_pg_rca_fa35_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_fa817_y2 = f_s_dadda_pg_rca32_fa817_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_fa875_y2 = f_s_dadda_pg_rca32_fa875_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_u_pg_rca_or35_y0 = f_s_dadda_pg_rca32_u_pg_rca_or35_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa36_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_fa817_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_fa875_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa36_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_fa817_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_fa875_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa36_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa36_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa36_f_s_dadda_pg_rca32_u_pg_rca_or35_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and36_f_s_dadda_pg_rca32_u_pg_rca_or35_y0 = f_s_dadda_pg_rca32_u_pg_rca_or35_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and36_f_s_dadda_pg_rca32_u_pg_rca_fa36_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa36_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and36_y0 = f_s_dadda_pg_rca32_u_pg_rca_and36_f_s_dadda_pg_rca32_u_pg_rca_or35_y0 & f_s_dadda_pg_rca32_u_pg_rca_and36_f_s_dadda_pg_rca32_u_pg_rca_fa36_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or36_f_s_dadda_pg_rca32_u_pg_rca_and36_y0 = f_s_dadda_pg_rca32_u_pg_rca_and36_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or36_f_s_dadda_pg_rca32_u_pg_rca_fa36_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa36_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or36_y0 = f_s_dadda_pg_rca32_u_pg_rca_or36_f_s_dadda_pg_rca32_u_pg_rca_and36_y0 | f_s_dadda_pg_rca32_u_pg_rca_or36_f_s_dadda_pg_rca32_u_pg_rca_fa36_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_fa818_y2 = f_s_dadda_pg_rca32_fa818_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_fa876_y2 = f_s_dadda_pg_rca32_fa876_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_u_pg_rca_or36_y0 = f_s_dadda_pg_rca32_u_pg_rca_or36_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa37_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_fa818_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_fa876_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa37_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_fa818_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_fa876_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa37_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa37_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa37_f_s_dadda_pg_rca32_u_pg_rca_or36_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and37_f_s_dadda_pg_rca32_u_pg_rca_or36_y0 = f_s_dadda_pg_rca32_u_pg_rca_or36_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and37_f_s_dadda_pg_rca32_u_pg_rca_fa37_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa37_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and37_y0 = f_s_dadda_pg_rca32_u_pg_rca_and37_f_s_dadda_pg_rca32_u_pg_rca_or36_y0 & f_s_dadda_pg_rca32_u_pg_rca_and37_f_s_dadda_pg_rca32_u_pg_rca_fa37_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or37_f_s_dadda_pg_rca32_u_pg_rca_and37_y0 = f_s_dadda_pg_rca32_u_pg_rca_and37_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or37_f_s_dadda_pg_rca32_u_pg_rca_fa37_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa37_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or37_y0 = f_s_dadda_pg_rca32_u_pg_rca_or37_f_s_dadda_pg_rca32_u_pg_rca_and37_y0 | f_s_dadda_pg_rca32_u_pg_rca_or37_f_s_dadda_pg_rca32_u_pg_rca_fa37_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_fa819_y2 = f_s_dadda_pg_rca32_fa819_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_fa877_y2 = f_s_dadda_pg_rca32_fa877_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_u_pg_rca_or37_y0 = f_s_dadda_pg_rca32_u_pg_rca_or37_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa38_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_fa819_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_fa877_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa38_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_fa819_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_fa877_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa38_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa38_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa38_f_s_dadda_pg_rca32_u_pg_rca_or37_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and38_f_s_dadda_pg_rca32_u_pg_rca_or37_y0 = f_s_dadda_pg_rca32_u_pg_rca_or37_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and38_f_s_dadda_pg_rca32_u_pg_rca_fa38_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa38_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and38_y0 = f_s_dadda_pg_rca32_u_pg_rca_and38_f_s_dadda_pg_rca32_u_pg_rca_or37_y0 & f_s_dadda_pg_rca32_u_pg_rca_and38_f_s_dadda_pg_rca32_u_pg_rca_fa38_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or38_f_s_dadda_pg_rca32_u_pg_rca_and38_y0 = f_s_dadda_pg_rca32_u_pg_rca_and38_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or38_f_s_dadda_pg_rca32_u_pg_rca_fa38_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa38_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or38_y0 = f_s_dadda_pg_rca32_u_pg_rca_or38_f_s_dadda_pg_rca32_u_pg_rca_and38_y0 | f_s_dadda_pg_rca32_u_pg_rca_or38_f_s_dadda_pg_rca32_u_pg_rca_fa38_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_fa820_y2 = f_s_dadda_pg_rca32_fa820_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_fa878_y2 = f_s_dadda_pg_rca32_fa878_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_u_pg_rca_or38_y0 = f_s_dadda_pg_rca32_u_pg_rca_or38_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa39_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_fa820_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_fa878_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa39_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_fa820_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_fa878_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa39_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa39_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa39_f_s_dadda_pg_rca32_u_pg_rca_or38_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and39_f_s_dadda_pg_rca32_u_pg_rca_or38_y0 = f_s_dadda_pg_rca32_u_pg_rca_or38_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and39_f_s_dadda_pg_rca32_u_pg_rca_fa39_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa39_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and39_y0 = f_s_dadda_pg_rca32_u_pg_rca_and39_f_s_dadda_pg_rca32_u_pg_rca_or38_y0 & f_s_dadda_pg_rca32_u_pg_rca_and39_f_s_dadda_pg_rca32_u_pg_rca_fa39_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or39_f_s_dadda_pg_rca32_u_pg_rca_and39_y0 = f_s_dadda_pg_rca32_u_pg_rca_and39_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or39_f_s_dadda_pg_rca32_u_pg_rca_fa39_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa39_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or39_y0 = f_s_dadda_pg_rca32_u_pg_rca_or39_f_s_dadda_pg_rca32_u_pg_rca_and39_y0 | f_s_dadda_pg_rca32_u_pg_rca_or39_f_s_dadda_pg_rca32_u_pg_rca_fa39_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_fa821_y2 = f_s_dadda_pg_rca32_fa821_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_fa879_y2 = f_s_dadda_pg_rca32_fa879_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_u_pg_rca_or39_y0 = f_s_dadda_pg_rca32_u_pg_rca_or39_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa40_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_fa821_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_fa879_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa40_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_fa821_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_fa879_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa40_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa40_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa40_f_s_dadda_pg_rca32_u_pg_rca_or39_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and40_f_s_dadda_pg_rca32_u_pg_rca_or39_y0 = f_s_dadda_pg_rca32_u_pg_rca_or39_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and40_f_s_dadda_pg_rca32_u_pg_rca_fa40_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa40_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and40_y0 = f_s_dadda_pg_rca32_u_pg_rca_and40_f_s_dadda_pg_rca32_u_pg_rca_or39_y0 & f_s_dadda_pg_rca32_u_pg_rca_and40_f_s_dadda_pg_rca32_u_pg_rca_fa40_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or40_f_s_dadda_pg_rca32_u_pg_rca_and40_y0 = f_s_dadda_pg_rca32_u_pg_rca_and40_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or40_f_s_dadda_pg_rca32_u_pg_rca_fa40_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa40_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or40_y0 = f_s_dadda_pg_rca32_u_pg_rca_or40_f_s_dadda_pg_rca32_u_pg_rca_and40_y0 | f_s_dadda_pg_rca32_u_pg_rca_or40_f_s_dadda_pg_rca32_u_pg_rca_fa40_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_fa822_y2 = f_s_dadda_pg_rca32_fa822_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_fa880_y2 = f_s_dadda_pg_rca32_fa880_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_u_pg_rca_or40_y0 = f_s_dadda_pg_rca32_u_pg_rca_or40_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa41_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_fa822_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_fa880_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa41_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_fa822_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_fa880_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa41_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa41_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa41_f_s_dadda_pg_rca32_u_pg_rca_or40_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and41_f_s_dadda_pg_rca32_u_pg_rca_or40_y0 = f_s_dadda_pg_rca32_u_pg_rca_or40_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and41_f_s_dadda_pg_rca32_u_pg_rca_fa41_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa41_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and41_y0 = f_s_dadda_pg_rca32_u_pg_rca_and41_f_s_dadda_pg_rca32_u_pg_rca_or40_y0 & f_s_dadda_pg_rca32_u_pg_rca_and41_f_s_dadda_pg_rca32_u_pg_rca_fa41_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or41_f_s_dadda_pg_rca32_u_pg_rca_and41_y0 = f_s_dadda_pg_rca32_u_pg_rca_and41_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or41_f_s_dadda_pg_rca32_u_pg_rca_fa41_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa41_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or41_y0 = f_s_dadda_pg_rca32_u_pg_rca_or41_f_s_dadda_pg_rca32_u_pg_rca_and41_y0 | f_s_dadda_pg_rca32_u_pg_rca_or41_f_s_dadda_pg_rca32_u_pg_rca_fa41_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_fa823_y2 = f_s_dadda_pg_rca32_fa823_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_fa881_y2 = f_s_dadda_pg_rca32_fa881_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_u_pg_rca_or41_y0 = f_s_dadda_pg_rca32_u_pg_rca_or41_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa42_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_fa823_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_fa881_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa42_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_fa823_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_fa881_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa42_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa42_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa42_f_s_dadda_pg_rca32_u_pg_rca_or41_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and42_f_s_dadda_pg_rca32_u_pg_rca_or41_y0 = f_s_dadda_pg_rca32_u_pg_rca_or41_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and42_f_s_dadda_pg_rca32_u_pg_rca_fa42_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa42_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and42_y0 = f_s_dadda_pg_rca32_u_pg_rca_and42_f_s_dadda_pg_rca32_u_pg_rca_or41_y0 & f_s_dadda_pg_rca32_u_pg_rca_and42_f_s_dadda_pg_rca32_u_pg_rca_fa42_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or42_f_s_dadda_pg_rca32_u_pg_rca_and42_y0 = f_s_dadda_pg_rca32_u_pg_rca_and42_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or42_f_s_dadda_pg_rca32_u_pg_rca_fa42_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa42_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or42_y0 = f_s_dadda_pg_rca32_u_pg_rca_or42_f_s_dadda_pg_rca32_u_pg_rca_and42_y0 | f_s_dadda_pg_rca32_u_pg_rca_or42_f_s_dadda_pg_rca32_u_pg_rca_fa42_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_fa824_y2 = f_s_dadda_pg_rca32_fa824_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_fa882_y2 = f_s_dadda_pg_rca32_fa882_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_u_pg_rca_or42_y0 = f_s_dadda_pg_rca32_u_pg_rca_or42_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa43_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_fa824_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_fa882_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa43_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_fa824_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_fa882_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa43_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa43_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa43_f_s_dadda_pg_rca32_u_pg_rca_or42_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and43_f_s_dadda_pg_rca32_u_pg_rca_or42_y0 = f_s_dadda_pg_rca32_u_pg_rca_or42_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and43_f_s_dadda_pg_rca32_u_pg_rca_fa43_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa43_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and43_y0 = f_s_dadda_pg_rca32_u_pg_rca_and43_f_s_dadda_pg_rca32_u_pg_rca_or42_y0 & f_s_dadda_pg_rca32_u_pg_rca_and43_f_s_dadda_pg_rca32_u_pg_rca_fa43_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or43_f_s_dadda_pg_rca32_u_pg_rca_and43_y0 = f_s_dadda_pg_rca32_u_pg_rca_and43_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or43_f_s_dadda_pg_rca32_u_pg_rca_fa43_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa43_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or43_y0 = f_s_dadda_pg_rca32_u_pg_rca_or43_f_s_dadda_pg_rca32_u_pg_rca_and43_y0 | f_s_dadda_pg_rca32_u_pg_rca_or43_f_s_dadda_pg_rca32_u_pg_rca_fa43_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_fa825_y2 = f_s_dadda_pg_rca32_fa825_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_fa883_y2 = f_s_dadda_pg_rca32_fa883_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_u_pg_rca_or43_y0 = f_s_dadda_pg_rca32_u_pg_rca_or43_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa44_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_fa825_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_fa883_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa44_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_fa825_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_fa883_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa44_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa44_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa44_f_s_dadda_pg_rca32_u_pg_rca_or43_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and44_f_s_dadda_pg_rca32_u_pg_rca_or43_y0 = f_s_dadda_pg_rca32_u_pg_rca_or43_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and44_f_s_dadda_pg_rca32_u_pg_rca_fa44_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa44_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and44_y0 = f_s_dadda_pg_rca32_u_pg_rca_and44_f_s_dadda_pg_rca32_u_pg_rca_or43_y0 & f_s_dadda_pg_rca32_u_pg_rca_and44_f_s_dadda_pg_rca32_u_pg_rca_fa44_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or44_f_s_dadda_pg_rca32_u_pg_rca_and44_y0 = f_s_dadda_pg_rca32_u_pg_rca_and44_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or44_f_s_dadda_pg_rca32_u_pg_rca_fa44_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa44_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or44_y0 = f_s_dadda_pg_rca32_u_pg_rca_or44_f_s_dadda_pg_rca32_u_pg_rca_and44_y0 | f_s_dadda_pg_rca32_u_pg_rca_or44_f_s_dadda_pg_rca32_u_pg_rca_fa44_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_fa826_y2 = f_s_dadda_pg_rca32_fa826_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_fa884_y2 = f_s_dadda_pg_rca32_fa884_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_u_pg_rca_or44_y0 = f_s_dadda_pg_rca32_u_pg_rca_or44_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa45_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_fa826_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_fa884_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa45_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_fa826_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_fa884_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa45_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa45_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa45_f_s_dadda_pg_rca32_u_pg_rca_or44_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and45_f_s_dadda_pg_rca32_u_pg_rca_or44_y0 = f_s_dadda_pg_rca32_u_pg_rca_or44_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and45_f_s_dadda_pg_rca32_u_pg_rca_fa45_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa45_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and45_y0 = f_s_dadda_pg_rca32_u_pg_rca_and45_f_s_dadda_pg_rca32_u_pg_rca_or44_y0 & f_s_dadda_pg_rca32_u_pg_rca_and45_f_s_dadda_pg_rca32_u_pg_rca_fa45_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or45_f_s_dadda_pg_rca32_u_pg_rca_and45_y0 = f_s_dadda_pg_rca32_u_pg_rca_and45_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or45_f_s_dadda_pg_rca32_u_pg_rca_fa45_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa45_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or45_y0 = f_s_dadda_pg_rca32_u_pg_rca_or45_f_s_dadda_pg_rca32_u_pg_rca_and45_y0 | f_s_dadda_pg_rca32_u_pg_rca_or45_f_s_dadda_pg_rca32_u_pg_rca_fa45_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_fa827_y2 = f_s_dadda_pg_rca32_fa827_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_fa885_y2 = f_s_dadda_pg_rca32_fa885_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_u_pg_rca_or45_y0 = f_s_dadda_pg_rca32_u_pg_rca_or45_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa46_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_fa827_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_fa885_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa46_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_fa827_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_fa885_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa46_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa46_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa46_f_s_dadda_pg_rca32_u_pg_rca_or45_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and46_f_s_dadda_pg_rca32_u_pg_rca_or45_y0 = f_s_dadda_pg_rca32_u_pg_rca_or45_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and46_f_s_dadda_pg_rca32_u_pg_rca_fa46_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa46_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and46_y0 = f_s_dadda_pg_rca32_u_pg_rca_and46_f_s_dadda_pg_rca32_u_pg_rca_or45_y0 & f_s_dadda_pg_rca32_u_pg_rca_and46_f_s_dadda_pg_rca32_u_pg_rca_fa46_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or46_f_s_dadda_pg_rca32_u_pg_rca_and46_y0 = f_s_dadda_pg_rca32_u_pg_rca_and46_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or46_f_s_dadda_pg_rca32_u_pg_rca_fa46_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa46_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or46_y0 = f_s_dadda_pg_rca32_u_pg_rca_or46_f_s_dadda_pg_rca32_u_pg_rca_and46_y0 | f_s_dadda_pg_rca32_u_pg_rca_or46_f_s_dadda_pg_rca32_u_pg_rca_fa46_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_fa828_y2 = f_s_dadda_pg_rca32_fa828_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_fa886_y2 = f_s_dadda_pg_rca32_fa886_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_u_pg_rca_or46_y0 = f_s_dadda_pg_rca32_u_pg_rca_or46_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa47_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_fa828_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_fa886_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa47_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_fa828_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_fa886_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa47_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa47_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa47_f_s_dadda_pg_rca32_u_pg_rca_or46_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and47_f_s_dadda_pg_rca32_u_pg_rca_or46_y0 = f_s_dadda_pg_rca32_u_pg_rca_or46_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and47_f_s_dadda_pg_rca32_u_pg_rca_fa47_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa47_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and47_y0 = f_s_dadda_pg_rca32_u_pg_rca_and47_f_s_dadda_pg_rca32_u_pg_rca_or46_y0 & f_s_dadda_pg_rca32_u_pg_rca_and47_f_s_dadda_pg_rca32_u_pg_rca_fa47_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or47_f_s_dadda_pg_rca32_u_pg_rca_and47_y0 = f_s_dadda_pg_rca32_u_pg_rca_and47_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or47_f_s_dadda_pg_rca32_u_pg_rca_fa47_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa47_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or47_y0 = f_s_dadda_pg_rca32_u_pg_rca_or47_f_s_dadda_pg_rca32_u_pg_rca_and47_y0 | f_s_dadda_pg_rca32_u_pg_rca_or47_f_s_dadda_pg_rca32_u_pg_rca_fa47_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_fa829_y2 = f_s_dadda_pg_rca32_fa829_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_fa887_y2 = f_s_dadda_pg_rca32_fa887_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_u_pg_rca_or47_y0 = f_s_dadda_pg_rca32_u_pg_rca_or47_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa48_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_fa829_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_fa887_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa48_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_fa829_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_fa887_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa48_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa48_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa48_f_s_dadda_pg_rca32_u_pg_rca_or47_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and48_f_s_dadda_pg_rca32_u_pg_rca_or47_y0 = f_s_dadda_pg_rca32_u_pg_rca_or47_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and48_f_s_dadda_pg_rca32_u_pg_rca_fa48_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa48_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and48_y0 = f_s_dadda_pg_rca32_u_pg_rca_and48_f_s_dadda_pg_rca32_u_pg_rca_or47_y0 & f_s_dadda_pg_rca32_u_pg_rca_and48_f_s_dadda_pg_rca32_u_pg_rca_fa48_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or48_f_s_dadda_pg_rca32_u_pg_rca_and48_y0 = f_s_dadda_pg_rca32_u_pg_rca_and48_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or48_f_s_dadda_pg_rca32_u_pg_rca_fa48_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa48_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or48_y0 = f_s_dadda_pg_rca32_u_pg_rca_or48_f_s_dadda_pg_rca32_u_pg_rca_and48_y0 | f_s_dadda_pg_rca32_u_pg_rca_or48_f_s_dadda_pg_rca32_u_pg_rca_fa48_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_fa830_y2 = f_s_dadda_pg_rca32_fa830_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_fa888_y2 = f_s_dadda_pg_rca32_fa888_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_u_pg_rca_or48_y0 = f_s_dadda_pg_rca32_u_pg_rca_or48_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa49_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_fa830_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_fa888_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa49_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_fa830_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_fa888_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa49_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa49_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa49_f_s_dadda_pg_rca32_u_pg_rca_or48_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and49_f_s_dadda_pg_rca32_u_pg_rca_or48_y0 = f_s_dadda_pg_rca32_u_pg_rca_or48_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and49_f_s_dadda_pg_rca32_u_pg_rca_fa49_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa49_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and49_y0 = f_s_dadda_pg_rca32_u_pg_rca_and49_f_s_dadda_pg_rca32_u_pg_rca_or48_y0 & f_s_dadda_pg_rca32_u_pg_rca_and49_f_s_dadda_pg_rca32_u_pg_rca_fa49_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or49_f_s_dadda_pg_rca32_u_pg_rca_and49_y0 = f_s_dadda_pg_rca32_u_pg_rca_and49_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or49_f_s_dadda_pg_rca32_u_pg_rca_fa49_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa49_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or49_y0 = f_s_dadda_pg_rca32_u_pg_rca_or49_f_s_dadda_pg_rca32_u_pg_rca_and49_y0 | f_s_dadda_pg_rca32_u_pg_rca_or49_f_s_dadda_pg_rca32_u_pg_rca_fa49_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_fa831_y2 = f_s_dadda_pg_rca32_fa831_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_fa889_y2 = f_s_dadda_pg_rca32_fa889_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_u_pg_rca_or49_y0 = f_s_dadda_pg_rca32_u_pg_rca_or49_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa50_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_fa831_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_fa889_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa50_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_fa831_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_fa889_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa50_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa50_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa50_f_s_dadda_pg_rca32_u_pg_rca_or49_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and50_f_s_dadda_pg_rca32_u_pg_rca_or49_y0 = f_s_dadda_pg_rca32_u_pg_rca_or49_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and50_f_s_dadda_pg_rca32_u_pg_rca_fa50_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa50_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and50_y0 = f_s_dadda_pg_rca32_u_pg_rca_and50_f_s_dadda_pg_rca32_u_pg_rca_or49_y0 & f_s_dadda_pg_rca32_u_pg_rca_and50_f_s_dadda_pg_rca32_u_pg_rca_fa50_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or50_f_s_dadda_pg_rca32_u_pg_rca_and50_y0 = f_s_dadda_pg_rca32_u_pg_rca_and50_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or50_f_s_dadda_pg_rca32_u_pg_rca_fa50_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa50_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or50_y0 = f_s_dadda_pg_rca32_u_pg_rca_or50_f_s_dadda_pg_rca32_u_pg_rca_and50_y0 | f_s_dadda_pg_rca32_u_pg_rca_or50_f_s_dadda_pg_rca32_u_pg_rca_fa50_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_fa832_y2 = f_s_dadda_pg_rca32_fa832_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_fa890_y2 = f_s_dadda_pg_rca32_fa890_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_u_pg_rca_or50_y0 = f_s_dadda_pg_rca32_u_pg_rca_or50_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa51_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_fa832_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_fa890_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa51_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_fa832_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_fa890_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa51_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa51_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa51_f_s_dadda_pg_rca32_u_pg_rca_or50_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and51_f_s_dadda_pg_rca32_u_pg_rca_or50_y0 = f_s_dadda_pg_rca32_u_pg_rca_or50_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and51_f_s_dadda_pg_rca32_u_pg_rca_fa51_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa51_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and51_y0 = f_s_dadda_pg_rca32_u_pg_rca_and51_f_s_dadda_pg_rca32_u_pg_rca_or50_y0 & f_s_dadda_pg_rca32_u_pg_rca_and51_f_s_dadda_pg_rca32_u_pg_rca_fa51_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or51_f_s_dadda_pg_rca32_u_pg_rca_and51_y0 = f_s_dadda_pg_rca32_u_pg_rca_and51_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or51_f_s_dadda_pg_rca32_u_pg_rca_fa51_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa51_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or51_y0 = f_s_dadda_pg_rca32_u_pg_rca_or51_f_s_dadda_pg_rca32_u_pg_rca_and51_y0 | f_s_dadda_pg_rca32_u_pg_rca_or51_f_s_dadda_pg_rca32_u_pg_rca_fa51_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_fa833_y2 = f_s_dadda_pg_rca32_fa833_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_fa891_y2 = f_s_dadda_pg_rca32_fa891_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_u_pg_rca_or51_y0 = f_s_dadda_pg_rca32_u_pg_rca_or51_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa52_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_fa833_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_fa891_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa52_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_fa833_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_fa891_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa52_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa52_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa52_f_s_dadda_pg_rca32_u_pg_rca_or51_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and52_f_s_dadda_pg_rca32_u_pg_rca_or51_y0 = f_s_dadda_pg_rca32_u_pg_rca_or51_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and52_f_s_dadda_pg_rca32_u_pg_rca_fa52_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa52_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and52_y0 = f_s_dadda_pg_rca32_u_pg_rca_and52_f_s_dadda_pg_rca32_u_pg_rca_or51_y0 & f_s_dadda_pg_rca32_u_pg_rca_and52_f_s_dadda_pg_rca32_u_pg_rca_fa52_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or52_f_s_dadda_pg_rca32_u_pg_rca_and52_y0 = f_s_dadda_pg_rca32_u_pg_rca_and52_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or52_f_s_dadda_pg_rca32_u_pg_rca_fa52_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa52_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or52_y0 = f_s_dadda_pg_rca32_u_pg_rca_or52_f_s_dadda_pg_rca32_u_pg_rca_and52_y0 | f_s_dadda_pg_rca32_u_pg_rca_or52_f_s_dadda_pg_rca32_u_pg_rca_fa52_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_fa834_y2 = f_s_dadda_pg_rca32_fa834_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_fa892_y2 = f_s_dadda_pg_rca32_fa892_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_u_pg_rca_or52_y0 = f_s_dadda_pg_rca32_u_pg_rca_or52_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa53_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_fa834_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_fa892_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa53_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_fa834_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_fa892_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa53_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa53_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa53_f_s_dadda_pg_rca32_u_pg_rca_or52_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and53_f_s_dadda_pg_rca32_u_pg_rca_or52_y0 = f_s_dadda_pg_rca32_u_pg_rca_or52_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and53_f_s_dadda_pg_rca32_u_pg_rca_fa53_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa53_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and53_y0 = f_s_dadda_pg_rca32_u_pg_rca_and53_f_s_dadda_pg_rca32_u_pg_rca_or52_y0 & f_s_dadda_pg_rca32_u_pg_rca_and53_f_s_dadda_pg_rca32_u_pg_rca_fa53_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or53_f_s_dadda_pg_rca32_u_pg_rca_and53_y0 = f_s_dadda_pg_rca32_u_pg_rca_and53_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or53_f_s_dadda_pg_rca32_u_pg_rca_fa53_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa53_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or53_y0 = f_s_dadda_pg_rca32_u_pg_rca_or53_f_s_dadda_pg_rca32_u_pg_rca_and53_y0 | f_s_dadda_pg_rca32_u_pg_rca_or53_f_s_dadda_pg_rca32_u_pg_rca_fa53_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_fa835_y2 = f_s_dadda_pg_rca32_fa835_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_fa893_y2 = f_s_dadda_pg_rca32_fa893_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_u_pg_rca_or53_y0 = f_s_dadda_pg_rca32_u_pg_rca_or53_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa54_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_fa835_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_fa893_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa54_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_fa835_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_fa893_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa54_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa54_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa54_f_s_dadda_pg_rca32_u_pg_rca_or53_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and54_f_s_dadda_pg_rca32_u_pg_rca_or53_y0 = f_s_dadda_pg_rca32_u_pg_rca_or53_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and54_f_s_dadda_pg_rca32_u_pg_rca_fa54_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa54_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and54_y0 = f_s_dadda_pg_rca32_u_pg_rca_and54_f_s_dadda_pg_rca32_u_pg_rca_or53_y0 & f_s_dadda_pg_rca32_u_pg_rca_and54_f_s_dadda_pg_rca32_u_pg_rca_fa54_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or54_f_s_dadda_pg_rca32_u_pg_rca_and54_y0 = f_s_dadda_pg_rca32_u_pg_rca_and54_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or54_f_s_dadda_pg_rca32_u_pg_rca_fa54_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa54_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or54_y0 = f_s_dadda_pg_rca32_u_pg_rca_or54_f_s_dadda_pg_rca32_u_pg_rca_and54_y0 | f_s_dadda_pg_rca32_u_pg_rca_or54_f_s_dadda_pg_rca32_u_pg_rca_fa54_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_fa836_y2 = f_s_dadda_pg_rca32_fa836_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_fa894_y2 = f_s_dadda_pg_rca32_fa894_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_u_pg_rca_or54_y0 = f_s_dadda_pg_rca32_u_pg_rca_or54_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa55_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_fa836_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_fa894_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa55_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_fa836_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_fa894_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa55_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa55_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa55_f_s_dadda_pg_rca32_u_pg_rca_or54_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and55_f_s_dadda_pg_rca32_u_pg_rca_or54_y0 = f_s_dadda_pg_rca32_u_pg_rca_or54_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and55_f_s_dadda_pg_rca32_u_pg_rca_fa55_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa55_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and55_y0 = f_s_dadda_pg_rca32_u_pg_rca_and55_f_s_dadda_pg_rca32_u_pg_rca_or54_y0 & f_s_dadda_pg_rca32_u_pg_rca_and55_f_s_dadda_pg_rca32_u_pg_rca_fa55_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or55_f_s_dadda_pg_rca32_u_pg_rca_and55_y0 = f_s_dadda_pg_rca32_u_pg_rca_and55_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or55_f_s_dadda_pg_rca32_u_pg_rca_fa55_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa55_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or55_y0 = f_s_dadda_pg_rca32_u_pg_rca_or55_f_s_dadda_pg_rca32_u_pg_rca_and55_y0 | f_s_dadda_pg_rca32_u_pg_rca_or55_f_s_dadda_pg_rca32_u_pg_rca_fa55_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_fa837_y2 = f_s_dadda_pg_rca32_fa837_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_fa895_y2 = f_s_dadda_pg_rca32_fa895_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_u_pg_rca_or55_y0 = f_s_dadda_pg_rca32_u_pg_rca_or55_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa56_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_fa837_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_fa895_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa56_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_fa837_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_fa895_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa56_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa56_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa56_f_s_dadda_pg_rca32_u_pg_rca_or55_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and56_f_s_dadda_pg_rca32_u_pg_rca_or55_y0 = f_s_dadda_pg_rca32_u_pg_rca_or55_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and56_f_s_dadda_pg_rca32_u_pg_rca_fa56_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa56_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and56_y0 = f_s_dadda_pg_rca32_u_pg_rca_and56_f_s_dadda_pg_rca32_u_pg_rca_or55_y0 & f_s_dadda_pg_rca32_u_pg_rca_and56_f_s_dadda_pg_rca32_u_pg_rca_fa56_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or56_f_s_dadda_pg_rca32_u_pg_rca_and56_y0 = f_s_dadda_pg_rca32_u_pg_rca_and56_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or56_f_s_dadda_pg_rca32_u_pg_rca_fa56_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa56_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or56_y0 = f_s_dadda_pg_rca32_u_pg_rca_or56_f_s_dadda_pg_rca32_u_pg_rca_and56_y0 | f_s_dadda_pg_rca32_u_pg_rca_or56_f_s_dadda_pg_rca32_u_pg_rca_fa56_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_fa838_y2 = f_s_dadda_pg_rca32_fa838_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_fa896_y2 = f_s_dadda_pg_rca32_fa896_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_u_pg_rca_or56_y0 = f_s_dadda_pg_rca32_u_pg_rca_or56_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa57_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_fa838_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_fa896_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa57_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_fa838_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_fa896_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa57_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa57_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa57_f_s_dadda_pg_rca32_u_pg_rca_or56_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and57_f_s_dadda_pg_rca32_u_pg_rca_or56_y0 = f_s_dadda_pg_rca32_u_pg_rca_or56_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and57_f_s_dadda_pg_rca32_u_pg_rca_fa57_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa57_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and57_y0 = f_s_dadda_pg_rca32_u_pg_rca_and57_f_s_dadda_pg_rca32_u_pg_rca_or56_y0 & f_s_dadda_pg_rca32_u_pg_rca_and57_f_s_dadda_pg_rca32_u_pg_rca_fa57_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or57_f_s_dadda_pg_rca32_u_pg_rca_and57_y0 = f_s_dadda_pg_rca32_u_pg_rca_and57_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or57_f_s_dadda_pg_rca32_u_pg_rca_fa57_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa57_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or57_y0 = f_s_dadda_pg_rca32_u_pg_rca_or57_f_s_dadda_pg_rca32_u_pg_rca_and57_y0 | f_s_dadda_pg_rca32_u_pg_rca_or57_f_s_dadda_pg_rca32_u_pg_rca_fa57_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_fa839_y2 = f_s_dadda_pg_rca32_fa839_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_fa897_y2 = f_s_dadda_pg_rca32_fa897_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_u_pg_rca_or57_y0 = f_s_dadda_pg_rca32_u_pg_rca_or57_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa58_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_fa839_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_fa897_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa58_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_fa839_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_fa897_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa58_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa58_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa58_f_s_dadda_pg_rca32_u_pg_rca_or57_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and58_f_s_dadda_pg_rca32_u_pg_rca_or57_y0 = f_s_dadda_pg_rca32_u_pg_rca_or57_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and58_f_s_dadda_pg_rca32_u_pg_rca_fa58_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa58_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and58_y0 = f_s_dadda_pg_rca32_u_pg_rca_and58_f_s_dadda_pg_rca32_u_pg_rca_or57_y0 & f_s_dadda_pg_rca32_u_pg_rca_and58_f_s_dadda_pg_rca32_u_pg_rca_fa58_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or58_f_s_dadda_pg_rca32_u_pg_rca_and58_y0 = f_s_dadda_pg_rca32_u_pg_rca_and58_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or58_f_s_dadda_pg_rca32_u_pg_rca_fa58_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa58_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or58_y0 = f_s_dadda_pg_rca32_u_pg_rca_or58_f_s_dadda_pg_rca32_u_pg_rca_and58_y0 | f_s_dadda_pg_rca32_u_pg_rca_or58_f_s_dadda_pg_rca32_u_pg_rca_fa58_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_fa840_y2 = f_s_dadda_pg_rca32_fa840_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_fa898_y2 = f_s_dadda_pg_rca32_fa898_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_u_pg_rca_or58_y0 = f_s_dadda_pg_rca32_u_pg_rca_or58_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa59_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_fa840_y2 ^ f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_fa898_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa59_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_fa840_y2 & f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_fa898_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa59_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa59_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa59_f_s_dadda_pg_rca32_u_pg_rca_or58_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and59_f_s_dadda_pg_rca32_u_pg_rca_or58_y0 = f_s_dadda_pg_rca32_u_pg_rca_or58_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and59_f_s_dadda_pg_rca32_u_pg_rca_fa59_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa59_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and59_y0 = f_s_dadda_pg_rca32_u_pg_rca_and59_f_s_dadda_pg_rca32_u_pg_rca_or58_y0 & f_s_dadda_pg_rca32_u_pg_rca_and59_f_s_dadda_pg_rca32_u_pg_rca_fa59_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or59_f_s_dadda_pg_rca32_u_pg_rca_and59_y0 = f_s_dadda_pg_rca32_u_pg_rca_and59_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or59_f_s_dadda_pg_rca32_u_pg_rca_fa59_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa59_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or59_y0 = f_s_dadda_pg_rca32_u_pg_rca_or59_f_s_dadda_pg_rca32_u_pg_rca_and59_y0 | f_s_dadda_pg_rca32_u_pg_rca_or59_f_s_dadda_pg_rca32_u_pg_rca_fa59_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_nand_30_31_y0 = f_s_dadda_pg_rca32_nand_30_31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_fa899_y2 = f_s_dadda_pg_rca32_fa899_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_u_pg_rca_or59_y0 = f_s_dadda_pg_rca32_u_pg_rca_or59_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa60_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_nand_30_31_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_fa899_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa60_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_nand_30_31_y0 & f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_fa899_y2;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa60_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa60_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa60_f_s_dadda_pg_rca32_u_pg_rca_or59_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and60_f_s_dadda_pg_rca32_u_pg_rca_or59_y0 = f_s_dadda_pg_rca32_u_pg_rca_or59_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and60_f_s_dadda_pg_rca32_u_pg_rca_fa60_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa60_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and60_y0 = f_s_dadda_pg_rca32_u_pg_rca_and60_f_s_dadda_pg_rca32_u_pg_rca_or59_y0 & f_s_dadda_pg_rca32_u_pg_rca_and60_f_s_dadda_pg_rca32_u_pg_rca_fa60_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or60_f_s_dadda_pg_rca32_u_pg_rca_and60_y0 = f_s_dadda_pg_rca32_u_pg_rca_and60_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or60_f_s_dadda_pg_rca32_u_pg_rca_fa60_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa60_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or60_y0 = f_s_dadda_pg_rca32_u_pg_rca_or60_f_s_dadda_pg_rca32_u_pg_rca_and60_y0 | f_s_dadda_pg_rca32_u_pg_rca_or60_f_s_dadda_pg_rca32_u_pg_rca_fa60_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_fa899_y4 = f_s_dadda_pg_rca32_fa899_y4;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_and_31_31_y0 = f_s_dadda_pg_rca32_and_31_31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_u_pg_rca_or60_y0 = f_s_dadda_pg_rca32_u_pg_rca_or60_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa61_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_fa899_y4 ^ f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_and_31_31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa61_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_fa899_y4 & f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_and_31_31_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_fa61_y2 = f_s_dadda_pg_rca32_u_pg_rca_fa61_y0 ^ f_s_dadda_pg_rca32_u_pg_rca_fa61_f_s_dadda_pg_rca32_u_pg_rca_or60_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and61_f_s_dadda_pg_rca32_u_pg_rca_or60_y0 = f_s_dadda_pg_rca32_u_pg_rca_or60_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and61_f_s_dadda_pg_rca32_u_pg_rca_fa61_y0 = f_s_dadda_pg_rca32_u_pg_rca_fa61_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_and61_y0 = f_s_dadda_pg_rca32_u_pg_rca_and61_f_s_dadda_pg_rca32_u_pg_rca_or60_y0 & f_s_dadda_pg_rca32_u_pg_rca_and61_f_s_dadda_pg_rca32_u_pg_rca_fa61_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or61_f_s_dadda_pg_rca32_u_pg_rca_and61_y0 = f_s_dadda_pg_rca32_u_pg_rca_and61_y0;
  assign f_s_dadda_pg_rca32_u_pg_rca_or61_f_s_dadda_pg_rca32_u_pg_rca_fa61_y1 = f_s_dadda_pg_rca32_u_pg_rca_fa61_y1;
  assign f_s_dadda_pg_rca32_u_pg_rca_or61_y0 = f_s_dadda_pg_rca32_u_pg_rca_or61_f_s_dadda_pg_rca32_u_pg_rca_and61_y0 | f_s_dadda_pg_rca32_u_pg_rca_or61_f_s_dadda_pg_rca32_u_pg_rca_fa61_y1;
  assign f_s_dadda_pg_rca32_xor0_constant_wire_1 = constant_wire_1;
  assign f_s_dadda_pg_rca32_xor0_f_s_dadda_pg_rca32_u_pg_rca_or61_y0 = f_s_dadda_pg_rca32_u_pg_rca_or61_y0;
  assign f_s_dadda_pg_rca32_xor0_y0 = f_s_dadda_pg_rca32_xor0_constant_wire_1 ^ f_s_dadda_pg_rca32_xor0_f_s_dadda_pg_rca32_u_pg_rca_or61_y0;

  assign out[0] = f_s_dadda_pg_rca32_and_0_0_y0;
  assign out[1] = f_s_dadda_pg_rca32_u_pg_rca_fa0_y2;
  assign out[2] = f_s_dadda_pg_rca32_u_pg_rca_fa1_y2;
  assign out[3] = f_s_dadda_pg_rca32_u_pg_rca_fa2_y2;
  assign out[4] = f_s_dadda_pg_rca32_u_pg_rca_fa3_y2;
  assign out[5] = f_s_dadda_pg_rca32_u_pg_rca_fa4_y2;
  assign out[6] = f_s_dadda_pg_rca32_u_pg_rca_fa5_y2;
  assign out[7] = f_s_dadda_pg_rca32_u_pg_rca_fa6_y2;
  assign out[8] = f_s_dadda_pg_rca32_u_pg_rca_fa7_y2;
  assign out[9] = f_s_dadda_pg_rca32_u_pg_rca_fa8_y2;
  assign out[10] = f_s_dadda_pg_rca32_u_pg_rca_fa9_y2;
  assign out[11] = f_s_dadda_pg_rca32_u_pg_rca_fa10_y2;
  assign out[12] = f_s_dadda_pg_rca32_u_pg_rca_fa11_y2;
  assign out[13] = f_s_dadda_pg_rca32_u_pg_rca_fa12_y2;
  assign out[14] = f_s_dadda_pg_rca32_u_pg_rca_fa13_y2;
  assign out[15] = f_s_dadda_pg_rca32_u_pg_rca_fa14_y2;
  assign out[16] = f_s_dadda_pg_rca32_u_pg_rca_fa15_y2;
  assign out[17] = f_s_dadda_pg_rca32_u_pg_rca_fa16_y2;
  assign out[18] = f_s_dadda_pg_rca32_u_pg_rca_fa17_y2;
  assign out[19] = f_s_dadda_pg_rca32_u_pg_rca_fa18_y2;
  assign out[20] = f_s_dadda_pg_rca32_u_pg_rca_fa19_y2;
  assign out[21] = f_s_dadda_pg_rca32_u_pg_rca_fa20_y2;
  assign out[22] = f_s_dadda_pg_rca32_u_pg_rca_fa21_y2;
  assign out[23] = f_s_dadda_pg_rca32_u_pg_rca_fa22_y2;
  assign out[24] = f_s_dadda_pg_rca32_u_pg_rca_fa23_y2;
  assign out[25] = f_s_dadda_pg_rca32_u_pg_rca_fa24_y2;
  assign out[26] = f_s_dadda_pg_rca32_u_pg_rca_fa25_y2;
  assign out[27] = f_s_dadda_pg_rca32_u_pg_rca_fa26_y2;
  assign out[28] = f_s_dadda_pg_rca32_u_pg_rca_fa27_y2;
  assign out[29] = f_s_dadda_pg_rca32_u_pg_rca_fa28_y2;
  assign out[30] = f_s_dadda_pg_rca32_u_pg_rca_fa29_y2;
  assign out[31] = f_s_dadda_pg_rca32_u_pg_rca_fa30_y2;
  assign out[32] = f_s_dadda_pg_rca32_u_pg_rca_fa31_y2;
  assign out[33] = f_s_dadda_pg_rca32_u_pg_rca_fa32_y2;
  assign out[34] = f_s_dadda_pg_rca32_u_pg_rca_fa33_y2;
  assign out[35] = f_s_dadda_pg_rca32_u_pg_rca_fa34_y2;
  assign out[36] = f_s_dadda_pg_rca32_u_pg_rca_fa35_y2;
  assign out[37] = f_s_dadda_pg_rca32_u_pg_rca_fa36_y2;
  assign out[38] = f_s_dadda_pg_rca32_u_pg_rca_fa37_y2;
  assign out[39] = f_s_dadda_pg_rca32_u_pg_rca_fa38_y2;
  assign out[40] = f_s_dadda_pg_rca32_u_pg_rca_fa39_y2;
  assign out[41] = f_s_dadda_pg_rca32_u_pg_rca_fa40_y2;
  assign out[42] = f_s_dadda_pg_rca32_u_pg_rca_fa41_y2;
  assign out[43] = f_s_dadda_pg_rca32_u_pg_rca_fa42_y2;
  assign out[44] = f_s_dadda_pg_rca32_u_pg_rca_fa43_y2;
  assign out[45] = f_s_dadda_pg_rca32_u_pg_rca_fa44_y2;
  assign out[46] = f_s_dadda_pg_rca32_u_pg_rca_fa45_y2;
  assign out[47] = f_s_dadda_pg_rca32_u_pg_rca_fa46_y2;
  assign out[48] = f_s_dadda_pg_rca32_u_pg_rca_fa47_y2;
  assign out[49] = f_s_dadda_pg_rca32_u_pg_rca_fa48_y2;
  assign out[50] = f_s_dadda_pg_rca32_u_pg_rca_fa49_y2;
  assign out[51] = f_s_dadda_pg_rca32_u_pg_rca_fa50_y2;
  assign out[52] = f_s_dadda_pg_rca32_u_pg_rca_fa51_y2;
  assign out[53] = f_s_dadda_pg_rca32_u_pg_rca_fa52_y2;
  assign out[54] = f_s_dadda_pg_rca32_u_pg_rca_fa53_y2;
  assign out[55] = f_s_dadda_pg_rca32_u_pg_rca_fa54_y2;
  assign out[56] = f_s_dadda_pg_rca32_u_pg_rca_fa55_y2;
  assign out[57] = f_s_dadda_pg_rca32_u_pg_rca_fa56_y2;
  assign out[58] = f_s_dadda_pg_rca32_u_pg_rca_fa57_y2;
  assign out[59] = f_s_dadda_pg_rca32_u_pg_rca_fa58_y2;
  assign out[60] = f_s_dadda_pg_rca32_u_pg_rca_fa59_y2;
  assign out[61] = f_s_dadda_pg_rca32_u_pg_rca_fa60_y2;
  assign out[62] = f_s_dadda_pg_rca32_u_pg_rca_fa61_y2;
  assign out[63] = f_s_dadda_pg_rca32_xor0_y0;
endmodule