module f_s_pg_rca24(input [23:0] a, input [23:0] b, output [24:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire constant_wire_value_0_a_0;
  wire constant_wire_value_0_b_0;
  wire constant_wire_value_0_y0;
  wire constant_wire_value_0_y1;
  wire constant_wire_0;
  wire f_s_pg_rca24_fa0_a_0;
  wire f_s_pg_rca24_fa0_b_0;
  wire f_s_pg_rca24_fa0_y0;
  wire f_s_pg_rca24_fa0_y1;
  wire f_s_pg_rca24_fa0_constant_wire_0;
  wire f_s_pg_rca24_fa0_y2;
  wire f_s_pg_rca24_and0_constant_wire_0;
  wire f_s_pg_rca24_and0_f_s_pg_rca24_fa0_y0;
  wire f_s_pg_rca24_and0_y0;
  wire f_s_pg_rca24_or0_f_s_pg_rca24_and0_y0;
  wire f_s_pg_rca24_or0_f_s_pg_rca24_fa0_y1;
  wire f_s_pg_rca24_or0_y0;
  wire f_s_pg_rca24_fa1_a_1;
  wire f_s_pg_rca24_fa1_b_1;
  wire f_s_pg_rca24_fa1_y0;
  wire f_s_pg_rca24_fa1_y1;
  wire f_s_pg_rca24_fa1_f_s_pg_rca24_or0_y0;
  wire f_s_pg_rca24_fa1_y2;
  wire f_s_pg_rca24_and1_f_s_pg_rca24_or0_y0;
  wire f_s_pg_rca24_and1_f_s_pg_rca24_fa1_y0;
  wire f_s_pg_rca24_and1_y0;
  wire f_s_pg_rca24_or1_f_s_pg_rca24_and1_y0;
  wire f_s_pg_rca24_or1_f_s_pg_rca24_fa1_y1;
  wire f_s_pg_rca24_or1_y0;
  wire f_s_pg_rca24_fa2_a_2;
  wire f_s_pg_rca24_fa2_b_2;
  wire f_s_pg_rca24_fa2_y0;
  wire f_s_pg_rca24_fa2_y1;
  wire f_s_pg_rca24_fa2_f_s_pg_rca24_or1_y0;
  wire f_s_pg_rca24_fa2_y2;
  wire f_s_pg_rca24_and2_f_s_pg_rca24_or1_y0;
  wire f_s_pg_rca24_and2_f_s_pg_rca24_fa2_y0;
  wire f_s_pg_rca24_and2_y0;
  wire f_s_pg_rca24_or2_f_s_pg_rca24_and2_y0;
  wire f_s_pg_rca24_or2_f_s_pg_rca24_fa2_y1;
  wire f_s_pg_rca24_or2_y0;
  wire f_s_pg_rca24_fa3_a_3;
  wire f_s_pg_rca24_fa3_b_3;
  wire f_s_pg_rca24_fa3_y0;
  wire f_s_pg_rca24_fa3_y1;
  wire f_s_pg_rca24_fa3_f_s_pg_rca24_or2_y0;
  wire f_s_pg_rca24_fa3_y2;
  wire f_s_pg_rca24_and3_f_s_pg_rca24_or2_y0;
  wire f_s_pg_rca24_and3_f_s_pg_rca24_fa3_y0;
  wire f_s_pg_rca24_and3_y0;
  wire f_s_pg_rca24_or3_f_s_pg_rca24_and3_y0;
  wire f_s_pg_rca24_or3_f_s_pg_rca24_fa3_y1;
  wire f_s_pg_rca24_or3_y0;
  wire f_s_pg_rca24_fa4_a_4;
  wire f_s_pg_rca24_fa4_b_4;
  wire f_s_pg_rca24_fa4_y0;
  wire f_s_pg_rca24_fa4_y1;
  wire f_s_pg_rca24_fa4_f_s_pg_rca24_or3_y0;
  wire f_s_pg_rca24_fa4_y2;
  wire f_s_pg_rca24_and4_f_s_pg_rca24_or3_y0;
  wire f_s_pg_rca24_and4_f_s_pg_rca24_fa4_y0;
  wire f_s_pg_rca24_and4_y0;
  wire f_s_pg_rca24_or4_f_s_pg_rca24_and4_y0;
  wire f_s_pg_rca24_or4_f_s_pg_rca24_fa4_y1;
  wire f_s_pg_rca24_or4_y0;
  wire f_s_pg_rca24_fa5_a_5;
  wire f_s_pg_rca24_fa5_b_5;
  wire f_s_pg_rca24_fa5_y0;
  wire f_s_pg_rca24_fa5_y1;
  wire f_s_pg_rca24_fa5_f_s_pg_rca24_or4_y0;
  wire f_s_pg_rca24_fa5_y2;
  wire f_s_pg_rca24_and5_f_s_pg_rca24_or4_y0;
  wire f_s_pg_rca24_and5_f_s_pg_rca24_fa5_y0;
  wire f_s_pg_rca24_and5_y0;
  wire f_s_pg_rca24_or5_f_s_pg_rca24_and5_y0;
  wire f_s_pg_rca24_or5_f_s_pg_rca24_fa5_y1;
  wire f_s_pg_rca24_or5_y0;
  wire f_s_pg_rca24_fa6_a_6;
  wire f_s_pg_rca24_fa6_b_6;
  wire f_s_pg_rca24_fa6_y0;
  wire f_s_pg_rca24_fa6_y1;
  wire f_s_pg_rca24_fa6_f_s_pg_rca24_or5_y0;
  wire f_s_pg_rca24_fa6_y2;
  wire f_s_pg_rca24_and6_f_s_pg_rca24_or5_y0;
  wire f_s_pg_rca24_and6_f_s_pg_rca24_fa6_y0;
  wire f_s_pg_rca24_and6_y0;
  wire f_s_pg_rca24_or6_f_s_pg_rca24_and6_y0;
  wire f_s_pg_rca24_or6_f_s_pg_rca24_fa6_y1;
  wire f_s_pg_rca24_or6_y0;
  wire f_s_pg_rca24_fa7_a_7;
  wire f_s_pg_rca24_fa7_b_7;
  wire f_s_pg_rca24_fa7_y0;
  wire f_s_pg_rca24_fa7_y1;
  wire f_s_pg_rca24_fa7_f_s_pg_rca24_or6_y0;
  wire f_s_pg_rca24_fa7_y2;
  wire f_s_pg_rca24_and7_f_s_pg_rca24_or6_y0;
  wire f_s_pg_rca24_and7_f_s_pg_rca24_fa7_y0;
  wire f_s_pg_rca24_and7_y0;
  wire f_s_pg_rca24_or7_f_s_pg_rca24_and7_y0;
  wire f_s_pg_rca24_or7_f_s_pg_rca24_fa7_y1;
  wire f_s_pg_rca24_or7_y0;
  wire f_s_pg_rca24_fa8_a_8;
  wire f_s_pg_rca24_fa8_b_8;
  wire f_s_pg_rca24_fa8_y0;
  wire f_s_pg_rca24_fa8_y1;
  wire f_s_pg_rca24_fa8_f_s_pg_rca24_or7_y0;
  wire f_s_pg_rca24_fa8_y2;
  wire f_s_pg_rca24_and8_f_s_pg_rca24_or7_y0;
  wire f_s_pg_rca24_and8_f_s_pg_rca24_fa8_y0;
  wire f_s_pg_rca24_and8_y0;
  wire f_s_pg_rca24_or8_f_s_pg_rca24_and8_y0;
  wire f_s_pg_rca24_or8_f_s_pg_rca24_fa8_y1;
  wire f_s_pg_rca24_or8_y0;
  wire f_s_pg_rca24_fa9_a_9;
  wire f_s_pg_rca24_fa9_b_9;
  wire f_s_pg_rca24_fa9_y0;
  wire f_s_pg_rca24_fa9_y1;
  wire f_s_pg_rca24_fa9_f_s_pg_rca24_or8_y0;
  wire f_s_pg_rca24_fa9_y2;
  wire f_s_pg_rca24_and9_f_s_pg_rca24_or8_y0;
  wire f_s_pg_rca24_and9_f_s_pg_rca24_fa9_y0;
  wire f_s_pg_rca24_and9_y0;
  wire f_s_pg_rca24_or9_f_s_pg_rca24_and9_y0;
  wire f_s_pg_rca24_or9_f_s_pg_rca24_fa9_y1;
  wire f_s_pg_rca24_or9_y0;
  wire f_s_pg_rca24_fa10_a_10;
  wire f_s_pg_rca24_fa10_b_10;
  wire f_s_pg_rca24_fa10_y0;
  wire f_s_pg_rca24_fa10_y1;
  wire f_s_pg_rca24_fa10_f_s_pg_rca24_or9_y0;
  wire f_s_pg_rca24_fa10_y2;
  wire f_s_pg_rca24_and10_f_s_pg_rca24_or9_y0;
  wire f_s_pg_rca24_and10_f_s_pg_rca24_fa10_y0;
  wire f_s_pg_rca24_and10_y0;
  wire f_s_pg_rca24_or10_f_s_pg_rca24_and10_y0;
  wire f_s_pg_rca24_or10_f_s_pg_rca24_fa10_y1;
  wire f_s_pg_rca24_or10_y0;
  wire f_s_pg_rca24_fa11_a_11;
  wire f_s_pg_rca24_fa11_b_11;
  wire f_s_pg_rca24_fa11_y0;
  wire f_s_pg_rca24_fa11_y1;
  wire f_s_pg_rca24_fa11_f_s_pg_rca24_or10_y0;
  wire f_s_pg_rca24_fa11_y2;
  wire f_s_pg_rca24_and11_f_s_pg_rca24_or10_y0;
  wire f_s_pg_rca24_and11_f_s_pg_rca24_fa11_y0;
  wire f_s_pg_rca24_and11_y0;
  wire f_s_pg_rca24_or11_f_s_pg_rca24_and11_y0;
  wire f_s_pg_rca24_or11_f_s_pg_rca24_fa11_y1;
  wire f_s_pg_rca24_or11_y0;
  wire f_s_pg_rca24_fa12_a_12;
  wire f_s_pg_rca24_fa12_b_12;
  wire f_s_pg_rca24_fa12_y0;
  wire f_s_pg_rca24_fa12_y1;
  wire f_s_pg_rca24_fa12_f_s_pg_rca24_or11_y0;
  wire f_s_pg_rca24_fa12_y2;
  wire f_s_pg_rca24_and12_f_s_pg_rca24_or11_y0;
  wire f_s_pg_rca24_and12_f_s_pg_rca24_fa12_y0;
  wire f_s_pg_rca24_and12_y0;
  wire f_s_pg_rca24_or12_f_s_pg_rca24_and12_y0;
  wire f_s_pg_rca24_or12_f_s_pg_rca24_fa12_y1;
  wire f_s_pg_rca24_or12_y0;
  wire f_s_pg_rca24_fa13_a_13;
  wire f_s_pg_rca24_fa13_b_13;
  wire f_s_pg_rca24_fa13_y0;
  wire f_s_pg_rca24_fa13_y1;
  wire f_s_pg_rca24_fa13_f_s_pg_rca24_or12_y0;
  wire f_s_pg_rca24_fa13_y2;
  wire f_s_pg_rca24_and13_f_s_pg_rca24_or12_y0;
  wire f_s_pg_rca24_and13_f_s_pg_rca24_fa13_y0;
  wire f_s_pg_rca24_and13_y0;
  wire f_s_pg_rca24_or13_f_s_pg_rca24_and13_y0;
  wire f_s_pg_rca24_or13_f_s_pg_rca24_fa13_y1;
  wire f_s_pg_rca24_or13_y0;
  wire f_s_pg_rca24_fa14_a_14;
  wire f_s_pg_rca24_fa14_b_14;
  wire f_s_pg_rca24_fa14_y0;
  wire f_s_pg_rca24_fa14_y1;
  wire f_s_pg_rca24_fa14_f_s_pg_rca24_or13_y0;
  wire f_s_pg_rca24_fa14_y2;
  wire f_s_pg_rca24_and14_f_s_pg_rca24_or13_y0;
  wire f_s_pg_rca24_and14_f_s_pg_rca24_fa14_y0;
  wire f_s_pg_rca24_and14_y0;
  wire f_s_pg_rca24_or14_f_s_pg_rca24_and14_y0;
  wire f_s_pg_rca24_or14_f_s_pg_rca24_fa14_y1;
  wire f_s_pg_rca24_or14_y0;
  wire f_s_pg_rca24_fa15_a_15;
  wire f_s_pg_rca24_fa15_b_15;
  wire f_s_pg_rca24_fa15_y0;
  wire f_s_pg_rca24_fa15_y1;
  wire f_s_pg_rca24_fa15_f_s_pg_rca24_or14_y0;
  wire f_s_pg_rca24_fa15_y2;
  wire f_s_pg_rca24_and15_f_s_pg_rca24_or14_y0;
  wire f_s_pg_rca24_and15_f_s_pg_rca24_fa15_y0;
  wire f_s_pg_rca24_and15_y0;
  wire f_s_pg_rca24_or15_f_s_pg_rca24_and15_y0;
  wire f_s_pg_rca24_or15_f_s_pg_rca24_fa15_y1;
  wire f_s_pg_rca24_or15_y0;
  wire f_s_pg_rca24_fa16_a_16;
  wire f_s_pg_rca24_fa16_b_16;
  wire f_s_pg_rca24_fa16_y0;
  wire f_s_pg_rca24_fa16_y1;
  wire f_s_pg_rca24_fa16_f_s_pg_rca24_or15_y0;
  wire f_s_pg_rca24_fa16_y2;
  wire f_s_pg_rca24_and16_f_s_pg_rca24_or15_y0;
  wire f_s_pg_rca24_and16_f_s_pg_rca24_fa16_y0;
  wire f_s_pg_rca24_and16_y0;
  wire f_s_pg_rca24_or16_f_s_pg_rca24_and16_y0;
  wire f_s_pg_rca24_or16_f_s_pg_rca24_fa16_y1;
  wire f_s_pg_rca24_or16_y0;
  wire f_s_pg_rca24_fa17_a_17;
  wire f_s_pg_rca24_fa17_b_17;
  wire f_s_pg_rca24_fa17_y0;
  wire f_s_pg_rca24_fa17_y1;
  wire f_s_pg_rca24_fa17_f_s_pg_rca24_or16_y0;
  wire f_s_pg_rca24_fa17_y2;
  wire f_s_pg_rca24_and17_f_s_pg_rca24_or16_y0;
  wire f_s_pg_rca24_and17_f_s_pg_rca24_fa17_y0;
  wire f_s_pg_rca24_and17_y0;
  wire f_s_pg_rca24_or17_f_s_pg_rca24_and17_y0;
  wire f_s_pg_rca24_or17_f_s_pg_rca24_fa17_y1;
  wire f_s_pg_rca24_or17_y0;
  wire f_s_pg_rca24_fa18_a_18;
  wire f_s_pg_rca24_fa18_b_18;
  wire f_s_pg_rca24_fa18_y0;
  wire f_s_pg_rca24_fa18_y1;
  wire f_s_pg_rca24_fa18_f_s_pg_rca24_or17_y0;
  wire f_s_pg_rca24_fa18_y2;
  wire f_s_pg_rca24_and18_f_s_pg_rca24_or17_y0;
  wire f_s_pg_rca24_and18_f_s_pg_rca24_fa18_y0;
  wire f_s_pg_rca24_and18_y0;
  wire f_s_pg_rca24_or18_f_s_pg_rca24_and18_y0;
  wire f_s_pg_rca24_or18_f_s_pg_rca24_fa18_y1;
  wire f_s_pg_rca24_or18_y0;
  wire f_s_pg_rca24_fa19_a_19;
  wire f_s_pg_rca24_fa19_b_19;
  wire f_s_pg_rca24_fa19_y0;
  wire f_s_pg_rca24_fa19_y1;
  wire f_s_pg_rca24_fa19_f_s_pg_rca24_or18_y0;
  wire f_s_pg_rca24_fa19_y2;
  wire f_s_pg_rca24_and19_f_s_pg_rca24_or18_y0;
  wire f_s_pg_rca24_and19_f_s_pg_rca24_fa19_y0;
  wire f_s_pg_rca24_and19_y0;
  wire f_s_pg_rca24_or19_f_s_pg_rca24_and19_y0;
  wire f_s_pg_rca24_or19_f_s_pg_rca24_fa19_y1;
  wire f_s_pg_rca24_or19_y0;
  wire f_s_pg_rca24_fa20_a_20;
  wire f_s_pg_rca24_fa20_b_20;
  wire f_s_pg_rca24_fa20_y0;
  wire f_s_pg_rca24_fa20_y1;
  wire f_s_pg_rca24_fa20_f_s_pg_rca24_or19_y0;
  wire f_s_pg_rca24_fa20_y2;
  wire f_s_pg_rca24_and20_f_s_pg_rca24_or19_y0;
  wire f_s_pg_rca24_and20_f_s_pg_rca24_fa20_y0;
  wire f_s_pg_rca24_and20_y0;
  wire f_s_pg_rca24_or20_f_s_pg_rca24_and20_y0;
  wire f_s_pg_rca24_or20_f_s_pg_rca24_fa20_y1;
  wire f_s_pg_rca24_or20_y0;
  wire f_s_pg_rca24_fa21_a_21;
  wire f_s_pg_rca24_fa21_b_21;
  wire f_s_pg_rca24_fa21_y0;
  wire f_s_pg_rca24_fa21_y1;
  wire f_s_pg_rca24_fa21_f_s_pg_rca24_or20_y0;
  wire f_s_pg_rca24_fa21_y2;
  wire f_s_pg_rca24_and21_f_s_pg_rca24_or20_y0;
  wire f_s_pg_rca24_and21_f_s_pg_rca24_fa21_y0;
  wire f_s_pg_rca24_and21_y0;
  wire f_s_pg_rca24_or21_f_s_pg_rca24_and21_y0;
  wire f_s_pg_rca24_or21_f_s_pg_rca24_fa21_y1;
  wire f_s_pg_rca24_or21_y0;
  wire f_s_pg_rca24_fa22_a_22;
  wire f_s_pg_rca24_fa22_b_22;
  wire f_s_pg_rca24_fa22_y0;
  wire f_s_pg_rca24_fa22_y1;
  wire f_s_pg_rca24_fa22_f_s_pg_rca24_or21_y0;
  wire f_s_pg_rca24_fa22_y2;
  wire f_s_pg_rca24_and22_f_s_pg_rca24_or21_y0;
  wire f_s_pg_rca24_and22_f_s_pg_rca24_fa22_y0;
  wire f_s_pg_rca24_and22_y0;
  wire f_s_pg_rca24_or22_f_s_pg_rca24_and22_y0;
  wire f_s_pg_rca24_or22_f_s_pg_rca24_fa22_y1;
  wire f_s_pg_rca24_or22_y0;
  wire f_s_pg_rca24_fa23_a_23;
  wire f_s_pg_rca24_fa23_b_23;
  wire f_s_pg_rca24_fa23_y0;
  wire f_s_pg_rca24_fa23_y1;
  wire f_s_pg_rca24_fa23_f_s_pg_rca24_or22_y0;
  wire f_s_pg_rca24_fa23_y2;
  wire f_s_pg_rca24_and23_f_s_pg_rca24_or22_y0;
  wire f_s_pg_rca24_and23_f_s_pg_rca24_fa23_y0;
  wire f_s_pg_rca24_and23_y0;
  wire f_s_pg_rca24_or23_f_s_pg_rca24_and23_y0;
  wire f_s_pg_rca24_or23_f_s_pg_rca24_fa23_y1;
  wire f_s_pg_rca24_or23_y0;
  wire f_s_pg_rca24_xor0_a_23;
  wire f_s_pg_rca24_xor0_b_23;
  wire f_s_pg_rca24_xor0_y0;
  wire f_s_pg_rca24_xor1_f_s_pg_rca24_xor0_y0;
  wire f_s_pg_rca24_xor1_f_s_pg_rca24_or23_y0;
  wire f_s_pg_rca24_xor1_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign constant_wire_value_0_a_0 = a_0;
  assign constant_wire_value_0_b_0 = b_0;
  assign constant_wire_value_0_y0 = constant_wire_value_0_a_0 ^ constant_wire_value_0_b_0;
  assign constant_wire_value_0_y1 = ~(constant_wire_value_0_a_0 ^ constant_wire_value_0_b_0);
  assign constant_wire_0 = ~(constant_wire_value_0_y0 | constant_wire_value_0_y1);
  assign f_s_pg_rca24_fa0_a_0 = a_0;
  assign f_s_pg_rca24_fa0_b_0 = b_0;
  assign f_s_pg_rca24_fa0_constant_wire_0 = constant_wire_0;
  assign f_s_pg_rca24_fa0_y0 = f_s_pg_rca24_fa0_a_0 ^ f_s_pg_rca24_fa0_b_0;
  assign f_s_pg_rca24_fa0_y1 = f_s_pg_rca24_fa0_a_0 & f_s_pg_rca24_fa0_b_0;
  assign f_s_pg_rca24_fa0_y2 = f_s_pg_rca24_fa0_y0 ^ f_s_pg_rca24_fa0_constant_wire_0;
  assign f_s_pg_rca24_and0_constant_wire_0 = constant_wire_0;
  assign f_s_pg_rca24_and0_f_s_pg_rca24_fa0_y0 = f_s_pg_rca24_fa0_y0;
  assign f_s_pg_rca24_and0_y0 = f_s_pg_rca24_and0_constant_wire_0 & f_s_pg_rca24_and0_f_s_pg_rca24_fa0_y0;
  assign f_s_pg_rca24_or0_f_s_pg_rca24_and0_y0 = f_s_pg_rca24_and0_y0;
  assign f_s_pg_rca24_or0_f_s_pg_rca24_fa0_y1 = f_s_pg_rca24_fa0_y1;
  assign f_s_pg_rca24_or0_y0 = f_s_pg_rca24_or0_f_s_pg_rca24_and0_y0 | f_s_pg_rca24_or0_f_s_pg_rca24_fa0_y1;
  assign f_s_pg_rca24_fa1_a_1 = a_1;
  assign f_s_pg_rca24_fa1_b_1 = b_1;
  assign f_s_pg_rca24_fa1_f_s_pg_rca24_or0_y0 = f_s_pg_rca24_or0_y0;
  assign f_s_pg_rca24_fa1_y0 = f_s_pg_rca24_fa1_a_1 ^ f_s_pg_rca24_fa1_b_1;
  assign f_s_pg_rca24_fa1_y1 = f_s_pg_rca24_fa1_a_1 & f_s_pg_rca24_fa1_b_1;
  assign f_s_pg_rca24_fa1_y2 = f_s_pg_rca24_fa1_y0 ^ f_s_pg_rca24_fa1_f_s_pg_rca24_or0_y0;
  assign f_s_pg_rca24_and1_f_s_pg_rca24_or0_y0 = f_s_pg_rca24_or0_y0;
  assign f_s_pg_rca24_and1_f_s_pg_rca24_fa1_y0 = f_s_pg_rca24_fa1_y0;
  assign f_s_pg_rca24_and1_y0 = f_s_pg_rca24_and1_f_s_pg_rca24_or0_y0 & f_s_pg_rca24_and1_f_s_pg_rca24_fa1_y0;
  assign f_s_pg_rca24_or1_f_s_pg_rca24_and1_y0 = f_s_pg_rca24_and1_y0;
  assign f_s_pg_rca24_or1_f_s_pg_rca24_fa1_y1 = f_s_pg_rca24_fa1_y1;
  assign f_s_pg_rca24_or1_y0 = f_s_pg_rca24_or1_f_s_pg_rca24_and1_y0 | f_s_pg_rca24_or1_f_s_pg_rca24_fa1_y1;
  assign f_s_pg_rca24_fa2_a_2 = a_2;
  assign f_s_pg_rca24_fa2_b_2 = b_2;
  assign f_s_pg_rca24_fa2_f_s_pg_rca24_or1_y0 = f_s_pg_rca24_or1_y0;
  assign f_s_pg_rca24_fa2_y0 = f_s_pg_rca24_fa2_a_2 ^ f_s_pg_rca24_fa2_b_2;
  assign f_s_pg_rca24_fa2_y1 = f_s_pg_rca24_fa2_a_2 & f_s_pg_rca24_fa2_b_2;
  assign f_s_pg_rca24_fa2_y2 = f_s_pg_rca24_fa2_y0 ^ f_s_pg_rca24_fa2_f_s_pg_rca24_or1_y0;
  assign f_s_pg_rca24_and2_f_s_pg_rca24_or1_y0 = f_s_pg_rca24_or1_y0;
  assign f_s_pg_rca24_and2_f_s_pg_rca24_fa2_y0 = f_s_pg_rca24_fa2_y0;
  assign f_s_pg_rca24_and2_y0 = f_s_pg_rca24_and2_f_s_pg_rca24_or1_y0 & f_s_pg_rca24_and2_f_s_pg_rca24_fa2_y0;
  assign f_s_pg_rca24_or2_f_s_pg_rca24_and2_y0 = f_s_pg_rca24_and2_y0;
  assign f_s_pg_rca24_or2_f_s_pg_rca24_fa2_y1 = f_s_pg_rca24_fa2_y1;
  assign f_s_pg_rca24_or2_y0 = f_s_pg_rca24_or2_f_s_pg_rca24_and2_y0 | f_s_pg_rca24_or2_f_s_pg_rca24_fa2_y1;
  assign f_s_pg_rca24_fa3_a_3 = a_3;
  assign f_s_pg_rca24_fa3_b_3 = b_3;
  assign f_s_pg_rca24_fa3_f_s_pg_rca24_or2_y0 = f_s_pg_rca24_or2_y0;
  assign f_s_pg_rca24_fa3_y0 = f_s_pg_rca24_fa3_a_3 ^ f_s_pg_rca24_fa3_b_3;
  assign f_s_pg_rca24_fa3_y1 = f_s_pg_rca24_fa3_a_3 & f_s_pg_rca24_fa3_b_3;
  assign f_s_pg_rca24_fa3_y2 = f_s_pg_rca24_fa3_y0 ^ f_s_pg_rca24_fa3_f_s_pg_rca24_or2_y0;
  assign f_s_pg_rca24_and3_f_s_pg_rca24_or2_y0 = f_s_pg_rca24_or2_y0;
  assign f_s_pg_rca24_and3_f_s_pg_rca24_fa3_y0 = f_s_pg_rca24_fa3_y0;
  assign f_s_pg_rca24_and3_y0 = f_s_pg_rca24_and3_f_s_pg_rca24_or2_y0 & f_s_pg_rca24_and3_f_s_pg_rca24_fa3_y0;
  assign f_s_pg_rca24_or3_f_s_pg_rca24_and3_y0 = f_s_pg_rca24_and3_y0;
  assign f_s_pg_rca24_or3_f_s_pg_rca24_fa3_y1 = f_s_pg_rca24_fa3_y1;
  assign f_s_pg_rca24_or3_y0 = f_s_pg_rca24_or3_f_s_pg_rca24_and3_y0 | f_s_pg_rca24_or3_f_s_pg_rca24_fa3_y1;
  assign f_s_pg_rca24_fa4_a_4 = a_4;
  assign f_s_pg_rca24_fa4_b_4 = b_4;
  assign f_s_pg_rca24_fa4_f_s_pg_rca24_or3_y0 = f_s_pg_rca24_or3_y0;
  assign f_s_pg_rca24_fa4_y0 = f_s_pg_rca24_fa4_a_4 ^ f_s_pg_rca24_fa4_b_4;
  assign f_s_pg_rca24_fa4_y1 = f_s_pg_rca24_fa4_a_4 & f_s_pg_rca24_fa4_b_4;
  assign f_s_pg_rca24_fa4_y2 = f_s_pg_rca24_fa4_y0 ^ f_s_pg_rca24_fa4_f_s_pg_rca24_or3_y0;
  assign f_s_pg_rca24_and4_f_s_pg_rca24_or3_y0 = f_s_pg_rca24_or3_y0;
  assign f_s_pg_rca24_and4_f_s_pg_rca24_fa4_y0 = f_s_pg_rca24_fa4_y0;
  assign f_s_pg_rca24_and4_y0 = f_s_pg_rca24_and4_f_s_pg_rca24_or3_y0 & f_s_pg_rca24_and4_f_s_pg_rca24_fa4_y0;
  assign f_s_pg_rca24_or4_f_s_pg_rca24_and4_y0 = f_s_pg_rca24_and4_y0;
  assign f_s_pg_rca24_or4_f_s_pg_rca24_fa4_y1 = f_s_pg_rca24_fa4_y1;
  assign f_s_pg_rca24_or4_y0 = f_s_pg_rca24_or4_f_s_pg_rca24_and4_y0 | f_s_pg_rca24_or4_f_s_pg_rca24_fa4_y1;
  assign f_s_pg_rca24_fa5_a_5 = a_5;
  assign f_s_pg_rca24_fa5_b_5 = b_5;
  assign f_s_pg_rca24_fa5_f_s_pg_rca24_or4_y0 = f_s_pg_rca24_or4_y0;
  assign f_s_pg_rca24_fa5_y0 = f_s_pg_rca24_fa5_a_5 ^ f_s_pg_rca24_fa5_b_5;
  assign f_s_pg_rca24_fa5_y1 = f_s_pg_rca24_fa5_a_5 & f_s_pg_rca24_fa5_b_5;
  assign f_s_pg_rca24_fa5_y2 = f_s_pg_rca24_fa5_y0 ^ f_s_pg_rca24_fa5_f_s_pg_rca24_or4_y0;
  assign f_s_pg_rca24_and5_f_s_pg_rca24_or4_y0 = f_s_pg_rca24_or4_y0;
  assign f_s_pg_rca24_and5_f_s_pg_rca24_fa5_y0 = f_s_pg_rca24_fa5_y0;
  assign f_s_pg_rca24_and5_y0 = f_s_pg_rca24_and5_f_s_pg_rca24_or4_y0 & f_s_pg_rca24_and5_f_s_pg_rca24_fa5_y0;
  assign f_s_pg_rca24_or5_f_s_pg_rca24_and5_y0 = f_s_pg_rca24_and5_y0;
  assign f_s_pg_rca24_or5_f_s_pg_rca24_fa5_y1 = f_s_pg_rca24_fa5_y1;
  assign f_s_pg_rca24_or5_y0 = f_s_pg_rca24_or5_f_s_pg_rca24_and5_y0 | f_s_pg_rca24_or5_f_s_pg_rca24_fa5_y1;
  assign f_s_pg_rca24_fa6_a_6 = a_6;
  assign f_s_pg_rca24_fa6_b_6 = b_6;
  assign f_s_pg_rca24_fa6_f_s_pg_rca24_or5_y0 = f_s_pg_rca24_or5_y0;
  assign f_s_pg_rca24_fa6_y0 = f_s_pg_rca24_fa6_a_6 ^ f_s_pg_rca24_fa6_b_6;
  assign f_s_pg_rca24_fa6_y1 = f_s_pg_rca24_fa6_a_6 & f_s_pg_rca24_fa6_b_6;
  assign f_s_pg_rca24_fa6_y2 = f_s_pg_rca24_fa6_y0 ^ f_s_pg_rca24_fa6_f_s_pg_rca24_or5_y0;
  assign f_s_pg_rca24_and6_f_s_pg_rca24_or5_y0 = f_s_pg_rca24_or5_y0;
  assign f_s_pg_rca24_and6_f_s_pg_rca24_fa6_y0 = f_s_pg_rca24_fa6_y0;
  assign f_s_pg_rca24_and6_y0 = f_s_pg_rca24_and6_f_s_pg_rca24_or5_y0 & f_s_pg_rca24_and6_f_s_pg_rca24_fa6_y0;
  assign f_s_pg_rca24_or6_f_s_pg_rca24_and6_y0 = f_s_pg_rca24_and6_y0;
  assign f_s_pg_rca24_or6_f_s_pg_rca24_fa6_y1 = f_s_pg_rca24_fa6_y1;
  assign f_s_pg_rca24_or6_y0 = f_s_pg_rca24_or6_f_s_pg_rca24_and6_y0 | f_s_pg_rca24_or6_f_s_pg_rca24_fa6_y1;
  assign f_s_pg_rca24_fa7_a_7 = a_7;
  assign f_s_pg_rca24_fa7_b_7 = b_7;
  assign f_s_pg_rca24_fa7_f_s_pg_rca24_or6_y0 = f_s_pg_rca24_or6_y0;
  assign f_s_pg_rca24_fa7_y0 = f_s_pg_rca24_fa7_a_7 ^ f_s_pg_rca24_fa7_b_7;
  assign f_s_pg_rca24_fa7_y1 = f_s_pg_rca24_fa7_a_7 & f_s_pg_rca24_fa7_b_7;
  assign f_s_pg_rca24_fa7_y2 = f_s_pg_rca24_fa7_y0 ^ f_s_pg_rca24_fa7_f_s_pg_rca24_or6_y0;
  assign f_s_pg_rca24_and7_f_s_pg_rca24_or6_y0 = f_s_pg_rca24_or6_y0;
  assign f_s_pg_rca24_and7_f_s_pg_rca24_fa7_y0 = f_s_pg_rca24_fa7_y0;
  assign f_s_pg_rca24_and7_y0 = f_s_pg_rca24_and7_f_s_pg_rca24_or6_y0 & f_s_pg_rca24_and7_f_s_pg_rca24_fa7_y0;
  assign f_s_pg_rca24_or7_f_s_pg_rca24_and7_y0 = f_s_pg_rca24_and7_y0;
  assign f_s_pg_rca24_or7_f_s_pg_rca24_fa7_y1 = f_s_pg_rca24_fa7_y1;
  assign f_s_pg_rca24_or7_y0 = f_s_pg_rca24_or7_f_s_pg_rca24_and7_y0 | f_s_pg_rca24_or7_f_s_pg_rca24_fa7_y1;
  assign f_s_pg_rca24_fa8_a_8 = a_8;
  assign f_s_pg_rca24_fa8_b_8 = b_8;
  assign f_s_pg_rca24_fa8_f_s_pg_rca24_or7_y0 = f_s_pg_rca24_or7_y0;
  assign f_s_pg_rca24_fa8_y0 = f_s_pg_rca24_fa8_a_8 ^ f_s_pg_rca24_fa8_b_8;
  assign f_s_pg_rca24_fa8_y1 = f_s_pg_rca24_fa8_a_8 & f_s_pg_rca24_fa8_b_8;
  assign f_s_pg_rca24_fa8_y2 = f_s_pg_rca24_fa8_y0 ^ f_s_pg_rca24_fa8_f_s_pg_rca24_or7_y0;
  assign f_s_pg_rca24_and8_f_s_pg_rca24_or7_y0 = f_s_pg_rca24_or7_y0;
  assign f_s_pg_rca24_and8_f_s_pg_rca24_fa8_y0 = f_s_pg_rca24_fa8_y0;
  assign f_s_pg_rca24_and8_y0 = f_s_pg_rca24_and8_f_s_pg_rca24_or7_y0 & f_s_pg_rca24_and8_f_s_pg_rca24_fa8_y0;
  assign f_s_pg_rca24_or8_f_s_pg_rca24_and8_y0 = f_s_pg_rca24_and8_y0;
  assign f_s_pg_rca24_or8_f_s_pg_rca24_fa8_y1 = f_s_pg_rca24_fa8_y1;
  assign f_s_pg_rca24_or8_y0 = f_s_pg_rca24_or8_f_s_pg_rca24_and8_y0 | f_s_pg_rca24_or8_f_s_pg_rca24_fa8_y1;
  assign f_s_pg_rca24_fa9_a_9 = a_9;
  assign f_s_pg_rca24_fa9_b_9 = b_9;
  assign f_s_pg_rca24_fa9_f_s_pg_rca24_or8_y0 = f_s_pg_rca24_or8_y0;
  assign f_s_pg_rca24_fa9_y0 = f_s_pg_rca24_fa9_a_9 ^ f_s_pg_rca24_fa9_b_9;
  assign f_s_pg_rca24_fa9_y1 = f_s_pg_rca24_fa9_a_9 & f_s_pg_rca24_fa9_b_9;
  assign f_s_pg_rca24_fa9_y2 = f_s_pg_rca24_fa9_y0 ^ f_s_pg_rca24_fa9_f_s_pg_rca24_or8_y0;
  assign f_s_pg_rca24_and9_f_s_pg_rca24_or8_y0 = f_s_pg_rca24_or8_y0;
  assign f_s_pg_rca24_and9_f_s_pg_rca24_fa9_y0 = f_s_pg_rca24_fa9_y0;
  assign f_s_pg_rca24_and9_y0 = f_s_pg_rca24_and9_f_s_pg_rca24_or8_y0 & f_s_pg_rca24_and9_f_s_pg_rca24_fa9_y0;
  assign f_s_pg_rca24_or9_f_s_pg_rca24_and9_y0 = f_s_pg_rca24_and9_y0;
  assign f_s_pg_rca24_or9_f_s_pg_rca24_fa9_y1 = f_s_pg_rca24_fa9_y1;
  assign f_s_pg_rca24_or9_y0 = f_s_pg_rca24_or9_f_s_pg_rca24_and9_y0 | f_s_pg_rca24_or9_f_s_pg_rca24_fa9_y1;
  assign f_s_pg_rca24_fa10_a_10 = a_10;
  assign f_s_pg_rca24_fa10_b_10 = b_10;
  assign f_s_pg_rca24_fa10_f_s_pg_rca24_or9_y0 = f_s_pg_rca24_or9_y0;
  assign f_s_pg_rca24_fa10_y0 = f_s_pg_rca24_fa10_a_10 ^ f_s_pg_rca24_fa10_b_10;
  assign f_s_pg_rca24_fa10_y1 = f_s_pg_rca24_fa10_a_10 & f_s_pg_rca24_fa10_b_10;
  assign f_s_pg_rca24_fa10_y2 = f_s_pg_rca24_fa10_y0 ^ f_s_pg_rca24_fa10_f_s_pg_rca24_or9_y0;
  assign f_s_pg_rca24_and10_f_s_pg_rca24_or9_y0 = f_s_pg_rca24_or9_y0;
  assign f_s_pg_rca24_and10_f_s_pg_rca24_fa10_y0 = f_s_pg_rca24_fa10_y0;
  assign f_s_pg_rca24_and10_y0 = f_s_pg_rca24_and10_f_s_pg_rca24_or9_y0 & f_s_pg_rca24_and10_f_s_pg_rca24_fa10_y0;
  assign f_s_pg_rca24_or10_f_s_pg_rca24_and10_y0 = f_s_pg_rca24_and10_y0;
  assign f_s_pg_rca24_or10_f_s_pg_rca24_fa10_y1 = f_s_pg_rca24_fa10_y1;
  assign f_s_pg_rca24_or10_y0 = f_s_pg_rca24_or10_f_s_pg_rca24_and10_y0 | f_s_pg_rca24_or10_f_s_pg_rca24_fa10_y1;
  assign f_s_pg_rca24_fa11_a_11 = a_11;
  assign f_s_pg_rca24_fa11_b_11 = b_11;
  assign f_s_pg_rca24_fa11_f_s_pg_rca24_or10_y0 = f_s_pg_rca24_or10_y0;
  assign f_s_pg_rca24_fa11_y0 = f_s_pg_rca24_fa11_a_11 ^ f_s_pg_rca24_fa11_b_11;
  assign f_s_pg_rca24_fa11_y1 = f_s_pg_rca24_fa11_a_11 & f_s_pg_rca24_fa11_b_11;
  assign f_s_pg_rca24_fa11_y2 = f_s_pg_rca24_fa11_y0 ^ f_s_pg_rca24_fa11_f_s_pg_rca24_or10_y0;
  assign f_s_pg_rca24_and11_f_s_pg_rca24_or10_y0 = f_s_pg_rca24_or10_y0;
  assign f_s_pg_rca24_and11_f_s_pg_rca24_fa11_y0 = f_s_pg_rca24_fa11_y0;
  assign f_s_pg_rca24_and11_y0 = f_s_pg_rca24_and11_f_s_pg_rca24_or10_y0 & f_s_pg_rca24_and11_f_s_pg_rca24_fa11_y0;
  assign f_s_pg_rca24_or11_f_s_pg_rca24_and11_y0 = f_s_pg_rca24_and11_y0;
  assign f_s_pg_rca24_or11_f_s_pg_rca24_fa11_y1 = f_s_pg_rca24_fa11_y1;
  assign f_s_pg_rca24_or11_y0 = f_s_pg_rca24_or11_f_s_pg_rca24_and11_y0 | f_s_pg_rca24_or11_f_s_pg_rca24_fa11_y1;
  assign f_s_pg_rca24_fa12_a_12 = a_12;
  assign f_s_pg_rca24_fa12_b_12 = b_12;
  assign f_s_pg_rca24_fa12_f_s_pg_rca24_or11_y0 = f_s_pg_rca24_or11_y0;
  assign f_s_pg_rca24_fa12_y0 = f_s_pg_rca24_fa12_a_12 ^ f_s_pg_rca24_fa12_b_12;
  assign f_s_pg_rca24_fa12_y1 = f_s_pg_rca24_fa12_a_12 & f_s_pg_rca24_fa12_b_12;
  assign f_s_pg_rca24_fa12_y2 = f_s_pg_rca24_fa12_y0 ^ f_s_pg_rca24_fa12_f_s_pg_rca24_or11_y0;
  assign f_s_pg_rca24_and12_f_s_pg_rca24_or11_y0 = f_s_pg_rca24_or11_y0;
  assign f_s_pg_rca24_and12_f_s_pg_rca24_fa12_y0 = f_s_pg_rca24_fa12_y0;
  assign f_s_pg_rca24_and12_y0 = f_s_pg_rca24_and12_f_s_pg_rca24_or11_y0 & f_s_pg_rca24_and12_f_s_pg_rca24_fa12_y0;
  assign f_s_pg_rca24_or12_f_s_pg_rca24_and12_y0 = f_s_pg_rca24_and12_y0;
  assign f_s_pg_rca24_or12_f_s_pg_rca24_fa12_y1 = f_s_pg_rca24_fa12_y1;
  assign f_s_pg_rca24_or12_y0 = f_s_pg_rca24_or12_f_s_pg_rca24_and12_y0 | f_s_pg_rca24_or12_f_s_pg_rca24_fa12_y1;
  assign f_s_pg_rca24_fa13_a_13 = a_13;
  assign f_s_pg_rca24_fa13_b_13 = b_13;
  assign f_s_pg_rca24_fa13_f_s_pg_rca24_or12_y0 = f_s_pg_rca24_or12_y0;
  assign f_s_pg_rca24_fa13_y0 = f_s_pg_rca24_fa13_a_13 ^ f_s_pg_rca24_fa13_b_13;
  assign f_s_pg_rca24_fa13_y1 = f_s_pg_rca24_fa13_a_13 & f_s_pg_rca24_fa13_b_13;
  assign f_s_pg_rca24_fa13_y2 = f_s_pg_rca24_fa13_y0 ^ f_s_pg_rca24_fa13_f_s_pg_rca24_or12_y0;
  assign f_s_pg_rca24_and13_f_s_pg_rca24_or12_y0 = f_s_pg_rca24_or12_y0;
  assign f_s_pg_rca24_and13_f_s_pg_rca24_fa13_y0 = f_s_pg_rca24_fa13_y0;
  assign f_s_pg_rca24_and13_y0 = f_s_pg_rca24_and13_f_s_pg_rca24_or12_y0 & f_s_pg_rca24_and13_f_s_pg_rca24_fa13_y0;
  assign f_s_pg_rca24_or13_f_s_pg_rca24_and13_y0 = f_s_pg_rca24_and13_y0;
  assign f_s_pg_rca24_or13_f_s_pg_rca24_fa13_y1 = f_s_pg_rca24_fa13_y1;
  assign f_s_pg_rca24_or13_y0 = f_s_pg_rca24_or13_f_s_pg_rca24_and13_y0 | f_s_pg_rca24_or13_f_s_pg_rca24_fa13_y1;
  assign f_s_pg_rca24_fa14_a_14 = a_14;
  assign f_s_pg_rca24_fa14_b_14 = b_14;
  assign f_s_pg_rca24_fa14_f_s_pg_rca24_or13_y0 = f_s_pg_rca24_or13_y0;
  assign f_s_pg_rca24_fa14_y0 = f_s_pg_rca24_fa14_a_14 ^ f_s_pg_rca24_fa14_b_14;
  assign f_s_pg_rca24_fa14_y1 = f_s_pg_rca24_fa14_a_14 & f_s_pg_rca24_fa14_b_14;
  assign f_s_pg_rca24_fa14_y2 = f_s_pg_rca24_fa14_y0 ^ f_s_pg_rca24_fa14_f_s_pg_rca24_or13_y0;
  assign f_s_pg_rca24_and14_f_s_pg_rca24_or13_y0 = f_s_pg_rca24_or13_y0;
  assign f_s_pg_rca24_and14_f_s_pg_rca24_fa14_y0 = f_s_pg_rca24_fa14_y0;
  assign f_s_pg_rca24_and14_y0 = f_s_pg_rca24_and14_f_s_pg_rca24_or13_y0 & f_s_pg_rca24_and14_f_s_pg_rca24_fa14_y0;
  assign f_s_pg_rca24_or14_f_s_pg_rca24_and14_y0 = f_s_pg_rca24_and14_y0;
  assign f_s_pg_rca24_or14_f_s_pg_rca24_fa14_y1 = f_s_pg_rca24_fa14_y1;
  assign f_s_pg_rca24_or14_y0 = f_s_pg_rca24_or14_f_s_pg_rca24_and14_y0 | f_s_pg_rca24_or14_f_s_pg_rca24_fa14_y1;
  assign f_s_pg_rca24_fa15_a_15 = a_15;
  assign f_s_pg_rca24_fa15_b_15 = b_15;
  assign f_s_pg_rca24_fa15_f_s_pg_rca24_or14_y0 = f_s_pg_rca24_or14_y0;
  assign f_s_pg_rca24_fa15_y0 = f_s_pg_rca24_fa15_a_15 ^ f_s_pg_rca24_fa15_b_15;
  assign f_s_pg_rca24_fa15_y1 = f_s_pg_rca24_fa15_a_15 & f_s_pg_rca24_fa15_b_15;
  assign f_s_pg_rca24_fa15_y2 = f_s_pg_rca24_fa15_y0 ^ f_s_pg_rca24_fa15_f_s_pg_rca24_or14_y0;
  assign f_s_pg_rca24_and15_f_s_pg_rca24_or14_y0 = f_s_pg_rca24_or14_y0;
  assign f_s_pg_rca24_and15_f_s_pg_rca24_fa15_y0 = f_s_pg_rca24_fa15_y0;
  assign f_s_pg_rca24_and15_y0 = f_s_pg_rca24_and15_f_s_pg_rca24_or14_y0 & f_s_pg_rca24_and15_f_s_pg_rca24_fa15_y0;
  assign f_s_pg_rca24_or15_f_s_pg_rca24_and15_y0 = f_s_pg_rca24_and15_y0;
  assign f_s_pg_rca24_or15_f_s_pg_rca24_fa15_y1 = f_s_pg_rca24_fa15_y1;
  assign f_s_pg_rca24_or15_y0 = f_s_pg_rca24_or15_f_s_pg_rca24_and15_y0 | f_s_pg_rca24_or15_f_s_pg_rca24_fa15_y1;
  assign f_s_pg_rca24_fa16_a_16 = a_16;
  assign f_s_pg_rca24_fa16_b_16 = b_16;
  assign f_s_pg_rca24_fa16_f_s_pg_rca24_or15_y0 = f_s_pg_rca24_or15_y0;
  assign f_s_pg_rca24_fa16_y0 = f_s_pg_rca24_fa16_a_16 ^ f_s_pg_rca24_fa16_b_16;
  assign f_s_pg_rca24_fa16_y1 = f_s_pg_rca24_fa16_a_16 & f_s_pg_rca24_fa16_b_16;
  assign f_s_pg_rca24_fa16_y2 = f_s_pg_rca24_fa16_y0 ^ f_s_pg_rca24_fa16_f_s_pg_rca24_or15_y0;
  assign f_s_pg_rca24_and16_f_s_pg_rca24_or15_y0 = f_s_pg_rca24_or15_y0;
  assign f_s_pg_rca24_and16_f_s_pg_rca24_fa16_y0 = f_s_pg_rca24_fa16_y0;
  assign f_s_pg_rca24_and16_y0 = f_s_pg_rca24_and16_f_s_pg_rca24_or15_y0 & f_s_pg_rca24_and16_f_s_pg_rca24_fa16_y0;
  assign f_s_pg_rca24_or16_f_s_pg_rca24_and16_y0 = f_s_pg_rca24_and16_y0;
  assign f_s_pg_rca24_or16_f_s_pg_rca24_fa16_y1 = f_s_pg_rca24_fa16_y1;
  assign f_s_pg_rca24_or16_y0 = f_s_pg_rca24_or16_f_s_pg_rca24_and16_y0 | f_s_pg_rca24_or16_f_s_pg_rca24_fa16_y1;
  assign f_s_pg_rca24_fa17_a_17 = a_17;
  assign f_s_pg_rca24_fa17_b_17 = b_17;
  assign f_s_pg_rca24_fa17_f_s_pg_rca24_or16_y0 = f_s_pg_rca24_or16_y0;
  assign f_s_pg_rca24_fa17_y0 = f_s_pg_rca24_fa17_a_17 ^ f_s_pg_rca24_fa17_b_17;
  assign f_s_pg_rca24_fa17_y1 = f_s_pg_rca24_fa17_a_17 & f_s_pg_rca24_fa17_b_17;
  assign f_s_pg_rca24_fa17_y2 = f_s_pg_rca24_fa17_y0 ^ f_s_pg_rca24_fa17_f_s_pg_rca24_or16_y0;
  assign f_s_pg_rca24_and17_f_s_pg_rca24_or16_y0 = f_s_pg_rca24_or16_y0;
  assign f_s_pg_rca24_and17_f_s_pg_rca24_fa17_y0 = f_s_pg_rca24_fa17_y0;
  assign f_s_pg_rca24_and17_y0 = f_s_pg_rca24_and17_f_s_pg_rca24_or16_y0 & f_s_pg_rca24_and17_f_s_pg_rca24_fa17_y0;
  assign f_s_pg_rca24_or17_f_s_pg_rca24_and17_y0 = f_s_pg_rca24_and17_y0;
  assign f_s_pg_rca24_or17_f_s_pg_rca24_fa17_y1 = f_s_pg_rca24_fa17_y1;
  assign f_s_pg_rca24_or17_y0 = f_s_pg_rca24_or17_f_s_pg_rca24_and17_y0 | f_s_pg_rca24_or17_f_s_pg_rca24_fa17_y1;
  assign f_s_pg_rca24_fa18_a_18 = a_18;
  assign f_s_pg_rca24_fa18_b_18 = b_18;
  assign f_s_pg_rca24_fa18_f_s_pg_rca24_or17_y0 = f_s_pg_rca24_or17_y0;
  assign f_s_pg_rca24_fa18_y0 = f_s_pg_rca24_fa18_a_18 ^ f_s_pg_rca24_fa18_b_18;
  assign f_s_pg_rca24_fa18_y1 = f_s_pg_rca24_fa18_a_18 & f_s_pg_rca24_fa18_b_18;
  assign f_s_pg_rca24_fa18_y2 = f_s_pg_rca24_fa18_y0 ^ f_s_pg_rca24_fa18_f_s_pg_rca24_or17_y0;
  assign f_s_pg_rca24_and18_f_s_pg_rca24_or17_y0 = f_s_pg_rca24_or17_y0;
  assign f_s_pg_rca24_and18_f_s_pg_rca24_fa18_y0 = f_s_pg_rca24_fa18_y0;
  assign f_s_pg_rca24_and18_y0 = f_s_pg_rca24_and18_f_s_pg_rca24_or17_y0 & f_s_pg_rca24_and18_f_s_pg_rca24_fa18_y0;
  assign f_s_pg_rca24_or18_f_s_pg_rca24_and18_y0 = f_s_pg_rca24_and18_y0;
  assign f_s_pg_rca24_or18_f_s_pg_rca24_fa18_y1 = f_s_pg_rca24_fa18_y1;
  assign f_s_pg_rca24_or18_y0 = f_s_pg_rca24_or18_f_s_pg_rca24_and18_y0 | f_s_pg_rca24_or18_f_s_pg_rca24_fa18_y1;
  assign f_s_pg_rca24_fa19_a_19 = a_19;
  assign f_s_pg_rca24_fa19_b_19 = b_19;
  assign f_s_pg_rca24_fa19_f_s_pg_rca24_or18_y0 = f_s_pg_rca24_or18_y0;
  assign f_s_pg_rca24_fa19_y0 = f_s_pg_rca24_fa19_a_19 ^ f_s_pg_rca24_fa19_b_19;
  assign f_s_pg_rca24_fa19_y1 = f_s_pg_rca24_fa19_a_19 & f_s_pg_rca24_fa19_b_19;
  assign f_s_pg_rca24_fa19_y2 = f_s_pg_rca24_fa19_y0 ^ f_s_pg_rca24_fa19_f_s_pg_rca24_or18_y0;
  assign f_s_pg_rca24_and19_f_s_pg_rca24_or18_y0 = f_s_pg_rca24_or18_y0;
  assign f_s_pg_rca24_and19_f_s_pg_rca24_fa19_y0 = f_s_pg_rca24_fa19_y0;
  assign f_s_pg_rca24_and19_y0 = f_s_pg_rca24_and19_f_s_pg_rca24_or18_y0 & f_s_pg_rca24_and19_f_s_pg_rca24_fa19_y0;
  assign f_s_pg_rca24_or19_f_s_pg_rca24_and19_y0 = f_s_pg_rca24_and19_y0;
  assign f_s_pg_rca24_or19_f_s_pg_rca24_fa19_y1 = f_s_pg_rca24_fa19_y1;
  assign f_s_pg_rca24_or19_y0 = f_s_pg_rca24_or19_f_s_pg_rca24_and19_y0 | f_s_pg_rca24_or19_f_s_pg_rca24_fa19_y1;
  assign f_s_pg_rca24_fa20_a_20 = a_20;
  assign f_s_pg_rca24_fa20_b_20 = b_20;
  assign f_s_pg_rca24_fa20_f_s_pg_rca24_or19_y0 = f_s_pg_rca24_or19_y0;
  assign f_s_pg_rca24_fa20_y0 = f_s_pg_rca24_fa20_a_20 ^ f_s_pg_rca24_fa20_b_20;
  assign f_s_pg_rca24_fa20_y1 = f_s_pg_rca24_fa20_a_20 & f_s_pg_rca24_fa20_b_20;
  assign f_s_pg_rca24_fa20_y2 = f_s_pg_rca24_fa20_y0 ^ f_s_pg_rca24_fa20_f_s_pg_rca24_or19_y0;
  assign f_s_pg_rca24_and20_f_s_pg_rca24_or19_y0 = f_s_pg_rca24_or19_y0;
  assign f_s_pg_rca24_and20_f_s_pg_rca24_fa20_y0 = f_s_pg_rca24_fa20_y0;
  assign f_s_pg_rca24_and20_y0 = f_s_pg_rca24_and20_f_s_pg_rca24_or19_y0 & f_s_pg_rca24_and20_f_s_pg_rca24_fa20_y0;
  assign f_s_pg_rca24_or20_f_s_pg_rca24_and20_y0 = f_s_pg_rca24_and20_y0;
  assign f_s_pg_rca24_or20_f_s_pg_rca24_fa20_y1 = f_s_pg_rca24_fa20_y1;
  assign f_s_pg_rca24_or20_y0 = f_s_pg_rca24_or20_f_s_pg_rca24_and20_y0 | f_s_pg_rca24_or20_f_s_pg_rca24_fa20_y1;
  assign f_s_pg_rca24_fa21_a_21 = a_21;
  assign f_s_pg_rca24_fa21_b_21 = b_21;
  assign f_s_pg_rca24_fa21_f_s_pg_rca24_or20_y0 = f_s_pg_rca24_or20_y0;
  assign f_s_pg_rca24_fa21_y0 = f_s_pg_rca24_fa21_a_21 ^ f_s_pg_rca24_fa21_b_21;
  assign f_s_pg_rca24_fa21_y1 = f_s_pg_rca24_fa21_a_21 & f_s_pg_rca24_fa21_b_21;
  assign f_s_pg_rca24_fa21_y2 = f_s_pg_rca24_fa21_y0 ^ f_s_pg_rca24_fa21_f_s_pg_rca24_or20_y0;
  assign f_s_pg_rca24_and21_f_s_pg_rca24_or20_y0 = f_s_pg_rca24_or20_y0;
  assign f_s_pg_rca24_and21_f_s_pg_rca24_fa21_y0 = f_s_pg_rca24_fa21_y0;
  assign f_s_pg_rca24_and21_y0 = f_s_pg_rca24_and21_f_s_pg_rca24_or20_y0 & f_s_pg_rca24_and21_f_s_pg_rca24_fa21_y0;
  assign f_s_pg_rca24_or21_f_s_pg_rca24_and21_y0 = f_s_pg_rca24_and21_y0;
  assign f_s_pg_rca24_or21_f_s_pg_rca24_fa21_y1 = f_s_pg_rca24_fa21_y1;
  assign f_s_pg_rca24_or21_y0 = f_s_pg_rca24_or21_f_s_pg_rca24_and21_y0 | f_s_pg_rca24_or21_f_s_pg_rca24_fa21_y1;
  assign f_s_pg_rca24_fa22_a_22 = a_22;
  assign f_s_pg_rca24_fa22_b_22 = b_22;
  assign f_s_pg_rca24_fa22_f_s_pg_rca24_or21_y0 = f_s_pg_rca24_or21_y0;
  assign f_s_pg_rca24_fa22_y0 = f_s_pg_rca24_fa22_a_22 ^ f_s_pg_rca24_fa22_b_22;
  assign f_s_pg_rca24_fa22_y1 = f_s_pg_rca24_fa22_a_22 & f_s_pg_rca24_fa22_b_22;
  assign f_s_pg_rca24_fa22_y2 = f_s_pg_rca24_fa22_y0 ^ f_s_pg_rca24_fa22_f_s_pg_rca24_or21_y0;
  assign f_s_pg_rca24_and22_f_s_pg_rca24_or21_y0 = f_s_pg_rca24_or21_y0;
  assign f_s_pg_rca24_and22_f_s_pg_rca24_fa22_y0 = f_s_pg_rca24_fa22_y0;
  assign f_s_pg_rca24_and22_y0 = f_s_pg_rca24_and22_f_s_pg_rca24_or21_y0 & f_s_pg_rca24_and22_f_s_pg_rca24_fa22_y0;
  assign f_s_pg_rca24_or22_f_s_pg_rca24_and22_y0 = f_s_pg_rca24_and22_y0;
  assign f_s_pg_rca24_or22_f_s_pg_rca24_fa22_y1 = f_s_pg_rca24_fa22_y1;
  assign f_s_pg_rca24_or22_y0 = f_s_pg_rca24_or22_f_s_pg_rca24_and22_y0 | f_s_pg_rca24_or22_f_s_pg_rca24_fa22_y1;
  assign f_s_pg_rca24_fa23_a_23 = a_23;
  assign f_s_pg_rca24_fa23_b_23 = b_23;
  assign f_s_pg_rca24_fa23_f_s_pg_rca24_or22_y0 = f_s_pg_rca24_or22_y0;
  assign f_s_pg_rca24_fa23_y0 = f_s_pg_rca24_fa23_a_23 ^ f_s_pg_rca24_fa23_b_23;
  assign f_s_pg_rca24_fa23_y1 = f_s_pg_rca24_fa23_a_23 & f_s_pg_rca24_fa23_b_23;
  assign f_s_pg_rca24_fa23_y2 = f_s_pg_rca24_fa23_y0 ^ f_s_pg_rca24_fa23_f_s_pg_rca24_or22_y0;
  assign f_s_pg_rca24_and23_f_s_pg_rca24_or22_y0 = f_s_pg_rca24_or22_y0;
  assign f_s_pg_rca24_and23_f_s_pg_rca24_fa23_y0 = f_s_pg_rca24_fa23_y0;
  assign f_s_pg_rca24_and23_y0 = f_s_pg_rca24_and23_f_s_pg_rca24_or22_y0 & f_s_pg_rca24_and23_f_s_pg_rca24_fa23_y0;
  assign f_s_pg_rca24_or23_f_s_pg_rca24_and23_y0 = f_s_pg_rca24_and23_y0;
  assign f_s_pg_rca24_or23_f_s_pg_rca24_fa23_y1 = f_s_pg_rca24_fa23_y1;
  assign f_s_pg_rca24_or23_y0 = f_s_pg_rca24_or23_f_s_pg_rca24_and23_y0 | f_s_pg_rca24_or23_f_s_pg_rca24_fa23_y1;
  assign f_s_pg_rca24_xor0_a_23 = a_23;
  assign f_s_pg_rca24_xor0_b_23 = b_23;
  assign f_s_pg_rca24_xor0_y0 = f_s_pg_rca24_xor0_a_23 ^ f_s_pg_rca24_xor0_b_23;
  assign f_s_pg_rca24_xor1_f_s_pg_rca24_xor0_y0 = f_s_pg_rca24_xor0_y0;
  assign f_s_pg_rca24_xor1_f_s_pg_rca24_or23_y0 = f_s_pg_rca24_or23_y0;
  assign f_s_pg_rca24_xor1_y0 = f_s_pg_rca24_xor1_f_s_pg_rca24_xor0_y0 ^ f_s_pg_rca24_xor1_f_s_pg_rca24_or23_y0;

  assign out[0] = f_s_pg_rca24_fa0_y2;
  assign out[1] = f_s_pg_rca24_fa1_y2;
  assign out[2] = f_s_pg_rca24_fa2_y2;
  assign out[3] = f_s_pg_rca24_fa3_y2;
  assign out[4] = f_s_pg_rca24_fa4_y2;
  assign out[5] = f_s_pg_rca24_fa5_y2;
  assign out[6] = f_s_pg_rca24_fa6_y2;
  assign out[7] = f_s_pg_rca24_fa7_y2;
  assign out[8] = f_s_pg_rca24_fa8_y2;
  assign out[9] = f_s_pg_rca24_fa9_y2;
  assign out[10] = f_s_pg_rca24_fa10_y2;
  assign out[11] = f_s_pg_rca24_fa11_y2;
  assign out[12] = f_s_pg_rca24_fa12_y2;
  assign out[13] = f_s_pg_rca24_fa13_y2;
  assign out[14] = f_s_pg_rca24_fa14_y2;
  assign out[15] = f_s_pg_rca24_fa15_y2;
  assign out[16] = f_s_pg_rca24_fa16_y2;
  assign out[17] = f_s_pg_rca24_fa17_y2;
  assign out[18] = f_s_pg_rca24_fa18_y2;
  assign out[19] = f_s_pg_rca24_fa19_y2;
  assign out[20] = f_s_pg_rca24_fa20_y2;
  assign out[21] = f_s_pg_rca24_fa21_y2;
  assign out[22] = f_s_pg_rca24_fa22_y2;
  assign out[23] = f_s_pg_rca24_fa23_y2;
  assign out[24] = f_s_pg_rca24_xor1_y0;
endmodule