module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module nand_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a & _b);
endmodule

module constant_wire_value_1(input a, input b, output constant_wire_1);
  wire constant_wire_value_1_a;
  wire constant_wire_value_1_b;

  assign constant_wire_value_1_a = a;
  assign constant_wire_value_1_b = b;

  xor_gate xor_gate_constant_wire_value_1_y0(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y0);
  xnor_gate xnor_gate_constant_wire_value_1_y1(constant_wire_value_1_a, constant_wire_value_1_b, constant_wire_value_1_y1);
  or_gate or_gate_constant_wire_1(constant_wire_value_1_y0, constant_wire_value_1_y1, constant_wire_1);
endmodule

module ha(input a, input b, output ha_y0, output ha_y1);
  wire ha_a;
  wire ha_b;

  assign ha_a = a;
  assign ha_b = b;

  xor_gate xor_gate_ha_y0(ha_a, ha_b, ha_y0);
  and_gate and_gate_ha_y1(ha_a, ha_b, ha_y1);
endmodule

module fa(input a, input b, input cin, output fa_y2, output fa_y4);
  wire fa_a;
  wire fa_b;
  wire fa_cin;

  assign fa_a = a;
  assign fa_b = b;
  assign fa_cin = cin;

  xor_gate xor_gate_fa_y0(fa_a, fa_b, fa_y0);
  and_gate and_gate_fa_y1(fa_a, fa_b, fa_y1);
  xor_gate xor_gate_fa_y2(fa_y0, fa_cin, fa_y2);
  and_gate and_gate_fa_y3(fa_y0, fa_cin, fa_y3);
  or_gate or_gate_fa_y4(fa_y1, fa_y3, fa_y4);
endmodule

module h_s_arrmul24(input [23:0] a, input [23:0] b, output [47:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire constant_wire_1;
  wire h_s_arrmul24_and0_0_y0;
  wire h_s_arrmul24_and1_0_y0;
  wire h_s_arrmul24_and2_0_y0;
  wire h_s_arrmul24_and3_0_y0;
  wire h_s_arrmul24_and4_0_y0;
  wire h_s_arrmul24_and5_0_y0;
  wire h_s_arrmul24_and6_0_y0;
  wire h_s_arrmul24_and7_0_y0;
  wire h_s_arrmul24_and8_0_y0;
  wire h_s_arrmul24_and9_0_y0;
  wire h_s_arrmul24_and10_0_y0;
  wire h_s_arrmul24_and11_0_y0;
  wire h_s_arrmul24_and12_0_y0;
  wire h_s_arrmul24_and13_0_y0;
  wire h_s_arrmul24_and14_0_y0;
  wire h_s_arrmul24_and15_0_y0;
  wire h_s_arrmul24_and16_0_y0;
  wire h_s_arrmul24_and17_0_y0;
  wire h_s_arrmul24_and18_0_y0;
  wire h_s_arrmul24_and19_0_y0;
  wire h_s_arrmul24_and20_0_y0;
  wire h_s_arrmul24_and21_0_y0;
  wire h_s_arrmul24_and22_0_y0;
  wire h_s_arrmul24_nand23_0_y0;
  wire h_s_arrmul24_and0_1_y0;
  wire h_s_arrmul24_ha0_1_y0;
  wire h_s_arrmul24_ha0_1_y1;
  wire h_s_arrmul24_and1_1_y0;
  wire h_s_arrmul24_fa1_1_y2;
  wire h_s_arrmul24_fa1_1_y4;
  wire h_s_arrmul24_and2_1_y0;
  wire h_s_arrmul24_fa2_1_y2;
  wire h_s_arrmul24_fa2_1_y4;
  wire h_s_arrmul24_and3_1_y0;
  wire h_s_arrmul24_fa3_1_y2;
  wire h_s_arrmul24_fa3_1_y4;
  wire h_s_arrmul24_and4_1_y0;
  wire h_s_arrmul24_fa4_1_y2;
  wire h_s_arrmul24_fa4_1_y4;
  wire h_s_arrmul24_and5_1_y0;
  wire h_s_arrmul24_fa5_1_y2;
  wire h_s_arrmul24_fa5_1_y4;
  wire h_s_arrmul24_and6_1_y0;
  wire h_s_arrmul24_fa6_1_y2;
  wire h_s_arrmul24_fa6_1_y4;
  wire h_s_arrmul24_and7_1_y0;
  wire h_s_arrmul24_fa7_1_y2;
  wire h_s_arrmul24_fa7_1_y4;
  wire h_s_arrmul24_and8_1_y0;
  wire h_s_arrmul24_fa8_1_y2;
  wire h_s_arrmul24_fa8_1_y4;
  wire h_s_arrmul24_and9_1_y0;
  wire h_s_arrmul24_fa9_1_y2;
  wire h_s_arrmul24_fa9_1_y4;
  wire h_s_arrmul24_and10_1_y0;
  wire h_s_arrmul24_fa10_1_y2;
  wire h_s_arrmul24_fa10_1_y4;
  wire h_s_arrmul24_and11_1_y0;
  wire h_s_arrmul24_fa11_1_y2;
  wire h_s_arrmul24_fa11_1_y4;
  wire h_s_arrmul24_and12_1_y0;
  wire h_s_arrmul24_fa12_1_y2;
  wire h_s_arrmul24_fa12_1_y4;
  wire h_s_arrmul24_and13_1_y0;
  wire h_s_arrmul24_fa13_1_y2;
  wire h_s_arrmul24_fa13_1_y4;
  wire h_s_arrmul24_and14_1_y0;
  wire h_s_arrmul24_fa14_1_y2;
  wire h_s_arrmul24_fa14_1_y4;
  wire h_s_arrmul24_and15_1_y0;
  wire h_s_arrmul24_fa15_1_y2;
  wire h_s_arrmul24_fa15_1_y4;
  wire h_s_arrmul24_and16_1_y0;
  wire h_s_arrmul24_fa16_1_y2;
  wire h_s_arrmul24_fa16_1_y4;
  wire h_s_arrmul24_and17_1_y0;
  wire h_s_arrmul24_fa17_1_y2;
  wire h_s_arrmul24_fa17_1_y4;
  wire h_s_arrmul24_and18_1_y0;
  wire h_s_arrmul24_fa18_1_y2;
  wire h_s_arrmul24_fa18_1_y4;
  wire h_s_arrmul24_and19_1_y0;
  wire h_s_arrmul24_fa19_1_y2;
  wire h_s_arrmul24_fa19_1_y4;
  wire h_s_arrmul24_and20_1_y0;
  wire h_s_arrmul24_fa20_1_y2;
  wire h_s_arrmul24_fa20_1_y4;
  wire h_s_arrmul24_and21_1_y0;
  wire h_s_arrmul24_fa21_1_y2;
  wire h_s_arrmul24_fa21_1_y4;
  wire h_s_arrmul24_and22_1_y0;
  wire h_s_arrmul24_fa22_1_y2;
  wire h_s_arrmul24_fa22_1_y4;
  wire h_s_arrmul24_nand23_1_y0;
  wire h_s_arrmul24_fa23_1_y2;
  wire h_s_arrmul24_fa23_1_y4;
  wire h_s_arrmul24_and0_2_y0;
  wire h_s_arrmul24_ha0_2_y0;
  wire h_s_arrmul24_ha0_2_y1;
  wire h_s_arrmul24_and1_2_y0;
  wire h_s_arrmul24_fa1_2_y2;
  wire h_s_arrmul24_fa1_2_y4;
  wire h_s_arrmul24_and2_2_y0;
  wire h_s_arrmul24_fa2_2_y2;
  wire h_s_arrmul24_fa2_2_y4;
  wire h_s_arrmul24_and3_2_y0;
  wire h_s_arrmul24_fa3_2_y2;
  wire h_s_arrmul24_fa3_2_y4;
  wire h_s_arrmul24_and4_2_y0;
  wire h_s_arrmul24_fa4_2_y2;
  wire h_s_arrmul24_fa4_2_y4;
  wire h_s_arrmul24_and5_2_y0;
  wire h_s_arrmul24_fa5_2_y2;
  wire h_s_arrmul24_fa5_2_y4;
  wire h_s_arrmul24_and6_2_y0;
  wire h_s_arrmul24_fa6_2_y2;
  wire h_s_arrmul24_fa6_2_y4;
  wire h_s_arrmul24_and7_2_y0;
  wire h_s_arrmul24_fa7_2_y2;
  wire h_s_arrmul24_fa7_2_y4;
  wire h_s_arrmul24_and8_2_y0;
  wire h_s_arrmul24_fa8_2_y2;
  wire h_s_arrmul24_fa8_2_y4;
  wire h_s_arrmul24_and9_2_y0;
  wire h_s_arrmul24_fa9_2_y2;
  wire h_s_arrmul24_fa9_2_y4;
  wire h_s_arrmul24_and10_2_y0;
  wire h_s_arrmul24_fa10_2_y2;
  wire h_s_arrmul24_fa10_2_y4;
  wire h_s_arrmul24_and11_2_y0;
  wire h_s_arrmul24_fa11_2_y2;
  wire h_s_arrmul24_fa11_2_y4;
  wire h_s_arrmul24_and12_2_y0;
  wire h_s_arrmul24_fa12_2_y2;
  wire h_s_arrmul24_fa12_2_y4;
  wire h_s_arrmul24_and13_2_y0;
  wire h_s_arrmul24_fa13_2_y2;
  wire h_s_arrmul24_fa13_2_y4;
  wire h_s_arrmul24_and14_2_y0;
  wire h_s_arrmul24_fa14_2_y2;
  wire h_s_arrmul24_fa14_2_y4;
  wire h_s_arrmul24_and15_2_y0;
  wire h_s_arrmul24_fa15_2_y2;
  wire h_s_arrmul24_fa15_2_y4;
  wire h_s_arrmul24_and16_2_y0;
  wire h_s_arrmul24_fa16_2_y2;
  wire h_s_arrmul24_fa16_2_y4;
  wire h_s_arrmul24_and17_2_y0;
  wire h_s_arrmul24_fa17_2_y2;
  wire h_s_arrmul24_fa17_2_y4;
  wire h_s_arrmul24_and18_2_y0;
  wire h_s_arrmul24_fa18_2_y2;
  wire h_s_arrmul24_fa18_2_y4;
  wire h_s_arrmul24_and19_2_y0;
  wire h_s_arrmul24_fa19_2_y2;
  wire h_s_arrmul24_fa19_2_y4;
  wire h_s_arrmul24_and20_2_y0;
  wire h_s_arrmul24_fa20_2_y2;
  wire h_s_arrmul24_fa20_2_y4;
  wire h_s_arrmul24_and21_2_y0;
  wire h_s_arrmul24_fa21_2_y2;
  wire h_s_arrmul24_fa21_2_y4;
  wire h_s_arrmul24_and22_2_y0;
  wire h_s_arrmul24_fa22_2_y2;
  wire h_s_arrmul24_fa22_2_y4;
  wire h_s_arrmul24_nand23_2_y0;
  wire h_s_arrmul24_fa23_2_y2;
  wire h_s_arrmul24_fa23_2_y4;
  wire h_s_arrmul24_and0_3_y0;
  wire h_s_arrmul24_ha0_3_y0;
  wire h_s_arrmul24_ha0_3_y1;
  wire h_s_arrmul24_and1_3_y0;
  wire h_s_arrmul24_fa1_3_y2;
  wire h_s_arrmul24_fa1_3_y4;
  wire h_s_arrmul24_and2_3_y0;
  wire h_s_arrmul24_fa2_3_y2;
  wire h_s_arrmul24_fa2_3_y4;
  wire h_s_arrmul24_and3_3_y0;
  wire h_s_arrmul24_fa3_3_y2;
  wire h_s_arrmul24_fa3_3_y4;
  wire h_s_arrmul24_and4_3_y0;
  wire h_s_arrmul24_fa4_3_y2;
  wire h_s_arrmul24_fa4_3_y4;
  wire h_s_arrmul24_and5_3_y0;
  wire h_s_arrmul24_fa5_3_y2;
  wire h_s_arrmul24_fa5_3_y4;
  wire h_s_arrmul24_and6_3_y0;
  wire h_s_arrmul24_fa6_3_y2;
  wire h_s_arrmul24_fa6_3_y4;
  wire h_s_arrmul24_and7_3_y0;
  wire h_s_arrmul24_fa7_3_y2;
  wire h_s_arrmul24_fa7_3_y4;
  wire h_s_arrmul24_and8_3_y0;
  wire h_s_arrmul24_fa8_3_y2;
  wire h_s_arrmul24_fa8_3_y4;
  wire h_s_arrmul24_and9_3_y0;
  wire h_s_arrmul24_fa9_3_y2;
  wire h_s_arrmul24_fa9_3_y4;
  wire h_s_arrmul24_and10_3_y0;
  wire h_s_arrmul24_fa10_3_y2;
  wire h_s_arrmul24_fa10_3_y4;
  wire h_s_arrmul24_and11_3_y0;
  wire h_s_arrmul24_fa11_3_y2;
  wire h_s_arrmul24_fa11_3_y4;
  wire h_s_arrmul24_and12_3_y0;
  wire h_s_arrmul24_fa12_3_y2;
  wire h_s_arrmul24_fa12_3_y4;
  wire h_s_arrmul24_and13_3_y0;
  wire h_s_arrmul24_fa13_3_y2;
  wire h_s_arrmul24_fa13_3_y4;
  wire h_s_arrmul24_and14_3_y0;
  wire h_s_arrmul24_fa14_3_y2;
  wire h_s_arrmul24_fa14_3_y4;
  wire h_s_arrmul24_and15_3_y0;
  wire h_s_arrmul24_fa15_3_y2;
  wire h_s_arrmul24_fa15_3_y4;
  wire h_s_arrmul24_and16_3_y0;
  wire h_s_arrmul24_fa16_3_y2;
  wire h_s_arrmul24_fa16_3_y4;
  wire h_s_arrmul24_and17_3_y0;
  wire h_s_arrmul24_fa17_3_y2;
  wire h_s_arrmul24_fa17_3_y4;
  wire h_s_arrmul24_and18_3_y0;
  wire h_s_arrmul24_fa18_3_y2;
  wire h_s_arrmul24_fa18_3_y4;
  wire h_s_arrmul24_and19_3_y0;
  wire h_s_arrmul24_fa19_3_y2;
  wire h_s_arrmul24_fa19_3_y4;
  wire h_s_arrmul24_and20_3_y0;
  wire h_s_arrmul24_fa20_3_y2;
  wire h_s_arrmul24_fa20_3_y4;
  wire h_s_arrmul24_and21_3_y0;
  wire h_s_arrmul24_fa21_3_y2;
  wire h_s_arrmul24_fa21_3_y4;
  wire h_s_arrmul24_and22_3_y0;
  wire h_s_arrmul24_fa22_3_y2;
  wire h_s_arrmul24_fa22_3_y4;
  wire h_s_arrmul24_nand23_3_y0;
  wire h_s_arrmul24_fa23_3_y2;
  wire h_s_arrmul24_fa23_3_y4;
  wire h_s_arrmul24_and0_4_y0;
  wire h_s_arrmul24_ha0_4_y0;
  wire h_s_arrmul24_ha0_4_y1;
  wire h_s_arrmul24_and1_4_y0;
  wire h_s_arrmul24_fa1_4_y2;
  wire h_s_arrmul24_fa1_4_y4;
  wire h_s_arrmul24_and2_4_y0;
  wire h_s_arrmul24_fa2_4_y2;
  wire h_s_arrmul24_fa2_4_y4;
  wire h_s_arrmul24_and3_4_y0;
  wire h_s_arrmul24_fa3_4_y2;
  wire h_s_arrmul24_fa3_4_y4;
  wire h_s_arrmul24_and4_4_y0;
  wire h_s_arrmul24_fa4_4_y2;
  wire h_s_arrmul24_fa4_4_y4;
  wire h_s_arrmul24_and5_4_y0;
  wire h_s_arrmul24_fa5_4_y2;
  wire h_s_arrmul24_fa5_4_y4;
  wire h_s_arrmul24_and6_4_y0;
  wire h_s_arrmul24_fa6_4_y2;
  wire h_s_arrmul24_fa6_4_y4;
  wire h_s_arrmul24_and7_4_y0;
  wire h_s_arrmul24_fa7_4_y2;
  wire h_s_arrmul24_fa7_4_y4;
  wire h_s_arrmul24_and8_4_y0;
  wire h_s_arrmul24_fa8_4_y2;
  wire h_s_arrmul24_fa8_4_y4;
  wire h_s_arrmul24_and9_4_y0;
  wire h_s_arrmul24_fa9_4_y2;
  wire h_s_arrmul24_fa9_4_y4;
  wire h_s_arrmul24_and10_4_y0;
  wire h_s_arrmul24_fa10_4_y2;
  wire h_s_arrmul24_fa10_4_y4;
  wire h_s_arrmul24_and11_4_y0;
  wire h_s_arrmul24_fa11_4_y2;
  wire h_s_arrmul24_fa11_4_y4;
  wire h_s_arrmul24_and12_4_y0;
  wire h_s_arrmul24_fa12_4_y2;
  wire h_s_arrmul24_fa12_4_y4;
  wire h_s_arrmul24_and13_4_y0;
  wire h_s_arrmul24_fa13_4_y2;
  wire h_s_arrmul24_fa13_4_y4;
  wire h_s_arrmul24_and14_4_y0;
  wire h_s_arrmul24_fa14_4_y2;
  wire h_s_arrmul24_fa14_4_y4;
  wire h_s_arrmul24_and15_4_y0;
  wire h_s_arrmul24_fa15_4_y2;
  wire h_s_arrmul24_fa15_4_y4;
  wire h_s_arrmul24_and16_4_y0;
  wire h_s_arrmul24_fa16_4_y2;
  wire h_s_arrmul24_fa16_4_y4;
  wire h_s_arrmul24_and17_4_y0;
  wire h_s_arrmul24_fa17_4_y2;
  wire h_s_arrmul24_fa17_4_y4;
  wire h_s_arrmul24_and18_4_y0;
  wire h_s_arrmul24_fa18_4_y2;
  wire h_s_arrmul24_fa18_4_y4;
  wire h_s_arrmul24_and19_4_y0;
  wire h_s_arrmul24_fa19_4_y2;
  wire h_s_arrmul24_fa19_4_y4;
  wire h_s_arrmul24_and20_4_y0;
  wire h_s_arrmul24_fa20_4_y2;
  wire h_s_arrmul24_fa20_4_y4;
  wire h_s_arrmul24_and21_4_y0;
  wire h_s_arrmul24_fa21_4_y2;
  wire h_s_arrmul24_fa21_4_y4;
  wire h_s_arrmul24_and22_4_y0;
  wire h_s_arrmul24_fa22_4_y2;
  wire h_s_arrmul24_fa22_4_y4;
  wire h_s_arrmul24_nand23_4_y0;
  wire h_s_arrmul24_fa23_4_y2;
  wire h_s_arrmul24_fa23_4_y4;
  wire h_s_arrmul24_and0_5_y0;
  wire h_s_arrmul24_ha0_5_y0;
  wire h_s_arrmul24_ha0_5_y1;
  wire h_s_arrmul24_and1_5_y0;
  wire h_s_arrmul24_fa1_5_y2;
  wire h_s_arrmul24_fa1_5_y4;
  wire h_s_arrmul24_and2_5_y0;
  wire h_s_arrmul24_fa2_5_y2;
  wire h_s_arrmul24_fa2_5_y4;
  wire h_s_arrmul24_and3_5_y0;
  wire h_s_arrmul24_fa3_5_y2;
  wire h_s_arrmul24_fa3_5_y4;
  wire h_s_arrmul24_and4_5_y0;
  wire h_s_arrmul24_fa4_5_y2;
  wire h_s_arrmul24_fa4_5_y4;
  wire h_s_arrmul24_and5_5_y0;
  wire h_s_arrmul24_fa5_5_y2;
  wire h_s_arrmul24_fa5_5_y4;
  wire h_s_arrmul24_and6_5_y0;
  wire h_s_arrmul24_fa6_5_y2;
  wire h_s_arrmul24_fa6_5_y4;
  wire h_s_arrmul24_and7_5_y0;
  wire h_s_arrmul24_fa7_5_y2;
  wire h_s_arrmul24_fa7_5_y4;
  wire h_s_arrmul24_and8_5_y0;
  wire h_s_arrmul24_fa8_5_y2;
  wire h_s_arrmul24_fa8_5_y4;
  wire h_s_arrmul24_and9_5_y0;
  wire h_s_arrmul24_fa9_5_y2;
  wire h_s_arrmul24_fa9_5_y4;
  wire h_s_arrmul24_and10_5_y0;
  wire h_s_arrmul24_fa10_5_y2;
  wire h_s_arrmul24_fa10_5_y4;
  wire h_s_arrmul24_and11_5_y0;
  wire h_s_arrmul24_fa11_5_y2;
  wire h_s_arrmul24_fa11_5_y4;
  wire h_s_arrmul24_and12_5_y0;
  wire h_s_arrmul24_fa12_5_y2;
  wire h_s_arrmul24_fa12_5_y4;
  wire h_s_arrmul24_and13_5_y0;
  wire h_s_arrmul24_fa13_5_y2;
  wire h_s_arrmul24_fa13_5_y4;
  wire h_s_arrmul24_and14_5_y0;
  wire h_s_arrmul24_fa14_5_y2;
  wire h_s_arrmul24_fa14_5_y4;
  wire h_s_arrmul24_and15_5_y0;
  wire h_s_arrmul24_fa15_5_y2;
  wire h_s_arrmul24_fa15_5_y4;
  wire h_s_arrmul24_and16_5_y0;
  wire h_s_arrmul24_fa16_5_y2;
  wire h_s_arrmul24_fa16_5_y4;
  wire h_s_arrmul24_and17_5_y0;
  wire h_s_arrmul24_fa17_5_y2;
  wire h_s_arrmul24_fa17_5_y4;
  wire h_s_arrmul24_and18_5_y0;
  wire h_s_arrmul24_fa18_5_y2;
  wire h_s_arrmul24_fa18_5_y4;
  wire h_s_arrmul24_and19_5_y0;
  wire h_s_arrmul24_fa19_5_y2;
  wire h_s_arrmul24_fa19_5_y4;
  wire h_s_arrmul24_and20_5_y0;
  wire h_s_arrmul24_fa20_5_y2;
  wire h_s_arrmul24_fa20_5_y4;
  wire h_s_arrmul24_and21_5_y0;
  wire h_s_arrmul24_fa21_5_y2;
  wire h_s_arrmul24_fa21_5_y4;
  wire h_s_arrmul24_and22_5_y0;
  wire h_s_arrmul24_fa22_5_y2;
  wire h_s_arrmul24_fa22_5_y4;
  wire h_s_arrmul24_nand23_5_y0;
  wire h_s_arrmul24_fa23_5_y2;
  wire h_s_arrmul24_fa23_5_y4;
  wire h_s_arrmul24_and0_6_y0;
  wire h_s_arrmul24_ha0_6_y0;
  wire h_s_arrmul24_ha0_6_y1;
  wire h_s_arrmul24_and1_6_y0;
  wire h_s_arrmul24_fa1_6_y2;
  wire h_s_arrmul24_fa1_6_y4;
  wire h_s_arrmul24_and2_6_y0;
  wire h_s_arrmul24_fa2_6_y2;
  wire h_s_arrmul24_fa2_6_y4;
  wire h_s_arrmul24_and3_6_y0;
  wire h_s_arrmul24_fa3_6_y2;
  wire h_s_arrmul24_fa3_6_y4;
  wire h_s_arrmul24_and4_6_y0;
  wire h_s_arrmul24_fa4_6_y2;
  wire h_s_arrmul24_fa4_6_y4;
  wire h_s_arrmul24_and5_6_y0;
  wire h_s_arrmul24_fa5_6_y2;
  wire h_s_arrmul24_fa5_6_y4;
  wire h_s_arrmul24_and6_6_y0;
  wire h_s_arrmul24_fa6_6_y2;
  wire h_s_arrmul24_fa6_6_y4;
  wire h_s_arrmul24_and7_6_y0;
  wire h_s_arrmul24_fa7_6_y2;
  wire h_s_arrmul24_fa7_6_y4;
  wire h_s_arrmul24_and8_6_y0;
  wire h_s_arrmul24_fa8_6_y2;
  wire h_s_arrmul24_fa8_6_y4;
  wire h_s_arrmul24_and9_6_y0;
  wire h_s_arrmul24_fa9_6_y2;
  wire h_s_arrmul24_fa9_6_y4;
  wire h_s_arrmul24_and10_6_y0;
  wire h_s_arrmul24_fa10_6_y2;
  wire h_s_arrmul24_fa10_6_y4;
  wire h_s_arrmul24_and11_6_y0;
  wire h_s_arrmul24_fa11_6_y2;
  wire h_s_arrmul24_fa11_6_y4;
  wire h_s_arrmul24_and12_6_y0;
  wire h_s_arrmul24_fa12_6_y2;
  wire h_s_arrmul24_fa12_6_y4;
  wire h_s_arrmul24_and13_6_y0;
  wire h_s_arrmul24_fa13_6_y2;
  wire h_s_arrmul24_fa13_6_y4;
  wire h_s_arrmul24_and14_6_y0;
  wire h_s_arrmul24_fa14_6_y2;
  wire h_s_arrmul24_fa14_6_y4;
  wire h_s_arrmul24_and15_6_y0;
  wire h_s_arrmul24_fa15_6_y2;
  wire h_s_arrmul24_fa15_6_y4;
  wire h_s_arrmul24_and16_6_y0;
  wire h_s_arrmul24_fa16_6_y2;
  wire h_s_arrmul24_fa16_6_y4;
  wire h_s_arrmul24_and17_6_y0;
  wire h_s_arrmul24_fa17_6_y2;
  wire h_s_arrmul24_fa17_6_y4;
  wire h_s_arrmul24_and18_6_y0;
  wire h_s_arrmul24_fa18_6_y2;
  wire h_s_arrmul24_fa18_6_y4;
  wire h_s_arrmul24_and19_6_y0;
  wire h_s_arrmul24_fa19_6_y2;
  wire h_s_arrmul24_fa19_6_y4;
  wire h_s_arrmul24_and20_6_y0;
  wire h_s_arrmul24_fa20_6_y2;
  wire h_s_arrmul24_fa20_6_y4;
  wire h_s_arrmul24_and21_6_y0;
  wire h_s_arrmul24_fa21_6_y2;
  wire h_s_arrmul24_fa21_6_y4;
  wire h_s_arrmul24_and22_6_y0;
  wire h_s_arrmul24_fa22_6_y2;
  wire h_s_arrmul24_fa22_6_y4;
  wire h_s_arrmul24_nand23_6_y0;
  wire h_s_arrmul24_fa23_6_y2;
  wire h_s_arrmul24_fa23_6_y4;
  wire h_s_arrmul24_and0_7_y0;
  wire h_s_arrmul24_ha0_7_y0;
  wire h_s_arrmul24_ha0_7_y1;
  wire h_s_arrmul24_and1_7_y0;
  wire h_s_arrmul24_fa1_7_y2;
  wire h_s_arrmul24_fa1_7_y4;
  wire h_s_arrmul24_and2_7_y0;
  wire h_s_arrmul24_fa2_7_y2;
  wire h_s_arrmul24_fa2_7_y4;
  wire h_s_arrmul24_and3_7_y0;
  wire h_s_arrmul24_fa3_7_y2;
  wire h_s_arrmul24_fa3_7_y4;
  wire h_s_arrmul24_and4_7_y0;
  wire h_s_arrmul24_fa4_7_y2;
  wire h_s_arrmul24_fa4_7_y4;
  wire h_s_arrmul24_and5_7_y0;
  wire h_s_arrmul24_fa5_7_y2;
  wire h_s_arrmul24_fa5_7_y4;
  wire h_s_arrmul24_and6_7_y0;
  wire h_s_arrmul24_fa6_7_y2;
  wire h_s_arrmul24_fa6_7_y4;
  wire h_s_arrmul24_and7_7_y0;
  wire h_s_arrmul24_fa7_7_y2;
  wire h_s_arrmul24_fa7_7_y4;
  wire h_s_arrmul24_and8_7_y0;
  wire h_s_arrmul24_fa8_7_y2;
  wire h_s_arrmul24_fa8_7_y4;
  wire h_s_arrmul24_and9_7_y0;
  wire h_s_arrmul24_fa9_7_y2;
  wire h_s_arrmul24_fa9_7_y4;
  wire h_s_arrmul24_and10_7_y0;
  wire h_s_arrmul24_fa10_7_y2;
  wire h_s_arrmul24_fa10_7_y4;
  wire h_s_arrmul24_and11_7_y0;
  wire h_s_arrmul24_fa11_7_y2;
  wire h_s_arrmul24_fa11_7_y4;
  wire h_s_arrmul24_and12_7_y0;
  wire h_s_arrmul24_fa12_7_y2;
  wire h_s_arrmul24_fa12_7_y4;
  wire h_s_arrmul24_and13_7_y0;
  wire h_s_arrmul24_fa13_7_y2;
  wire h_s_arrmul24_fa13_7_y4;
  wire h_s_arrmul24_and14_7_y0;
  wire h_s_arrmul24_fa14_7_y2;
  wire h_s_arrmul24_fa14_7_y4;
  wire h_s_arrmul24_and15_7_y0;
  wire h_s_arrmul24_fa15_7_y2;
  wire h_s_arrmul24_fa15_7_y4;
  wire h_s_arrmul24_and16_7_y0;
  wire h_s_arrmul24_fa16_7_y2;
  wire h_s_arrmul24_fa16_7_y4;
  wire h_s_arrmul24_and17_7_y0;
  wire h_s_arrmul24_fa17_7_y2;
  wire h_s_arrmul24_fa17_7_y4;
  wire h_s_arrmul24_and18_7_y0;
  wire h_s_arrmul24_fa18_7_y2;
  wire h_s_arrmul24_fa18_7_y4;
  wire h_s_arrmul24_and19_7_y0;
  wire h_s_arrmul24_fa19_7_y2;
  wire h_s_arrmul24_fa19_7_y4;
  wire h_s_arrmul24_and20_7_y0;
  wire h_s_arrmul24_fa20_7_y2;
  wire h_s_arrmul24_fa20_7_y4;
  wire h_s_arrmul24_and21_7_y0;
  wire h_s_arrmul24_fa21_7_y2;
  wire h_s_arrmul24_fa21_7_y4;
  wire h_s_arrmul24_and22_7_y0;
  wire h_s_arrmul24_fa22_7_y2;
  wire h_s_arrmul24_fa22_7_y4;
  wire h_s_arrmul24_nand23_7_y0;
  wire h_s_arrmul24_fa23_7_y2;
  wire h_s_arrmul24_fa23_7_y4;
  wire h_s_arrmul24_and0_8_y0;
  wire h_s_arrmul24_ha0_8_y0;
  wire h_s_arrmul24_ha0_8_y1;
  wire h_s_arrmul24_and1_8_y0;
  wire h_s_arrmul24_fa1_8_y2;
  wire h_s_arrmul24_fa1_8_y4;
  wire h_s_arrmul24_and2_8_y0;
  wire h_s_arrmul24_fa2_8_y2;
  wire h_s_arrmul24_fa2_8_y4;
  wire h_s_arrmul24_and3_8_y0;
  wire h_s_arrmul24_fa3_8_y2;
  wire h_s_arrmul24_fa3_8_y4;
  wire h_s_arrmul24_and4_8_y0;
  wire h_s_arrmul24_fa4_8_y2;
  wire h_s_arrmul24_fa4_8_y4;
  wire h_s_arrmul24_and5_8_y0;
  wire h_s_arrmul24_fa5_8_y2;
  wire h_s_arrmul24_fa5_8_y4;
  wire h_s_arrmul24_and6_8_y0;
  wire h_s_arrmul24_fa6_8_y2;
  wire h_s_arrmul24_fa6_8_y4;
  wire h_s_arrmul24_and7_8_y0;
  wire h_s_arrmul24_fa7_8_y2;
  wire h_s_arrmul24_fa7_8_y4;
  wire h_s_arrmul24_and8_8_y0;
  wire h_s_arrmul24_fa8_8_y2;
  wire h_s_arrmul24_fa8_8_y4;
  wire h_s_arrmul24_and9_8_y0;
  wire h_s_arrmul24_fa9_8_y2;
  wire h_s_arrmul24_fa9_8_y4;
  wire h_s_arrmul24_and10_8_y0;
  wire h_s_arrmul24_fa10_8_y2;
  wire h_s_arrmul24_fa10_8_y4;
  wire h_s_arrmul24_and11_8_y0;
  wire h_s_arrmul24_fa11_8_y2;
  wire h_s_arrmul24_fa11_8_y4;
  wire h_s_arrmul24_and12_8_y0;
  wire h_s_arrmul24_fa12_8_y2;
  wire h_s_arrmul24_fa12_8_y4;
  wire h_s_arrmul24_and13_8_y0;
  wire h_s_arrmul24_fa13_8_y2;
  wire h_s_arrmul24_fa13_8_y4;
  wire h_s_arrmul24_and14_8_y0;
  wire h_s_arrmul24_fa14_8_y2;
  wire h_s_arrmul24_fa14_8_y4;
  wire h_s_arrmul24_and15_8_y0;
  wire h_s_arrmul24_fa15_8_y2;
  wire h_s_arrmul24_fa15_8_y4;
  wire h_s_arrmul24_and16_8_y0;
  wire h_s_arrmul24_fa16_8_y2;
  wire h_s_arrmul24_fa16_8_y4;
  wire h_s_arrmul24_and17_8_y0;
  wire h_s_arrmul24_fa17_8_y2;
  wire h_s_arrmul24_fa17_8_y4;
  wire h_s_arrmul24_and18_8_y0;
  wire h_s_arrmul24_fa18_8_y2;
  wire h_s_arrmul24_fa18_8_y4;
  wire h_s_arrmul24_and19_8_y0;
  wire h_s_arrmul24_fa19_8_y2;
  wire h_s_arrmul24_fa19_8_y4;
  wire h_s_arrmul24_and20_8_y0;
  wire h_s_arrmul24_fa20_8_y2;
  wire h_s_arrmul24_fa20_8_y4;
  wire h_s_arrmul24_and21_8_y0;
  wire h_s_arrmul24_fa21_8_y2;
  wire h_s_arrmul24_fa21_8_y4;
  wire h_s_arrmul24_and22_8_y0;
  wire h_s_arrmul24_fa22_8_y2;
  wire h_s_arrmul24_fa22_8_y4;
  wire h_s_arrmul24_nand23_8_y0;
  wire h_s_arrmul24_fa23_8_y2;
  wire h_s_arrmul24_fa23_8_y4;
  wire h_s_arrmul24_and0_9_y0;
  wire h_s_arrmul24_ha0_9_y0;
  wire h_s_arrmul24_ha0_9_y1;
  wire h_s_arrmul24_and1_9_y0;
  wire h_s_arrmul24_fa1_9_y2;
  wire h_s_arrmul24_fa1_9_y4;
  wire h_s_arrmul24_and2_9_y0;
  wire h_s_arrmul24_fa2_9_y2;
  wire h_s_arrmul24_fa2_9_y4;
  wire h_s_arrmul24_and3_9_y0;
  wire h_s_arrmul24_fa3_9_y2;
  wire h_s_arrmul24_fa3_9_y4;
  wire h_s_arrmul24_and4_9_y0;
  wire h_s_arrmul24_fa4_9_y2;
  wire h_s_arrmul24_fa4_9_y4;
  wire h_s_arrmul24_and5_9_y0;
  wire h_s_arrmul24_fa5_9_y2;
  wire h_s_arrmul24_fa5_9_y4;
  wire h_s_arrmul24_and6_9_y0;
  wire h_s_arrmul24_fa6_9_y2;
  wire h_s_arrmul24_fa6_9_y4;
  wire h_s_arrmul24_and7_9_y0;
  wire h_s_arrmul24_fa7_9_y2;
  wire h_s_arrmul24_fa7_9_y4;
  wire h_s_arrmul24_and8_9_y0;
  wire h_s_arrmul24_fa8_9_y2;
  wire h_s_arrmul24_fa8_9_y4;
  wire h_s_arrmul24_and9_9_y0;
  wire h_s_arrmul24_fa9_9_y2;
  wire h_s_arrmul24_fa9_9_y4;
  wire h_s_arrmul24_and10_9_y0;
  wire h_s_arrmul24_fa10_9_y2;
  wire h_s_arrmul24_fa10_9_y4;
  wire h_s_arrmul24_and11_9_y0;
  wire h_s_arrmul24_fa11_9_y2;
  wire h_s_arrmul24_fa11_9_y4;
  wire h_s_arrmul24_and12_9_y0;
  wire h_s_arrmul24_fa12_9_y2;
  wire h_s_arrmul24_fa12_9_y4;
  wire h_s_arrmul24_and13_9_y0;
  wire h_s_arrmul24_fa13_9_y2;
  wire h_s_arrmul24_fa13_9_y4;
  wire h_s_arrmul24_and14_9_y0;
  wire h_s_arrmul24_fa14_9_y2;
  wire h_s_arrmul24_fa14_9_y4;
  wire h_s_arrmul24_and15_9_y0;
  wire h_s_arrmul24_fa15_9_y2;
  wire h_s_arrmul24_fa15_9_y4;
  wire h_s_arrmul24_and16_9_y0;
  wire h_s_arrmul24_fa16_9_y2;
  wire h_s_arrmul24_fa16_9_y4;
  wire h_s_arrmul24_and17_9_y0;
  wire h_s_arrmul24_fa17_9_y2;
  wire h_s_arrmul24_fa17_9_y4;
  wire h_s_arrmul24_and18_9_y0;
  wire h_s_arrmul24_fa18_9_y2;
  wire h_s_arrmul24_fa18_9_y4;
  wire h_s_arrmul24_and19_9_y0;
  wire h_s_arrmul24_fa19_9_y2;
  wire h_s_arrmul24_fa19_9_y4;
  wire h_s_arrmul24_and20_9_y0;
  wire h_s_arrmul24_fa20_9_y2;
  wire h_s_arrmul24_fa20_9_y4;
  wire h_s_arrmul24_and21_9_y0;
  wire h_s_arrmul24_fa21_9_y2;
  wire h_s_arrmul24_fa21_9_y4;
  wire h_s_arrmul24_and22_9_y0;
  wire h_s_arrmul24_fa22_9_y2;
  wire h_s_arrmul24_fa22_9_y4;
  wire h_s_arrmul24_nand23_9_y0;
  wire h_s_arrmul24_fa23_9_y2;
  wire h_s_arrmul24_fa23_9_y4;
  wire h_s_arrmul24_and0_10_y0;
  wire h_s_arrmul24_ha0_10_y0;
  wire h_s_arrmul24_ha0_10_y1;
  wire h_s_arrmul24_and1_10_y0;
  wire h_s_arrmul24_fa1_10_y2;
  wire h_s_arrmul24_fa1_10_y4;
  wire h_s_arrmul24_and2_10_y0;
  wire h_s_arrmul24_fa2_10_y2;
  wire h_s_arrmul24_fa2_10_y4;
  wire h_s_arrmul24_and3_10_y0;
  wire h_s_arrmul24_fa3_10_y2;
  wire h_s_arrmul24_fa3_10_y4;
  wire h_s_arrmul24_and4_10_y0;
  wire h_s_arrmul24_fa4_10_y2;
  wire h_s_arrmul24_fa4_10_y4;
  wire h_s_arrmul24_and5_10_y0;
  wire h_s_arrmul24_fa5_10_y2;
  wire h_s_arrmul24_fa5_10_y4;
  wire h_s_arrmul24_and6_10_y0;
  wire h_s_arrmul24_fa6_10_y2;
  wire h_s_arrmul24_fa6_10_y4;
  wire h_s_arrmul24_and7_10_y0;
  wire h_s_arrmul24_fa7_10_y2;
  wire h_s_arrmul24_fa7_10_y4;
  wire h_s_arrmul24_and8_10_y0;
  wire h_s_arrmul24_fa8_10_y2;
  wire h_s_arrmul24_fa8_10_y4;
  wire h_s_arrmul24_and9_10_y0;
  wire h_s_arrmul24_fa9_10_y2;
  wire h_s_arrmul24_fa9_10_y4;
  wire h_s_arrmul24_and10_10_y0;
  wire h_s_arrmul24_fa10_10_y2;
  wire h_s_arrmul24_fa10_10_y4;
  wire h_s_arrmul24_and11_10_y0;
  wire h_s_arrmul24_fa11_10_y2;
  wire h_s_arrmul24_fa11_10_y4;
  wire h_s_arrmul24_and12_10_y0;
  wire h_s_arrmul24_fa12_10_y2;
  wire h_s_arrmul24_fa12_10_y4;
  wire h_s_arrmul24_and13_10_y0;
  wire h_s_arrmul24_fa13_10_y2;
  wire h_s_arrmul24_fa13_10_y4;
  wire h_s_arrmul24_and14_10_y0;
  wire h_s_arrmul24_fa14_10_y2;
  wire h_s_arrmul24_fa14_10_y4;
  wire h_s_arrmul24_and15_10_y0;
  wire h_s_arrmul24_fa15_10_y2;
  wire h_s_arrmul24_fa15_10_y4;
  wire h_s_arrmul24_and16_10_y0;
  wire h_s_arrmul24_fa16_10_y2;
  wire h_s_arrmul24_fa16_10_y4;
  wire h_s_arrmul24_and17_10_y0;
  wire h_s_arrmul24_fa17_10_y2;
  wire h_s_arrmul24_fa17_10_y4;
  wire h_s_arrmul24_and18_10_y0;
  wire h_s_arrmul24_fa18_10_y2;
  wire h_s_arrmul24_fa18_10_y4;
  wire h_s_arrmul24_and19_10_y0;
  wire h_s_arrmul24_fa19_10_y2;
  wire h_s_arrmul24_fa19_10_y4;
  wire h_s_arrmul24_and20_10_y0;
  wire h_s_arrmul24_fa20_10_y2;
  wire h_s_arrmul24_fa20_10_y4;
  wire h_s_arrmul24_and21_10_y0;
  wire h_s_arrmul24_fa21_10_y2;
  wire h_s_arrmul24_fa21_10_y4;
  wire h_s_arrmul24_and22_10_y0;
  wire h_s_arrmul24_fa22_10_y2;
  wire h_s_arrmul24_fa22_10_y4;
  wire h_s_arrmul24_nand23_10_y0;
  wire h_s_arrmul24_fa23_10_y2;
  wire h_s_arrmul24_fa23_10_y4;
  wire h_s_arrmul24_and0_11_y0;
  wire h_s_arrmul24_ha0_11_y0;
  wire h_s_arrmul24_ha0_11_y1;
  wire h_s_arrmul24_and1_11_y0;
  wire h_s_arrmul24_fa1_11_y2;
  wire h_s_arrmul24_fa1_11_y4;
  wire h_s_arrmul24_and2_11_y0;
  wire h_s_arrmul24_fa2_11_y2;
  wire h_s_arrmul24_fa2_11_y4;
  wire h_s_arrmul24_and3_11_y0;
  wire h_s_arrmul24_fa3_11_y2;
  wire h_s_arrmul24_fa3_11_y4;
  wire h_s_arrmul24_and4_11_y0;
  wire h_s_arrmul24_fa4_11_y2;
  wire h_s_arrmul24_fa4_11_y4;
  wire h_s_arrmul24_and5_11_y0;
  wire h_s_arrmul24_fa5_11_y2;
  wire h_s_arrmul24_fa5_11_y4;
  wire h_s_arrmul24_and6_11_y0;
  wire h_s_arrmul24_fa6_11_y2;
  wire h_s_arrmul24_fa6_11_y4;
  wire h_s_arrmul24_and7_11_y0;
  wire h_s_arrmul24_fa7_11_y2;
  wire h_s_arrmul24_fa7_11_y4;
  wire h_s_arrmul24_and8_11_y0;
  wire h_s_arrmul24_fa8_11_y2;
  wire h_s_arrmul24_fa8_11_y4;
  wire h_s_arrmul24_and9_11_y0;
  wire h_s_arrmul24_fa9_11_y2;
  wire h_s_arrmul24_fa9_11_y4;
  wire h_s_arrmul24_and10_11_y0;
  wire h_s_arrmul24_fa10_11_y2;
  wire h_s_arrmul24_fa10_11_y4;
  wire h_s_arrmul24_and11_11_y0;
  wire h_s_arrmul24_fa11_11_y2;
  wire h_s_arrmul24_fa11_11_y4;
  wire h_s_arrmul24_and12_11_y0;
  wire h_s_arrmul24_fa12_11_y2;
  wire h_s_arrmul24_fa12_11_y4;
  wire h_s_arrmul24_and13_11_y0;
  wire h_s_arrmul24_fa13_11_y2;
  wire h_s_arrmul24_fa13_11_y4;
  wire h_s_arrmul24_and14_11_y0;
  wire h_s_arrmul24_fa14_11_y2;
  wire h_s_arrmul24_fa14_11_y4;
  wire h_s_arrmul24_and15_11_y0;
  wire h_s_arrmul24_fa15_11_y2;
  wire h_s_arrmul24_fa15_11_y4;
  wire h_s_arrmul24_and16_11_y0;
  wire h_s_arrmul24_fa16_11_y2;
  wire h_s_arrmul24_fa16_11_y4;
  wire h_s_arrmul24_and17_11_y0;
  wire h_s_arrmul24_fa17_11_y2;
  wire h_s_arrmul24_fa17_11_y4;
  wire h_s_arrmul24_and18_11_y0;
  wire h_s_arrmul24_fa18_11_y2;
  wire h_s_arrmul24_fa18_11_y4;
  wire h_s_arrmul24_and19_11_y0;
  wire h_s_arrmul24_fa19_11_y2;
  wire h_s_arrmul24_fa19_11_y4;
  wire h_s_arrmul24_and20_11_y0;
  wire h_s_arrmul24_fa20_11_y2;
  wire h_s_arrmul24_fa20_11_y4;
  wire h_s_arrmul24_and21_11_y0;
  wire h_s_arrmul24_fa21_11_y2;
  wire h_s_arrmul24_fa21_11_y4;
  wire h_s_arrmul24_and22_11_y0;
  wire h_s_arrmul24_fa22_11_y2;
  wire h_s_arrmul24_fa22_11_y4;
  wire h_s_arrmul24_nand23_11_y0;
  wire h_s_arrmul24_fa23_11_y2;
  wire h_s_arrmul24_fa23_11_y4;
  wire h_s_arrmul24_and0_12_y0;
  wire h_s_arrmul24_ha0_12_y0;
  wire h_s_arrmul24_ha0_12_y1;
  wire h_s_arrmul24_and1_12_y0;
  wire h_s_arrmul24_fa1_12_y2;
  wire h_s_arrmul24_fa1_12_y4;
  wire h_s_arrmul24_and2_12_y0;
  wire h_s_arrmul24_fa2_12_y2;
  wire h_s_arrmul24_fa2_12_y4;
  wire h_s_arrmul24_and3_12_y0;
  wire h_s_arrmul24_fa3_12_y2;
  wire h_s_arrmul24_fa3_12_y4;
  wire h_s_arrmul24_and4_12_y0;
  wire h_s_arrmul24_fa4_12_y2;
  wire h_s_arrmul24_fa4_12_y4;
  wire h_s_arrmul24_and5_12_y0;
  wire h_s_arrmul24_fa5_12_y2;
  wire h_s_arrmul24_fa5_12_y4;
  wire h_s_arrmul24_and6_12_y0;
  wire h_s_arrmul24_fa6_12_y2;
  wire h_s_arrmul24_fa6_12_y4;
  wire h_s_arrmul24_and7_12_y0;
  wire h_s_arrmul24_fa7_12_y2;
  wire h_s_arrmul24_fa7_12_y4;
  wire h_s_arrmul24_and8_12_y0;
  wire h_s_arrmul24_fa8_12_y2;
  wire h_s_arrmul24_fa8_12_y4;
  wire h_s_arrmul24_and9_12_y0;
  wire h_s_arrmul24_fa9_12_y2;
  wire h_s_arrmul24_fa9_12_y4;
  wire h_s_arrmul24_and10_12_y0;
  wire h_s_arrmul24_fa10_12_y2;
  wire h_s_arrmul24_fa10_12_y4;
  wire h_s_arrmul24_and11_12_y0;
  wire h_s_arrmul24_fa11_12_y2;
  wire h_s_arrmul24_fa11_12_y4;
  wire h_s_arrmul24_and12_12_y0;
  wire h_s_arrmul24_fa12_12_y2;
  wire h_s_arrmul24_fa12_12_y4;
  wire h_s_arrmul24_and13_12_y0;
  wire h_s_arrmul24_fa13_12_y2;
  wire h_s_arrmul24_fa13_12_y4;
  wire h_s_arrmul24_and14_12_y0;
  wire h_s_arrmul24_fa14_12_y2;
  wire h_s_arrmul24_fa14_12_y4;
  wire h_s_arrmul24_and15_12_y0;
  wire h_s_arrmul24_fa15_12_y2;
  wire h_s_arrmul24_fa15_12_y4;
  wire h_s_arrmul24_and16_12_y0;
  wire h_s_arrmul24_fa16_12_y2;
  wire h_s_arrmul24_fa16_12_y4;
  wire h_s_arrmul24_and17_12_y0;
  wire h_s_arrmul24_fa17_12_y2;
  wire h_s_arrmul24_fa17_12_y4;
  wire h_s_arrmul24_and18_12_y0;
  wire h_s_arrmul24_fa18_12_y2;
  wire h_s_arrmul24_fa18_12_y4;
  wire h_s_arrmul24_and19_12_y0;
  wire h_s_arrmul24_fa19_12_y2;
  wire h_s_arrmul24_fa19_12_y4;
  wire h_s_arrmul24_and20_12_y0;
  wire h_s_arrmul24_fa20_12_y2;
  wire h_s_arrmul24_fa20_12_y4;
  wire h_s_arrmul24_and21_12_y0;
  wire h_s_arrmul24_fa21_12_y2;
  wire h_s_arrmul24_fa21_12_y4;
  wire h_s_arrmul24_and22_12_y0;
  wire h_s_arrmul24_fa22_12_y2;
  wire h_s_arrmul24_fa22_12_y4;
  wire h_s_arrmul24_nand23_12_y0;
  wire h_s_arrmul24_fa23_12_y2;
  wire h_s_arrmul24_fa23_12_y4;
  wire h_s_arrmul24_and0_13_y0;
  wire h_s_arrmul24_ha0_13_y0;
  wire h_s_arrmul24_ha0_13_y1;
  wire h_s_arrmul24_and1_13_y0;
  wire h_s_arrmul24_fa1_13_y2;
  wire h_s_arrmul24_fa1_13_y4;
  wire h_s_arrmul24_and2_13_y0;
  wire h_s_arrmul24_fa2_13_y2;
  wire h_s_arrmul24_fa2_13_y4;
  wire h_s_arrmul24_and3_13_y0;
  wire h_s_arrmul24_fa3_13_y2;
  wire h_s_arrmul24_fa3_13_y4;
  wire h_s_arrmul24_and4_13_y0;
  wire h_s_arrmul24_fa4_13_y2;
  wire h_s_arrmul24_fa4_13_y4;
  wire h_s_arrmul24_and5_13_y0;
  wire h_s_arrmul24_fa5_13_y2;
  wire h_s_arrmul24_fa5_13_y4;
  wire h_s_arrmul24_and6_13_y0;
  wire h_s_arrmul24_fa6_13_y2;
  wire h_s_arrmul24_fa6_13_y4;
  wire h_s_arrmul24_and7_13_y0;
  wire h_s_arrmul24_fa7_13_y2;
  wire h_s_arrmul24_fa7_13_y4;
  wire h_s_arrmul24_and8_13_y0;
  wire h_s_arrmul24_fa8_13_y2;
  wire h_s_arrmul24_fa8_13_y4;
  wire h_s_arrmul24_and9_13_y0;
  wire h_s_arrmul24_fa9_13_y2;
  wire h_s_arrmul24_fa9_13_y4;
  wire h_s_arrmul24_and10_13_y0;
  wire h_s_arrmul24_fa10_13_y2;
  wire h_s_arrmul24_fa10_13_y4;
  wire h_s_arrmul24_and11_13_y0;
  wire h_s_arrmul24_fa11_13_y2;
  wire h_s_arrmul24_fa11_13_y4;
  wire h_s_arrmul24_and12_13_y0;
  wire h_s_arrmul24_fa12_13_y2;
  wire h_s_arrmul24_fa12_13_y4;
  wire h_s_arrmul24_and13_13_y0;
  wire h_s_arrmul24_fa13_13_y2;
  wire h_s_arrmul24_fa13_13_y4;
  wire h_s_arrmul24_and14_13_y0;
  wire h_s_arrmul24_fa14_13_y2;
  wire h_s_arrmul24_fa14_13_y4;
  wire h_s_arrmul24_and15_13_y0;
  wire h_s_arrmul24_fa15_13_y2;
  wire h_s_arrmul24_fa15_13_y4;
  wire h_s_arrmul24_and16_13_y0;
  wire h_s_arrmul24_fa16_13_y2;
  wire h_s_arrmul24_fa16_13_y4;
  wire h_s_arrmul24_and17_13_y0;
  wire h_s_arrmul24_fa17_13_y2;
  wire h_s_arrmul24_fa17_13_y4;
  wire h_s_arrmul24_and18_13_y0;
  wire h_s_arrmul24_fa18_13_y2;
  wire h_s_arrmul24_fa18_13_y4;
  wire h_s_arrmul24_and19_13_y0;
  wire h_s_arrmul24_fa19_13_y2;
  wire h_s_arrmul24_fa19_13_y4;
  wire h_s_arrmul24_and20_13_y0;
  wire h_s_arrmul24_fa20_13_y2;
  wire h_s_arrmul24_fa20_13_y4;
  wire h_s_arrmul24_and21_13_y0;
  wire h_s_arrmul24_fa21_13_y2;
  wire h_s_arrmul24_fa21_13_y4;
  wire h_s_arrmul24_and22_13_y0;
  wire h_s_arrmul24_fa22_13_y2;
  wire h_s_arrmul24_fa22_13_y4;
  wire h_s_arrmul24_nand23_13_y0;
  wire h_s_arrmul24_fa23_13_y2;
  wire h_s_arrmul24_fa23_13_y4;
  wire h_s_arrmul24_and0_14_y0;
  wire h_s_arrmul24_ha0_14_y0;
  wire h_s_arrmul24_ha0_14_y1;
  wire h_s_arrmul24_and1_14_y0;
  wire h_s_arrmul24_fa1_14_y2;
  wire h_s_arrmul24_fa1_14_y4;
  wire h_s_arrmul24_and2_14_y0;
  wire h_s_arrmul24_fa2_14_y2;
  wire h_s_arrmul24_fa2_14_y4;
  wire h_s_arrmul24_and3_14_y0;
  wire h_s_arrmul24_fa3_14_y2;
  wire h_s_arrmul24_fa3_14_y4;
  wire h_s_arrmul24_and4_14_y0;
  wire h_s_arrmul24_fa4_14_y2;
  wire h_s_arrmul24_fa4_14_y4;
  wire h_s_arrmul24_and5_14_y0;
  wire h_s_arrmul24_fa5_14_y2;
  wire h_s_arrmul24_fa5_14_y4;
  wire h_s_arrmul24_and6_14_y0;
  wire h_s_arrmul24_fa6_14_y2;
  wire h_s_arrmul24_fa6_14_y4;
  wire h_s_arrmul24_and7_14_y0;
  wire h_s_arrmul24_fa7_14_y2;
  wire h_s_arrmul24_fa7_14_y4;
  wire h_s_arrmul24_and8_14_y0;
  wire h_s_arrmul24_fa8_14_y2;
  wire h_s_arrmul24_fa8_14_y4;
  wire h_s_arrmul24_and9_14_y0;
  wire h_s_arrmul24_fa9_14_y2;
  wire h_s_arrmul24_fa9_14_y4;
  wire h_s_arrmul24_and10_14_y0;
  wire h_s_arrmul24_fa10_14_y2;
  wire h_s_arrmul24_fa10_14_y4;
  wire h_s_arrmul24_and11_14_y0;
  wire h_s_arrmul24_fa11_14_y2;
  wire h_s_arrmul24_fa11_14_y4;
  wire h_s_arrmul24_and12_14_y0;
  wire h_s_arrmul24_fa12_14_y2;
  wire h_s_arrmul24_fa12_14_y4;
  wire h_s_arrmul24_and13_14_y0;
  wire h_s_arrmul24_fa13_14_y2;
  wire h_s_arrmul24_fa13_14_y4;
  wire h_s_arrmul24_and14_14_y0;
  wire h_s_arrmul24_fa14_14_y2;
  wire h_s_arrmul24_fa14_14_y4;
  wire h_s_arrmul24_and15_14_y0;
  wire h_s_arrmul24_fa15_14_y2;
  wire h_s_arrmul24_fa15_14_y4;
  wire h_s_arrmul24_and16_14_y0;
  wire h_s_arrmul24_fa16_14_y2;
  wire h_s_arrmul24_fa16_14_y4;
  wire h_s_arrmul24_and17_14_y0;
  wire h_s_arrmul24_fa17_14_y2;
  wire h_s_arrmul24_fa17_14_y4;
  wire h_s_arrmul24_and18_14_y0;
  wire h_s_arrmul24_fa18_14_y2;
  wire h_s_arrmul24_fa18_14_y4;
  wire h_s_arrmul24_and19_14_y0;
  wire h_s_arrmul24_fa19_14_y2;
  wire h_s_arrmul24_fa19_14_y4;
  wire h_s_arrmul24_and20_14_y0;
  wire h_s_arrmul24_fa20_14_y2;
  wire h_s_arrmul24_fa20_14_y4;
  wire h_s_arrmul24_and21_14_y0;
  wire h_s_arrmul24_fa21_14_y2;
  wire h_s_arrmul24_fa21_14_y4;
  wire h_s_arrmul24_and22_14_y0;
  wire h_s_arrmul24_fa22_14_y2;
  wire h_s_arrmul24_fa22_14_y4;
  wire h_s_arrmul24_nand23_14_y0;
  wire h_s_arrmul24_fa23_14_y2;
  wire h_s_arrmul24_fa23_14_y4;
  wire h_s_arrmul24_and0_15_y0;
  wire h_s_arrmul24_ha0_15_y0;
  wire h_s_arrmul24_ha0_15_y1;
  wire h_s_arrmul24_and1_15_y0;
  wire h_s_arrmul24_fa1_15_y2;
  wire h_s_arrmul24_fa1_15_y4;
  wire h_s_arrmul24_and2_15_y0;
  wire h_s_arrmul24_fa2_15_y2;
  wire h_s_arrmul24_fa2_15_y4;
  wire h_s_arrmul24_and3_15_y0;
  wire h_s_arrmul24_fa3_15_y2;
  wire h_s_arrmul24_fa3_15_y4;
  wire h_s_arrmul24_and4_15_y0;
  wire h_s_arrmul24_fa4_15_y2;
  wire h_s_arrmul24_fa4_15_y4;
  wire h_s_arrmul24_and5_15_y0;
  wire h_s_arrmul24_fa5_15_y2;
  wire h_s_arrmul24_fa5_15_y4;
  wire h_s_arrmul24_and6_15_y0;
  wire h_s_arrmul24_fa6_15_y2;
  wire h_s_arrmul24_fa6_15_y4;
  wire h_s_arrmul24_and7_15_y0;
  wire h_s_arrmul24_fa7_15_y2;
  wire h_s_arrmul24_fa7_15_y4;
  wire h_s_arrmul24_and8_15_y0;
  wire h_s_arrmul24_fa8_15_y2;
  wire h_s_arrmul24_fa8_15_y4;
  wire h_s_arrmul24_and9_15_y0;
  wire h_s_arrmul24_fa9_15_y2;
  wire h_s_arrmul24_fa9_15_y4;
  wire h_s_arrmul24_and10_15_y0;
  wire h_s_arrmul24_fa10_15_y2;
  wire h_s_arrmul24_fa10_15_y4;
  wire h_s_arrmul24_and11_15_y0;
  wire h_s_arrmul24_fa11_15_y2;
  wire h_s_arrmul24_fa11_15_y4;
  wire h_s_arrmul24_and12_15_y0;
  wire h_s_arrmul24_fa12_15_y2;
  wire h_s_arrmul24_fa12_15_y4;
  wire h_s_arrmul24_and13_15_y0;
  wire h_s_arrmul24_fa13_15_y2;
  wire h_s_arrmul24_fa13_15_y4;
  wire h_s_arrmul24_and14_15_y0;
  wire h_s_arrmul24_fa14_15_y2;
  wire h_s_arrmul24_fa14_15_y4;
  wire h_s_arrmul24_and15_15_y0;
  wire h_s_arrmul24_fa15_15_y2;
  wire h_s_arrmul24_fa15_15_y4;
  wire h_s_arrmul24_and16_15_y0;
  wire h_s_arrmul24_fa16_15_y2;
  wire h_s_arrmul24_fa16_15_y4;
  wire h_s_arrmul24_and17_15_y0;
  wire h_s_arrmul24_fa17_15_y2;
  wire h_s_arrmul24_fa17_15_y4;
  wire h_s_arrmul24_and18_15_y0;
  wire h_s_arrmul24_fa18_15_y2;
  wire h_s_arrmul24_fa18_15_y4;
  wire h_s_arrmul24_and19_15_y0;
  wire h_s_arrmul24_fa19_15_y2;
  wire h_s_arrmul24_fa19_15_y4;
  wire h_s_arrmul24_and20_15_y0;
  wire h_s_arrmul24_fa20_15_y2;
  wire h_s_arrmul24_fa20_15_y4;
  wire h_s_arrmul24_and21_15_y0;
  wire h_s_arrmul24_fa21_15_y2;
  wire h_s_arrmul24_fa21_15_y4;
  wire h_s_arrmul24_and22_15_y0;
  wire h_s_arrmul24_fa22_15_y2;
  wire h_s_arrmul24_fa22_15_y4;
  wire h_s_arrmul24_nand23_15_y0;
  wire h_s_arrmul24_fa23_15_y2;
  wire h_s_arrmul24_fa23_15_y4;
  wire h_s_arrmul24_and0_16_y0;
  wire h_s_arrmul24_ha0_16_y0;
  wire h_s_arrmul24_ha0_16_y1;
  wire h_s_arrmul24_and1_16_y0;
  wire h_s_arrmul24_fa1_16_y2;
  wire h_s_arrmul24_fa1_16_y4;
  wire h_s_arrmul24_and2_16_y0;
  wire h_s_arrmul24_fa2_16_y2;
  wire h_s_arrmul24_fa2_16_y4;
  wire h_s_arrmul24_and3_16_y0;
  wire h_s_arrmul24_fa3_16_y2;
  wire h_s_arrmul24_fa3_16_y4;
  wire h_s_arrmul24_and4_16_y0;
  wire h_s_arrmul24_fa4_16_y2;
  wire h_s_arrmul24_fa4_16_y4;
  wire h_s_arrmul24_and5_16_y0;
  wire h_s_arrmul24_fa5_16_y2;
  wire h_s_arrmul24_fa5_16_y4;
  wire h_s_arrmul24_and6_16_y0;
  wire h_s_arrmul24_fa6_16_y2;
  wire h_s_arrmul24_fa6_16_y4;
  wire h_s_arrmul24_and7_16_y0;
  wire h_s_arrmul24_fa7_16_y2;
  wire h_s_arrmul24_fa7_16_y4;
  wire h_s_arrmul24_and8_16_y0;
  wire h_s_arrmul24_fa8_16_y2;
  wire h_s_arrmul24_fa8_16_y4;
  wire h_s_arrmul24_and9_16_y0;
  wire h_s_arrmul24_fa9_16_y2;
  wire h_s_arrmul24_fa9_16_y4;
  wire h_s_arrmul24_and10_16_y0;
  wire h_s_arrmul24_fa10_16_y2;
  wire h_s_arrmul24_fa10_16_y4;
  wire h_s_arrmul24_and11_16_y0;
  wire h_s_arrmul24_fa11_16_y2;
  wire h_s_arrmul24_fa11_16_y4;
  wire h_s_arrmul24_and12_16_y0;
  wire h_s_arrmul24_fa12_16_y2;
  wire h_s_arrmul24_fa12_16_y4;
  wire h_s_arrmul24_and13_16_y0;
  wire h_s_arrmul24_fa13_16_y2;
  wire h_s_arrmul24_fa13_16_y4;
  wire h_s_arrmul24_and14_16_y0;
  wire h_s_arrmul24_fa14_16_y2;
  wire h_s_arrmul24_fa14_16_y4;
  wire h_s_arrmul24_and15_16_y0;
  wire h_s_arrmul24_fa15_16_y2;
  wire h_s_arrmul24_fa15_16_y4;
  wire h_s_arrmul24_and16_16_y0;
  wire h_s_arrmul24_fa16_16_y2;
  wire h_s_arrmul24_fa16_16_y4;
  wire h_s_arrmul24_and17_16_y0;
  wire h_s_arrmul24_fa17_16_y2;
  wire h_s_arrmul24_fa17_16_y4;
  wire h_s_arrmul24_and18_16_y0;
  wire h_s_arrmul24_fa18_16_y2;
  wire h_s_arrmul24_fa18_16_y4;
  wire h_s_arrmul24_and19_16_y0;
  wire h_s_arrmul24_fa19_16_y2;
  wire h_s_arrmul24_fa19_16_y4;
  wire h_s_arrmul24_and20_16_y0;
  wire h_s_arrmul24_fa20_16_y2;
  wire h_s_arrmul24_fa20_16_y4;
  wire h_s_arrmul24_and21_16_y0;
  wire h_s_arrmul24_fa21_16_y2;
  wire h_s_arrmul24_fa21_16_y4;
  wire h_s_arrmul24_and22_16_y0;
  wire h_s_arrmul24_fa22_16_y2;
  wire h_s_arrmul24_fa22_16_y4;
  wire h_s_arrmul24_nand23_16_y0;
  wire h_s_arrmul24_fa23_16_y2;
  wire h_s_arrmul24_fa23_16_y4;
  wire h_s_arrmul24_and0_17_y0;
  wire h_s_arrmul24_ha0_17_y0;
  wire h_s_arrmul24_ha0_17_y1;
  wire h_s_arrmul24_and1_17_y0;
  wire h_s_arrmul24_fa1_17_y2;
  wire h_s_arrmul24_fa1_17_y4;
  wire h_s_arrmul24_and2_17_y0;
  wire h_s_arrmul24_fa2_17_y2;
  wire h_s_arrmul24_fa2_17_y4;
  wire h_s_arrmul24_and3_17_y0;
  wire h_s_arrmul24_fa3_17_y2;
  wire h_s_arrmul24_fa3_17_y4;
  wire h_s_arrmul24_and4_17_y0;
  wire h_s_arrmul24_fa4_17_y2;
  wire h_s_arrmul24_fa4_17_y4;
  wire h_s_arrmul24_and5_17_y0;
  wire h_s_arrmul24_fa5_17_y2;
  wire h_s_arrmul24_fa5_17_y4;
  wire h_s_arrmul24_and6_17_y0;
  wire h_s_arrmul24_fa6_17_y2;
  wire h_s_arrmul24_fa6_17_y4;
  wire h_s_arrmul24_and7_17_y0;
  wire h_s_arrmul24_fa7_17_y2;
  wire h_s_arrmul24_fa7_17_y4;
  wire h_s_arrmul24_and8_17_y0;
  wire h_s_arrmul24_fa8_17_y2;
  wire h_s_arrmul24_fa8_17_y4;
  wire h_s_arrmul24_and9_17_y0;
  wire h_s_arrmul24_fa9_17_y2;
  wire h_s_arrmul24_fa9_17_y4;
  wire h_s_arrmul24_and10_17_y0;
  wire h_s_arrmul24_fa10_17_y2;
  wire h_s_arrmul24_fa10_17_y4;
  wire h_s_arrmul24_and11_17_y0;
  wire h_s_arrmul24_fa11_17_y2;
  wire h_s_arrmul24_fa11_17_y4;
  wire h_s_arrmul24_and12_17_y0;
  wire h_s_arrmul24_fa12_17_y2;
  wire h_s_arrmul24_fa12_17_y4;
  wire h_s_arrmul24_and13_17_y0;
  wire h_s_arrmul24_fa13_17_y2;
  wire h_s_arrmul24_fa13_17_y4;
  wire h_s_arrmul24_and14_17_y0;
  wire h_s_arrmul24_fa14_17_y2;
  wire h_s_arrmul24_fa14_17_y4;
  wire h_s_arrmul24_and15_17_y0;
  wire h_s_arrmul24_fa15_17_y2;
  wire h_s_arrmul24_fa15_17_y4;
  wire h_s_arrmul24_and16_17_y0;
  wire h_s_arrmul24_fa16_17_y2;
  wire h_s_arrmul24_fa16_17_y4;
  wire h_s_arrmul24_and17_17_y0;
  wire h_s_arrmul24_fa17_17_y2;
  wire h_s_arrmul24_fa17_17_y4;
  wire h_s_arrmul24_and18_17_y0;
  wire h_s_arrmul24_fa18_17_y2;
  wire h_s_arrmul24_fa18_17_y4;
  wire h_s_arrmul24_and19_17_y0;
  wire h_s_arrmul24_fa19_17_y2;
  wire h_s_arrmul24_fa19_17_y4;
  wire h_s_arrmul24_and20_17_y0;
  wire h_s_arrmul24_fa20_17_y2;
  wire h_s_arrmul24_fa20_17_y4;
  wire h_s_arrmul24_and21_17_y0;
  wire h_s_arrmul24_fa21_17_y2;
  wire h_s_arrmul24_fa21_17_y4;
  wire h_s_arrmul24_and22_17_y0;
  wire h_s_arrmul24_fa22_17_y2;
  wire h_s_arrmul24_fa22_17_y4;
  wire h_s_arrmul24_nand23_17_y0;
  wire h_s_arrmul24_fa23_17_y2;
  wire h_s_arrmul24_fa23_17_y4;
  wire h_s_arrmul24_and0_18_y0;
  wire h_s_arrmul24_ha0_18_y0;
  wire h_s_arrmul24_ha0_18_y1;
  wire h_s_arrmul24_and1_18_y0;
  wire h_s_arrmul24_fa1_18_y2;
  wire h_s_arrmul24_fa1_18_y4;
  wire h_s_arrmul24_and2_18_y0;
  wire h_s_arrmul24_fa2_18_y2;
  wire h_s_arrmul24_fa2_18_y4;
  wire h_s_arrmul24_and3_18_y0;
  wire h_s_arrmul24_fa3_18_y2;
  wire h_s_arrmul24_fa3_18_y4;
  wire h_s_arrmul24_and4_18_y0;
  wire h_s_arrmul24_fa4_18_y2;
  wire h_s_arrmul24_fa4_18_y4;
  wire h_s_arrmul24_and5_18_y0;
  wire h_s_arrmul24_fa5_18_y2;
  wire h_s_arrmul24_fa5_18_y4;
  wire h_s_arrmul24_and6_18_y0;
  wire h_s_arrmul24_fa6_18_y2;
  wire h_s_arrmul24_fa6_18_y4;
  wire h_s_arrmul24_and7_18_y0;
  wire h_s_arrmul24_fa7_18_y2;
  wire h_s_arrmul24_fa7_18_y4;
  wire h_s_arrmul24_and8_18_y0;
  wire h_s_arrmul24_fa8_18_y2;
  wire h_s_arrmul24_fa8_18_y4;
  wire h_s_arrmul24_and9_18_y0;
  wire h_s_arrmul24_fa9_18_y2;
  wire h_s_arrmul24_fa9_18_y4;
  wire h_s_arrmul24_and10_18_y0;
  wire h_s_arrmul24_fa10_18_y2;
  wire h_s_arrmul24_fa10_18_y4;
  wire h_s_arrmul24_and11_18_y0;
  wire h_s_arrmul24_fa11_18_y2;
  wire h_s_arrmul24_fa11_18_y4;
  wire h_s_arrmul24_and12_18_y0;
  wire h_s_arrmul24_fa12_18_y2;
  wire h_s_arrmul24_fa12_18_y4;
  wire h_s_arrmul24_and13_18_y0;
  wire h_s_arrmul24_fa13_18_y2;
  wire h_s_arrmul24_fa13_18_y4;
  wire h_s_arrmul24_and14_18_y0;
  wire h_s_arrmul24_fa14_18_y2;
  wire h_s_arrmul24_fa14_18_y4;
  wire h_s_arrmul24_and15_18_y0;
  wire h_s_arrmul24_fa15_18_y2;
  wire h_s_arrmul24_fa15_18_y4;
  wire h_s_arrmul24_and16_18_y0;
  wire h_s_arrmul24_fa16_18_y2;
  wire h_s_arrmul24_fa16_18_y4;
  wire h_s_arrmul24_and17_18_y0;
  wire h_s_arrmul24_fa17_18_y2;
  wire h_s_arrmul24_fa17_18_y4;
  wire h_s_arrmul24_and18_18_y0;
  wire h_s_arrmul24_fa18_18_y2;
  wire h_s_arrmul24_fa18_18_y4;
  wire h_s_arrmul24_and19_18_y0;
  wire h_s_arrmul24_fa19_18_y2;
  wire h_s_arrmul24_fa19_18_y4;
  wire h_s_arrmul24_and20_18_y0;
  wire h_s_arrmul24_fa20_18_y2;
  wire h_s_arrmul24_fa20_18_y4;
  wire h_s_arrmul24_and21_18_y0;
  wire h_s_arrmul24_fa21_18_y2;
  wire h_s_arrmul24_fa21_18_y4;
  wire h_s_arrmul24_and22_18_y0;
  wire h_s_arrmul24_fa22_18_y2;
  wire h_s_arrmul24_fa22_18_y4;
  wire h_s_arrmul24_nand23_18_y0;
  wire h_s_arrmul24_fa23_18_y2;
  wire h_s_arrmul24_fa23_18_y4;
  wire h_s_arrmul24_and0_19_y0;
  wire h_s_arrmul24_ha0_19_y0;
  wire h_s_arrmul24_ha0_19_y1;
  wire h_s_arrmul24_and1_19_y0;
  wire h_s_arrmul24_fa1_19_y2;
  wire h_s_arrmul24_fa1_19_y4;
  wire h_s_arrmul24_and2_19_y0;
  wire h_s_arrmul24_fa2_19_y2;
  wire h_s_arrmul24_fa2_19_y4;
  wire h_s_arrmul24_and3_19_y0;
  wire h_s_arrmul24_fa3_19_y2;
  wire h_s_arrmul24_fa3_19_y4;
  wire h_s_arrmul24_and4_19_y0;
  wire h_s_arrmul24_fa4_19_y2;
  wire h_s_arrmul24_fa4_19_y4;
  wire h_s_arrmul24_and5_19_y0;
  wire h_s_arrmul24_fa5_19_y2;
  wire h_s_arrmul24_fa5_19_y4;
  wire h_s_arrmul24_and6_19_y0;
  wire h_s_arrmul24_fa6_19_y2;
  wire h_s_arrmul24_fa6_19_y4;
  wire h_s_arrmul24_and7_19_y0;
  wire h_s_arrmul24_fa7_19_y2;
  wire h_s_arrmul24_fa7_19_y4;
  wire h_s_arrmul24_and8_19_y0;
  wire h_s_arrmul24_fa8_19_y2;
  wire h_s_arrmul24_fa8_19_y4;
  wire h_s_arrmul24_and9_19_y0;
  wire h_s_arrmul24_fa9_19_y2;
  wire h_s_arrmul24_fa9_19_y4;
  wire h_s_arrmul24_and10_19_y0;
  wire h_s_arrmul24_fa10_19_y2;
  wire h_s_arrmul24_fa10_19_y4;
  wire h_s_arrmul24_and11_19_y0;
  wire h_s_arrmul24_fa11_19_y2;
  wire h_s_arrmul24_fa11_19_y4;
  wire h_s_arrmul24_and12_19_y0;
  wire h_s_arrmul24_fa12_19_y2;
  wire h_s_arrmul24_fa12_19_y4;
  wire h_s_arrmul24_and13_19_y0;
  wire h_s_arrmul24_fa13_19_y2;
  wire h_s_arrmul24_fa13_19_y4;
  wire h_s_arrmul24_and14_19_y0;
  wire h_s_arrmul24_fa14_19_y2;
  wire h_s_arrmul24_fa14_19_y4;
  wire h_s_arrmul24_and15_19_y0;
  wire h_s_arrmul24_fa15_19_y2;
  wire h_s_arrmul24_fa15_19_y4;
  wire h_s_arrmul24_and16_19_y0;
  wire h_s_arrmul24_fa16_19_y2;
  wire h_s_arrmul24_fa16_19_y4;
  wire h_s_arrmul24_and17_19_y0;
  wire h_s_arrmul24_fa17_19_y2;
  wire h_s_arrmul24_fa17_19_y4;
  wire h_s_arrmul24_and18_19_y0;
  wire h_s_arrmul24_fa18_19_y2;
  wire h_s_arrmul24_fa18_19_y4;
  wire h_s_arrmul24_and19_19_y0;
  wire h_s_arrmul24_fa19_19_y2;
  wire h_s_arrmul24_fa19_19_y4;
  wire h_s_arrmul24_and20_19_y0;
  wire h_s_arrmul24_fa20_19_y2;
  wire h_s_arrmul24_fa20_19_y4;
  wire h_s_arrmul24_and21_19_y0;
  wire h_s_arrmul24_fa21_19_y2;
  wire h_s_arrmul24_fa21_19_y4;
  wire h_s_arrmul24_and22_19_y0;
  wire h_s_arrmul24_fa22_19_y2;
  wire h_s_arrmul24_fa22_19_y4;
  wire h_s_arrmul24_nand23_19_y0;
  wire h_s_arrmul24_fa23_19_y2;
  wire h_s_arrmul24_fa23_19_y4;
  wire h_s_arrmul24_and0_20_y0;
  wire h_s_arrmul24_ha0_20_y0;
  wire h_s_arrmul24_ha0_20_y1;
  wire h_s_arrmul24_and1_20_y0;
  wire h_s_arrmul24_fa1_20_y2;
  wire h_s_arrmul24_fa1_20_y4;
  wire h_s_arrmul24_and2_20_y0;
  wire h_s_arrmul24_fa2_20_y2;
  wire h_s_arrmul24_fa2_20_y4;
  wire h_s_arrmul24_and3_20_y0;
  wire h_s_arrmul24_fa3_20_y2;
  wire h_s_arrmul24_fa3_20_y4;
  wire h_s_arrmul24_and4_20_y0;
  wire h_s_arrmul24_fa4_20_y2;
  wire h_s_arrmul24_fa4_20_y4;
  wire h_s_arrmul24_and5_20_y0;
  wire h_s_arrmul24_fa5_20_y2;
  wire h_s_arrmul24_fa5_20_y4;
  wire h_s_arrmul24_and6_20_y0;
  wire h_s_arrmul24_fa6_20_y2;
  wire h_s_arrmul24_fa6_20_y4;
  wire h_s_arrmul24_and7_20_y0;
  wire h_s_arrmul24_fa7_20_y2;
  wire h_s_arrmul24_fa7_20_y4;
  wire h_s_arrmul24_and8_20_y0;
  wire h_s_arrmul24_fa8_20_y2;
  wire h_s_arrmul24_fa8_20_y4;
  wire h_s_arrmul24_and9_20_y0;
  wire h_s_arrmul24_fa9_20_y2;
  wire h_s_arrmul24_fa9_20_y4;
  wire h_s_arrmul24_and10_20_y0;
  wire h_s_arrmul24_fa10_20_y2;
  wire h_s_arrmul24_fa10_20_y4;
  wire h_s_arrmul24_and11_20_y0;
  wire h_s_arrmul24_fa11_20_y2;
  wire h_s_arrmul24_fa11_20_y4;
  wire h_s_arrmul24_and12_20_y0;
  wire h_s_arrmul24_fa12_20_y2;
  wire h_s_arrmul24_fa12_20_y4;
  wire h_s_arrmul24_and13_20_y0;
  wire h_s_arrmul24_fa13_20_y2;
  wire h_s_arrmul24_fa13_20_y4;
  wire h_s_arrmul24_and14_20_y0;
  wire h_s_arrmul24_fa14_20_y2;
  wire h_s_arrmul24_fa14_20_y4;
  wire h_s_arrmul24_and15_20_y0;
  wire h_s_arrmul24_fa15_20_y2;
  wire h_s_arrmul24_fa15_20_y4;
  wire h_s_arrmul24_and16_20_y0;
  wire h_s_arrmul24_fa16_20_y2;
  wire h_s_arrmul24_fa16_20_y4;
  wire h_s_arrmul24_and17_20_y0;
  wire h_s_arrmul24_fa17_20_y2;
  wire h_s_arrmul24_fa17_20_y4;
  wire h_s_arrmul24_and18_20_y0;
  wire h_s_arrmul24_fa18_20_y2;
  wire h_s_arrmul24_fa18_20_y4;
  wire h_s_arrmul24_and19_20_y0;
  wire h_s_arrmul24_fa19_20_y2;
  wire h_s_arrmul24_fa19_20_y4;
  wire h_s_arrmul24_and20_20_y0;
  wire h_s_arrmul24_fa20_20_y2;
  wire h_s_arrmul24_fa20_20_y4;
  wire h_s_arrmul24_and21_20_y0;
  wire h_s_arrmul24_fa21_20_y2;
  wire h_s_arrmul24_fa21_20_y4;
  wire h_s_arrmul24_and22_20_y0;
  wire h_s_arrmul24_fa22_20_y2;
  wire h_s_arrmul24_fa22_20_y4;
  wire h_s_arrmul24_nand23_20_y0;
  wire h_s_arrmul24_fa23_20_y2;
  wire h_s_arrmul24_fa23_20_y4;
  wire h_s_arrmul24_and0_21_y0;
  wire h_s_arrmul24_ha0_21_y0;
  wire h_s_arrmul24_ha0_21_y1;
  wire h_s_arrmul24_and1_21_y0;
  wire h_s_arrmul24_fa1_21_y2;
  wire h_s_arrmul24_fa1_21_y4;
  wire h_s_arrmul24_and2_21_y0;
  wire h_s_arrmul24_fa2_21_y2;
  wire h_s_arrmul24_fa2_21_y4;
  wire h_s_arrmul24_and3_21_y0;
  wire h_s_arrmul24_fa3_21_y2;
  wire h_s_arrmul24_fa3_21_y4;
  wire h_s_arrmul24_and4_21_y0;
  wire h_s_arrmul24_fa4_21_y2;
  wire h_s_arrmul24_fa4_21_y4;
  wire h_s_arrmul24_and5_21_y0;
  wire h_s_arrmul24_fa5_21_y2;
  wire h_s_arrmul24_fa5_21_y4;
  wire h_s_arrmul24_and6_21_y0;
  wire h_s_arrmul24_fa6_21_y2;
  wire h_s_arrmul24_fa6_21_y4;
  wire h_s_arrmul24_and7_21_y0;
  wire h_s_arrmul24_fa7_21_y2;
  wire h_s_arrmul24_fa7_21_y4;
  wire h_s_arrmul24_and8_21_y0;
  wire h_s_arrmul24_fa8_21_y2;
  wire h_s_arrmul24_fa8_21_y4;
  wire h_s_arrmul24_and9_21_y0;
  wire h_s_arrmul24_fa9_21_y2;
  wire h_s_arrmul24_fa9_21_y4;
  wire h_s_arrmul24_and10_21_y0;
  wire h_s_arrmul24_fa10_21_y2;
  wire h_s_arrmul24_fa10_21_y4;
  wire h_s_arrmul24_and11_21_y0;
  wire h_s_arrmul24_fa11_21_y2;
  wire h_s_arrmul24_fa11_21_y4;
  wire h_s_arrmul24_and12_21_y0;
  wire h_s_arrmul24_fa12_21_y2;
  wire h_s_arrmul24_fa12_21_y4;
  wire h_s_arrmul24_and13_21_y0;
  wire h_s_arrmul24_fa13_21_y2;
  wire h_s_arrmul24_fa13_21_y4;
  wire h_s_arrmul24_and14_21_y0;
  wire h_s_arrmul24_fa14_21_y2;
  wire h_s_arrmul24_fa14_21_y4;
  wire h_s_arrmul24_and15_21_y0;
  wire h_s_arrmul24_fa15_21_y2;
  wire h_s_arrmul24_fa15_21_y4;
  wire h_s_arrmul24_and16_21_y0;
  wire h_s_arrmul24_fa16_21_y2;
  wire h_s_arrmul24_fa16_21_y4;
  wire h_s_arrmul24_and17_21_y0;
  wire h_s_arrmul24_fa17_21_y2;
  wire h_s_arrmul24_fa17_21_y4;
  wire h_s_arrmul24_and18_21_y0;
  wire h_s_arrmul24_fa18_21_y2;
  wire h_s_arrmul24_fa18_21_y4;
  wire h_s_arrmul24_and19_21_y0;
  wire h_s_arrmul24_fa19_21_y2;
  wire h_s_arrmul24_fa19_21_y4;
  wire h_s_arrmul24_and20_21_y0;
  wire h_s_arrmul24_fa20_21_y2;
  wire h_s_arrmul24_fa20_21_y4;
  wire h_s_arrmul24_and21_21_y0;
  wire h_s_arrmul24_fa21_21_y2;
  wire h_s_arrmul24_fa21_21_y4;
  wire h_s_arrmul24_and22_21_y0;
  wire h_s_arrmul24_fa22_21_y2;
  wire h_s_arrmul24_fa22_21_y4;
  wire h_s_arrmul24_nand23_21_y0;
  wire h_s_arrmul24_fa23_21_y2;
  wire h_s_arrmul24_fa23_21_y4;
  wire h_s_arrmul24_and0_22_y0;
  wire h_s_arrmul24_ha0_22_y0;
  wire h_s_arrmul24_ha0_22_y1;
  wire h_s_arrmul24_and1_22_y0;
  wire h_s_arrmul24_fa1_22_y2;
  wire h_s_arrmul24_fa1_22_y4;
  wire h_s_arrmul24_and2_22_y0;
  wire h_s_arrmul24_fa2_22_y2;
  wire h_s_arrmul24_fa2_22_y4;
  wire h_s_arrmul24_and3_22_y0;
  wire h_s_arrmul24_fa3_22_y2;
  wire h_s_arrmul24_fa3_22_y4;
  wire h_s_arrmul24_and4_22_y0;
  wire h_s_arrmul24_fa4_22_y2;
  wire h_s_arrmul24_fa4_22_y4;
  wire h_s_arrmul24_and5_22_y0;
  wire h_s_arrmul24_fa5_22_y2;
  wire h_s_arrmul24_fa5_22_y4;
  wire h_s_arrmul24_and6_22_y0;
  wire h_s_arrmul24_fa6_22_y2;
  wire h_s_arrmul24_fa6_22_y4;
  wire h_s_arrmul24_and7_22_y0;
  wire h_s_arrmul24_fa7_22_y2;
  wire h_s_arrmul24_fa7_22_y4;
  wire h_s_arrmul24_and8_22_y0;
  wire h_s_arrmul24_fa8_22_y2;
  wire h_s_arrmul24_fa8_22_y4;
  wire h_s_arrmul24_and9_22_y0;
  wire h_s_arrmul24_fa9_22_y2;
  wire h_s_arrmul24_fa9_22_y4;
  wire h_s_arrmul24_and10_22_y0;
  wire h_s_arrmul24_fa10_22_y2;
  wire h_s_arrmul24_fa10_22_y4;
  wire h_s_arrmul24_and11_22_y0;
  wire h_s_arrmul24_fa11_22_y2;
  wire h_s_arrmul24_fa11_22_y4;
  wire h_s_arrmul24_and12_22_y0;
  wire h_s_arrmul24_fa12_22_y2;
  wire h_s_arrmul24_fa12_22_y4;
  wire h_s_arrmul24_and13_22_y0;
  wire h_s_arrmul24_fa13_22_y2;
  wire h_s_arrmul24_fa13_22_y4;
  wire h_s_arrmul24_and14_22_y0;
  wire h_s_arrmul24_fa14_22_y2;
  wire h_s_arrmul24_fa14_22_y4;
  wire h_s_arrmul24_and15_22_y0;
  wire h_s_arrmul24_fa15_22_y2;
  wire h_s_arrmul24_fa15_22_y4;
  wire h_s_arrmul24_and16_22_y0;
  wire h_s_arrmul24_fa16_22_y2;
  wire h_s_arrmul24_fa16_22_y4;
  wire h_s_arrmul24_and17_22_y0;
  wire h_s_arrmul24_fa17_22_y2;
  wire h_s_arrmul24_fa17_22_y4;
  wire h_s_arrmul24_and18_22_y0;
  wire h_s_arrmul24_fa18_22_y2;
  wire h_s_arrmul24_fa18_22_y4;
  wire h_s_arrmul24_and19_22_y0;
  wire h_s_arrmul24_fa19_22_y2;
  wire h_s_arrmul24_fa19_22_y4;
  wire h_s_arrmul24_and20_22_y0;
  wire h_s_arrmul24_fa20_22_y2;
  wire h_s_arrmul24_fa20_22_y4;
  wire h_s_arrmul24_and21_22_y0;
  wire h_s_arrmul24_fa21_22_y2;
  wire h_s_arrmul24_fa21_22_y4;
  wire h_s_arrmul24_and22_22_y0;
  wire h_s_arrmul24_fa22_22_y2;
  wire h_s_arrmul24_fa22_22_y4;
  wire h_s_arrmul24_nand23_22_y0;
  wire h_s_arrmul24_fa23_22_y2;
  wire h_s_arrmul24_fa23_22_y4;
  wire h_s_arrmul24_nand0_23_y0;
  wire h_s_arrmul24_ha0_23_y0;
  wire h_s_arrmul24_ha0_23_y1;
  wire h_s_arrmul24_nand1_23_y0;
  wire h_s_arrmul24_fa1_23_y2;
  wire h_s_arrmul24_fa1_23_y4;
  wire h_s_arrmul24_nand2_23_y0;
  wire h_s_arrmul24_fa2_23_y2;
  wire h_s_arrmul24_fa2_23_y4;
  wire h_s_arrmul24_nand3_23_y0;
  wire h_s_arrmul24_fa3_23_y2;
  wire h_s_arrmul24_fa3_23_y4;
  wire h_s_arrmul24_nand4_23_y0;
  wire h_s_arrmul24_fa4_23_y2;
  wire h_s_arrmul24_fa4_23_y4;
  wire h_s_arrmul24_nand5_23_y0;
  wire h_s_arrmul24_fa5_23_y2;
  wire h_s_arrmul24_fa5_23_y4;
  wire h_s_arrmul24_nand6_23_y0;
  wire h_s_arrmul24_fa6_23_y2;
  wire h_s_arrmul24_fa6_23_y4;
  wire h_s_arrmul24_nand7_23_y0;
  wire h_s_arrmul24_fa7_23_y2;
  wire h_s_arrmul24_fa7_23_y4;
  wire h_s_arrmul24_nand8_23_y0;
  wire h_s_arrmul24_fa8_23_y2;
  wire h_s_arrmul24_fa8_23_y4;
  wire h_s_arrmul24_nand9_23_y0;
  wire h_s_arrmul24_fa9_23_y2;
  wire h_s_arrmul24_fa9_23_y4;
  wire h_s_arrmul24_nand10_23_y0;
  wire h_s_arrmul24_fa10_23_y2;
  wire h_s_arrmul24_fa10_23_y4;
  wire h_s_arrmul24_nand11_23_y0;
  wire h_s_arrmul24_fa11_23_y2;
  wire h_s_arrmul24_fa11_23_y4;
  wire h_s_arrmul24_nand12_23_y0;
  wire h_s_arrmul24_fa12_23_y2;
  wire h_s_arrmul24_fa12_23_y4;
  wire h_s_arrmul24_nand13_23_y0;
  wire h_s_arrmul24_fa13_23_y2;
  wire h_s_arrmul24_fa13_23_y4;
  wire h_s_arrmul24_nand14_23_y0;
  wire h_s_arrmul24_fa14_23_y2;
  wire h_s_arrmul24_fa14_23_y4;
  wire h_s_arrmul24_nand15_23_y0;
  wire h_s_arrmul24_fa15_23_y2;
  wire h_s_arrmul24_fa15_23_y4;
  wire h_s_arrmul24_nand16_23_y0;
  wire h_s_arrmul24_fa16_23_y2;
  wire h_s_arrmul24_fa16_23_y4;
  wire h_s_arrmul24_nand17_23_y0;
  wire h_s_arrmul24_fa17_23_y2;
  wire h_s_arrmul24_fa17_23_y4;
  wire h_s_arrmul24_nand18_23_y0;
  wire h_s_arrmul24_fa18_23_y2;
  wire h_s_arrmul24_fa18_23_y4;
  wire h_s_arrmul24_nand19_23_y0;
  wire h_s_arrmul24_fa19_23_y2;
  wire h_s_arrmul24_fa19_23_y4;
  wire h_s_arrmul24_nand20_23_y0;
  wire h_s_arrmul24_fa20_23_y2;
  wire h_s_arrmul24_fa20_23_y4;
  wire h_s_arrmul24_nand21_23_y0;
  wire h_s_arrmul24_fa21_23_y2;
  wire h_s_arrmul24_fa21_23_y4;
  wire h_s_arrmul24_nand22_23_y0;
  wire h_s_arrmul24_fa22_23_y2;
  wire h_s_arrmul24_fa22_23_y4;
  wire h_s_arrmul24_and23_23_y0;
  wire h_s_arrmul24_fa23_23_y2;
  wire h_s_arrmul24_fa23_23_y4;
  wire h_s_arrmul24_xor24_23_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  constant_wire_value_1 constant_wire_value_1_constant_wire_1(a_0, b_0, constant_wire_1);
  and_gate and_gate_h_s_arrmul24_and0_0_y0(a_0, b_0, h_s_arrmul24_and0_0_y0);
  and_gate and_gate_h_s_arrmul24_and1_0_y0(a_1, b_0, h_s_arrmul24_and1_0_y0);
  and_gate and_gate_h_s_arrmul24_and2_0_y0(a_2, b_0, h_s_arrmul24_and2_0_y0);
  and_gate and_gate_h_s_arrmul24_and3_0_y0(a_3, b_0, h_s_arrmul24_and3_0_y0);
  and_gate and_gate_h_s_arrmul24_and4_0_y0(a_4, b_0, h_s_arrmul24_and4_0_y0);
  and_gate and_gate_h_s_arrmul24_and5_0_y0(a_5, b_0, h_s_arrmul24_and5_0_y0);
  and_gate and_gate_h_s_arrmul24_and6_0_y0(a_6, b_0, h_s_arrmul24_and6_0_y0);
  and_gate and_gate_h_s_arrmul24_and7_0_y0(a_7, b_0, h_s_arrmul24_and7_0_y0);
  and_gate and_gate_h_s_arrmul24_and8_0_y0(a_8, b_0, h_s_arrmul24_and8_0_y0);
  and_gate and_gate_h_s_arrmul24_and9_0_y0(a_9, b_0, h_s_arrmul24_and9_0_y0);
  and_gate and_gate_h_s_arrmul24_and10_0_y0(a_10, b_0, h_s_arrmul24_and10_0_y0);
  and_gate and_gate_h_s_arrmul24_and11_0_y0(a_11, b_0, h_s_arrmul24_and11_0_y0);
  and_gate and_gate_h_s_arrmul24_and12_0_y0(a_12, b_0, h_s_arrmul24_and12_0_y0);
  and_gate and_gate_h_s_arrmul24_and13_0_y0(a_13, b_0, h_s_arrmul24_and13_0_y0);
  and_gate and_gate_h_s_arrmul24_and14_0_y0(a_14, b_0, h_s_arrmul24_and14_0_y0);
  and_gate and_gate_h_s_arrmul24_and15_0_y0(a_15, b_0, h_s_arrmul24_and15_0_y0);
  and_gate and_gate_h_s_arrmul24_and16_0_y0(a_16, b_0, h_s_arrmul24_and16_0_y0);
  and_gate and_gate_h_s_arrmul24_and17_0_y0(a_17, b_0, h_s_arrmul24_and17_0_y0);
  and_gate and_gate_h_s_arrmul24_and18_0_y0(a_18, b_0, h_s_arrmul24_and18_0_y0);
  and_gate and_gate_h_s_arrmul24_and19_0_y0(a_19, b_0, h_s_arrmul24_and19_0_y0);
  and_gate and_gate_h_s_arrmul24_and20_0_y0(a_20, b_0, h_s_arrmul24_and20_0_y0);
  and_gate and_gate_h_s_arrmul24_and21_0_y0(a_21, b_0, h_s_arrmul24_and21_0_y0);
  and_gate and_gate_h_s_arrmul24_and22_0_y0(a_22, b_0, h_s_arrmul24_and22_0_y0);
  nand_gate nand_gate_h_s_arrmul24_nand23_0_y0(a_23, b_0, h_s_arrmul24_nand23_0_y0);
  and_gate and_gate_h_s_arrmul24_and0_1_y0(a_0, b_1, h_s_arrmul24_and0_1_y0);
  ha ha_h_s_arrmul24_ha0_1_y0(h_s_arrmul24_and0_1_y0, h_s_arrmul24_and1_0_y0, h_s_arrmul24_ha0_1_y0, h_s_arrmul24_ha0_1_y1);
  and_gate and_gate_h_s_arrmul24_and1_1_y0(a_1, b_1, h_s_arrmul24_and1_1_y0);
  fa fa_h_s_arrmul24_fa1_1_y2(h_s_arrmul24_and1_1_y0, h_s_arrmul24_and2_0_y0, h_s_arrmul24_ha0_1_y1, h_s_arrmul24_fa1_1_y2, h_s_arrmul24_fa1_1_y4);
  and_gate and_gate_h_s_arrmul24_and2_1_y0(a_2, b_1, h_s_arrmul24_and2_1_y0);
  fa fa_h_s_arrmul24_fa2_1_y2(h_s_arrmul24_and2_1_y0, h_s_arrmul24_and3_0_y0, h_s_arrmul24_fa1_1_y4, h_s_arrmul24_fa2_1_y2, h_s_arrmul24_fa2_1_y4);
  and_gate and_gate_h_s_arrmul24_and3_1_y0(a_3, b_1, h_s_arrmul24_and3_1_y0);
  fa fa_h_s_arrmul24_fa3_1_y2(h_s_arrmul24_and3_1_y0, h_s_arrmul24_and4_0_y0, h_s_arrmul24_fa2_1_y4, h_s_arrmul24_fa3_1_y2, h_s_arrmul24_fa3_1_y4);
  and_gate and_gate_h_s_arrmul24_and4_1_y0(a_4, b_1, h_s_arrmul24_and4_1_y0);
  fa fa_h_s_arrmul24_fa4_1_y2(h_s_arrmul24_and4_1_y0, h_s_arrmul24_and5_0_y0, h_s_arrmul24_fa3_1_y4, h_s_arrmul24_fa4_1_y2, h_s_arrmul24_fa4_1_y4);
  and_gate and_gate_h_s_arrmul24_and5_1_y0(a_5, b_1, h_s_arrmul24_and5_1_y0);
  fa fa_h_s_arrmul24_fa5_1_y2(h_s_arrmul24_and5_1_y0, h_s_arrmul24_and6_0_y0, h_s_arrmul24_fa4_1_y4, h_s_arrmul24_fa5_1_y2, h_s_arrmul24_fa5_1_y4);
  and_gate and_gate_h_s_arrmul24_and6_1_y0(a_6, b_1, h_s_arrmul24_and6_1_y0);
  fa fa_h_s_arrmul24_fa6_1_y2(h_s_arrmul24_and6_1_y0, h_s_arrmul24_and7_0_y0, h_s_arrmul24_fa5_1_y4, h_s_arrmul24_fa6_1_y2, h_s_arrmul24_fa6_1_y4);
  and_gate and_gate_h_s_arrmul24_and7_1_y0(a_7, b_1, h_s_arrmul24_and7_1_y0);
  fa fa_h_s_arrmul24_fa7_1_y2(h_s_arrmul24_and7_1_y0, h_s_arrmul24_and8_0_y0, h_s_arrmul24_fa6_1_y4, h_s_arrmul24_fa7_1_y2, h_s_arrmul24_fa7_1_y4);
  and_gate and_gate_h_s_arrmul24_and8_1_y0(a_8, b_1, h_s_arrmul24_and8_1_y0);
  fa fa_h_s_arrmul24_fa8_1_y2(h_s_arrmul24_and8_1_y0, h_s_arrmul24_and9_0_y0, h_s_arrmul24_fa7_1_y4, h_s_arrmul24_fa8_1_y2, h_s_arrmul24_fa8_1_y4);
  and_gate and_gate_h_s_arrmul24_and9_1_y0(a_9, b_1, h_s_arrmul24_and9_1_y0);
  fa fa_h_s_arrmul24_fa9_1_y2(h_s_arrmul24_and9_1_y0, h_s_arrmul24_and10_0_y0, h_s_arrmul24_fa8_1_y4, h_s_arrmul24_fa9_1_y2, h_s_arrmul24_fa9_1_y4);
  and_gate and_gate_h_s_arrmul24_and10_1_y0(a_10, b_1, h_s_arrmul24_and10_1_y0);
  fa fa_h_s_arrmul24_fa10_1_y2(h_s_arrmul24_and10_1_y0, h_s_arrmul24_and11_0_y0, h_s_arrmul24_fa9_1_y4, h_s_arrmul24_fa10_1_y2, h_s_arrmul24_fa10_1_y4);
  and_gate and_gate_h_s_arrmul24_and11_1_y0(a_11, b_1, h_s_arrmul24_and11_1_y0);
  fa fa_h_s_arrmul24_fa11_1_y2(h_s_arrmul24_and11_1_y0, h_s_arrmul24_and12_0_y0, h_s_arrmul24_fa10_1_y4, h_s_arrmul24_fa11_1_y2, h_s_arrmul24_fa11_1_y4);
  and_gate and_gate_h_s_arrmul24_and12_1_y0(a_12, b_1, h_s_arrmul24_and12_1_y0);
  fa fa_h_s_arrmul24_fa12_1_y2(h_s_arrmul24_and12_1_y0, h_s_arrmul24_and13_0_y0, h_s_arrmul24_fa11_1_y4, h_s_arrmul24_fa12_1_y2, h_s_arrmul24_fa12_1_y4);
  and_gate and_gate_h_s_arrmul24_and13_1_y0(a_13, b_1, h_s_arrmul24_and13_1_y0);
  fa fa_h_s_arrmul24_fa13_1_y2(h_s_arrmul24_and13_1_y0, h_s_arrmul24_and14_0_y0, h_s_arrmul24_fa12_1_y4, h_s_arrmul24_fa13_1_y2, h_s_arrmul24_fa13_1_y4);
  and_gate and_gate_h_s_arrmul24_and14_1_y0(a_14, b_1, h_s_arrmul24_and14_1_y0);
  fa fa_h_s_arrmul24_fa14_1_y2(h_s_arrmul24_and14_1_y0, h_s_arrmul24_and15_0_y0, h_s_arrmul24_fa13_1_y4, h_s_arrmul24_fa14_1_y2, h_s_arrmul24_fa14_1_y4);
  and_gate and_gate_h_s_arrmul24_and15_1_y0(a_15, b_1, h_s_arrmul24_and15_1_y0);
  fa fa_h_s_arrmul24_fa15_1_y2(h_s_arrmul24_and15_1_y0, h_s_arrmul24_and16_0_y0, h_s_arrmul24_fa14_1_y4, h_s_arrmul24_fa15_1_y2, h_s_arrmul24_fa15_1_y4);
  and_gate and_gate_h_s_arrmul24_and16_1_y0(a_16, b_1, h_s_arrmul24_and16_1_y0);
  fa fa_h_s_arrmul24_fa16_1_y2(h_s_arrmul24_and16_1_y0, h_s_arrmul24_and17_0_y0, h_s_arrmul24_fa15_1_y4, h_s_arrmul24_fa16_1_y2, h_s_arrmul24_fa16_1_y4);
  and_gate and_gate_h_s_arrmul24_and17_1_y0(a_17, b_1, h_s_arrmul24_and17_1_y0);
  fa fa_h_s_arrmul24_fa17_1_y2(h_s_arrmul24_and17_1_y0, h_s_arrmul24_and18_0_y0, h_s_arrmul24_fa16_1_y4, h_s_arrmul24_fa17_1_y2, h_s_arrmul24_fa17_1_y4);
  and_gate and_gate_h_s_arrmul24_and18_1_y0(a_18, b_1, h_s_arrmul24_and18_1_y0);
  fa fa_h_s_arrmul24_fa18_1_y2(h_s_arrmul24_and18_1_y0, h_s_arrmul24_and19_0_y0, h_s_arrmul24_fa17_1_y4, h_s_arrmul24_fa18_1_y2, h_s_arrmul24_fa18_1_y4);
  and_gate and_gate_h_s_arrmul24_and19_1_y0(a_19, b_1, h_s_arrmul24_and19_1_y0);
  fa fa_h_s_arrmul24_fa19_1_y2(h_s_arrmul24_and19_1_y0, h_s_arrmul24_and20_0_y0, h_s_arrmul24_fa18_1_y4, h_s_arrmul24_fa19_1_y2, h_s_arrmul24_fa19_1_y4);
  and_gate and_gate_h_s_arrmul24_and20_1_y0(a_20, b_1, h_s_arrmul24_and20_1_y0);
  fa fa_h_s_arrmul24_fa20_1_y2(h_s_arrmul24_and20_1_y0, h_s_arrmul24_and21_0_y0, h_s_arrmul24_fa19_1_y4, h_s_arrmul24_fa20_1_y2, h_s_arrmul24_fa20_1_y4);
  and_gate and_gate_h_s_arrmul24_and21_1_y0(a_21, b_1, h_s_arrmul24_and21_1_y0);
  fa fa_h_s_arrmul24_fa21_1_y2(h_s_arrmul24_and21_1_y0, h_s_arrmul24_and22_0_y0, h_s_arrmul24_fa20_1_y4, h_s_arrmul24_fa21_1_y2, h_s_arrmul24_fa21_1_y4);
  and_gate and_gate_h_s_arrmul24_and22_1_y0(a_22, b_1, h_s_arrmul24_and22_1_y0);
  fa fa_h_s_arrmul24_fa22_1_y2(h_s_arrmul24_and22_1_y0, h_s_arrmul24_nand23_0_y0, h_s_arrmul24_fa21_1_y4, h_s_arrmul24_fa22_1_y2, h_s_arrmul24_fa22_1_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_1_y0(a_23, b_1, h_s_arrmul24_nand23_1_y0);
  fa fa_h_s_arrmul24_fa23_1_y2(h_s_arrmul24_nand23_1_y0, constant_wire_1, h_s_arrmul24_fa22_1_y4, h_s_arrmul24_fa23_1_y2, h_s_arrmul24_fa23_1_y4);
  and_gate and_gate_h_s_arrmul24_and0_2_y0(a_0, b_2, h_s_arrmul24_and0_2_y0);
  ha ha_h_s_arrmul24_ha0_2_y0(h_s_arrmul24_and0_2_y0, h_s_arrmul24_fa1_1_y2, h_s_arrmul24_ha0_2_y0, h_s_arrmul24_ha0_2_y1);
  and_gate and_gate_h_s_arrmul24_and1_2_y0(a_1, b_2, h_s_arrmul24_and1_2_y0);
  fa fa_h_s_arrmul24_fa1_2_y2(h_s_arrmul24_and1_2_y0, h_s_arrmul24_fa2_1_y2, h_s_arrmul24_ha0_2_y1, h_s_arrmul24_fa1_2_y2, h_s_arrmul24_fa1_2_y4);
  and_gate and_gate_h_s_arrmul24_and2_2_y0(a_2, b_2, h_s_arrmul24_and2_2_y0);
  fa fa_h_s_arrmul24_fa2_2_y2(h_s_arrmul24_and2_2_y0, h_s_arrmul24_fa3_1_y2, h_s_arrmul24_fa1_2_y4, h_s_arrmul24_fa2_2_y2, h_s_arrmul24_fa2_2_y4);
  and_gate and_gate_h_s_arrmul24_and3_2_y0(a_3, b_2, h_s_arrmul24_and3_2_y0);
  fa fa_h_s_arrmul24_fa3_2_y2(h_s_arrmul24_and3_2_y0, h_s_arrmul24_fa4_1_y2, h_s_arrmul24_fa2_2_y4, h_s_arrmul24_fa3_2_y2, h_s_arrmul24_fa3_2_y4);
  and_gate and_gate_h_s_arrmul24_and4_2_y0(a_4, b_2, h_s_arrmul24_and4_2_y0);
  fa fa_h_s_arrmul24_fa4_2_y2(h_s_arrmul24_and4_2_y0, h_s_arrmul24_fa5_1_y2, h_s_arrmul24_fa3_2_y4, h_s_arrmul24_fa4_2_y2, h_s_arrmul24_fa4_2_y4);
  and_gate and_gate_h_s_arrmul24_and5_2_y0(a_5, b_2, h_s_arrmul24_and5_2_y0);
  fa fa_h_s_arrmul24_fa5_2_y2(h_s_arrmul24_and5_2_y0, h_s_arrmul24_fa6_1_y2, h_s_arrmul24_fa4_2_y4, h_s_arrmul24_fa5_2_y2, h_s_arrmul24_fa5_2_y4);
  and_gate and_gate_h_s_arrmul24_and6_2_y0(a_6, b_2, h_s_arrmul24_and6_2_y0);
  fa fa_h_s_arrmul24_fa6_2_y2(h_s_arrmul24_and6_2_y0, h_s_arrmul24_fa7_1_y2, h_s_arrmul24_fa5_2_y4, h_s_arrmul24_fa6_2_y2, h_s_arrmul24_fa6_2_y4);
  and_gate and_gate_h_s_arrmul24_and7_2_y0(a_7, b_2, h_s_arrmul24_and7_2_y0);
  fa fa_h_s_arrmul24_fa7_2_y2(h_s_arrmul24_and7_2_y0, h_s_arrmul24_fa8_1_y2, h_s_arrmul24_fa6_2_y4, h_s_arrmul24_fa7_2_y2, h_s_arrmul24_fa7_2_y4);
  and_gate and_gate_h_s_arrmul24_and8_2_y0(a_8, b_2, h_s_arrmul24_and8_2_y0);
  fa fa_h_s_arrmul24_fa8_2_y2(h_s_arrmul24_and8_2_y0, h_s_arrmul24_fa9_1_y2, h_s_arrmul24_fa7_2_y4, h_s_arrmul24_fa8_2_y2, h_s_arrmul24_fa8_2_y4);
  and_gate and_gate_h_s_arrmul24_and9_2_y0(a_9, b_2, h_s_arrmul24_and9_2_y0);
  fa fa_h_s_arrmul24_fa9_2_y2(h_s_arrmul24_and9_2_y0, h_s_arrmul24_fa10_1_y2, h_s_arrmul24_fa8_2_y4, h_s_arrmul24_fa9_2_y2, h_s_arrmul24_fa9_2_y4);
  and_gate and_gate_h_s_arrmul24_and10_2_y0(a_10, b_2, h_s_arrmul24_and10_2_y0);
  fa fa_h_s_arrmul24_fa10_2_y2(h_s_arrmul24_and10_2_y0, h_s_arrmul24_fa11_1_y2, h_s_arrmul24_fa9_2_y4, h_s_arrmul24_fa10_2_y2, h_s_arrmul24_fa10_2_y4);
  and_gate and_gate_h_s_arrmul24_and11_2_y0(a_11, b_2, h_s_arrmul24_and11_2_y0);
  fa fa_h_s_arrmul24_fa11_2_y2(h_s_arrmul24_and11_2_y0, h_s_arrmul24_fa12_1_y2, h_s_arrmul24_fa10_2_y4, h_s_arrmul24_fa11_2_y2, h_s_arrmul24_fa11_2_y4);
  and_gate and_gate_h_s_arrmul24_and12_2_y0(a_12, b_2, h_s_arrmul24_and12_2_y0);
  fa fa_h_s_arrmul24_fa12_2_y2(h_s_arrmul24_and12_2_y0, h_s_arrmul24_fa13_1_y2, h_s_arrmul24_fa11_2_y4, h_s_arrmul24_fa12_2_y2, h_s_arrmul24_fa12_2_y4);
  and_gate and_gate_h_s_arrmul24_and13_2_y0(a_13, b_2, h_s_arrmul24_and13_2_y0);
  fa fa_h_s_arrmul24_fa13_2_y2(h_s_arrmul24_and13_2_y0, h_s_arrmul24_fa14_1_y2, h_s_arrmul24_fa12_2_y4, h_s_arrmul24_fa13_2_y2, h_s_arrmul24_fa13_2_y4);
  and_gate and_gate_h_s_arrmul24_and14_2_y0(a_14, b_2, h_s_arrmul24_and14_2_y0);
  fa fa_h_s_arrmul24_fa14_2_y2(h_s_arrmul24_and14_2_y0, h_s_arrmul24_fa15_1_y2, h_s_arrmul24_fa13_2_y4, h_s_arrmul24_fa14_2_y2, h_s_arrmul24_fa14_2_y4);
  and_gate and_gate_h_s_arrmul24_and15_2_y0(a_15, b_2, h_s_arrmul24_and15_2_y0);
  fa fa_h_s_arrmul24_fa15_2_y2(h_s_arrmul24_and15_2_y0, h_s_arrmul24_fa16_1_y2, h_s_arrmul24_fa14_2_y4, h_s_arrmul24_fa15_2_y2, h_s_arrmul24_fa15_2_y4);
  and_gate and_gate_h_s_arrmul24_and16_2_y0(a_16, b_2, h_s_arrmul24_and16_2_y0);
  fa fa_h_s_arrmul24_fa16_2_y2(h_s_arrmul24_and16_2_y0, h_s_arrmul24_fa17_1_y2, h_s_arrmul24_fa15_2_y4, h_s_arrmul24_fa16_2_y2, h_s_arrmul24_fa16_2_y4);
  and_gate and_gate_h_s_arrmul24_and17_2_y0(a_17, b_2, h_s_arrmul24_and17_2_y0);
  fa fa_h_s_arrmul24_fa17_2_y2(h_s_arrmul24_and17_2_y0, h_s_arrmul24_fa18_1_y2, h_s_arrmul24_fa16_2_y4, h_s_arrmul24_fa17_2_y2, h_s_arrmul24_fa17_2_y4);
  and_gate and_gate_h_s_arrmul24_and18_2_y0(a_18, b_2, h_s_arrmul24_and18_2_y0);
  fa fa_h_s_arrmul24_fa18_2_y2(h_s_arrmul24_and18_2_y0, h_s_arrmul24_fa19_1_y2, h_s_arrmul24_fa17_2_y4, h_s_arrmul24_fa18_2_y2, h_s_arrmul24_fa18_2_y4);
  and_gate and_gate_h_s_arrmul24_and19_2_y0(a_19, b_2, h_s_arrmul24_and19_2_y0);
  fa fa_h_s_arrmul24_fa19_2_y2(h_s_arrmul24_and19_2_y0, h_s_arrmul24_fa20_1_y2, h_s_arrmul24_fa18_2_y4, h_s_arrmul24_fa19_2_y2, h_s_arrmul24_fa19_2_y4);
  and_gate and_gate_h_s_arrmul24_and20_2_y0(a_20, b_2, h_s_arrmul24_and20_2_y0);
  fa fa_h_s_arrmul24_fa20_2_y2(h_s_arrmul24_and20_2_y0, h_s_arrmul24_fa21_1_y2, h_s_arrmul24_fa19_2_y4, h_s_arrmul24_fa20_2_y2, h_s_arrmul24_fa20_2_y4);
  and_gate and_gate_h_s_arrmul24_and21_2_y0(a_21, b_2, h_s_arrmul24_and21_2_y0);
  fa fa_h_s_arrmul24_fa21_2_y2(h_s_arrmul24_and21_2_y0, h_s_arrmul24_fa22_1_y2, h_s_arrmul24_fa20_2_y4, h_s_arrmul24_fa21_2_y2, h_s_arrmul24_fa21_2_y4);
  and_gate and_gate_h_s_arrmul24_and22_2_y0(a_22, b_2, h_s_arrmul24_and22_2_y0);
  fa fa_h_s_arrmul24_fa22_2_y2(h_s_arrmul24_and22_2_y0, h_s_arrmul24_fa23_1_y2, h_s_arrmul24_fa21_2_y4, h_s_arrmul24_fa22_2_y2, h_s_arrmul24_fa22_2_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_2_y0(a_23, b_2, h_s_arrmul24_nand23_2_y0);
  fa fa_h_s_arrmul24_fa23_2_y2(h_s_arrmul24_nand23_2_y0, h_s_arrmul24_fa23_1_y4, h_s_arrmul24_fa22_2_y4, h_s_arrmul24_fa23_2_y2, h_s_arrmul24_fa23_2_y4);
  and_gate and_gate_h_s_arrmul24_and0_3_y0(a_0, b_3, h_s_arrmul24_and0_3_y0);
  ha ha_h_s_arrmul24_ha0_3_y0(h_s_arrmul24_and0_3_y0, h_s_arrmul24_fa1_2_y2, h_s_arrmul24_ha0_3_y0, h_s_arrmul24_ha0_3_y1);
  and_gate and_gate_h_s_arrmul24_and1_3_y0(a_1, b_3, h_s_arrmul24_and1_3_y0);
  fa fa_h_s_arrmul24_fa1_3_y2(h_s_arrmul24_and1_3_y0, h_s_arrmul24_fa2_2_y2, h_s_arrmul24_ha0_3_y1, h_s_arrmul24_fa1_3_y2, h_s_arrmul24_fa1_3_y4);
  and_gate and_gate_h_s_arrmul24_and2_3_y0(a_2, b_3, h_s_arrmul24_and2_3_y0);
  fa fa_h_s_arrmul24_fa2_3_y2(h_s_arrmul24_and2_3_y0, h_s_arrmul24_fa3_2_y2, h_s_arrmul24_fa1_3_y4, h_s_arrmul24_fa2_3_y2, h_s_arrmul24_fa2_3_y4);
  and_gate and_gate_h_s_arrmul24_and3_3_y0(a_3, b_3, h_s_arrmul24_and3_3_y0);
  fa fa_h_s_arrmul24_fa3_3_y2(h_s_arrmul24_and3_3_y0, h_s_arrmul24_fa4_2_y2, h_s_arrmul24_fa2_3_y4, h_s_arrmul24_fa3_3_y2, h_s_arrmul24_fa3_3_y4);
  and_gate and_gate_h_s_arrmul24_and4_3_y0(a_4, b_3, h_s_arrmul24_and4_3_y0);
  fa fa_h_s_arrmul24_fa4_3_y2(h_s_arrmul24_and4_3_y0, h_s_arrmul24_fa5_2_y2, h_s_arrmul24_fa3_3_y4, h_s_arrmul24_fa4_3_y2, h_s_arrmul24_fa4_3_y4);
  and_gate and_gate_h_s_arrmul24_and5_3_y0(a_5, b_3, h_s_arrmul24_and5_3_y0);
  fa fa_h_s_arrmul24_fa5_3_y2(h_s_arrmul24_and5_3_y0, h_s_arrmul24_fa6_2_y2, h_s_arrmul24_fa4_3_y4, h_s_arrmul24_fa5_3_y2, h_s_arrmul24_fa5_3_y4);
  and_gate and_gate_h_s_arrmul24_and6_3_y0(a_6, b_3, h_s_arrmul24_and6_3_y0);
  fa fa_h_s_arrmul24_fa6_3_y2(h_s_arrmul24_and6_3_y0, h_s_arrmul24_fa7_2_y2, h_s_arrmul24_fa5_3_y4, h_s_arrmul24_fa6_3_y2, h_s_arrmul24_fa6_3_y4);
  and_gate and_gate_h_s_arrmul24_and7_3_y0(a_7, b_3, h_s_arrmul24_and7_3_y0);
  fa fa_h_s_arrmul24_fa7_3_y2(h_s_arrmul24_and7_3_y0, h_s_arrmul24_fa8_2_y2, h_s_arrmul24_fa6_3_y4, h_s_arrmul24_fa7_3_y2, h_s_arrmul24_fa7_3_y4);
  and_gate and_gate_h_s_arrmul24_and8_3_y0(a_8, b_3, h_s_arrmul24_and8_3_y0);
  fa fa_h_s_arrmul24_fa8_3_y2(h_s_arrmul24_and8_3_y0, h_s_arrmul24_fa9_2_y2, h_s_arrmul24_fa7_3_y4, h_s_arrmul24_fa8_3_y2, h_s_arrmul24_fa8_3_y4);
  and_gate and_gate_h_s_arrmul24_and9_3_y0(a_9, b_3, h_s_arrmul24_and9_3_y0);
  fa fa_h_s_arrmul24_fa9_3_y2(h_s_arrmul24_and9_3_y0, h_s_arrmul24_fa10_2_y2, h_s_arrmul24_fa8_3_y4, h_s_arrmul24_fa9_3_y2, h_s_arrmul24_fa9_3_y4);
  and_gate and_gate_h_s_arrmul24_and10_3_y0(a_10, b_3, h_s_arrmul24_and10_3_y0);
  fa fa_h_s_arrmul24_fa10_3_y2(h_s_arrmul24_and10_3_y0, h_s_arrmul24_fa11_2_y2, h_s_arrmul24_fa9_3_y4, h_s_arrmul24_fa10_3_y2, h_s_arrmul24_fa10_3_y4);
  and_gate and_gate_h_s_arrmul24_and11_3_y0(a_11, b_3, h_s_arrmul24_and11_3_y0);
  fa fa_h_s_arrmul24_fa11_3_y2(h_s_arrmul24_and11_3_y0, h_s_arrmul24_fa12_2_y2, h_s_arrmul24_fa10_3_y4, h_s_arrmul24_fa11_3_y2, h_s_arrmul24_fa11_3_y4);
  and_gate and_gate_h_s_arrmul24_and12_3_y0(a_12, b_3, h_s_arrmul24_and12_3_y0);
  fa fa_h_s_arrmul24_fa12_3_y2(h_s_arrmul24_and12_3_y0, h_s_arrmul24_fa13_2_y2, h_s_arrmul24_fa11_3_y4, h_s_arrmul24_fa12_3_y2, h_s_arrmul24_fa12_3_y4);
  and_gate and_gate_h_s_arrmul24_and13_3_y0(a_13, b_3, h_s_arrmul24_and13_3_y0);
  fa fa_h_s_arrmul24_fa13_3_y2(h_s_arrmul24_and13_3_y0, h_s_arrmul24_fa14_2_y2, h_s_arrmul24_fa12_3_y4, h_s_arrmul24_fa13_3_y2, h_s_arrmul24_fa13_3_y4);
  and_gate and_gate_h_s_arrmul24_and14_3_y0(a_14, b_3, h_s_arrmul24_and14_3_y0);
  fa fa_h_s_arrmul24_fa14_3_y2(h_s_arrmul24_and14_3_y0, h_s_arrmul24_fa15_2_y2, h_s_arrmul24_fa13_3_y4, h_s_arrmul24_fa14_3_y2, h_s_arrmul24_fa14_3_y4);
  and_gate and_gate_h_s_arrmul24_and15_3_y0(a_15, b_3, h_s_arrmul24_and15_3_y0);
  fa fa_h_s_arrmul24_fa15_3_y2(h_s_arrmul24_and15_3_y0, h_s_arrmul24_fa16_2_y2, h_s_arrmul24_fa14_3_y4, h_s_arrmul24_fa15_3_y2, h_s_arrmul24_fa15_3_y4);
  and_gate and_gate_h_s_arrmul24_and16_3_y0(a_16, b_3, h_s_arrmul24_and16_3_y0);
  fa fa_h_s_arrmul24_fa16_3_y2(h_s_arrmul24_and16_3_y0, h_s_arrmul24_fa17_2_y2, h_s_arrmul24_fa15_3_y4, h_s_arrmul24_fa16_3_y2, h_s_arrmul24_fa16_3_y4);
  and_gate and_gate_h_s_arrmul24_and17_3_y0(a_17, b_3, h_s_arrmul24_and17_3_y0);
  fa fa_h_s_arrmul24_fa17_3_y2(h_s_arrmul24_and17_3_y0, h_s_arrmul24_fa18_2_y2, h_s_arrmul24_fa16_3_y4, h_s_arrmul24_fa17_3_y2, h_s_arrmul24_fa17_3_y4);
  and_gate and_gate_h_s_arrmul24_and18_3_y0(a_18, b_3, h_s_arrmul24_and18_3_y0);
  fa fa_h_s_arrmul24_fa18_3_y2(h_s_arrmul24_and18_3_y0, h_s_arrmul24_fa19_2_y2, h_s_arrmul24_fa17_3_y4, h_s_arrmul24_fa18_3_y2, h_s_arrmul24_fa18_3_y4);
  and_gate and_gate_h_s_arrmul24_and19_3_y0(a_19, b_3, h_s_arrmul24_and19_3_y0);
  fa fa_h_s_arrmul24_fa19_3_y2(h_s_arrmul24_and19_3_y0, h_s_arrmul24_fa20_2_y2, h_s_arrmul24_fa18_3_y4, h_s_arrmul24_fa19_3_y2, h_s_arrmul24_fa19_3_y4);
  and_gate and_gate_h_s_arrmul24_and20_3_y0(a_20, b_3, h_s_arrmul24_and20_3_y0);
  fa fa_h_s_arrmul24_fa20_3_y2(h_s_arrmul24_and20_3_y0, h_s_arrmul24_fa21_2_y2, h_s_arrmul24_fa19_3_y4, h_s_arrmul24_fa20_3_y2, h_s_arrmul24_fa20_3_y4);
  and_gate and_gate_h_s_arrmul24_and21_3_y0(a_21, b_3, h_s_arrmul24_and21_3_y0);
  fa fa_h_s_arrmul24_fa21_3_y2(h_s_arrmul24_and21_3_y0, h_s_arrmul24_fa22_2_y2, h_s_arrmul24_fa20_3_y4, h_s_arrmul24_fa21_3_y2, h_s_arrmul24_fa21_3_y4);
  and_gate and_gate_h_s_arrmul24_and22_3_y0(a_22, b_3, h_s_arrmul24_and22_3_y0);
  fa fa_h_s_arrmul24_fa22_3_y2(h_s_arrmul24_and22_3_y0, h_s_arrmul24_fa23_2_y2, h_s_arrmul24_fa21_3_y4, h_s_arrmul24_fa22_3_y2, h_s_arrmul24_fa22_3_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_3_y0(a_23, b_3, h_s_arrmul24_nand23_3_y0);
  fa fa_h_s_arrmul24_fa23_3_y2(h_s_arrmul24_nand23_3_y0, h_s_arrmul24_fa23_2_y4, h_s_arrmul24_fa22_3_y4, h_s_arrmul24_fa23_3_y2, h_s_arrmul24_fa23_3_y4);
  and_gate and_gate_h_s_arrmul24_and0_4_y0(a_0, b_4, h_s_arrmul24_and0_4_y0);
  ha ha_h_s_arrmul24_ha0_4_y0(h_s_arrmul24_and0_4_y0, h_s_arrmul24_fa1_3_y2, h_s_arrmul24_ha0_4_y0, h_s_arrmul24_ha0_4_y1);
  and_gate and_gate_h_s_arrmul24_and1_4_y0(a_1, b_4, h_s_arrmul24_and1_4_y0);
  fa fa_h_s_arrmul24_fa1_4_y2(h_s_arrmul24_and1_4_y0, h_s_arrmul24_fa2_3_y2, h_s_arrmul24_ha0_4_y1, h_s_arrmul24_fa1_4_y2, h_s_arrmul24_fa1_4_y4);
  and_gate and_gate_h_s_arrmul24_and2_4_y0(a_2, b_4, h_s_arrmul24_and2_4_y0);
  fa fa_h_s_arrmul24_fa2_4_y2(h_s_arrmul24_and2_4_y0, h_s_arrmul24_fa3_3_y2, h_s_arrmul24_fa1_4_y4, h_s_arrmul24_fa2_4_y2, h_s_arrmul24_fa2_4_y4);
  and_gate and_gate_h_s_arrmul24_and3_4_y0(a_3, b_4, h_s_arrmul24_and3_4_y0);
  fa fa_h_s_arrmul24_fa3_4_y2(h_s_arrmul24_and3_4_y0, h_s_arrmul24_fa4_3_y2, h_s_arrmul24_fa2_4_y4, h_s_arrmul24_fa3_4_y2, h_s_arrmul24_fa3_4_y4);
  and_gate and_gate_h_s_arrmul24_and4_4_y0(a_4, b_4, h_s_arrmul24_and4_4_y0);
  fa fa_h_s_arrmul24_fa4_4_y2(h_s_arrmul24_and4_4_y0, h_s_arrmul24_fa5_3_y2, h_s_arrmul24_fa3_4_y4, h_s_arrmul24_fa4_4_y2, h_s_arrmul24_fa4_4_y4);
  and_gate and_gate_h_s_arrmul24_and5_4_y0(a_5, b_4, h_s_arrmul24_and5_4_y0);
  fa fa_h_s_arrmul24_fa5_4_y2(h_s_arrmul24_and5_4_y0, h_s_arrmul24_fa6_3_y2, h_s_arrmul24_fa4_4_y4, h_s_arrmul24_fa5_4_y2, h_s_arrmul24_fa5_4_y4);
  and_gate and_gate_h_s_arrmul24_and6_4_y0(a_6, b_4, h_s_arrmul24_and6_4_y0);
  fa fa_h_s_arrmul24_fa6_4_y2(h_s_arrmul24_and6_4_y0, h_s_arrmul24_fa7_3_y2, h_s_arrmul24_fa5_4_y4, h_s_arrmul24_fa6_4_y2, h_s_arrmul24_fa6_4_y4);
  and_gate and_gate_h_s_arrmul24_and7_4_y0(a_7, b_4, h_s_arrmul24_and7_4_y0);
  fa fa_h_s_arrmul24_fa7_4_y2(h_s_arrmul24_and7_4_y0, h_s_arrmul24_fa8_3_y2, h_s_arrmul24_fa6_4_y4, h_s_arrmul24_fa7_4_y2, h_s_arrmul24_fa7_4_y4);
  and_gate and_gate_h_s_arrmul24_and8_4_y0(a_8, b_4, h_s_arrmul24_and8_4_y0);
  fa fa_h_s_arrmul24_fa8_4_y2(h_s_arrmul24_and8_4_y0, h_s_arrmul24_fa9_3_y2, h_s_arrmul24_fa7_4_y4, h_s_arrmul24_fa8_4_y2, h_s_arrmul24_fa8_4_y4);
  and_gate and_gate_h_s_arrmul24_and9_4_y0(a_9, b_4, h_s_arrmul24_and9_4_y0);
  fa fa_h_s_arrmul24_fa9_4_y2(h_s_arrmul24_and9_4_y0, h_s_arrmul24_fa10_3_y2, h_s_arrmul24_fa8_4_y4, h_s_arrmul24_fa9_4_y2, h_s_arrmul24_fa9_4_y4);
  and_gate and_gate_h_s_arrmul24_and10_4_y0(a_10, b_4, h_s_arrmul24_and10_4_y0);
  fa fa_h_s_arrmul24_fa10_4_y2(h_s_arrmul24_and10_4_y0, h_s_arrmul24_fa11_3_y2, h_s_arrmul24_fa9_4_y4, h_s_arrmul24_fa10_4_y2, h_s_arrmul24_fa10_4_y4);
  and_gate and_gate_h_s_arrmul24_and11_4_y0(a_11, b_4, h_s_arrmul24_and11_4_y0);
  fa fa_h_s_arrmul24_fa11_4_y2(h_s_arrmul24_and11_4_y0, h_s_arrmul24_fa12_3_y2, h_s_arrmul24_fa10_4_y4, h_s_arrmul24_fa11_4_y2, h_s_arrmul24_fa11_4_y4);
  and_gate and_gate_h_s_arrmul24_and12_4_y0(a_12, b_4, h_s_arrmul24_and12_4_y0);
  fa fa_h_s_arrmul24_fa12_4_y2(h_s_arrmul24_and12_4_y0, h_s_arrmul24_fa13_3_y2, h_s_arrmul24_fa11_4_y4, h_s_arrmul24_fa12_4_y2, h_s_arrmul24_fa12_4_y4);
  and_gate and_gate_h_s_arrmul24_and13_4_y0(a_13, b_4, h_s_arrmul24_and13_4_y0);
  fa fa_h_s_arrmul24_fa13_4_y2(h_s_arrmul24_and13_4_y0, h_s_arrmul24_fa14_3_y2, h_s_arrmul24_fa12_4_y4, h_s_arrmul24_fa13_4_y2, h_s_arrmul24_fa13_4_y4);
  and_gate and_gate_h_s_arrmul24_and14_4_y0(a_14, b_4, h_s_arrmul24_and14_4_y0);
  fa fa_h_s_arrmul24_fa14_4_y2(h_s_arrmul24_and14_4_y0, h_s_arrmul24_fa15_3_y2, h_s_arrmul24_fa13_4_y4, h_s_arrmul24_fa14_4_y2, h_s_arrmul24_fa14_4_y4);
  and_gate and_gate_h_s_arrmul24_and15_4_y0(a_15, b_4, h_s_arrmul24_and15_4_y0);
  fa fa_h_s_arrmul24_fa15_4_y2(h_s_arrmul24_and15_4_y0, h_s_arrmul24_fa16_3_y2, h_s_arrmul24_fa14_4_y4, h_s_arrmul24_fa15_4_y2, h_s_arrmul24_fa15_4_y4);
  and_gate and_gate_h_s_arrmul24_and16_4_y0(a_16, b_4, h_s_arrmul24_and16_4_y0);
  fa fa_h_s_arrmul24_fa16_4_y2(h_s_arrmul24_and16_4_y0, h_s_arrmul24_fa17_3_y2, h_s_arrmul24_fa15_4_y4, h_s_arrmul24_fa16_4_y2, h_s_arrmul24_fa16_4_y4);
  and_gate and_gate_h_s_arrmul24_and17_4_y0(a_17, b_4, h_s_arrmul24_and17_4_y0);
  fa fa_h_s_arrmul24_fa17_4_y2(h_s_arrmul24_and17_4_y0, h_s_arrmul24_fa18_3_y2, h_s_arrmul24_fa16_4_y4, h_s_arrmul24_fa17_4_y2, h_s_arrmul24_fa17_4_y4);
  and_gate and_gate_h_s_arrmul24_and18_4_y0(a_18, b_4, h_s_arrmul24_and18_4_y0);
  fa fa_h_s_arrmul24_fa18_4_y2(h_s_arrmul24_and18_4_y0, h_s_arrmul24_fa19_3_y2, h_s_arrmul24_fa17_4_y4, h_s_arrmul24_fa18_4_y2, h_s_arrmul24_fa18_4_y4);
  and_gate and_gate_h_s_arrmul24_and19_4_y0(a_19, b_4, h_s_arrmul24_and19_4_y0);
  fa fa_h_s_arrmul24_fa19_4_y2(h_s_arrmul24_and19_4_y0, h_s_arrmul24_fa20_3_y2, h_s_arrmul24_fa18_4_y4, h_s_arrmul24_fa19_4_y2, h_s_arrmul24_fa19_4_y4);
  and_gate and_gate_h_s_arrmul24_and20_4_y0(a_20, b_4, h_s_arrmul24_and20_4_y0);
  fa fa_h_s_arrmul24_fa20_4_y2(h_s_arrmul24_and20_4_y0, h_s_arrmul24_fa21_3_y2, h_s_arrmul24_fa19_4_y4, h_s_arrmul24_fa20_4_y2, h_s_arrmul24_fa20_4_y4);
  and_gate and_gate_h_s_arrmul24_and21_4_y0(a_21, b_4, h_s_arrmul24_and21_4_y0);
  fa fa_h_s_arrmul24_fa21_4_y2(h_s_arrmul24_and21_4_y0, h_s_arrmul24_fa22_3_y2, h_s_arrmul24_fa20_4_y4, h_s_arrmul24_fa21_4_y2, h_s_arrmul24_fa21_4_y4);
  and_gate and_gate_h_s_arrmul24_and22_4_y0(a_22, b_4, h_s_arrmul24_and22_4_y0);
  fa fa_h_s_arrmul24_fa22_4_y2(h_s_arrmul24_and22_4_y0, h_s_arrmul24_fa23_3_y2, h_s_arrmul24_fa21_4_y4, h_s_arrmul24_fa22_4_y2, h_s_arrmul24_fa22_4_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_4_y0(a_23, b_4, h_s_arrmul24_nand23_4_y0);
  fa fa_h_s_arrmul24_fa23_4_y2(h_s_arrmul24_nand23_4_y0, h_s_arrmul24_fa23_3_y4, h_s_arrmul24_fa22_4_y4, h_s_arrmul24_fa23_4_y2, h_s_arrmul24_fa23_4_y4);
  and_gate and_gate_h_s_arrmul24_and0_5_y0(a_0, b_5, h_s_arrmul24_and0_5_y0);
  ha ha_h_s_arrmul24_ha0_5_y0(h_s_arrmul24_and0_5_y0, h_s_arrmul24_fa1_4_y2, h_s_arrmul24_ha0_5_y0, h_s_arrmul24_ha0_5_y1);
  and_gate and_gate_h_s_arrmul24_and1_5_y0(a_1, b_5, h_s_arrmul24_and1_5_y0);
  fa fa_h_s_arrmul24_fa1_5_y2(h_s_arrmul24_and1_5_y0, h_s_arrmul24_fa2_4_y2, h_s_arrmul24_ha0_5_y1, h_s_arrmul24_fa1_5_y2, h_s_arrmul24_fa1_5_y4);
  and_gate and_gate_h_s_arrmul24_and2_5_y0(a_2, b_5, h_s_arrmul24_and2_5_y0);
  fa fa_h_s_arrmul24_fa2_5_y2(h_s_arrmul24_and2_5_y0, h_s_arrmul24_fa3_4_y2, h_s_arrmul24_fa1_5_y4, h_s_arrmul24_fa2_5_y2, h_s_arrmul24_fa2_5_y4);
  and_gate and_gate_h_s_arrmul24_and3_5_y0(a_3, b_5, h_s_arrmul24_and3_5_y0);
  fa fa_h_s_arrmul24_fa3_5_y2(h_s_arrmul24_and3_5_y0, h_s_arrmul24_fa4_4_y2, h_s_arrmul24_fa2_5_y4, h_s_arrmul24_fa3_5_y2, h_s_arrmul24_fa3_5_y4);
  and_gate and_gate_h_s_arrmul24_and4_5_y0(a_4, b_5, h_s_arrmul24_and4_5_y0);
  fa fa_h_s_arrmul24_fa4_5_y2(h_s_arrmul24_and4_5_y0, h_s_arrmul24_fa5_4_y2, h_s_arrmul24_fa3_5_y4, h_s_arrmul24_fa4_5_y2, h_s_arrmul24_fa4_5_y4);
  and_gate and_gate_h_s_arrmul24_and5_5_y0(a_5, b_5, h_s_arrmul24_and5_5_y0);
  fa fa_h_s_arrmul24_fa5_5_y2(h_s_arrmul24_and5_5_y0, h_s_arrmul24_fa6_4_y2, h_s_arrmul24_fa4_5_y4, h_s_arrmul24_fa5_5_y2, h_s_arrmul24_fa5_5_y4);
  and_gate and_gate_h_s_arrmul24_and6_5_y0(a_6, b_5, h_s_arrmul24_and6_5_y0);
  fa fa_h_s_arrmul24_fa6_5_y2(h_s_arrmul24_and6_5_y0, h_s_arrmul24_fa7_4_y2, h_s_arrmul24_fa5_5_y4, h_s_arrmul24_fa6_5_y2, h_s_arrmul24_fa6_5_y4);
  and_gate and_gate_h_s_arrmul24_and7_5_y0(a_7, b_5, h_s_arrmul24_and7_5_y0);
  fa fa_h_s_arrmul24_fa7_5_y2(h_s_arrmul24_and7_5_y0, h_s_arrmul24_fa8_4_y2, h_s_arrmul24_fa6_5_y4, h_s_arrmul24_fa7_5_y2, h_s_arrmul24_fa7_5_y4);
  and_gate and_gate_h_s_arrmul24_and8_5_y0(a_8, b_5, h_s_arrmul24_and8_5_y0);
  fa fa_h_s_arrmul24_fa8_5_y2(h_s_arrmul24_and8_5_y0, h_s_arrmul24_fa9_4_y2, h_s_arrmul24_fa7_5_y4, h_s_arrmul24_fa8_5_y2, h_s_arrmul24_fa8_5_y4);
  and_gate and_gate_h_s_arrmul24_and9_5_y0(a_9, b_5, h_s_arrmul24_and9_5_y0);
  fa fa_h_s_arrmul24_fa9_5_y2(h_s_arrmul24_and9_5_y0, h_s_arrmul24_fa10_4_y2, h_s_arrmul24_fa8_5_y4, h_s_arrmul24_fa9_5_y2, h_s_arrmul24_fa9_5_y4);
  and_gate and_gate_h_s_arrmul24_and10_5_y0(a_10, b_5, h_s_arrmul24_and10_5_y0);
  fa fa_h_s_arrmul24_fa10_5_y2(h_s_arrmul24_and10_5_y0, h_s_arrmul24_fa11_4_y2, h_s_arrmul24_fa9_5_y4, h_s_arrmul24_fa10_5_y2, h_s_arrmul24_fa10_5_y4);
  and_gate and_gate_h_s_arrmul24_and11_5_y0(a_11, b_5, h_s_arrmul24_and11_5_y0);
  fa fa_h_s_arrmul24_fa11_5_y2(h_s_arrmul24_and11_5_y0, h_s_arrmul24_fa12_4_y2, h_s_arrmul24_fa10_5_y4, h_s_arrmul24_fa11_5_y2, h_s_arrmul24_fa11_5_y4);
  and_gate and_gate_h_s_arrmul24_and12_5_y0(a_12, b_5, h_s_arrmul24_and12_5_y0);
  fa fa_h_s_arrmul24_fa12_5_y2(h_s_arrmul24_and12_5_y0, h_s_arrmul24_fa13_4_y2, h_s_arrmul24_fa11_5_y4, h_s_arrmul24_fa12_5_y2, h_s_arrmul24_fa12_5_y4);
  and_gate and_gate_h_s_arrmul24_and13_5_y0(a_13, b_5, h_s_arrmul24_and13_5_y0);
  fa fa_h_s_arrmul24_fa13_5_y2(h_s_arrmul24_and13_5_y0, h_s_arrmul24_fa14_4_y2, h_s_arrmul24_fa12_5_y4, h_s_arrmul24_fa13_5_y2, h_s_arrmul24_fa13_5_y4);
  and_gate and_gate_h_s_arrmul24_and14_5_y0(a_14, b_5, h_s_arrmul24_and14_5_y0);
  fa fa_h_s_arrmul24_fa14_5_y2(h_s_arrmul24_and14_5_y0, h_s_arrmul24_fa15_4_y2, h_s_arrmul24_fa13_5_y4, h_s_arrmul24_fa14_5_y2, h_s_arrmul24_fa14_5_y4);
  and_gate and_gate_h_s_arrmul24_and15_5_y0(a_15, b_5, h_s_arrmul24_and15_5_y0);
  fa fa_h_s_arrmul24_fa15_5_y2(h_s_arrmul24_and15_5_y0, h_s_arrmul24_fa16_4_y2, h_s_arrmul24_fa14_5_y4, h_s_arrmul24_fa15_5_y2, h_s_arrmul24_fa15_5_y4);
  and_gate and_gate_h_s_arrmul24_and16_5_y0(a_16, b_5, h_s_arrmul24_and16_5_y0);
  fa fa_h_s_arrmul24_fa16_5_y2(h_s_arrmul24_and16_5_y0, h_s_arrmul24_fa17_4_y2, h_s_arrmul24_fa15_5_y4, h_s_arrmul24_fa16_5_y2, h_s_arrmul24_fa16_5_y4);
  and_gate and_gate_h_s_arrmul24_and17_5_y0(a_17, b_5, h_s_arrmul24_and17_5_y0);
  fa fa_h_s_arrmul24_fa17_5_y2(h_s_arrmul24_and17_5_y0, h_s_arrmul24_fa18_4_y2, h_s_arrmul24_fa16_5_y4, h_s_arrmul24_fa17_5_y2, h_s_arrmul24_fa17_5_y4);
  and_gate and_gate_h_s_arrmul24_and18_5_y0(a_18, b_5, h_s_arrmul24_and18_5_y0);
  fa fa_h_s_arrmul24_fa18_5_y2(h_s_arrmul24_and18_5_y0, h_s_arrmul24_fa19_4_y2, h_s_arrmul24_fa17_5_y4, h_s_arrmul24_fa18_5_y2, h_s_arrmul24_fa18_5_y4);
  and_gate and_gate_h_s_arrmul24_and19_5_y0(a_19, b_5, h_s_arrmul24_and19_5_y0);
  fa fa_h_s_arrmul24_fa19_5_y2(h_s_arrmul24_and19_5_y0, h_s_arrmul24_fa20_4_y2, h_s_arrmul24_fa18_5_y4, h_s_arrmul24_fa19_5_y2, h_s_arrmul24_fa19_5_y4);
  and_gate and_gate_h_s_arrmul24_and20_5_y0(a_20, b_5, h_s_arrmul24_and20_5_y0);
  fa fa_h_s_arrmul24_fa20_5_y2(h_s_arrmul24_and20_5_y0, h_s_arrmul24_fa21_4_y2, h_s_arrmul24_fa19_5_y4, h_s_arrmul24_fa20_5_y2, h_s_arrmul24_fa20_5_y4);
  and_gate and_gate_h_s_arrmul24_and21_5_y0(a_21, b_5, h_s_arrmul24_and21_5_y0);
  fa fa_h_s_arrmul24_fa21_5_y2(h_s_arrmul24_and21_5_y0, h_s_arrmul24_fa22_4_y2, h_s_arrmul24_fa20_5_y4, h_s_arrmul24_fa21_5_y2, h_s_arrmul24_fa21_5_y4);
  and_gate and_gate_h_s_arrmul24_and22_5_y0(a_22, b_5, h_s_arrmul24_and22_5_y0);
  fa fa_h_s_arrmul24_fa22_5_y2(h_s_arrmul24_and22_5_y0, h_s_arrmul24_fa23_4_y2, h_s_arrmul24_fa21_5_y4, h_s_arrmul24_fa22_5_y2, h_s_arrmul24_fa22_5_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_5_y0(a_23, b_5, h_s_arrmul24_nand23_5_y0);
  fa fa_h_s_arrmul24_fa23_5_y2(h_s_arrmul24_nand23_5_y0, h_s_arrmul24_fa23_4_y4, h_s_arrmul24_fa22_5_y4, h_s_arrmul24_fa23_5_y2, h_s_arrmul24_fa23_5_y4);
  and_gate and_gate_h_s_arrmul24_and0_6_y0(a_0, b_6, h_s_arrmul24_and0_6_y0);
  ha ha_h_s_arrmul24_ha0_6_y0(h_s_arrmul24_and0_6_y0, h_s_arrmul24_fa1_5_y2, h_s_arrmul24_ha0_6_y0, h_s_arrmul24_ha0_6_y1);
  and_gate and_gate_h_s_arrmul24_and1_6_y0(a_1, b_6, h_s_arrmul24_and1_6_y0);
  fa fa_h_s_arrmul24_fa1_6_y2(h_s_arrmul24_and1_6_y0, h_s_arrmul24_fa2_5_y2, h_s_arrmul24_ha0_6_y1, h_s_arrmul24_fa1_6_y2, h_s_arrmul24_fa1_6_y4);
  and_gate and_gate_h_s_arrmul24_and2_6_y0(a_2, b_6, h_s_arrmul24_and2_6_y0);
  fa fa_h_s_arrmul24_fa2_6_y2(h_s_arrmul24_and2_6_y0, h_s_arrmul24_fa3_5_y2, h_s_arrmul24_fa1_6_y4, h_s_arrmul24_fa2_6_y2, h_s_arrmul24_fa2_6_y4);
  and_gate and_gate_h_s_arrmul24_and3_6_y0(a_3, b_6, h_s_arrmul24_and3_6_y0);
  fa fa_h_s_arrmul24_fa3_6_y2(h_s_arrmul24_and3_6_y0, h_s_arrmul24_fa4_5_y2, h_s_arrmul24_fa2_6_y4, h_s_arrmul24_fa3_6_y2, h_s_arrmul24_fa3_6_y4);
  and_gate and_gate_h_s_arrmul24_and4_6_y0(a_4, b_6, h_s_arrmul24_and4_6_y0);
  fa fa_h_s_arrmul24_fa4_6_y2(h_s_arrmul24_and4_6_y0, h_s_arrmul24_fa5_5_y2, h_s_arrmul24_fa3_6_y4, h_s_arrmul24_fa4_6_y2, h_s_arrmul24_fa4_6_y4);
  and_gate and_gate_h_s_arrmul24_and5_6_y0(a_5, b_6, h_s_arrmul24_and5_6_y0);
  fa fa_h_s_arrmul24_fa5_6_y2(h_s_arrmul24_and5_6_y0, h_s_arrmul24_fa6_5_y2, h_s_arrmul24_fa4_6_y4, h_s_arrmul24_fa5_6_y2, h_s_arrmul24_fa5_6_y4);
  and_gate and_gate_h_s_arrmul24_and6_6_y0(a_6, b_6, h_s_arrmul24_and6_6_y0);
  fa fa_h_s_arrmul24_fa6_6_y2(h_s_arrmul24_and6_6_y0, h_s_arrmul24_fa7_5_y2, h_s_arrmul24_fa5_6_y4, h_s_arrmul24_fa6_6_y2, h_s_arrmul24_fa6_6_y4);
  and_gate and_gate_h_s_arrmul24_and7_6_y0(a_7, b_6, h_s_arrmul24_and7_6_y0);
  fa fa_h_s_arrmul24_fa7_6_y2(h_s_arrmul24_and7_6_y0, h_s_arrmul24_fa8_5_y2, h_s_arrmul24_fa6_6_y4, h_s_arrmul24_fa7_6_y2, h_s_arrmul24_fa7_6_y4);
  and_gate and_gate_h_s_arrmul24_and8_6_y0(a_8, b_6, h_s_arrmul24_and8_6_y0);
  fa fa_h_s_arrmul24_fa8_6_y2(h_s_arrmul24_and8_6_y0, h_s_arrmul24_fa9_5_y2, h_s_arrmul24_fa7_6_y4, h_s_arrmul24_fa8_6_y2, h_s_arrmul24_fa8_6_y4);
  and_gate and_gate_h_s_arrmul24_and9_6_y0(a_9, b_6, h_s_arrmul24_and9_6_y0);
  fa fa_h_s_arrmul24_fa9_6_y2(h_s_arrmul24_and9_6_y0, h_s_arrmul24_fa10_5_y2, h_s_arrmul24_fa8_6_y4, h_s_arrmul24_fa9_6_y2, h_s_arrmul24_fa9_6_y4);
  and_gate and_gate_h_s_arrmul24_and10_6_y0(a_10, b_6, h_s_arrmul24_and10_6_y0);
  fa fa_h_s_arrmul24_fa10_6_y2(h_s_arrmul24_and10_6_y0, h_s_arrmul24_fa11_5_y2, h_s_arrmul24_fa9_6_y4, h_s_arrmul24_fa10_6_y2, h_s_arrmul24_fa10_6_y4);
  and_gate and_gate_h_s_arrmul24_and11_6_y0(a_11, b_6, h_s_arrmul24_and11_6_y0);
  fa fa_h_s_arrmul24_fa11_6_y2(h_s_arrmul24_and11_6_y0, h_s_arrmul24_fa12_5_y2, h_s_arrmul24_fa10_6_y4, h_s_arrmul24_fa11_6_y2, h_s_arrmul24_fa11_6_y4);
  and_gate and_gate_h_s_arrmul24_and12_6_y0(a_12, b_6, h_s_arrmul24_and12_6_y0);
  fa fa_h_s_arrmul24_fa12_6_y2(h_s_arrmul24_and12_6_y0, h_s_arrmul24_fa13_5_y2, h_s_arrmul24_fa11_6_y4, h_s_arrmul24_fa12_6_y2, h_s_arrmul24_fa12_6_y4);
  and_gate and_gate_h_s_arrmul24_and13_6_y0(a_13, b_6, h_s_arrmul24_and13_6_y0);
  fa fa_h_s_arrmul24_fa13_6_y2(h_s_arrmul24_and13_6_y0, h_s_arrmul24_fa14_5_y2, h_s_arrmul24_fa12_6_y4, h_s_arrmul24_fa13_6_y2, h_s_arrmul24_fa13_6_y4);
  and_gate and_gate_h_s_arrmul24_and14_6_y0(a_14, b_6, h_s_arrmul24_and14_6_y0);
  fa fa_h_s_arrmul24_fa14_6_y2(h_s_arrmul24_and14_6_y0, h_s_arrmul24_fa15_5_y2, h_s_arrmul24_fa13_6_y4, h_s_arrmul24_fa14_6_y2, h_s_arrmul24_fa14_6_y4);
  and_gate and_gate_h_s_arrmul24_and15_6_y0(a_15, b_6, h_s_arrmul24_and15_6_y0);
  fa fa_h_s_arrmul24_fa15_6_y2(h_s_arrmul24_and15_6_y0, h_s_arrmul24_fa16_5_y2, h_s_arrmul24_fa14_6_y4, h_s_arrmul24_fa15_6_y2, h_s_arrmul24_fa15_6_y4);
  and_gate and_gate_h_s_arrmul24_and16_6_y0(a_16, b_6, h_s_arrmul24_and16_6_y0);
  fa fa_h_s_arrmul24_fa16_6_y2(h_s_arrmul24_and16_6_y0, h_s_arrmul24_fa17_5_y2, h_s_arrmul24_fa15_6_y4, h_s_arrmul24_fa16_6_y2, h_s_arrmul24_fa16_6_y4);
  and_gate and_gate_h_s_arrmul24_and17_6_y0(a_17, b_6, h_s_arrmul24_and17_6_y0);
  fa fa_h_s_arrmul24_fa17_6_y2(h_s_arrmul24_and17_6_y0, h_s_arrmul24_fa18_5_y2, h_s_arrmul24_fa16_6_y4, h_s_arrmul24_fa17_6_y2, h_s_arrmul24_fa17_6_y4);
  and_gate and_gate_h_s_arrmul24_and18_6_y0(a_18, b_6, h_s_arrmul24_and18_6_y0);
  fa fa_h_s_arrmul24_fa18_6_y2(h_s_arrmul24_and18_6_y0, h_s_arrmul24_fa19_5_y2, h_s_arrmul24_fa17_6_y4, h_s_arrmul24_fa18_6_y2, h_s_arrmul24_fa18_6_y4);
  and_gate and_gate_h_s_arrmul24_and19_6_y0(a_19, b_6, h_s_arrmul24_and19_6_y0);
  fa fa_h_s_arrmul24_fa19_6_y2(h_s_arrmul24_and19_6_y0, h_s_arrmul24_fa20_5_y2, h_s_arrmul24_fa18_6_y4, h_s_arrmul24_fa19_6_y2, h_s_arrmul24_fa19_6_y4);
  and_gate and_gate_h_s_arrmul24_and20_6_y0(a_20, b_6, h_s_arrmul24_and20_6_y0);
  fa fa_h_s_arrmul24_fa20_6_y2(h_s_arrmul24_and20_6_y0, h_s_arrmul24_fa21_5_y2, h_s_arrmul24_fa19_6_y4, h_s_arrmul24_fa20_6_y2, h_s_arrmul24_fa20_6_y4);
  and_gate and_gate_h_s_arrmul24_and21_6_y0(a_21, b_6, h_s_arrmul24_and21_6_y0);
  fa fa_h_s_arrmul24_fa21_6_y2(h_s_arrmul24_and21_6_y0, h_s_arrmul24_fa22_5_y2, h_s_arrmul24_fa20_6_y4, h_s_arrmul24_fa21_6_y2, h_s_arrmul24_fa21_6_y4);
  and_gate and_gate_h_s_arrmul24_and22_6_y0(a_22, b_6, h_s_arrmul24_and22_6_y0);
  fa fa_h_s_arrmul24_fa22_6_y2(h_s_arrmul24_and22_6_y0, h_s_arrmul24_fa23_5_y2, h_s_arrmul24_fa21_6_y4, h_s_arrmul24_fa22_6_y2, h_s_arrmul24_fa22_6_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_6_y0(a_23, b_6, h_s_arrmul24_nand23_6_y0);
  fa fa_h_s_arrmul24_fa23_6_y2(h_s_arrmul24_nand23_6_y0, h_s_arrmul24_fa23_5_y4, h_s_arrmul24_fa22_6_y4, h_s_arrmul24_fa23_6_y2, h_s_arrmul24_fa23_6_y4);
  and_gate and_gate_h_s_arrmul24_and0_7_y0(a_0, b_7, h_s_arrmul24_and0_7_y0);
  ha ha_h_s_arrmul24_ha0_7_y0(h_s_arrmul24_and0_7_y0, h_s_arrmul24_fa1_6_y2, h_s_arrmul24_ha0_7_y0, h_s_arrmul24_ha0_7_y1);
  and_gate and_gate_h_s_arrmul24_and1_7_y0(a_1, b_7, h_s_arrmul24_and1_7_y0);
  fa fa_h_s_arrmul24_fa1_7_y2(h_s_arrmul24_and1_7_y0, h_s_arrmul24_fa2_6_y2, h_s_arrmul24_ha0_7_y1, h_s_arrmul24_fa1_7_y2, h_s_arrmul24_fa1_7_y4);
  and_gate and_gate_h_s_arrmul24_and2_7_y0(a_2, b_7, h_s_arrmul24_and2_7_y0);
  fa fa_h_s_arrmul24_fa2_7_y2(h_s_arrmul24_and2_7_y0, h_s_arrmul24_fa3_6_y2, h_s_arrmul24_fa1_7_y4, h_s_arrmul24_fa2_7_y2, h_s_arrmul24_fa2_7_y4);
  and_gate and_gate_h_s_arrmul24_and3_7_y0(a_3, b_7, h_s_arrmul24_and3_7_y0);
  fa fa_h_s_arrmul24_fa3_7_y2(h_s_arrmul24_and3_7_y0, h_s_arrmul24_fa4_6_y2, h_s_arrmul24_fa2_7_y4, h_s_arrmul24_fa3_7_y2, h_s_arrmul24_fa3_7_y4);
  and_gate and_gate_h_s_arrmul24_and4_7_y0(a_4, b_7, h_s_arrmul24_and4_7_y0);
  fa fa_h_s_arrmul24_fa4_7_y2(h_s_arrmul24_and4_7_y0, h_s_arrmul24_fa5_6_y2, h_s_arrmul24_fa3_7_y4, h_s_arrmul24_fa4_7_y2, h_s_arrmul24_fa4_7_y4);
  and_gate and_gate_h_s_arrmul24_and5_7_y0(a_5, b_7, h_s_arrmul24_and5_7_y0);
  fa fa_h_s_arrmul24_fa5_7_y2(h_s_arrmul24_and5_7_y0, h_s_arrmul24_fa6_6_y2, h_s_arrmul24_fa4_7_y4, h_s_arrmul24_fa5_7_y2, h_s_arrmul24_fa5_7_y4);
  and_gate and_gate_h_s_arrmul24_and6_7_y0(a_6, b_7, h_s_arrmul24_and6_7_y0);
  fa fa_h_s_arrmul24_fa6_7_y2(h_s_arrmul24_and6_7_y0, h_s_arrmul24_fa7_6_y2, h_s_arrmul24_fa5_7_y4, h_s_arrmul24_fa6_7_y2, h_s_arrmul24_fa6_7_y4);
  and_gate and_gate_h_s_arrmul24_and7_7_y0(a_7, b_7, h_s_arrmul24_and7_7_y0);
  fa fa_h_s_arrmul24_fa7_7_y2(h_s_arrmul24_and7_7_y0, h_s_arrmul24_fa8_6_y2, h_s_arrmul24_fa6_7_y4, h_s_arrmul24_fa7_7_y2, h_s_arrmul24_fa7_7_y4);
  and_gate and_gate_h_s_arrmul24_and8_7_y0(a_8, b_7, h_s_arrmul24_and8_7_y0);
  fa fa_h_s_arrmul24_fa8_7_y2(h_s_arrmul24_and8_7_y0, h_s_arrmul24_fa9_6_y2, h_s_arrmul24_fa7_7_y4, h_s_arrmul24_fa8_7_y2, h_s_arrmul24_fa8_7_y4);
  and_gate and_gate_h_s_arrmul24_and9_7_y0(a_9, b_7, h_s_arrmul24_and9_7_y0);
  fa fa_h_s_arrmul24_fa9_7_y2(h_s_arrmul24_and9_7_y0, h_s_arrmul24_fa10_6_y2, h_s_arrmul24_fa8_7_y4, h_s_arrmul24_fa9_7_y2, h_s_arrmul24_fa9_7_y4);
  and_gate and_gate_h_s_arrmul24_and10_7_y0(a_10, b_7, h_s_arrmul24_and10_7_y0);
  fa fa_h_s_arrmul24_fa10_7_y2(h_s_arrmul24_and10_7_y0, h_s_arrmul24_fa11_6_y2, h_s_arrmul24_fa9_7_y4, h_s_arrmul24_fa10_7_y2, h_s_arrmul24_fa10_7_y4);
  and_gate and_gate_h_s_arrmul24_and11_7_y0(a_11, b_7, h_s_arrmul24_and11_7_y0);
  fa fa_h_s_arrmul24_fa11_7_y2(h_s_arrmul24_and11_7_y0, h_s_arrmul24_fa12_6_y2, h_s_arrmul24_fa10_7_y4, h_s_arrmul24_fa11_7_y2, h_s_arrmul24_fa11_7_y4);
  and_gate and_gate_h_s_arrmul24_and12_7_y0(a_12, b_7, h_s_arrmul24_and12_7_y0);
  fa fa_h_s_arrmul24_fa12_7_y2(h_s_arrmul24_and12_7_y0, h_s_arrmul24_fa13_6_y2, h_s_arrmul24_fa11_7_y4, h_s_arrmul24_fa12_7_y2, h_s_arrmul24_fa12_7_y4);
  and_gate and_gate_h_s_arrmul24_and13_7_y0(a_13, b_7, h_s_arrmul24_and13_7_y0);
  fa fa_h_s_arrmul24_fa13_7_y2(h_s_arrmul24_and13_7_y0, h_s_arrmul24_fa14_6_y2, h_s_arrmul24_fa12_7_y4, h_s_arrmul24_fa13_7_y2, h_s_arrmul24_fa13_7_y4);
  and_gate and_gate_h_s_arrmul24_and14_7_y0(a_14, b_7, h_s_arrmul24_and14_7_y0);
  fa fa_h_s_arrmul24_fa14_7_y2(h_s_arrmul24_and14_7_y0, h_s_arrmul24_fa15_6_y2, h_s_arrmul24_fa13_7_y4, h_s_arrmul24_fa14_7_y2, h_s_arrmul24_fa14_7_y4);
  and_gate and_gate_h_s_arrmul24_and15_7_y0(a_15, b_7, h_s_arrmul24_and15_7_y0);
  fa fa_h_s_arrmul24_fa15_7_y2(h_s_arrmul24_and15_7_y0, h_s_arrmul24_fa16_6_y2, h_s_arrmul24_fa14_7_y4, h_s_arrmul24_fa15_7_y2, h_s_arrmul24_fa15_7_y4);
  and_gate and_gate_h_s_arrmul24_and16_7_y0(a_16, b_7, h_s_arrmul24_and16_7_y0);
  fa fa_h_s_arrmul24_fa16_7_y2(h_s_arrmul24_and16_7_y0, h_s_arrmul24_fa17_6_y2, h_s_arrmul24_fa15_7_y4, h_s_arrmul24_fa16_7_y2, h_s_arrmul24_fa16_7_y4);
  and_gate and_gate_h_s_arrmul24_and17_7_y0(a_17, b_7, h_s_arrmul24_and17_7_y0);
  fa fa_h_s_arrmul24_fa17_7_y2(h_s_arrmul24_and17_7_y0, h_s_arrmul24_fa18_6_y2, h_s_arrmul24_fa16_7_y4, h_s_arrmul24_fa17_7_y2, h_s_arrmul24_fa17_7_y4);
  and_gate and_gate_h_s_arrmul24_and18_7_y0(a_18, b_7, h_s_arrmul24_and18_7_y0);
  fa fa_h_s_arrmul24_fa18_7_y2(h_s_arrmul24_and18_7_y0, h_s_arrmul24_fa19_6_y2, h_s_arrmul24_fa17_7_y4, h_s_arrmul24_fa18_7_y2, h_s_arrmul24_fa18_7_y4);
  and_gate and_gate_h_s_arrmul24_and19_7_y0(a_19, b_7, h_s_arrmul24_and19_7_y0);
  fa fa_h_s_arrmul24_fa19_7_y2(h_s_arrmul24_and19_7_y0, h_s_arrmul24_fa20_6_y2, h_s_arrmul24_fa18_7_y4, h_s_arrmul24_fa19_7_y2, h_s_arrmul24_fa19_7_y4);
  and_gate and_gate_h_s_arrmul24_and20_7_y0(a_20, b_7, h_s_arrmul24_and20_7_y0);
  fa fa_h_s_arrmul24_fa20_7_y2(h_s_arrmul24_and20_7_y0, h_s_arrmul24_fa21_6_y2, h_s_arrmul24_fa19_7_y4, h_s_arrmul24_fa20_7_y2, h_s_arrmul24_fa20_7_y4);
  and_gate and_gate_h_s_arrmul24_and21_7_y0(a_21, b_7, h_s_arrmul24_and21_7_y0);
  fa fa_h_s_arrmul24_fa21_7_y2(h_s_arrmul24_and21_7_y0, h_s_arrmul24_fa22_6_y2, h_s_arrmul24_fa20_7_y4, h_s_arrmul24_fa21_7_y2, h_s_arrmul24_fa21_7_y4);
  and_gate and_gate_h_s_arrmul24_and22_7_y0(a_22, b_7, h_s_arrmul24_and22_7_y0);
  fa fa_h_s_arrmul24_fa22_7_y2(h_s_arrmul24_and22_7_y0, h_s_arrmul24_fa23_6_y2, h_s_arrmul24_fa21_7_y4, h_s_arrmul24_fa22_7_y2, h_s_arrmul24_fa22_7_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_7_y0(a_23, b_7, h_s_arrmul24_nand23_7_y0);
  fa fa_h_s_arrmul24_fa23_7_y2(h_s_arrmul24_nand23_7_y0, h_s_arrmul24_fa23_6_y4, h_s_arrmul24_fa22_7_y4, h_s_arrmul24_fa23_7_y2, h_s_arrmul24_fa23_7_y4);
  and_gate and_gate_h_s_arrmul24_and0_8_y0(a_0, b_8, h_s_arrmul24_and0_8_y0);
  ha ha_h_s_arrmul24_ha0_8_y0(h_s_arrmul24_and0_8_y0, h_s_arrmul24_fa1_7_y2, h_s_arrmul24_ha0_8_y0, h_s_arrmul24_ha0_8_y1);
  and_gate and_gate_h_s_arrmul24_and1_8_y0(a_1, b_8, h_s_arrmul24_and1_8_y0);
  fa fa_h_s_arrmul24_fa1_8_y2(h_s_arrmul24_and1_8_y0, h_s_arrmul24_fa2_7_y2, h_s_arrmul24_ha0_8_y1, h_s_arrmul24_fa1_8_y2, h_s_arrmul24_fa1_8_y4);
  and_gate and_gate_h_s_arrmul24_and2_8_y0(a_2, b_8, h_s_arrmul24_and2_8_y0);
  fa fa_h_s_arrmul24_fa2_8_y2(h_s_arrmul24_and2_8_y0, h_s_arrmul24_fa3_7_y2, h_s_arrmul24_fa1_8_y4, h_s_arrmul24_fa2_8_y2, h_s_arrmul24_fa2_8_y4);
  and_gate and_gate_h_s_arrmul24_and3_8_y0(a_3, b_8, h_s_arrmul24_and3_8_y0);
  fa fa_h_s_arrmul24_fa3_8_y2(h_s_arrmul24_and3_8_y0, h_s_arrmul24_fa4_7_y2, h_s_arrmul24_fa2_8_y4, h_s_arrmul24_fa3_8_y2, h_s_arrmul24_fa3_8_y4);
  and_gate and_gate_h_s_arrmul24_and4_8_y0(a_4, b_8, h_s_arrmul24_and4_8_y0);
  fa fa_h_s_arrmul24_fa4_8_y2(h_s_arrmul24_and4_8_y0, h_s_arrmul24_fa5_7_y2, h_s_arrmul24_fa3_8_y4, h_s_arrmul24_fa4_8_y2, h_s_arrmul24_fa4_8_y4);
  and_gate and_gate_h_s_arrmul24_and5_8_y0(a_5, b_8, h_s_arrmul24_and5_8_y0);
  fa fa_h_s_arrmul24_fa5_8_y2(h_s_arrmul24_and5_8_y0, h_s_arrmul24_fa6_7_y2, h_s_arrmul24_fa4_8_y4, h_s_arrmul24_fa5_8_y2, h_s_arrmul24_fa5_8_y4);
  and_gate and_gate_h_s_arrmul24_and6_8_y0(a_6, b_8, h_s_arrmul24_and6_8_y0);
  fa fa_h_s_arrmul24_fa6_8_y2(h_s_arrmul24_and6_8_y0, h_s_arrmul24_fa7_7_y2, h_s_arrmul24_fa5_8_y4, h_s_arrmul24_fa6_8_y2, h_s_arrmul24_fa6_8_y4);
  and_gate and_gate_h_s_arrmul24_and7_8_y0(a_7, b_8, h_s_arrmul24_and7_8_y0);
  fa fa_h_s_arrmul24_fa7_8_y2(h_s_arrmul24_and7_8_y0, h_s_arrmul24_fa8_7_y2, h_s_arrmul24_fa6_8_y4, h_s_arrmul24_fa7_8_y2, h_s_arrmul24_fa7_8_y4);
  and_gate and_gate_h_s_arrmul24_and8_8_y0(a_8, b_8, h_s_arrmul24_and8_8_y0);
  fa fa_h_s_arrmul24_fa8_8_y2(h_s_arrmul24_and8_8_y0, h_s_arrmul24_fa9_7_y2, h_s_arrmul24_fa7_8_y4, h_s_arrmul24_fa8_8_y2, h_s_arrmul24_fa8_8_y4);
  and_gate and_gate_h_s_arrmul24_and9_8_y0(a_9, b_8, h_s_arrmul24_and9_8_y0);
  fa fa_h_s_arrmul24_fa9_8_y2(h_s_arrmul24_and9_8_y0, h_s_arrmul24_fa10_7_y2, h_s_arrmul24_fa8_8_y4, h_s_arrmul24_fa9_8_y2, h_s_arrmul24_fa9_8_y4);
  and_gate and_gate_h_s_arrmul24_and10_8_y0(a_10, b_8, h_s_arrmul24_and10_8_y0);
  fa fa_h_s_arrmul24_fa10_8_y2(h_s_arrmul24_and10_8_y0, h_s_arrmul24_fa11_7_y2, h_s_arrmul24_fa9_8_y4, h_s_arrmul24_fa10_8_y2, h_s_arrmul24_fa10_8_y4);
  and_gate and_gate_h_s_arrmul24_and11_8_y0(a_11, b_8, h_s_arrmul24_and11_8_y0);
  fa fa_h_s_arrmul24_fa11_8_y2(h_s_arrmul24_and11_8_y0, h_s_arrmul24_fa12_7_y2, h_s_arrmul24_fa10_8_y4, h_s_arrmul24_fa11_8_y2, h_s_arrmul24_fa11_8_y4);
  and_gate and_gate_h_s_arrmul24_and12_8_y0(a_12, b_8, h_s_arrmul24_and12_8_y0);
  fa fa_h_s_arrmul24_fa12_8_y2(h_s_arrmul24_and12_8_y0, h_s_arrmul24_fa13_7_y2, h_s_arrmul24_fa11_8_y4, h_s_arrmul24_fa12_8_y2, h_s_arrmul24_fa12_8_y4);
  and_gate and_gate_h_s_arrmul24_and13_8_y0(a_13, b_8, h_s_arrmul24_and13_8_y0);
  fa fa_h_s_arrmul24_fa13_8_y2(h_s_arrmul24_and13_8_y0, h_s_arrmul24_fa14_7_y2, h_s_arrmul24_fa12_8_y4, h_s_arrmul24_fa13_8_y2, h_s_arrmul24_fa13_8_y4);
  and_gate and_gate_h_s_arrmul24_and14_8_y0(a_14, b_8, h_s_arrmul24_and14_8_y0);
  fa fa_h_s_arrmul24_fa14_8_y2(h_s_arrmul24_and14_8_y0, h_s_arrmul24_fa15_7_y2, h_s_arrmul24_fa13_8_y4, h_s_arrmul24_fa14_8_y2, h_s_arrmul24_fa14_8_y4);
  and_gate and_gate_h_s_arrmul24_and15_8_y0(a_15, b_8, h_s_arrmul24_and15_8_y0);
  fa fa_h_s_arrmul24_fa15_8_y2(h_s_arrmul24_and15_8_y0, h_s_arrmul24_fa16_7_y2, h_s_arrmul24_fa14_8_y4, h_s_arrmul24_fa15_8_y2, h_s_arrmul24_fa15_8_y4);
  and_gate and_gate_h_s_arrmul24_and16_8_y0(a_16, b_8, h_s_arrmul24_and16_8_y0);
  fa fa_h_s_arrmul24_fa16_8_y2(h_s_arrmul24_and16_8_y0, h_s_arrmul24_fa17_7_y2, h_s_arrmul24_fa15_8_y4, h_s_arrmul24_fa16_8_y2, h_s_arrmul24_fa16_8_y4);
  and_gate and_gate_h_s_arrmul24_and17_8_y0(a_17, b_8, h_s_arrmul24_and17_8_y0);
  fa fa_h_s_arrmul24_fa17_8_y2(h_s_arrmul24_and17_8_y0, h_s_arrmul24_fa18_7_y2, h_s_arrmul24_fa16_8_y4, h_s_arrmul24_fa17_8_y2, h_s_arrmul24_fa17_8_y4);
  and_gate and_gate_h_s_arrmul24_and18_8_y0(a_18, b_8, h_s_arrmul24_and18_8_y0);
  fa fa_h_s_arrmul24_fa18_8_y2(h_s_arrmul24_and18_8_y0, h_s_arrmul24_fa19_7_y2, h_s_arrmul24_fa17_8_y4, h_s_arrmul24_fa18_8_y2, h_s_arrmul24_fa18_8_y4);
  and_gate and_gate_h_s_arrmul24_and19_8_y0(a_19, b_8, h_s_arrmul24_and19_8_y0);
  fa fa_h_s_arrmul24_fa19_8_y2(h_s_arrmul24_and19_8_y0, h_s_arrmul24_fa20_7_y2, h_s_arrmul24_fa18_8_y4, h_s_arrmul24_fa19_8_y2, h_s_arrmul24_fa19_8_y4);
  and_gate and_gate_h_s_arrmul24_and20_8_y0(a_20, b_8, h_s_arrmul24_and20_8_y0);
  fa fa_h_s_arrmul24_fa20_8_y2(h_s_arrmul24_and20_8_y0, h_s_arrmul24_fa21_7_y2, h_s_arrmul24_fa19_8_y4, h_s_arrmul24_fa20_8_y2, h_s_arrmul24_fa20_8_y4);
  and_gate and_gate_h_s_arrmul24_and21_8_y0(a_21, b_8, h_s_arrmul24_and21_8_y0);
  fa fa_h_s_arrmul24_fa21_8_y2(h_s_arrmul24_and21_8_y0, h_s_arrmul24_fa22_7_y2, h_s_arrmul24_fa20_8_y4, h_s_arrmul24_fa21_8_y2, h_s_arrmul24_fa21_8_y4);
  and_gate and_gate_h_s_arrmul24_and22_8_y0(a_22, b_8, h_s_arrmul24_and22_8_y0);
  fa fa_h_s_arrmul24_fa22_8_y2(h_s_arrmul24_and22_8_y0, h_s_arrmul24_fa23_7_y2, h_s_arrmul24_fa21_8_y4, h_s_arrmul24_fa22_8_y2, h_s_arrmul24_fa22_8_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_8_y0(a_23, b_8, h_s_arrmul24_nand23_8_y0);
  fa fa_h_s_arrmul24_fa23_8_y2(h_s_arrmul24_nand23_8_y0, h_s_arrmul24_fa23_7_y4, h_s_arrmul24_fa22_8_y4, h_s_arrmul24_fa23_8_y2, h_s_arrmul24_fa23_8_y4);
  and_gate and_gate_h_s_arrmul24_and0_9_y0(a_0, b_9, h_s_arrmul24_and0_9_y0);
  ha ha_h_s_arrmul24_ha0_9_y0(h_s_arrmul24_and0_9_y0, h_s_arrmul24_fa1_8_y2, h_s_arrmul24_ha0_9_y0, h_s_arrmul24_ha0_9_y1);
  and_gate and_gate_h_s_arrmul24_and1_9_y0(a_1, b_9, h_s_arrmul24_and1_9_y0);
  fa fa_h_s_arrmul24_fa1_9_y2(h_s_arrmul24_and1_9_y0, h_s_arrmul24_fa2_8_y2, h_s_arrmul24_ha0_9_y1, h_s_arrmul24_fa1_9_y2, h_s_arrmul24_fa1_9_y4);
  and_gate and_gate_h_s_arrmul24_and2_9_y0(a_2, b_9, h_s_arrmul24_and2_9_y0);
  fa fa_h_s_arrmul24_fa2_9_y2(h_s_arrmul24_and2_9_y0, h_s_arrmul24_fa3_8_y2, h_s_arrmul24_fa1_9_y4, h_s_arrmul24_fa2_9_y2, h_s_arrmul24_fa2_9_y4);
  and_gate and_gate_h_s_arrmul24_and3_9_y0(a_3, b_9, h_s_arrmul24_and3_9_y0);
  fa fa_h_s_arrmul24_fa3_9_y2(h_s_arrmul24_and3_9_y0, h_s_arrmul24_fa4_8_y2, h_s_arrmul24_fa2_9_y4, h_s_arrmul24_fa3_9_y2, h_s_arrmul24_fa3_9_y4);
  and_gate and_gate_h_s_arrmul24_and4_9_y0(a_4, b_9, h_s_arrmul24_and4_9_y0);
  fa fa_h_s_arrmul24_fa4_9_y2(h_s_arrmul24_and4_9_y0, h_s_arrmul24_fa5_8_y2, h_s_arrmul24_fa3_9_y4, h_s_arrmul24_fa4_9_y2, h_s_arrmul24_fa4_9_y4);
  and_gate and_gate_h_s_arrmul24_and5_9_y0(a_5, b_9, h_s_arrmul24_and5_9_y0);
  fa fa_h_s_arrmul24_fa5_9_y2(h_s_arrmul24_and5_9_y0, h_s_arrmul24_fa6_8_y2, h_s_arrmul24_fa4_9_y4, h_s_arrmul24_fa5_9_y2, h_s_arrmul24_fa5_9_y4);
  and_gate and_gate_h_s_arrmul24_and6_9_y0(a_6, b_9, h_s_arrmul24_and6_9_y0);
  fa fa_h_s_arrmul24_fa6_9_y2(h_s_arrmul24_and6_9_y0, h_s_arrmul24_fa7_8_y2, h_s_arrmul24_fa5_9_y4, h_s_arrmul24_fa6_9_y2, h_s_arrmul24_fa6_9_y4);
  and_gate and_gate_h_s_arrmul24_and7_9_y0(a_7, b_9, h_s_arrmul24_and7_9_y0);
  fa fa_h_s_arrmul24_fa7_9_y2(h_s_arrmul24_and7_9_y0, h_s_arrmul24_fa8_8_y2, h_s_arrmul24_fa6_9_y4, h_s_arrmul24_fa7_9_y2, h_s_arrmul24_fa7_9_y4);
  and_gate and_gate_h_s_arrmul24_and8_9_y0(a_8, b_9, h_s_arrmul24_and8_9_y0);
  fa fa_h_s_arrmul24_fa8_9_y2(h_s_arrmul24_and8_9_y0, h_s_arrmul24_fa9_8_y2, h_s_arrmul24_fa7_9_y4, h_s_arrmul24_fa8_9_y2, h_s_arrmul24_fa8_9_y4);
  and_gate and_gate_h_s_arrmul24_and9_9_y0(a_9, b_9, h_s_arrmul24_and9_9_y0);
  fa fa_h_s_arrmul24_fa9_9_y2(h_s_arrmul24_and9_9_y0, h_s_arrmul24_fa10_8_y2, h_s_arrmul24_fa8_9_y4, h_s_arrmul24_fa9_9_y2, h_s_arrmul24_fa9_9_y4);
  and_gate and_gate_h_s_arrmul24_and10_9_y0(a_10, b_9, h_s_arrmul24_and10_9_y0);
  fa fa_h_s_arrmul24_fa10_9_y2(h_s_arrmul24_and10_9_y0, h_s_arrmul24_fa11_8_y2, h_s_arrmul24_fa9_9_y4, h_s_arrmul24_fa10_9_y2, h_s_arrmul24_fa10_9_y4);
  and_gate and_gate_h_s_arrmul24_and11_9_y0(a_11, b_9, h_s_arrmul24_and11_9_y0);
  fa fa_h_s_arrmul24_fa11_9_y2(h_s_arrmul24_and11_9_y0, h_s_arrmul24_fa12_8_y2, h_s_arrmul24_fa10_9_y4, h_s_arrmul24_fa11_9_y2, h_s_arrmul24_fa11_9_y4);
  and_gate and_gate_h_s_arrmul24_and12_9_y0(a_12, b_9, h_s_arrmul24_and12_9_y0);
  fa fa_h_s_arrmul24_fa12_9_y2(h_s_arrmul24_and12_9_y0, h_s_arrmul24_fa13_8_y2, h_s_arrmul24_fa11_9_y4, h_s_arrmul24_fa12_9_y2, h_s_arrmul24_fa12_9_y4);
  and_gate and_gate_h_s_arrmul24_and13_9_y0(a_13, b_9, h_s_arrmul24_and13_9_y0);
  fa fa_h_s_arrmul24_fa13_9_y2(h_s_arrmul24_and13_9_y0, h_s_arrmul24_fa14_8_y2, h_s_arrmul24_fa12_9_y4, h_s_arrmul24_fa13_9_y2, h_s_arrmul24_fa13_9_y4);
  and_gate and_gate_h_s_arrmul24_and14_9_y0(a_14, b_9, h_s_arrmul24_and14_9_y0);
  fa fa_h_s_arrmul24_fa14_9_y2(h_s_arrmul24_and14_9_y0, h_s_arrmul24_fa15_8_y2, h_s_arrmul24_fa13_9_y4, h_s_arrmul24_fa14_9_y2, h_s_arrmul24_fa14_9_y4);
  and_gate and_gate_h_s_arrmul24_and15_9_y0(a_15, b_9, h_s_arrmul24_and15_9_y0);
  fa fa_h_s_arrmul24_fa15_9_y2(h_s_arrmul24_and15_9_y0, h_s_arrmul24_fa16_8_y2, h_s_arrmul24_fa14_9_y4, h_s_arrmul24_fa15_9_y2, h_s_arrmul24_fa15_9_y4);
  and_gate and_gate_h_s_arrmul24_and16_9_y0(a_16, b_9, h_s_arrmul24_and16_9_y0);
  fa fa_h_s_arrmul24_fa16_9_y2(h_s_arrmul24_and16_9_y0, h_s_arrmul24_fa17_8_y2, h_s_arrmul24_fa15_9_y4, h_s_arrmul24_fa16_9_y2, h_s_arrmul24_fa16_9_y4);
  and_gate and_gate_h_s_arrmul24_and17_9_y0(a_17, b_9, h_s_arrmul24_and17_9_y0);
  fa fa_h_s_arrmul24_fa17_9_y2(h_s_arrmul24_and17_9_y0, h_s_arrmul24_fa18_8_y2, h_s_arrmul24_fa16_9_y4, h_s_arrmul24_fa17_9_y2, h_s_arrmul24_fa17_9_y4);
  and_gate and_gate_h_s_arrmul24_and18_9_y0(a_18, b_9, h_s_arrmul24_and18_9_y0);
  fa fa_h_s_arrmul24_fa18_9_y2(h_s_arrmul24_and18_9_y0, h_s_arrmul24_fa19_8_y2, h_s_arrmul24_fa17_9_y4, h_s_arrmul24_fa18_9_y2, h_s_arrmul24_fa18_9_y4);
  and_gate and_gate_h_s_arrmul24_and19_9_y0(a_19, b_9, h_s_arrmul24_and19_9_y0);
  fa fa_h_s_arrmul24_fa19_9_y2(h_s_arrmul24_and19_9_y0, h_s_arrmul24_fa20_8_y2, h_s_arrmul24_fa18_9_y4, h_s_arrmul24_fa19_9_y2, h_s_arrmul24_fa19_9_y4);
  and_gate and_gate_h_s_arrmul24_and20_9_y0(a_20, b_9, h_s_arrmul24_and20_9_y0);
  fa fa_h_s_arrmul24_fa20_9_y2(h_s_arrmul24_and20_9_y0, h_s_arrmul24_fa21_8_y2, h_s_arrmul24_fa19_9_y4, h_s_arrmul24_fa20_9_y2, h_s_arrmul24_fa20_9_y4);
  and_gate and_gate_h_s_arrmul24_and21_9_y0(a_21, b_9, h_s_arrmul24_and21_9_y0);
  fa fa_h_s_arrmul24_fa21_9_y2(h_s_arrmul24_and21_9_y0, h_s_arrmul24_fa22_8_y2, h_s_arrmul24_fa20_9_y4, h_s_arrmul24_fa21_9_y2, h_s_arrmul24_fa21_9_y4);
  and_gate and_gate_h_s_arrmul24_and22_9_y0(a_22, b_9, h_s_arrmul24_and22_9_y0);
  fa fa_h_s_arrmul24_fa22_9_y2(h_s_arrmul24_and22_9_y0, h_s_arrmul24_fa23_8_y2, h_s_arrmul24_fa21_9_y4, h_s_arrmul24_fa22_9_y2, h_s_arrmul24_fa22_9_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_9_y0(a_23, b_9, h_s_arrmul24_nand23_9_y0);
  fa fa_h_s_arrmul24_fa23_9_y2(h_s_arrmul24_nand23_9_y0, h_s_arrmul24_fa23_8_y4, h_s_arrmul24_fa22_9_y4, h_s_arrmul24_fa23_9_y2, h_s_arrmul24_fa23_9_y4);
  and_gate and_gate_h_s_arrmul24_and0_10_y0(a_0, b_10, h_s_arrmul24_and0_10_y0);
  ha ha_h_s_arrmul24_ha0_10_y0(h_s_arrmul24_and0_10_y0, h_s_arrmul24_fa1_9_y2, h_s_arrmul24_ha0_10_y0, h_s_arrmul24_ha0_10_y1);
  and_gate and_gate_h_s_arrmul24_and1_10_y0(a_1, b_10, h_s_arrmul24_and1_10_y0);
  fa fa_h_s_arrmul24_fa1_10_y2(h_s_arrmul24_and1_10_y0, h_s_arrmul24_fa2_9_y2, h_s_arrmul24_ha0_10_y1, h_s_arrmul24_fa1_10_y2, h_s_arrmul24_fa1_10_y4);
  and_gate and_gate_h_s_arrmul24_and2_10_y0(a_2, b_10, h_s_arrmul24_and2_10_y0);
  fa fa_h_s_arrmul24_fa2_10_y2(h_s_arrmul24_and2_10_y0, h_s_arrmul24_fa3_9_y2, h_s_arrmul24_fa1_10_y4, h_s_arrmul24_fa2_10_y2, h_s_arrmul24_fa2_10_y4);
  and_gate and_gate_h_s_arrmul24_and3_10_y0(a_3, b_10, h_s_arrmul24_and3_10_y0);
  fa fa_h_s_arrmul24_fa3_10_y2(h_s_arrmul24_and3_10_y0, h_s_arrmul24_fa4_9_y2, h_s_arrmul24_fa2_10_y4, h_s_arrmul24_fa3_10_y2, h_s_arrmul24_fa3_10_y4);
  and_gate and_gate_h_s_arrmul24_and4_10_y0(a_4, b_10, h_s_arrmul24_and4_10_y0);
  fa fa_h_s_arrmul24_fa4_10_y2(h_s_arrmul24_and4_10_y0, h_s_arrmul24_fa5_9_y2, h_s_arrmul24_fa3_10_y4, h_s_arrmul24_fa4_10_y2, h_s_arrmul24_fa4_10_y4);
  and_gate and_gate_h_s_arrmul24_and5_10_y0(a_5, b_10, h_s_arrmul24_and5_10_y0);
  fa fa_h_s_arrmul24_fa5_10_y2(h_s_arrmul24_and5_10_y0, h_s_arrmul24_fa6_9_y2, h_s_arrmul24_fa4_10_y4, h_s_arrmul24_fa5_10_y2, h_s_arrmul24_fa5_10_y4);
  and_gate and_gate_h_s_arrmul24_and6_10_y0(a_6, b_10, h_s_arrmul24_and6_10_y0);
  fa fa_h_s_arrmul24_fa6_10_y2(h_s_arrmul24_and6_10_y0, h_s_arrmul24_fa7_9_y2, h_s_arrmul24_fa5_10_y4, h_s_arrmul24_fa6_10_y2, h_s_arrmul24_fa6_10_y4);
  and_gate and_gate_h_s_arrmul24_and7_10_y0(a_7, b_10, h_s_arrmul24_and7_10_y0);
  fa fa_h_s_arrmul24_fa7_10_y2(h_s_arrmul24_and7_10_y0, h_s_arrmul24_fa8_9_y2, h_s_arrmul24_fa6_10_y4, h_s_arrmul24_fa7_10_y2, h_s_arrmul24_fa7_10_y4);
  and_gate and_gate_h_s_arrmul24_and8_10_y0(a_8, b_10, h_s_arrmul24_and8_10_y0);
  fa fa_h_s_arrmul24_fa8_10_y2(h_s_arrmul24_and8_10_y0, h_s_arrmul24_fa9_9_y2, h_s_arrmul24_fa7_10_y4, h_s_arrmul24_fa8_10_y2, h_s_arrmul24_fa8_10_y4);
  and_gate and_gate_h_s_arrmul24_and9_10_y0(a_9, b_10, h_s_arrmul24_and9_10_y0);
  fa fa_h_s_arrmul24_fa9_10_y2(h_s_arrmul24_and9_10_y0, h_s_arrmul24_fa10_9_y2, h_s_arrmul24_fa8_10_y4, h_s_arrmul24_fa9_10_y2, h_s_arrmul24_fa9_10_y4);
  and_gate and_gate_h_s_arrmul24_and10_10_y0(a_10, b_10, h_s_arrmul24_and10_10_y0);
  fa fa_h_s_arrmul24_fa10_10_y2(h_s_arrmul24_and10_10_y0, h_s_arrmul24_fa11_9_y2, h_s_arrmul24_fa9_10_y4, h_s_arrmul24_fa10_10_y2, h_s_arrmul24_fa10_10_y4);
  and_gate and_gate_h_s_arrmul24_and11_10_y0(a_11, b_10, h_s_arrmul24_and11_10_y0);
  fa fa_h_s_arrmul24_fa11_10_y2(h_s_arrmul24_and11_10_y0, h_s_arrmul24_fa12_9_y2, h_s_arrmul24_fa10_10_y4, h_s_arrmul24_fa11_10_y2, h_s_arrmul24_fa11_10_y4);
  and_gate and_gate_h_s_arrmul24_and12_10_y0(a_12, b_10, h_s_arrmul24_and12_10_y0);
  fa fa_h_s_arrmul24_fa12_10_y2(h_s_arrmul24_and12_10_y0, h_s_arrmul24_fa13_9_y2, h_s_arrmul24_fa11_10_y4, h_s_arrmul24_fa12_10_y2, h_s_arrmul24_fa12_10_y4);
  and_gate and_gate_h_s_arrmul24_and13_10_y0(a_13, b_10, h_s_arrmul24_and13_10_y0);
  fa fa_h_s_arrmul24_fa13_10_y2(h_s_arrmul24_and13_10_y0, h_s_arrmul24_fa14_9_y2, h_s_arrmul24_fa12_10_y4, h_s_arrmul24_fa13_10_y2, h_s_arrmul24_fa13_10_y4);
  and_gate and_gate_h_s_arrmul24_and14_10_y0(a_14, b_10, h_s_arrmul24_and14_10_y0);
  fa fa_h_s_arrmul24_fa14_10_y2(h_s_arrmul24_and14_10_y0, h_s_arrmul24_fa15_9_y2, h_s_arrmul24_fa13_10_y4, h_s_arrmul24_fa14_10_y2, h_s_arrmul24_fa14_10_y4);
  and_gate and_gate_h_s_arrmul24_and15_10_y0(a_15, b_10, h_s_arrmul24_and15_10_y0);
  fa fa_h_s_arrmul24_fa15_10_y2(h_s_arrmul24_and15_10_y0, h_s_arrmul24_fa16_9_y2, h_s_arrmul24_fa14_10_y4, h_s_arrmul24_fa15_10_y2, h_s_arrmul24_fa15_10_y4);
  and_gate and_gate_h_s_arrmul24_and16_10_y0(a_16, b_10, h_s_arrmul24_and16_10_y0);
  fa fa_h_s_arrmul24_fa16_10_y2(h_s_arrmul24_and16_10_y0, h_s_arrmul24_fa17_9_y2, h_s_arrmul24_fa15_10_y4, h_s_arrmul24_fa16_10_y2, h_s_arrmul24_fa16_10_y4);
  and_gate and_gate_h_s_arrmul24_and17_10_y0(a_17, b_10, h_s_arrmul24_and17_10_y0);
  fa fa_h_s_arrmul24_fa17_10_y2(h_s_arrmul24_and17_10_y0, h_s_arrmul24_fa18_9_y2, h_s_arrmul24_fa16_10_y4, h_s_arrmul24_fa17_10_y2, h_s_arrmul24_fa17_10_y4);
  and_gate and_gate_h_s_arrmul24_and18_10_y0(a_18, b_10, h_s_arrmul24_and18_10_y0);
  fa fa_h_s_arrmul24_fa18_10_y2(h_s_arrmul24_and18_10_y0, h_s_arrmul24_fa19_9_y2, h_s_arrmul24_fa17_10_y4, h_s_arrmul24_fa18_10_y2, h_s_arrmul24_fa18_10_y4);
  and_gate and_gate_h_s_arrmul24_and19_10_y0(a_19, b_10, h_s_arrmul24_and19_10_y0);
  fa fa_h_s_arrmul24_fa19_10_y2(h_s_arrmul24_and19_10_y0, h_s_arrmul24_fa20_9_y2, h_s_arrmul24_fa18_10_y4, h_s_arrmul24_fa19_10_y2, h_s_arrmul24_fa19_10_y4);
  and_gate and_gate_h_s_arrmul24_and20_10_y0(a_20, b_10, h_s_arrmul24_and20_10_y0);
  fa fa_h_s_arrmul24_fa20_10_y2(h_s_arrmul24_and20_10_y0, h_s_arrmul24_fa21_9_y2, h_s_arrmul24_fa19_10_y4, h_s_arrmul24_fa20_10_y2, h_s_arrmul24_fa20_10_y4);
  and_gate and_gate_h_s_arrmul24_and21_10_y0(a_21, b_10, h_s_arrmul24_and21_10_y0);
  fa fa_h_s_arrmul24_fa21_10_y2(h_s_arrmul24_and21_10_y0, h_s_arrmul24_fa22_9_y2, h_s_arrmul24_fa20_10_y4, h_s_arrmul24_fa21_10_y2, h_s_arrmul24_fa21_10_y4);
  and_gate and_gate_h_s_arrmul24_and22_10_y0(a_22, b_10, h_s_arrmul24_and22_10_y0);
  fa fa_h_s_arrmul24_fa22_10_y2(h_s_arrmul24_and22_10_y0, h_s_arrmul24_fa23_9_y2, h_s_arrmul24_fa21_10_y4, h_s_arrmul24_fa22_10_y2, h_s_arrmul24_fa22_10_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_10_y0(a_23, b_10, h_s_arrmul24_nand23_10_y0);
  fa fa_h_s_arrmul24_fa23_10_y2(h_s_arrmul24_nand23_10_y0, h_s_arrmul24_fa23_9_y4, h_s_arrmul24_fa22_10_y4, h_s_arrmul24_fa23_10_y2, h_s_arrmul24_fa23_10_y4);
  and_gate and_gate_h_s_arrmul24_and0_11_y0(a_0, b_11, h_s_arrmul24_and0_11_y0);
  ha ha_h_s_arrmul24_ha0_11_y0(h_s_arrmul24_and0_11_y0, h_s_arrmul24_fa1_10_y2, h_s_arrmul24_ha0_11_y0, h_s_arrmul24_ha0_11_y1);
  and_gate and_gate_h_s_arrmul24_and1_11_y0(a_1, b_11, h_s_arrmul24_and1_11_y0);
  fa fa_h_s_arrmul24_fa1_11_y2(h_s_arrmul24_and1_11_y0, h_s_arrmul24_fa2_10_y2, h_s_arrmul24_ha0_11_y1, h_s_arrmul24_fa1_11_y2, h_s_arrmul24_fa1_11_y4);
  and_gate and_gate_h_s_arrmul24_and2_11_y0(a_2, b_11, h_s_arrmul24_and2_11_y0);
  fa fa_h_s_arrmul24_fa2_11_y2(h_s_arrmul24_and2_11_y0, h_s_arrmul24_fa3_10_y2, h_s_arrmul24_fa1_11_y4, h_s_arrmul24_fa2_11_y2, h_s_arrmul24_fa2_11_y4);
  and_gate and_gate_h_s_arrmul24_and3_11_y0(a_3, b_11, h_s_arrmul24_and3_11_y0);
  fa fa_h_s_arrmul24_fa3_11_y2(h_s_arrmul24_and3_11_y0, h_s_arrmul24_fa4_10_y2, h_s_arrmul24_fa2_11_y4, h_s_arrmul24_fa3_11_y2, h_s_arrmul24_fa3_11_y4);
  and_gate and_gate_h_s_arrmul24_and4_11_y0(a_4, b_11, h_s_arrmul24_and4_11_y0);
  fa fa_h_s_arrmul24_fa4_11_y2(h_s_arrmul24_and4_11_y0, h_s_arrmul24_fa5_10_y2, h_s_arrmul24_fa3_11_y4, h_s_arrmul24_fa4_11_y2, h_s_arrmul24_fa4_11_y4);
  and_gate and_gate_h_s_arrmul24_and5_11_y0(a_5, b_11, h_s_arrmul24_and5_11_y0);
  fa fa_h_s_arrmul24_fa5_11_y2(h_s_arrmul24_and5_11_y0, h_s_arrmul24_fa6_10_y2, h_s_arrmul24_fa4_11_y4, h_s_arrmul24_fa5_11_y2, h_s_arrmul24_fa5_11_y4);
  and_gate and_gate_h_s_arrmul24_and6_11_y0(a_6, b_11, h_s_arrmul24_and6_11_y0);
  fa fa_h_s_arrmul24_fa6_11_y2(h_s_arrmul24_and6_11_y0, h_s_arrmul24_fa7_10_y2, h_s_arrmul24_fa5_11_y4, h_s_arrmul24_fa6_11_y2, h_s_arrmul24_fa6_11_y4);
  and_gate and_gate_h_s_arrmul24_and7_11_y0(a_7, b_11, h_s_arrmul24_and7_11_y0);
  fa fa_h_s_arrmul24_fa7_11_y2(h_s_arrmul24_and7_11_y0, h_s_arrmul24_fa8_10_y2, h_s_arrmul24_fa6_11_y4, h_s_arrmul24_fa7_11_y2, h_s_arrmul24_fa7_11_y4);
  and_gate and_gate_h_s_arrmul24_and8_11_y0(a_8, b_11, h_s_arrmul24_and8_11_y0);
  fa fa_h_s_arrmul24_fa8_11_y2(h_s_arrmul24_and8_11_y0, h_s_arrmul24_fa9_10_y2, h_s_arrmul24_fa7_11_y4, h_s_arrmul24_fa8_11_y2, h_s_arrmul24_fa8_11_y4);
  and_gate and_gate_h_s_arrmul24_and9_11_y0(a_9, b_11, h_s_arrmul24_and9_11_y0);
  fa fa_h_s_arrmul24_fa9_11_y2(h_s_arrmul24_and9_11_y0, h_s_arrmul24_fa10_10_y2, h_s_arrmul24_fa8_11_y4, h_s_arrmul24_fa9_11_y2, h_s_arrmul24_fa9_11_y4);
  and_gate and_gate_h_s_arrmul24_and10_11_y0(a_10, b_11, h_s_arrmul24_and10_11_y0);
  fa fa_h_s_arrmul24_fa10_11_y2(h_s_arrmul24_and10_11_y0, h_s_arrmul24_fa11_10_y2, h_s_arrmul24_fa9_11_y4, h_s_arrmul24_fa10_11_y2, h_s_arrmul24_fa10_11_y4);
  and_gate and_gate_h_s_arrmul24_and11_11_y0(a_11, b_11, h_s_arrmul24_and11_11_y0);
  fa fa_h_s_arrmul24_fa11_11_y2(h_s_arrmul24_and11_11_y0, h_s_arrmul24_fa12_10_y2, h_s_arrmul24_fa10_11_y4, h_s_arrmul24_fa11_11_y2, h_s_arrmul24_fa11_11_y4);
  and_gate and_gate_h_s_arrmul24_and12_11_y0(a_12, b_11, h_s_arrmul24_and12_11_y0);
  fa fa_h_s_arrmul24_fa12_11_y2(h_s_arrmul24_and12_11_y0, h_s_arrmul24_fa13_10_y2, h_s_arrmul24_fa11_11_y4, h_s_arrmul24_fa12_11_y2, h_s_arrmul24_fa12_11_y4);
  and_gate and_gate_h_s_arrmul24_and13_11_y0(a_13, b_11, h_s_arrmul24_and13_11_y0);
  fa fa_h_s_arrmul24_fa13_11_y2(h_s_arrmul24_and13_11_y0, h_s_arrmul24_fa14_10_y2, h_s_arrmul24_fa12_11_y4, h_s_arrmul24_fa13_11_y2, h_s_arrmul24_fa13_11_y4);
  and_gate and_gate_h_s_arrmul24_and14_11_y0(a_14, b_11, h_s_arrmul24_and14_11_y0);
  fa fa_h_s_arrmul24_fa14_11_y2(h_s_arrmul24_and14_11_y0, h_s_arrmul24_fa15_10_y2, h_s_arrmul24_fa13_11_y4, h_s_arrmul24_fa14_11_y2, h_s_arrmul24_fa14_11_y4);
  and_gate and_gate_h_s_arrmul24_and15_11_y0(a_15, b_11, h_s_arrmul24_and15_11_y0);
  fa fa_h_s_arrmul24_fa15_11_y2(h_s_arrmul24_and15_11_y0, h_s_arrmul24_fa16_10_y2, h_s_arrmul24_fa14_11_y4, h_s_arrmul24_fa15_11_y2, h_s_arrmul24_fa15_11_y4);
  and_gate and_gate_h_s_arrmul24_and16_11_y0(a_16, b_11, h_s_arrmul24_and16_11_y0);
  fa fa_h_s_arrmul24_fa16_11_y2(h_s_arrmul24_and16_11_y0, h_s_arrmul24_fa17_10_y2, h_s_arrmul24_fa15_11_y4, h_s_arrmul24_fa16_11_y2, h_s_arrmul24_fa16_11_y4);
  and_gate and_gate_h_s_arrmul24_and17_11_y0(a_17, b_11, h_s_arrmul24_and17_11_y0);
  fa fa_h_s_arrmul24_fa17_11_y2(h_s_arrmul24_and17_11_y0, h_s_arrmul24_fa18_10_y2, h_s_arrmul24_fa16_11_y4, h_s_arrmul24_fa17_11_y2, h_s_arrmul24_fa17_11_y4);
  and_gate and_gate_h_s_arrmul24_and18_11_y0(a_18, b_11, h_s_arrmul24_and18_11_y0);
  fa fa_h_s_arrmul24_fa18_11_y2(h_s_arrmul24_and18_11_y0, h_s_arrmul24_fa19_10_y2, h_s_arrmul24_fa17_11_y4, h_s_arrmul24_fa18_11_y2, h_s_arrmul24_fa18_11_y4);
  and_gate and_gate_h_s_arrmul24_and19_11_y0(a_19, b_11, h_s_arrmul24_and19_11_y0);
  fa fa_h_s_arrmul24_fa19_11_y2(h_s_arrmul24_and19_11_y0, h_s_arrmul24_fa20_10_y2, h_s_arrmul24_fa18_11_y4, h_s_arrmul24_fa19_11_y2, h_s_arrmul24_fa19_11_y4);
  and_gate and_gate_h_s_arrmul24_and20_11_y0(a_20, b_11, h_s_arrmul24_and20_11_y0);
  fa fa_h_s_arrmul24_fa20_11_y2(h_s_arrmul24_and20_11_y0, h_s_arrmul24_fa21_10_y2, h_s_arrmul24_fa19_11_y4, h_s_arrmul24_fa20_11_y2, h_s_arrmul24_fa20_11_y4);
  and_gate and_gate_h_s_arrmul24_and21_11_y0(a_21, b_11, h_s_arrmul24_and21_11_y0);
  fa fa_h_s_arrmul24_fa21_11_y2(h_s_arrmul24_and21_11_y0, h_s_arrmul24_fa22_10_y2, h_s_arrmul24_fa20_11_y4, h_s_arrmul24_fa21_11_y2, h_s_arrmul24_fa21_11_y4);
  and_gate and_gate_h_s_arrmul24_and22_11_y0(a_22, b_11, h_s_arrmul24_and22_11_y0);
  fa fa_h_s_arrmul24_fa22_11_y2(h_s_arrmul24_and22_11_y0, h_s_arrmul24_fa23_10_y2, h_s_arrmul24_fa21_11_y4, h_s_arrmul24_fa22_11_y2, h_s_arrmul24_fa22_11_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_11_y0(a_23, b_11, h_s_arrmul24_nand23_11_y0);
  fa fa_h_s_arrmul24_fa23_11_y2(h_s_arrmul24_nand23_11_y0, h_s_arrmul24_fa23_10_y4, h_s_arrmul24_fa22_11_y4, h_s_arrmul24_fa23_11_y2, h_s_arrmul24_fa23_11_y4);
  and_gate and_gate_h_s_arrmul24_and0_12_y0(a_0, b_12, h_s_arrmul24_and0_12_y0);
  ha ha_h_s_arrmul24_ha0_12_y0(h_s_arrmul24_and0_12_y0, h_s_arrmul24_fa1_11_y2, h_s_arrmul24_ha0_12_y0, h_s_arrmul24_ha0_12_y1);
  and_gate and_gate_h_s_arrmul24_and1_12_y0(a_1, b_12, h_s_arrmul24_and1_12_y0);
  fa fa_h_s_arrmul24_fa1_12_y2(h_s_arrmul24_and1_12_y0, h_s_arrmul24_fa2_11_y2, h_s_arrmul24_ha0_12_y1, h_s_arrmul24_fa1_12_y2, h_s_arrmul24_fa1_12_y4);
  and_gate and_gate_h_s_arrmul24_and2_12_y0(a_2, b_12, h_s_arrmul24_and2_12_y0);
  fa fa_h_s_arrmul24_fa2_12_y2(h_s_arrmul24_and2_12_y0, h_s_arrmul24_fa3_11_y2, h_s_arrmul24_fa1_12_y4, h_s_arrmul24_fa2_12_y2, h_s_arrmul24_fa2_12_y4);
  and_gate and_gate_h_s_arrmul24_and3_12_y0(a_3, b_12, h_s_arrmul24_and3_12_y0);
  fa fa_h_s_arrmul24_fa3_12_y2(h_s_arrmul24_and3_12_y0, h_s_arrmul24_fa4_11_y2, h_s_arrmul24_fa2_12_y4, h_s_arrmul24_fa3_12_y2, h_s_arrmul24_fa3_12_y4);
  and_gate and_gate_h_s_arrmul24_and4_12_y0(a_4, b_12, h_s_arrmul24_and4_12_y0);
  fa fa_h_s_arrmul24_fa4_12_y2(h_s_arrmul24_and4_12_y0, h_s_arrmul24_fa5_11_y2, h_s_arrmul24_fa3_12_y4, h_s_arrmul24_fa4_12_y2, h_s_arrmul24_fa4_12_y4);
  and_gate and_gate_h_s_arrmul24_and5_12_y0(a_5, b_12, h_s_arrmul24_and5_12_y0);
  fa fa_h_s_arrmul24_fa5_12_y2(h_s_arrmul24_and5_12_y0, h_s_arrmul24_fa6_11_y2, h_s_arrmul24_fa4_12_y4, h_s_arrmul24_fa5_12_y2, h_s_arrmul24_fa5_12_y4);
  and_gate and_gate_h_s_arrmul24_and6_12_y0(a_6, b_12, h_s_arrmul24_and6_12_y0);
  fa fa_h_s_arrmul24_fa6_12_y2(h_s_arrmul24_and6_12_y0, h_s_arrmul24_fa7_11_y2, h_s_arrmul24_fa5_12_y4, h_s_arrmul24_fa6_12_y2, h_s_arrmul24_fa6_12_y4);
  and_gate and_gate_h_s_arrmul24_and7_12_y0(a_7, b_12, h_s_arrmul24_and7_12_y0);
  fa fa_h_s_arrmul24_fa7_12_y2(h_s_arrmul24_and7_12_y0, h_s_arrmul24_fa8_11_y2, h_s_arrmul24_fa6_12_y4, h_s_arrmul24_fa7_12_y2, h_s_arrmul24_fa7_12_y4);
  and_gate and_gate_h_s_arrmul24_and8_12_y0(a_8, b_12, h_s_arrmul24_and8_12_y0);
  fa fa_h_s_arrmul24_fa8_12_y2(h_s_arrmul24_and8_12_y0, h_s_arrmul24_fa9_11_y2, h_s_arrmul24_fa7_12_y4, h_s_arrmul24_fa8_12_y2, h_s_arrmul24_fa8_12_y4);
  and_gate and_gate_h_s_arrmul24_and9_12_y0(a_9, b_12, h_s_arrmul24_and9_12_y0);
  fa fa_h_s_arrmul24_fa9_12_y2(h_s_arrmul24_and9_12_y0, h_s_arrmul24_fa10_11_y2, h_s_arrmul24_fa8_12_y4, h_s_arrmul24_fa9_12_y2, h_s_arrmul24_fa9_12_y4);
  and_gate and_gate_h_s_arrmul24_and10_12_y0(a_10, b_12, h_s_arrmul24_and10_12_y0);
  fa fa_h_s_arrmul24_fa10_12_y2(h_s_arrmul24_and10_12_y0, h_s_arrmul24_fa11_11_y2, h_s_arrmul24_fa9_12_y4, h_s_arrmul24_fa10_12_y2, h_s_arrmul24_fa10_12_y4);
  and_gate and_gate_h_s_arrmul24_and11_12_y0(a_11, b_12, h_s_arrmul24_and11_12_y0);
  fa fa_h_s_arrmul24_fa11_12_y2(h_s_arrmul24_and11_12_y0, h_s_arrmul24_fa12_11_y2, h_s_arrmul24_fa10_12_y4, h_s_arrmul24_fa11_12_y2, h_s_arrmul24_fa11_12_y4);
  and_gate and_gate_h_s_arrmul24_and12_12_y0(a_12, b_12, h_s_arrmul24_and12_12_y0);
  fa fa_h_s_arrmul24_fa12_12_y2(h_s_arrmul24_and12_12_y0, h_s_arrmul24_fa13_11_y2, h_s_arrmul24_fa11_12_y4, h_s_arrmul24_fa12_12_y2, h_s_arrmul24_fa12_12_y4);
  and_gate and_gate_h_s_arrmul24_and13_12_y0(a_13, b_12, h_s_arrmul24_and13_12_y0);
  fa fa_h_s_arrmul24_fa13_12_y2(h_s_arrmul24_and13_12_y0, h_s_arrmul24_fa14_11_y2, h_s_arrmul24_fa12_12_y4, h_s_arrmul24_fa13_12_y2, h_s_arrmul24_fa13_12_y4);
  and_gate and_gate_h_s_arrmul24_and14_12_y0(a_14, b_12, h_s_arrmul24_and14_12_y0);
  fa fa_h_s_arrmul24_fa14_12_y2(h_s_arrmul24_and14_12_y0, h_s_arrmul24_fa15_11_y2, h_s_arrmul24_fa13_12_y4, h_s_arrmul24_fa14_12_y2, h_s_arrmul24_fa14_12_y4);
  and_gate and_gate_h_s_arrmul24_and15_12_y0(a_15, b_12, h_s_arrmul24_and15_12_y0);
  fa fa_h_s_arrmul24_fa15_12_y2(h_s_arrmul24_and15_12_y0, h_s_arrmul24_fa16_11_y2, h_s_arrmul24_fa14_12_y4, h_s_arrmul24_fa15_12_y2, h_s_arrmul24_fa15_12_y4);
  and_gate and_gate_h_s_arrmul24_and16_12_y0(a_16, b_12, h_s_arrmul24_and16_12_y0);
  fa fa_h_s_arrmul24_fa16_12_y2(h_s_arrmul24_and16_12_y0, h_s_arrmul24_fa17_11_y2, h_s_arrmul24_fa15_12_y4, h_s_arrmul24_fa16_12_y2, h_s_arrmul24_fa16_12_y4);
  and_gate and_gate_h_s_arrmul24_and17_12_y0(a_17, b_12, h_s_arrmul24_and17_12_y0);
  fa fa_h_s_arrmul24_fa17_12_y2(h_s_arrmul24_and17_12_y0, h_s_arrmul24_fa18_11_y2, h_s_arrmul24_fa16_12_y4, h_s_arrmul24_fa17_12_y2, h_s_arrmul24_fa17_12_y4);
  and_gate and_gate_h_s_arrmul24_and18_12_y0(a_18, b_12, h_s_arrmul24_and18_12_y0);
  fa fa_h_s_arrmul24_fa18_12_y2(h_s_arrmul24_and18_12_y0, h_s_arrmul24_fa19_11_y2, h_s_arrmul24_fa17_12_y4, h_s_arrmul24_fa18_12_y2, h_s_arrmul24_fa18_12_y4);
  and_gate and_gate_h_s_arrmul24_and19_12_y0(a_19, b_12, h_s_arrmul24_and19_12_y0);
  fa fa_h_s_arrmul24_fa19_12_y2(h_s_arrmul24_and19_12_y0, h_s_arrmul24_fa20_11_y2, h_s_arrmul24_fa18_12_y4, h_s_arrmul24_fa19_12_y2, h_s_arrmul24_fa19_12_y4);
  and_gate and_gate_h_s_arrmul24_and20_12_y0(a_20, b_12, h_s_arrmul24_and20_12_y0);
  fa fa_h_s_arrmul24_fa20_12_y2(h_s_arrmul24_and20_12_y0, h_s_arrmul24_fa21_11_y2, h_s_arrmul24_fa19_12_y4, h_s_arrmul24_fa20_12_y2, h_s_arrmul24_fa20_12_y4);
  and_gate and_gate_h_s_arrmul24_and21_12_y0(a_21, b_12, h_s_arrmul24_and21_12_y0);
  fa fa_h_s_arrmul24_fa21_12_y2(h_s_arrmul24_and21_12_y0, h_s_arrmul24_fa22_11_y2, h_s_arrmul24_fa20_12_y4, h_s_arrmul24_fa21_12_y2, h_s_arrmul24_fa21_12_y4);
  and_gate and_gate_h_s_arrmul24_and22_12_y0(a_22, b_12, h_s_arrmul24_and22_12_y0);
  fa fa_h_s_arrmul24_fa22_12_y2(h_s_arrmul24_and22_12_y0, h_s_arrmul24_fa23_11_y2, h_s_arrmul24_fa21_12_y4, h_s_arrmul24_fa22_12_y2, h_s_arrmul24_fa22_12_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_12_y0(a_23, b_12, h_s_arrmul24_nand23_12_y0);
  fa fa_h_s_arrmul24_fa23_12_y2(h_s_arrmul24_nand23_12_y0, h_s_arrmul24_fa23_11_y4, h_s_arrmul24_fa22_12_y4, h_s_arrmul24_fa23_12_y2, h_s_arrmul24_fa23_12_y4);
  and_gate and_gate_h_s_arrmul24_and0_13_y0(a_0, b_13, h_s_arrmul24_and0_13_y0);
  ha ha_h_s_arrmul24_ha0_13_y0(h_s_arrmul24_and0_13_y0, h_s_arrmul24_fa1_12_y2, h_s_arrmul24_ha0_13_y0, h_s_arrmul24_ha0_13_y1);
  and_gate and_gate_h_s_arrmul24_and1_13_y0(a_1, b_13, h_s_arrmul24_and1_13_y0);
  fa fa_h_s_arrmul24_fa1_13_y2(h_s_arrmul24_and1_13_y0, h_s_arrmul24_fa2_12_y2, h_s_arrmul24_ha0_13_y1, h_s_arrmul24_fa1_13_y2, h_s_arrmul24_fa1_13_y4);
  and_gate and_gate_h_s_arrmul24_and2_13_y0(a_2, b_13, h_s_arrmul24_and2_13_y0);
  fa fa_h_s_arrmul24_fa2_13_y2(h_s_arrmul24_and2_13_y0, h_s_arrmul24_fa3_12_y2, h_s_arrmul24_fa1_13_y4, h_s_arrmul24_fa2_13_y2, h_s_arrmul24_fa2_13_y4);
  and_gate and_gate_h_s_arrmul24_and3_13_y0(a_3, b_13, h_s_arrmul24_and3_13_y0);
  fa fa_h_s_arrmul24_fa3_13_y2(h_s_arrmul24_and3_13_y0, h_s_arrmul24_fa4_12_y2, h_s_arrmul24_fa2_13_y4, h_s_arrmul24_fa3_13_y2, h_s_arrmul24_fa3_13_y4);
  and_gate and_gate_h_s_arrmul24_and4_13_y0(a_4, b_13, h_s_arrmul24_and4_13_y0);
  fa fa_h_s_arrmul24_fa4_13_y2(h_s_arrmul24_and4_13_y0, h_s_arrmul24_fa5_12_y2, h_s_arrmul24_fa3_13_y4, h_s_arrmul24_fa4_13_y2, h_s_arrmul24_fa4_13_y4);
  and_gate and_gate_h_s_arrmul24_and5_13_y0(a_5, b_13, h_s_arrmul24_and5_13_y0);
  fa fa_h_s_arrmul24_fa5_13_y2(h_s_arrmul24_and5_13_y0, h_s_arrmul24_fa6_12_y2, h_s_arrmul24_fa4_13_y4, h_s_arrmul24_fa5_13_y2, h_s_arrmul24_fa5_13_y4);
  and_gate and_gate_h_s_arrmul24_and6_13_y0(a_6, b_13, h_s_arrmul24_and6_13_y0);
  fa fa_h_s_arrmul24_fa6_13_y2(h_s_arrmul24_and6_13_y0, h_s_arrmul24_fa7_12_y2, h_s_arrmul24_fa5_13_y4, h_s_arrmul24_fa6_13_y2, h_s_arrmul24_fa6_13_y4);
  and_gate and_gate_h_s_arrmul24_and7_13_y0(a_7, b_13, h_s_arrmul24_and7_13_y0);
  fa fa_h_s_arrmul24_fa7_13_y2(h_s_arrmul24_and7_13_y0, h_s_arrmul24_fa8_12_y2, h_s_arrmul24_fa6_13_y4, h_s_arrmul24_fa7_13_y2, h_s_arrmul24_fa7_13_y4);
  and_gate and_gate_h_s_arrmul24_and8_13_y0(a_8, b_13, h_s_arrmul24_and8_13_y0);
  fa fa_h_s_arrmul24_fa8_13_y2(h_s_arrmul24_and8_13_y0, h_s_arrmul24_fa9_12_y2, h_s_arrmul24_fa7_13_y4, h_s_arrmul24_fa8_13_y2, h_s_arrmul24_fa8_13_y4);
  and_gate and_gate_h_s_arrmul24_and9_13_y0(a_9, b_13, h_s_arrmul24_and9_13_y0);
  fa fa_h_s_arrmul24_fa9_13_y2(h_s_arrmul24_and9_13_y0, h_s_arrmul24_fa10_12_y2, h_s_arrmul24_fa8_13_y4, h_s_arrmul24_fa9_13_y2, h_s_arrmul24_fa9_13_y4);
  and_gate and_gate_h_s_arrmul24_and10_13_y0(a_10, b_13, h_s_arrmul24_and10_13_y0);
  fa fa_h_s_arrmul24_fa10_13_y2(h_s_arrmul24_and10_13_y0, h_s_arrmul24_fa11_12_y2, h_s_arrmul24_fa9_13_y4, h_s_arrmul24_fa10_13_y2, h_s_arrmul24_fa10_13_y4);
  and_gate and_gate_h_s_arrmul24_and11_13_y0(a_11, b_13, h_s_arrmul24_and11_13_y0);
  fa fa_h_s_arrmul24_fa11_13_y2(h_s_arrmul24_and11_13_y0, h_s_arrmul24_fa12_12_y2, h_s_arrmul24_fa10_13_y4, h_s_arrmul24_fa11_13_y2, h_s_arrmul24_fa11_13_y4);
  and_gate and_gate_h_s_arrmul24_and12_13_y0(a_12, b_13, h_s_arrmul24_and12_13_y0);
  fa fa_h_s_arrmul24_fa12_13_y2(h_s_arrmul24_and12_13_y0, h_s_arrmul24_fa13_12_y2, h_s_arrmul24_fa11_13_y4, h_s_arrmul24_fa12_13_y2, h_s_arrmul24_fa12_13_y4);
  and_gate and_gate_h_s_arrmul24_and13_13_y0(a_13, b_13, h_s_arrmul24_and13_13_y0);
  fa fa_h_s_arrmul24_fa13_13_y2(h_s_arrmul24_and13_13_y0, h_s_arrmul24_fa14_12_y2, h_s_arrmul24_fa12_13_y4, h_s_arrmul24_fa13_13_y2, h_s_arrmul24_fa13_13_y4);
  and_gate and_gate_h_s_arrmul24_and14_13_y0(a_14, b_13, h_s_arrmul24_and14_13_y0);
  fa fa_h_s_arrmul24_fa14_13_y2(h_s_arrmul24_and14_13_y0, h_s_arrmul24_fa15_12_y2, h_s_arrmul24_fa13_13_y4, h_s_arrmul24_fa14_13_y2, h_s_arrmul24_fa14_13_y4);
  and_gate and_gate_h_s_arrmul24_and15_13_y0(a_15, b_13, h_s_arrmul24_and15_13_y0);
  fa fa_h_s_arrmul24_fa15_13_y2(h_s_arrmul24_and15_13_y0, h_s_arrmul24_fa16_12_y2, h_s_arrmul24_fa14_13_y4, h_s_arrmul24_fa15_13_y2, h_s_arrmul24_fa15_13_y4);
  and_gate and_gate_h_s_arrmul24_and16_13_y0(a_16, b_13, h_s_arrmul24_and16_13_y0);
  fa fa_h_s_arrmul24_fa16_13_y2(h_s_arrmul24_and16_13_y0, h_s_arrmul24_fa17_12_y2, h_s_arrmul24_fa15_13_y4, h_s_arrmul24_fa16_13_y2, h_s_arrmul24_fa16_13_y4);
  and_gate and_gate_h_s_arrmul24_and17_13_y0(a_17, b_13, h_s_arrmul24_and17_13_y0);
  fa fa_h_s_arrmul24_fa17_13_y2(h_s_arrmul24_and17_13_y0, h_s_arrmul24_fa18_12_y2, h_s_arrmul24_fa16_13_y4, h_s_arrmul24_fa17_13_y2, h_s_arrmul24_fa17_13_y4);
  and_gate and_gate_h_s_arrmul24_and18_13_y0(a_18, b_13, h_s_arrmul24_and18_13_y0);
  fa fa_h_s_arrmul24_fa18_13_y2(h_s_arrmul24_and18_13_y0, h_s_arrmul24_fa19_12_y2, h_s_arrmul24_fa17_13_y4, h_s_arrmul24_fa18_13_y2, h_s_arrmul24_fa18_13_y4);
  and_gate and_gate_h_s_arrmul24_and19_13_y0(a_19, b_13, h_s_arrmul24_and19_13_y0);
  fa fa_h_s_arrmul24_fa19_13_y2(h_s_arrmul24_and19_13_y0, h_s_arrmul24_fa20_12_y2, h_s_arrmul24_fa18_13_y4, h_s_arrmul24_fa19_13_y2, h_s_arrmul24_fa19_13_y4);
  and_gate and_gate_h_s_arrmul24_and20_13_y0(a_20, b_13, h_s_arrmul24_and20_13_y0);
  fa fa_h_s_arrmul24_fa20_13_y2(h_s_arrmul24_and20_13_y0, h_s_arrmul24_fa21_12_y2, h_s_arrmul24_fa19_13_y4, h_s_arrmul24_fa20_13_y2, h_s_arrmul24_fa20_13_y4);
  and_gate and_gate_h_s_arrmul24_and21_13_y0(a_21, b_13, h_s_arrmul24_and21_13_y0);
  fa fa_h_s_arrmul24_fa21_13_y2(h_s_arrmul24_and21_13_y0, h_s_arrmul24_fa22_12_y2, h_s_arrmul24_fa20_13_y4, h_s_arrmul24_fa21_13_y2, h_s_arrmul24_fa21_13_y4);
  and_gate and_gate_h_s_arrmul24_and22_13_y0(a_22, b_13, h_s_arrmul24_and22_13_y0);
  fa fa_h_s_arrmul24_fa22_13_y2(h_s_arrmul24_and22_13_y0, h_s_arrmul24_fa23_12_y2, h_s_arrmul24_fa21_13_y4, h_s_arrmul24_fa22_13_y2, h_s_arrmul24_fa22_13_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_13_y0(a_23, b_13, h_s_arrmul24_nand23_13_y0);
  fa fa_h_s_arrmul24_fa23_13_y2(h_s_arrmul24_nand23_13_y0, h_s_arrmul24_fa23_12_y4, h_s_arrmul24_fa22_13_y4, h_s_arrmul24_fa23_13_y2, h_s_arrmul24_fa23_13_y4);
  and_gate and_gate_h_s_arrmul24_and0_14_y0(a_0, b_14, h_s_arrmul24_and0_14_y0);
  ha ha_h_s_arrmul24_ha0_14_y0(h_s_arrmul24_and0_14_y0, h_s_arrmul24_fa1_13_y2, h_s_arrmul24_ha0_14_y0, h_s_arrmul24_ha0_14_y1);
  and_gate and_gate_h_s_arrmul24_and1_14_y0(a_1, b_14, h_s_arrmul24_and1_14_y0);
  fa fa_h_s_arrmul24_fa1_14_y2(h_s_arrmul24_and1_14_y0, h_s_arrmul24_fa2_13_y2, h_s_arrmul24_ha0_14_y1, h_s_arrmul24_fa1_14_y2, h_s_arrmul24_fa1_14_y4);
  and_gate and_gate_h_s_arrmul24_and2_14_y0(a_2, b_14, h_s_arrmul24_and2_14_y0);
  fa fa_h_s_arrmul24_fa2_14_y2(h_s_arrmul24_and2_14_y0, h_s_arrmul24_fa3_13_y2, h_s_arrmul24_fa1_14_y4, h_s_arrmul24_fa2_14_y2, h_s_arrmul24_fa2_14_y4);
  and_gate and_gate_h_s_arrmul24_and3_14_y0(a_3, b_14, h_s_arrmul24_and3_14_y0);
  fa fa_h_s_arrmul24_fa3_14_y2(h_s_arrmul24_and3_14_y0, h_s_arrmul24_fa4_13_y2, h_s_arrmul24_fa2_14_y4, h_s_arrmul24_fa3_14_y2, h_s_arrmul24_fa3_14_y4);
  and_gate and_gate_h_s_arrmul24_and4_14_y0(a_4, b_14, h_s_arrmul24_and4_14_y0);
  fa fa_h_s_arrmul24_fa4_14_y2(h_s_arrmul24_and4_14_y0, h_s_arrmul24_fa5_13_y2, h_s_arrmul24_fa3_14_y4, h_s_arrmul24_fa4_14_y2, h_s_arrmul24_fa4_14_y4);
  and_gate and_gate_h_s_arrmul24_and5_14_y0(a_5, b_14, h_s_arrmul24_and5_14_y0);
  fa fa_h_s_arrmul24_fa5_14_y2(h_s_arrmul24_and5_14_y0, h_s_arrmul24_fa6_13_y2, h_s_arrmul24_fa4_14_y4, h_s_arrmul24_fa5_14_y2, h_s_arrmul24_fa5_14_y4);
  and_gate and_gate_h_s_arrmul24_and6_14_y0(a_6, b_14, h_s_arrmul24_and6_14_y0);
  fa fa_h_s_arrmul24_fa6_14_y2(h_s_arrmul24_and6_14_y0, h_s_arrmul24_fa7_13_y2, h_s_arrmul24_fa5_14_y4, h_s_arrmul24_fa6_14_y2, h_s_arrmul24_fa6_14_y4);
  and_gate and_gate_h_s_arrmul24_and7_14_y0(a_7, b_14, h_s_arrmul24_and7_14_y0);
  fa fa_h_s_arrmul24_fa7_14_y2(h_s_arrmul24_and7_14_y0, h_s_arrmul24_fa8_13_y2, h_s_arrmul24_fa6_14_y4, h_s_arrmul24_fa7_14_y2, h_s_arrmul24_fa7_14_y4);
  and_gate and_gate_h_s_arrmul24_and8_14_y0(a_8, b_14, h_s_arrmul24_and8_14_y0);
  fa fa_h_s_arrmul24_fa8_14_y2(h_s_arrmul24_and8_14_y0, h_s_arrmul24_fa9_13_y2, h_s_arrmul24_fa7_14_y4, h_s_arrmul24_fa8_14_y2, h_s_arrmul24_fa8_14_y4);
  and_gate and_gate_h_s_arrmul24_and9_14_y0(a_9, b_14, h_s_arrmul24_and9_14_y0);
  fa fa_h_s_arrmul24_fa9_14_y2(h_s_arrmul24_and9_14_y0, h_s_arrmul24_fa10_13_y2, h_s_arrmul24_fa8_14_y4, h_s_arrmul24_fa9_14_y2, h_s_arrmul24_fa9_14_y4);
  and_gate and_gate_h_s_arrmul24_and10_14_y0(a_10, b_14, h_s_arrmul24_and10_14_y0);
  fa fa_h_s_arrmul24_fa10_14_y2(h_s_arrmul24_and10_14_y0, h_s_arrmul24_fa11_13_y2, h_s_arrmul24_fa9_14_y4, h_s_arrmul24_fa10_14_y2, h_s_arrmul24_fa10_14_y4);
  and_gate and_gate_h_s_arrmul24_and11_14_y0(a_11, b_14, h_s_arrmul24_and11_14_y0);
  fa fa_h_s_arrmul24_fa11_14_y2(h_s_arrmul24_and11_14_y0, h_s_arrmul24_fa12_13_y2, h_s_arrmul24_fa10_14_y4, h_s_arrmul24_fa11_14_y2, h_s_arrmul24_fa11_14_y4);
  and_gate and_gate_h_s_arrmul24_and12_14_y0(a_12, b_14, h_s_arrmul24_and12_14_y0);
  fa fa_h_s_arrmul24_fa12_14_y2(h_s_arrmul24_and12_14_y0, h_s_arrmul24_fa13_13_y2, h_s_arrmul24_fa11_14_y4, h_s_arrmul24_fa12_14_y2, h_s_arrmul24_fa12_14_y4);
  and_gate and_gate_h_s_arrmul24_and13_14_y0(a_13, b_14, h_s_arrmul24_and13_14_y0);
  fa fa_h_s_arrmul24_fa13_14_y2(h_s_arrmul24_and13_14_y0, h_s_arrmul24_fa14_13_y2, h_s_arrmul24_fa12_14_y4, h_s_arrmul24_fa13_14_y2, h_s_arrmul24_fa13_14_y4);
  and_gate and_gate_h_s_arrmul24_and14_14_y0(a_14, b_14, h_s_arrmul24_and14_14_y0);
  fa fa_h_s_arrmul24_fa14_14_y2(h_s_arrmul24_and14_14_y0, h_s_arrmul24_fa15_13_y2, h_s_arrmul24_fa13_14_y4, h_s_arrmul24_fa14_14_y2, h_s_arrmul24_fa14_14_y4);
  and_gate and_gate_h_s_arrmul24_and15_14_y0(a_15, b_14, h_s_arrmul24_and15_14_y0);
  fa fa_h_s_arrmul24_fa15_14_y2(h_s_arrmul24_and15_14_y0, h_s_arrmul24_fa16_13_y2, h_s_arrmul24_fa14_14_y4, h_s_arrmul24_fa15_14_y2, h_s_arrmul24_fa15_14_y4);
  and_gate and_gate_h_s_arrmul24_and16_14_y0(a_16, b_14, h_s_arrmul24_and16_14_y0);
  fa fa_h_s_arrmul24_fa16_14_y2(h_s_arrmul24_and16_14_y0, h_s_arrmul24_fa17_13_y2, h_s_arrmul24_fa15_14_y4, h_s_arrmul24_fa16_14_y2, h_s_arrmul24_fa16_14_y4);
  and_gate and_gate_h_s_arrmul24_and17_14_y0(a_17, b_14, h_s_arrmul24_and17_14_y0);
  fa fa_h_s_arrmul24_fa17_14_y2(h_s_arrmul24_and17_14_y0, h_s_arrmul24_fa18_13_y2, h_s_arrmul24_fa16_14_y4, h_s_arrmul24_fa17_14_y2, h_s_arrmul24_fa17_14_y4);
  and_gate and_gate_h_s_arrmul24_and18_14_y0(a_18, b_14, h_s_arrmul24_and18_14_y0);
  fa fa_h_s_arrmul24_fa18_14_y2(h_s_arrmul24_and18_14_y0, h_s_arrmul24_fa19_13_y2, h_s_arrmul24_fa17_14_y4, h_s_arrmul24_fa18_14_y2, h_s_arrmul24_fa18_14_y4);
  and_gate and_gate_h_s_arrmul24_and19_14_y0(a_19, b_14, h_s_arrmul24_and19_14_y0);
  fa fa_h_s_arrmul24_fa19_14_y2(h_s_arrmul24_and19_14_y0, h_s_arrmul24_fa20_13_y2, h_s_arrmul24_fa18_14_y4, h_s_arrmul24_fa19_14_y2, h_s_arrmul24_fa19_14_y4);
  and_gate and_gate_h_s_arrmul24_and20_14_y0(a_20, b_14, h_s_arrmul24_and20_14_y0);
  fa fa_h_s_arrmul24_fa20_14_y2(h_s_arrmul24_and20_14_y0, h_s_arrmul24_fa21_13_y2, h_s_arrmul24_fa19_14_y4, h_s_arrmul24_fa20_14_y2, h_s_arrmul24_fa20_14_y4);
  and_gate and_gate_h_s_arrmul24_and21_14_y0(a_21, b_14, h_s_arrmul24_and21_14_y0);
  fa fa_h_s_arrmul24_fa21_14_y2(h_s_arrmul24_and21_14_y0, h_s_arrmul24_fa22_13_y2, h_s_arrmul24_fa20_14_y4, h_s_arrmul24_fa21_14_y2, h_s_arrmul24_fa21_14_y4);
  and_gate and_gate_h_s_arrmul24_and22_14_y0(a_22, b_14, h_s_arrmul24_and22_14_y0);
  fa fa_h_s_arrmul24_fa22_14_y2(h_s_arrmul24_and22_14_y0, h_s_arrmul24_fa23_13_y2, h_s_arrmul24_fa21_14_y4, h_s_arrmul24_fa22_14_y2, h_s_arrmul24_fa22_14_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_14_y0(a_23, b_14, h_s_arrmul24_nand23_14_y0);
  fa fa_h_s_arrmul24_fa23_14_y2(h_s_arrmul24_nand23_14_y0, h_s_arrmul24_fa23_13_y4, h_s_arrmul24_fa22_14_y4, h_s_arrmul24_fa23_14_y2, h_s_arrmul24_fa23_14_y4);
  and_gate and_gate_h_s_arrmul24_and0_15_y0(a_0, b_15, h_s_arrmul24_and0_15_y0);
  ha ha_h_s_arrmul24_ha0_15_y0(h_s_arrmul24_and0_15_y0, h_s_arrmul24_fa1_14_y2, h_s_arrmul24_ha0_15_y0, h_s_arrmul24_ha0_15_y1);
  and_gate and_gate_h_s_arrmul24_and1_15_y0(a_1, b_15, h_s_arrmul24_and1_15_y0);
  fa fa_h_s_arrmul24_fa1_15_y2(h_s_arrmul24_and1_15_y0, h_s_arrmul24_fa2_14_y2, h_s_arrmul24_ha0_15_y1, h_s_arrmul24_fa1_15_y2, h_s_arrmul24_fa1_15_y4);
  and_gate and_gate_h_s_arrmul24_and2_15_y0(a_2, b_15, h_s_arrmul24_and2_15_y0);
  fa fa_h_s_arrmul24_fa2_15_y2(h_s_arrmul24_and2_15_y0, h_s_arrmul24_fa3_14_y2, h_s_arrmul24_fa1_15_y4, h_s_arrmul24_fa2_15_y2, h_s_arrmul24_fa2_15_y4);
  and_gate and_gate_h_s_arrmul24_and3_15_y0(a_3, b_15, h_s_arrmul24_and3_15_y0);
  fa fa_h_s_arrmul24_fa3_15_y2(h_s_arrmul24_and3_15_y0, h_s_arrmul24_fa4_14_y2, h_s_arrmul24_fa2_15_y4, h_s_arrmul24_fa3_15_y2, h_s_arrmul24_fa3_15_y4);
  and_gate and_gate_h_s_arrmul24_and4_15_y0(a_4, b_15, h_s_arrmul24_and4_15_y0);
  fa fa_h_s_arrmul24_fa4_15_y2(h_s_arrmul24_and4_15_y0, h_s_arrmul24_fa5_14_y2, h_s_arrmul24_fa3_15_y4, h_s_arrmul24_fa4_15_y2, h_s_arrmul24_fa4_15_y4);
  and_gate and_gate_h_s_arrmul24_and5_15_y0(a_5, b_15, h_s_arrmul24_and5_15_y0);
  fa fa_h_s_arrmul24_fa5_15_y2(h_s_arrmul24_and5_15_y0, h_s_arrmul24_fa6_14_y2, h_s_arrmul24_fa4_15_y4, h_s_arrmul24_fa5_15_y2, h_s_arrmul24_fa5_15_y4);
  and_gate and_gate_h_s_arrmul24_and6_15_y0(a_6, b_15, h_s_arrmul24_and6_15_y0);
  fa fa_h_s_arrmul24_fa6_15_y2(h_s_arrmul24_and6_15_y0, h_s_arrmul24_fa7_14_y2, h_s_arrmul24_fa5_15_y4, h_s_arrmul24_fa6_15_y2, h_s_arrmul24_fa6_15_y4);
  and_gate and_gate_h_s_arrmul24_and7_15_y0(a_7, b_15, h_s_arrmul24_and7_15_y0);
  fa fa_h_s_arrmul24_fa7_15_y2(h_s_arrmul24_and7_15_y0, h_s_arrmul24_fa8_14_y2, h_s_arrmul24_fa6_15_y4, h_s_arrmul24_fa7_15_y2, h_s_arrmul24_fa7_15_y4);
  and_gate and_gate_h_s_arrmul24_and8_15_y0(a_8, b_15, h_s_arrmul24_and8_15_y0);
  fa fa_h_s_arrmul24_fa8_15_y2(h_s_arrmul24_and8_15_y0, h_s_arrmul24_fa9_14_y2, h_s_arrmul24_fa7_15_y4, h_s_arrmul24_fa8_15_y2, h_s_arrmul24_fa8_15_y4);
  and_gate and_gate_h_s_arrmul24_and9_15_y0(a_9, b_15, h_s_arrmul24_and9_15_y0);
  fa fa_h_s_arrmul24_fa9_15_y2(h_s_arrmul24_and9_15_y0, h_s_arrmul24_fa10_14_y2, h_s_arrmul24_fa8_15_y4, h_s_arrmul24_fa9_15_y2, h_s_arrmul24_fa9_15_y4);
  and_gate and_gate_h_s_arrmul24_and10_15_y0(a_10, b_15, h_s_arrmul24_and10_15_y0);
  fa fa_h_s_arrmul24_fa10_15_y2(h_s_arrmul24_and10_15_y0, h_s_arrmul24_fa11_14_y2, h_s_arrmul24_fa9_15_y4, h_s_arrmul24_fa10_15_y2, h_s_arrmul24_fa10_15_y4);
  and_gate and_gate_h_s_arrmul24_and11_15_y0(a_11, b_15, h_s_arrmul24_and11_15_y0);
  fa fa_h_s_arrmul24_fa11_15_y2(h_s_arrmul24_and11_15_y0, h_s_arrmul24_fa12_14_y2, h_s_arrmul24_fa10_15_y4, h_s_arrmul24_fa11_15_y2, h_s_arrmul24_fa11_15_y4);
  and_gate and_gate_h_s_arrmul24_and12_15_y0(a_12, b_15, h_s_arrmul24_and12_15_y0);
  fa fa_h_s_arrmul24_fa12_15_y2(h_s_arrmul24_and12_15_y0, h_s_arrmul24_fa13_14_y2, h_s_arrmul24_fa11_15_y4, h_s_arrmul24_fa12_15_y2, h_s_arrmul24_fa12_15_y4);
  and_gate and_gate_h_s_arrmul24_and13_15_y0(a_13, b_15, h_s_arrmul24_and13_15_y0);
  fa fa_h_s_arrmul24_fa13_15_y2(h_s_arrmul24_and13_15_y0, h_s_arrmul24_fa14_14_y2, h_s_arrmul24_fa12_15_y4, h_s_arrmul24_fa13_15_y2, h_s_arrmul24_fa13_15_y4);
  and_gate and_gate_h_s_arrmul24_and14_15_y0(a_14, b_15, h_s_arrmul24_and14_15_y0);
  fa fa_h_s_arrmul24_fa14_15_y2(h_s_arrmul24_and14_15_y0, h_s_arrmul24_fa15_14_y2, h_s_arrmul24_fa13_15_y4, h_s_arrmul24_fa14_15_y2, h_s_arrmul24_fa14_15_y4);
  and_gate and_gate_h_s_arrmul24_and15_15_y0(a_15, b_15, h_s_arrmul24_and15_15_y0);
  fa fa_h_s_arrmul24_fa15_15_y2(h_s_arrmul24_and15_15_y0, h_s_arrmul24_fa16_14_y2, h_s_arrmul24_fa14_15_y4, h_s_arrmul24_fa15_15_y2, h_s_arrmul24_fa15_15_y4);
  and_gate and_gate_h_s_arrmul24_and16_15_y0(a_16, b_15, h_s_arrmul24_and16_15_y0);
  fa fa_h_s_arrmul24_fa16_15_y2(h_s_arrmul24_and16_15_y0, h_s_arrmul24_fa17_14_y2, h_s_arrmul24_fa15_15_y4, h_s_arrmul24_fa16_15_y2, h_s_arrmul24_fa16_15_y4);
  and_gate and_gate_h_s_arrmul24_and17_15_y0(a_17, b_15, h_s_arrmul24_and17_15_y0);
  fa fa_h_s_arrmul24_fa17_15_y2(h_s_arrmul24_and17_15_y0, h_s_arrmul24_fa18_14_y2, h_s_arrmul24_fa16_15_y4, h_s_arrmul24_fa17_15_y2, h_s_arrmul24_fa17_15_y4);
  and_gate and_gate_h_s_arrmul24_and18_15_y0(a_18, b_15, h_s_arrmul24_and18_15_y0);
  fa fa_h_s_arrmul24_fa18_15_y2(h_s_arrmul24_and18_15_y0, h_s_arrmul24_fa19_14_y2, h_s_arrmul24_fa17_15_y4, h_s_arrmul24_fa18_15_y2, h_s_arrmul24_fa18_15_y4);
  and_gate and_gate_h_s_arrmul24_and19_15_y0(a_19, b_15, h_s_arrmul24_and19_15_y0);
  fa fa_h_s_arrmul24_fa19_15_y2(h_s_arrmul24_and19_15_y0, h_s_arrmul24_fa20_14_y2, h_s_arrmul24_fa18_15_y4, h_s_arrmul24_fa19_15_y2, h_s_arrmul24_fa19_15_y4);
  and_gate and_gate_h_s_arrmul24_and20_15_y0(a_20, b_15, h_s_arrmul24_and20_15_y0);
  fa fa_h_s_arrmul24_fa20_15_y2(h_s_arrmul24_and20_15_y0, h_s_arrmul24_fa21_14_y2, h_s_arrmul24_fa19_15_y4, h_s_arrmul24_fa20_15_y2, h_s_arrmul24_fa20_15_y4);
  and_gate and_gate_h_s_arrmul24_and21_15_y0(a_21, b_15, h_s_arrmul24_and21_15_y0);
  fa fa_h_s_arrmul24_fa21_15_y2(h_s_arrmul24_and21_15_y0, h_s_arrmul24_fa22_14_y2, h_s_arrmul24_fa20_15_y4, h_s_arrmul24_fa21_15_y2, h_s_arrmul24_fa21_15_y4);
  and_gate and_gate_h_s_arrmul24_and22_15_y0(a_22, b_15, h_s_arrmul24_and22_15_y0);
  fa fa_h_s_arrmul24_fa22_15_y2(h_s_arrmul24_and22_15_y0, h_s_arrmul24_fa23_14_y2, h_s_arrmul24_fa21_15_y4, h_s_arrmul24_fa22_15_y2, h_s_arrmul24_fa22_15_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_15_y0(a_23, b_15, h_s_arrmul24_nand23_15_y0);
  fa fa_h_s_arrmul24_fa23_15_y2(h_s_arrmul24_nand23_15_y0, h_s_arrmul24_fa23_14_y4, h_s_arrmul24_fa22_15_y4, h_s_arrmul24_fa23_15_y2, h_s_arrmul24_fa23_15_y4);
  and_gate and_gate_h_s_arrmul24_and0_16_y0(a_0, b_16, h_s_arrmul24_and0_16_y0);
  ha ha_h_s_arrmul24_ha0_16_y0(h_s_arrmul24_and0_16_y0, h_s_arrmul24_fa1_15_y2, h_s_arrmul24_ha0_16_y0, h_s_arrmul24_ha0_16_y1);
  and_gate and_gate_h_s_arrmul24_and1_16_y0(a_1, b_16, h_s_arrmul24_and1_16_y0);
  fa fa_h_s_arrmul24_fa1_16_y2(h_s_arrmul24_and1_16_y0, h_s_arrmul24_fa2_15_y2, h_s_arrmul24_ha0_16_y1, h_s_arrmul24_fa1_16_y2, h_s_arrmul24_fa1_16_y4);
  and_gate and_gate_h_s_arrmul24_and2_16_y0(a_2, b_16, h_s_arrmul24_and2_16_y0);
  fa fa_h_s_arrmul24_fa2_16_y2(h_s_arrmul24_and2_16_y0, h_s_arrmul24_fa3_15_y2, h_s_arrmul24_fa1_16_y4, h_s_arrmul24_fa2_16_y2, h_s_arrmul24_fa2_16_y4);
  and_gate and_gate_h_s_arrmul24_and3_16_y0(a_3, b_16, h_s_arrmul24_and3_16_y0);
  fa fa_h_s_arrmul24_fa3_16_y2(h_s_arrmul24_and3_16_y0, h_s_arrmul24_fa4_15_y2, h_s_arrmul24_fa2_16_y4, h_s_arrmul24_fa3_16_y2, h_s_arrmul24_fa3_16_y4);
  and_gate and_gate_h_s_arrmul24_and4_16_y0(a_4, b_16, h_s_arrmul24_and4_16_y0);
  fa fa_h_s_arrmul24_fa4_16_y2(h_s_arrmul24_and4_16_y0, h_s_arrmul24_fa5_15_y2, h_s_arrmul24_fa3_16_y4, h_s_arrmul24_fa4_16_y2, h_s_arrmul24_fa4_16_y4);
  and_gate and_gate_h_s_arrmul24_and5_16_y0(a_5, b_16, h_s_arrmul24_and5_16_y0);
  fa fa_h_s_arrmul24_fa5_16_y2(h_s_arrmul24_and5_16_y0, h_s_arrmul24_fa6_15_y2, h_s_arrmul24_fa4_16_y4, h_s_arrmul24_fa5_16_y2, h_s_arrmul24_fa5_16_y4);
  and_gate and_gate_h_s_arrmul24_and6_16_y0(a_6, b_16, h_s_arrmul24_and6_16_y0);
  fa fa_h_s_arrmul24_fa6_16_y2(h_s_arrmul24_and6_16_y0, h_s_arrmul24_fa7_15_y2, h_s_arrmul24_fa5_16_y4, h_s_arrmul24_fa6_16_y2, h_s_arrmul24_fa6_16_y4);
  and_gate and_gate_h_s_arrmul24_and7_16_y0(a_7, b_16, h_s_arrmul24_and7_16_y0);
  fa fa_h_s_arrmul24_fa7_16_y2(h_s_arrmul24_and7_16_y0, h_s_arrmul24_fa8_15_y2, h_s_arrmul24_fa6_16_y4, h_s_arrmul24_fa7_16_y2, h_s_arrmul24_fa7_16_y4);
  and_gate and_gate_h_s_arrmul24_and8_16_y0(a_8, b_16, h_s_arrmul24_and8_16_y0);
  fa fa_h_s_arrmul24_fa8_16_y2(h_s_arrmul24_and8_16_y0, h_s_arrmul24_fa9_15_y2, h_s_arrmul24_fa7_16_y4, h_s_arrmul24_fa8_16_y2, h_s_arrmul24_fa8_16_y4);
  and_gate and_gate_h_s_arrmul24_and9_16_y0(a_9, b_16, h_s_arrmul24_and9_16_y0);
  fa fa_h_s_arrmul24_fa9_16_y2(h_s_arrmul24_and9_16_y0, h_s_arrmul24_fa10_15_y2, h_s_arrmul24_fa8_16_y4, h_s_arrmul24_fa9_16_y2, h_s_arrmul24_fa9_16_y4);
  and_gate and_gate_h_s_arrmul24_and10_16_y0(a_10, b_16, h_s_arrmul24_and10_16_y0);
  fa fa_h_s_arrmul24_fa10_16_y2(h_s_arrmul24_and10_16_y0, h_s_arrmul24_fa11_15_y2, h_s_arrmul24_fa9_16_y4, h_s_arrmul24_fa10_16_y2, h_s_arrmul24_fa10_16_y4);
  and_gate and_gate_h_s_arrmul24_and11_16_y0(a_11, b_16, h_s_arrmul24_and11_16_y0);
  fa fa_h_s_arrmul24_fa11_16_y2(h_s_arrmul24_and11_16_y0, h_s_arrmul24_fa12_15_y2, h_s_arrmul24_fa10_16_y4, h_s_arrmul24_fa11_16_y2, h_s_arrmul24_fa11_16_y4);
  and_gate and_gate_h_s_arrmul24_and12_16_y0(a_12, b_16, h_s_arrmul24_and12_16_y0);
  fa fa_h_s_arrmul24_fa12_16_y2(h_s_arrmul24_and12_16_y0, h_s_arrmul24_fa13_15_y2, h_s_arrmul24_fa11_16_y4, h_s_arrmul24_fa12_16_y2, h_s_arrmul24_fa12_16_y4);
  and_gate and_gate_h_s_arrmul24_and13_16_y0(a_13, b_16, h_s_arrmul24_and13_16_y0);
  fa fa_h_s_arrmul24_fa13_16_y2(h_s_arrmul24_and13_16_y0, h_s_arrmul24_fa14_15_y2, h_s_arrmul24_fa12_16_y4, h_s_arrmul24_fa13_16_y2, h_s_arrmul24_fa13_16_y4);
  and_gate and_gate_h_s_arrmul24_and14_16_y0(a_14, b_16, h_s_arrmul24_and14_16_y0);
  fa fa_h_s_arrmul24_fa14_16_y2(h_s_arrmul24_and14_16_y0, h_s_arrmul24_fa15_15_y2, h_s_arrmul24_fa13_16_y4, h_s_arrmul24_fa14_16_y2, h_s_arrmul24_fa14_16_y4);
  and_gate and_gate_h_s_arrmul24_and15_16_y0(a_15, b_16, h_s_arrmul24_and15_16_y0);
  fa fa_h_s_arrmul24_fa15_16_y2(h_s_arrmul24_and15_16_y0, h_s_arrmul24_fa16_15_y2, h_s_arrmul24_fa14_16_y4, h_s_arrmul24_fa15_16_y2, h_s_arrmul24_fa15_16_y4);
  and_gate and_gate_h_s_arrmul24_and16_16_y0(a_16, b_16, h_s_arrmul24_and16_16_y0);
  fa fa_h_s_arrmul24_fa16_16_y2(h_s_arrmul24_and16_16_y0, h_s_arrmul24_fa17_15_y2, h_s_arrmul24_fa15_16_y4, h_s_arrmul24_fa16_16_y2, h_s_arrmul24_fa16_16_y4);
  and_gate and_gate_h_s_arrmul24_and17_16_y0(a_17, b_16, h_s_arrmul24_and17_16_y0);
  fa fa_h_s_arrmul24_fa17_16_y2(h_s_arrmul24_and17_16_y0, h_s_arrmul24_fa18_15_y2, h_s_arrmul24_fa16_16_y4, h_s_arrmul24_fa17_16_y2, h_s_arrmul24_fa17_16_y4);
  and_gate and_gate_h_s_arrmul24_and18_16_y0(a_18, b_16, h_s_arrmul24_and18_16_y0);
  fa fa_h_s_arrmul24_fa18_16_y2(h_s_arrmul24_and18_16_y0, h_s_arrmul24_fa19_15_y2, h_s_arrmul24_fa17_16_y4, h_s_arrmul24_fa18_16_y2, h_s_arrmul24_fa18_16_y4);
  and_gate and_gate_h_s_arrmul24_and19_16_y0(a_19, b_16, h_s_arrmul24_and19_16_y0);
  fa fa_h_s_arrmul24_fa19_16_y2(h_s_arrmul24_and19_16_y0, h_s_arrmul24_fa20_15_y2, h_s_arrmul24_fa18_16_y4, h_s_arrmul24_fa19_16_y2, h_s_arrmul24_fa19_16_y4);
  and_gate and_gate_h_s_arrmul24_and20_16_y0(a_20, b_16, h_s_arrmul24_and20_16_y0);
  fa fa_h_s_arrmul24_fa20_16_y2(h_s_arrmul24_and20_16_y0, h_s_arrmul24_fa21_15_y2, h_s_arrmul24_fa19_16_y4, h_s_arrmul24_fa20_16_y2, h_s_arrmul24_fa20_16_y4);
  and_gate and_gate_h_s_arrmul24_and21_16_y0(a_21, b_16, h_s_arrmul24_and21_16_y0);
  fa fa_h_s_arrmul24_fa21_16_y2(h_s_arrmul24_and21_16_y0, h_s_arrmul24_fa22_15_y2, h_s_arrmul24_fa20_16_y4, h_s_arrmul24_fa21_16_y2, h_s_arrmul24_fa21_16_y4);
  and_gate and_gate_h_s_arrmul24_and22_16_y0(a_22, b_16, h_s_arrmul24_and22_16_y0);
  fa fa_h_s_arrmul24_fa22_16_y2(h_s_arrmul24_and22_16_y0, h_s_arrmul24_fa23_15_y2, h_s_arrmul24_fa21_16_y4, h_s_arrmul24_fa22_16_y2, h_s_arrmul24_fa22_16_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_16_y0(a_23, b_16, h_s_arrmul24_nand23_16_y0);
  fa fa_h_s_arrmul24_fa23_16_y2(h_s_arrmul24_nand23_16_y0, h_s_arrmul24_fa23_15_y4, h_s_arrmul24_fa22_16_y4, h_s_arrmul24_fa23_16_y2, h_s_arrmul24_fa23_16_y4);
  and_gate and_gate_h_s_arrmul24_and0_17_y0(a_0, b_17, h_s_arrmul24_and0_17_y0);
  ha ha_h_s_arrmul24_ha0_17_y0(h_s_arrmul24_and0_17_y0, h_s_arrmul24_fa1_16_y2, h_s_arrmul24_ha0_17_y0, h_s_arrmul24_ha0_17_y1);
  and_gate and_gate_h_s_arrmul24_and1_17_y0(a_1, b_17, h_s_arrmul24_and1_17_y0);
  fa fa_h_s_arrmul24_fa1_17_y2(h_s_arrmul24_and1_17_y0, h_s_arrmul24_fa2_16_y2, h_s_arrmul24_ha0_17_y1, h_s_arrmul24_fa1_17_y2, h_s_arrmul24_fa1_17_y4);
  and_gate and_gate_h_s_arrmul24_and2_17_y0(a_2, b_17, h_s_arrmul24_and2_17_y0);
  fa fa_h_s_arrmul24_fa2_17_y2(h_s_arrmul24_and2_17_y0, h_s_arrmul24_fa3_16_y2, h_s_arrmul24_fa1_17_y4, h_s_arrmul24_fa2_17_y2, h_s_arrmul24_fa2_17_y4);
  and_gate and_gate_h_s_arrmul24_and3_17_y0(a_3, b_17, h_s_arrmul24_and3_17_y0);
  fa fa_h_s_arrmul24_fa3_17_y2(h_s_arrmul24_and3_17_y0, h_s_arrmul24_fa4_16_y2, h_s_arrmul24_fa2_17_y4, h_s_arrmul24_fa3_17_y2, h_s_arrmul24_fa3_17_y4);
  and_gate and_gate_h_s_arrmul24_and4_17_y0(a_4, b_17, h_s_arrmul24_and4_17_y0);
  fa fa_h_s_arrmul24_fa4_17_y2(h_s_arrmul24_and4_17_y0, h_s_arrmul24_fa5_16_y2, h_s_arrmul24_fa3_17_y4, h_s_arrmul24_fa4_17_y2, h_s_arrmul24_fa4_17_y4);
  and_gate and_gate_h_s_arrmul24_and5_17_y0(a_5, b_17, h_s_arrmul24_and5_17_y0);
  fa fa_h_s_arrmul24_fa5_17_y2(h_s_arrmul24_and5_17_y0, h_s_arrmul24_fa6_16_y2, h_s_arrmul24_fa4_17_y4, h_s_arrmul24_fa5_17_y2, h_s_arrmul24_fa5_17_y4);
  and_gate and_gate_h_s_arrmul24_and6_17_y0(a_6, b_17, h_s_arrmul24_and6_17_y0);
  fa fa_h_s_arrmul24_fa6_17_y2(h_s_arrmul24_and6_17_y0, h_s_arrmul24_fa7_16_y2, h_s_arrmul24_fa5_17_y4, h_s_arrmul24_fa6_17_y2, h_s_arrmul24_fa6_17_y4);
  and_gate and_gate_h_s_arrmul24_and7_17_y0(a_7, b_17, h_s_arrmul24_and7_17_y0);
  fa fa_h_s_arrmul24_fa7_17_y2(h_s_arrmul24_and7_17_y0, h_s_arrmul24_fa8_16_y2, h_s_arrmul24_fa6_17_y4, h_s_arrmul24_fa7_17_y2, h_s_arrmul24_fa7_17_y4);
  and_gate and_gate_h_s_arrmul24_and8_17_y0(a_8, b_17, h_s_arrmul24_and8_17_y0);
  fa fa_h_s_arrmul24_fa8_17_y2(h_s_arrmul24_and8_17_y0, h_s_arrmul24_fa9_16_y2, h_s_arrmul24_fa7_17_y4, h_s_arrmul24_fa8_17_y2, h_s_arrmul24_fa8_17_y4);
  and_gate and_gate_h_s_arrmul24_and9_17_y0(a_9, b_17, h_s_arrmul24_and9_17_y0);
  fa fa_h_s_arrmul24_fa9_17_y2(h_s_arrmul24_and9_17_y0, h_s_arrmul24_fa10_16_y2, h_s_arrmul24_fa8_17_y4, h_s_arrmul24_fa9_17_y2, h_s_arrmul24_fa9_17_y4);
  and_gate and_gate_h_s_arrmul24_and10_17_y0(a_10, b_17, h_s_arrmul24_and10_17_y0);
  fa fa_h_s_arrmul24_fa10_17_y2(h_s_arrmul24_and10_17_y0, h_s_arrmul24_fa11_16_y2, h_s_arrmul24_fa9_17_y4, h_s_arrmul24_fa10_17_y2, h_s_arrmul24_fa10_17_y4);
  and_gate and_gate_h_s_arrmul24_and11_17_y0(a_11, b_17, h_s_arrmul24_and11_17_y0);
  fa fa_h_s_arrmul24_fa11_17_y2(h_s_arrmul24_and11_17_y0, h_s_arrmul24_fa12_16_y2, h_s_arrmul24_fa10_17_y4, h_s_arrmul24_fa11_17_y2, h_s_arrmul24_fa11_17_y4);
  and_gate and_gate_h_s_arrmul24_and12_17_y0(a_12, b_17, h_s_arrmul24_and12_17_y0);
  fa fa_h_s_arrmul24_fa12_17_y2(h_s_arrmul24_and12_17_y0, h_s_arrmul24_fa13_16_y2, h_s_arrmul24_fa11_17_y4, h_s_arrmul24_fa12_17_y2, h_s_arrmul24_fa12_17_y4);
  and_gate and_gate_h_s_arrmul24_and13_17_y0(a_13, b_17, h_s_arrmul24_and13_17_y0);
  fa fa_h_s_arrmul24_fa13_17_y2(h_s_arrmul24_and13_17_y0, h_s_arrmul24_fa14_16_y2, h_s_arrmul24_fa12_17_y4, h_s_arrmul24_fa13_17_y2, h_s_arrmul24_fa13_17_y4);
  and_gate and_gate_h_s_arrmul24_and14_17_y0(a_14, b_17, h_s_arrmul24_and14_17_y0);
  fa fa_h_s_arrmul24_fa14_17_y2(h_s_arrmul24_and14_17_y0, h_s_arrmul24_fa15_16_y2, h_s_arrmul24_fa13_17_y4, h_s_arrmul24_fa14_17_y2, h_s_arrmul24_fa14_17_y4);
  and_gate and_gate_h_s_arrmul24_and15_17_y0(a_15, b_17, h_s_arrmul24_and15_17_y0);
  fa fa_h_s_arrmul24_fa15_17_y2(h_s_arrmul24_and15_17_y0, h_s_arrmul24_fa16_16_y2, h_s_arrmul24_fa14_17_y4, h_s_arrmul24_fa15_17_y2, h_s_arrmul24_fa15_17_y4);
  and_gate and_gate_h_s_arrmul24_and16_17_y0(a_16, b_17, h_s_arrmul24_and16_17_y0);
  fa fa_h_s_arrmul24_fa16_17_y2(h_s_arrmul24_and16_17_y0, h_s_arrmul24_fa17_16_y2, h_s_arrmul24_fa15_17_y4, h_s_arrmul24_fa16_17_y2, h_s_arrmul24_fa16_17_y4);
  and_gate and_gate_h_s_arrmul24_and17_17_y0(a_17, b_17, h_s_arrmul24_and17_17_y0);
  fa fa_h_s_arrmul24_fa17_17_y2(h_s_arrmul24_and17_17_y0, h_s_arrmul24_fa18_16_y2, h_s_arrmul24_fa16_17_y4, h_s_arrmul24_fa17_17_y2, h_s_arrmul24_fa17_17_y4);
  and_gate and_gate_h_s_arrmul24_and18_17_y0(a_18, b_17, h_s_arrmul24_and18_17_y0);
  fa fa_h_s_arrmul24_fa18_17_y2(h_s_arrmul24_and18_17_y0, h_s_arrmul24_fa19_16_y2, h_s_arrmul24_fa17_17_y4, h_s_arrmul24_fa18_17_y2, h_s_arrmul24_fa18_17_y4);
  and_gate and_gate_h_s_arrmul24_and19_17_y0(a_19, b_17, h_s_arrmul24_and19_17_y0);
  fa fa_h_s_arrmul24_fa19_17_y2(h_s_arrmul24_and19_17_y0, h_s_arrmul24_fa20_16_y2, h_s_arrmul24_fa18_17_y4, h_s_arrmul24_fa19_17_y2, h_s_arrmul24_fa19_17_y4);
  and_gate and_gate_h_s_arrmul24_and20_17_y0(a_20, b_17, h_s_arrmul24_and20_17_y0);
  fa fa_h_s_arrmul24_fa20_17_y2(h_s_arrmul24_and20_17_y0, h_s_arrmul24_fa21_16_y2, h_s_arrmul24_fa19_17_y4, h_s_arrmul24_fa20_17_y2, h_s_arrmul24_fa20_17_y4);
  and_gate and_gate_h_s_arrmul24_and21_17_y0(a_21, b_17, h_s_arrmul24_and21_17_y0);
  fa fa_h_s_arrmul24_fa21_17_y2(h_s_arrmul24_and21_17_y0, h_s_arrmul24_fa22_16_y2, h_s_arrmul24_fa20_17_y4, h_s_arrmul24_fa21_17_y2, h_s_arrmul24_fa21_17_y4);
  and_gate and_gate_h_s_arrmul24_and22_17_y0(a_22, b_17, h_s_arrmul24_and22_17_y0);
  fa fa_h_s_arrmul24_fa22_17_y2(h_s_arrmul24_and22_17_y0, h_s_arrmul24_fa23_16_y2, h_s_arrmul24_fa21_17_y4, h_s_arrmul24_fa22_17_y2, h_s_arrmul24_fa22_17_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_17_y0(a_23, b_17, h_s_arrmul24_nand23_17_y0);
  fa fa_h_s_arrmul24_fa23_17_y2(h_s_arrmul24_nand23_17_y0, h_s_arrmul24_fa23_16_y4, h_s_arrmul24_fa22_17_y4, h_s_arrmul24_fa23_17_y2, h_s_arrmul24_fa23_17_y4);
  and_gate and_gate_h_s_arrmul24_and0_18_y0(a_0, b_18, h_s_arrmul24_and0_18_y0);
  ha ha_h_s_arrmul24_ha0_18_y0(h_s_arrmul24_and0_18_y0, h_s_arrmul24_fa1_17_y2, h_s_arrmul24_ha0_18_y0, h_s_arrmul24_ha0_18_y1);
  and_gate and_gate_h_s_arrmul24_and1_18_y0(a_1, b_18, h_s_arrmul24_and1_18_y0);
  fa fa_h_s_arrmul24_fa1_18_y2(h_s_arrmul24_and1_18_y0, h_s_arrmul24_fa2_17_y2, h_s_arrmul24_ha0_18_y1, h_s_arrmul24_fa1_18_y2, h_s_arrmul24_fa1_18_y4);
  and_gate and_gate_h_s_arrmul24_and2_18_y0(a_2, b_18, h_s_arrmul24_and2_18_y0);
  fa fa_h_s_arrmul24_fa2_18_y2(h_s_arrmul24_and2_18_y0, h_s_arrmul24_fa3_17_y2, h_s_arrmul24_fa1_18_y4, h_s_arrmul24_fa2_18_y2, h_s_arrmul24_fa2_18_y4);
  and_gate and_gate_h_s_arrmul24_and3_18_y0(a_3, b_18, h_s_arrmul24_and3_18_y0);
  fa fa_h_s_arrmul24_fa3_18_y2(h_s_arrmul24_and3_18_y0, h_s_arrmul24_fa4_17_y2, h_s_arrmul24_fa2_18_y4, h_s_arrmul24_fa3_18_y2, h_s_arrmul24_fa3_18_y4);
  and_gate and_gate_h_s_arrmul24_and4_18_y0(a_4, b_18, h_s_arrmul24_and4_18_y0);
  fa fa_h_s_arrmul24_fa4_18_y2(h_s_arrmul24_and4_18_y0, h_s_arrmul24_fa5_17_y2, h_s_arrmul24_fa3_18_y4, h_s_arrmul24_fa4_18_y2, h_s_arrmul24_fa4_18_y4);
  and_gate and_gate_h_s_arrmul24_and5_18_y0(a_5, b_18, h_s_arrmul24_and5_18_y0);
  fa fa_h_s_arrmul24_fa5_18_y2(h_s_arrmul24_and5_18_y0, h_s_arrmul24_fa6_17_y2, h_s_arrmul24_fa4_18_y4, h_s_arrmul24_fa5_18_y2, h_s_arrmul24_fa5_18_y4);
  and_gate and_gate_h_s_arrmul24_and6_18_y0(a_6, b_18, h_s_arrmul24_and6_18_y0);
  fa fa_h_s_arrmul24_fa6_18_y2(h_s_arrmul24_and6_18_y0, h_s_arrmul24_fa7_17_y2, h_s_arrmul24_fa5_18_y4, h_s_arrmul24_fa6_18_y2, h_s_arrmul24_fa6_18_y4);
  and_gate and_gate_h_s_arrmul24_and7_18_y0(a_7, b_18, h_s_arrmul24_and7_18_y0);
  fa fa_h_s_arrmul24_fa7_18_y2(h_s_arrmul24_and7_18_y0, h_s_arrmul24_fa8_17_y2, h_s_arrmul24_fa6_18_y4, h_s_arrmul24_fa7_18_y2, h_s_arrmul24_fa7_18_y4);
  and_gate and_gate_h_s_arrmul24_and8_18_y0(a_8, b_18, h_s_arrmul24_and8_18_y0);
  fa fa_h_s_arrmul24_fa8_18_y2(h_s_arrmul24_and8_18_y0, h_s_arrmul24_fa9_17_y2, h_s_arrmul24_fa7_18_y4, h_s_arrmul24_fa8_18_y2, h_s_arrmul24_fa8_18_y4);
  and_gate and_gate_h_s_arrmul24_and9_18_y0(a_9, b_18, h_s_arrmul24_and9_18_y0);
  fa fa_h_s_arrmul24_fa9_18_y2(h_s_arrmul24_and9_18_y0, h_s_arrmul24_fa10_17_y2, h_s_arrmul24_fa8_18_y4, h_s_arrmul24_fa9_18_y2, h_s_arrmul24_fa9_18_y4);
  and_gate and_gate_h_s_arrmul24_and10_18_y0(a_10, b_18, h_s_arrmul24_and10_18_y0);
  fa fa_h_s_arrmul24_fa10_18_y2(h_s_arrmul24_and10_18_y0, h_s_arrmul24_fa11_17_y2, h_s_arrmul24_fa9_18_y4, h_s_arrmul24_fa10_18_y2, h_s_arrmul24_fa10_18_y4);
  and_gate and_gate_h_s_arrmul24_and11_18_y0(a_11, b_18, h_s_arrmul24_and11_18_y0);
  fa fa_h_s_arrmul24_fa11_18_y2(h_s_arrmul24_and11_18_y0, h_s_arrmul24_fa12_17_y2, h_s_arrmul24_fa10_18_y4, h_s_arrmul24_fa11_18_y2, h_s_arrmul24_fa11_18_y4);
  and_gate and_gate_h_s_arrmul24_and12_18_y0(a_12, b_18, h_s_arrmul24_and12_18_y0);
  fa fa_h_s_arrmul24_fa12_18_y2(h_s_arrmul24_and12_18_y0, h_s_arrmul24_fa13_17_y2, h_s_arrmul24_fa11_18_y4, h_s_arrmul24_fa12_18_y2, h_s_arrmul24_fa12_18_y4);
  and_gate and_gate_h_s_arrmul24_and13_18_y0(a_13, b_18, h_s_arrmul24_and13_18_y0);
  fa fa_h_s_arrmul24_fa13_18_y2(h_s_arrmul24_and13_18_y0, h_s_arrmul24_fa14_17_y2, h_s_arrmul24_fa12_18_y4, h_s_arrmul24_fa13_18_y2, h_s_arrmul24_fa13_18_y4);
  and_gate and_gate_h_s_arrmul24_and14_18_y0(a_14, b_18, h_s_arrmul24_and14_18_y0);
  fa fa_h_s_arrmul24_fa14_18_y2(h_s_arrmul24_and14_18_y0, h_s_arrmul24_fa15_17_y2, h_s_arrmul24_fa13_18_y4, h_s_arrmul24_fa14_18_y2, h_s_arrmul24_fa14_18_y4);
  and_gate and_gate_h_s_arrmul24_and15_18_y0(a_15, b_18, h_s_arrmul24_and15_18_y0);
  fa fa_h_s_arrmul24_fa15_18_y2(h_s_arrmul24_and15_18_y0, h_s_arrmul24_fa16_17_y2, h_s_arrmul24_fa14_18_y4, h_s_arrmul24_fa15_18_y2, h_s_arrmul24_fa15_18_y4);
  and_gate and_gate_h_s_arrmul24_and16_18_y0(a_16, b_18, h_s_arrmul24_and16_18_y0);
  fa fa_h_s_arrmul24_fa16_18_y2(h_s_arrmul24_and16_18_y0, h_s_arrmul24_fa17_17_y2, h_s_arrmul24_fa15_18_y4, h_s_arrmul24_fa16_18_y2, h_s_arrmul24_fa16_18_y4);
  and_gate and_gate_h_s_arrmul24_and17_18_y0(a_17, b_18, h_s_arrmul24_and17_18_y0);
  fa fa_h_s_arrmul24_fa17_18_y2(h_s_arrmul24_and17_18_y0, h_s_arrmul24_fa18_17_y2, h_s_arrmul24_fa16_18_y4, h_s_arrmul24_fa17_18_y2, h_s_arrmul24_fa17_18_y4);
  and_gate and_gate_h_s_arrmul24_and18_18_y0(a_18, b_18, h_s_arrmul24_and18_18_y0);
  fa fa_h_s_arrmul24_fa18_18_y2(h_s_arrmul24_and18_18_y0, h_s_arrmul24_fa19_17_y2, h_s_arrmul24_fa17_18_y4, h_s_arrmul24_fa18_18_y2, h_s_arrmul24_fa18_18_y4);
  and_gate and_gate_h_s_arrmul24_and19_18_y0(a_19, b_18, h_s_arrmul24_and19_18_y0);
  fa fa_h_s_arrmul24_fa19_18_y2(h_s_arrmul24_and19_18_y0, h_s_arrmul24_fa20_17_y2, h_s_arrmul24_fa18_18_y4, h_s_arrmul24_fa19_18_y2, h_s_arrmul24_fa19_18_y4);
  and_gate and_gate_h_s_arrmul24_and20_18_y0(a_20, b_18, h_s_arrmul24_and20_18_y0);
  fa fa_h_s_arrmul24_fa20_18_y2(h_s_arrmul24_and20_18_y0, h_s_arrmul24_fa21_17_y2, h_s_arrmul24_fa19_18_y4, h_s_arrmul24_fa20_18_y2, h_s_arrmul24_fa20_18_y4);
  and_gate and_gate_h_s_arrmul24_and21_18_y0(a_21, b_18, h_s_arrmul24_and21_18_y0);
  fa fa_h_s_arrmul24_fa21_18_y2(h_s_arrmul24_and21_18_y0, h_s_arrmul24_fa22_17_y2, h_s_arrmul24_fa20_18_y4, h_s_arrmul24_fa21_18_y2, h_s_arrmul24_fa21_18_y4);
  and_gate and_gate_h_s_arrmul24_and22_18_y0(a_22, b_18, h_s_arrmul24_and22_18_y0);
  fa fa_h_s_arrmul24_fa22_18_y2(h_s_arrmul24_and22_18_y0, h_s_arrmul24_fa23_17_y2, h_s_arrmul24_fa21_18_y4, h_s_arrmul24_fa22_18_y2, h_s_arrmul24_fa22_18_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_18_y0(a_23, b_18, h_s_arrmul24_nand23_18_y0);
  fa fa_h_s_arrmul24_fa23_18_y2(h_s_arrmul24_nand23_18_y0, h_s_arrmul24_fa23_17_y4, h_s_arrmul24_fa22_18_y4, h_s_arrmul24_fa23_18_y2, h_s_arrmul24_fa23_18_y4);
  and_gate and_gate_h_s_arrmul24_and0_19_y0(a_0, b_19, h_s_arrmul24_and0_19_y0);
  ha ha_h_s_arrmul24_ha0_19_y0(h_s_arrmul24_and0_19_y0, h_s_arrmul24_fa1_18_y2, h_s_arrmul24_ha0_19_y0, h_s_arrmul24_ha0_19_y1);
  and_gate and_gate_h_s_arrmul24_and1_19_y0(a_1, b_19, h_s_arrmul24_and1_19_y0);
  fa fa_h_s_arrmul24_fa1_19_y2(h_s_arrmul24_and1_19_y0, h_s_arrmul24_fa2_18_y2, h_s_arrmul24_ha0_19_y1, h_s_arrmul24_fa1_19_y2, h_s_arrmul24_fa1_19_y4);
  and_gate and_gate_h_s_arrmul24_and2_19_y0(a_2, b_19, h_s_arrmul24_and2_19_y0);
  fa fa_h_s_arrmul24_fa2_19_y2(h_s_arrmul24_and2_19_y0, h_s_arrmul24_fa3_18_y2, h_s_arrmul24_fa1_19_y4, h_s_arrmul24_fa2_19_y2, h_s_arrmul24_fa2_19_y4);
  and_gate and_gate_h_s_arrmul24_and3_19_y0(a_3, b_19, h_s_arrmul24_and3_19_y0);
  fa fa_h_s_arrmul24_fa3_19_y2(h_s_arrmul24_and3_19_y0, h_s_arrmul24_fa4_18_y2, h_s_arrmul24_fa2_19_y4, h_s_arrmul24_fa3_19_y2, h_s_arrmul24_fa3_19_y4);
  and_gate and_gate_h_s_arrmul24_and4_19_y0(a_4, b_19, h_s_arrmul24_and4_19_y0);
  fa fa_h_s_arrmul24_fa4_19_y2(h_s_arrmul24_and4_19_y0, h_s_arrmul24_fa5_18_y2, h_s_arrmul24_fa3_19_y4, h_s_arrmul24_fa4_19_y2, h_s_arrmul24_fa4_19_y4);
  and_gate and_gate_h_s_arrmul24_and5_19_y0(a_5, b_19, h_s_arrmul24_and5_19_y0);
  fa fa_h_s_arrmul24_fa5_19_y2(h_s_arrmul24_and5_19_y0, h_s_arrmul24_fa6_18_y2, h_s_arrmul24_fa4_19_y4, h_s_arrmul24_fa5_19_y2, h_s_arrmul24_fa5_19_y4);
  and_gate and_gate_h_s_arrmul24_and6_19_y0(a_6, b_19, h_s_arrmul24_and6_19_y0);
  fa fa_h_s_arrmul24_fa6_19_y2(h_s_arrmul24_and6_19_y0, h_s_arrmul24_fa7_18_y2, h_s_arrmul24_fa5_19_y4, h_s_arrmul24_fa6_19_y2, h_s_arrmul24_fa6_19_y4);
  and_gate and_gate_h_s_arrmul24_and7_19_y0(a_7, b_19, h_s_arrmul24_and7_19_y0);
  fa fa_h_s_arrmul24_fa7_19_y2(h_s_arrmul24_and7_19_y0, h_s_arrmul24_fa8_18_y2, h_s_arrmul24_fa6_19_y4, h_s_arrmul24_fa7_19_y2, h_s_arrmul24_fa7_19_y4);
  and_gate and_gate_h_s_arrmul24_and8_19_y0(a_8, b_19, h_s_arrmul24_and8_19_y0);
  fa fa_h_s_arrmul24_fa8_19_y2(h_s_arrmul24_and8_19_y0, h_s_arrmul24_fa9_18_y2, h_s_arrmul24_fa7_19_y4, h_s_arrmul24_fa8_19_y2, h_s_arrmul24_fa8_19_y4);
  and_gate and_gate_h_s_arrmul24_and9_19_y0(a_9, b_19, h_s_arrmul24_and9_19_y0);
  fa fa_h_s_arrmul24_fa9_19_y2(h_s_arrmul24_and9_19_y0, h_s_arrmul24_fa10_18_y2, h_s_arrmul24_fa8_19_y4, h_s_arrmul24_fa9_19_y2, h_s_arrmul24_fa9_19_y4);
  and_gate and_gate_h_s_arrmul24_and10_19_y0(a_10, b_19, h_s_arrmul24_and10_19_y0);
  fa fa_h_s_arrmul24_fa10_19_y2(h_s_arrmul24_and10_19_y0, h_s_arrmul24_fa11_18_y2, h_s_arrmul24_fa9_19_y4, h_s_arrmul24_fa10_19_y2, h_s_arrmul24_fa10_19_y4);
  and_gate and_gate_h_s_arrmul24_and11_19_y0(a_11, b_19, h_s_arrmul24_and11_19_y0);
  fa fa_h_s_arrmul24_fa11_19_y2(h_s_arrmul24_and11_19_y0, h_s_arrmul24_fa12_18_y2, h_s_arrmul24_fa10_19_y4, h_s_arrmul24_fa11_19_y2, h_s_arrmul24_fa11_19_y4);
  and_gate and_gate_h_s_arrmul24_and12_19_y0(a_12, b_19, h_s_arrmul24_and12_19_y0);
  fa fa_h_s_arrmul24_fa12_19_y2(h_s_arrmul24_and12_19_y0, h_s_arrmul24_fa13_18_y2, h_s_arrmul24_fa11_19_y4, h_s_arrmul24_fa12_19_y2, h_s_arrmul24_fa12_19_y4);
  and_gate and_gate_h_s_arrmul24_and13_19_y0(a_13, b_19, h_s_arrmul24_and13_19_y0);
  fa fa_h_s_arrmul24_fa13_19_y2(h_s_arrmul24_and13_19_y0, h_s_arrmul24_fa14_18_y2, h_s_arrmul24_fa12_19_y4, h_s_arrmul24_fa13_19_y2, h_s_arrmul24_fa13_19_y4);
  and_gate and_gate_h_s_arrmul24_and14_19_y0(a_14, b_19, h_s_arrmul24_and14_19_y0);
  fa fa_h_s_arrmul24_fa14_19_y2(h_s_arrmul24_and14_19_y0, h_s_arrmul24_fa15_18_y2, h_s_arrmul24_fa13_19_y4, h_s_arrmul24_fa14_19_y2, h_s_arrmul24_fa14_19_y4);
  and_gate and_gate_h_s_arrmul24_and15_19_y0(a_15, b_19, h_s_arrmul24_and15_19_y0);
  fa fa_h_s_arrmul24_fa15_19_y2(h_s_arrmul24_and15_19_y0, h_s_arrmul24_fa16_18_y2, h_s_arrmul24_fa14_19_y4, h_s_arrmul24_fa15_19_y2, h_s_arrmul24_fa15_19_y4);
  and_gate and_gate_h_s_arrmul24_and16_19_y0(a_16, b_19, h_s_arrmul24_and16_19_y0);
  fa fa_h_s_arrmul24_fa16_19_y2(h_s_arrmul24_and16_19_y0, h_s_arrmul24_fa17_18_y2, h_s_arrmul24_fa15_19_y4, h_s_arrmul24_fa16_19_y2, h_s_arrmul24_fa16_19_y4);
  and_gate and_gate_h_s_arrmul24_and17_19_y0(a_17, b_19, h_s_arrmul24_and17_19_y0);
  fa fa_h_s_arrmul24_fa17_19_y2(h_s_arrmul24_and17_19_y0, h_s_arrmul24_fa18_18_y2, h_s_arrmul24_fa16_19_y4, h_s_arrmul24_fa17_19_y2, h_s_arrmul24_fa17_19_y4);
  and_gate and_gate_h_s_arrmul24_and18_19_y0(a_18, b_19, h_s_arrmul24_and18_19_y0);
  fa fa_h_s_arrmul24_fa18_19_y2(h_s_arrmul24_and18_19_y0, h_s_arrmul24_fa19_18_y2, h_s_arrmul24_fa17_19_y4, h_s_arrmul24_fa18_19_y2, h_s_arrmul24_fa18_19_y4);
  and_gate and_gate_h_s_arrmul24_and19_19_y0(a_19, b_19, h_s_arrmul24_and19_19_y0);
  fa fa_h_s_arrmul24_fa19_19_y2(h_s_arrmul24_and19_19_y0, h_s_arrmul24_fa20_18_y2, h_s_arrmul24_fa18_19_y4, h_s_arrmul24_fa19_19_y2, h_s_arrmul24_fa19_19_y4);
  and_gate and_gate_h_s_arrmul24_and20_19_y0(a_20, b_19, h_s_arrmul24_and20_19_y0);
  fa fa_h_s_arrmul24_fa20_19_y2(h_s_arrmul24_and20_19_y0, h_s_arrmul24_fa21_18_y2, h_s_arrmul24_fa19_19_y4, h_s_arrmul24_fa20_19_y2, h_s_arrmul24_fa20_19_y4);
  and_gate and_gate_h_s_arrmul24_and21_19_y0(a_21, b_19, h_s_arrmul24_and21_19_y0);
  fa fa_h_s_arrmul24_fa21_19_y2(h_s_arrmul24_and21_19_y0, h_s_arrmul24_fa22_18_y2, h_s_arrmul24_fa20_19_y4, h_s_arrmul24_fa21_19_y2, h_s_arrmul24_fa21_19_y4);
  and_gate and_gate_h_s_arrmul24_and22_19_y0(a_22, b_19, h_s_arrmul24_and22_19_y0);
  fa fa_h_s_arrmul24_fa22_19_y2(h_s_arrmul24_and22_19_y0, h_s_arrmul24_fa23_18_y2, h_s_arrmul24_fa21_19_y4, h_s_arrmul24_fa22_19_y2, h_s_arrmul24_fa22_19_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_19_y0(a_23, b_19, h_s_arrmul24_nand23_19_y0);
  fa fa_h_s_arrmul24_fa23_19_y2(h_s_arrmul24_nand23_19_y0, h_s_arrmul24_fa23_18_y4, h_s_arrmul24_fa22_19_y4, h_s_arrmul24_fa23_19_y2, h_s_arrmul24_fa23_19_y4);
  and_gate and_gate_h_s_arrmul24_and0_20_y0(a_0, b_20, h_s_arrmul24_and0_20_y0);
  ha ha_h_s_arrmul24_ha0_20_y0(h_s_arrmul24_and0_20_y0, h_s_arrmul24_fa1_19_y2, h_s_arrmul24_ha0_20_y0, h_s_arrmul24_ha0_20_y1);
  and_gate and_gate_h_s_arrmul24_and1_20_y0(a_1, b_20, h_s_arrmul24_and1_20_y0);
  fa fa_h_s_arrmul24_fa1_20_y2(h_s_arrmul24_and1_20_y0, h_s_arrmul24_fa2_19_y2, h_s_arrmul24_ha0_20_y1, h_s_arrmul24_fa1_20_y2, h_s_arrmul24_fa1_20_y4);
  and_gate and_gate_h_s_arrmul24_and2_20_y0(a_2, b_20, h_s_arrmul24_and2_20_y0);
  fa fa_h_s_arrmul24_fa2_20_y2(h_s_arrmul24_and2_20_y0, h_s_arrmul24_fa3_19_y2, h_s_arrmul24_fa1_20_y4, h_s_arrmul24_fa2_20_y2, h_s_arrmul24_fa2_20_y4);
  and_gate and_gate_h_s_arrmul24_and3_20_y0(a_3, b_20, h_s_arrmul24_and3_20_y0);
  fa fa_h_s_arrmul24_fa3_20_y2(h_s_arrmul24_and3_20_y0, h_s_arrmul24_fa4_19_y2, h_s_arrmul24_fa2_20_y4, h_s_arrmul24_fa3_20_y2, h_s_arrmul24_fa3_20_y4);
  and_gate and_gate_h_s_arrmul24_and4_20_y0(a_4, b_20, h_s_arrmul24_and4_20_y0);
  fa fa_h_s_arrmul24_fa4_20_y2(h_s_arrmul24_and4_20_y0, h_s_arrmul24_fa5_19_y2, h_s_arrmul24_fa3_20_y4, h_s_arrmul24_fa4_20_y2, h_s_arrmul24_fa4_20_y4);
  and_gate and_gate_h_s_arrmul24_and5_20_y0(a_5, b_20, h_s_arrmul24_and5_20_y0);
  fa fa_h_s_arrmul24_fa5_20_y2(h_s_arrmul24_and5_20_y0, h_s_arrmul24_fa6_19_y2, h_s_arrmul24_fa4_20_y4, h_s_arrmul24_fa5_20_y2, h_s_arrmul24_fa5_20_y4);
  and_gate and_gate_h_s_arrmul24_and6_20_y0(a_6, b_20, h_s_arrmul24_and6_20_y0);
  fa fa_h_s_arrmul24_fa6_20_y2(h_s_arrmul24_and6_20_y0, h_s_arrmul24_fa7_19_y2, h_s_arrmul24_fa5_20_y4, h_s_arrmul24_fa6_20_y2, h_s_arrmul24_fa6_20_y4);
  and_gate and_gate_h_s_arrmul24_and7_20_y0(a_7, b_20, h_s_arrmul24_and7_20_y0);
  fa fa_h_s_arrmul24_fa7_20_y2(h_s_arrmul24_and7_20_y0, h_s_arrmul24_fa8_19_y2, h_s_arrmul24_fa6_20_y4, h_s_arrmul24_fa7_20_y2, h_s_arrmul24_fa7_20_y4);
  and_gate and_gate_h_s_arrmul24_and8_20_y0(a_8, b_20, h_s_arrmul24_and8_20_y0);
  fa fa_h_s_arrmul24_fa8_20_y2(h_s_arrmul24_and8_20_y0, h_s_arrmul24_fa9_19_y2, h_s_arrmul24_fa7_20_y4, h_s_arrmul24_fa8_20_y2, h_s_arrmul24_fa8_20_y4);
  and_gate and_gate_h_s_arrmul24_and9_20_y0(a_9, b_20, h_s_arrmul24_and9_20_y0);
  fa fa_h_s_arrmul24_fa9_20_y2(h_s_arrmul24_and9_20_y0, h_s_arrmul24_fa10_19_y2, h_s_arrmul24_fa8_20_y4, h_s_arrmul24_fa9_20_y2, h_s_arrmul24_fa9_20_y4);
  and_gate and_gate_h_s_arrmul24_and10_20_y0(a_10, b_20, h_s_arrmul24_and10_20_y0);
  fa fa_h_s_arrmul24_fa10_20_y2(h_s_arrmul24_and10_20_y0, h_s_arrmul24_fa11_19_y2, h_s_arrmul24_fa9_20_y4, h_s_arrmul24_fa10_20_y2, h_s_arrmul24_fa10_20_y4);
  and_gate and_gate_h_s_arrmul24_and11_20_y0(a_11, b_20, h_s_arrmul24_and11_20_y0);
  fa fa_h_s_arrmul24_fa11_20_y2(h_s_arrmul24_and11_20_y0, h_s_arrmul24_fa12_19_y2, h_s_arrmul24_fa10_20_y4, h_s_arrmul24_fa11_20_y2, h_s_arrmul24_fa11_20_y4);
  and_gate and_gate_h_s_arrmul24_and12_20_y0(a_12, b_20, h_s_arrmul24_and12_20_y0);
  fa fa_h_s_arrmul24_fa12_20_y2(h_s_arrmul24_and12_20_y0, h_s_arrmul24_fa13_19_y2, h_s_arrmul24_fa11_20_y4, h_s_arrmul24_fa12_20_y2, h_s_arrmul24_fa12_20_y4);
  and_gate and_gate_h_s_arrmul24_and13_20_y0(a_13, b_20, h_s_arrmul24_and13_20_y0);
  fa fa_h_s_arrmul24_fa13_20_y2(h_s_arrmul24_and13_20_y0, h_s_arrmul24_fa14_19_y2, h_s_arrmul24_fa12_20_y4, h_s_arrmul24_fa13_20_y2, h_s_arrmul24_fa13_20_y4);
  and_gate and_gate_h_s_arrmul24_and14_20_y0(a_14, b_20, h_s_arrmul24_and14_20_y0);
  fa fa_h_s_arrmul24_fa14_20_y2(h_s_arrmul24_and14_20_y0, h_s_arrmul24_fa15_19_y2, h_s_arrmul24_fa13_20_y4, h_s_arrmul24_fa14_20_y2, h_s_arrmul24_fa14_20_y4);
  and_gate and_gate_h_s_arrmul24_and15_20_y0(a_15, b_20, h_s_arrmul24_and15_20_y0);
  fa fa_h_s_arrmul24_fa15_20_y2(h_s_arrmul24_and15_20_y0, h_s_arrmul24_fa16_19_y2, h_s_arrmul24_fa14_20_y4, h_s_arrmul24_fa15_20_y2, h_s_arrmul24_fa15_20_y4);
  and_gate and_gate_h_s_arrmul24_and16_20_y0(a_16, b_20, h_s_arrmul24_and16_20_y0);
  fa fa_h_s_arrmul24_fa16_20_y2(h_s_arrmul24_and16_20_y0, h_s_arrmul24_fa17_19_y2, h_s_arrmul24_fa15_20_y4, h_s_arrmul24_fa16_20_y2, h_s_arrmul24_fa16_20_y4);
  and_gate and_gate_h_s_arrmul24_and17_20_y0(a_17, b_20, h_s_arrmul24_and17_20_y0);
  fa fa_h_s_arrmul24_fa17_20_y2(h_s_arrmul24_and17_20_y0, h_s_arrmul24_fa18_19_y2, h_s_arrmul24_fa16_20_y4, h_s_arrmul24_fa17_20_y2, h_s_arrmul24_fa17_20_y4);
  and_gate and_gate_h_s_arrmul24_and18_20_y0(a_18, b_20, h_s_arrmul24_and18_20_y0);
  fa fa_h_s_arrmul24_fa18_20_y2(h_s_arrmul24_and18_20_y0, h_s_arrmul24_fa19_19_y2, h_s_arrmul24_fa17_20_y4, h_s_arrmul24_fa18_20_y2, h_s_arrmul24_fa18_20_y4);
  and_gate and_gate_h_s_arrmul24_and19_20_y0(a_19, b_20, h_s_arrmul24_and19_20_y0);
  fa fa_h_s_arrmul24_fa19_20_y2(h_s_arrmul24_and19_20_y0, h_s_arrmul24_fa20_19_y2, h_s_arrmul24_fa18_20_y4, h_s_arrmul24_fa19_20_y2, h_s_arrmul24_fa19_20_y4);
  and_gate and_gate_h_s_arrmul24_and20_20_y0(a_20, b_20, h_s_arrmul24_and20_20_y0);
  fa fa_h_s_arrmul24_fa20_20_y2(h_s_arrmul24_and20_20_y0, h_s_arrmul24_fa21_19_y2, h_s_arrmul24_fa19_20_y4, h_s_arrmul24_fa20_20_y2, h_s_arrmul24_fa20_20_y4);
  and_gate and_gate_h_s_arrmul24_and21_20_y0(a_21, b_20, h_s_arrmul24_and21_20_y0);
  fa fa_h_s_arrmul24_fa21_20_y2(h_s_arrmul24_and21_20_y0, h_s_arrmul24_fa22_19_y2, h_s_arrmul24_fa20_20_y4, h_s_arrmul24_fa21_20_y2, h_s_arrmul24_fa21_20_y4);
  and_gate and_gate_h_s_arrmul24_and22_20_y0(a_22, b_20, h_s_arrmul24_and22_20_y0);
  fa fa_h_s_arrmul24_fa22_20_y2(h_s_arrmul24_and22_20_y0, h_s_arrmul24_fa23_19_y2, h_s_arrmul24_fa21_20_y4, h_s_arrmul24_fa22_20_y2, h_s_arrmul24_fa22_20_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_20_y0(a_23, b_20, h_s_arrmul24_nand23_20_y0);
  fa fa_h_s_arrmul24_fa23_20_y2(h_s_arrmul24_nand23_20_y0, h_s_arrmul24_fa23_19_y4, h_s_arrmul24_fa22_20_y4, h_s_arrmul24_fa23_20_y2, h_s_arrmul24_fa23_20_y4);
  and_gate and_gate_h_s_arrmul24_and0_21_y0(a_0, b_21, h_s_arrmul24_and0_21_y0);
  ha ha_h_s_arrmul24_ha0_21_y0(h_s_arrmul24_and0_21_y0, h_s_arrmul24_fa1_20_y2, h_s_arrmul24_ha0_21_y0, h_s_arrmul24_ha0_21_y1);
  and_gate and_gate_h_s_arrmul24_and1_21_y0(a_1, b_21, h_s_arrmul24_and1_21_y0);
  fa fa_h_s_arrmul24_fa1_21_y2(h_s_arrmul24_and1_21_y0, h_s_arrmul24_fa2_20_y2, h_s_arrmul24_ha0_21_y1, h_s_arrmul24_fa1_21_y2, h_s_arrmul24_fa1_21_y4);
  and_gate and_gate_h_s_arrmul24_and2_21_y0(a_2, b_21, h_s_arrmul24_and2_21_y0);
  fa fa_h_s_arrmul24_fa2_21_y2(h_s_arrmul24_and2_21_y0, h_s_arrmul24_fa3_20_y2, h_s_arrmul24_fa1_21_y4, h_s_arrmul24_fa2_21_y2, h_s_arrmul24_fa2_21_y4);
  and_gate and_gate_h_s_arrmul24_and3_21_y0(a_3, b_21, h_s_arrmul24_and3_21_y0);
  fa fa_h_s_arrmul24_fa3_21_y2(h_s_arrmul24_and3_21_y0, h_s_arrmul24_fa4_20_y2, h_s_arrmul24_fa2_21_y4, h_s_arrmul24_fa3_21_y2, h_s_arrmul24_fa3_21_y4);
  and_gate and_gate_h_s_arrmul24_and4_21_y0(a_4, b_21, h_s_arrmul24_and4_21_y0);
  fa fa_h_s_arrmul24_fa4_21_y2(h_s_arrmul24_and4_21_y0, h_s_arrmul24_fa5_20_y2, h_s_arrmul24_fa3_21_y4, h_s_arrmul24_fa4_21_y2, h_s_arrmul24_fa4_21_y4);
  and_gate and_gate_h_s_arrmul24_and5_21_y0(a_5, b_21, h_s_arrmul24_and5_21_y0);
  fa fa_h_s_arrmul24_fa5_21_y2(h_s_arrmul24_and5_21_y0, h_s_arrmul24_fa6_20_y2, h_s_arrmul24_fa4_21_y4, h_s_arrmul24_fa5_21_y2, h_s_arrmul24_fa5_21_y4);
  and_gate and_gate_h_s_arrmul24_and6_21_y0(a_6, b_21, h_s_arrmul24_and6_21_y0);
  fa fa_h_s_arrmul24_fa6_21_y2(h_s_arrmul24_and6_21_y0, h_s_arrmul24_fa7_20_y2, h_s_arrmul24_fa5_21_y4, h_s_arrmul24_fa6_21_y2, h_s_arrmul24_fa6_21_y4);
  and_gate and_gate_h_s_arrmul24_and7_21_y0(a_7, b_21, h_s_arrmul24_and7_21_y0);
  fa fa_h_s_arrmul24_fa7_21_y2(h_s_arrmul24_and7_21_y0, h_s_arrmul24_fa8_20_y2, h_s_arrmul24_fa6_21_y4, h_s_arrmul24_fa7_21_y2, h_s_arrmul24_fa7_21_y4);
  and_gate and_gate_h_s_arrmul24_and8_21_y0(a_8, b_21, h_s_arrmul24_and8_21_y0);
  fa fa_h_s_arrmul24_fa8_21_y2(h_s_arrmul24_and8_21_y0, h_s_arrmul24_fa9_20_y2, h_s_arrmul24_fa7_21_y4, h_s_arrmul24_fa8_21_y2, h_s_arrmul24_fa8_21_y4);
  and_gate and_gate_h_s_arrmul24_and9_21_y0(a_9, b_21, h_s_arrmul24_and9_21_y0);
  fa fa_h_s_arrmul24_fa9_21_y2(h_s_arrmul24_and9_21_y0, h_s_arrmul24_fa10_20_y2, h_s_arrmul24_fa8_21_y4, h_s_arrmul24_fa9_21_y2, h_s_arrmul24_fa9_21_y4);
  and_gate and_gate_h_s_arrmul24_and10_21_y0(a_10, b_21, h_s_arrmul24_and10_21_y0);
  fa fa_h_s_arrmul24_fa10_21_y2(h_s_arrmul24_and10_21_y0, h_s_arrmul24_fa11_20_y2, h_s_arrmul24_fa9_21_y4, h_s_arrmul24_fa10_21_y2, h_s_arrmul24_fa10_21_y4);
  and_gate and_gate_h_s_arrmul24_and11_21_y0(a_11, b_21, h_s_arrmul24_and11_21_y0);
  fa fa_h_s_arrmul24_fa11_21_y2(h_s_arrmul24_and11_21_y0, h_s_arrmul24_fa12_20_y2, h_s_arrmul24_fa10_21_y4, h_s_arrmul24_fa11_21_y2, h_s_arrmul24_fa11_21_y4);
  and_gate and_gate_h_s_arrmul24_and12_21_y0(a_12, b_21, h_s_arrmul24_and12_21_y0);
  fa fa_h_s_arrmul24_fa12_21_y2(h_s_arrmul24_and12_21_y0, h_s_arrmul24_fa13_20_y2, h_s_arrmul24_fa11_21_y4, h_s_arrmul24_fa12_21_y2, h_s_arrmul24_fa12_21_y4);
  and_gate and_gate_h_s_arrmul24_and13_21_y0(a_13, b_21, h_s_arrmul24_and13_21_y0);
  fa fa_h_s_arrmul24_fa13_21_y2(h_s_arrmul24_and13_21_y0, h_s_arrmul24_fa14_20_y2, h_s_arrmul24_fa12_21_y4, h_s_arrmul24_fa13_21_y2, h_s_arrmul24_fa13_21_y4);
  and_gate and_gate_h_s_arrmul24_and14_21_y0(a_14, b_21, h_s_arrmul24_and14_21_y0);
  fa fa_h_s_arrmul24_fa14_21_y2(h_s_arrmul24_and14_21_y0, h_s_arrmul24_fa15_20_y2, h_s_arrmul24_fa13_21_y4, h_s_arrmul24_fa14_21_y2, h_s_arrmul24_fa14_21_y4);
  and_gate and_gate_h_s_arrmul24_and15_21_y0(a_15, b_21, h_s_arrmul24_and15_21_y0);
  fa fa_h_s_arrmul24_fa15_21_y2(h_s_arrmul24_and15_21_y0, h_s_arrmul24_fa16_20_y2, h_s_arrmul24_fa14_21_y4, h_s_arrmul24_fa15_21_y2, h_s_arrmul24_fa15_21_y4);
  and_gate and_gate_h_s_arrmul24_and16_21_y0(a_16, b_21, h_s_arrmul24_and16_21_y0);
  fa fa_h_s_arrmul24_fa16_21_y2(h_s_arrmul24_and16_21_y0, h_s_arrmul24_fa17_20_y2, h_s_arrmul24_fa15_21_y4, h_s_arrmul24_fa16_21_y2, h_s_arrmul24_fa16_21_y4);
  and_gate and_gate_h_s_arrmul24_and17_21_y0(a_17, b_21, h_s_arrmul24_and17_21_y0);
  fa fa_h_s_arrmul24_fa17_21_y2(h_s_arrmul24_and17_21_y0, h_s_arrmul24_fa18_20_y2, h_s_arrmul24_fa16_21_y4, h_s_arrmul24_fa17_21_y2, h_s_arrmul24_fa17_21_y4);
  and_gate and_gate_h_s_arrmul24_and18_21_y0(a_18, b_21, h_s_arrmul24_and18_21_y0);
  fa fa_h_s_arrmul24_fa18_21_y2(h_s_arrmul24_and18_21_y0, h_s_arrmul24_fa19_20_y2, h_s_arrmul24_fa17_21_y4, h_s_arrmul24_fa18_21_y2, h_s_arrmul24_fa18_21_y4);
  and_gate and_gate_h_s_arrmul24_and19_21_y0(a_19, b_21, h_s_arrmul24_and19_21_y0);
  fa fa_h_s_arrmul24_fa19_21_y2(h_s_arrmul24_and19_21_y0, h_s_arrmul24_fa20_20_y2, h_s_arrmul24_fa18_21_y4, h_s_arrmul24_fa19_21_y2, h_s_arrmul24_fa19_21_y4);
  and_gate and_gate_h_s_arrmul24_and20_21_y0(a_20, b_21, h_s_arrmul24_and20_21_y0);
  fa fa_h_s_arrmul24_fa20_21_y2(h_s_arrmul24_and20_21_y0, h_s_arrmul24_fa21_20_y2, h_s_arrmul24_fa19_21_y4, h_s_arrmul24_fa20_21_y2, h_s_arrmul24_fa20_21_y4);
  and_gate and_gate_h_s_arrmul24_and21_21_y0(a_21, b_21, h_s_arrmul24_and21_21_y0);
  fa fa_h_s_arrmul24_fa21_21_y2(h_s_arrmul24_and21_21_y0, h_s_arrmul24_fa22_20_y2, h_s_arrmul24_fa20_21_y4, h_s_arrmul24_fa21_21_y2, h_s_arrmul24_fa21_21_y4);
  and_gate and_gate_h_s_arrmul24_and22_21_y0(a_22, b_21, h_s_arrmul24_and22_21_y0);
  fa fa_h_s_arrmul24_fa22_21_y2(h_s_arrmul24_and22_21_y0, h_s_arrmul24_fa23_20_y2, h_s_arrmul24_fa21_21_y4, h_s_arrmul24_fa22_21_y2, h_s_arrmul24_fa22_21_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_21_y0(a_23, b_21, h_s_arrmul24_nand23_21_y0);
  fa fa_h_s_arrmul24_fa23_21_y2(h_s_arrmul24_nand23_21_y0, h_s_arrmul24_fa23_20_y4, h_s_arrmul24_fa22_21_y4, h_s_arrmul24_fa23_21_y2, h_s_arrmul24_fa23_21_y4);
  and_gate and_gate_h_s_arrmul24_and0_22_y0(a_0, b_22, h_s_arrmul24_and0_22_y0);
  ha ha_h_s_arrmul24_ha0_22_y0(h_s_arrmul24_and0_22_y0, h_s_arrmul24_fa1_21_y2, h_s_arrmul24_ha0_22_y0, h_s_arrmul24_ha0_22_y1);
  and_gate and_gate_h_s_arrmul24_and1_22_y0(a_1, b_22, h_s_arrmul24_and1_22_y0);
  fa fa_h_s_arrmul24_fa1_22_y2(h_s_arrmul24_and1_22_y0, h_s_arrmul24_fa2_21_y2, h_s_arrmul24_ha0_22_y1, h_s_arrmul24_fa1_22_y2, h_s_arrmul24_fa1_22_y4);
  and_gate and_gate_h_s_arrmul24_and2_22_y0(a_2, b_22, h_s_arrmul24_and2_22_y0);
  fa fa_h_s_arrmul24_fa2_22_y2(h_s_arrmul24_and2_22_y0, h_s_arrmul24_fa3_21_y2, h_s_arrmul24_fa1_22_y4, h_s_arrmul24_fa2_22_y2, h_s_arrmul24_fa2_22_y4);
  and_gate and_gate_h_s_arrmul24_and3_22_y0(a_3, b_22, h_s_arrmul24_and3_22_y0);
  fa fa_h_s_arrmul24_fa3_22_y2(h_s_arrmul24_and3_22_y0, h_s_arrmul24_fa4_21_y2, h_s_arrmul24_fa2_22_y4, h_s_arrmul24_fa3_22_y2, h_s_arrmul24_fa3_22_y4);
  and_gate and_gate_h_s_arrmul24_and4_22_y0(a_4, b_22, h_s_arrmul24_and4_22_y0);
  fa fa_h_s_arrmul24_fa4_22_y2(h_s_arrmul24_and4_22_y0, h_s_arrmul24_fa5_21_y2, h_s_arrmul24_fa3_22_y4, h_s_arrmul24_fa4_22_y2, h_s_arrmul24_fa4_22_y4);
  and_gate and_gate_h_s_arrmul24_and5_22_y0(a_5, b_22, h_s_arrmul24_and5_22_y0);
  fa fa_h_s_arrmul24_fa5_22_y2(h_s_arrmul24_and5_22_y0, h_s_arrmul24_fa6_21_y2, h_s_arrmul24_fa4_22_y4, h_s_arrmul24_fa5_22_y2, h_s_arrmul24_fa5_22_y4);
  and_gate and_gate_h_s_arrmul24_and6_22_y0(a_6, b_22, h_s_arrmul24_and6_22_y0);
  fa fa_h_s_arrmul24_fa6_22_y2(h_s_arrmul24_and6_22_y0, h_s_arrmul24_fa7_21_y2, h_s_arrmul24_fa5_22_y4, h_s_arrmul24_fa6_22_y2, h_s_arrmul24_fa6_22_y4);
  and_gate and_gate_h_s_arrmul24_and7_22_y0(a_7, b_22, h_s_arrmul24_and7_22_y0);
  fa fa_h_s_arrmul24_fa7_22_y2(h_s_arrmul24_and7_22_y0, h_s_arrmul24_fa8_21_y2, h_s_arrmul24_fa6_22_y4, h_s_arrmul24_fa7_22_y2, h_s_arrmul24_fa7_22_y4);
  and_gate and_gate_h_s_arrmul24_and8_22_y0(a_8, b_22, h_s_arrmul24_and8_22_y0);
  fa fa_h_s_arrmul24_fa8_22_y2(h_s_arrmul24_and8_22_y0, h_s_arrmul24_fa9_21_y2, h_s_arrmul24_fa7_22_y4, h_s_arrmul24_fa8_22_y2, h_s_arrmul24_fa8_22_y4);
  and_gate and_gate_h_s_arrmul24_and9_22_y0(a_9, b_22, h_s_arrmul24_and9_22_y0);
  fa fa_h_s_arrmul24_fa9_22_y2(h_s_arrmul24_and9_22_y0, h_s_arrmul24_fa10_21_y2, h_s_arrmul24_fa8_22_y4, h_s_arrmul24_fa9_22_y2, h_s_arrmul24_fa9_22_y4);
  and_gate and_gate_h_s_arrmul24_and10_22_y0(a_10, b_22, h_s_arrmul24_and10_22_y0);
  fa fa_h_s_arrmul24_fa10_22_y2(h_s_arrmul24_and10_22_y0, h_s_arrmul24_fa11_21_y2, h_s_arrmul24_fa9_22_y4, h_s_arrmul24_fa10_22_y2, h_s_arrmul24_fa10_22_y4);
  and_gate and_gate_h_s_arrmul24_and11_22_y0(a_11, b_22, h_s_arrmul24_and11_22_y0);
  fa fa_h_s_arrmul24_fa11_22_y2(h_s_arrmul24_and11_22_y0, h_s_arrmul24_fa12_21_y2, h_s_arrmul24_fa10_22_y4, h_s_arrmul24_fa11_22_y2, h_s_arrmul24_fa11_22_y4);
  and_gate and_gate_h_s_arrmul24_and12_22_y0(a_12, b_22, h_s_arrmul24_and12_22_y0);
  fa fa_h_s_arrmul24_fa12_22_y2(h_s_arrmul24_and12_22_y0, h_s_arrmul24_fa13_21_y2, h_s_arrmul24_fa11_22_y4, h_s_arrmul24_fa12_22_y2, h_s_arrmul24_fa12_22_y4);
  and_gate and_gate_h_s_arrmul24_and13_22_y0(a_13, b_22, h_s_arrmul24_and13_22_y0);
  fa fa_h_s_arrmul24_fa13_22_y2(h_s_arrmul24_and13_22_y0, h_s_arrmul24_fa14_21_y2, h_s_arrmul24_fa12_22_y4, h_s_arrmul24_fa13_22_y2, h_s_arrmul24_fa13_22_y4);
  and_gate and_gate_h_s_arrmul24_and14_22_y0(a_14, b_22, h_s_arrmul24_and14_22_y0);
  fa fa_h_s_arrmul24_fa14_22_y2(h_s_arrmul24_and14_22_y0, h_s_arrmul24_fa15_21_y2, h_s_arrmul24_fa13_22_y4, h_s_arrmul24_fa14_22_y2, h_s_arrmul24_fa14_22_y4);
  and_gate and_gate_h_s_arrmul24_and15_22_y0(a_15, b_22, h_s_arrmul24_and15_22_y0);
  fa fa_h_s_arrmul24_fa15_22_y2(h_s_arrmul24_and15_22_y0, h_s_arrmul24_fa16_21_y2, h_s_arrmul24_fa14_22_y4, h_s_arrmul24_fa15_22_y2, h_s_arrmul24_fa15_22_y4);
  and_gate and_gate_h_s_arrmul24_and16_22_y0(a_16, b_22, h_s_arrmul24_and16_22_y0);
  fa fa_h_s_arrmul24_fa16_22_y2(h_s_arrmul24_and16_22_y0, h_s_arrmul24_fa17_21_y2, h_s_arrmul24_fa15_22_y4, h_s_arrmul24_fa16_22_y2, h_s_arrmul24_fa16_22_y4);
  and_gate and_gate_h_s_arrmul24_and17_22_y0(a_17, b_22, h_s_arrmul24_and17_22_y0);
  fa fa_h_s_arrmul24_fa17_22_y2(h_s_arrmul24_and17_22_y0, h_s_arrmul24_fa18_21_y2, h_s_arrmul24_fa16_22_y4, h_s_arrmul24_fa17_22_y2, h_s_arrmul24_fa17_22_y4);
  and_gate and_gate_h_s_arrmul24_and18_22_y0(a_18, b_22, h_s_arrmul24_and18_22_y0);
  fa fa_h_s_arrmul24_fa18_22_y2(h_s_arrmul24_and18_22_y0, h_s_arrmul24_fa19_21_y2, h_s_arrmul24_fa17_22_y4, h_s_arrmul24_fa18_22_y2, h_s_arrmul24_fa18_22_y4);
  and_gate and_gate_h_s_arrmul24_and19_22_y0(a_19, b_22, h_s_arrmul24_and19_22_y0);
  fa fa_h_s_arrmul24_fa19_22_y2(h_s_arrmul24_and19_22_y0, h_s_arrmul24_fa20_21_y2, h_s_arrmul24_fa18_22_y4, h_s_arrmul24_fa19_22_y2, h_s_arrmul24_fa19_22_y4);
  and_gate and_gate_h_s_arrmul24_and20_22_y0(a_20, b_22, h_s_arrmul24_and20_22_y0);
  fa fa_h_s_arrmul24_fa20_22_y2(h_s_arrmul24_and20_22_y0, h_s_arrmul24_fa21_21_y2, h_s_arrmul24_fa19_22_y4, h_s_arrmul24_fa20_22_y2, h_s_arrmul24_fa20_22_y4);
  and_gate and_gate_h_s_arrmul24_and21_22_y0(a_21, b_22, h_s_arrmul24_and21_22_y0);
  fa fa_h_s_arrmul24_fa21_22_y2(h_s_arrmul24_and21_22_y0, h_s_arrmul24_fa22_21_y2, h_s_arrmul24_fa20_22_y4, h_s_arrmul24_fa21_22_y2, h_s_arrmul24_fa21_22_y4);
  and_gate and_gate_h_s_arrmul24_and22_22_y0(a_22, b_22, h_s_arrmul24_and22_22_y0);
  fa fa_h_s_arrmul24_fa22_22_y2(h_s_arrmul24_and22_22_y0, h_s_arrmul24_fa23_21_y2, h_s_arrmul24_fa21_22_y4, h_s_arrmul24_fa22_22_y2, h_s_arrmul24_fa22_22_y4);
  nand_gate nand_gate_h_s_arrmul24_nand23_22_y0(a_23, b_22, h_s_arrmul24_nand23_22_y0);
  fa fa_h_s_arrmul24_fa23_22_y2(h_s_arrmul24_nand23_22_y0, h_s_arrmul24_fa23_21_y4, h_s_arrmul24_fa22_22_y4, h_s_arrmul24_fa23_22_y2, h_s_arrmul24_fa23_22_y4);
  nand_gate nand_gate_h_s_arrmul24_nand0_23_y0(a_0, b_23, h_s_arrmul24_nand0_23_y0);
  ha ha_h_s_arrmul24_ha0_23_y0(h_s_arrmul24_nand0_23_y0, h_s_arrmul24_fa1_22_y2, h_s_arrmul24_ha0_23_y0, h_s_arrmul24_ha0_23_y1);
  nand_gate nand_gate_h_s_arrmul24_nand1_23_y0(a_1, b_23, h_s_arrmul24_nand1_23_y0);
  fa fa_h_s_arrmul24_fa1_23_y2(h_s_arrmul24_nand1_23_y0, h_s_arrmul24_fa2_22_y2, h_s_arrmul24_ha0_23_y1, h_s_arrmul24_fa1_23_y2, h_s_arrmul24_fa1_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand2_23_y0(a_2, b_23, h_s_arrmul24_nand2_23_y0);
  fa fa_h_s_arrmul24_fa2_23_y2(h_s_arrmul24_nand2_23_y0, h_s_arrmul24_fa3_22_y2, h_s_arrmul24_fa1_23_y4, h_s_arrmul24_fa2_23_y2, h_s_arrmul24_fa2_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand3_23_y0(a_3, b_23, h_s_arrmul24_nand3_23_y0);
  fa fa_h_s_arrmul24_fa3_23_y2(h_s_arrmul24_nand3_23_y0, h_s_arrmul24_fa4_22_y2, h_s_arrmul24_fa2_23_y4, h_s_arrmul24_fa3_23_y2, h_s_arrmul24_fa3_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand4_23_y0(a_4, b_23, h_s_arrmul24_nand4_23_y0);
  fa fa_h_s_arrmul24_fa4_23_y2(h_s_arrmul24_nand4_23_y0, h_s_arrmul24_fa5_22_y2, h_s_arrmul24_fa3_23_y4, h_s_arrmul24_fa4_23_y2, h_s_arrmul24_fa4_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand5_23_y0(a_5, b_23, h_s_arrmul24_nand5_23_y0);
  fa fa_h_s_arrmul24_fa5_23_y2(h_s_arrmul24_nand5_23_y0, h_s_arrmul24_fa6_22_y2, h_s_arrmul24_fa4_23_y4, h_s_arrmul24_fa5_23_y2, h_s_arrmul24_fa5_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand6_23_y0(a_6, b_23, h_s_arrmul24_nand6_23_y0);
  fa fa_h_s_arrmul24_fa6_23_y2(h_s_arrmul24_nand6_23_y0, h_s_arrmul24_fa7_22_y2, h_s_arrmul24_fa5_23_y4, h_s_arrmul24_fa6_23_y2, h_s_arrmul24_fa6_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand7_23_y0(a_7, b_23, h_s_arrmul24_nand7_23_y0);
  fa fa_h_s_arrmul24_fa7_23_y2(h_s_arrmul24_nand7_23_y0, h_s_arrmul24_fa8_22_y2, h_s_arrmul24_fa6_23_y4, h_s_arrmul24_fa7_23_y2, h_s_arrmul24_fa7_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand8_23_y0(a_8, b_23, h_s_arrmul24_nand8_23_y0);
  fa fa_h_s_arrmul24_fa8_23_y2(h_s_arrmul24_nand8_23_y0, h_s_arrmul24_fa9_22_y2, h_s_arrmul24_fa7_23_y4, h_s_arrmul24_fa8_23_y2, h_s_arrmul24_fa8_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand9_23_y0(a_9, b_23, h_s_arrmul24_nand9_23_y0);
  fa fa_h_s_arrmul24_fa9_23_y2(h_s_arrmul24_nand9_23_y0, h_s_arrmul24_fa10_22_y2, h_s_arrmul24_fa8_23_y4, h_s_arrmul24_fa9_23_y2, h_s_arrmul24_fa9_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand10_23_y0(a_10, b_23, h_s_arrmul24_nand10_23_y0);
  fa fa_h_s_arrmul24_fa10_23_y2(h_s_arrmul24_nand10_23_y0, h_s_arrmul24_fa11_22_y2, h_s_arrmul24_fa9_23_y4, h_s_arrmul24_fa10_23_y2, h_s_arrmul24_fa10_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand11_23_y0(a_11, b_23, h_s_arrmul24_nand11_23_y0);
  fa fa_h_s_arrmul24_fa11_23_y2(h_s_arrmul24_nand11_23_y0, h_s_arrmul24_fa12_22_y2, h_s_arrmul24_fa10_23_y4, h_s_arrmul24_fa11_23_y2, h_s_arrmul24_fa11_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand12_23_y0(a_12, b_23, h_s_arrmul24_nand12_23_y0);
  fa fa_h_s_arrmul24_fa12_23_y2(h_s_arrmul24_nand12_23_y0, h_s_arrmul24_fa13_22_y2, h_s_arrmul24_fa11_23_y4, h_s_arrmul24_fa12_23_y2, h_s_arrmul24_fa12_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand13_23_y0(a_13, b_23, h_s_arrmul24_nand13_23_y0);
  fa fa_h_s_arrmul24_fa13_23_y2(h_s_arrmul24_nand13_23_y0, h_s_arrmul24_fa14_22_y2, h_s_arrmul24_fa12_23_y4, h_s_arrmul24_fa13_23_y2, h_s_arrmul24_fa13_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand14_23_y0(a_14, b_23, h_s_arrmul24_nand14_23_y0);
  fa fa_h_s_arrmul24_fa14_23_y2(h_s_arrmul24_nand14_23_y0, h_s_arrmul24_fa15_22_y2, h_s_arrmul24_fa13_23_y4, h_s_arrmul24_fa14_23_y2, h_s_arrmul24_fa14_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand15_23_y0(a_15, b_23, h_s_arrmul24_nand15_23_y0);
  fa fa_h_s_arrmul24_fa15_23_y2(h_s_arrmul24_nand15_23_y0, h_s_arrmul24_fa16_22_y2, h_s_arrmul24_fa14_23_y4, h_s_arrmul24_fa15_23_y2, h_s_arrmul24_fa15_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand16_23_y0(a_16, b_23, h_s_arrmul24_nand16_23_y0);
  fa fa_h_s_arrmul24_fa16_23_y2(h_s_arrmul24_nand16_23_y0, h_s_arrmul24_fa17_22_y2, h_s_arrmul24_fa15_23_y4, h_s_arrmul24_fa16_23_y2, h_s_arrmul24_fa16_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand17_23_y0(a_17, b_23, h_s_arrmul24_nand17_23_y0);
  fa fa_h_s_arrmul24_fa17_23_y2(h_s_arrmul24_nand17_23_y0, h_s_arrmul24_fa18_22_y2, h_s_arrmul24_fa16_23_y4, h_s_arrmul24_fa17_23_y2, h_s_arrmul24_fa17_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand18_23_y0(a_18, b_23, h_s_arrmul24_nand18_23_y0);
  fa fa_h_s_arrmul24_fa18_23_y2(h_s_arrmul24_nand18_23_y0, h_s_arrmul24_fa19_22_y2, h_s_arrmul24_fa17_23_y4, h_s_arrmul24_fa18_23_y2, h_s_arrmul24_fa18_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand19_23_y0(a_19, b_23, h_s_arrmul24_nand19_23_y0);
  fa fa_h_s_arrmul24_fa19_23_y2(h_s_arrmul24_nand19_23_y0, h_s_arrmul24_fa20_22_y2, h_s_arrmul24_fa18_23_y4, h_s_arrmul24_fa19_23_y2, h_s_arrmul24_fa19_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand20_23_y0(a_20, b_23, h_s_arrmul24_nand20_23_y0);
  fa fa_h_s_arrmul24_fa20_23_y2(h_s_arrmul24_nand20_23_y0, h_s_arrmul24_fa21_22_y2, h_s_arrmul24_fa19_23_y4, h_s_arrmul24_fa20_23_y2, h_s_arrmul24_fa20_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand21_23_y0(a_21, b_23, h_s_arrmul24_nand21_23_y0);
  fa fa_h_s_arrmul24_fa21_23_y2(h_s_arrmul24_nand21_23_y0, h_s_arrmul24_fa22_22_y2, h_s_arrmul24_fa20_23_y4, h_s_arrmul24_fa21_23_y2, h_s_arrmul24_fa21_23_y4);
  nand_gate nand_gate_h_s_arrmul24_nand22_23_y0(a_22, b_23, h_s_arrmul24_nand22_23_y0);
  fa fa_h_s_arrmul24_fa22_23_y2(h_s_arrmul24_nand22_23_y0, h_s_arrmul24_fa23_22_y2, h_s_arrmul24_fa21_23_y4, h_s_arrmul24_fa22_23_y2, h_s_arrmul24_fa22_23_y4);
  and_gate and_gate_h_s_arrmul24_and23_23_y0(a_23, b_23, h_s_arrmul24_and23_23_y0);
  fa fa_h_s_arrmul24_fa23_23_y2(h_s_arrmul24_and23_23_y0, h_s_arrmul24_fa23_22_y4, h_s_arrmul24_fa22_23_y4, h_s_arrmul24_fa23_23_y2, h_s_arrmul24_fa23_23_y4);
  xor_gate xor_gate_h_s_arrmul24_xor24_23_y0(h_s_arrmul24_fa23_23_y4, constant_wire_1, h_s_arrmul24_xor24_23_y0);

  assign out[0] = h_s_arrmul24_and0_0_y0;
  assign out[1] = h_s_arrmul24_ha0_1_y0;
  assign out[2] = h_s_arrmul24_ha0_2_y0;
  assign out[3] = h_s_arrmul24_ha0_3_y0;
  assign out[4] = h_s_arrmul24_ha0_4_y0;
  assign out[5] = h_s_arrmul24_ha0_5_y0;
  assign out[6] = h_s_arrmul24_ha0_6_y0;
  assign out[7] = h_s_arrmul24_ha0_7_y0;
  assign out[8] = h_s_arrmul24_ha0_8_y0;
  assign out[9] = h_s_arrmul24_ha0_9_y0;
  assign out[10] = h_s_arrmul24_ha0_10_y0;
  assign out[11] = h_s_arrmul24_ha0_11_y0;
  assign out[12] = h_s_arrmul24_ha0_12_y0;
  assign out[13] = h_s_arrmul24_ha0_13_y0;
  assign out[14] = h_s_arrmul24_ha0_14_y0;
  assign out[15] = h_s_arrmul24_ha0_15_y0;
  assign out[16] = h_s_arrmul24_ha0_16_y0;
  assign out[17] = h_s_arrmul24_ha0_17_y0;
  assign out[18] = h_s_arrmul24_ha0_18_y0;
  assign out[19] = h_s_arrmul24_ha0_19_y0;
  assign out[20] = h_s_arrmul24_ha0_20_y0;
  assign out[21] = h_s_arrmul24_ha0_21_y0;
  assign out[22] = h_s_arrmul24_ha0_22_y0;
  assign out[23] = h_s_arrmul24_ha0_23_y0;
  assign out[24] = h_s_arrmul24_fa1_23_y2;
  assign out[25] = h_s_arrmul24_fa2_23_y2;
  assign out[26] = h_s_arrmul24_fa3_23_y2;
  assign out[27] = h_s_arrmul24_fa4_23_y2;
  assign out[28] = h_s_arrmul24_fa5_23_y2;
  assign out[29] = h_s_arrmul24_fa6_23_y2;
  assign out[30] = h_s_arrmul24_fa7_23_y2;
  assign out[31] = h_s_arrmul24_fa8_23_y2;
  assign out[32] = h_s_arrmul24_fa9_23_y2;
  assign out[33] = h_s_arrmul24_fa10_23_y2;
  assign out[34] = h_s_arrmul24_fa11_23_y2;
  assign out[35] = h_s_arrmul24_fa12_23_y2;
  assign out[36] = h_s_arrmul24_fa13_23_y2;
  assign out[37] = h_s_arrmul24_fa14_23_y2;
  assign out[38] = h_s_arrmul24_fa15_23_y2;
  assign out[39] = h_s_arrmul24_fa16_23_y2;
  assign out[40] = h_s_arrmul24_fa17_23_y2;
  assign out[41] = h_s_arrmul24_fa18_23_y2;
  assign out[42] = h_s_arrmul24_fa19_23_y2;
  assign out[43] = h_s_arrmul24_fa20_23_y2;
  assign out[44] = h_s_arrmul24_fa21_23_y2;
  assign out[45] = h_s_arrmul24_fa22_23_y2;
  assign out[46] = h_s_arrmul24_fa23_23_y2;
  assign out[47] = h_s_arrmul24_xor24_23_y0;
endmodule