module f_s_dadda_rca24(input [23:0] a, input [23:0] b, output [47:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire a_16;
  wire a_17;
  wire a_18;
  wire a_19;
  wire a_20;
  wire a_21;
  wire a_22;
  wire a_23;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire b_16;
  wire b_17;
  wire b_18;
  wire b_19;
  wire b_20;
  wire b_21;
  wire b_22;
  wire b_23;
  wire constant_wire_value_1_a_0;
  wire constant_wire_value_1_b_0;
  wire constant_wire_value_1_y0;
  wire constant_wire_value_1_y1;
  wire constant_wire_1;
  wire f_s_dadda_rca24_and_19_0_a_19;
  wire f_s_dadda_rca24_and_19_0_b_0;
  wire f_s_dadda_rca24_and_19_0_y0;
  wire f_s_dadda_rca24_and_18_1_a_18;
  wire f_s_dadda_rca24_and_18_1_b_1;
  wire f_s_dadda_rca24_and_18_1_y0;
  wire f_s_dadda_rca24_ha0_f_s_dadda_rca24_and_19_0_y0;
  wire f_s_dadda_rca24_ha0_f_s_dadda_rca24_and_18_1_y0;
  wire f_s_dadda_rca24_ha0_y0;
  wire f_s_dadda_rca24_ha0_y1;
  wire f_s_dadda_rca24_and_20_0_a_20;
  wire f_s_dadda_rca24_and_20_0_b_0;
  wire f_s_dadda_rca24_and_20_0_y0;
  wire f_s_dadda_rca24_and_19_1_a_19;
  wire f_s_dadda_rca24_and_19_1_b_1;
  wire f_s_dadda_rca24_and_19_1_y0;
  wire f_s_dadda_rca24_fa0_f_s_dadda_rca24_ha0_y1;
  wire f_s_dadda_rca24_fa0_f_s_dadda_rca24_and_20_0_y0;
  wire f_s_dadda_rca24_fa0_y0;
  wire f_s_dadda_rca24_fa0_y1;
  wire f_s_dadda_rca24_fa0_f_s_dadda_rca24_and_19_1_y0;
  wire f_s_dadda_rca24_fa0_y2;
  wire f_s_dadda_rca24_fa0_y3;
  wire f_s_dadda_rca24_fa0_y4;
  wire f_s_dadda_rca24_and_18_2_a_18;
  wire f_s_dadda_rca24_and_18_2_b_2;
  wire f_s_dadda_rca24_and_18_2_y0;
  wire f_s_dadda_rca24_and_17_3_a_17;
  wire f_s_dadda_rca24_and_17_3_b_3;
  wire f_s_dadda_rca24_and_17_3_y0;
  wire f_s_dadda_rca24_ha1_f_s_dadda_rca24_and_18_2_y0;
  wire f_s_dadda_rca24_ha1_f_s_dadda_rca24_and_17_3_y0;
  wire f_s_dadda_rca24_ha1_y0;
  wire f_s_dadda_rca24_ha1_y1;
  wire f_s_dadda_rca24_and_21_0_a_21;
  wire f_s_dadda_rca24_and_21_0_b_0;
  wire f_s_dadda_rca24_and_21_0_y0;
  wire f_s_dadda_rca24_fa1_f_s_dadda_rca24_ha1_y1;
  wire f_s_dadda_rca24_fa1_f_s_dadda_rca24_fa0_y4;
  wire f_s_dadda_rca24_fa1_y0;
  wire f_s_dadda_rca24_fa1_y1;
  wire f_s_dadda_rca24_fa1_f_s_dadda_rca24_and_21_0_y0;
  wire f_s_dadda_rca24_fa1_y2;
  wire f_s_dadda_rca24_fa1_y3;
  wire f_s_dadda_rca24_fa1_y4;
  wire f_s_dadda_rca24_and_20_1_a_20;
  wire f_s_dadda_rca24_and_20_1_b_1;
  wire f_s_dadda_rca24_and_20_1_y0;
  wire f_s_dadda_rca24_and_19_2_a_19;
  wire f_s_dadda_rca24_and_19_2_b_2;
  wire f_s_dadda_rca24_and_19_2_y0;
  wire f_s_dadda_rca24_and_18_3_a_18;
  wire f_s_dadda_rca24_and_18_3_b_3;
  wire f_s_dadda_rca24_and_18_3_y0;
  wire f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_20_1_y0;
  wire f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_19_2_y0;
  wire f_s_dadda_rca24_fa2_y0;
  wire f_s_dadda_rca24_fa2_y1;
  wire f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_18_3_y0;
  wire f_s_dadda_rca24_fa2_y2;
  wire f_s_dadda_rca24_fa2_y3;
  wire f_s_dadda_rca24_fa2_y4;
  wire f_s_dadda_rca24_and_17_4_a_17;
  wire f_s_dadda_rca24_and_17_4_b_4;
  wire f_s_dadda_rca24_and_17_4_y0;
  wire f_s_dadda_rca24_and_16_5_a_16;
  wire f_s_dadda_rca24_and_16_5_b_5;
  wire f_s_dadda_rca24_and_16_5_y0;
  wire f_s_dadda_rca24_ha2_f_s_dadda_rca24_and_17_4_y0;
  wire f_s_dadda_rca24_ha2_f_s_dadda_rca24_and_16_5_y0;
  wire f_s_dadda_rca24_ha2_y0;
  wire f_s_dadda_rca24_ha2_y1;
  wire f_s_dadda_rca24_fa3_f_s_dadda_rca24_ha2_y1;
  wire f_s_dadda_rca24_fa3_f_s_dadda_rca24_fa2_y4;
  wire f_s_dadda_rca24_fa3_y0;
  wire f_s_dadda_rca24_fa3_y1;
  wire f_s_dadda_rca24_fa3_f_s_dadda_rca24_fa1_y4;
  wire f_s_dadda_rca24_fa3_y2;
  wire f_s_dadda_rca24_fa3_y3;
  wire f_s_dadda_rca24_fa3_y4;
  wire f_s_dadda_rca24_and_22_0_a_22;
  wire f_s_dadda_rca24_and_22_0_b_0;
  wire f_s_dadda_rca24_and_22_0_y0;
  wire f_s_dadda_rca24_and_21_1_a_21;
  wire f_s_dadda_rca24_and_21_1_b_1;
  wire f_s_dadda_rca24_and_21_1_y0;
  wire f_s_dadda_rca24_and_20_2_a_20;
  wire f_s_dadda_rca24_and_20_2_b_2;
  wire f_s_dadda_rca24_and_20_2_y0;
  wire f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_22_0_y0;
  wire f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_21_1_y0;
  wire f_s_dadda_rca24_fa4_y0;
  wire f_s_dadda_rca24_fa4_y1;
  wire f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_20_2_y0;
  wire f_s_dadda_rca24_fa4_y2;
  wire f_s_dadda_rca24_fa4_y3;
  wire f_s_dadda_rca24_fa4_y4;
  wire f_s_dadda_rca24_and_19_3_a_19;
  wire f_s_dadda_rca24_and_19_3_b_3;
  wire f_s_dadda_rca24_and_19_3_y0;
  wire f_s_dadda_rca24_and_18_4_a_18;
  wire f_s_dadda_rca24_and_18_4_b_4;
  wire f_s_dadda_rca24_and_18_4_y0;
  wire f_s_dadda_rca24_and_17_5_a_17;
  wire f_s_dadda_rca24_and_17_5_b_5;
  wire f_s_dadda_rca24_and_17_5_y0;
  wire f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_19_3_y0;
  wire f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_18_4_y0;
  wire f_s_dadda_rca24_fa5_y0;
  wire f_s_dadda_rca24_fa5_y1;
  wire f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_17_5_y0;
  wire f_s_dadda_rca24_fa5_y2;
  wire f_s_dadda_rca24_fa5_y3;
  wire f_s_dadda_rca24_fa5_y4;
  wire f_s_dadda_rca24_and_16_6_a_16;
  wire f_s_dadda_rca24_and_16_6_b_6;
  wire f_s_dadda_rca24_and_16_6_y0;
  wire f_s_dadda_rca24_and_15_7_a_15;
  wire f_s_dadda_rca24_and_15_7_b_7;
  wire f_s_dadda_rca24_and_15_7_y0;
  wire f_s_dadda_rca24_ha3_f_s_dadda_rca24_and_16_6_y0;
  wire f_s_dadda_rca24_ha3_f_s_dadda_rca24_and_15_7_y0;
  wire f_s_dadda_rca24_ha3_y0;
  wire f_s_dadda_rca24_ha3_y1;
  wire f_s_dadda_rca24_fa6_f_s_dadda_rca24_ha3_y1;
  wire f_s_dadda_rca24_fa6_f_s_dadda_rca24_fa5_y4;
  wire f_s_dadda_rca24_fa6_y0;
  wire f_s_dadda_rca24_fa6_y1;
  wire f_s_dadda_rca24_fa6_f_s_dadda_rca24_fa4_y4;
  wire f_s_dadda_rca24_fa6_y2;
  wire f_s_dadda_rca24_fa6_y3;
  wire f_s_dadda_rca24_fa6_y4;
  wire f_s_dadda_rca24_nand_23_0_a_23;
  wire f_s_dadda_rca24_nand_23_0_b_0;
  wire f_s_dadda_rca24_nand_23_0_y0;
  wire f_s_dadda_rca24_and_22_1_a_22;
  wire f_s_dadda_rca24_and_22_1_b_1;
  wire f_s_dadda_rca24_and_22_1_y0;
  wire f_s_dadda_rca24_fa7_f_s_dadda_rca24_fa3_y4;
  wire f_s_dadda_rca24_fa7_f_s_dadda_rca24_nand_23_0_y0;
  wire f_s_dadda_rca24_fa7_y0;
  wire f_s_dadda_rca24_fa7_y1;
  wire f_s_dadda_rca24_fa7_f_s_dadda_rca24_and_22_1_y0;
  wire f_s_dadda_rca24_fa7_y2;
  wire f_s_dadda_rca24_fa7_y3;
  wire f_s_dadda_rca24_fa7_y4;
  wire f_s_dadda_rca24_and_21_2_a_21;
  wire f_s_dadda_rca24_and_21_2_b_2;
  wire f_s_dadda_rca24_and_21_2_y0;
  wire f_s_dadda_rca24_and_20_3_a_20;
  wire f_s_dadda_rca24_and_20_3_b_3;
  wire f_s_dadda_rca24_and_20_3_y0;
  wire f_s_dadda_rca24_and_19_4_a_19;
  wire f_s_dadda_rca24_and_19_4_b_4;
  wire f_s_dadda_rca24_and_19_4_y0;
  wire f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_21_2_y0;
  wire f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_20_3_y0;
  wire f_s_dadda_rca24_fa8_y0;
  wire f_s_dadda_rca24_fa8_y1;
  wire f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_19_4_y0;
  wire f_s_dadda_rca24_fa8_y2;
  wire f_s_dadda_rca24_fa8_y3;
  wire f_s_dadda_rca24_fa8_y4;
  wire f_s_dadda_rca24_and_18_5_a_18;
  wire f_s_dadda_rca24_and_18_5_b_5;
  wire f_s_dadda_rca24_and_18_5_y0;
  wire f_s_dadda_rca24_and_17_6_a_17;
  wire f_s_dadda_rca24_and_17_6_b_6;
  wire f_s_dadda_rca24_and_17_6_y0;
  wire f_s_dadda_rca24_and_16_7_a_16;
  wire f_s_dadda_rca24_and_16_7_b_7;
  wire f_s_dadda_rca24_and_16_7_y0;
  wire f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_18_5_y0;
  wire f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_17_6_y0;
  wire f_s_dadda_rca24_fa9_y0;
  wire f_s_dadda_rca24_fa9_y1;
  wire f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_16_7_y0;
  wire f_s_dadda_rca24_fa9_y2;
  wire f_s_dadda_rca24_fa9_y3;
  wire f_s_dadda_rca24_fa9_y4;
  wire f_s_dadda_rca24_and_15_8_a_15;
  wire f_s_dadda_rca24_and_15_8_b_8;
  wire f_s_dadda_rca24_and_15_8_y0;
  wire f_s_dadda_rca24_and_14_9_a_14;
  wire f_s_dadda_rca24_and_14_9_b_9;
  wire f_s_dadda_rca24_and_14_9_y0;
  wire f_s_dadda_rca24_ha4_f_s_dadda_rca24_and_15_8_y0;
  wire f_s_dadda_rca24_ha4_f_s_dadda_rca24_and_14_9_y0;
  wire f_s_dadda_rca24_ha4_y0;
  wire f_s_dadda_rca24_ha4_y1;
  wire f_s_dadda_rca24_fa10_f_s_dadda_rca24_ha4_y1;
  wire f_s_dadda_rca24_fa10_f_s_dadda_rca24_fa9_y4;
  wire f_s_dadda_rca24_fa10_y0;
  wire f_s_dadda_rca24_fa10_y1;
  wire f_s_dadda_rca24_fa10_f_s_dadda_rca24_fa8_y4;
  wire f_s_dadda_rca24_fa10_y2;
  wire f_s_dadda_rca24_fa10_y3;
  wire f_s_dadda_rca24_fa10_y4;
  wire f_s_dadda_rca24_fa11_f_s_dadda_rca24_fa7_y4;
  wire f_s_dadda_rca24_fa11_f_s_dadda_rca24_fa6_y4;
  wire f_s_dadda_rca24_fa11_y0;
  wire f_s_dadda_rca24_fa11_y1;
  wire f_s_dadda_rca24_fa11_constant_wire_1;
  wire f_s_dadda_rca24_fa11_y2;
  wire f_s_dadda_rca24_fa11_y3;
  wire f_s_dadda_rca24_fa11_y4;
  wire f_s_dadda_rca24_nand_23_1_a_23;
  wire f_s_dadda_rca24_nand_23_1_b_1;
  wire f_s_dadda_rca24_nand_23_1_y0;
  wire f_s_dadda_rca24_and_22_2_a_22;
  wire f_s_dadda_rca24_and_22_2_b_2;
  wire f_s_dadda_rca24_and_22_2_y0;
  wire f_s_dadda_rca24_and_21_3_a_21;
  wire f_s_dadda_rca24_and_21_3_b_3;
  wire f_s_dadda_rca24_and_21_3_y0;
  wire f_s_dadda_rca24_fa12_f_s_dadda_rca24_nand_23_1_y0;
  wire f_s_dadda_rca24_fa12_f_s_dadda_rca24_and_22_2_y0;
  wire f_s_dadda_rca24_fa12_y0;
  wire f_s_dadda_rca24_fa12_y1;
  wire f_s_dadda_rca24_fa12_f_s_dadda_rca24_and_21_3_y0;
  wire f_s_dadda_rca24_fa12_y2;
  wire f_s_dadda_rca24_fa12_y3;
  wire f_s_dadda_rca24_fa12_y4;
  wire f_s_dadda_rca24_and_20_4_a_20;
  wire f_s_dadda_rca24_and_20_4_b_4;
  wire f_s_dadda_rca24_and_20_4_y0;
  wire f_s_dadda_rca24_and_19_5_a_19;
  wire f_s_dadda_rca24_and_19_5_b_5;
  wire f_s_dadda_rca24_and_19_5_y0;
  wire f_s_dadda_rca24_and_18_6_a_18;
  wire f_s_dadda_rca24_and_18_6_b_6;
  wire f_s_dadda_rca24_and_18_6_y0;
  wire f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_20_4_y0;
  wire f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_19_5_y0;
  wire f_s_dadda_rca24_fa13_y0;
  wire f_s_dadda_rca24_fa13_y1;
  wire f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_18_6_y0;
  wire f_s_dadda_rca24_fa13_y2;
  wire f_s_dadda_rca24_fa13_y3;
  wire f_s_dadda_rca24_fa13_y4;
  wire f_s_dadda_rca24_and_17_7_a_17;
  wire f_s_dadda_rca24_and_17_7_b_7;
  wire f_s_dadda_rca24_and_17_7_y0;
  wire f_s_dadda_rca24_and_16_8_a_16;
  wire f_s_dadda_rca24_and_16_8_b_8;
  wire f_s_dadda_rca24_and_16_8_y0;
  wire f_s_dadda_rca24_and_15_9_a_15;
  wire f_s_dadda_rca24_and_15_9_b_9;
  wire f_s_dadda_rca24_and_15_9_y0;
  wire f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_17_7_y0;
  wire f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_16_8_y0;
  wire f_s_dadda_rca24_fa14_y0;
  wire f_s_dadda_rca24_fa14_y1;
  wire f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_15_9_y0;
  wire f_s_dadda_rca24_fa14_y2;
  wire f_s_dadda_rca24_fa14_y3;
  wire f_s_dadda_rca24_fa14_y4;
  wire f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa14_y4;
  wire f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa13_y4;
  wire f_s_dadda_rca24_fa15_y0;
  wire f_s_dadda_rca24_fa15_y1;
  wire f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa12_y4;
  wire f_s_dadda_rca24_fa15_y2;
  wire f_s_dadda_rca24_fa15_y3;
  wire f_s_dadda_rca24_fa15_y4;
  wire f_s_dadda_rca24_nand_23_2_a_23;
  wire f_s_dadda_rca24_nand_23_2_b_2;
  wire f_s_dadda_rca24_nand_23_2_y0;
  wire f_s_dadda_rca24_fa16_f_s_dadda_rca24_fa11_y4;
  wire f_s_dadda_rca24_fa16_f_s_dadda_rca24_fa10_y4;
  wire f_s_dadda_rca24_fa16_y0;
  wire f_s_dadda_rca24_fa16_y1;
  wire f_s_dadda_rca24_fa16_f_s_dadda_rca24_nand_23_2_y0;
  wire f_s_dadda_rca24_fa16_y2;
  wire f_s_dadda_rca24_fa16_y3;
  wire f_s_dadda_rca24_fa16_y4;
  wire f_s_dadda_rca24_and_22_3_a_22;
  wire f_s_dadda_rca24_and_22_3_b_3;
  wire f_s_dadda_rca24_and_22_3_y0;
  wire f_s_dadda_rca24_and_21_4_a_21;
  wire f_s_dadda_rca24_and_21_4_b_4;
  wire f_s_dadda_rca24_and_21_4_y0;
  wire f_s_dadda_rca24_and_20_5_a_20;
  wire f_s_dadda_rca24_and_20_5_b_5;
  wire f_s_dadda_rca24_and_20_5_y0;
  wire f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_22_3_y0;
  wire f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_21_4_y0;
  wire f_s_dadda_rca24_fa17_y0;
  wire f_s_dadda_rca24_fa17_y1;
  wire f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_20_5_y0;
  wire f_s_dadda_rca24_fa17_y2;
  wire f_s_dadda_rca24_fa17_y3;
  wire f_s_dadda_rca24_fa17_y4;
  wire f_s_dadda_rca24_and_19_6_a_19;
  wire f_s_dadda_rca24_and_19_6_b_6;
  wire f_s_dadda_rca24_and_19_6_y0;
  wire f_s_dadda_rca24_and_18_7_a_18;
  wire f_s_dadda_rca24_and_18_7_b_7;
  wire f_s_dadda_rca24_and_18_7_y0;
  wire f_s_dadda_rca24_and_17_8_a_17;
  wire f_s_dadda_rca24_and_17_8_b_8;
  wire f_s_dadda_rca24_and_17_8_y0;
  wire f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_19_6_y0;
  wire f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_18_7_y0;
  wire f_s_dadda_rca24_fa18_y0;
  wire f_s_dadda_rca24_fa18_y1;
  wire f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_17_8_y0;
  wire f_s_dadda_rca24_fa18_y2;
  wire f_s_dadda_rca24_fa18_y3;
  wire f_s_dadda_rca24_fa18_y4;
  wire f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa18_y4;
  wire f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa17_y4;
  wire f_s_dadda_rca24_fa19_y0;
  wire f_s_dadda_rca24_fa19_y1;
  wire f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa16_y4;
  wire f_s_dadda_rca24_fa19_y2;
  wire f_s_dadda_rca24_fa19_y3;
  wire f_s_dadda_rca24_fa19_y4;
  wire f_s_dadda_rca24_nand_23_3_a_23;
  wire f_s_dadda_rca24_nand_23_3_b_3;
  wire f_s_dadda_rca24_nand_23_3_y0;
  wire f_s_dadda_rca24_and_22_4_a_22;
  wire f_s_dadda_rca24_and_22_4_b_4;
  wire f_s_dadda_rca24_and_22_4_y0;
  wire f_s_dadda_rca24_fa20_f_s_dadda_rca24_fa15_y4;
  wire f_s_dadda_rca24_fa20_f_s_dadda_rca24_nand_23_3_y0;
  wire f_s_dadda_rca24_fa20_y0;
  wire f_s_dadda_rca24_fa20_y1;
  wire f_s_dadda_rca24_fa20_f_s_dadda_rca24_and_22_4_y0;
  wire f_s_dadda_rca24_fa20_y2;
  wire f_s_dadda_rca24_fa20_y3;
  wire f_s_dadda_rca24_fa20_y4;
  wire f_s_dadda_rca24_and_21_5_a_21;
  wire f_s_dadda_rca24_and_21_5_b_5;
  wire f_s_dadda_rca24_and_21_5_y0;
  wire f_s_dadda_rca24_and_20_6_a_20;
  wire f_s_dadda_rca24_and_20_6_b_6;
  wire f_s_dadda_rca24_and_20_6_y0;
  wire f_s_dadda_rca24_and_19_7_a_19;
  wire f_s_dadda_rca24_and_19_7_b_7;
  wire f_s_dadda_rca24_and_19_7_y0;
  wire f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_21_5_y0;
  wire f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_20_6_y0;
  wire f_s_dadda_rca24_fa21_y0;
  wire f_s_dadda_rca24_fa21_y1;
  wire f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_19_7_y0;
  wire f_s_dadda_rca24_fa21_y2;
  wire f_s_dadda_rca24_fa21_y3;
  wire f_s_dadda_rca24_fa21_y4;
  wire f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa21_y4;
  wire f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa20_y4;
  wire f_s_dadda_rca24_fa22_y0;
  wire f_s_dadda_rca24_fa22_y1;
  wire f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa19_y4;
  wire f_s_dadda_rca24_fa22_y2;
  wire f_s_dadda_rca24_fa22_y3;
  wire f_s_dadda_rca24_fa22_y4;
  wire f_s_dadda_rca24_nand_23_4_a_23;
  wire f_s_dadda_rca24_nand_23_4_b_4;
  wire f_s_dadda_rca24_nand_23_4_y0;
  wire f_s_dadda_rca24_and_22_5_a_22;
  wire f_s_dadda_rca24_and_22_5_b_5;
  wire f_s_dadda_rca24_and_22_5_y0;
  wire f_s_dadda_rca24_and_21_6_a_21;
  wire f_s_dadda_rca24_and_21_6_b_6;
  wire f_s_dadda_rca24_and_21_6_y0;
  wire f_s_dadda_rca24_fa23_f_s_dadda_rca24_nand_23_4_y0;
  wire f_s_dadda_rca24_fa23_f_s_dadda_rca24_and_22_5_y0;
  wire f_s_dadda_rca24_fa23_y0;
  wire f_s_dadda_rca24_fa23_y1;
  wire f_s_dadda_rca24_fa23_f_s_dadda_rca24_and_21_6_y0;
  wire f_s_dadda_rca24_fa23_y2;
  wire f_s_dadda_rca24_fa23_y3;
  wire f_s_dadda_rca24_fa23_y4;
  wire f_s_dadda_rca24_nand_23_5_a_23;
  wire f_s_dadda_rca24_nand_23_5_b_5;
  wire f_s_dadda_rca24_nand_23_5_y0;
  wire f_s_dadda_rca24_fa24_f_s_dadda_rca24_fa23_y4;
  wire f_s_dadda_rca24_fa24_f_s_dadda_rca24_fa22_y4;
  wire f_s_dadda_rca24_fa24_y0;
  wire f_s_dadda_rca24_fa24_y1;
  wire f_s_dadda_rca24_fa24_f_s_dadda_rca24_nand_23_5_y0;
  wire f_s_dadda_rca24_fa24_y2;
  wire f_s_dadda_rca24_fa24_y3;
  wire f_s_dadda_rca24_fa24_y4;
  wire f_s_dadda_rca24_and_6_0_a_6;
  wire f_s_dadda_rca24_and_6_0_b_0;
  wire f_s_dadda_rca24_and_6_0_y0;
  wire f_s_dadda_rca24_and_5_1_a_5;
  wire f_s_dadda_rca24_and_5_1_b_1;
  wire f_s_dadda_rca24_and_5_1_y0;
  wire f_s_dadda_rca24_ha5_f_s_dadda_rca24_and_6_0_y0;
  wire f_s_dadda_rca24_ha5_f_s_dadda_rca24_and_5_1_y0;
  wire f_s_dadda_rca24_ha5_y0;
  wire f_s_dadda_rca24_ha5_y1;
  wire f_s_dadda_rca24_and_7_0_a_7;
  wire f_s_dadda_rca24_and_7_0_b_0;
  wire f_s_dadda_rca24_and_7_0_y0;
  wire f_s_dadda_rca24_and_6_1_a_6;
  wire f_s_dadda_rca24_and_6_1_b_1;
  wire f_s_dadda_rca24_and_6_1_y0;
  wire f_s_dadda_rca24_fa25_f_s_dadda_rca24_ha5_y1;
  wire f_s_dadda_rca24_fa25_f_s_dadda_rca24_and_7_0_y0;
  wire f_s_dadda_rca24_fa25_y0;
  wire f_s_dadda_rca24_fa25_y1;
  wire f_s_dadda_rca24_fa25_f_s_dadda_rca24_and_6_1_y0;
  wire f_s_dadda_rca24_fa25_y2;
  wire f_s_dadda_rca24_fa25_y3;
  wire f_s_dadda_rca24_fa25_y4;
  wire f_s_dadda_rca24_and_5_2_a_5;
  wire f_s_dadda_rca24_and_5_2_b_2;
  wire f_s_dadda_rca24_and_5_2_y0;
  wire f_s_dadda_rca24_and_4_3_a_4;
  wire f_s_dadda_rca24_and_4_3_b_3;
  wire f_s_dadda_rca24_and_4_3_y0;
  wire f_s_dadda_rca24_ha6_f_s_dadda_rca24_and_5_2_y0;
  wire f_s_dadda_rca24_ha6_f_s_dadda_rca24_and_4_3_y0;
  wire f_s_dadda_rca24_ha6_y0;
  wire f_s_dadda_rca24_ha6_y1;
  wire f_s_dadda_rca24_and_8_0_a_8;
  wire f_s_dadda_rca24_and_8_0_b_0;
  wire f_s_dadda_rca24_and_8_0_y0;
  wire f_s_dadda_rca24_fa26_f_s_dadda_rca24_ha6_y1;
  wire f_s_dadda_rca24_fa26_f_s_dadda_rca24_fa25_y4;
  wire f_s_dadda_rca24_fa26_y0;
  wire f_s_dadda_rca24_fa26_y1;
  wire f_s_dadda_rca24_fa26_f_s_dadda_rca24_and_8_0_y0;
  wire f_s_dadda_rca24_fa26_y2;
  wire f_s_dadda_rca24_fa26_y3;
  wire f_s_dadda_rca24_fa26_y4;
  wire f_s_dadda_rca24_and_7_1_a_7;
  wire f_s_dadda_rca24_and_7_1_b_1;
  wire f_s_dadda_rca24_and_7_1_y0;
  wire f_s_dadda_rca24_and_6_2_a_6;
  wire f_s_dadda_rca24_and_6_2_b_2;
  wire f_s_dadda_rca24_and_6_2_y0;
  wire f_s_dadda_rca24_and_5_3_a_5;
  wire f_s_dadda_rca24_and_5_3_b_3;
  wire f_s_dadda_rca24_and_5_3_y0;
  wire f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_7_1_y0;
  wire f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_6_2_y0;
  wire f_s_dadda_rca24_fa27_y0;
  wire f_s_dadda_rca24_fa27_y1;
  wire f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_5_3_y0;
  wire f_s_dadda_rca24_fa27_y2;
  wire f_s_dadda_rca24_fa27_y3;
  wire f_s_dadda_rca24_fa27_y4;
  wire f_s_dadda_rca24_and_4_4_a_4;
  wire f_s_dadda_rca24_and_4_4_b_4;
  wire f_s_dadda_rca24_and_4_4_y0;
  wire f_s_dadda_rca24_and_3_5_a_3;
  wire f_s_dadda_rca24_and_3_5_b_5;
  wire f_s_dadda_rca24_and_3_5_y0;
  wire f_s_dadda_rca24_ha7_f_s_dadda_rca24_and_4_4_y0;
  wire f_s_dadda_rca24_ha7_f_s_dadda_rca24_and_3_5_y0;
  wire f_s_dadda_rca24_ha7_y0;
  wire f_s_dadda_rca24_ha7_y1;
  wire f_s_dadda_rca24_fa28_f_s_dadda_rca24_ha7_y1;
  wire f_s_dadda_rca24_fa28_f_s_dadda_rca24_fa27_y4;
  wire f_s_dadda_rca24_fa28_y0;
  wire f_s_dadda_rca24_fa28_y1;
  wire f_s_dadda_rca24_fa28_f_s_dadda_rca24_fa26_y4;
  wire f_s_dadda_rca24_fa28_y2;
  wire f_s_dadda_rca24_fa28_y3;
  wire f_s_dadda_rca24_fa28_y4;
  wire f_s_dadda_rca24_and_9_0_a_9;
  wire f_s_dadda_rca24_and_9_0_b_0;
  wire f_s_dadda_rca24_and_9_0_y0;
  wire f_s_dadda_rca24_and_8_1_a_8;
  wire f_s_dadda_rca24_and_8_1_b_1;
  wire f_s_dadda_rca24_and_8_1_y0;
  wire f_s_dadda_rca24_and_7_2_a_7;
  wire f_s_dadda_rca24_and_7_2_b_2;
  wire f_s_dadda_rca24_and_7_2_y0;
  wire f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_9_0_y0;
  wire f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_8_1_y0;
  wire f_s_dadda_rca24_fa29_y0;
  wire f_s_dadda_rca24_fa29_y1;
  wire f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_7_2_y0;
  wire f_s_dadda_rca24_fa29_y2;
  wire f_s_dadda_rca24_fa29_y3;
  wire f_s_dadda_rca24_fa29_y4;
  wire f_s_dadda_rca24_and_6_3_a_6;
  wire f_s_dadda_rca24_and_6_3_b_3;
  wire f_s_dadda_rca24_and_6_3_y0;
  wire f_s_dadda_rca24_and_5_4_a_5;
  wire f_s_dadda_rca24_and_5_4_b_4;
  wire f_s_dadda_rca24_and_5_4_y0;
  wire f_s_dadda_rca24_and_4_5_a_4;
  wire f_s_dadda_rca24_and_4_5_b_5;
  wire f_s_dadda_rca24_and_4_5_y0;
  wire f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_6_3_y0;
  wire f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_5_4_y0;
  wire f_s_dadda_rca24_fa30_y0;
  wire f_s_dadda_rca24_fa30_y1;
  wire f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_4_5_y0;
  wire f_s_dadda_rca24_fa30_y2;
  wire f_s_dadda_rca24_fa30_y3;
  wire f_s_dadda_rca24_fa30_y4;
  wire f_s_dadda_rca24_and_3_6_a_3;
  wire f_s_dadda_rca24_and_3_6_b_6;
  wire f_s_dadda_rca24_and_3_6_y0;
  wire f_s_dadda_rca24_and_2_7_a_2;
  wire f_s_dadda_rca24_and_2_7_b_7;
  wire f_s_dadda_rca24_and_2_7_y0;
  wire f_s_dadda_rca24_ha8_f_s_dadda_rca24_and_3_6_y0;
  wire f_s_dadda_rca24_ha8_f_s_dadda_rca24_and_2_7_y0;
  wire f_s_dadda_rca24_ha8_y0;
  wire f_s_dadda_rca24_ha8_y1;
  wire f_s_dadda_rca24_fa31_f_s_dadda_rca24_ha8_y1;
  wire f_s_dadda_rca24_fa31_f_s_dadda_rca24_fa30_y4;
  wire f_s_dadda_rca24_fa31_y0;
  wire f_s_dadda_rca24_fa31_y1;
  wire f_s_dadda_rca24_fa31_f_s_dadda_rca24_fa29_y4;
  wire f_s_dadda_rca24_fa31_y2;
  wire f_s_dadda_rca24_fa31_y3;
  wire f_s_dadda_rca24_fa31_y4;
  wire f_s_dadda_rca24_and_10_0_a_10;
  wire f_s_dadda_rca24_and_10_0_b_0;
  wire f_s_dadda_rca24_and_10_0_y0;
  wire f_s_dadda_rca24_and_9_1_a_9;
  wire f_s_dadda_rca24_and_9_1_b_1;
  wire f_s_dadda_rca24_and_9_1_y0;
  wire f_s_dadda_rca24_fa32_f_s_dadda_rca24_fa28_y4;
  wire f_s_dadda_rca24_fa32_f_s_dadda_rca24_and_10_0_y0;
  wire f_s_dadda_rca24_fa32_y0;
  wire f_s_dadda_rca24_fa32_y1;
  wire f_s_dadda_rca24_fa32_f_s_dadda_rca24_and_9_1_y0;
  wire f_s_dadda_rca24_fa32_y2;
  wire f_s_dadda_rca24_fa32_y3;
  wire f_s_dadda_rca24_fa32_y4;
  wire f_s_dadda_rca24_and_8_2_a_8;
  wire f_s_dadda_rca24_and_8_2_b_2;
  wire f_s_dadda_rca24_and_8_2_y0;
  wire f_s_dadda_rca24_and_7_3_a_7;
  wire f_s_dadda_rca24_and_7_3_b_3;
  wire f_s_dadda_rca24_and_7_3_y0;
  wire f_s_dadda_rca24_and_6_4_a_6;
  wire f_s_dadda_rca24_and_6_4_b_4;
  wire f_s_dadda_rca24_and_6_4_y0;
  wire f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_8_2_y0;
  wire f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_7_3_y0;
  wire f_s_dadda_rca24_fa33_y0;
  wire f_s_dadda_rca24_fa33_y1;
  wire f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_6_4_y0;
  wire f_s_dadda_rca24_fa33_y2;
  wire f_s_dadda_rca24_fa33_y3;
  wire f_s_dadda_rca24_fa33_y4;
  wire f_s_dadda_rca24_and_5_5_a_5;
  wire f_s_dadda_rca24_and_5_5_b_5;
  wire f_s_dadda_rca24_and_5_5_y0;
  wire f_s_dadda_rca24_and_4_6_a_4;
  wire f_s_dadda_rca24_and_4_6_b_6;
  wire f_s_dadda_rca24_and_4_6_y0;
  wire f_s_dadda_rca24_and_3_7_a_3;
  wire f_s_dadda_rca24_and_3_7_b_7;
  wire f_s_dadda_rca24_and_3_7_y0;
  wire f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_5_5_y0;
  wire f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_4_6_y0;
  wire f_s_dadda_rca24_fa34_y0;
  wire f_s_dadda_rca24_fa34_y1;
  wire f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_3_7_y0;
  wire f_s_dadda_rca24_fa34_y2;
  wire f_s_dadda_rca24_fa34_y3;
  wire f_s_dadda_rca24_fa34_y4;
  wire f_s_dadda_rca24_and_2_8_a_2;
  wire f_s_dadda_rca24_and_2_8_b_8;
  wire f_s_dadda_rca24_and_2_8_y0;
  wire f_s_dadda_rca24_and_1_9_a_1;
  wire f_s_dadda_rca24_and_1_9_b_9;
  wire f_s_dadda_rca24_and_1_9_y0;
  wire f_s_dadda_rca24_ha9_f_s_dadda_rca24_and_2_8_y0;
  wire f_s_dadda_rca24_ha9_f_s_dadda_rca24_and_1_9_y0;
  wire f_s_dadda_rca24_ha9_y0;
  wire f_s_dadda_rca24_ha9_y1;
  wire f_s_dadda_rca24_fa35_f_s_dadda_rca24_ha9_y1;
  wire f_s_dadda_rca24_fa35_f_s_dadda_rca24_fa34_y4;
  wire f_s_dadda_rca24_fa35_y0;
  wire f_s_dadda_rca24_fa35_y1;
  wire f_s_dadda_rca24_fa35_f_s_dadda_rca24_fa33_y4;
  wire f_s_dadda_rca24_fa35_y2;
  wire f_s_dadda_rca24_fa35_y3;
  wire f_s_dadda_rca24_fa35_y4;
  wire f_s_dadda_rca24_and_11_0_a_11;
  wire f_s_dadda_rca24_and_11_0_b_0;
  wire f_s_dadda_rca24_and_11_0_y0;
  wire f_s_dadda_rca24_fa36_f_s_dadda_rca24_fa32_y4;
  wire f_s_dadda_rca24_fa36_f_s_dadda_rca24_fa31_y4;
  wire f_s_dadda_rca24_fa36_y0;
  wire f_s_dadda_rca24_fa36_y1;
  wire f_s_dadda_rca24_fa36_f_s_dadda_rca24_and_11_0_y0;
  wire f_s_dadda_rca24_fa36_y2;
  wire f_s_dadda_rca24_fa36_y3;
  wire f_s_dadda_rca24_fa36_y4;
  wire f_s_dadda_rca24_and_10_1_a_10;
  wire f_s_dadda_rca24_and_10_1_b_1;
  wire f_s_dadda_rca24_and_10_1_y0;
  wire f_s_dadda_rca24_and_9_2_a_9;
  wire f_s_dadda_rca24_and_9_2_b_2;
  wire f_s_dadda_rca24_and_9_2_y0;
  wire f_s_dadda_rca24_and_8_3_a_8;
  wire f_s_dadda_rca24_and_8_3_b_3;
  wire f_s_dadda_rca24_and_8_3_y0;
  wire f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_10_1_y0;
  wire f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_9_2_y0;
  wire f_s_dadda_rca24_fa37_y0;
  wire f_s_dadda_rca24_fa37_y1;
  wire f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_8_3_y0;
  wire f_s_dadda_rca24_fa37_y2;
  wire f_s_dadda_rca24_fa37_y3;
  wire f_s_dadda_rca24_fa37_y4;
  wire f_s_dadda_rca24_and_7_4_a_7;
  wire f_s_dadda_rca24_and_7_4_b_4;
  wire f_s_dadda_rca24_and_7_4_y0;
  wire f_s_dadda_rca24_and_6_5_a_6;
  wire f_s_dadda_rca24_and_6_5_b_5;
  wire f_s_dadda_rca24_and_6_5_y0;
  wire f_s_dadda_rca24_and_5_6_a_5;
  wire f_s_dadda_rca24_and_5_6_b_6;
  wire f_s_dadda_rca24_and_5_6_y0;
  wire f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_7_4_y0;
  wire f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_6_5_y0;
  wire f_s_dadda_rca24_fa38_y0;
  wire f_s_dadda_rca24_fa38_y1;
  wire f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_5_6_y0;
  wire f_s_dadda_rca24_fa38_y2;
  wire f_s_dadda_rca24_fa38_y3;
  wire f_s_dadda_rca24_fa38_y4;
  wire f_s_dadda_rca24_and_4_7_a_4;
  wire f_s_dadda_rca24_and_4_7_b_7;
  wire f_s_dadda_rca24_and_4_7_y0;
  wire f_s_dadda_rca24_and_3_8_a_3;
  wire f_s_dadda_rca24_and_3_8_b_8;
  wire f_s_dadda_rca24_and_3_8_y0;
  wire f_s_dadda_rca24_and_2_9_a_2;
  wire f_s_dadda_rca24_and_2_9_b_9;
  wire f_s_dadda_rca24_and_2_9_y0;
  wire f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_4_7_y0;
  wire f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_3_8_y0;
  wire f_s_dadda_rca24_fa39_y0;
  wire f_s_dadda_rca24_fa39_y1;
  wire f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_2_9_y0;
  wire f_s_dadda_rca24_fa39_y2;
  wire f_s_dadda_rca24_fa39_y3;
  wire f_s_dadda_rca24_fa39_y4;
  wire f_s_dadda_rca24_and_1_10_a_1;
  wire f_s_dadda_rca24_and_1_10_b_10;
  wire f_s_dadda_rca24_and_1_10_y0;
  wire f_s_dadda_rca24_and_0_11_a_0;
  wire f_s_dadda_rca24_and_0_11_b_11;
  wire f_s_dadda_rca24_and_0_11_y0;
  wire f_s_dadda_rca24_ha10_f_s_dadda_rca24_and_1_10_y0;
  wire f_s_dadda_rca24_ha10_f_s_dadda_rca24_and_0_11_y0;
  wire f_s_dadda_rca24_ha10_y0;
  wire f_s_dadda_rca24_ha10_y1;
  wire f_s_dadda_rca24_fa40_f_s_dadda_rca24_ha10_y1;
  wire f_s_dadda_rca24_fa40_f_s_dadda_rca24_fa39_y4;
  wire f_s_dadda_rca24_fa40_y0;
  wire f_s_dadda_rca24_fa40_y1;
  wire f_s_dadda_rca24_fa40_f_s_dadda_rca24_fa38_y4;
  wire f_s_dadda_rca24_fa40_y2;
  wire f_s_dadda_rca24_fa40_y3;
  wire f_s_dadda_rca24_fa40_y4;
  wire f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa37_y4;
  wire f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa36_y4;
  wire f_s_dadda_rca24_fa41_y0;
  wire f_s_dadda_rca24_fa41_y1;
  wire f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa35_y4;
  wire f_s_dadda_rca24_fa41_y2;
  wire f_s_dadda_rca24_fa41_y3;
  wire f_s_dadda_rca24_fa41_y4;
  wire f_s_dadda_rca24_and_12_0_a_12;
  wire f_s_dadda_rca24_and_12_0_b_0;
  wire f_s_dadda_rca24_and_12_0_y0;
  wire f_s_dadda_rca24_and_11_1_a_11;
  wire f_s_dadda_rca24_and_11_1_b_1;
  wire f_s_dadda_rca24_and_11_1_y0;
  wire f_s_dadda_rca24_and_10_2_a_10;
  wire f_s_dadda_rca24_and_10_2_b_2;
  wire f_s_dadda_rca24_and_10_2_y0;
  wire f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_12_0_y0;
  wire f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_11_1_y0;
  wire f_s_dadda_rca24_fa42_y0;
  wire f_s_dadda_rca24_fa42_y1;
  wire f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_10_2_y0;
  wire f_s_dadda_rca24_fa42_y2;
  wire f_s_dadda_rca24_fa42_y3;
  wire f_s_dadda_rca24_fa42_y4;
  wire f_s_dadda_rca24_and_9_3_a_9;
  wire f_s_dadda_rca24_and_9_3_b_3;
  wire f_s_dadda_rca24_and_9_3_y0;
  wire f_s_dadda_rca24_and_8_4_a_8;
  wire f_s_dadda_rca24_and_8_4_b_4;
  wire f_s_dadda_rca24_and_8_4_y0;
  wire f_s_dadda_rca24_and_7_5_a_7;
  wire f_s_dadda_rca24_and_7_5_b_5;
  wire f_s_dadda_rca24_and_7_5_y0;
  wire f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_9_3_y0;
  wire f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_8_4_y0;
  wire f_s_dadda_rca24_fa43_y0;
  wire f_s_dadda_rca24_fa43_y1;
  wire f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_7_5_y0;
  wire f_s_dadda_rca24_fa43_y2;
  wire f_s_dadda_rca24_fa43_y3;
  wire f_s_dadda_rca24_fa43_y4;
  wire f_s_dadda_rca24_and_6_6_a_6;
  wire f_s_dadda_rca24_and_6_6_b_6;
  wire f_s_dadda_rca24_and_6_6_y0;
  wire f_s_dadda_rca24_and_5_7_a_5;
  wire f_s_dadda_rca24_and_5_7_b_7;
  wire f_s_dadda_rca24_and_5_7_y0;
  wire f_s_dadda_rca24_and_4_8_a_4;
  wire f_s_dadda_rca24_and_4_8_b_8;
  wire f_s_dadda_rca24_and_4_8_y0;
  wire f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_6_6_y0;
  wire f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_5_7_y0;
  wire f_s_dadda_rca24_fa44_y0;
  wire f_s_dadda_rca24_fa44_y1;
  wire f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_4_8_y0;
  wire f_s_dadda_rca24_fa44_y2;
  wire f_s_dadda_rca24_fa44_y3;
  wire f_s_dadda_rca24_fa44_y4;
  wire f_s_dadda_rca24_and_3_9_a_3;
  wire f_s_dadda_rca24_and_3_9_b_9;
  wire f_s_dadda_rca24_and_3_9_y0;
  wire f_s_dadda_rca24_and_2_10_a_2;
  wire f_s_dadda_rca24_and_2_10_b_10;
  wire f_s_dadda_rca24_and_2_10_y0;
  wire f_s_dadda_rca24_and_1_11_a_1;
  wire f_s_dadda_rca24_and_1_11_b_11;
  wire f_s_dadda_rca24_and_1_11_y0;
  wire f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_3_9_y0;
  wire f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_2_10_y0;
  wire f_s_dadda_rca24_fa45_y0;
  wire f_s_dadda_rca24_fa45_y1;
  wire f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_1_11_y0;
  wire f_s_dadda_rca24_fa45_y2;
  wire f_s_dadda_rca24_fa45_y3;
  wire f_s_dadda_rca24_fa45_y4;
  wire f_s_dadda_rca24_and_0_12_a_0;
  wire f_s_dadda_rca24_and_0_12_b_12;
  wire f_s_dadda_rca24_and_0_12_y0;
  wire f_s_dadda_rca24_ha11_f_s_dadda_rca24_and_0_12_y0;
  wire f_s_dadda_rca24_ha11_f_s_dadda_rca24_fa40_y2;
  wire f_s_dadda_rca24_ha11_y0;
  wire f_s_dadda_rca24_ha11_y1;
  wire f_s_dadda_rca24_fa46_f_s_dadda_rca24_ha11_y1;
  wire f_s_dadda_rca24_fa46_f_s_dadda_rca24_fa45_y4;
  wire f_s_dadda_rca24_fa46_y0;
  wire f_s_dadda_rca24_fa46_y1;
  wire f_s_dadda_rca24_fa46_f_s_dadda_rca24_fa44_y4;
  wire f_s_dadda_rca24_fa46_y2;
  wire f_s_dadda_rca24_fa46_y3;
  wire f_s_dadda_rca24_fa46_y4;
  wire f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa43_y4;
  wire f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa42_y4;
  wire f_s_dadda_rca24_fa47_y0;
  wire f_s_dadda_rca24_fa47_y1;
  wire f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa41_y4;
  wire f_s_dadda_rca24_fa47_y2;
  wire f_s_dadda_rca24_fa47_y3;
  wire f_s_dadda_rca24_fa47_y4;
  wire f_s_dadda_rca24_and_13_0_a_13;
  wire f_s_dadda_rca24_and_13_0_b_0;
  wire f_s_dadda_rca24_and_13_0_y0;
  wire f_s_dadda_rca24_and_12_1_a_12;
  wire f_s_dadda_rca24_and_12_1_b_1;
  wire f_s_dadda_rca24_and_12_1_y0;
  wire f_s_dadda_rca24_fa48_f_s_dadda_rca24_fa40_y4;
  wire f_s_dadda_rca24_fa48_f_s_dadda_rca24_and_13_0_y0;
  wire f_s_dadda_rca24_fa48_y0;
  wire f_s_dadda_rca24_fa48_y1;
  wire f_s_dadda_rca24_fa48_f_s_dadda_rca24_and_12_1_y0;
  wire f_s_dadda_rca24_fa48_y2;
  wire f_s_dadda_rca24_fa48_y3;
  wire f_s_dadda_rca24_fa48_y4;
  wire f_s_dadda_rca24_and_11_2_a_11;
  wire f_s_dadda_rca24_and_11_2_b_2;
  wire f_s_dadda_rca24_and_11_2_y0;
  wire f_s_dadda_rca24_and_10_3_a_10;
  wire f_s_dadda_rca24_and_10_3_b_3;
  wire f_s_dadda_rca24_and_10_3_y0;
  wire f_s_dadda_rca24_and_9_4_a_9;
  wire f_s_dadda_rca24_and_9_4_b_4;
  wire f_s_dadda_rca24_and_9_4_y0;
  wire f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_11_2_y0;
  wire f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_10_3_y0;
  wire f_s_dadda_rca24_fa49_y0;
  wire f_s_dadda_rca24_fa49_y1;
  wire f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_9_4_y0;
  wire f_s_dadda_rca24_fa49_y2;
  wire f_s_dadda_rca24_fa49_y3;
  wire f_s_dadda_rca24_fa49_y4;
  wire f_s_dadda_rca24_and_8_5_a_8;
  wire f_s_dadda_rca24_and_8_5_b_5;
  wire f_s_dadda_rca24_and_8_5_y0;
  wire f_s_dadda_rca24_and_7_6_a_7;
  wire f_s_dadda_rca24_and_7_6_b_6;
  wire f_s_dadda_rca24_and_7_6_y0;
  wire f_s_dadda_rca24_and_6_7_a_6;
  wire f_s_dadda_rca24_and_6_7_b_7;
  wire f_s_dadda_rca24_and_6_7_y0;
  wire f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_8_5_y0;
  wire f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_7_6_y0;
  wire f_s_dadda_rca24_fa50_y0;
  wire f_s_dadda_rca24_fa50_y1;
  wire f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_6_7_y0;
  wire f_s_dadda_rca24_fa50_y2;
  wire f_s_dadda_rca24_fa50_y3;
  wire f_s_dadda_rca24_fa50_y4;
  wire f_s_dadda_rca24_and_5_8_a_5;
  wire f_s_dadda_rca24_and_5_8_b_8;
  wire f_s_dadda_rca24_and_5_8_y0;
  wire f_s_dadda_rca24_and_4_9_a_4;
  wire f_s_dadda_rca24_and_4_9_b_9;
  wire f_s_dadda_rca24_and_4_9_y0;
  wire f_s_dadda_rca24_and_3_10_a_3;
  wire f_s_dadda_rca24_and_3_10_b_10;
  wire f_s_dadda_rca24_and_3_10_y0;
  wire f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_5_8_y0;
  wire f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_4_9_y0;
  wire f_s_dadda_rca24_fa51_y0;
  wire f_s_dadda_rca24_fa51_y1;
  wire f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_3_10_y0;
  wire f_s_dadda_rca24_fa51_y2;
  wire f_s_dadda_rca24_fa51_y3;
  wire f_s_dadda_rca24_fa51_y4;
  wire f_s_dadda_rca24_and_2_11_a_2;
  wire f_s_dadda_rca24_and_2_11_b_11;
  wire f_s_dadda_rca24_and_2_11_y0;
  wire f_s_dadda_rca24_and_1_12_a_1;
  wire f_s_dadda_rca24_and_1_12_b_12;
  wire f_s_dadda_rca24_and_1_12_y0;
  wire f_s_dadda_rca24_and_0_13_a_0;
  wire f_s_dadda_rca24_and_0_13_b_13;
  wire f_s_dadda_rca24_and_0_13_y0;
  wire f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_2_11_y0;
  wire f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_1_12_y0;
  wire f_s_dadda_rca24_fa52_y0;
  wire f_s_dadda_rca24_fa52_y1;
  wire f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_0_13_y0;
  wire f_s_dadda_rca24_fa52_y2;
  wire f_s_dadda_rca24_fa52_y3;
  wire f_s_dadda_rca24_fa52_y4;
  wire f_s_dadda_rca24_ha12_f_s_dadda_rca24_fa46_y2;
  wire f_s_dadda_rca24_ha12_f_s_dadda_rca24_fa47_y2;
  wire f_s_dadda_rca24_ha12_y0;
  wire f_s_dadda_rca24_ha12_y1;
  wire f_s_dadda_rca24_fa53_f_s_dadda_rca24_ha12_y1;
  wire f_s_dadda_rca24_fa53_f_s_dadda_rca24_fa52_y4;
  wire f_s_dadda_rca24_fa53_y0;
  wire f_s_dadda_rca24_fa53_y1;
  wire f_s_dadda_rca24_fa53_f_s_dadda_rca24_fa51_y4;
  wire f_s_dadda_rca24_fa53_y2;
  wire f_s_dadda_rca24_fa53_y3;
  wire f_s_dadda_rca24_fa53_y4;
  wire f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa50_y4;
  wire f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa49_y4;
  wire f_s_dadda_rca24_fa54_y0;
  wire f_s_dadda_rca24_fa54_y1;
  wire f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa48_y4;
  wire f_s_dadda_rca24_fa54_y2;
  wire f_s_dadda_rca24_fa54_y3;
  wire f_s_dadda_rca24_fa54_y4;
  wire f_s_dadda_rca24_and_14_0_a_14;
  wire f_s_dadda_rca24_and_14_0_b_0;
  wire f_s_dadda_rca24_and_14_0_y0;
  wire f_s_dadda_rca24_fa55_f_s_dadda_rca24_fa47_y4;
  wire f_s_dadda_rca24_fa55_f_s_dadda_rca24_fa46_y4;
  wire f_s_dadda_rca24_fa55_y0;
  wire f_s_dadda_rca24_fa55_y1;
  wire f_s_dadda_rca24_fa55_f_s_dadda_rca24_and_14_0_y0;
  wire f_s_dadda_rca24_fa55_y2;
  wire f_s_dadda_rca24_fa55_y3;
  wire f_s_dadda_rca24_fa55_y4;
  wire f_s_dadda_rca24_and_13_1_a_13;
  wire f_s_dadda_rca24_and_13_1_b_1;
  wire f_s_dadda_rca24_and_13_1_y0;
  wire f_s_dadda_rca24_and_12_2_a_12;
  wire f_s_dadda_rca24_and_12_2_b_2;
  wire f_s_dadda_rca24_and_12_2_y0;
  wire f_s_dadda_rca24_and_11_3_a_11;
  wire f_s_dadda_rca24_and_11_3_b_3;
  wire f_s_dadda_rca24_and_11_3_y0;
  wire f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_13_1_y0;
  wire f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_12_2_y0;
  wire f_s_dadda_rca24_fa56_y0;
  wire f_s_dadda_rca24_fa56_y1;
  wire f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_11_3_y0;
  wire f_s_dadda_rca24_fa56_y2;
  wire f_s_dadda_rca24_fa56_y3;
  wire f_s_dadda_rca24_fa56_y4;
  wire f_s_dadda_rca24_and_10_4_a_10;
  wire f_s_dadda_rca24_and_10_4_b_4;
  wire f_s_dadda_rca24_and_10_4_y0;
  wire f_s_dadda_rca24_and_9_5_a_9;
  wire f_s_dadda_rca24_and_9_5_b_5;
  wire f_s_dadda_rca24_and_9_5_y0;
  wire f_s_dadda_rca24_and_8_6_a_8;
  wire f_s_dadda_rca24_and_8_6_b_6;
  wire f_s_dadda_rca24_and_8_6_y0;
  wire f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_10_4_y0;
  wire f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_9_5_y0;
  wire f_s_dadda_rca24_fa57_y0;
  wire f_s_dadda_rca24_fa57_y1;
  wire f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_8_6_y0;
  wire f_s_dadda_rca24_fa57_y2;
  wire f_s_dadda_rca24_fa57_y3;
  wire f_s_dadda_rca24_fa57_y4;
  wire f_s_dadda_rca24_and_7_7_a_7;
  wire f_s_dadda_rca24_and_7_7_b_7;
  wire f_s_dadda_rca24_and_7_7_y0;
  wire f_s_dadda_rca24_and_6_8_a_6;
  wire f_s_dadda_rca24_and_6_8_b_8;
  wire f_s_dadda_rca24_and_6_8_y0;
  wire f_s_dadda_rca24_and_5_9_a_5;
  wire f_s_dadda_rca24_and_5_9_b_9;
  wire f_s_dadda_rca24_and_5_9_y0;
  wire f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_7_7_y0;
  wire f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_6_8_y0;
  wire f_s_dadda_rca24_fa58_y0;
  wire f_s_dadda_rca24_fa58_y1;
  wire f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_5_9_y0;
  wire f_s_dadda_rca24_fa58_y2;
  wire f_s_dadda_rca24_fa58_y3;
  wire f_s_dadda_rca24_fa58_y4;
  wire f_s_dadda_rca24_and_4_10_a_4;
  wire f_s_dadda_rca24_and_4_10_b_10;
  wire f_s_dadda_rca24_and_4_10_y0;
  wire f_s_dadda_rca24_and_3_11_a_3;
  wire f_s_dadda_rca24_and_3_11_b_11;
  wire f_s_dadda_rca24_and_3_11_y0;
  wire f_s_dadda_rca24_and_2_12_a_2;
  wire f_s_dadda_rca24_and_2_12_b_12;
  wire f_s_dadda_rca24_and_2_12_y0;
  wire f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_4_10_y0;
  wire f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_3_11_y0;
  wire f_s_dadda_rca24_fa59_y0;
  wire f_s_dadda_rca24_fa59_y1;
  wire f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_2_12_y0;
  wire f_s_dadda_rca24_fa59_y2;
  wire f_s_dadda_rca24_fa59_y3;
  wire f_s_dadda_rca24_fa59_y4;
  wire f_s_dadda_rca24_and_1_13_a_1;
  wire f_s_dadda_rca24_and_1_13_b_13;
  wire f_s_dadda_rca24_and_1_13_y0;
  wire f_s_dadda_rca24_and_0_14_a_0;
  wire f_s_dadda_rca24_and_0_14_b_14;
  wire f_s_dadda_rca24_and_0_14_y0;
  wire f_s_dadda_rca24_fa60_f_s_dadda_rca24_and_1_13_y0;
  wire f_s_dadda_rca24_fa60_f_s_dadda_rca24_and_0_14_y0;
  wire f_s_dadda_rca24_fa60_y0;
  wire f_s_dadda_rca24_fa60_y1;
  wire f_s_dadda_rca24_fa60_f_s_dadda_rca24_fa53_y2;
  wire f_s_dadda_rca24_fa60_y2;
  wire f_s_dadda_rca24_fa60_y3;
  wire f_s_dadda_rca24_fa60_y4;
  wire f_s_dadda_rca24_ha13_f_s_dadda_rca24_fa54_y2;
  wire f_s_dadda_rca24_ha13_f_s_dadda_rca24_fa55_y2;
  wire f_s_dadda_rca24_ha13_y0;
  wire f_s_dadda_rca24_ha13_y1;
  wire f_s_dadda_rca24_fa61_f_s_dadda_rca24_ha13_y1;
  wire f_s_dadda_rca24_fa61_f_s_dadda_rca24_fa60_y4;
  wire f_s_dadda_rca24_fa61_y0;
  wire f_s_dadda_rca24_fa61_y1;
  wire f_s_dadda_rca24_fa61_f_s_dadda_rca24_fa59_y4;
  wire f_s_dadda_rca24_fa61_y2;
  wire f_s_dadda_rca24_fa61_y3;
  wire f_s_dadda_rca24_fa61_y4;
  wire f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa58_y4;
  wire f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa57_y4;
  wire f_s_dadda_rca24_fa62_y0;
  wire f_s_dadda_rca24_fa62_y1;
  wire f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa56_y4;
  wire f_s_dadda_rca24_fa62_y2;
  wire f_s_dadda_rca24_fa62_y3;
  wire f_s_dadda_rca24_fa62_y4;
  wire f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa55_y4;
  wire f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa54_y4;
  wire f_s_dadda_rca24_fa63_y0;
  wire f_s_dadda_rca24_fa63_y1;
  wire f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa53_y4;
  wire f_s_dadda_rca24_fa63_y2;
  wire f_s_dadda_rca24_fa63_y3;
  wire f_s_dadda_rca24_fa63_y4;
  wire f_s_dadda_rca24_and_15_0_a_15;
  wire f_s_dadda_rca24_and_15_0_b_0;
  wire f_s_dadda_rca24_and_15_0_y0;
  wire f_s_dadda_rca24_and_14_1_a_14;
  wire f_s_dadda_rca24_and_14_1_b_1;
  wire f_s_dadda_rca24_and_14_1_y0;
  wire f_s_dadda_rca24_and_13_2_a_13;
  wire f_s_dadda_rca24_and_13_2_b_2;
  wire f_s_dadda_rca24_and_13_2_y0;
  wire f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_15_0_y0;
  wire f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_14_1_y0;
  wire f_s_dadda_rca24_fa64_y0;
  wire f_s_dadda_rca24_fa64_y1;
  wire f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_13_2_y0;
  wire f_s_dadda_rca24_fa64_y2;
  wire f_s_dadda_rca24_fa64_y3;
  wire f_s_dadda_rca24_fa64_y4;
  wire f_s_dadda_rca24_and_12_3_a_12;
  wire f_s_dadda_rca24_and_12_3_b_3;
  wire f_s_dadda_rca24_and_12_3_y0;
  wire f_s_dadda_rca24_and_11_4_a_11;
  wire f_s_dadda_rca24_and_11_4_b_4;
  wire f_s_dadda_rca24_and_11_4_y0;
  wire f_s_dadda_rca24_and_10_5_a_10;
  wire f_s_dadda_rca24_and_10_5_b_5;
  wire f_s_dadda_rca24_and_10_5_y0;
  wire f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_12_3_y0;
  wire f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_11_4_y0;
  wire f_s_dadda_rca24_fa65_y0;
  wire f_s_dadda_rca24_fa65_y1;
  wire f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_10_5_y0;
  wire f_s_dadda_rca24_fa65_y2;
  wire f_s_dadda_rca24_fa65_y3;
  wire f_s_dadda_rca24_fa65_y4;
  wire f_s_dadda_rca24_and_9_6_a_9;
  wire f_s_dadda_rca24_and_9_6_b_6;
  wire f_s_dadda_rca24_and_9_6_y0;
  wire f_s_dadda_rca24_and_8_7_a_8;
  wire f_s_dadda_rca24_and_8_7_b_7;
  wire f_s_dadda_rca24_and_8_7_y0;
  wire f_s_dadda_rca24_and_7_8_a_7;
  wire f_s_dadda_rca24_and_7_8_b_8;
  wire f_s_dadda_rca24_and_7_8_y0;
  wire f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_9_6_y0;
  wire f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_8_7_y0;
  wire f_s_dadda_rca24_fa66_y0;
  wire f_s_dadda_rca24_fa66_y1;
  wire f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_7_8_y0;
  wire f_s_dadda_rca24_fa66_y2;
  wire f_s_dadda_rca24_fa66_y3;
  wire f_s_dadda_rca24_fa66_y4;
  wire f_s_dadda_rca24_and_6_9_a_6;
  wire f_s_dadda_rca24_and_6_9_b_9;
  wire f_s_dadda_rca24_and_6_9_y0;
  wire f_s_dadda_rca24_and_5_10_a_5;
  wire f_s_dadda_rca24_and_5_10_b_10;
  wire f_s_dadda_rca24_and_5_10_y0;
  wire f_s_dadda_rca24_and_4_11_a_4;
  wire f_s_dadda_rca24_and_4_11_b_11;
  wire f_s_dadda_rca24_and_4_11_y0;
  wire f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_6_9_y0;
  wire f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_5_10_y0;
  wire f_s_dadda_rca24_fa67_y0;
  wire f_s_dadda_rca24_fa67_y1;
  wire f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_4_11_y0;
  wire f_s_dadda_rca24_fa67_y2;
  wire f_s_dadda_rca24_fa67_y3;
  wire f_s_dadda_rca24_fa67_y4;
  wire f_s_dadda_rca24_and_3_12_a_3;
  wire f_s_dadda_rca24_and_3_12_b_12;
  wire f_s_dadda_rca24_and_3_12_y0;
  wire f_s_dadda_rca24_and_2_13_a_2;
  wire f_s_dadda_rca24_and_2_13_b_13;
  wire f_s_dadda_rca24_and_2_13_y0;
  wire f_s_dadda_rca24_and_1_14_a_1;
  wire f_s_dadda_rca24_and_1_14_b_14;
  wire f_s_dadda_rca24_and_1_14_y0;
  wire f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_3_12_y0;
  wire f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_2_13_y0;
  wire f_s_dadda_rca24_fa68_y0;
  wire f_s_dadda_rca24_fa68_y1;
  wire f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_1_14_y0;
  wire f_s_dadda_rca24_fa68_y2;
  wire f_s_dadda_rca24_fa68_y3;
  wire f_s_dadda_rca24_fa68_y4;
  wire f_s_dadda_rca24_and_0_15_a_0;
  wire f_s_dadda_rca24_and_0_15_b_15;
  wire f_s_dadda_rca24_and_0_15_y0;
  wire f_s_dadda_rca24_fa69_f_s_dadda_rca24_and_0_15_y0;
  wire f_s_dadda_rca24_fa69_f_s_dadda_rca24_fa61_y2;
  wire f_s_dadda_rca24_fa69_y0;
  wire f_s_dadda_rca24_fa69_y1;
  wire f_s_dadda_rca24_fa69_f_s_dadda_rca24_fa62_y2;
  wire f_s_dadda_rca24_fa69_y2;
  wire f_s_dadda_rca24_fa69_y3;
  wire f_s_dadda_rca24_fa69_y4;
  wire f_s_dadda_rca24_ha14_f_s_dadda_rca24_fa63_y2;
  wire f_s_dadda_rca24_ha14_f_s_dadda_rca24_fa64_y2;
  wire f_s_dadda_rca24_ha14_y0;
  wire f_s_dadda_rca24_ha14_y1;
  wire f_s_dadda_rca24_fa70_f_s_dadda_rca24_ha14_y1;
  wire f_s_dadda_rca24_fa70_f_s_dadda_rca24_fa69_y4;
  wire f_s_dadda_rca24_fa70_y0;
  wire f_s_dadda_rca24_fa70_y1;
  wire f_s_dadda_rca24_fa70_f_s_dadda_rca24_fa68_y4;
  wire f_s_dadda_rca24_fa70_y2;
  wire f_s_dadda_rca24_fa70_y3;
  wire f_s_dadda_rca24_fa70_y4;
  wire f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa67_y4;
  wire f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa66_y4;
  wire f_s_dadda_rca24_fa71_y0;
  wire f_s_dadda_rca24_fa71_y1;
  wire f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa65_y4;
  wire f_s_dadda_rca24_fa71_y2;
  wire f_s_dadda_rca24_fa71_y3;
  wire f_s_dadda_rca24_fa71_y4;
  wire f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa64_y4;
  wire f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa63_y4;
  wire f_s_dadda_rca24_fa72_y0;
  wire f_s_dadda_rca24_fa72_y1;
  wire f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa62_y4;
  wire f_s_dadda_rca24_fa72_y2;
  wire f_s_dadda_rca24_fa72_y3;
  wire f_s_dadda_rca24_fa72_y4;
  wire f_s_dadda_rca24_and_16_0_a_16;
  wire f_s_dadda_rca24_and_16_0_b_0;
  wire f_s_dadda_rca24_and_16_0_y0;
  wire f_s_dadda_rca24_and_15_1_a_15;
  wire f_s_dadda_rca24_and_15_1_b_1;
  wire f_s_dadda_rca24_and_15_1_y0;
  wire f_s_dadda_rca24_fa73_f_s_dadda_rca24_fa61_y4;
  wire f_s_dadda_rca24_fa73_f_s_dadda_rca24_and_16_0_y0;
  wire f_s_dadda_rca24_fa73_y0;
  wire f_s_dadda_rca24_fa73_y1;
  wire f_s_dadda_rca24_fa73_f_s_dadda_rca24_and_15_1_y0;
  wire f_s_dadda_rca24_fa73_y2;
  wire f_s_dadda_rca24_fa73_y3;
  wire f_s_dadda_rca24_fa73_y4;
  wire f_s_dadda_rca24_and_14_2_a_14;
  wire f_s_dadda_rca24_and_14_2_b_2;
  wire f_s_dadda_rca24_and_14_2_y0;
  wire f_s_dadda_rca24_and_13_3_a_13;
  wire f_s_dadda_rca24_and_13_3_b_3;
  wire f_s_dadda_rca24_and_13_3_y0;
  wire f_s_dadda_rca24_and_12_4_a_12;
  wire f_s_dadda_rca24_and_12_4_b_4;
  wire f_s_dadda_rca24_and_12_4_y0;
  wire f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_14_2_y0;
  wire f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_13_3_y0;
  wire f_s_dadda_rca24_fa74_y0;
  wire f_s_dadda_rca24_fa74_y1;
  wire f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_12_4_y0;
  wire f_s_dadda_rca24_fa74_y2;
  wire f_s_dadda_rca24_fa74_y3;
  wire f_s_dadda_rca24_fa74_y4;
  wire f_s_dadda_rca24_and_11_5_a_11;
  wire f_s_dadda_rca24_and_11_5_b_5;
  wire f_s_dadda_rca24_and_11_5_y0;
  wire f_s_dadda_rca24_and_10_6_a_10;
  wire f_s_dadda_rca24_and_10_6_b_6;
  wire f_s_dadda_rca24_and_10_6_y0;
  wire f_s_dadda_rca24_and_9_7_a_9;
  wire f_s_dadda_rca24_and_9_7_b_7;
  wire f_s_dadda_rca24_and_9_7_y0;
  wire f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_11_5_y0;
  wire f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_10_6_y0;
  wire f_s_dadda_rca24_fa75_y0;
  wire f_s_dadda_rca24_fa75_y1;
  wire f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_9_7_y0;
  wire f_s_dadda_rca24_fa75_y2;
  wire f_s_dadda_rca24_fa75_y3;
  wire f_s_dadda_rca24_fa75_y4;
  wire f_s_dadda_rca24_and_8_8_a_8;
  wire f_s_dadda_rca24_and_8_8_b_8;
  wire f_s_dadda_rca24_and_8_8_y0;
  wire f_s_dadda_rca24_and_7_9_a_7;
  wire f_s_dadda_rca24_and_7_9_b_9;
  wire f_s_dadda_rca24_and_7_9_y0;
  wire f_s_dadda_rca24_and_6_10_a_6;
  wire f_s_dadda_rca24_and_6_10_b_10;
  wire f_s_dadda_rca24_and_6_10_y0;
  wire f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_8_8_y0;
  wire f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_7_9_y0;
  wire f_s_dadda_rca24_fa76_y0;
  wire f_s_dadda_rca24_fa76_y1;
  wire f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_6_10_y0;
  wire f_s_dadda_rca24_fa76_y2;
  wire f_s_dadda_rca24_fa76_y3;
  wire f_s_dadda_rca24_fa76_y4;
  wire f_s_dadda_rca24_and_5_11_a_5;
  wire f_s_dadda_rca24_and_5_11_b_11;
  wire f_s_dadda_rca24_and_5_11_y0;
  wire f_s_dadda_rca24_and_4_12_a_4;
  wire f_s_dadda_rca24_and_4_12_b_12;
  wire f_s_dadda_rca24_and_4_12_y0;
  wire f_s_dadda_rca24_and_3_13_a_3;
  wire f_s_dadda_rca24_and_3_13_b_13;
  wire f_s_dadda_rca24_and_3_13_y0;
  wire f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_5_11_y0;
  wire f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_4_12_y0;
  wire f_s_dadda_rca24_fa77_y0;
  wire f_s_dadda_rca24_fa77_y1;
  wire f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_3_13_y0;
  wire f_s_dadda_rca24_fa77_y2;
  wire f_s_dadda_rca24_fa77_y3;
  wire f_s_dadda_rca24_fa77_y4;
  wire f_s_dadda_rca24_and_2_14_a_2;
  wire f_s_dadda_rca24_and_2_14_b_14;
  wire f_s_dadda_rca24_and_2_14_y0;
  wire f_s_dadda_rca24_and_1_15_a_1;
  wire f_s_dadda_rca24_and_1_15_b_15;
  wire f_s_dadda_rca24_and_1_15_y0;
  wire f_s_dadda_rca24_and_0_16_a_0;
  wire f_s_dadda_rca24_and_0_16_b_16;
  wire f_s_dadda_rca24_and_0_16_y0;
  wire f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_2_14_y0;
  wire f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_1_15_y0;
  wire f_s_dadda_rca24_fa78_y0;
  wire f_s_dadda_rca24_fa78_y1;
  wire f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_0_16_y0;
  wire f_s_dadda_rca24_fa78_y2;
  wire f_s_dadda_rca24_fa78_y3;
  wire f_s_dadda_rca24_fa78_y4;
  wire f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa70_y2;
  wire f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa71_y2;
  wire f_s_dadda_rca24_fa79_y0;
  wire f_s_dadda_rca24_fa79_y1;
  wire f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa72_y2;
  wire f_s_dadda_rca24_fa79_y2;
  wire f_s_dadda_rca24_fa79_y3;
  wire f_s_dadda_rca24_fa79_y4;
  wire f_s_dadda_rca24_ha15_f_s_dadda_rca24_fa73_y2;
  wire f_s_dadda_rca24_ha15_f_s_dadda_rca24_fa74_y2;
  wire f_s_dadda_rca24_ha15_y0;
  wire f_s_dadda_rca24_ha15_y1;
  wire f_s_dadda_rca24_fa80_f_s_dadda_rca24_ha15_y1;
  wire f_s_dadda_rca24_fa80_f_s_dadda_rca24_fa79_y4;
  wire f_s_dadda_rca24_fa80_y0;
  wire f_s_dadda_rca24_fa80_y1;
  wire f_s_dadda_rca24_fa80_f_s_dadda_rca24_fa78_y4;
  wire f_s_dadda_rca24_fa80_y2;
  wire f_s_dadda_rca24_fa80_y3;
  wire f_s_dadda_rca24_fa80_y4;
  wire f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa77_y4;
  wire f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa76_y4;
  wire f_s_dadda_rca24_fa81_y0;
  wire f_s_dadda_rca24_fa81_y1;
  wire f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa75_y4;
  wire f_s_dadda_rca24_fa81_y2;
  wire f_s_dadda_rca24_fa81_y3;
  wire f_s_dadda_rca24_fa81_y4;
  wire f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa74_y4;
  wire f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa73_y4;
  wire f_s_dadda_rca24_fa82_y0;
  wire f_s_dadda_rca24_fa82_y1;
  wire f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa72_y4;
  wire f_s_dadda_rca24_fa82_y2;
  wire f_s_dadda_rca24_fa82_y3;
  wire f_s_dadda_rca24_fa82_y4;
  wire f_s_dadda_rca24_and_17_0_a_17;
  wire f_s_dadda_rca24_and_17_0_b_0;
  wire f_s_dadda_rca24_and_17_0_y0;
  wire f_s_dadda_rca24_fa83_f_s_dadda_rca24_fa71_y4;
  wire f_s_dadda_rca24_fa83_f_s_dadda_rca24_fa70_y4;
  wire f_s_dadda_rca24_fa83_y0;
  wire f_s_dadda_rca24_fa83_y1;
  wire f_s_dadda_rca24_fa83_f_s_dadda_rca24_and_17_0_y0;
  wire f_s_dadda_rca24_fa83_y2;
  wire f_s_dadda_rca24_fa83_y3;
  wire f_s_dadda_rca24_fa83_y4;
  wire f_s_dadda_rca24_and_16_1_a_16;
  wire f_s_dadda_rca24_and_16_1_b_1;
  wire f_s_dadda_rca24_and_16_1_y0;
  wire f_s_dadda_rca24_and_15_2_a_15;
  wire f_s_dadda_rca24_and_15_2_b_2;
  wire f_s_dadda_rca24_and_15_2_y0;
  wire f_s_dadda_rca24_and_14_3_a_14;
  wire f_s_dadda_rca24_and_14_3_b_3;
  wire f_s_dadda_rca24_and_14_3_y0;
  wire f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_16_1_y0;
  wire f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_15_2_y0;
  wire f_s_dadda_rca24_fa84_y0;
  wire f_s_dadda_rca24_fa84_y1;
  wire f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_14_3_y0;
  wire f_s_dadda_rca24_fa84_y2;
  wire f_s_dadda_rca24_fa84_y3;
  wire f_s_dadda_rca24_fa84_y4;
  wire f_s_dadda_rca24_and_13_4_a_13;
  wire f_s_dadda_rca24_and_13_4_b_4;
  wire f_s_dadda_rca24_and_13_4_y0;
  wire f_s_dadda_rca24_and_12_5_a_12;
  wire f_s_dadda_rca24_and_12_5_b_5;
  wire f_s_dadda_rca24_and_12_5_y0;
  wire f_s_dadda_rca24_and_11_6_a_11;
  wire f_s_dadda_rca24_and_11_6_b_6;
  wire f_s_dadda_rca24_and_11_6_y0;
  wire f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_13_4_y0;
  wire f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_12_5_y0;
  wire f_s_dadda_rca24_fa85_y0;
  wire f_s_dadda_rca24_fa85_y1;
  wire f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_11_6_y0;
  wire f_s_dadda_rca24_fa85_y2;
  wire f_s_dadda_rca24_fa85_y3;
  wire f_s_dadda_rca24_fa85_y4;
  wire f_s_dadda_rca24_and_10_7_a_10;
  wire f_s_dadda_rca24_and_10_7_b_7;
  wire f_s_dadda_rca24_and_10_7_y0;
  wire f_s_dadda_rca24_and_9_8_a_9;
  wire f_s_dadda_rca24_and_9_8_b_8;
  wire f_s_dadda_rca24_and_9_8_y0;
  wire f_s_dadda_rca24_and_8_9_a_8;
  wire f_s_dadda_rca24_and_8_9_b_9;
  wire f_s_dadda_rca24_and_8_9_y0;
  wire f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_10_7_y0;
  wire f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_9_8_y0;
  wire f_s_dadda_rca24_fa86_y0;
  wire f_s_dadda_rca24_fa86_y1;
  wire f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_8_9_y0;
  wire f_s_dadda_rca24_fa86_y2;
  wire f_s_dadda_rca24_fa86_y3;
  wire f_s_dadda_rca24_fa86_y4;
  wire f_s_dadda_rca24_and_7_10_a_7;
  wire f_s_dadda_rca24_and_7_10_b_10;
  wire f_s_dadda_rca24_and_7_10_y0;
  wire f_s_dadda_rca24_and_6_11_a_6;
  wire f_s_dadda_rca24_and_6_11_b_11;
  wire f_s_dadda_rca24_and_6_11_y0;
  wire f_s_dadda_rca24_and_5_12_a_5;
  wire f_s_dadda_rca24_and_5_12_b_12;
  wire f_s_dadda_rca24_and_5_12_y0;
  wire f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_7_10_y0;
  wire f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_6_11_y0;
  wire f_s_dadda_rca24_fa87_y0;
  wire f_s_dadda_rca24_fa87_y1;
  wire f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_5_12_y0;
  wire f_s_dadda_rca24_fa87_y2;
  wire f_s_dadda_rca24_fa87_y3;
  wire f_s_dadda_rca24_fa87_y4;
  wire f_s_dadda_rca24_and_4_13_a_4;
  wire f_s_dadda_rca24_and_4_13_b_13;
  wire f_s_dadda_rca24_and_4_13_y0;
  wire f_s_dadda_rca24_and_3_14_a_3;
  wire f_s_dadda_rca24_and_3_14_b_14;
  wire f_s_dadda_rca24_and_3_14_y0;
  wire f_s_dadda_rca24_and_2_15_a_2;
  wire f_s_dadda_rca24_and_2_15_b_15;
  wire f_s_dadda_rca24_and_2_15_y0;
  wire f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_4_13_y0;
  wire f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_3_14_y0;
  wire f_s_dadda_rca24_fa88_y0;
  wire f_s_dadda_rca24_fa88_y1;
  wire f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_2_15_y0;
  wire f_s_dadda_rca24_fa88_y2;
  wire f_s_dadda_rca24_fa88_y3;
  wire f_s_dadda_rca24_fa88_y4;
  wire f_s_dadda_rca24_and_1_16_a_1;
  wire f_s_dadda_rca24_and_1_16_b_16;
  wire f_s_dadda_rca24_and_1_16_y0;
  wire f_s_dadda_rca24_and_0_17_a_0;
  wire f_s_dadda_rca24_and_0_17_b_17;
  wire f_s_dadda_rca24_and_0_17_y0;
  wire f_s_dadda_rca24_fa89_f_s_dadda_rca24_and_1_16_y0;
  wire f_s_dadda_rca24_fa89_f_s_dadda_rca24_and_0_17_y0;
  wire f_s_dadda_rca24_fa89_y0;
  wire f_s_dadda_rca24_fa89_y1;
  wire f_s_dadda_rca24_fa89_f_s_dadda_rca24_fa80_y2;
  wire f_s_dadda_rca24_fa89_y2;
  wire f_s_dadda_rca24_fa89_y3;
  wire f_s_dadda_rca24_fa89_y4;
  wire f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa81_y2;
  wire f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa82_y2;
  wire f_s_dadda_rca24_fa90_y0;
  wire f_s_dadda_rca24_fa90_y1;
  wire f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa83_y2;
  wire f_s_dadda_rca24_fa90_y2;
  wire f_s_dadda_rca24_fa90_y3;
  wire f_s_dadda_rca24_fa90_y4;
  wire f_s_dadda_rca24_ha16_f_s_dadda_rca24_fa84_y2;
  wire f_s_dadda_rca24_ha16_f_s_dadda_rca24_fa85_y2;
  wire f_s_dadda_rca24_ha16_y0;
  wire f_s_dadda_rca24_ha16_y1;
  wire f_s_dadda_rca24_fa91_f_s_dadda_rca24_ha16_y1;
  wire f_s_dadda_rca24_fa91_f_s_dadda_rca24_fa90_y4;
  wire f_s_dadda_rca24_fa91_y0;
  wire f_s_dadda_rca24_fa91_y1;
  wire f_s_dadda_rca24_fa91_f_s_dadda_rca24_fa89_y4;
  wire f_s_dadda_rca24_fa91_y2;
  wire f_s_dadda_rca24_fa91_y3;
  wire f_s_dadda_rca24_fa91_y4;
  wire f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa88_y4;
  wire f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa87_y4;
  wire f_s_dadda_rca24_fa92_y0;
  wire f_s_dadda_rca24_fa92_y1;
  wire f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa86_y4;
  wire f_s_dadda_rca24_fa92_y2;
  wire f_s_dadda_rca24_fa92_y3;
  wire f_s_dadda_rca24_fa92_y4;
  wire f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa85_y4;
  wire f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa84_y4;
  wire f_s_dadda_rca24_fa93_y0;
  wire f_s_dadda_rca24_fa93_y1;
  wire f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa83_y4;
  wire f_s_dadda_rca24_fa93_y2;
  wire f_s_dadda_rca24_fa93_y3;
  wire f_s_dadda_rca24_fa93_y4;
  wire f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa82_y4;
  wire f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa81_y4;
  wire f_s_dadda_rca24_fa94_y0;
  wire f_s_dadda_rca24_fa94_y1;
  wire f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa80_y4;
  wire f_s_dadda_rca24_fa94_y2;
  wire f_s_dadda_rca24_fa94_y3;
  wire f_s_dadda_rca24_fa94_y4;
  wire f_s_dadda_rca24_and_18_0_a_18;
  wire f_s_dadda_rca24_and_18_0_b_0;
  wire f_s_dadda_rca24_and_18_0_y0;
  wire f_s_dadda_rca24_and_17_1_a_17;
  wire f_s_dadda_rca24_and_17_1_b_1;
  wire f_s_dadda_rca24_and_17_1_y0;
  wire f_s_dadda_rca24_and_16_2_a_16;
  wire f_s_dadda_rca24_and_16_2_b_2;
  wire f_s_dadda_rca24_and_16_2_y0;
  wire f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_18_0_y0;
  wire f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_17_1_y0;
  wire f_s_dadda_rca24_fa95_y0;
  wire f_s_dadda_rca24_fa95_y1;
  wire f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_16_2_y0;
  wire f_s_dadda_rca24_fa95_y2;
  wire f_s_dadda_rca24_fa95_y3;
  wire f_s_dadda_rca24_fa95_y4;
  wire f_s_dadda_rca24_and_15_3_a_15;
  wire f_s_dadda_rca24_and_15_3_b_3;
  wire f_s_dadda_rca24_and_15_3_y0;
  wire f_s_dadda_rca24_and_14_4_a_14;
  wire f_s_dadda_rca24_and_14_4_b_4;
  wire f_s_dadda_rca24_and_14_4_y0;
  wire f_s_dadda_rca24_and_13_5_a_13;
  wire f_s_dadda_rca24_and_13_5_b_5;
  wire f_s_dadda_rca24_and_13_5_y0;
  wire f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_15_3_y0;
  wire f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_14_4_y0;
  wire f_s_dadda_rca24_fa96_y0;
  wire f_s_dadda_rca24_fa96_y1;
  wire f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_13_5_y0;
  wire f_s_dadda_rca24_fa96_y2;
  wire f_s_dadda_rca24_fa96_y3;
  wire f_s_dadda_rca24_fa96_y4;
  wire f_s_dadda_rca24_and_12_6_a_12;
  wire f_s_dadda_rca24_and_12_6_b_6;
  wire f_s_dadda_rca24_and_12_6_y0;
  wire f_s_dadda_rca24_and_11_7_a_11;
  wire f_s_dadda_rca24_and_11_7_b_7;
  wire f_s_dadda_rca24_and_11_7_y0;
  wire f_s_dadda_rca24_and_10_8_a_10;
  wire f_s_dadda_rca24_and_10_8_b_8;
  wire f_s_dadda_rca24_and_10_8_y0;
  wire f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_12_6_y0;
  wire f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_11_7_y0;
  wire f_s_dadda_rca24_fa97_y0;
  wire f_s_dadda_rca24_fa97_y1;
  wire f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_10_8_y0;
  wire f_s_dadda_rca24_fa97_y2;
  wire f_s_dadda_rca24_fa97_y3;
  wire f_s_dadda_rca24_fa97_y4;
  wire f_s_dadda_rca24_and_9_9_a_9;
  wire f_s_dadda_rca24_and_9_9_b_9;
  wire f_s_dadda_rca24_and_9_9_y0;
  wire f_s_dadda_rca24_and_8_10_a_8;
  wire f_s_dadda_rca24_and_8_10_b_10;
  wire f_s_dadda_rca24_and_8_10_y0;
  wire f_s_dadda_rca24_and_7_11_a_7;
  wire f_s_dadda_rca24_and_7_11_b_11;
  wire f_s_dadda_rca24_and_7_11_y0;
  wire f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_9_9_y0;
  wire f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_8_10_y0;
  wire f_s_dadda_rca24_fa98_y0;
  wire f_s_dadda_rca24_fa98_y1;
  wire f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_7_11_y0;
  wire f_s_dadda_rca24_fa98_y2;
  wire f_s_dadda_rca24_fa98_y3;
  wire f_s_dadda_rca24_fa98_y4;
  wire f_s_dadda_rca24_and_6_12_a_6;
  wire f_s_dadda_rca24_and_6_12_b_12;
  wire f_s_dadda_rca24_and_6_12_y0;
  wire f_s_dadda_rca24_and_5_13_a_5;
  wire f_s_dadda_rca24_and_5_13_b_13;
  wire f_s_dadda_rca24_and_5_13_y0;
  wire f_s_dadda_rca24_and_4_14_a_4;
  wire f_s_dadda_rca24_and_4_14_b_14;
  wire f_s_dadda_rca24_and_4_14_y0;
  wire f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_6_12_y0;
  wire f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_5_13_y0;
  wire f_s_dadda_rca24_fa99_y0;
  wire f_s_dadda_rca24_fa99_y1;
  wire f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_4_14_y0;
  wire f_s_dadda_rca24_fa99_y2;
  wire f_s_dadda_rca24_fa99_y3;
  wire f_s_dadda_rca24_fa99_y4;
  wire f_s_dadda_rca24_and_3_15_a_3;
  wire f_s_dadda_rca24_and_3_15_b_15;
  wire f_s_dadda_rca24_and_3_15_y0;
  wire f_s_dadda_rca24_and_2_16_a_2;
  wire f_s_dadda_rca24_and_2_16_b_16;
  wire f_s_dadda_rca24_and_2_16_y0;
  wire f_s_dadda_rca24_and_1_17_a_1;
  wire f_s_dadda_rca24_and_1_17_b_17;
  wire f_s_dadda_rca24_and_1_17_y0;
  wire f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_3_15_y0;
  wire f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_2_16_y0;
  wire f_s_dadda_rca24_fa100_y0;
  wire f_s_dadda_rca24_fa100_y1;
  wire f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_1_17_y0;
  wire f_s_dadda_rca24_fa100_y2;
  wire f_s_dadda_rca24_fa100_y3;
  wire f_s_dadda_rca24_fa100_y4;
  wire f_s_dadda_rca24_and_0_18_a_0;
  wire f_s_dadda_rca24_and_0_18_b_18;
  wire f_s_dadda_rca24_and_0_18_y0;
  wire f_s_dadda_rca24_fa101_f_s_dadda_rca24_and_0_18_y0;
  wire f_s_dadda_rca24_fa101_f_s_dadda_rca24_fa91_y2;
  wire f_s_dadda_rca24_fa101_y0;
  wire f_s_dadda_rca24_fa101_y1;
  wire f_s_dadda_rca24_fa101_f_s_dadda_rca24_fa92_y2;
  wire f_s_dadda_rca24_fa101_y2;
  wire f_s_dadda_rca24_fa101_y3;
  wire f_s_dadda_rca24_fa101_y4;
  wire f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa93_y2;
  wire f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa94_y2;
  wire f_s_dadda_rca24_fa102_y0;
  wire f_s_dadda_rca24_fa102_y1;
  wire f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa95_y2;
  wire f_s_dadda_rca24_fa102_y2;
  wire f_s_dadda_rca24_fa102_y3;
  wire f_s_dadda_rca24_fa102_y4;
  wire f_s_dadda_rca24_ha17_f_s_dadda_rca24_fa96_y2;
  wire f_s_dadda_rca24_ha17_f_s_dadda_rca24_fa97_y2;
  wire f_s_dadda_rca24_ha17_y0;
  wire f_s_dadda_rca24_ha17_y1;
  wire f_s_dadda_rca24_fa103_f_s_dadda_rca24_ha17_y1;
  wire f_s_dadda_rca24_fa103_f_s_dadda_rca24_fa102_y4;
  wire f_s_dadda_rca24_fa103_y0;
  wire f_s_dadda_rca24_fa103_y1;
  wire f_s_dadda_rca24_fa103_f_s_dadda_rca24_fa101_y4;
  wire f_s_dadda_rca24_fa103_y2;
  wire f_s_dadda_rca24_fa103_y3;
  wire f_s_dadda_rca24_fa103_y4;
  wire f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa100_y4;
  wire f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa99_y4;
  wire f_s_dadda_rca24_fa104_y0;
  wire f_s_dadda_rca24_fa104_y1;
  wire f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa98_y4;
  wire f_s_dadda_rca24_fa104_y2;
  wire f_s_dadda_rca24_fa104_y3;
  wire f_s_dadda_rca24_fa104_y4;
  wire f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa97_y4;
  wire f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa96_y4;
  wire f_s_dadda_rca24_fa105_y0;
  wire f_s_dadda_rca24_fa105_y1;
  wire f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa95_y4;
  wire f_s_dadda_rca24_fa105_y2;
  wire f_s_dadda_rca24_fa105_y3;
  wire f_s_dadda_rca24_fa105_y4;
  wire f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa94_y4;
  wire f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa93_y4;
  wire f_s_dadda_rca24_fa106_y0;
  wire f_s_dadda_rca24_fa106_y1;
  wire f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa92_y4;
  wire f_s_dadda_rca24_fa106_y2;
  wire f_s_dadda_rca24_fa106_y3;
  wire f_s_dadda_rca24_fa106_y4;
  wire f_s_dadda_rca24_and_17_2_a_17;
  wire f_s_dadda_rca24_and_17_2_b_2;
  wire f_s_dadda_rca24_and_17_2_y0;
  wire f_s_dadda_rca24_and_16_3_a_16;
  wire f_s_dadda_rca24_and_16_3_b_3;
  wire f_s_dadda_rca24_and_16_3_y0;
  wire f_s_dadda_rca24_fa107_f_s_dadda_rca24_fa91_y4;
  wire f_s_dadda_rca24_fa107_f_s_dadda_rca24_and_17_2_y0;
  wire f_s_dadda_rca24_fa107_y0;
  wire f_s_dadda_rca24_fa107_y1;
  wire f_s_dadda_rca24_fa107_f_s_dadda_rca24_and_16_3_y0;
  wire f_s_dadda_rca24_fa107_y2;
  wire f_s_dadda_rca24_fa107_y3;
  wire f_s_dadda_rca24_fa107_y4;
  wire f_s_dadda_rca24_and_15_4_a_15;
  wire f_s_dadda_rca24_and_15_4_b_4;
  wire f_s_dadda_rca24_and_15_4_y0;
  wire f_s_dadda_rca24_and_14_5_a_14;
  wire f_s_dadda_rca24_and_14_5_b_5;
  wire f_s_dadda_rca24_and_14_5_y0;
  wire f_s_dadda_rca24_and_13_6_a_13;
  wire f_s_dadda_rca24_and_13_6_b_6;
  wire f_s_dadda_rca24_and_13_6_y0;
  wire f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_15_4_y0;
  wire f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_14_5_y0;
  wire f_s_dadda_rca24_fa108_y0;
  wire f_s_dadda_rca24_fa108_y1;
  wire f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_13_6_y0;
  wire f_s_dadda_rca24_fa108_y2;
  wire f_s_dadda_rca24_fa108_y3;
  wire f_s_dadda_rca24_fa108_y4;
  wire f_s_dadda_rca24_and_12_7_a_12;
  wire f_s_dadda_rca24_and_12_7_b_7;
  wire f_s_dadda_rca24_and_12_7_y0;
  wire f_s_dadda_rca24_and_11_8_a_11;
  wire f_s_dadda_rca24_and_11_8_b_8;
  wire f_s_dadda_rca24_and_11_8_y0;
  wire f_s_dadda_rca24_and_10_9_a_10;
  wire f_s_dadda_rca24_and_10_9_b_9;
  wire f_s_dadda_rca24_and_10_9_y0;
  wire f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_12_7_y0;
  wire f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_11_8_y0;
  wire f_s_dadda_rca24_fa109_y0;
  wire f_s_dadda_rca24_fa109_y1;
  wire f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_10_9_y0;
  wire f_s_dadda_rca24_fa109_y2;
  wire f_s_dadda_rca24_fa109_y3;
  wire f_s_dadda_rca24_fa109_y4;
  wire f_s_dadda_rca24_and_9_10_a_9;
  wire f_s_dadda_rca24_and_9_10_b_10;
  wire f_s_dadda_rca24_and_9_10_y0;
  wire f_s_dadda_rca24_and_8_11_a_8;
  wire f_s_dadda_rca24_and_8_11_b_11;
  wire f_s_dadda_rca24_and_8_11_y0;
  wire f_s_dadda_rca24_and_7_12_a_7;
  wire f_s_dadda_rca24_and_7_12_b_12;
  wire f_s_dadda_rca24_and_7_12_y0;
  wire f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_9_10_y0;
  wire f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_8_11_y0;
  wire f_s_dadda_rca24_fa110_y0;
  wire f_s_dadda_rca24_fa110_y1;
  wire f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_7_12_y0;
  wire f_s_dadda_rca24_fa110_y2;
  wire f_s_dadda_rca24_fa110_y3;
  wire f_s_dadda_rca24_fa110_y4;
  wire f_s_dadda_rca24_and_6_13_a_6;
  wire f_s_dadda_rca24_and_6_13_b_13;
  wire f_s_dadda_rca24_and_6_13_y0;
  wire f_s_dadda_rca24_and_5_14_a_5;
  wire f_s_dadda_rca24_and_5_14_b_14;
  wire f_s_dadda_rca24_and_5_14_y0;
  wire f_s_dadda_rca24_and_4_15_a_4;
  wire f_s_dadda_rca24_and_4_15_b_15;
  wire f_s_dadda_rca24_and_4_15_y0;
  wire f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_6_13_y0;
  wire f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_5_14_y0;
  wire f_s_dadda_rca24_fa111_y0;
  wire f_s_dadda_rca24_fa111_y1;
  wire f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_4_15_y0;
  wire f_s_dadda_rca24_fa111_y2;
  wire f_s_dadda_rca24_fa111_y3;
  wire f_s_dadda_rca24_fa111_y4;
  wire f_s_dadda_rca24_and_3_16_a_3;
  wire f_s_dadda_rca24_and_3_16_b_16;
  wire f_s_dadda_rca24_and_3_16_y0;
  wire f_s_dadda_rca24_and_2_17_a_2;
  wire f_s_dadda_rca24_and_2_17_b_17;
  wire f_s_dadda_rca24_and_2_17_y0;
  wire f_s_dadda_rca24_and_1_18_a_1;
  wire f_s_dadda_rca24_and_1_18_b_18;
  wire f_s_dadda_rca24_and_1_18_y0;
  wire f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_3_16_y0;
  wire f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_2_17_y0;
  wire f_s_dadda_rca24_fa112_y0;
  wire f_s_dadda_rca24_fa112_y1;
  wire f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_1_18_y0;
  wire f_s_dadda_rca24_fa112_y2;
  wire f_s_dadda_rca24_fa112_y3;
  wire f_s_dadda_rca24_fa112_y4;
  wire f_s_dadda_rca24_and_0_19_a_0;
  wire f_s_dadda_rca24_and_0_19_b_19;
  wire f_s_dadda_rca24_and_0_19_y0;
  wire f_s_dadda_rca24_fa113_f_s_dadda_rca24_and_0_19_y0;
  wire f_s_dadda_rca24_fa113_f_s_dadda_rca24_ha0_y0;
  wire f_s_dadda_rca24_fa113_y0;
  wire f_s_dadda_rca24_fa113_y1;
  wire f_s_dadda_rca24_fa113_f_s_dadda_rca24_fa103_y2;
  wire f_s_dadda_rca24_fa113_y2;
  wire f_s_dadda_rca24_fa113_y3;
  wire f_s_dadda_rca24_fa113_y4;
  wire f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa104_y2;
  wire f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa105_y2;
  wire f_s_dadda_rca24_fa114_y0;
  wire f_s_dadda_rca24_fa114_y1;
  wire f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa106_y2;
  wire f_s_dadda_rca24_fa114_y2;
  wire f_s_dadda_rca24_fa114_y3;
  wire f_s_dadda_rca24_fa114_y4;
  wire f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa107_y2;
  wire f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa108_y2;
  wire f_s_dadda_rca24_fa115_y0;
  wire f_s_dadda_rca24_fa115_y1;
  wire f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa109_y2;
  wire f_s_dadda_rca24_fa115_y2;
  wire f_s_dadda_rca24_fa115_y3;
  wire f_s_dadda_rca24_fa115_y4;
  wire f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa115_y4;
  wire f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa114_y4;
  wire f_s_dadda_rca24_fa116_y0;
  wire f_s_dadda_rca24_fa116_y1;
  wire f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa113_y4;
  wire f_s_dadda_rca24_fa116_y2;
  wire f_s_dadda_rca24_fa116_y3;
  wire f_s_dadda_rca24_fa116_y4;
  wire f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa112_y4;
  wire f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa111_y4;
  wire f_s_dadda_rca24_fa117_y0;
  wire f_s_dadda_rca24_fa117_y1;
  wire f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa110_y4;
  wire f_s_dadda_rca24_fa117_y2;
  wire f_s_dadda_rca24_fa117_y3;
  wire f_s_dadda_rca24_fa117_y4;
  wire f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa109_y4;
  wire f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa108_y4;
  wire f_s_dadda_rca24_fa118_y0;
  wire f_s_dadda_rca24_fa118_y1;
  wire f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa107_y4;
  wire f_s_dadda_rca24_fa118_y2;
  wire f_s_dadda_rca24_fa118_y3;
  wire f_s_dadda_rca24_fa118_y4;
  wire f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa106_y4;
  wire f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa105_y4;
  wire f_s_dadda_rca24_fa119_y0;
  wire f_s_dadda_rca24_fa119_y1;
  wire f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa104_y4;
  wire f_s_dadda_rca24_fa119_y2;
  wire f_s_dadda_rca24_fa119_y3;
  wire f_s_dadda_rca24_fa119_y4;
  wire f_s_dadda_rca24_and_16_4_a_16;
  wire f_s_dadda_rca24_and_16_4_b_4;
  wire f_s_dadda_rca24_and_16_4_y0;
  wire f_s_dadda_rca24_and_15_5_a_15;
  wire f_s_dadda_rca24_and_15_5_b_5;
  wire f_s_dadda_rca24_and_15_5_y0;
  wire f_s_dadda_rca24_fa120_f_s_dadda_rca24_fa103_y4;
  wire f_s_dadda_rca24_fa120_f_s_dadda_rca24_and_16_4_y0;
  wire f_s_dadda_rca24_fa120_y0;
  wire f_s_dadda_rca24_fa120_y1;
  wire f_s_dadda_rca24_fa120_f_s_dadda_rca24_and_15_5_y0;
  wire f_s_dadda_rca24_fa120_y2;
  wire f_s_dadda_rca24_fa120_y3;
  wire f_s_dadda_rca24_fa120_y4;
  wire f_s_dadda_rca24_and_14_6_a_14;
  wire f_s_dadda_rca24_and_14_6_b_6;
  wire f_s_dadda_rca24_and_14_6_y0;
  wire f_s_dadda_rca24_and_13_7_a_13;
  wire f_s_dadda_rca24_and_13_7_b_7;
  wire f_s_dadda_rca24_and_13_7_y0;
  wire f_s_dadda_rca24_and_12_8_a_12;
  wire f_s_dadda_rca24_and_12_8_b_8;
  wire f_s_dadda_rca24_and_12_8_y0;
  wire f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_14_6_y0;
  wire f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_13_7_y0;
  wire f_s_dadda_rca24_fa121_y0;
  wire f_s_dadda_rca24_fa121_y1;
  wire f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_12_8_y0;
  wire f_s_dadda_rca24_fa121_y2;
  wire f_s_dadda_rca24_fa121_y3;
  wire f_s_dadda_rca24_fa121_y4;
  wire f_s_dadda_rca24_and_11_9_a_11;
  wire f_s_dadda_rca24_and_11_9_b_9;
  wire f_s_dadda_rca24_and_11_9_y0;
  wire f_s_dadda_rca24_and_10_10_a_10;
  wire f_s_dadda_rca24_and_10_10_b_10;
  wire f_s_dadda_rca24_and_10_10_y0;
  wire f_s_dadda_rca24_and_9_11_a_9;
  wire f_s_dadda_rca24_and_9_11_b_11;
  wire f_s_dadda_rca24_and_9_11_y0;
  wire f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_11_9_y0;
  wire f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_10_10_y0;
  wire f_s_dadda_rca24_fa122_y0;
  wire f_s_dadda_rca24_fa122_y1;
  wire f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_9_11_y0;
  wire f_s_dadda_rca24_fa122_y2;
  wire f_s_dadda_rca24_fa122_y3;
  wire f_s_dadda_rca24_fa122_y4;
  wire f_s_dadda_rca24_and_8_12_a_8;
  wire f_s_dadda_rca24_and_8_12_b_12;
  wire f_s_dadda_rca24_and_8_12_y0;
  wire f_s_dadda_rca24_and_7_13_a_7;
  wire f_s_dadda_rca24_and_7_13_b_13;
  wire f_s_dadda_rca24_and_7_13_y0;
  wire f_s_dadda_rca24_and_6_14_a_6;
  wire f_s_dadda_rca24_and_6_14_b_14;
  wire f_s_dadda_rca24_and_6_14_y0;
  wire f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_8_12_y0;
  wire f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_7_13_y0;
  wire f_s_dadda_rca24_fa123_y0;
  wire f_s_dadda_rca24_fa123_y1;
  wire f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_6_14_y0;
  wire f_s_dadda_rca24_fa123_y2;
  wire f_s_dadda_rca24_fa123_y3;
  wire f_s_dadda_rca24_fa123_y4;
  wire f_s_dadda_rca24_and_5_15_a_5;
  wire f_s_dadda_rca24_and_5_15_b_15;
  wire f_s_dadda_rca24_and_5_15_y0;
  wire f_s_dadda_rca24_and_4_16_a_4;
  wire f_s_dadda_rca24_and_4_16_b_16;
  wire f_s_dadda_rca24_and_4_16_y0;
  wire f_s_dadda_rca24_and_3_17_a_3;
  wire f_s_dadda_rca24_and_3_17_b_17;
  wire f_s_dadda_rca24_and_3_17_y0;
  wire f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_5_15_y0;
  wire f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_4_16_y0;
  wire f_s_dadda_rca24_fa124_y0;
  wire f_s_dadda_rca24_fa124_y1;
  wire f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_3_17_y0;
  wire f_s_dadda_rca24_fa124_y2;
  wire f_s_dadda_rca24_fa124_y3;
  wire f_s_dadda_rca24_fa124_y4;
  wire f_s_dadda_rca24_and_2_18_a_2;
  wire f_s_dadda_rca24_and_2_18_b_18;
  wire f_s_dadda_rca24_and_2_18_y0;
  wire f_s_dadda_rca24_and_1_19_a_1;
  wire f_s_dadda_rca24_and_1_19_b_19;
  wire f_s_dadda_rca24_and_1_19_y0;
  wire f_s_dadda_rca24_and_0_20_a_0;
  wire f_s_dadda_rca24_and_0_20_b_20;
  wire f_s_dadda_rca24_and_0_20_y0;
  wire f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_2_18_y0;
  wire f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_1_19_y0;
  wire f_s_dadda_rca24_fa125_y0;
  wire f_s_dadda_rca24_fa125_y1;
  wire f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_0_20_y0;
  wire f_s_dadda_rca24_fa125_y2;
  wire f_s_dadda_rca24_fa125_y3;
  wire f_s_dadda_rca24_fa125_y4;
  wire f_s_dadda_rca24_fa126_f_s_dadda_rca24_fa0_y2;
  wire f_s_dadda_rca24_fa126_f_s_dadda_rca24_ha1_y0;
  wire f_s_dadda_rca24_fa126_y0;
  wire f_s_dadda_rca24_fa126_y1;
  wire f_s_dadda_rca24_fa126_f_s_dadda_rca24_fa116_y2;
  wire f_s_dadda_rca24_fa126_y2;
  wire f_s_dadda_rca24_fa126_y3;
  wire f_s_dadda_rca24_fa126_y4;
  wire f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa117_y2;
  wire f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa118_y2;
  wire f_s_dadda_rca24_fa127_y0;
  wire f_s_dadda_rca24_fa127_y1;
  wire f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa119_y2;
  wire f_s_dadda_rca24_fa127_y2;
  wire f_s_dadda_rca24_fa127_y3;
  wire f_s_dadda_rca24_fa127_y4;
  wire f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa120_y2;
  wire f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa121_y2;
  wire f_s_dadda_rca24_fa128_y0;
  wire f_s_dadda_rca24_fa128_y1;
  wire f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa122_y2;
  wire f_s_dadda_rca24_fa128_y2;
  wire f_s_dadda_rca24_fa128_y3;
  wire f_s_dadda_rca24_fa128_y4;
  wire f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa128_y4;
  wire f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa127_y4;
  wire f_s_dadda_rca24_fa129_y0;
  wire f_s_dadda_rca24_fa129_y1;
  wire f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa126_y4;
  wire f_s_dadda_rca24_fa129_y2;
  wire f_s_dadda_rca24_fa129_y3;
  wire f_s_dadda_rca24_fa129_y4;
  wire f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa125_y4;
  wire f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa124_y4;
  wire f_s_dadda_rca24_fa130_y0;
  wire f_s_dadda_rca24_fa130_y1;
  wire f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa123_y4;
  wire f_s_dadda_rca24_fa130_y2;
  wire f_s_dadda_rca24_fa130_y3;
  wire f_s_dadda_rca24_fa130_y4;
  wire f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa122_y4;
  wire f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa121_y4;
  wire f_s_dadda_rca24_fa131_y0;
  wire f_s_dadda_rca24_fa131_y1;
  wire f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa120_y4;
  wire f_s_dadda_rca24_fa131_y2;
  wire f_s_dadda_rca24_fa131_y3;
  wire f_s_dadda_rca24_fa131_y4;
  wire f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa119_y4;
  wire f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa118_y4;
  wire f_s_dadda_rca24_fa132_y0;
  wire f_s_dadda_rca24_fa132_y1;
  wire f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa117_y4;
  wire f_s_dadda_rca24_fa132_y2;
  wire f_s_dadda_rca24_fa132_y3;
  wire f_s_dadda_rca24_fa132_y4;
  wire f_s_dadda_rca24_and_15_6_a_15;
  wire f_s_dadda_rca24_and_15_6_b_6;
  wire f_s_dadda_rca24_and_15_6_y0;
  wire f_s_dadda_rca24_and_14_7_a_14;
  wire f_s_dadda_rca24_and_14_7_b_7;
  wire f_s_dadda_rca24_and_14_7_y0;
  wire f_s_dadda_rca24_fa133_f_s_dadda_rca24_fa116_y4;
  wire f_s_dadda_rca24_fa133_f_s_dadda_rca24_and_15_6_y0;
  wire f_s_dadda_rca24_fa133_y0;
  wire f_s_dadda_rca24_fa133_y1;
  wire f_s_dadda_rca24_fa133_f_s_dadda_rca24_and_14_7_y0;
  wire f_s_dadda_rca24_fa133_y2;
  wire f_s_dadda_rca24_fa133_y3;
  wire f_s_dadda_rca24_fa133_y4;
  wire f_s_dadda_rca24_and_13_8_a_13;
  wire f_s_dadda_rca24_and_13_8_b_8;
  wire f_s_dadda_rca24_and_13_8_y0;
  wire f_s_dadda_rca24_and_12_9_a_12;
  wire f_s_dadda_rca24_and_12_9_b_9;
  wire f_s_dadda_rca24_and_12_9_y0;
  wire f_s_dadda_rca24_and_11_10_a_11;
  wire f_s_dadda_rca24_and_11_10_b_10;
  wire f_s_dadda_rca24_and_11_10_y0;
  wire f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_13_8_y0;
  wire f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_12_9_y0;
  wire f_s_dadda_rca24_fa134_y0;
  wire f_s_dadda_rca24_fa134_y1;
  wire f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_11_10_y0;
  wire f_s_dadda_rca24_fa134_y2;
  wire f_s_dadda_rca24_fa134_y3;
  wire f_s_dadda_rca24_fa134_y4;
  wire f_s_dadda_rca24_and_10_11_a_10;
  wire f_s_dadda_rca24_and_10_11_b_11;
  wire f_s_dadda_rca24_and_10_11_y0;
  wire f_s_dadda_rca24_and_9_12_a_9;
  wire f_s_dadda_rca24_and_9_12_b_12;
  wire f_s_dadda_rca24_and_9_12_y0;
  wire f_s_dadda_rca24_and_8_13_a_8;
  wire f_s_dadda_rca24_and_8_13_b_13;
  wire f_s_dadda_rca24_and_8_13_y0;
  wire f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_10_11_y0;
  wire f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_9_12_y0;
  wire f_s_dadda_rca24_fa135_y0;
  wire f_s_dadda_rca24_fa135_y1;
  wire f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_8_13_y0;
  wire f_s_dadda_rca24_fa135_y2;
  wire f_s_dadda_rca24_fa135_y3;
  wire f_s_dadda_rca24_fa135_y4;
  wire f_s_dadda_rca24_and_7_14_a_7;
  wire f_s_dadda_rca24_and_7_14_b_14;
  wire f_s_dadda_rca24_and_7_14_y0;
  wire f_s_dadda_rca24_and_6_15_a_6;
  wire f_s_dadda_rca24_and_6_15_b_15;
  wire f_s_dadda_rca24_and_6_15_y0;
  wire f_s_dadda_rca24_and_5_16_a_5;
  wire f_s_dadda_rca24_and_5_16_b_16;
  wire f_s_dadda_rca24_and_5_16_y0;
  wire f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_7_14_y0;
  wire f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_6_15_y0;
  wire f_s_dadda_rca24_fa136_y0;
  wire f_s_dadda_rca24_fa136_y1;
  wire f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_5_16_y0;
  wire f_s_dadda_rca24_fa136_y2;
  wire f_s_dadda_rca24_fa136_y3;
  wire f_s_dadda_rca24_fa136_y4;
  wire f_s_dadda_rca24_and_4_17_a_4;
  wire f_s_dadda_rca24_and_4_17_b_17;
  wire f_s_dadda_rca24_and_4_17_y0;
  wire f_s_dadda_rca24_and_3_18_a_3;
  wire f_s_dadda_rca24_and_3_18_b_18;
  wire f_s_dadda_rca24_and_3_18_y0;
  wire f_s_dadda_rca24_and_2_19_a_2;
  wire f_s_dadda_rca24_and_2_19_b_19;
  wire f_s_dadda_rca24_and_2_19_y0;
  wire f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_4_17_y0;
  wire f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_3_18_y0;
  wire f_s_dadda_rca24_fa137_y0;
  wire f_s_dadda_rca24_fa137_y1;
  wire f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_2_19_y0;
  wire f_s_dadda_rca24_fa137_y2;
  wire f_s_dadda_rca24_fa137_y3;
  wire f_s_dadda_rca24_fa137_y4;
  wire f_s_dadda_rca24_and_1_20_a_1;
  wire f_s_dadda_rca24_and_1_20_b_20;
  wire f_s_dadda_rca24_and_1_20_y0;
  wire f_s_dadda_rca24_and_0_21_a_0;
  wire f_s_dadda_rca24_and_0_21_b_21;
  wire f_s_dadda_rca24_and_0_21_y0;
  wire f_s_dadda_rca24_fa138_f_s_dadda_rca24_and_1_20_y0;
  wire f_s_dadda_rca24_fa138_f_s_dadda_rca24_and_0_21_y0;
  wire f_s_dadda_rca24_fa138_y0;
  wire f_s_dadda_rca24_fa138_y1;
  wire f_s_dadda_rca24_fa138_f_s_dadda_rca24_fa1_y2;
  wire f_s_dadda_rca24_fa138_y2;
  wire f_s_dadda_rca24_fa138_y3;
  wire f_s_dadda_rca24_fa138_y4;
  wire f_s_dadda_rca24_fa139_f_s_dadda_rca24_fa2_y2;
  wire f_s_dadda_rca24_fa139_f_s_dadda_rca24_ha2_y0;
  wire f_s_dadda_rca24_fa139_y0;
  wire f_s_dadda_rca24_fa139_y1;
  wire f_s_dadda_rca24_fa139_f_s_dadda_rca24_fa129_y2;
  wire f_s_dadda_rca24_fa139_y2;
  wire f_s_dadda_rca24_fa139_y3;
  wire f_s_dadda_rca24_fa139_y4;
  wire f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa130_y2;
  wire f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa131_y2;
  wire f_s_dadda_rca24_fa140_y0;
  wire f_s_dadda_rca24_fa140_y1;
  wire f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa132_y2;
  wire f_s_dadda_rca24_fa140_y2;
  wire f_s_dadda_rca24_fa140_y3;
  wire f_s_dadda_rca24_fa140_y4;
  wire f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa133_y2;
  wire f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa134_y2;
  wire f_s_dadda_rca24_fa141_y0;
  wire f_s_dadda_rca24_fa141_y1;
  wire f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa135_y2;
  wire f_s_dadda_rca24_fa141_y2;
  wire f_s_dadda_rca24_fa141_y3;
  wire f_s_dadda_rca24_fa141_y4;
  wire f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa141_y4;
  wire f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa140_y4;
  wire f_s_dadda_rca24_fa142_y0;
  wire f_s_dadda_rca24_fa142_y1;
  wire f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa139_y4;
  wire f_s_dadda_rca24_fa142_y2;
  wire f_s_dadda_rca24_fa142_y3;
  wire f_s_dadda_rca24_fa142_y4;
  wire f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa138_y4;
  wire f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa137_y4;
  wire f_s_dadda_rca24_fa143_y0;
  wire f_s_dadda_rca24_fa143_y1;
  wire f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa136_y4;
  wire f_s_dadda_rca24_fa143_y2;
  wire f_s_dadda_rca24_fa143_y3;
  wire f_s_dadda_rca24_fa143_y4;
  wire f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa135_y4;
  wire f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa134_y4;
  wire f_s_dadda_rca24_fa144_y0;
  wire f_s_dadda_rca24_fa144_y1;
  wire f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa133_y4;
  wire f_s_dadda_rca24_fa144_y2;
  wire f_s_dadda_rca24_fa144_y3;
  wire f_s_dadda_rca24_fa144_y4;
  wire f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa132_y4;
  wire f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa131_y4;
  wire f_s_dadda_rca24_fa145_y0;
  wire f_s_dadda_rca24_fa145_y1;
  wire f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa130_y4;
  wire f_s_dadda_rca24_fa145_y2;
  wire f_s_dadda_rca24_fa145_y3;
  wire f_s_dadda_rca24_fa145_y4;
  wire f_s_dadda_rca24_and_14_8_a_14;
  wire f_s_dadda_rca24_and_14_8_b_8;
  wire f_s_dadda_rca24_and_14_8_y0;
  wire f_s_dadda_rca24_and_13_9_a_13;
  wire f_s_dadda_rca24_and_13_9_b_9;
  wire f_s_dadda_rca24_and_13_9_y0;
  wire f_s_dadda_rca24_fa146_f_s_dadda_rca24_fa129_y4;
  wire f_s_dadda_rca24_fa146_f_s_dadda_rca24_and_14_8_y0;
  wire f_s_dadda_rca24_fa146_y0;
  wire f_s_dadda_rca24_fa146_y1;
  wire f_s_dadda_rca24_fa146_f_s_dadda_rca24_and_13_9_y0;
  wire f_s_dadda_rca24_fa146_y2;
  wire f_s_dadda_rca24_fa146_y3;
  wire f_s_dadda_rca24_fa146_y4;
  wire f_s_dadda_rca24_and_12_10_a_12;
  wire f_s_dadda_rca24_and_12_10_b_10;
  wire f_s_dadda_rca24_and_12_10_y0;
  wire f_s_dadda_rca24_and_11_11_a_11;
  wire f_s_dadda_rca24_and_11_11_b_11;
  wire f_s_dadda_rca24_and_11_11_y0;
  wire f_s_dadda_rca24_and_10_12_a_10;
  wire f_s_dadda_rca24_and_10_12_b_12;
  wire f_s_dadda_rca24_and_10_12_y0;
  wire f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_12_10_y0;
  wire f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_11_11_y0;
  wire f_s_dadda_rca24_fa147_y0;
  wire f_s_dadda_rca24_fa147_y1;
  wire f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_10_12_y0;
  wire f_s_dadda_rca24_fa147_y2;
  wire f_s_dadda_rca24_fa147_y3;
  wire f_s_dadda_rca24_fa147_y4;
  wire f_s_dadda_rca24_and_9_13_a_9;
  wire f_s_dadda_rca24_and_9_13_b_13;
  wire f_s_dadda_rca24_and_9_13_y0;
  wire f_s_dadda_rca24_and_8_14_a_8;
  wire f_s_dadda_rca24_and_8_14_b_14;
  wire f_s_dadda_rca24_and_8_14_y0;
  wire f_s_dadda_rca24_and_7_15_a_7;
  wire f_s_dadda_rca24_and_7_15_b_15;
  wire f_s_dadda_rca24_and_7_15_y0;
  wire f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_9_13_y0;
  wire f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_8_14_y0;
  wire f_s_dadda_rca24_fa148_y0;
  wire f_s_dadda_rca24_fa148_y1;
  wire f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_7_15_y0;
  wire f_s_dadda_rca24_fa148_y2;
  wire f_s_dadda_rca24_fa148_y3;
  wire f_s_dadda_rca24_fa148_y4;
  wire f_s_dadda_rca24_and_6_16_a_6;
  wire f_s_dadda_rca24_and_6_16_b_16;
  wire f_s_dadda_rca24_and_6_16_y0;
  wire f_s_dadda_rca24_and_5_17_a_5;
  wire f_s_dadda_rca24_and_5_17_b_17;
  wire f_s_dadda_rca24_and_5_17_y0;
  wire f_s_dadda_rca24_and_4_18_a_4;
  wire f_s_dadda_rca24_and_4_18_b_18;
  wire f_s_dadda_rca24_and_4_18_y0;
  wire f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_6_16_y0;
  wire f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_5_17_y0;
  wire f_s_dadda_rca24_fa149_y0;
  wire f_s_dadda_rca24_fa149_y1;
  wire f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_4_18_y0;
  wire f_s_dadda_rca24_fa149_y2;
  wire f_s_dadda_rca24_fa149_y3;
  wire f_s_dadda_rca24_fa149_y4;
  wire f_s_dadda_rca24_and_3_19_a_3;
  wire f_s_dadda_rca24_and_3_19_b_19;
  wire f_s_dadda_rca24_and_3_19_y0;
  wire f_s_dadda_rca24_and_2_20_a_2;
  wire f_s_dadda_rca24_and_2_20_b_20;
  wire f_s_dadda_rca24_and_2_20_y0;
  wire f_s_dadda_rca24_and_1_21_a_1;
  wire f_s_dadda_rca24_and_1_21_b_21;
  wire f_s_dadda_rca24_and_1_21_y0;
  wire f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_3_19_y0;
  wire f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_2_20_y0;
  wire f_s_dadda_rca24_fa150_y0;
  wire f_s_dadda_rca24_fa150_y1;
  wire f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_1_21_y0;
  wire f_s_dadda_rca24_fa150_y2;
  wire f_s_dadda_rca24_fa150_y3;
  wire f_s_dadda_rca24_fa150_y4;
  wire f_s_dadda_rca24_and_0_22_a_0;
  wire f_s_dadda_rca24_and_0_22_b_22;
  wire f_s_dadda_rca24_and_0_22_y0;
  wire f_s_dadda_rca24_fa151_f_s_dadda_rca24_and_0_22_y0;
  wire f_s_dadda_rca24_fa151_f_s_dadda_rca24_fa3_y2;
  wire f_s_dadda_rca24_fa151_y0;
  wire f_s_dadda_rca24_fa151_y1;
  wire f_s_dadda_rca24_fa151_f_s_dadda_rca24_fa4_y2;
  wire f_s_dadda_rca24_fa151_y2;
  wire f_s_dadda_rca24_fa151_y3;
  wire f_s_dadda_rca24_fa151_y4;
  wire f_s_dadda_rca24_fa152_f_s_dadda_rca24_fa5_y2;
  wire f_s_dadda_rca24_fa152_f_s_dadda_rca24_ha3_y0;
  wire f_s_dadda_rca24_fa152_y0;
  wire f_s_dadda_rca24_fa152_y1;
  wire f_s_dadda_rca24_fa152_f_s_dadda_rca24_fa142_y2;
  wire f_s_dadda_rca24_fa152_y2;
  wire f_s_dadda_rca24_fa152_y3;
  wire f_s_dadda_rca24_fa152_y4;
  wire f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa143_y2;
  wire f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa144_y2;
  wire f_s_dadda_rca24_fa153_y0;
  wire f_s_dadda_rca24_fa153_y1;
  wire f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa145_y2;
  wire f_s_dadda_rca24_fa153_y2;
  wire f_s_dadda_rca24_fa153_y3;
  wire f_s_dadda_rca24_fa153_y4;
  wire f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa146_y2;
  wire f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa147_y2;
  wire f_s_dadda_rca24_fa154_y0;
  wire f_s_dadda_rca24_fa154_y1;
  wire f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa148_y2;
  wire f_s_dadda_rca24_fa154_y2;
  wire f_s_dadda_rca24_fa154_y3;
  wire f_s_dadda_rca24_fa154_y4;
  wire f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa154_y4;
  wire f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa153_y4;
  wire f_s_dadda_rca24_fa155_y0;
  wire f_s_dadda_rca24_fa155_y1;
  wire f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa152_y4;
  wire f_s_dadda_rca24_fa155_y2;
  wire f_s_dadda_rca24_fa155_y3;
  wire f_s_dadda_rca24_fa155_y4;
  wire f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa151_y4;
  wire f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa150_y4;
  wire f_s_dadda_rca24_fa156_y0;
  wire f_s_dadda_rca24_fa156_y1;
  wire f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa149_y4;
  wire f_s_dadda_rca24_fa156_y2;
  wire f_s_dadda_rca24_fa156_y3;
  wire f_s_dadda_rca24_fa156_y4;
  wire f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa148_y4;
  wire f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa147_y4;
  wire f_s_dadda_rca24_fa157_y0;
  wire f_s_dadda_rca24_fa157_y1;
  wire f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa146_y4;
  wire f_s_dadda_rca24_fa157_y2;
  wire f_s_dadda_rca24_fa157_y3;
  wire f_s_dadda_rca24_fa157_y4;
  wire f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa145_y4;
  wire f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa144_y4;
  wire f_s_dadda_rca24_fa158_y0;
  wire f_s_dadda_rca24_fa158_y1;
  wire f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa143_y4;
  wire f_s_dadda_rca24_fa158_y2;
  wire f_s_dadda_rca24_fa158_y3;
  wire f_s_dadda_rca24_fa158_y4;
  wire f_s_dadda_rca24_and_13_10_a_13;
  wire f_s_dadda_rca24_and_13_10_b_10;
  wire f_s_dadda_rca24_and_13_10_y0;
  wire f_s_dadda_rca24_and_12_11_a_12;
  wire f_s_dadda_rca24_and_12_11_b_11;
  wire f_s_dadda_rca24_and_12_11_y0;
  wire f_s_dadda_rca24_fa159_f_s_dadda_rca24_fa142_y4;
  wire f_s_dadda_rca24_fa159_f_s_dadda_rca24_and_13_10_y0;
  wire f_s_dadda_rca24_fa159_y0;
  wire f_s_dadda_rca24_fa159_y1;
  wire f_s_dadda_rca24_fa159_f_s_dadda_rca24_and_12_11_y0;
  wire f_s_dadda_rca24_fa159_y2;
  wire f_s_dadda_rca24_fa159_y3;
  wire f_s_dadda_rca24_fa159_y4;
  wire f_s_dadda_rca24_and_11_12_a_11;
  wire f_s_dadda_rca24_and_11_12_b_12;
  wire f_s_dadda_rca24_and_11_12_y0;
  wire f_s_dadda_rca24_and_10_13_a_10;
  wire f_s_dadda_rca24_and_10_13_b_13;
  wire f_s_dadda_rca24_and_10_13_y0;
  wire f_s_dadda_rca24_and_9_14_a_9;
  wire f_s_dadda_rca24_and_9_14_b_14;
  wire f_s_dadda_rca24_and_9_14_y0;
  wire f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_11_12_y0;
  wire f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_10_13_y0;
  wire f_s_dadda_rca24_fa160_y0;
  wire f_s_dadda_rca24_fa160_y1;
  wire f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_9_14_y0;
  wire f_s_dadda_rca24_fa160_y2;
  wire f_s_dadda_rca24_fa160_y3;
  wire f_s_dadda_rca24_fa160_y4;
  wire f_s_dadda_rca24_and_8_15_a_8;
  wire f_s_dadda_rca24_and_8_15_b_15;
  wire f_s_dadda_rca24_and_8_15_y0;
  wire f_s_dadda_rca24_and_7_16_a_7;
  wire f_s_dadda_rca24_and_7_16_b_16;
  wire f_s_dadda_rca24_and_7_16_y0;
  wire f_s_dadda_rca24_and_6_17_a_6;
  wire f_s_dadda_rca24_and_6_17_b_17;
  wire f_s_dadda_rca24_and_6_17_y0;
  wire f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_8_15_y0;
  wire f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_7_16_y0;
  wire f_s_dadda_rca24_fa161_y0;
  wire f_s_dadda_rca24_fa161_y1;
  wire f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_6_17_y0;
  wire f_s_dadda_rca24_fa161_y2;
  wire f_s_dadda_rca24_fa161_y3;
  wire f_s_dadda_rca24_fa161_y4;
  wire f_s_dadda_rca24_and_5_18_a_5;
  wire f_s_dadda_rca24_and_5_18_b_18;
  wire f_s_dadda_rca24_and_5_18_y0;
  wire f_s_dadda_rca24_and_4_19_a_4;
  wire f_s_dadda_rca24_and_4_19_b_19;
  wire f_s_dadda_rca24_and_4_19_y0;
  wire f_s_dadda_rca24_and_3_20_a_3;
  wire f_s_dadda_rca24_and_3_20_b_20;
  wire f_s_dadda_rca24_and_3_20_y0;
  wire f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_5_18_y0;
  wire f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_4_19_y0;
  wire f_s_dadda_rca24_fa162_y0;
  wire f_s_dadda_rca24_fa162_y1;
  wire f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_3_20_y0;
  wire f_s_dadda_rca24_fa162_y2;
  wire f_s_dadda_rca24_fa162_y3;
  wire f_s_dadda_rca24_fa162_y4;
  wire f_s_dadda_rca24_and_2_21_a_2;
  wire f_s_dadda_rca24_and_2_21_b_21;
  wire f_s_dadda_rca24_and_2_21_y0;
  wire f_s_dadda_rca24_and_1_22_a_1;
  wire f_s_dadda_rca24_and_1_22_b_22;
  wire f_s_dadda_rca24_and_1_22_y0;
  wire f_s_dadda_rca24_nand_0_23_a_0;
  wire f_s_dadda_rca24_nand_0_23_b_23;
  wire f_s_dadda_rca24_nand_0_23_y0;
  wire f_s_dadda_rca24_fa163_f_s_dadda_rca24_and_2_21_y0;
  wire f_s_dadda_rca24_fa163_f_s_dadda_rca24_and_1_22_y0;
  wire f_s_dadda_rca24_fa163_y0;
  wire f_s_dadda_rca24_fa163_y1;
  wire f_s_dadda_rca24_fa163_f_s_dadda_rca24_nand_0_23_y0;
  wire f_s_dadda_rca24_fa163_y2;
  wire f_s_dadda_rca24_fa163_y3;
  wire f_s_dadda_rca24_fa163_y4;
  wire f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa6_y2;
  wire f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa7_y2;
  wire f_s_dadda_rca24_fa164_y0;
  wire f_s_dadda_rca24_fa164_y1;
  wire f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa8_y2;
  wire f_s_dadda_rca24_fa164_y2;
  wire f_s_dadda_rca24_fa164_y3;
  wire f_s_dadda_rca24_fa164_y4;
  wire f_s_dadda_rca24_fa165_f_s_dadda_rca24_fa9_y2;
  wire f_s_dadda_rca24_fa165_f_s_dadda_rca24_ha4_y0;
  wire f_s_dadda_rca24_fa165_y0;
  wire f_s_dadda_rca24_fa165_y1;
  wire f_s_dadda_rca24_fa165_f_s_dadda_rca24_fa155_y2;
  wire f_s_dadda_rca24_fa165_y2;
  wire f_s_dadda_rca24_fa165_y3;
  wire f_s_dadda_rca24_fa165_y4;
  wire f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa156_y2;
  wire f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa157_y2;
  wire f_s_dadda_rca24_fa166_y0;
  wire f_s_dadda_rca24_fa166_y1;
  wire f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa158_y2;
  wire f_s_dadda_rca24_fa166_y2;
  wire f_s_dadda_rca24_fa166_y3;
  wire f_s_dadda_rca24_fa166_y4;
  wire f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa159_y2;
  wire f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa160_y2;
  wire f_s_dadda_rca24_fa167_y0;
  wire f_s_dadda_rca24_fa167_y1;
  wire f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa161_y2;
  wire f_s_dadda_rca24_fa167_y2;
  wire f_s_dadda_rca24_fa167_y3;
  wire f_s_dadda_rca24_fa167_y4;
  wire f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa167_y4;
  wire f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa166_y4;
  wire f_s_dadda_rca24_fa168_y0;
  wire f_s_dadda_rca24_fa168_y1;
  wire f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa165_y4;
  wire f_s_dadda_rca24_fa168_y2;
  wire f_s_dadda_rca24_fa168_y3;
  wire f_s_dadda_rca24_fa168_y4;
  wire f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa164_y4;
  wire f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa163_y4;
  wire f_s_dadda_rca24_fa169_y0;
  wire f_s_dadda_rca24_fa169_y1;
  wire f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa162_y4;
  wire f_s_dadda_rca24_fa169_y2;
  wire f_s_dadda_rca24_fa169_y3;
  wire f_s_dadda_rca24_fa169_y4;
  wire f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa161_y4;
  wire f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa160_y4;
  wire f_s_dadda_rca24_fa170_y0;
  wire f_s_dadda_rca24_fa170_y1;
  wire f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa159_y4;
  wire f_s_dadda_rca24_fa170_y2;
  wire f_s_dadda_rca24_fa170_y3;
  wire f_s_dadda_rca24_fa170_y4;
  wire f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa158_y4;
  wire f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa157_y4;
  wire f_s_dadda_rca24_fa171_y0;
  wire f_s_dadda_rca24_fa171_y1;
  wire f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa156_y4;
  wire f_s_dadda_rca24_fa171_y2;
  wire f_s_dadda_rca24_fa171_y3;
  wire f_s_dadda_rca24_fa171_y4;
  wire f_s_dadda_rca24_and_14_10_a_14;
  wire f_s_dadda_rca24_and_14_10_b_10;
  wire f_s_dadda_rca24_and_14_10_y0;
  wire f_s_dadda_rca24_and_13_11_a_13;
  wire f_s_dadda_rca24_and_13_11_b_11;
  wire f_s_dadda_rca24_and_13_11_y0;
  wire f_s_dadda_rca24_fa172_f_s_dadda_rca24_fa155_y4;
  wire f_s_dadda_rca24_fa172_f_s_dadda_rca24_and_14_10_y0;
  wire f_s_dadda_rca24_fa172_y0;
  wire f_s_dadda_rca24_fa172_y1;
  wire f_s_dadda_rca24_fa172_f_s_dadda_rca24_and_13_11_y0;
  wire f_s_dadda_rca24_fa172_y2;
  wire f_s_dadda_rca24_fa172_y3;
  wire f_s_dadda_rca24_fa172_y4;
  wire f_s_dadda_rca24_and_12_12_a_12;
  wire f_s_dadda_rca24_and_12_12_b_12;
  wire f_s_dadda_rca24_and_12_12_y0;
  wire f_s_dadda_rca24_and_11_13_a_11;
  wire f_s_dadda_rca24_and_11_13_b_13;
  wire f_s_dadda_rca24_and_11_13_y0;
  wire f_s_dadda_rca24_and_10_14_a_10;
  wire f_s_dadda_rca24_and_10_14_b_14;
  wire f_s_dadda_rca24_and_10_14_y0;
  wire f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_12_12_y0;
  wire f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_11_13_y0;
  wire f_s_dadda_rca24_fa173_y0;
  wire f_s_dadda_rca24_fa173_y1;
  wire f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_10_14_y0;
  wire f_s_dadda_rca24_fa173_y2;
  wire f_s_dadda_rca24_fa173_y3;
  wire f_s_dadda_rca24_fa173_y4;
  wire f_s_dadda_rca24_and_9_15_a_9;
  wire f_s_dadda_rca24_and_9_15_b_15;
  wire f_s_dadda_rca24_and_9_15_y0;
  wire f_s_dadda_rca24_and_8_16_a_8;
  wire f_s_dadda_rca24_and_8_16_b_16;
  wire f_s_dadda_rca24_and_8_16_y0;
  wire f_s_dadda_rca24_and_7_17_a_7;
  wire f_s_dadda_rca24_and_7_17_b_17;
  wire f_s_dadda_rca24_and_7_17_y0;
  wire f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_9_15_y0;
  wire f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_8_16_y0;
  wire f_s_dadda_rca24_fa174_y0;
  wire f_s_dadda_rca24_fa174_y1;
  wire f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_7_17_y0;
  wire f_s_dadda_rca24_fa174_y2;
  wire f_s_dadda_rca24_fa174_y3;
  wire f_s_dadda_rca24_fa174_y4;
  wire f_s_dadda_rca24_and_6_18_a_6;
  wire f_s_dadda_rca24_and_6_18_b_18;
  wire f_s_dadda_rca24_and_6_18_y0;
  wire f_s_dadda_rca24_and_5_19_a_5;
  wire f_s_dadda_rca24_and_5_19_b_19;
  wire f_s_dadda_rca24_and_5_19_y0;
  wire f_s_dadda_rca24_and_4_20_a_4;
  wire f_s_dadda_rca24_and_4_20_b_20;
  wire f_s_dadda_rca24_and_4_20_y0;
  wire f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_6_18_y0;
  wire f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_5_19_y0;
  wire f_s_dadda_rca24_fa175_y0;
  wire f_s_dadda_rca24_fa175_y1;
  wire f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_4_20_y0;
  wire f_s_dadda_rca24_fa175_y2;
  wire f_s_dadda_rca24_fa175_y3;
  wire f_s_dadda_rca24_fa175_y4;
  wire f_s_dadda_rca24_and_3_21_a_3;
  wire f_s_dadda_rca24_and_3_21_b_21;
  wire f_s_dadda_rca24_and_3_21_y0;
  wire f_s_dadda_rca24_and_2_22_a_2;
  wire f_s_dadda_rca24_and_2_22_b_22;
  wire f_s_dadda_rca24_and_2_22_y0;
  wire f_s_dadda_rca24_nand_1_23_a_1;
  wire f_s_dadda_rca24_nand_1_23_b_23;
  wire f_s_dadda_rca24_nand_1_23_y0;
  wire f_s_dadda_rca24_fa176_f_s_dadda_rca24_and_3_21_y0;
  wire f_s_dadda_rca24_fa176_f_s_dadda_rca24_and_2_22_y0;
  wire f_s_dadda_rca24_fa176_y0;
  wire f_s_dadda_rca24_fa176_y1;
  wire f_s_dadda_rca24_fa176_f_s_dadda_rca24_nand_1_23_y0;
  wire f_s_dadda_rca24_fa176_y2;
  wire f_s_dadda_rca24_fa176_y3;
  wire f_s_dadda_rca24_fa176_y4;
  wire f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa10_y2;
  wire f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa11_y2;
  wire f_s_dadda_rca24_fa177_y0;
  wire f_s_dadda_rca24_fa177_y1;
  wire f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa12_y2;
  wire f_s_dadda_rca24_fa177_y2;
  wire f_s_dadda_rca24_fa177_y3;
  wire f_s_dadda_rca24_fa177_y4;
  wire f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa13_y2;
  wire f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa14_y2;
  wire f_s_dadda_rca24_fa178_y0;
  wire f_s_dadda_rca24_fa178_y1;
  wire f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa168_y2;
  wire f_s_dadda_rca24_fa178_y2;
  wire f_s_dadda_rca24_fa178_y3;
  wire f_s_dadda_rca24_fa178_y4;
  wire f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa169_y2;
  wire f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa170_y2;
  wire f_s_dadda_rca24_fa179_y0;
  wire f_s_dadda_rca24_fa179_y1;
  wire f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa171_y2;
  wire f_s_dadda_rca24_fa179_y2;
  wire f_s_dadda_rca24_fa179_y3;
  wire f_s_dadda_rca24_fa179_y4;
  wire f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa172_y2;
  wire f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa173_y2;
  wire f_s_dadda_rca24_fa180_y0;
  wire f_s_dadda_rca24_fa180_y1;
  wire f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa174_y2;
  wire f_s_dadda_rca24_fa180_y2;
  wire f_s_dadda_rca24_fa180_y3;
  wire f_s_dadda_rca24_fa180_y4;
  wire f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa180_y4;
  wire f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa179_y4;
  wire f_s_dadda_rca24_fa181_y0;
  wire f_s_dadda_rca24_fa181_y1;
  wire f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa178_y4;
  wire f_s_dadda_rca24_fa181_y2;
  wire f_s_dadda_rca24_fa181_y3;
  wire f_s_dadda_rca24_fa181_y4;
  wire f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa177_y4;
  wire f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa176_y4;
  wire f_s_dadda_rca24_fa182_y0;
  wire f_s_dadda_rca24_fa182_y1;
  wire f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa175_y4;
  wire f_s_dadda_rca24_fa182_y2;
  wire f_s_dadda_rca24_fa182_y3;
  wire f_s_dadda_rca24_fa182_y4;
  wire f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa174_y4;
  wire f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa173_y4;
  wire f_s_dadda_rca24_fa183_y0;
  wire f_s_dadda_rca24_fa183_y1;
  wire f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa172_y4;
  wire f_s_dadda_rca24_fa183_y2;
  wire f_s_dadda_rca24_fa183_y3;
  wire f_s_dadda_rca24_fa183_y4;
  wire f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa171_y4;
  wire f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa170_y4;
  wire f_s_dadda_rca24_fa184_y0;
  wire f_s_dadda_rca24_fa184_y1;
  wire f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa169_y4;
  wire f_s_dadda_rca24_fa184_y2;
  wire f_s_dadda_rca24_fa184_y3;
  wire f_s_dadda_rca24_fa184_y4;
  wire f_s_dadda_rca24_and_16_9_a_16;
  wire f_s_dadda_rca24_and_16_9_b_9;
  wire f_s_dadda_rca24_and_16_9_y0;
  wire f_s_dadda_rca24_and_15_10_a_15;
  wire f_s_dadda_rca24_and_15_10_b_10;
  wire f_s_dadda_rca24_and_15_10_y0;
  wire f_s_dadda_rca24_fa185_f_s_dadda_rca24_fa168_y4;
  wire f_s_dadda_rca24_fa185_f_s_dadda_rca24_and_16_9_y0;
  wire f_s_dadda_rca24_fa185_y0;
  wire f_s_dadda_rca24_fa185_y1;
  wire f_s_dadda_rca24_fa185_f_s_dadda_rca24_and_15_10_y0;
  wire f_s_dadda_rca24_fa185_y2;
  wire f_s_dadda_rca24_fa185_y3;
  wire f_s_dadda_rca24_fa185_y4;
  wire f_s_dadda_rca24_and_14_11_a_14;
  wire f_s_dadda_rca24_and_14_11_b_11;
  wire f_s_dadda_rca24_and_14_11_y0;
  wire f_s_dadda_rca24_and_13_12_a_13;
  wire f_s_dadda_rca24_and_13_12_b_12;
  wire f_s_dadda_rca24_and_13_12_y0;
  wire f_s_dadda_rca24_and_12_13_a_12;
  wire f_s_dadda_rca24_and_12_13_b_13;
  wire f_s_dadda_rca24_and_12_13_y0;
  wire f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_14_11_y0;
  wire f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_13_12_y0;
  wire f_s_dadda_rca24_fa186_y0;
  wire f_s_dadda_rca24_fa186_y1;
  wire f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_12_13_y0;
  wire f_s_dadda_rca24_fa186_y2;
  wire f_s_dadda_rca24_fa186_y3;
  wire f_s_dadda_rca24_fa186_y4;
  wire f_s_dadda_rca24_and_11_14_a_11;
  wire f_s_dadda_rca24_and_11_14_b_14;
  wire f_s_dadda_rca24_and_11_14_y0;
  wire f_s_dadda_rca24_and_10_15_a_10;
  wire f_s_dadda_rca24_and_10_15_b_15;
  wire f_s_dadda_rca24_and_10_15_y0;
  wire f_s_dadda_rca24_and_9_16_a_9;
  wire f_s_dadda_rca24_and_9_16_b_16;
  wire f_s_dadda_rca24_and_9_16_y0;
  wire f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_11_14_y0;
  wire f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_10_15_y0;
  wire f_s_dadda_rca24_fa187_y0;
  wire f_s_dadda_rca24_fa187_y1;
  wire f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_9_16_y0;
  wire f_s_dadda_rca24_fa187_y2;
  wire f_s_dadda_rca24_fa187_y3;
  wire f_s_dadda_rca24_fa187_y4;
  wire f_s_dadda_rca24_and_8_17_a_8;
  wire f_s_dadda_rca24_and_8_17_b_17;
  wire f_s_dadda_rca24_and_8_17_y0;
  wire f_s_dadda_rca24_and_7_18_a_7;
  wire f_s_dadda_rca24_and_7_18_b_18;
  wire f_s_dadda_rca24_and_7_18_y0;
  wire f_s_dadda_rca24_and_6_19_a_6;
  wire f_s_dadda_rca24_and_6_19_b_19;
  wire f_s_dadda_rca24_and_6_19_y0;
  wire f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_8_17_y0;
  wire f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_7_18_y0;
  wire f_s_dadda_rca24_fa188_y0;
  wire f_s_dadda_rca24_fa188_y1;
  wire f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_6_19_y0;
  wire f_s_dadda_rca24_fa188_y2;
  wire f_s_dadda_rca24_fa188_y3;
  wire f_s_dadda_rca24_fa188_y4;
  wire f_s_dadda_rca24_and_5_20_a_5;
  wire f_s_dadda_rca24_and_5_20_b_20;
  wire f_s_dadda_rca24_and_5_20_y0;
  wire f_s_dadda_rca24_and_4_21_a_4;
  wire f_s_dadda_rca24_and_4_21_b_21;
  wire f_s_dadda_rca24_and_4_21_y0;
  wire f_s_dadda_rca24_and_3_22_a_3;
  wire f_s_dadda_rca24_and_3_22_b_22;
  wire f_s_dadda_rca24_and_3_22_y0;
  wire f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_5_20_y0;
  wire f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_4_21_y0;
  wire f_s_dadda_rca24_fa189_y0;
  wire f_s_dadda_rca24_fa189_y1;
  wire f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_3_22_y0;
  wire f_s_dadda_rca24_fa189_y2;
  wire f_s_dadda_rca24_fa189_y3;
  wire f_s_dadda_rca24_fa189_y4;
  wire f_s_dadda_rca24_nand_2_23_a_2;
  wire f_s_dadda_rca24_nand_2_23_b_23;
  wire f_s_dadda_rca24_nand_2_23_y0;
  wire f_s_dadda_rca24_fa190_f_s_dadda_rca24_nand_2_23_y0;
  wire f_s_dadda_rca24_fa190_f_s_dadda_rca24_fa15_y2;
  wire f_s_dadda_rca24_fa190_y0;
  wire f_s_dadda_rca24_fa190_y1;
  wire f_s_dadda_rca24_fa190_f_s_dadda_rca24_fa16_y2;
  wire f_s_dadda_rca24_fa190_y2;
  wire f_s_dadda_rca24_fa190_y3;
  wire f_s_dadda_rca24_fa190_y4;
  wire f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa17_y2;
  wire f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa18_y2;
  wire f_s_dadda_rca24_fa191_y0;
  wire f_s_dadda_rca24_fa191_y1;
  wire f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa181_y2;
  wire f_s_dadda_rca24_fa191_y2;
  wire f_s_dadda_rca24_fa191_y3;
  wire f_s_dadda_rca24_fa191_y4;
  wire f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa182_y2;
  wire f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa183_y2;
  wire f_s_dadda_rca24_fa192_y0;
  wire f_s_dadda_rca24_fa192_y1;
  wire f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa184_y2;
  wire f_s_dadda_rca24_fa192_y2;
  wire f_s_dadda_rca24_fa192_y3;
  wire f_s_dadda_rca24_fa192_y4;
  wire f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa185_y2;
  wire f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa186_y2;
  wire f_s_dadda_rca24_fa193_y0;
  wire f_s_dadda_rca24_fa193_y1;
  wire f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa187_y2;
  wire f_s_dadda_rca24_fa193_y2;
  wire f_s_dadda_rca24_fa193_y3;
  wire f_s_dadda_rca24_fa193_y4;
  wire f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa193_y4;
  wire f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa192_y4;
  wire f_s_dadda_rca24_fa194_y0;
  wire f_s_dadda_rca24_fa194_y1;
  wire f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa191_y4;
  wire f_s_dadda_rca24_fa194_y2;
  wire f_s_dadda_rca24_fa194_y3;
  wire f_s_dadda_rca24_fa194_y4;
  wire f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa190_y4;
  wire f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa189_y4;
  wire f_s_dadda_rca24_fa195_y0;
  wire f_s_dadda_rca24_fa195_y1;
  wire f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa188_y4;
  wire f_s_dadda_rca24_fa195_y2;
  wire f_s_dadda_rca24_fa195_y3;
  wire f_s_dadda_rca24_fa195_y4;
  wire f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa187_y4;
  wire f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa186_y4;
  wire f_s_dadda_rca24_fa196_y0;
  wire f_s_dadda_rca24_fa196_y1;
  wire f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa185_y4;
  wire f_s_dadda_rca24_fa196_y2;
  wire f_s_dadda_rca24_fa196_y3;
  wire f_s_dadda_rca24_fa196_y4;
  wire f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa184_y4;
  wire f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa183_y4;
  wire f_s_dadda_rca24_fa197_y0;
  wire f_s_dadda_rca24_fa197_y1;
  wire f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa182_y4;
  wire f_s_dadda_rca24_fa197_y2;
  wire f_s_dadda_rca24_fa197_y3;
  wire f_s_dadda_rca24_fa197_y4;
  wire f_s_dadda_rca24_and_18_8_a_18;
  wire f_s_dadda_rca24_and_18_8_b_8;
  wire f_s_dadda_rca24_and_18_8_y0;
  wire f_s_dadda_rca24_and_17_9_a_17;
  wire f_s_dadda_rca24_and_17_9_b_9;
  wire f_s_dadda_rca24_and_17_9_y0;
  wire f_s_dadda_rca24_fa198_f_s_dadda_rca24_fa181_y4;
  wire f_s_dadda_rca24_fa198_f_s_dadda_rca24_and_18_8_y0;
  wire f_s_dadda_rca24_fa198_y0;
  wire f_s_dadda_rca24_fa198_y1;
  wire f_s_dadda_rca24_fa198_f_s_dadda_rca24_and_17_9_y0;
  wire f_s_dadda_rca24_fa198_y2;
  wire f_s_dadda_rca24_fa198_y3;
  wire f_s_dadda_rca24_fa198_y4;
  wire f_s_dadda_rca24_and_16_10_a_16;
  wire f_s_dadda_rca24_and_16_10_b_10;
  wire f_s_dadda_rca24_and_16_10_y0;
  wire f_s_dadda_rca24_and_15_11_a_15;
  wire f_s_dadda_rca24_and_15_11_b_11;
  wire f_s_dadda_rca24_and_15_11_y0;
  wire f_s_dadda_rca24_and_14_12_a_14;
  wire f_s_dadda_rca24_and_14_12_b_12;
  wire f_s_dadda_rca24_and_14_12_y0;
  wire f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_16_10_y0;
  wire f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_15_11_y0;
  wire f_s_dadda_rca24_fa199_y0;
  wire f_s_dadda_rca24_fa199_y1;
  wire f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_14_12_y0;
  wire f_s_dadda_rca24_fa199_y2;
  wire f_s_dadda_rca24_fa199_y3;
  wire f_s_dadda_rca24_fa199_y4;
  wire f_s_dadda_rca24_and_13_13_a_13;
  wire f_s_dadda_rca24_and_13_13_b_13;
  wire f_s_dadda_rca24_and_13_13_y0;
  wire f_s_dadda_rca24_and_12_14_a_12;
  wire f_s_dadda_rca24_and_12_14_b_14;
  wire f_s_dadda_rca24_and_12_14_y0;
  wire f_s_dadda_rca24_and_11_15_a_11;
  wire f_s_dadda_rca24_and_11_15_b_15;
  wire f_s_dadda_rca24_and_11_15_y0;
  wire f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_13_13_y0;
  wire f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_12_14_y0;
  wire f_s_dadda_rca24_fa200_y0;
  wire f_s_dadda_rca24_fa200_y1;
  wire f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_11_15_y0;
  wire f_s_dadda_rca24_fa200_y2;
  wire f_s_dadda_rca24_fa200_y3;
  wire f_s_dadda_rca24_fa200_y4;
  wire f_s_dadda_rca24_and_10_16_a_10;
  wire f_s_dadda_rca24_and_10_16_b_16;
  wire f_s_dadda_rca24_and_10_16_y0;
  wire f_s_dadda_rca24_and_9_17_a_9;
  wire f_s_dadda_rca24_and_9_17_b_17;
  wire f_s_dadda_rca24_and_9_17_y0;
  wire f_s_dadda_rca24_and_8_18_a_8;
  wire f_s_dadda_rca24_and_8_18_b_18;
  wire f_s_dadda_rca24_and_8_18_y0;
  wire f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_10_16_y0;
  wire f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_9_17_y0;
  wire f_s_dadda_rca24_fa201_y0;
  wire f_s_dadda_rca24_fa201_y1;
  wire f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_8_18_y0;
  wire f_s_dadda_rca24_fa201_y2;
  wire f_s_dadda_rca24_fa201_y3;
  wire f_s_dadda_rca24_fa201_y4;
  wire f_s_dadda_rca24_and_7_19_a_7;
  wire f_s_dadda_rca24_and_7_19_b_19;
  wire f_s_dadda_rca24_and_7_19_y0;
  wire f_s_dadda_rca24_and_6_20_a_6;
  wire f_s_dadda_rca24_and_6_20_b_20;
  wire f_s_dadda_rca24_and_6_20_y0;
  wire f_s_dadda_rca24_and_5_21_a_5;
  wire f_s_dadda_rca24_and_5_21_b_21;
  wire f_s_dadda_rca24_and_5_21_y0;
  wire f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_7_19_y0;
  wire f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_6_20_y0;
  wire f_s_dadda_rca24_fa202_y0;
  wire f_s_dadda_rca24_fa202_y1;
  wire f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_5_21_y0;
  wire f_s_dadda_rca24_fa202_y2;
  wire f_s_dadda_rca24_fa202_y3;
  wire f_s_dadda_rca24_fa202_y4;
  wire f_s_dadda_rca24_and_4_22_a_4;
  wire f_s_dadda_rca24_and_4_22_b_22;
  wire f_s_dadda_rca24_and_4_22_y0;
  wire f_s_dadda_rca24_nand_3_23_a_3;
  wire f_s_dadda_rca24_nand_3_23_b_23;
  wire f_s_dadda_rca24_nand_3_23_y0;
  wire f_s_dadda_rca24_fa203_f_s_dadda_rca24_and_4_22_y0;
  wire f_s_dadda_rca24_fa203_f_s_dadda_rca24_nand_3_23_y0;
  wire f_s_dadda_rca24_fa203_y0;
  wire f_s_dadda_rca24_fa203_y1;
  wire f_s_dadda_rca24_fa203_f_s_dadda_rca24_fa19_y2;
  wire f_s_dadda_rca24_fa203_y2;
  wire f_s_dadda_rca24_fa203_y3;
  wire f_s_dadda_rca24_fa203_y4;
  wire f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa20_y2;
  wire f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa21_y2;
  wire f_s_dadda_rca24_fa204_y0;
  wire f_s_dadda_rca24_fa204_y1;
  wire f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa194_y2;
  wire f_s_dadda_rca24_fa204_y2;
  wire f_s_dadda_rca24_fa204_y3;
  wire f_s_dadda_rca24_fa204_y4;
  wire f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa195_y2;
  wire f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa196_y2;
  wire f_s_dadda_rca24_fa205_y0;
  wire f_s_dadda_rca24_fa205_y1;
  wire f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa197_y2;
  wire f_s_dadda_rca24_fa205_y2;
  wire f_s_dadda_rca24_fa205_y3;
  wire f_s_dadda_rca24_fa205_y4;
  wire f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa198_y2;
  wire f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa199_y2;
  wire f_s_dadda_rca24_fa206_y0;
  wire f_s_dadda_rca24_fa206_y1;
  wire f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa200_y2;
  wire f_s_dadda_rca24_fa206_y2;
  wire f_s_dadda_rca24_fa206_y3;
  wire f_s_dadda_rca24_fa206_y4;
  wire f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa206_y4;
  wire f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa205_y4;
  wire f_s_dadda_rca24_fa207_y0;
  wire f_s_dadda_rca24_fa207_y1;
  wire f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa204_y4;
  wire f_s_dadda_rca24_fa207_y2;
  wire f_s_dadda_rca24_fa207_y3;
  wire f_s_dadda_rca24_fa207_y4;
  wire f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa203_y4;
  wire f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa202_y4;
  wire f_s_dadda_rca24_fa208_y0;
  wire f_s_dadda_rca24_fa208_y1;
  wire f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa201_y4;
  wire f_s_dadda_rca24_fa208_y2;
  wire f_s_dadda_rca24_fa208_y3;
  wire f_s_dadda_rca24_fa208_y4;
  wire f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa200_y4;
  wire f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa199_y4;
  wire f_s_dadda_rca24_fa209_y0;
  wire f_s_dadda_rca24_fa209_y1;
  wire f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa198_y4;
  wire f_s_dadda_rca24_fa209_y2;
  wire f_s_dadda_rca24_fa209_y3;
  wire f_s_dadda_rca24_fa209_y4;
  wire f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa197_y4;
  wire f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa196_y4;
  wire f_s_dadda_rca24_fa210_y0;
  wire f_s_dadda_rca24_fa210_y1;
  wire f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa195_y4;
  wire f_s_dadda_rca24_fa210_y2;
  wire f_s_dadda_rca24_fa210_y3;
  wire f_s_dadda_rca24_fa210_y4;
  wire f_s_dadda_rca24_and_20_7_a_20;
  wire f_s_dadda_rca24_and_20_7_b_7;
  wire f_s_dadda_rca24_and_20_7_y0;
  wire f_s_dadda_rca24_and_19_8_a_19;
  wire f_s_dadda_rca24_and_19_8_b_8;
  wire f_s_dadda_rca24_and_19_8_y0;
  wire f_s_dadda_rca24_fa211_f_s_dadda_rca24_fa194_y4;
  wire f_s_dadda_rca24_fa211_f_s_dadda_rca24_and_20_7_y0;
  wire f_s_dadda_rca24_fa211_y0;
  wire f_s_dadda_rca24_fa211_y1;
  wire f_s_dadda_rca24_fa211_f_s_dadda_rca24_and_19_8_y0;
  wire f_s_dadda_rca24_fa211_y2;
  wire f_s_dadda_rca24_fa211_y3;
  wire f_s_dadda_rca24_fa211_y4;
  wire f_s_dadda_rca24_and_18_9_a_18;
  wire f_s_dadda_rca24_and_18_9_b_9;
  wire f_s_dadda_rca24_and_18_9_y0;
  wire f_s_dadda_rca24_and_17_10_a_17;
  wire f_s_dadda_rca24_and_17_10_b_10;
  wire f_s_dadda_rca24_and_17_10_y0;
  wire f_s_dadda_rca24_and_16_11_a_16;
  wire f_s_dadda_rca24_and_16_11_b_11;
  wire f_s_dadda_rca24_and_16_11_y0;
  wire f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_18_9_y0;
  wire f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_17_10_y0;
  wire f_s_dadda_rca24_fa212_y0;
  wire f_s_dadda_rca24_fa212_y1;
  wire f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_16_11_y0;
  wire f_s_dadda_rca24_fa212_y2;
  wire f_s_dadda_rca24_fa212_y3;
  wire f_s_dadda_rca24_fa212_y4;
  wire f_s_dadda_rca24_and_15_12_a_15;
  wire f_s_dadda_rca24_and_15_12_b_12;
  wire f_s_dadda_rca24_and_15_12_y0;
  wire f_s_dadda_rca24_and_14_13_a_14;
  wire f_s_dadda_rca24_and_14_13_b_13;
  wire f_s_dadda_rca24_and_14_13_y0;
  wire f_s_dadda_rca24_and_13_14_a_13;
  wire f_s_dadda_rca24_and_13_14_b_14;
  wire f_s_dadda_rca24_and_13_14_y0;
  wire f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_15_12_y0;
  wire f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_14_13_y0;
  wire f_s_dadda_rca24_fa213_y0;
  wire f_s_dadda_rca24_fa213_y1;
  wire f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_13_14_y0;
  wire f_s_dadda_rca24_fa213_y2;
  wire f_s_dadda_rca24_fa213_y3;
  wire f_s_dadda_rca24_fa213_y4;
  wire f_s_dadda_rca24_and_12_15_a_12;
  wire f_s_dadda_rca24_and_12_15_b_15;
  wire f_s_dadda_rca24_and_12_15_y0;
  wire f_s_dadda_rca24_and_11_16_a_11;
  wire f_s_dadda_rca24_and_11_16_b_16;
  wire f_s_dadda_rca24_and_11_16_y0;
  wire f_s_dadda_rca24_and_10_17_a_10;
  wire f_s_dadda_rca24_and_10_17_b_17;
  wire f_s_dadda_rca24_and_10_17_y0;
  wire f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_12_15_y0;
  wire f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_11_16_y0;
  wire f_s_dadda_rca24_fa214_y0;
  wire f_s_dadda_rca24_fa214_y1;
  wire f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_10_17_y0;
  wire f_s_dadda_rca24_fa214_y2;
  wire f_s_dadda_rca24_fa214_y3;
  wire f_s_dadda_rca24_fa214_y4;
  wire f_s_dadda_rca24_and_9_18_a_9;
  wire f_s_dadda_rca24_and_9_18_b_18;
  wire f_s_dadda_rca24_and_9_18_y0;
  wire f_s_dadda_rca24_and_8_19_a_8;
  wire f_s_dadda_rca24_and_8_19_b_19;
  wire f_s_dadda_rca24_and_8_19_y0;
  wire f_s_dadda_rca24_and_7_20_a_7;
  wire f_s_dadda_rca24_and_7_20_b_20;
  wire f_s_dadda_rca24_and_7_20_y0;
  wire f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_9_18_y0;
  wire f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_8_19_y0;
  wire f_s_dadda_rca24_fa215_y0;
  wire f_s_dadda_rca24_fa215_y1;
  wire f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_7_20_y0;
  wire f_s_dadda_rca24_fa215_y2;
  wire f_s_dadda_rca24_fa215_y3;
  wire f_s_dadda_rca24_fa215_y4;
  wire f_s_dadda_rca24_and_6_21_a_6;
  wire f_s_dadda_rca24_and_6_21_b_21;
  wire f_s_dadda_rca24_and_6_21_y0;
  wire f_s_dadda_rca24_and_5_22_a_5;
  wire f_s_dadda_rca24_and_5_22_b_22;
  wire f_s_dadda_rca24_and_5_22_y0;
  wire f_s_dadda_rca24_nand_4_23_a_4;
  wire f_s_dadda_rca24_nand_4_23_b_23;
  wire f_s_dadda_rca24_nand_4_23_y0;
  wire f_s_dadda_rca24_fa216_f_s_dadda_rca24_and_6_21_y0;
  wire f_s_dadda_rca24_fa216_f_s_dadda_rca24_and_5_22_y0;
  wire f_s_dadda_rca24_fa216_y0;
  wire f_s_dadda_rca24_fa216_y1;
  wire f_s_dadda_rca24_fa216_f_s_dadda_rca24_nand_4_23_y0;
  wire f_s_dadda_rca24_fa216_y2;
  wire f_s_dadda_rca24_fa216_y3;
  wire f_s_dadda_rca24_fa216_y4;
  wire f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa22_y2;
  wire f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa23_y2;
  wire f_s_dadda_rca24_fa217_y0;
  wire f_s_dadda_rca24_fa217_y1;
  wire f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa207_y2;
  wire f_s_dadda_rca24_fa217_y2;
  wire f_s_dadda_rca24_fa217_y3;
  wire f_s_dadda_rca24_fa217_y4;
  wire f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa208_y2;
  wire f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa209_y2;
  wire f_s_dadda_rca24_fa218_y0;
  wire f_s_dadda_rca24_fa218_y1;
  wire f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa210_y2;
  wire f_s_dadda_rca24_fa218_y2;
  wire f_s_dadda_rca24_fa218_y3;
  wire f_s_dadda_rca24_fa218_y4;
  wire f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa211_y2;
  wire f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa212_y2;
  wire f_s_dadda_rca24_fa219_y0;
  wire f_s_dadda_rca24_fa219_y1;
  wire f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa213_y2;
  wire f_s_dadda_rca24_fa219_y2;
  wire f_s_dadda_rca24_fa219_y3;
  wire f_s_dadda_rca24_fa219_y4;
  wire f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa219_y4;
  wire f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa218_y4;
  wire f_s_dadda_rca24_fa220_y0;
  wire f_s_dadda_rca24_fa220_y1;
  wire f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa217_y4;
  wire f_s_dadda_rca24_fa220_y2;
  wire f_s_dadda_rca24_fa220_y3;
  wire f_s_dadda_rca24_fa220_y4;
  wire f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa216_y4;
  wire f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa215_y4;
  wire f_s_dadda_rca24_fa221_y0;
  wire f_s_dadda_rca24_fa221_y1;
  wire f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa214_y4;
  wire f_s_dadda_rca24_fa221_y2;
  wire f_s_dadda_rca24_fa221_y3;
  wire f_s_dadda_rca24_fa221_y4;
  wire f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa213_y4;
  wire f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa212_y4;
  wire f_s_dadda_rca24_fa222_y0;
  wire f_s_dadda_rca24_fa222_y1;
  wire f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa211_y4;
  wire f_s_dadda_rca24_fa222_y2;
  wire f_s_dadda_rca24_fa222_y3;
  wire f_s_dadda_rca24_fa222_y4;
  wire f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa210_y4;
  wire f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa209_y4;
  wire f_s_dadda_rca24_fa223_y0;
  wire f_s_dadda_rca24_fa223_y1;
  wire f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa208_y4;
  wire f_s_dadda_rca24_fa223_y2;
  wire f_s_dadda_rca24_fa223_y3;
  wire f_s_dadda_rca24_fa223_y4;
  wire f_s_dadda_rca24_and_22_6_a_22;
  wire f_s_dadda_rca24_and_22_6_b_6;
  wire f_s_dadda_rca24_and_22_6_y0;
  wire f_s_dadda_rca24_and_21_7_a_21;
  wire f_s_dadda_rca24_and_21_7_b_7;
  wire f_s_dadda_rca24_and_21_7_y0;
  wire f_s_dadda_rca24_fa224_f_s_dadda_rca24_fa207_y4;
  wire f_s_dadda_rca24_fa224_f_s_dadda_rca24_and_22_6_y0;
  wire f_s_dadda_rca24_fa224_y0;
  wire f_s_dadda_rca24_fa224_y1;
  wire f_s_dadda_rca24_fa224_f_s_dadda_rca24_and_21_7_y0;
  wire f_s_dadda_rca24_fa224_y2;
  wire f_s_dadda_rca24_fa224_y3;
  wire f_s_dadda_rca24_fa224_y4;
  wire f_s_dadda_rca24_and_20_8_a_20;
  wire f_s_dadda_rca24_and_20_8_b_8;
  wire f_s_dadda_rca24_and_20_8_y0;
  wire f_s_dadda_rca24_and_19_9_a_19;
  wire f_s_dadda_rca24_and_19_9_b_9;
  wire f_s_dadda_rca24_and_19_9_y0;
  wire f_s_dadda_rca24_and_18_10_a_18;
  wire f_s_dadda_rca24_and_18_10_b_10;
  wire f_s_dadda_rca24_and_18_10_y0;
  wire f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_20_8_y0;
  wire f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_19_9_y0;
  wire f_s_dadda_rca24_fa225_y0;
  wire f_s_dadda_rca24_fa225_y1;
  wire f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_18_10_y0;
  wire f_s_dadda_rca24_fa225_y2;
  wire f_s_dadda_rca24_fa225_y3;
  wire f_s_dadda_rca24_fa225_y4;
  wire f_s_dadda_rca24_and_17_11_a_17;
  wire f_s_dadda_rca24_and_17_11_b_11;
  wire f_s_dadda_rca24_and_17_11_y0;
  wire f_s_dadda_rca24_and_16_12_a_16;
  wire f_s_dadda_rca24_and_16_12_b_12;
  wire f_s_dadda_rca24_and_16_12_y0;
  wire f_s_dadda_rca24_and_15_13_a_15;
  wire f_s_dadda_rca24_and_15_13_b_13;
  wire f_s_dadda_rca24_and_15_13_y0;
  wire f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_17_11_y0;
  wire f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_16_12_y0;
  wire f_s_dadda_rca24_fa226_y0;
  wire f_s_dadda_rca24_fa226_y1;
  wire f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_15_13_y0;
  wire f_s_dadda_rca24_fa226_y2;
  wire f_s_dadda_rca24_fa226_y3;
  wire f_s_dadda_rca24_fa226_y4;
  wire f_s_dadda_rca24_and_14_14_a_14;
  wire f_s_dadda_rca24_and_14_14_b_14;
  wire f_s_dadda_rca24_and_14_14_y0;
  wire f_s_dadda_rca24_and_13_15_a_13;
  wire f_s_dadda_rca24_and_13_15_b_15;
  wire f_s_dadda_rca24_and_13_15_y0;
  wire f_s_dadda_rca24_and_12_16_a_12;
  wire f_s_dadda_rca24_and_12_16_b_16;
  wire f_s_dadda_rca24_and_12_16_y0;
  wire f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_14_14_y0;
  wire f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_13_15_y0;
  wire f_s_dadda_rca24_fa227_y0;
  wire f_s_dadda_rca24_fa227_y1;
  wire f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_12_16_y0;
  wire f_s_dadda_rca24_fa227_y2;
  wire f_s_dadda_rca24_fa227_y3;
  wire f_s_dadda_rca24_fa227_y4;
  wire f_s_dadda_rca24_and_11_17_a_11;
  wire f_s_dadda_rca24_and_11_17_b_17;
  wire f_s_dadda_rca24_and_11_17_y0;
  wire f_s_dadda_rca24_and_10_18_a_10;
  wire f_s_dadda_rca24_and_10_18_b_18;
  wire f_s_dadda_rca24_and_10_18_y0;
  wire f_s_dadda_rca24_and_9_19_a_9;
  wire f_s_dadda_rca24_and_9_19_b_19;
  wire f_s_dadda_rca24_and_9_19_y0;
  wire f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_11_17_y0;
  wire f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_10_18_y0;
  wire f_s_dadda_rca24_fa228_y0;
  wire f_s_dadda_rca24_fa228_y1;
  wire f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_9_19_y0;
  wire f_s_dadda_rca24_fa228_y2;
  wire f_s_dadda_rca24_fa228_y3;
  wire f_s_dadda_rca24_fa228_y4;
  wire f_s_dadda_rca24_and_8_20_a_8;
  wire f_s_dadda_rca24_and_8_20_b_20;
  wire f_s_dadda_rca24_and_8_20_y0;
  wire f_s_dadda_rca24_and_7_21_a_7;
  wire f_s_dadda_rca24_and_7_21_b_21;
  wire f_s_dadda_rca24_and_7_21_y0;
  wire f_s_dadda_rca24_and_6_22_a_6;
  wire f_s_dadda_rca24_and_6_22_b_22;
  wire f_s_dadda_rca24_and_6_22_y0;
  wire f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_8_20_y0;
  wire f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_7_21_y0;
  wire f_s_dadda_rca24_fa229_y0;
  wire f_s_dadda_rca24_fa229_y1;
  wire f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_6_22_y0;
  wire f_s_dadda_rca24_fa229_y2;
  wire f_s_dadda_rca24_fa229_y3;
  wire f_s_dadda_rca24_fa229_y4;
  wire f_s_dadda_rca24_nand_5_23_a_5;
  wire f_s_dadda_rca24_nand_5_23_b_23;
  wire f_s_dadda_rca24_nand_5_23_y0;
  wire f_s_dadda_rca24_fa230_f_s_dadda_rca24_nand_5_23_y0;
  wire f_s_dadda_rca24_fa230_f_s_dadda_rca24_fa24_y2;
  wire f_s_dadda_rca24_fa230_y0;
  wire f_s_dadda_rca24_fa230_y1;
  wire f_s_dadda_rca24_fa230_f_s_dadda_rca24_fa220_y2;
  wire f_s_dadda_rca24_fa230_y2;
  wire f_s_dadda_rca24_fa230_y3;
  wire f_s_dadda_rca24_fa230_y4;
  wire f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa221_y2;
  wire f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa222_y2;
  wire f_s_dadda_rca24_fa231_y0;
  wire f_s_dadda_rca24_fa231_y1;
  wire f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa223_y2;
  wire f_s_dadda_rca24_fa231_y2;
  wire f_s_dadda_rca24_fa231_y3;
  wire f_s_dadda_rca24_fa231_y4;
  wire f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa224_y2;
  wire f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa225_y2;
  wire f_s_dadda_rca24_fa232_y0;
  wire f_s_dadda_rca24_fa232_y1;
  wire f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa226_y2;
  wire f_s_dadda_rca24_fa232_y2;
  wire f_s_dadda_rca24_fa232_y3;
  wire f_s_dadda_rca24_fa232_y4;
  wire f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa232_y4;
  wire f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa231_y4;
  wire f_s_dadda_rca24_fa233_y0;
  wire f_s_dadda_rca24_fa233_y1;
  wire f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa230_y4;
  wire f_s_dadda_rca24_fa233_y2;
  wire f_s_dadda_rca24_fa233_y3;
  wire f_s_dadda_rca24_fa233_y4;
  wire f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa229_y4;
  wire f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa228_y4;
  wire f_s_dadda_rca24_fa234_y0;
  wire f_s_dadda_rca24_fa234_y1;
  wire f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa227_y4;
  wire f_s_dadda_rca24_fa234_y2;
  wire f_s_dadda_rca24_fa234_y3;
  wire f_s_dadda_rca24_fa234_y4;
  wire f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa226_y4;
  wire f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa225_y4;
  wire f_s_dadda_rca24_fa235_y0;
  wire f_s_dadda_rca24_fa235_y1;
  wire f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa224_y4;
  wire f_s_dadda_rca24_fa235_y2;
  wire f_s_dadda_rca24_fa235_y3;
  wire f_s_dadda_rca24_fa235_y4;
  wire f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa223_y4;
  wire f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa222_y4;
  wire f_s_dadda_rca24_fa236_y0;
  wire f_s_dadda_rca24_fa236_y1;
  wire f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa221_y4;
  wire f_s_dadda_rca24_fa236_y2;
  wire f_s_dadda_rca24_fa236_y3;
  wire f_s_dadda_rca24_fa236_y4;
  wire f_s_dadda_rca24_nand_23_6_a_23;
  wire f_s_dadda_rca24_nand_23_6_b_6;
  wire f_s_dadda_rca24_nand_23_6_y0;
  wire f_s_dadda_rca24_fa237_f_s_dadda_rca24_fa220_y4;
  wire f_s_dadda_rca24_fa237_f_s_dadda_rca24_fa24_y4;
  wire f_s_dadda_rca24_fa237_y0;
  wire f_s_dadda_rca24_fa237_y1;
  wire f_s_dadda_rca24_fa237_f_s_dadda_rca24_nand_23_6_y0;
  wire f_s_dadda_rca24_fa237_y2;
  wire f_s_dadda_rca24_fa237_y3;
  wire f_s_dadda_rca24_fa237_y4;
  wire f_s_dadda_rca24_and_22_7_a_22;
  wire f_s_dadda_rca24_and_22_7_b_7;
  wire f_s_dadda_rca24_and_22_7_y0;
  wire f_s_dadda_rca24_and_21_8_a_21;
  wire f_s_dadda_rca24_and_21_8_b_8;
  wire f_s_dadda_rca24_and_21_8_y0;
  wire f_s_dadda_rca24_and_20_9_a_20;
  wire f_s_dadda_rca24_and_20_9_b_9;
  wire f_s_dadda_rca24_and_20_9_y0;
  wire f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_22_7_y0;
  wire f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_21_8_y0;
  wire f_s_dadda_rca24_fa238_y0;
  wire f_s_dadda_rca24_fa238_y1;
  wire f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_20_9_y0;
  wire f_s_dadda_rca24_fa238_y2;
  wire f_s_dadda_rca24_fa238_y3;
  wire f_s_dadda_rca24_fa238_y4;
  wire f_s_dadda_rca24_and_19_10_a_19;
  wire f_s_dadda_rca24_and_19_10_b_10;
  wire f_s_dadda_rca24_and_19_10_y0;
  wire f_s_dadda_rca24_and_18_11_a_18;
  wire f_s_dadda_rca24_and_18_11_b_11;
  wire f_s_dadda_rca24_and_18_11_y0;
  wire f_s_dadda_rca24_and_17_12_a_17;
  wire f_s_dadda_rca24_and_17_12_b_12;
  wire f_s_dadda_rca24_and_17_12_y0;
  wire f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_19_10_y0;
  wire f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_18_11_y0;
  wire f_s_dadda_rca24_fa239_y0;
  wire f_s_dadda_rca24_fa239_y1;
  wire f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_17_12_y0;
  wire f_s_dadda_rca24_fa239_y2;
  wire f_s_dadda_rca24_fa239_y3;
  wire f_s_dadda_rca24_fa239_y4;
  wire f_s_dadda_rca24_and_16_13_a_16;
  wire f_s_dadda_rca24_and_16_13_b_13;
  wire f_s_dadda_rca24_and_16_13_y0;
  wire f_s_dadda_rca24_and_15_14_a_15;
  wire f_s_dadda_rca24_and_15_14_b_14;
  wire f_s_dadda_rca24_and_15_14_y0;
  wire f_s_dadda_rca24_and_14_15_a_14;
  wire f_s_dadda_rca24_and_14_15_b_15;
  wire f_s_dadda_rca24_and_14_15_y0;
  wire f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_16_13_y0;
  wire f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_15_14_y0;
  wire f_s_dadda_rca24_fa240_y0;
  wire f_s_dadda_rca24_fa240_y1;
  wire f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_14_15_y0;
  wire f_s_dadda_rca24_fa240_y2;
  wire f_s_dadda_rca24_fa240_y3;
  wire f_s_dadda_rca24_fa240_y4;
  wire f_s_dadda_rca24_and_13_16_a_13;
  wire f_s_dadda_rca24_and_13_16_b_16;
  wire f_s_dadda_rca24_and_13_16_y0;
  wire f_s_dadda_rca24_and_12_17_a_12;
  wire f_s_dadda_rca24_and_12_17_b_17;
  wire f_s_dadda_rca24_and_12_17_y0;
  wire f_s_dadda_rca24_and_11_18_a_11;
  wire f_s_dadda_rca24_and_11_18_b_18;
  wire f_s_dadda_rca24_and_11_18_y0;
  wire f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_13_16_y0;
  wire f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_12_17_y0;
  wire f_s_dadda_rca24_fa241_y0;
  wire f_s_dadda_rca24_fa241_y1;
  wire f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_11_18_y0;
  wire f_s_dadda_rca24_fa241_y2;
  wire f_s_dadda_rca24_fa241_y3;
  wire f_s_dadda_rca24_fa241_y4;
  wire f_s_dadda_rca24_and_10_19_a_10;
  wire f_s_dadda_rca24_and_10_19_b_19;
  wire f_s_dadda_rca24_and_10_19_y0;
  wire f_s_dadda_rca24_and_9_20_a_9;
  wire f_s_dadda_rca24_and_9_20_b_20;
  wire f_s_dadda_rca24_and_9_20_y0;
  wire f_s_dadda_rca24_and_8_21_a_8;
  wire f_s_dadda_rca24_and_8_21_b_21;
  wire f_s_dadda_rca24_and_8_21_y0;
  wire f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_10_19_y0;
  wire f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_9_20_y0;
  wire f_s_dadda_rca24_fa242_y0;
  wire f_s_dadda_rca24_fa242_y1;
  wire f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_8_21_y0;
  wire f_s_dadda_rca24_fa242_y2;
  wire f_s_dadda_rca24_fa242_y3;
  wire f_s_dadda_rca24_fa242_y4;
  wire f_s_dadda_rca24_and_7_22_a_7;
  wire f_s_dadda_rca24_and_7_22_b_22;
  wire f_s_dadda_rca24_and_7_22_y0;
  wire f_s_dadda_rca24_nand_6_23_a_6;
  wire f_s_dadda_rca24_nand_6_23_b_23;
  wire f_s_dadda_rca24_nand_6_23_y0;
  wire f_s_dadda_rca24_fa243_f_s_dadda_rca24_and_7_22_y0;
  wire f_s_dadda_rca24_fa243_f_s_dadda_rca24_nand_6_23_y0;
  wire f_s_dadda_rca24_fa243_y0;
  wire f_s_dadda_rca24_fa243_y1;
  wire f_s_dadda_rca24_fa243_f_s_dadda_rca24_fa233_y2;
  wire f_s_dadda_rca24_fa243_y2;
  wire f_s_dadda_rca24_fa243_y3;
  wire f_s_dadda_rca24_fa243_y4;
  wire f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa234_y2;
  wire f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa235_y2;
  wire f_s_dadda_rca24_fa244_y0;
  wire f_s_dadda_rca24_fa244_y1;
  wire f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa236_y2;
  wire f_s_dadda_rca24_fa244_y2;
  wire f_s_dadda_rca24_fa244_y3;
  wire f_s_dadda_rca24_fa244_y4;
  wire f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa237_y2;
  wire f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa238_y2;
  wire f_s_dadda_rca24_fa245_y0;
  wire f_s_dadda_rca24_fa245_y1;
  wire f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa239_y2;
  wire f_s_dadda_rca24_fa245_y2;
  wire f_s_dadda_rca24_fa245_y3;
  wire f_s_dadda_rca24_fa245_y4;
  wire f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa245_y4;
  wire f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa244_y4;
  wire f_s_dadda_rca24_fa246_y0;
  wire f_s_dadda_rca24_fa246_y1;
  wire f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa243_y4;
  wire f_s_dadda_rca24_fa246_y2;
  wire f_s_dadda_rca24_fa246_y3;
  wire f_s_dadda_rca24_fa246_y4;
  wire f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa242_y4;
  wire f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa241_y4;
  wire f_s_dadda_rca24_fa247_y0;
  wire f_s_dadda_rca24_fa247_y1;
  wire f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa240_y4;
  wire f_s_dadda_rca24_fa247_y2;
  wire f_s_dadda_rca24_fa247_y3;
  wire f_s_dadda_rca24_fa247_y4;
  wire f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa239_y4;
  wire f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa238_y4;
  wire f_s_dadda_rca24_fa248_y0;
  wire f_s_dadda_rca24_fa248_y1;
  wire f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa237_y4;
  wire f_s_dadda_rca24_fa248_y2;
  wire f_s_dadda_rca24_fa248_y3;
  wire f_s_dadda_rca24_fa248_y4;
  wire f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa236_y4;
  wire f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa235_y4;
  wire f_s_dadda_rca24_fa249_y0;
  wire f_s_dadda_rca24_fa249_y1;
  wire f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa234_y4;
  wire f_s_dadda_rca24_fa249_y2;
  wire f_s_dadda_rca24_fa249_y3;
  wire f_s_dadda_rca24_fa249_y4;
  wire f_s_dadda_rca24_nand_23_7_a_23;
  wire f_s_dadda_rca24_nand_23_7_b_7;
  wire f_s_dadda_rca24_nand_23_7_y0;
  wire f_s_dadda_rca24_and_22_8_a_22;
  wire f_s_dadda_rca24_and_22_8_b_8;
  wire f_s_dadda_rca24_and_22_8_y0;
  wire f_s_dadda_rca24_fa250_f_s_dadda_rca24_fa233_y4;
  wire f_s_dadda_rca24_fa250_f_s_dadda_rca24_nand_23_7_y0;
  wire f_s_dadda_rca24_fa250_y0;
  wire f_s_dadda_rca24_fa250_y1;
  wire f_s_dadda_rca24_fa250_f_s_dadda_rca24_and_22_8_y0;
  wire f_s_dadda_rca24_fa250_y2;
  wire f_s_dadda_rca24_fa250_y3;
  wire f_s_dadda_rca24_fa250_y4;
  wire f_s_dadda_rca24_and_21_9_a_21;
  wire f_s_dadda_rca24_and_21_9_b_9;
  wire f_s_dadda_rca24_and_21_9_y0;
  wire f_s_dadda_rca24_and_20_10_a_20;
  wire f_s_dadda_rca24_and_20_10_b_10;
  wire f_s_dadda_rca24_and_20_10_y0;
  wire f_s_dadda_rca24_and_19_11_a_19;
  wire f_s_dadda_rca24_and_19_11_b_11;
  wire f_s_dadda_rca24_and_19_11_y0;
  wire f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_21_9_y0;
  wire f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_20_10_y0;
  wire f_s_dadda_rca24_fa251_y0;
  wire f_s_dadda_rca24_fa251_y1;
  wire f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_19_11_y0;
  wire f_s_dadda_rca24_fa251_y2;
  wire f_s_dadda_rca24_fa251_y3;
  wire f_s_dadda_rca24_fa251_y4;
  wire f_s_dadda_rca24_and_18_12_a_18;
  wire f_s_dadda_rca24_and_18_12_b_12;
  wire f_s_dadda_rca24_and_18_12_y0;
  wire f_s_dadda_rca24_and_17_13_a_17;
  wire f_s_dadda_rca24_and_17_13_b_13;
  wire f_s_dadda_rca24_and_17_13_y0;
  wire f_s_dadda_rca24_and_16_14_a_16;
  wire f_s_dadda_rca24_and_16_14_b_14;
  wire f_s_dadda_rca24_and_16_14_y0;
  wire f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_18_12_y0;
  wire f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_17_13_y0;
  wire f_s_dadda_rca24_fa252_y0;
  wire f_s_dadda_rca24_fa252_y1;
  wire f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_16_14_y0;
  wire f_s_dadda_rca24_fa252_y2;
  wire f_s_dadda_rca24_fa252_y3;
  wire f_s_dadda_rca24_fa252_y4;
  wire f_s_dadda_rca24_and_15_15_a_15;
  wire f_s_dadda_rca24_and_15_15_b_15;
  wire f_s_dadda_rca24_and_15_15_y0;
  wire f_s_dadda_rca24_and_14_16_a_14;
  wire f_s_dadda_rca24_and_14_16_b_16;
  wire f_s_dadda_rca24_and_14_16_y0;
  wire f_s_dadda_rca24_and_13_17_a_13;
  wire f_s_dadda_rca24_and_13_17_b_17;
  wire f_s_dadda_rca24_and_13_17_y0;
  wire f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_15_15_y0;
  wire f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_14_16_y0;
  wire f_s_dadda_rca24_fa253_y0;
  wire f_s_dadda_rca24_fa253_y1;
  wire f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_13_17_y0;
  wire f_s_dadda_rca24_fa253_y2;
  wire f_s_dadda_rca24_fa253_y3;
  wire f_s_dadda_rca24_fa253_y4;
  wire f_s_dadda_rca24_and_12_18_a_12;
  wire f_s_dadda_rca24_and_12_18_b_18;
  wire f_s_dadda_rca24_and_12_18_y0;
  wire f_s_dadda_rca24_and_11_19_a_11;
  wire f_s_dadda_rca24_and_11_19_b_19;
  wire f_s_dadda_rca24_and_11_19_y0;
  wire f_s_dadda_rca24_and_10_20_a_10;
  wire f_s_dadda_rca24_and_10_20_b_20;
  wire f_s_dadda_rca24_and_10_20_y0;
  wire f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_12_18_y0;
  wire f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_11_19_y0;
  wire f_s_dadda_rca24_fa254_y0;
  wire f_s_dadda_rca24_fa254_y1;
  wire f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_10_20_y0;
  wire f_s_dadda_rca24_fa254_y2;
  wire f_s_dadda_rca24_fa254_y3;
  wire f_s_dadda_rca24_fa254_y4;
  wire f_s_dadda_rca24_and_9_21_a_9;
  wire f_s_dadda_rca24_and_9_21_b_21;
  wire f_s_dadda_rca24_and_9_21_y0;
  wire f_s_dadda_rca24_and_8_22_a_8;
  wire f_s_dadda_rca24_and_8_22_b_22;
  wire f_s_dadda_rca24_and_8_22_y0;
  wire f_s_dadda_rca24_nand_7_23_a_7;
  wire f_s_dadda_rca24_nand_7_23_b_23;
  wire f_s_dadda_rca24_nand_7_23_y0;
  wire f_s_dadda_rca24_fa255_f_s_dadda_rca24_and_9_21_y0;
  wire f_s_dadda_rca24_fa255_f_s_dadda_rca24_and_8_22_y0;
  wire f_s_dadda_rca24_fa255_y0;
  wire f_s_dadda_rca24_fa255_y1;
  wire f_s_dadda_rca24_fa255_f_s_dadda_rca24_nand_7_23_y0;
  wire f_s_dadda_rca24_fa255_y2;
  wire f_s_dadda_rca24_fa255_y3;
  wire f_s_dadda_rca24_fa255_y4;
  wire f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa246_y2;
  wire f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa247_y2;
  wire f_s_dadda_rca24_fa256_y0;
  wire f_s_dadda_rca24_fa256_y1;
  wire f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa248_y2;
  wire f_s_dadda_rca24_fa256_y2;
  wire f_s_dadda_rca24_fa256_y3;
  wire f_s_dadda_rca24_fa256_y4;
  wire f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa249_y2;
  wire f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa250_y2;
  wire f_s_dadda_rca24_fa257_y0;
  wire f_s_dadda_rca24_fa257_y1;
  wire f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa251_y2;
  wire f_s_dadda_rca24_fa257_y2;
  wire f_s_dadda_rca24_fa257_y3;
  wire f_s_dadda_rca24_fa257_y4;
  wire f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa257_y4;
  wire f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa256_y4;
  wire f_s_dadda_rca24_fa258_y0;
  wire f_s_dadda_rca24_fa258_y1;
  wire f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa255_y4;
  wire f_s_dadda_rca24_fa258_y2;
  wire f_s_dadda_rca24_fa258_y3;
  wire f_s_dadda_rca24_fa258_y4;
  wire f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa254_y4;
  wire f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa253_y4;
  wire f_s_dadda_rca24_fa259_y0;
  wire f_s_dadda_rca24_fa259_y1;
  wire f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa252_y4;
  wire f_s_dadda_rca24_fa259_y2;
  wire f_s_dadda_rca24_fa259_y3;
  wire f_s_dadda_rca24_fa259_y4;
  wire f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa251_y4;
  wire f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa250_y4;
  wire f_s_dadda_rca24_fa260_y0;
  wire f_s_dadda_rca24_fa260_y1;
  wire f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa249_y4;
  wire f_s_dadda_rca24_fa260_y2;
  wire f_s_dadda_rca24_fa260_y3;
  wire f_s_dadda_rca24_fa260_y4;
  wire f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa248_y4;
  wire f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa247_y4;
  wire f_s_dadda_rca24_fa261_y0;
  wire f_s_dadda_rca24_fa261_y1;
  wire f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa246_y4;
  wire f_s_dadda_rca24_fa261_y2;
  wire f_s_dadda_rca24_fa261_y3;
  wire f_s_dadda_rca24_fa261_y4;
  wire f_s_dadda_rca24_nand_23_8_a_23;
  wire f_s_dadda_rca24_nand_23_8_b_8;
  wire f_s_dadda_rca24_nand_23_8_y0;
  wire f_s_dadda_rca24_and_22_9_a_22;
  wire f_s_dadda_rca24_and_22_9_b_9;
  wire f_s_dadda_rca24_and_22_9_y0;
  wire f_s_dadda_rca24_and_21_10_a_21;
  wire f_s_dadda_rca24_and_21_10_b_10;
  wire f_s_dadda_rca24_and_21_10_y0;
  wire f_s_dadda_rca24_fa262_f_s_dadda_rca24_nand_23_8_y0;
  wire f_s_dadda_rca24_fa262_f_s_dadda_rca24_and_22_9_y0;
  wire f_s_dadda_rca24_fa262_y0;
  wire f_s_dadda_rca24_fa262_y1;
  wire f_s_dadda_rca24_fa262_f_s_dadda_rca24_and_21_10_y0;
  wire f_s_dadda_rca24_fa262_y2;
  wire f_s_dadda_rca24_fa262_y3;
  wire f_s_dadda_rca24_fa262_y4;
  wire f_s_dadda_rca24_and_20_11_a_20;
  wire f_s_dadda_rca24_and_20_11_b_11;
  wire f_s_dadda_rca24_and_20_11_y0;
  wire f_s_dadda_rca24_and_19_12_a_19;
  wire f_s_dadda_rca24_and_19_12_b_12;
  wire f_s_dadda_rca24_and_19_12_y0;
  wire f_s_dadda_rca24_and_18_13_a_18;
  wire f_s_dadda_rca24_and_18_13_b_13;
  wire f_s_dadda_rca24_and_18_13_y0;
  wire f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_20_11_y0;
  wire f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_19_12_y0;
  wire f_s_dadda_rca24_fa263_y0;
  wire f_s_dadda_rca24_fa263_y1;
  wire f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_18_13_y0;
  wire f_s_dadda_rca24_fa263_y2;
  wire f_s_dadda_rca24_fa263_y3;
  wire f_s_dadda_rca24_fa263_y4;
  wire f_s_dadda_rca24_and_17_14_a_17;
  wire f_s_dadda_rca24_and_17_14_b_14;
  wire f_s_dadda_rca24_and_17_14_y0;
  wire f_s_dadda_rca24_and_16_15_a_16;
  wire f_s_dadda_rca24_and_16_15_b_15;
  wire f_s_dadda_rca24_and_16_15_y0;
  wire f_s_dadda_rca24_and_15_16_a_15;
  wire f_s_dadda_rca24_and_15_16_b_16;
  wire f_s_dadda_rca24_and_15_16_y0;
  wire f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_17_14_y0;
  wire f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_16_15_y0;
  wire f_s_dadda_rca24_fa264_y0;
  wire f_s_dadda_rca24_fa264_y1;
  wire f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_15_16_y0;
  wire f_s_dadda_rca24_fa264_y2;
  wire f_s_dadda_rca24_fa264_y3;
  wire f_s_dadda_rca24_fa264_y4;
  wire f_s_dadda_rca24_and_14_17_a_14;
  wire f_s_dadda_rca24_and_14_17_b_17;
  wire f_s_dadda_rca24_and_14_17_y0;
  wire f_s_dadda_rca24_and_13_18_a_13;
  wire f_s_dadda_rca24_and_13_18_b_18;
  wire f_s_dadda_rca24_and_13_18_y0;
  wire f_s_dadda_rca24_and_12_19_a_12;
  wire f_s_dadda_rca24_and_12_19_b_19;
  wire f_s_dadda_rca24_and_12_19_y0;
  wire f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_14_17_y0;
  wire f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_13_18_y0;
  wire f_s_dadda_rca24_fa265_y0;
  wire f_s_dadda_rca24_fa265_y1;
  wire f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_12_19_y0;
  wire f_s_dadda_rca24_fa265_y2;
  wire f_s_dadda_rca24_fa265_y3;
  wire f_s_dadda_rca24_fa265_y4;
  wire f_s_dadda_rca24_and_11_20_a_11;
  wire f_s_dadda_rca24_and_11_20_b_20;
  wire f_s_dadda_rca24_and_11_20_y0;
  wire f_s_dadda_rca24_and_10_21_a_10;
  wire f_s_dadda_rca24_and_10_21_b_21;
  wire f_s_dadda_rca24_and_10_21_y0;
  wire f_s_dadda_rca24_and_9_22_a_9;
  wire f_s_dadda_rca24_and_9_22_b_22;
  wire f_s_dadda_rca24_and_9_22_y0;
  wire f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_11_20_y0;
  wire f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_10_21_y0;
  wire f_s_dadda_rca24_fa266_y0;
  wire f_s_dadda_rca24_fa266_y1;
  wire f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_9_22_y0;
  wire f_s_dadda_rca24_fa266_y2;
  wire f_s_dadda_rca24_fa266_y3;
  wire f_s_dadda_rca24_fa266_y4;
  wire f_s_dadda_rca24_nand_8_23_a_8;
  wire f_s_dadda_rca24_nand_8_23_b_23;
  wire f_s_dadda_rca24_nand_8_23_y0;
  wire f_s_dadda_rca24_fa267_f_s_dadda_rca24_nand_8_23_y0;
  wire f_s_dadda_rca24_fa267_f_s_dadda_rca24_fa258_y2;
  wire f_s_dadda_rca24_fa267_y0;
  wire f_s_dadda_rca24_fa267_y1;
  wire f_s_dadda_rca24_fa267_f_s_dadda_rca24_fa259_y2;
  wire f_s_dadda_rca24_fa267_y2;
  wire f_s_dadda_rca24_fa267_y3;
  wire f_s_dadda_rca24_fa267_y4;
  wire f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa260_y2;
  wire f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa261_y2;
  wire f_s_dadda_rca24_fa268_y0;
  wire f_s_dadda_rca24_fa268_y1;
  wire f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa262_y2;
  wire f_s_dadda_rca24_fa268_y2;
  wire f_s_dadda_rca24_fa268_y3;
  wire f_s_dadda_rca24_fa268_y4;
  wire f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa268_y4;
  wire f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa267_y4;
  wire f_s_dadda_rca24_fa269_y0;
  wire f_s_dadda_rca24_fa269_y1;
  wire f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa266_y4;
  wire f_s_dadda_rca24_fa269_y2;
  wire f_s_dadda_rca24_fa269_y3;
  wire f_s_dadda_rca24_fa269_y4;
  wire f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa265_y4;
  wire f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa264_y4;
  wire f_s_dadda_rca24_fa270_y0;
  wire f_s_dadda_rca24_fa270_y1;
  wire f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa263_y4;
  wire f_s_dadda_rca24_fa270_y2;
  wire f_s_dadda_rca24_fa270_y3;
  wire f_s_dadda_rca24_fa270_y4;
  wire f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa262_y4;
  wire f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa261_y4;
  wire f_s_dadda_rca24_fa271_y0;
  wire f_s_dadda_rca24_fa271_y1;
  wire f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa260_y4;
  wire f_s_dadda_rca24_fa271_y2;
  wire f_s_dadda_rca24_fa271_y3;
  wire f_s_dadda_rca24_fa271_y4;
  wire f_s_dadda_rca24_nand_23_9_a_23;
  wire f_s_dadda_rca24_nand_23_9_b_9;
  wire f_s_dadda_rca24_nand_23_9_y0;
  wire f_s_dadda_rca24_fa272_f_s_dadda_rca24_fa259_y4;
  wire f_s_dadda_rca24_fa272_f_s_dadda_rca24_fa258_y4;
  wire f_s_dadda_rca24_fa272_y0;
  wire f_s_dadda_rca24_fa272_y1;
  wire f_s_dadda_rca24_fa272_f_s_dadda_rca24_nand_23_9_y0;
  wire f_s_dadda_rca24_fa272_y2;
  wire f_s_dadda_rca24_fa272_y3;
  wire f_s_dadda_rca24_fa272_y4;
  wire f_s_dadda_rca24_and_22_10_a_22;
  wire f_s_dadda_rca24_and_22_10_b_10;
  wire f_s_dadda_rca24_and_22_10_y0;
  wire f_s_dadda_rca24_and_21_11_a_21;
  wire f_s_dadda_rca24_and_21_11_b_11;
  wire f_s_dadda_rca24_and_21_11_y0;
  wire f_s_dadda_rca24_and_20_12_a_20;
  wire f_s_dadda_rca24_and_20_12_b_12;
  wire f_s_dadda_rca24_and_20_12_y0;
  wire f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_22_10_y0;
  wire f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_21_11_y0;
  wire f_s_dadda_rca24_fa273_y0;
  wire f_s_dadda_rca24_fa273_y1;
  wire f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_20_12_y0;
  wire f_s_dadda_rca24_fa273_y2;
  wire f_s_dadda_rca24_fa273_y3;
  wire f_s_dadda_rca24_fa273_y4;
  wire f_s_dadda_rca24_and_19_13_a_19;
  wire f_s_dadda_rca24_and_19_13_b_13;
  wire f_s_dadda_rca24_and_19_13_y0;
  wire f_s_dadda_rca24_and_18_14_a_18;
  wire f_s_dadda_rca24_and_18_14_b_14;
  wire f_s_dadda_rca24_and_18_14_y0;
  wire f_s_dadda_rca24_and_17_15_a_17;
  wire f_s_dadda_rca24_and_17_15_b_15;
  wire f_s_dadda_rca24_and_17_15_y0;
  wire f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_19_13_y0;
  wire f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_18_14_y0;
  wire f_s_dadda_rca24_fa274_y0;
  wire f_s_dadda_rca24_fa274_y1;
  wire f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_17_15_y0;
  wire f_s_dadda_rca24_fa274_y2;
  wire f_s_dadda_rca24_fa274_y3;
  wire f_s_dadda_rca24_fa274_y4;
  wire f_s_dadda_rca24_and_16_16_a_16;
  wire f_s_dadda_rca24_and_16_16_b_16;
  wire f_s_dadda_rca24_and_16_16_y0;
  wire f_s_dadda_rca24_and_15_17_a_15;
  wire f_s_dadda_rca24_and_15_17_b_17;
  wire f_s_dadda_rca24_and_15_17_y0;
  wire f_s_dadda_rca24_and_14_18_a_14;
  wire f_s_dadda_rca24_and_14_18_b_18;
  wire f_s_dadda_rca24_and_14_18_y0;
  wire f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_16_16_y0;
  wire f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_15_17_y0;
  wire f_s_dadda_rca24_fa275_y0;
  wire f_s_dadda_rca24_fa275_y1;
  wire f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_14_18_y0;
  wire f_s_dadda_rca24_fa275_y2;
  wire f_s_dadda_rca24_fa275_y3;
  wire f_s_dadda_rca24_fa275_y4;
  wire f_s_dadda_rca24_and_13_19_a_13;
  wire f_s_dadda_rca24_and_13_19_b_19;
  wire f_s_dadda_rca24_and_13_19_y0;
  wire f_s_dadda_rca24_and_12_20_a_12;
  wire f_s_dadda_rca24_and_12_20_b_20;
  wire f_s_dadda_rca24_and_12_20_y0;
  wire f_s_dadda_rca24_and_11_21_a_11;
  wire f_s_dadda_rca24_and_11_21_b_21;
  wire f_s_dadda_rca24_and_11_21_y0;
  wire f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_13_19_y0;
  wire f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_12_20_y0;
  wire f_s_dadda_rca24_fa276_y0;
  wire f_s_dadda_rca24_fa276_y1;
  wire f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_11_21_y0;
  wire f_s_dadda_rca24_fa276_y2;
  wire f_s_dadda_rca24_fa276_y3;
  wire f_s_dadda_rca24_fa276_y4;
  wire f_s_dadda_rca24_and_10_22_a_10;
  wire f_s_dadda_rca24_and_10_22_b_22;
  wire f_s_dadda_rca24_and_10_22_y0;
  wire f_s_dadda_rca24_nand_9_23_a_9;
  wire f_s_dadda_rca24_nand_9_23_b_23;
  wire f_s_dadda_rca24_nand_9_23_y0;
  wire f_s_dadda_rca24_fa277_f_s_dadda_rca24_and_10_22_y0;
  wire f_s_dadda_rca24_fa277_f_s_dadda_rca24_nand_9_23_y0;
  wire f_s_dadda_rca24_fa277_y0;
  wire f_s_dadda_rca24_fa277_y1;
  wire f_s_dadda_rca24_fa277_f_s_dadda_rca24_fa269_y2;
  wire f_s_dadda_rca24_fa277_y2;
  wire f_s_dadda_rca24_fa277_y3;
  wire f_s_dadda_rca24_fa277_y4;
  wire f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa270_y2;
  wire f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa271_y2;
  wire f_s_dadda_rca24_fa278_y0;
  wire f_s_dadda_rca24_fa278_y1;
  wire f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa272_y2;
  wire f_s_dadda_rca24_fa278_y2;
  wire f_s_dadda_rca24_fa278_y3;
  wire f_s_dadda_rca24_fa278_y4;
  wire f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa278_y4;
  wire f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa277_y4;
  wire f_s_dadda_rca24_fa279_y0;
  wire f_s_dadda_rca24_fa279_y1;
  wire f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa276_y4;
  wire f_s_dadda_rca24_fa279_y2;
  wire f_s_dadda_rca24_fa279_y3;
  wire f_s_dadda_rca24_fa279_y4;
  wire f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa275_y4;
  wire f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa274_y4;
  wire f_s_dadda_rca24_fa280_y0;
  wire f_s_dadda_rca24_fa280_y1;
  wire f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa273_y4;
  wire f_s_dadda_rca24_fa280_y2;
  wire f_s_dadda_rca24_fa280_y3;
  wire f_s_dadda_rca24_fa280_y4;
  wire f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa272_y4;
  wire f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa271_y4;
  wire f_s_dadda_rca24_fa281_y0;
  wire f_s_dadda_rca24_fa281_y1;
  wire f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa270_y4;
  wire f_s_dadda_rca24_fa281_y2;
  wire f_s_dadda_rca24_fa281_y3;
  wire f_s_dadda_rca24_fa281_y4;
  wire f_s_dadda_rca24_nand_23_10_a_23;
  wire f_s_dadda_rca24_nand_23_10_b_10;
  wire f_s_dadda_rca24_nand_23_10_y0;
  wire f_s_dadda_rca24_and_22_11_a_22;
  wire f_s_dadda_rca24_and_22_11_b_11;
  wire f_s_dadda_rca24_and_22_11_y0;
  wire f_s_dadda_rca24_fa282_f_s_dadda_rca24_fa269_y4;
  wire f_s_dadda_rca24_fa282_f_s_dadda_rca24_nand_23_10_y0;
  wire f_s_dadda_rca24_fa282_y0;
  wire f_s_dadda_rca24_fa282_y1;
  wire f_s_dadda_rca24_fa282_f_s_dadda_rca24_and_22_11_y0;
  wire f_s_dadda_rca24_fa282_y2;
  wire f_s_dadda_rca24_fa282_y3;
  wire f_s_dadda_rca24_fa282_y4;
  wire f_s_dadda_rca24_and_21_12_a_21;
  wire f_s_dadda_rca24_and_21_12_b_12;
  wire f_s_dadda_rca24_and_21_12_y0;
  wire f_s_dadda_rca24_and_20_13_a_20;
  wire f_s_dadda_rca24_and_20_13_b_13;
  wire f_s_dadda_rca24_and_20_13_y0;
  wire f_s_dadda_rca24_and_19_14_a_19;
  wire f_s_dadda_rca24_and_19_14_b_14;
  wire f_s_dadda_rca24_and_19_14_y0;
  wire f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_21_12_y0;
  wire f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_20_13_y0;
  wire f_s_dadda_rca24_fa283_y0;
  wire f_s_dadda_rca24_fa283_y1;
  wire f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_19_14_y0;
  wire f_s_dadda_rca24_fa283_y2;
  wire f_s_dadda_rca24_fa283_y3;
  wire f_s_dadda_rca24_fa283_y4;
  wire f_s_dadda_rca24_and_18_15_a_18;
  wire f_s_dadda_rca24_and_18_15_b_15;
  wire f_s_dadda_rca24_and_18_15_y0;
  wire f_s_dadda_rca24_and_17_16_a_17;
  wire f_s_dadda_rca24_and_17_16_b_16;
  wire f_s_dadda_rca24_and_17_16_y0;
  wire f_s_dadda_rca24_and_16_17_a_16;
  wire f_s_dadda_rca24_and_16_17_b_17;
  wire f_s_dadda_rca24_and_16_17_y0;
  wire f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_18_15_y0;
  wire f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_17_16_y0;
  wire f_s_dadda_rca24_fa284_y0;
  wire f_s_dadda_rca24_fa284_y1;
  wire f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_16_17_y0;
  wire f_s_dadda_rca24_fa284_y2;
  wire f_s_dadda_rca24_fa284_y3;
  wire f_s_dadda_rca24_fa284_y4;
  wire f_s_dadda_rca24_and_15_18_a_15;
  wire f_s_dadda_rca24_and_15_18_b_18;
  wire f_s_dadda_rca24_and_15_18_y0;
  wire f_s_dadda_rca24_and_14_19_a_14;
  wire f_s_dadda_rca24_and_14_19_b_19;
  wire f_s_dadda_rca24_and_14_19_y0;
  wire f_s_dadda_rca24_and_13_20_a_13;
  wire f_s_dadda_rca24_and_13_20_b_20;
  wire f_s_dadda_rca24_and_13_20_y0;
  wire f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_15_18_y0;
  wire f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_14_19_y0;
  wire f_s_dadda_rca24_fa285_y0;
  wire f_s_dadda_rca24_fa285_y1;
  wire f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_13_20_y0;
  wire f_s_dadda_rca24_fa285_y2;
  wire f_s_dadda_rca24_fa285_y3;
  wire f_s_dadda_rca24_fa285_y4;
  wire f_s_dadda_rca24_and_12_21_a_12;
  wire f_s_dadda_rca24_and_12_21_b_21;
  wire f_s_dadda_rca24_and_12_21_y0;
  wire f_s_dadda_rca24_and_11_22_a_11;
  wire f_s_dadda_rca24_and_11_22_b_22;
  wire f_s_dadda_rca24_and_11_22_y0;
  wire f_s_dadda_rca24_nand_10_23_a_10;
  wire f_s_dadda_rca24_nand_10_23_b_23;
  wire f_s_dadda_rca24_nand_10_23_y0;
  wire f_s_dadda_rca24_fa286_f_s_dadda_rca24_and_12_21_y0;
  wire f_s_dadda_rca24_fa286_f_s_dadda_rca24_and_11_22_y0;
  wire f_s_dadda_rca24_fa286_y0;
  wire f_s_dadda_rca24_fa286_y1;
  wire f_s_dadda_rca24_fa286_f_s_dadda_rca24_nand_10_23_y0;
  wire f_s_dadda_rca24_fa286_y2;
  wire f_s_dadda_rca24_fa286_y3;
  wire f_s_dadda_rca24_fa286_y4;
  wire f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa279_y2;
  wire f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa280_y2;
  wire f_s_dadda_rca24_fa287_y0;
  wire f_s_dadda_rca24_fa287_y1;
  wire f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa281_y2;
  wire f_s_dadda_rca24_fa287_y2;
  wire f_s_dadda_rca24_fa287_y3;
  wire f_s_dadda_rca24_fa287_y4;
  wire f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa287_y4;
  wire f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa286_y4;
  wire f_s_dadda_rca24_fa288_y0;
  wire f_s_dadda_rca24_fa288_y1;
  wire f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa285_y4;
  wire f_s_dadda_rca24_fa288_y2;
  wire f_s_dadda_rca24_fa288_y3;
  wire f_s_dadda_rca24_fa288_y4;
  wire f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa284_y4;
  wire f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa283_y4;
  wire f_s_dadda_rca24_fa289_y0;
  wire f_s_dadda_rca24_fa289_y1;
  wire f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa282_y4;
  wire f_s_dadda_rca24_fa289_y2;
  wire f_s_dadda_rca24_fa289_y3;
  wire f_s_dadda_rca24_fa289_y4;
  wire f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa281_y4;
  wire f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa280_y4;
  wire f_s_dadda_rca24_fa290_y0;
  wire f_s_dadda_rca24_fa290_y1;
  wire f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa279_y4;
  wire f_s_dadda_rca24_fa290_y2;
  wire f_s_dadda_rca24_fa290_y3;
  wire f_s_dadda_rca24_fa290_y4;
  wire f_s_dadda_rca24_nand_23_11_a_23;
  wire f_s_dadda_rca24_nand_23_11_b_11;
  wire f_s_dadda_rca24_nand_23_11_y0;
  wire f_s_dadda_rca24_and_22_12_a_22;
  wire f_s_dadda_rca24_and_22_12_b_12;
  wire f_s_dadda_rca24_and_22_12_y0;
  wire f_s_dadda_rca24_and_21_13_a_21;
  wire f_s_dadda_rca24_and_21_13_b_13;
  wire f_s_dadda_rca24_and_21_13_y0;
  wire f_s_dadda_rca24_fa291_f_s_dadda_rca24_nand_23_11_y0;
  wire f_s_dadda_rca24_fa291_f_s_dadda_rca24_and_22_12_y0;
  wire f_s_dadda_rca24_fa291_y0;
  wire f_s_dadda_rca24_fa291_y1;
  wire f_s_dadda_rca24_fa291_f_s_dadda_rca24_and_21_13_y0;
  wire f_s_dadda_rca24_fa291_y2;
  wire f_s_dadda_rca24_fa291_y3;
  wire f_s_dadda_rca24_fa291_y4;
  wire f_s_dadda_rca24_and_20_14_a_20;
  wire f_s_dadda_rca24_and_20_14_b_14;
  wire f_s_dadda_rca24_and_20_14_y0;
  wire f_s_dadda_rca24_and_19_15_a_19;
  wire f_s_dadda_rca24_and_19_15_b_15;
  wire f_s_dadda_rca24_and_19_15_y0;
  wire f_s_dadda_rca24_and_18_16_a_18;
  wire f_s_dadda_rca24_and_18_16_b_16;
  wire f_s_dadda_rca24_and_18_16_y0;
  wire f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_20_14_y0;
  wire f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_19_15_y0;
  wire f_s_dadda_rca24_fa292_y0;
  wire f_s_dadda_rca24_fa292_y1;
  wire f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_18_16_y0;
  wire f_s_dadda_rca24_fa292_y2;
  wire f_s_dadda_rca24_fa292_y3;
  wire f_s_dadda_rca24_fa292_y4;
  wire f_s_dadda_rca24_and_17_17_a_17;
  wire f_s_dadda_rca24_and_17_17_b_17;
  wire f_s_dadda_rca24_and_17_17_y0;
  wire f_s_dadda_rca24_and_16_18_a_16;
  wire f_s_dadda_rca24_and_16_18_b_18;
  wire f_s_dadda_rca24_and_16_18_y0;
  wire f_s_dadda_rca24_and_15_19_a_15;
  wire f_s_dadda_rca24_and_15_19_b_19;
  wire f_s_dadda_rca24_and_15_19_y0;
  wire f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_17_17_y0;
  wire f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_16_18_y0;
  wire f_s_dadda_rca24_fa293_y0;
  wire f_s_dadda_rca24_fa293_y1;
  wire f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_15_19_y0;
  wire f_s_dadda_rca24_fa293_y2;
  wire f_s_dadda_rca24_fa293_y3;
  wire f_s_dadda_rca24_fa293_y4;
  wire f_s_dadda_rca24_and_14_20_a_14;
  wire f_s_dadda_rca24_and_14_20_b_20;
  wire f_s_dadda_rca24_and_14_20_y0;
  wire f_s_dadda_rca24_and_13_21_a_13;
  wire f_s_dadda_rca24_and_13_21_b_21;
  wire f_s_dadda_rca24_and_13_21_y0;
  wire f_s_dadda_rca24_and_12_22_a_12;
  wire f_s_dadda_rca24_and_12_22_b_22;
  wire f_s_dadda_rca24_and_12_22_y0;
  wire f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_14_20_y0;
  wire f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_13_21_y0;
  wire f_s_dadda_rca24_fa294_y0;
  wire f_s_dadda_rca24_fa294_y1;
  wire f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_12_22_y0;
  wire f_s_dadda_rca24_fa294_y2;
  wire f_s_dadda_rca24_fa294_y3;
  wire f_s_dadda_rca24_fa294_y4;
  wire f_s_dadda_rca24_nand_11_23_a_11;
  wire f_s_dadda_rca24_nand_11_23_b_23;
  wire f_s_dadda_rca24_nand_11_23_y0;
  wire f_s_dadda_rca24_fa295_f_s_dadda_rca24_nand_11_23_y0;
  wire f_s_dadda_rca24_fa295_f_s_dadda_rca24_fa288_y2;
  wire f_s_dadda_rca24_fa295_y0;
  wire f_s_dadda_rca24_fa295_y1;
  wire f_s_dadda_rca24_fa295_f_s_dadda_rca24_fa289_y2;
  wire f_s_dadda_rca24_fa295_y2;
  wire f_s_dadda_rca24_fa295_y3;
  wire f_s_dadda_rca24_fa295_y4;
  wire f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa295_y4;
  wire f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa294_y4;
  wire f_s_dadda_rca24_fa296_y0;
  wire f_s_dadda_rca24_fa296_y1;
  wire f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa293_y4;
  wire f_s_dadda_rca24_fa296_y2;
  wire f_s_dadda_rca24_fa296_y3;
  wire f_s_dadda_rca24_fa296_y4;
  wire f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa292_y4;
  wire f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa291_y4;
  wire f_s_dadda_rca24_fa297_y0;
  wire f_s_dadda_rca24_fa297_y1;
  wire f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa290_y4;
  wire f_s_dadda_rca24_fa297_y2;
  wire f_s_dadda_rca24_fa297_y3;
  wire f_s_dadda_rca24_fa297_y4;
  wire f_s_dadda_rca24_nand_23_12_a_23;
  wire f_s_dadda_rca24_nand_23_12_b_12;
  wire f_s_dadda_rca24_nand_23_12_y0;
  wire f_s_dadda_rca24_fa298_f_s_dadda_rca24_fa289_y4;
  wire f_s_dadda_rca24_fa298_f_s_dadda_rca24_fa288_y4;
  wire f_s_dadda_rca24_fa298_y0;
  wire f_s_dadda_rca24_fa298_y1;
  wire f_s_dadda_rca24_fa298_f_s_dadda_rca24_nand_23_12_y0;
  wire f_s_dadda_rca24_fa298_y2;
  wire f_s_dadda_rca24_fa298_y3;
  wire f_s_dadda_rca24_fa298_y4;
  wire f_s_dadda_rca24_and_22_13_a_22;
  wire f_s_dadda_rca24_and_22_13_b_13;
  wire f_s_dadda_rca24_and_22_13_y0;
  wire f_s_dadda_rca24_and_21_14_a_21;
  wire f_s_dadda_rca24_and_21_14_b_14;
  wire f_s_dadda_rca24_and_21_14_y0;
  wire f_s_dadda_rca24_and_20_15_a_20;
  wire f_s_dadda_rca24_and_20_15_b_15;
  wire f_s_dadda_rca24_and_20_15_y0;
  wire f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_22_13_y0;
  wire f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_21_14_y0;
  wire f_s_dadda_rca24_fa299_y0;
  wire f_s_dadda_rca24_fa299_y1;
  wire f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_20_15_y0;
  wire f_s_dadda_rca24_fa299_y2;
  wire f_s_dadda_rca24_fa299_y3;
  wire f_s_dadda_rca24_fa299_y4;
  wire f_s_dadda_rca24_and_19_16_a_19;
  wire f_s_dadda_rca24_and_19_16_b_16;
  wire f_s_dadda_rca24_and_19_16_y0;
  wire f_s_dadda_rca24_and_18_17_a_18;
  wire f_s_dadda_rca24_and_18_17_b_17;
  wire f_s_dadda_rca24_and_18_17_y0;
  wire f_s_dadda_rca24_and_17_18_a_17;
  wire f_s_dadda_rca24_and_17_18_b_18;
  wire f_s_dadda_rca24_and_17_18_y0;
  wire f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_19_16_y0;
  wire f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_18_17_y0;
  wire f_s_dadda_rca24_fa300_y0;
  wire f_s_dadda_rca24_fa300_y1;
  wire f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_17_18_y0;
  wire f_s_dadda_rca24_fa300_y2;
  wire f_s_dadda_rca24_fa300_y3;
  wire f_s_dadda_rca24_fa300_y4;
  wire f_s_dadda_rca24_and_16_19_a_16;
  wire f_s_dadda_rca24_and_16_19_b_19;
  wire f_s_dadda_rca24_and_16_19_y0;
  wire f_s_dadda_rca24_and_15_20_a_15;
  wire f_s_dadda_rca24_and_15_20_b_20;
  wire f_s_dadda_rca24_and_15_20_y0;
  wire f_s_dadda_rca24_and_14_21_a_14;
  wire f_s_dadda_rca24_and_14_21_b_21;
  wire f_s_dadda_rca24_and_14_21_y0;
  wire f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_16_19_y0;
  wire f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_15_20_y0;
  wire f_s_dadda_rca24_fa301_y0;
  wire f_s_dadda_rca24_fa301_y1;
  wire f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_14_21_y0;
  wire f_s_dadda_rca24_fa301_y2;
  wire f_s_dadda_rca24_fa301_y3;
  wire f_s_dadda_rca24_fa301_y4;
  wire f_s_dadda_rca24_and_13_22_a_13;
  wire f_s_dadda_rca24_and_13_22_b_22;
  wire f_s_dadda_rca24_and_13_22_y0;
  wire f_s_dadda_rca24_nand_12_23_a_12;
  wire f_s_dadda_rca24_nand_12_23_b_23;
  wire f_s_dadda_rca24_nand_12_23_y0;
  wire f_s_dadda_rca24_fa302_f_s_dadda_rca24_and_13_22_y0;
  wire f_s_dadda_rca24_fa302_f_s_dadda_rca24_nand_12_23_y0;
  wire f_s_dadda_rca24_fa302_y0;
  wire f_s_dadda_rca24_fa302_y1;
  wire f_s_dadda_rca24_fa302_f_s_dadda_rca24_fa296_y2;
  wire f_s_dadda_rca24_fa302_y2;
  wire f_s_dadda_rca24_fa302_y3;
  wire f_s_dadda_rca24_fa302_y4;
  wire f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa302_y4;
  wire f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa301_y4;
  wire f_s_dadda_rca24_fa303_y0;
  wire f_s_dadda_rca24_fa303_y1;
  wire f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa300_y4;
  wire f_s_dadda_rca24_fa303_y2;
  wire f_s_dadda_rca24_fa303_y3;
  wire f_s_dadda_rca24_fa303_y4;
  wire f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa299_y4;
  wire f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa298_y4;
  wire f_s_dadda_rca24_fa304_y0;
  wire f_s_dadda_rca24_fa304_y1;
  wire f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa297_y4;
  wire f_s_dadda_rca24_fa304_y2;
  wire f_s_dadda_rca24_fa304_y3;
  wire f_s_dadda_rca24_fa304_y4;
  wire f_s_dadda_rca24_nand_23_13_a_23;
  wire f_s_dadda_rca24_nand_23_13_b_13;
  wire f_s_dadda_rca24_nand_23_13_y0;
  wire f_s_dadda_rca24_and_22_14_a_22;
  wire f_s_dadda_rca24_and_22_14_b_14;
  wire f_s_dadda_rca24_and_22_14_y0;
  wire f_s_dadda_rca24_fa305_f_s_dadda_rca24_fa296_y4;
  wire f_s_dadda_rca24_fa305_f_s_dadda_rca24_nand_23_13_y0;
  wire f_s_dadda_rca24_fa305_y0;
  wire f_s_dadda_rca24_fa305_y1;
  wire f_s_dadda_rca24_fa305_f_s_dadda_rca24_and_22_14_y0;
  wire f_s_dadda_rca24_fa305_y2;
  wire f_s_dadda_rca24_fa305_y3;
  wire f_s_dadda_rca24_fa305_y4;
  wire f_s_dadda_rca24_and_21_15_a_21;
  wire f_s_dadda_rca24_and_21_15_b_15;
  wire f_s_dadda_rca24_and_21_15_y0;
  wire f_s_dadda_rca24_and_20_16_a_20;
  wire f_s_dadda_rca24_and_20_16_b_16;
  wire f_s_dadda_rca24_and_20_16_y0;
  wire f_s_dadda_rca24_and_19_17_a_19;
  wire f_s_dadda_rca24_and_19_17_b_17;
  wire f_s_dadda_rca24_and_19_17_y0;
  wire f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_21_15_y0;
  wire f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_20_16_y0;
  wire f_s_dadda_rca24_fa306_y0;
  wire f_s_dadda_rca24_fa306_y1;
  wire f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_19_17_y0;
  wire f_s_dadda_rca24_fa306_y2;
  wire f_s_dadda_rca24_fa306_y3;
  wire f_s_dadda_rca24_fa306_y4;
  wire f_s_dadda_rca24_and_18_18_a_18;
  wire f_s_dadda_rca24_and_18_18_b_18;
  wire f_s_dadda_rca24_and_18_18_y0;
  wire f_s_dadda_rca24_and_17_19_a_17;
  wire f_s_dadda_rca24_and_17_19_b_19;
  wire f_s_dadda_rca24_and_17_19_y0;
  wire f_s_dadda_rca24_and_16_20_a_16;
  wire f_s_dadda_rca24_and_16_20_b_20;
  wire f_s_dadda_rca24_and_16_20_y0;
  wire f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_18_18_y0;
  wire f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_17_19_y0;
  wire f_s_dadda_rca24_fa307_y0;
  wire f_s_dadda_rca24_fa307_y1;
  wire f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_16_20_y0;
  wire f_s_dadda_rca24_fa307_y2;
  wire f_s_dadda_rca24_fa307_y3;
  wire f_s_dadda_rca24_fa307_y4;
  wire f_s_dadda_rca24_and_15_21_a_15;
  wire f_s_dadda_rca24_and_15_21_b_21;
  wire f_s_dadda_rca24_and_15_21_y0;
  wire f_s_dadda_rca24_and_14_22_a_14;
  wire f_s_dadda_rca24_and_14_22_b_22;
  wire f_s_dadda_rca24_and_14_22_y0;
  wire f_s_dadda_rca24_nand_13_23_a_13;
  wire f_s_dadda_rca24_nand_13_23_b_23;
  wire f_s_dadda_rca24_nand_13_23_y0;
  wire f_s_dadda_rca24_fa308_f_s_dadda_rca24_and_15_21_y0;
  wire f_s_dadda_rca24_fa308_f_s_dadda_rca24_and_14_22_y0;
  wire f_s_dadda_rca24_fa308_y0;
  wire f_s_dadda_rca24_fa308_y1;
  wire f_s_dadda_rca24_fa308_f_s_dadda_rca24_nand_13_23_y0;
  wire f_s_dadda_rca24_fa308_y2;
  wire f_s_dadda_rca24_fa308_y3;
  wire f_s_dadda_rca24_fa308_y4;
  wire f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa308_y4;
  wire f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa307_y4;
  wire f_s_dadda_rca24_fa309_y0;
  wire f_s_dadda_rca24_fa309_y1;
  wire f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa306_y4;
  wire f_s_dadda_rca24_fa309_y2;
  wire f_s_dadda_rca24_fa309_y3;
  wire f_s_dadda_rca24_fa309_y4;
  wire f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa305_y4;
  wire f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa304_y4;
  wire f_s_dadda_rca24_fa310_y0;
  wire f_s_dadda_rca24_fa310_y1;
  wire f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa303_y4;
  wire f_s_dadda_rca24_fa310_y2;
  wire f_s_dadda_rca24_fa310_y3;
  wire f_s_dadda_rca24_fa310_y4;
  wire f_s_dadda_rca24_nand_23_14_a_23;
  wire f_s_dadda_rca24_nand_23_14_b_14;
  wire f_s_dadda_rca24_nand_23_14_y0;
  wire f_s_dadda_rca24_and_22_15_a_22;
  wire f_s_dadda_rca24_and_22_15_b_15;
  wire f_s_dadda_rca24_and_22_15_y0;
  wire f_s_dadda_rca24_and_21_16_a_21;
  wire f_s_dadda_rca24_and_21_16_b_16;
  wire f_s_dadda_rca24_and_21_16_y0;
  wire f_s_dadda_rca24_fa311_f_s_dadda_rca24_nand_23_14_y0;
  wire f_s_dadda_rca24_fa311_f_s_dadda_rca24_and_22_15_y0;
  wire f_s_dadda_rca24_fa311_y0;
  wire f_s_dadda_rca24_fa311_y1;
  wire f_s_dadda_rca24_fa311_f_s_dadda_rca24_and_21_16_y0;
  wire f_s_dadda_rca24_fa311_y2;
  wire f_s_dadda_rca24_fa311_y3;
  wire f_s_dadda_rca24_fa311_y4;
  wire f_s_dadda_rca24_and_20_17_a_20;
  wire f_s_dadda_rca24_and_20_17_b_17;
  wire f_s_dadda_rca24_and_20_17_y0;
  wire f_s_dadda_rca24_and_19_18_a_19;
  wire f_s_dadda_rca24_and_19_18_b_18;
  wire f_s_dadda_rca24_and_19_18_y0;
  wire f_s_dadda_rca24_and_18_19_a_18;
  wire f_s_dadda_rca24_and_18_19_b_19;
  wire f_s_dadda_rca24_and_18_19_y0;
  wire f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_20_17_y0;
  wire f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_19_18_y0;
  wire f_s_dadda_rca24_fa312_y0;
  wire f_s_dadda_rca24_fa312_y1;
  wire f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_18_19_y0;
  wire f_s_dadda_rca24_fa312_y2;
  wire f_s_dadda_rca24_fa312_y3;
  wire f_s_dadda_rca24_fa312_y4;
  wire f_s_dadda_rca24_and_17_20_a_17;
  wire f_s_dadda_rca24_and_17_20_b_20;
  wire f_s_dadda_rca24_and_17_20_y0;
  wire f_s_dadda_rca24_and_16_21_a_16;
  wire f_s_dadda_rca24_and_16_21_b_21;
  wire f_s_dadda_rca24_and_16_21_y0;
  wire f_s_dadda_rca24_and_15_22_a_15;
  wire f_s_dadda_rca24_and_15_22_b_22;
  wire f_s_dadda_rca24_and_15_22_y0;
  wire f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_17_20_y0;
  wire f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_16_21_y0;
  wire f_s_dadda_rca24_fa313_y0;
  wire f_s_dadda_rca24_fa313_y1;
  wire f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_15_22_y0;
  wire f_s_dadda_rca24_fa313_y2;
  wire f_s_dadda_rca24_fa313_y3;
  wire f_s_dadda_rca24_fa313_y4;
  wire f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa313_y4;
  wire f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa312_y4;
  wire f_s_dadda_rca24_fa314_y0;
  wire f_s_dadda_rca24_fa314_y1;
  wire f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa311_y4;
  wire f_s_dadda_rca24_fa314_y2;
  wire f_s_dadda_rca24_fa314_y3;
  wire f_s_dadda_rca24_fa314_y4;
  wire f_s_dadda_rca24_nand_23_15_a_23;
  wire f_s_dadda_rca24_nand_23_15_b_15;
  wire f_s_dadda_rca24_nand_23_15_y0;
  wire f_s_dadda_rca24_fa315_f_s_dadda_rca24_fa310_y4;
  wire f_s_dadda_rca24_fa315_f_s_dadda_rca24_fa309_y4;
  wire f_s_dadda_rca24_fa315_y0;
  wire f_s_dadda_rca24_fa315_y1;
  wire f_s_dadda_rca24_fa315_f_s_dadda_rca24_nand_23_15_y0;
  wire f_s_dadda_rca24_fa315_y2;
  wire f_s_dadda_rca24_fa315_y3;
  wire f_s_dadda_rca24_fa315_y4;
  wire f_s_dadda_rca24_and_22_16_a_22;
  wire f_s_dadda_rca24_and_22_16_b_16;
  wire f_s_dadda_rca24_and_22_16_y0;
  wire f_s_dadda_rca24_and_21_17_a_21;
  wire f_s_dadda_rca24_and_21_17_b_17;
  wire f_s_dadda_rca24_and_21_17_y0;
  wire f_s_dadda_rca24_and_20_18_a_20;
  wire f_s_dadda_rca24_and_20_18_b_18;
  wire f_s_dadda_rca24_and_20_18_y0;
  wire f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_22_16_y0;
  wire f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_21_17_y0;
  wire f_s_dadda_rca24_fa316_y0;
  wire f_s_dadda_rca24_fa316_y1;
  wire f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_20_18_y0;
  wire f_s_dadda_rca24_fa316_y2;
  wire f_s_dadda_rca24_fa316_y3;
  wire f_s_dadda_rca24_fa316_y4;
  wire f_s_dadda_rca24_and_19_19_a_19;
  wire f_s_dadda_rca24_and_19_19_b_19;
  wire f_s_dadda_rca24_and_19_19_y0;
  wire f_s_dadda_rca24_and_18_20_a_18;
  wire f_s_dadda_rca24_and_18_20_b_20;
  wire f_s_dadda_rca24_and_18_20_y0;
  wire f_s_dadda_rca24_and_17_21_a_17;
  wire f_s_dadda_rca24_and_17_21_b_21;
  wire f_s_dadda_rca24_and_17_21_y0;
  wire f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_19_19_y0;
  wire f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_18_20_y0;
  wire f_s_dadda_rca24_fa317_y0;
  wire f_s_dadda_rca24_fa317_y1;
  wire f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_17_21_y0;
  wire f_s_dadda_rca24_fa317_y2;
  wire f_s_dadda_rca24_fa317_y3;
  wire f_s_dadda_rca24_fa317_y4;
  wire f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa317_y4;
  wire f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa316_y4;
  wire f_s_dadda_rca24_fa318_y0;
  wire f_s_dadda_rca24_fa318_y1;
  wire f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa315_y4;
  wire f_s_dadda_rca24_fa318_y2;
  wire f_s_dadda_rca24_fa318_y3;
  wire f_s_dadda_rca24_fa318_y4;
  wire f_s_dadda_rca24_nand_23_16_a_23;
  wire f_s_dadda_rca24_nand_23_16_b_16;
  wire f_s_dadda_rca24_nand_23_16_y0;
  wire f_s_dadda_rca24_and_22_17_a_22;
  wire f_s_dadda_rca24_and_22_17_b_17;
  wire f_s_dadda_rca24_and_22_17_y0;
  wire f_s_dadda_rca24_fa319_f_s_dadda_rca24_fa314_y4;
  wire f_s_dadda_rca24_fa319_f_s_dadda_rca24_nand_23_16_y0;
  wire f_s_dadda_rca24_fa319_y0;
  wire f_s_dadda_rca24_fa319_y1;
  wire f_s_dadda_rca24_fa319_f_s_dadda_rca24_and_22_17_y0;
  wire f_s_dadda_rca24_fa319_y2;
  wire f_s_dadda_rca24_fa319_y3;
  wire f_s_dadda_rca24_fa319_y4;
  wire f_s_dadda_rca24_and_21_18_a_21;
  wire f_s_dadda_rca24_and_21_18_b_18;
  wire f_s_dadda_rca24_and_21_18_y0;
  wire f_s_dadda_rca24_and_20_19_a_20;
  wire f_s_dadda_rca24_and_20_19_b_19;
  wire f_s_dadda_rca24_and_20_19_y0;
  wire f_s_dadda_rca24_and_19_20_a_19;
  wire f_s_dadda_rca24_and_19_20_b_20;
  wire f_s_dadda_rca24_and_19_20_y0;
  wire f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_21_18_y0;
  wire f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_20_19_y0;
  wire f_s_dadda_rca24_fa320_y0;
  wire f_s_dadda_rca24_fa320_y1;
  wire f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_19_20_y0;
  wire f_s_dadda_rca24_fa320_y2;
  wire f_s_dadda_rca24_fa320_y3;
  wire f_s_dadda_rca24_fa320_y4;
  wire f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa320_y4;
  wire f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa319_y4;
  wire f_s_dadda_rca24_fa321_y0;
  wire f_s_dadda_rca24_fa321_y1;
  wire f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa318_y4;
  wire f_s_dadda_rca24_fa321_y2;
  wire f_s_dadda_rca24_fa321_y3;
  wire f_s_dadda_rca24_fa321_y4;
  wire f_s_dadda_rca24_nand_23_17_a_23;
  wire f_s_dadda_rca24_nand_23_17_b_17;
  wire f_s_dadda_rca24_nand_23_17_y0;
  wire f_s_dadda_rca24_and_22_18_a_22;
  wire f_s_dadda_rca24_and_22_18_b_18;
  wire f_s_dadda_rca24_and_22_18_y0;
  wire f_s_dadda_rca24_and_21_19_a_21;
  wire f_s_dadda_rca24_and_21_19_b_19;
  wire f_s_dadda_rca24_and_21_19_y0;
  wire f_s_dadda_rca24_fa322_f_s_dadda_rca24_nand_23_17_y0;
  wire f_s_dadda_rca24_fa322_f_s_dadda_rca24_and_22_18_y0;
  wire f_s_dadda_rca24_fa322_y0;
  wire f_s_dadda_rca24_fa322_y1;
  wire f_s_dadda_rca24_fa322_f_s_dadda_rca24_and_21_19_y0;
  wire f_s_dadda_rca24_fa322_y2;
  wire f_s_dadda_rca24_fa322_y3;
  wire f_s_dadda_rca24_fa322_y4;
  wire f_s_dadda_rca24_nand_23_18_a_23;
  wire f_s_dadda_rca24_nand_23_18_b_18;
  wire f_s_dadda_rca24_nand_23_18_y0;
  wire f_s_dadda_rca24_fa323_f_s_dadda_rca24_fa322_y4;
  wire f_s_dadda_rca24_fa323_f_s_dadda_rca24_fa321_y4;
  wire f_s_dadda_rca24_fa323_y0;
  wire f_s_dadda_rca24_fa323_y1;
  wire f_s_dadda_rca24_fa323_f_s_dadda_rca24_nand_23_18_y0;
  wire f_s_dadda_rca24_fa323_y2;
  wire f_s_dadda_rca24_fa323_y3;
  wire f_s_dadda_rca24_fa323_y4;
  wire f_s_dadda_rca24_and_4_0_a_4;
  wire f_s_dadda_rca24_and_4_0_b_0;
  wire f_s_dadda_rca24_and_4_0_y0;
  wire f_s_dadda_rca24_and_3_1_a_3;
  wire f_s_dadda_rca24_and_3_1_b_1;
  wire f_s_dadda_rca24_and_3_1_y0;
  wire f_s_dadda_rca24_ha18_f_s_dadda_rca24_and_4_0_y0;
  wire f_s_dadda_rca24_ha18_f_s_dadda_rca24_and_3_1_y0;
  wire f_s_dadda_rca24_ha18_y0;
  wire f_s_dadda_rca24_ha18_y1;
  wire f_s_dadda_rca24_and_5_0_a_5;
  wire f_s_dadda_rca24_and_5_0_b_0;
  wire f_s_dadda_rca24_and_5_0_y0;
  wire f_s_dadda_rca24_and_4_1_a_4;
  wire f_s_dadda_rca24_and_4_1_b_1;
  wire f_s_dadda_rca24_and_4_1_y0;
  wire f_s_dadda_rca24_fa324_f_s_dadda_rca24_ha18_y1;
  wire f_s_dadda_rca24_fa324_f_s_dadda_rca24_and_5_0_y0;
  wire f_s_dadda_rca24_fa324_y0;
  wire f_s_dadda_rca24_fa324_y1;
  wire f_s_dadda_rca24_fa324_f_s_dadda_rca24_and_4_1_y0;
  wire f_s_dadda_rca24_fa324_y2;
  wire f_s_dadda_rca24_fa324_y3;
  wire f_s_dadda_rca24_fa324_y4;
  wire f_s_dadda_rca24_and_3_2_a_3;
  wire f_s_dadda_rca24_and_3_2_b_2;
  wire f_s_dadda_rca24_and_3_2_y0;
  wire f_s_dadda_rca24_and_2_3_a_2;
  wire f_s_dadda_rca24_and_2_3_b_3;
  wire f_s_dadda_rca24_and_2_3_y0;
  wire f_s_dadda_rca24_ha19_f_s_dadda_rca24_and_3_2_y0;
  wire f_s_dadda_rca24_ha19_f_s_dadda_rca24_and_2_3_y0;
  wire f_s_dadda_rca24_ha19_y0;
  wire f_s_dadda_rca24_ha19_y1;
  wire f_s_dadda_rca24_and_4_2_a_4;
  wire f_s_dadda_rca24_and_4_2_b_2;
  wire f_s_dadda_rca24_and_4_2_y0;
  wire f_s_dadda_rca24_fa325_f_s_dadda_rca24_ha19_y1;
  wire f_s_dadda_rca24_fa325_f_s_dadda_rca24_fa324_y4;
  wire f_s_dadda_rca24_fa325_y0;
  wire f_s_dadda_rca24_fa325_y1;
  wire f_s_dadda_rca24_fa325_f_s_dadda_rca24_and_4_2_y0;
  wire f_s_dadda_rca24_fa325_y2;
  wire f_s_dadda_rca24_fa325_y3;
  wire f_s_dadda_rca24_fa325_y4;
  wire f_s_dadda_rca24_and_3_3_a_3;
  wire f_s_dadda_rca24_and_3_3_b_3;
  wire f_s_dadda_rca24_and_3_3_y0;
  wire f_s_dadda_rca24_and_2_4_a_2;
  wire f_s_dadda_rca24_and_2_4_b_4;
  wire f_s_dadda_rca24_and_2_4_y0;
  wire f_s_dadda_rca24_and_1_5_a_1;
  wire f_s_dadda_rca24_and_1_5_b_5;
  wire f_s_dadda_rca24_and_1_5_y0;
  wire f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_3_3_y0;
  wire f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_2_4_y0;
  wire f_s_dadda_rca24_fa326_y0;
  wire f_s_dadda_rca24_fa326_y1;
  wire f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_1_5_y0;
  wire f_s_dadda_rca24_fa326_y2;
  wire f_s_dadda_rca24_fa326_y3;
  wire f_s_dadda_rca24_fa326_y4;
  wire f_s_dadda_rca24_and_3_4_a_3;
  wire f_s_dadda_rca24_and_3_4_b_4;
  wire f_s_dadda_rca24_and_3_4_y0;
  wire f_s_dadda_rca24_fa327_f_s_dadda_rca24_fa326_y4;
  wire f_s_dadda_rca24_fa327_f_s_dadda_rca24_fa325_y4;
  wire f_s_dadda_rca24_fa327_y0;
  wire f_s_dadda_rca24_fa327_y1;
  wire f_s_dadda_rca24_fa327_f_s_dadda_rca24_and_3_4_y0;
  wire f_s_dadda_rca24_fa327_y2;
  wire f_s_dadda_rca24_fa327_y3;
  wire f_s_dadda_rca24_fa327_y4;
  wire f_s_dadda_rca24_and_2_5_a_2;
  wire f_s_dadda_rca24_and_2_5_b_5;
  wire f_s_dadda_rca24_and_2_5_y0;
  wire f_s_dadda_rca24_and_1_6_a_1;
  wire f_s_dadda_rca24_and_1_6_b_6;
  wire f_s_dadda_rca24_and_1_6_y0;
  wire f_s_dadda_rca24_and_0_7_a_0;
  wire f_s_dadda_rca24_and_0_7_b_7;
  wire f_s_dadda_rca24_and_0_7_y0;
  wire f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_2_5_y0;
  wire f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_1_6_y0;
  wire f_s_dadda_rca24_fa328_y0;
  wire f_s_dadda_rca24_fa328_y1;
  wire f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_0_7_y0;
  wire f_s_dadda_rca24_fa328_y2;
  wire f_s_dadda_rca24_fa328_y3;
  wire f_s_dadda_rca24_fa328_y4;
  wire f_s_dadda_rca24_and_2_6_a_2;
  wire f_s_dadda_rca24_and_2_6_b_6;
  wire f_s_dadda_rca24_and_2_6_y0;
  wire f_s_dadda_rca24_fa329_f_s_dadda_rca24_fa328_y4;
  wire f_s_dadda_rca24_fa329_f_s_dadda_rca24_fa327_y4;
  wire f_s_dadda_rca24_fa329_y0;
  wire f_s_dadda_rca24_fa329_y1;
  wire f_s_dadda_rca24_fa329_f_s_dadda_rca24_and_2_6_y0;
  wire f_s_dadda_rca24_fa329_y2;
  wire f_s_dadda_rca24_fa329_y3;
  wire f_s_dadda_rca24_fa329_y4;
  wire f_s_dadda_rca24_and_1_7_a_1;
  wire f_s_dadda_rca24_and_1_7_b_7;
  wire f_s_dadda_rca24_and_1_7_y0;
  wire f_s_dadda_rca24_and_0_8_a_0;
  wire f_s_dadda_rca24_and_0_8_b_8;
  wire f_s_dadda_rca24_and_0_8_y0;
  wire f_s_dadda_rca24_fa330_f_s_dadda_rca24_and_1_7_y0;
  wire f_s_dadda_rca24_fa330_f_s_dadda_rca24_and_0_8_y0;
  wire f_s_dadda_rca24_fa330_y0;
  wire f_s_dadda_rca24_fa330_y1;
  wire f_s_dadda_rca24_fa330_f_s_dadda_rca24_fa26_y2;
  wire f_s_dadda_rca24_fa330_y2;
  wire f_s_dadda_rca24_fa330_y3;
  wire f_s_dadda_rca24_fa330_y4;
  wire f_s_dadda_rca24_and_1_8_a_1;
  wire f_s_dadda_rca24_and_1_8_b_8;
  wire f_s_dadda_rca24_and_1_8_y0;
  wire f_s_dadda_rca24_fa331_f_s_dadda_rca24_fa330_y4;
  wire f_s_dadda_rca24_fa331_f_s_dadda_rca24_fa329_y4;
  wire f_s_dadda_rca24_fa331_y0;
  wire f_s_dadda_rca24_fa331_y1;
  wire f_s_dadda_rca24_fa331_f_s_dadda_rca24_and_1_8_y0;
  wire f_s_dadda_rca24_fa331_y2;
  wire f_s_dadda_rca24_fa331_y3;
  wire f_s_dadda_rca24_fa331_y4;
  wire f_s_dadda_rca24_and_0_9_a_0;
  wire f_s_dadda_rca24_and_0_9_b_9;
  wire f_s_dadda_rca24_and_0_9_y0;
  wire f_s_dadda_rca24_fa332_f_s_dadda_rca24_and_0_9_y0;
  wire f_s_dadda_rca24_fa332_f_s_dadda_rca24_fa28_y2;
  wire f_s_dadda_rca24_fa332_y0;
  wire f_s_dadda_rca24_fa332_y1;
  wire f_s_dadda_rca24_fa332_f_s_dadda_rca24_fa29_y2;
  wire f_s_dadda_rca24_fa332_y2;
  wire f_s_dadda_rca24_fa332_y3;
  wire f_s_dadda_rca24_fa332_y4;
  wire f_s_dadda_rca24_and_0_10_a_0;
  wire f_s_dadda_rca24_and_0_10_b_10;
  wire f_s_dadda_rca24_and_0_10_y0;
  wire f_s_dadda_rca24_fa333_f_s_dadda_rca24_fa332_y4;
  wire f_s_dadda_rca24_fa333_f_s_dadda_rca24_fa331_y4;
  wire f_s_dadda_rca24_fa333_y0;
  wire f_s_dadda_rca24_fa333_y1;
  wire f_s_dadda_rca24_fa333_f_s_dadda_rca24_and_0_10_y0;
  wire f_s_dadda_rca24_fa333_y2;
  wire f_s_dadda_rca24_fa333_y3;
  wire f_s_dadda_rca24_fa333_y4;
  wire f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa31_y2;
  wire f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa32_y2;
  wire f_s_dadda_rca24_fa334_y0;
  wire f_s_dadda_rca24_fa334_y1;
  wire f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa33_y2;
  wire f_s_dadda_rca24_fa334_y2;
  wire f_s_dadda_rca24_fa334_y3;
  wire f_s_dadda_rca24_fa334_y4;
  wire f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa334_y4;
  wire f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa333_y4;
  wire f_s_dadda_rca24_fa335_y0;
  wire f_s_dadda_rca24_fa335_y1;
  wire f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa35_y2;
  wire f_s_dadda_rca24_fa335_y2;
  wire f_s_dadda_rca24_fa335_y3;
  wire f_s_dadda_rca24_fa335_y4;
  wire f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa36_y2;
  wire f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa37_y2;
  wire f_s_dadda_rca24_fa336_y0;
  wire f_s_dadda_rca24_fa336_y1;
  wire f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa38_y2;
  wire f_s_dadda_rca24_fa336_y2;
  wire f_s_dadda_rca24_fa336_y3;
  wire f_s_dadda_rca24_fa336_y4;
  wire f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa336_y4;
  wire f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa335_y4;
  wire f_s_dadda_rca24_fa337_y0;
  wire f_s_dadda_rca24_fa337_y1;
  wire f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa41_y2;
  wire f_s_dadda_rca24_fa337_y2;
  wire f_s_dadda_rca24_fa337_y3;
  wire f_s_dadda_rca24_fa337_y4;
  wire f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa42_y2;
  wire f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa43_y2;
  wire f_s_dadda_rca24_fa338_y0;
  wire f_s_dadda_rca24_fa338_y1;
  wire f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa44_y2;
  wire f_s_dadda_rca24_fa338_y2;
  wire f_s_dadda_rca24_fa338_y3;
  wire f_s_dadda_rca24_fa338_y4;
  wire f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa338_y4;
  wire f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa337_y4;
  wire f_s_dadda_rca24_fa339_y0;
  wire f_s_dadda_rca24_fa339_y1;
  wire f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa48_y2;
  wire f_s_dadda_rca24_fa339_y2;
  wire f_s_dadda_rca24_fa339_y3;
  wire f_s_dadda_rca24_fa339_y4;
  wire f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa49_y2;
  wire f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa50_y2;
  wire f_s_dadda_rca24_fa340_y0;
  wire f_s_dadda_rca24_fa340_y1;
  wire f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa51_y2;
  wire f_s_dadda_rca24_fa340_y2;
  wire f_s_dadda_rca24_fa340_y3;
  wire f_s_dadda_rca24_fa340_y4;
  wire f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa340_y4;
  wire f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa339_y4;
  wire f_s_dadda_rca24_fa341_y0;
  wire f_s_dadda_rca24_fa341_y1;
  wire f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa56_y2;
  wire f_s_dadda_rca24_fa341_y2;
  wire f_s_dadda_rca24_fa341_y3;
  wire f_s_dadda_rca24_fa341_y4;
  wire f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa57_y2;
  wire f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa58_y2;
  wire f_s_dadda_rca24_fa342_y0;
  wire f_s_dadda_rca24_fa342_y1;
  wire f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa59_y2;
  wire f_s_dadda_rca24_fa342_y2;
  wire f_s_dadda_rca24_fa342_y3;
  wire f_s_dadda_rca24_fa342_y4;
  wire f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa342_y4;
  wire f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa341_y4;
  wire f_s_dadda_rca24_fa343_y0;
  wire f_s_dadda_rca24_fa343_y1;
  wire f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa65_y2;
  wire f_s_dadda_rca24_fa343_y2;
  wire f_s_dadda_rca24_fa343_y3;
  wire f_s_dadda_rca24_fa343_y4;
  wire f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa66_y2;
  wire f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa67_y2;
  wire f_s_dadda_rca24_fa344_y0;
  wire f_s_dadda_rca24_fa344_y1;
  wire f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa68_y2;
  wire f_s_dadda_rca24_fa344_y2;
  wire f_s_dadda_rca24_fa344_y3;
  wire f_s_dadda_rca24_fa344_y4;
  wire f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa344_y4;
  wire f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa343_y4;
  wire f_s_dadda_rca24_fa345_y0;
  wire f_s_dadda_rca24_fa345_y1;
  wire f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa75_y2;
  wire f_s_dadda_rca24_fa345_y2;
  wire f_s_dadda_rca24_fa345_y3;
  wire f_s_dadda_rca24_fa345_y4;
  wire f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa76_y2;
  wire f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa77_y2;
  wire f_s_dadda_rca24_fa346_y0;
  wire f_s_dadda_rca24_fa346_y1;
  wire f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa78_y2;
  wire f_s_dadda_rca24_fa346_y2;
  wire f_s_dadda_rca24_fa346_y3;
  wire f_s_dadda_rca24_fa346_y4;
  wire f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa346_y4;
  wire f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa345_y4;
  wire f_s_dadda_rca24_fa347_y0;
  wire f_s_dadda_rca24_fa347_y1;
  wire f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa86_y2;
  wire f_s_dadda_rca24_fa347_y2;
  wire f_s_dadda_rca24_fa347_y3;
  wire f_s_dadda_rca24_fa347_y4;
  wire f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa87_y2;
  wire f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa88_y2;
  wire f_s_dadda_rca24_fa348_y0;
  wire f_s_dadda_rca24_fa348_y1;
  wire f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa89_y2;
  wire f_s_dadda_rca24_fa348_y2;
  wire f_s_dadda_rca24_fa348_y3;
  wire f_s_dadda_rca24_fa348_y4;
  wire f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa348_y4;
  wire f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa347_y4;
  wire f_s_dadda_rca24_fa349_y0;
  wire f_s_dadda_rca24_fa349_y1;
  wire f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa98_y2;
  wire f_s_dadda_rca24_fa349_y2;
  wire f_s_dadda_rca24_fa349_y3;
  wire f_s_dadda_rca24_fa349_y4;
  wire f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa99_y2;
  wire f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa100_y2;
  wire f_s_dadda_rca24_fa350_y0;
  wire f_s_dadda_rca24_fa350_y1;
  wire f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa101_y2;
  wire f_s_dadda_rca24_fa350_y2;
  wire f_s_dadda_rca24_fa350_y3;
  wire f_s_dadda_rca24_fa350_y4;
  wire f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa350_y4;
  wire f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa349_y4;
  wire f_s_dadda_rca24_fa351_y0;
  wire f_s_dadda_rca24_fa351_y1;
  wire f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa110_y2;
  wire f_s_dadda_rca24_fa351_y2;
  wire f_s_dadda_rca24_fa351_y3;
  wire f_s_dadda_rca24_fa351_y4;
  wire f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa111_y2;
  wire f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa112_y2;
  wire f_s_dadda_rca24_fa352_y0;
  wire f_s_dadda_rca24_fa352_y1;
  wire f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa113_y2;
  wire f_s_dadda_rca24_fa352_y2;
  wire f_s_dadda_rca24_fa352_y3;
  wire f_s_dadda_rca24_fa352_y4;
  wire f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa352_y4;
  wire f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa351_y4;
  wire f_s_dadda_rca24_fa353_y0;
  wire f_s_dadda_rca24_fa353_y1;
  wire f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa123_y2;
  wire f_s_dadda_rca24_fa353_y2;
  wire f_s_dadda_rca24_fa353_y3;
  wire f_s_dadda_rca24_fa353_y4;
  wire f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa124_y2;
  wire f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa125_y2;
  wire f_s_dadda_rca24_fa354_y0;
  wire f_s_dadda_rca24_fa354_y1;
  wire f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa126_y2;
  wire f_s_dadda_rca24_fa354_y2;
  wire f_s_dadda_rca24_fa354_y3;
  wire f_s_dadda_rca24_fa354_y4;
  wire f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa354_y4;
  wire f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa353_y4;
  wire f_s_dadda_rca24_fa355_y0;
  wire f_s_dadda_rca24_fa355_y1;
  wire f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa136_y2;
  wire f_s_dadda_rca24_fa355_y2;
  wire f_s_dadda_rca24_fa355_y3;
  wire f_s_dadda_rca24_fa355_y4;
  wire f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa137_y2;
  wire f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa138_y2;
  wire f_s_dadda_rca24_fa356_y0;
  wire f_s_dadda_rca24_fa356_y1;
  wire f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa139_y2;
  wire f_s_dadda_rca24_fa356_y2;
  wire f_s_dadda_rca24_fa356_y3;
  wire f_s_dadda_rca24_fa356_y4;
  wire f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa356_y4;
  wire f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa355_y4;
  wire f_s_dadda_rca24_fa357_y0;
  wire f_s_dadda_rca24_fa357_y1;
  wire f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa149_y2;
  wire f_s_dadda_rca24_fa357_y2;
  wire f_s_dadda_rca24_fa357_y3;
  wire f_s_dadda_rca24_fa357_y4;
  wire f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa150_y2;
  wire f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa151_y2;
  wire f_s_dadda_rca24_fa358_y0;
  wire f_s_dadda_rca24_fa358_y1;
  wire f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa152_y2;
  wire f_s_dadda_rca24_fa358_y2;
  wire f_s_dadda_rca24_fa358_y3;
  wire f_s_dadda_rca24_fa358_y4;
  wire f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa358_y4;
  wire f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa357_y4;
  wire f_s_dadda_rca24_fa359_y0;
  wire f_s_dadda_rca24_fa359_y1;
  wire f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa162_y2;
  wire f_s_dadda_rca24_fa359_y2;
  wire f_s_dadda_rca24_fa359_y3;
  wire f_s_dadda_rca24_fa359_y4;
  wire f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa163_y2;
  wire f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa164_y2;
  wire f_s_dadda_rca24_fa360_y0;
  wire f_s_dadda_rca24_fa360_y1;
  wire f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa165_y2;
  wire f_s_dadda_rca24_fa360_y2;
  wire f_s_dadda_rca24_fa360_y3;
  wire f_s_dadda_rca24_fa360_y4;
  wire f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa360_y4;
  wire f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa359_y4;
  wire f_s_dadda_rca24_fa361_y0;
  wire f_s_dadda_rca24_fa361_y1;
  wire f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa175_y2;
  wire f_s_dadda_rca24_fa361_y2;
  wire f_s_dadda_rca24_fa361_y3;
  wire f_s_dadda_rca24_fa361_y4;
  wire f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa176_y2;
  wire f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa177_y2;
  wire f_s_dadda_rca24_fa362_y0;
  wire f_s_dadda_rca24_fa362_y1;
  wire f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa178_y2;
  wire f_s_dadda_rca24_fa362_y2;
  wire f_s_dadda_rca24_fa362_y3;
  wire f_s_dadda_rca24_fa362_y4;
  wire f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa362_y4;
  wire f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa361_y4;
  wire f_s_dadda_rca24_fa363_y0;
  wire f_s_dadda_rca24_fa363_y1;
  wire f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa188_y2;
  wire f_s_dadda_rca24_fa363_y2;
  wire f_s_dadda_rca24_fa363_y3;
  wire f_s_dadda_rca24_fa363_y4;
  wire f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa189_y2;
  wire f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa190_y2;
  wire f_s_dadda_rca24_fa364_y0;
  wire f_s_dadda_rca24_fa364_y1;
  wire f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa191_y2;
  wire f_s_dadda_rca24_fa364_y2;
  wire f_s_dadda_rca24_fa364_y3;
  wire f_s_dadda_rca24_fa364_y4;
  wire f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa364_y4;
  wire f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa363_y4;
  wire f_s_dadda_rca24_fa365_y0;
  wire f_s_dadda_rca24_fa365_y1;
  wire f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa201_y2;
  wire f_s_dadda_rca24_fa365_y2;
  wire f_s_dadda_rca24_fa365_y3;
  wire f_s_dadda_rca24_fa365_y4;
  wire f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa202_y2;
  wire f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa203_y2;
  wire f_s_dadda_rca24_fa366_y0;
  wire f_s_dadda_rca24_fa366_y1;
  wire f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa204_y2;
  wire f_s_dadda_rca24_fa366_y2;
  wire f_s_dadda_rca24_fa366_y3;
  wire f_s_dadda_rca24_fa366_y4;
  wire f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa366_y4;
  wire f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa365_y4;
  wire f_s_dadda_rca24_fa367_y0;
  wire f_s_dadda_rca24_fa367_y1;
  wire f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa214_y2;
  wire f_s_dadda_rca24_fa367_y2;
  wire f_s_dadda_rca24_fa367_y3;
  wire f_s_dadda_rca24_fa367_y4;
  wire f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa215_y2;
  wire f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa216_y2;
  wire f_s_dadda_rca24_fa368_y0;
  wire f_s_dadda_rca24_fa368_y1;
  wire f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa217_y2;
  wire f_s_dadda_rca24_fa368_y2;
  wire f_s_dadda_rca24_fa368_y3;
  wire f_s_dadda_rca24_fa368_y4;
  wire f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa368_y4;
  wire f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa367_y4;
  wire f_s_dadda_rca24_fa369_y0;
  wire f_s_dadda_rca24_fa369_y1;
  wire f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa227_y2;
  wire f_s_dadda_rca24_fa369_y2;
  wire f_s_dadda_rca24_fa369_y3;
  wire f_s_dadda_rca24_fa369_y4;
  wire f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa228_y2;
  wire f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa229_y2;
  wire f_s_dadda_rca24_fa370_y0;
  wire f_s_dadda_rca24_fa370_y1;
  wire f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa230_y2;
  wire f_s_dadda_rca24_fa370_y2;
  wire f_s_dadda_rca24_fa370_y3;
  wire f_s_dadda_rca24_fa370_y4;
  wire f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa370_y4;
  wire f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa369_y4;
  wire f_s_dadda_rca24_fa371_y0;
  wire f_s_dadda_rca24_fa371_y1;
  wire f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa240_y2;
  wire f_s_dadda_rca24_fa371_y2;
  wire f_s_dadda_rca24_fa371_y3;
  wire f_s_dadda_rca24_fa371_y4;
  wire f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa241_y2;
  wire f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa242_y2;
  wire f_s_dadda_rca24_fa372_y0;
  wire f_s_dadda_rca24_fa372_y1;
  wire f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa243_y2;
  wire f_s_dadda_rca24_fa372_y2;
  wire f_s_dadda_rca24_fa372_y3;
  wire f_s_dadda_rca24_fa372_y4;
  wire f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa372_y4;
  wire f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa371_y4;
  wire f_s_dadda_rca24_fa373_y0;
  wire f_s_dadda_rca24_fa373_y1;
  wire f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa252_y2;
  wire f_s_dadda_rca24_fa373_y2;
  wire f_s_dadda_rca24_fa373_y3;
  wire f_s_dadda_rca24_fa373_y4;
  wire f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa253_y2;
  wire f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa254_y2;
  wire f_s_dadda_rca24_fa374_y0;
  wire f_s_dadda_rca24_fa374_y1;
  wire f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa255_y2;
  wire f_s_dadda_rca24_fa374_y2;
  wire f_s_dadda_rca24_fa374_y3;
  wire f_s_dadda_rca24_fa374_y4;
  wire f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa374_y4;
  wire f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa373_y4;
  wire f_s_dadda_rca24_fa375_y0;
  wire f_s_dadda_rca24_fa375_y1;
  wire f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa263_y2;
  wire f_s_dadda_rca24_fa375_y2;
  wire f_s_dadda_rca24_fa375_y3;
  wire f_s_dadda_rca24_fa375_y4;
  wire f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa264_y2;
  wire f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa265_y2;
  wire f_s_dadda_rca24_fa376_y0;
  wire f_s_dadda_rca24_fa376_y1;
  wire f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa266_y2;
  wire f_s_dadda_rca24_fa376_y2;
  wire f_s_dadda_rca24_fa376_y3;
  wire f_s_dadda_rca24_fa376_y4;
  wire f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa376_y4;
  wire f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa375_y4;
  wire f_s_dadda_rca24_fa377_y0;
  wire f_s_dadda_rca24_fa377_y1;
  wire f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa273_y2;
  wire f_s_dadda_rca24_fa377_y2;
  wire f_s_dadda_rca24_fa377_y3;
  wire f_s_dadda_rca24_fa377_y4;
  wire f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa274_y2;
  wire f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa275_y2;
  wire f_s_dadda_rca24_fa378_y0;
  wire f_s_dadda_rca24_fa378_y1;
  wire f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa276_y2;
  wire f_s_dadda_rca24_fa378_y2;
  wire f_s_dadda_rca24_fa378_y3;
  wire f_s_dadda_rca24_fa378_y4;
  wire f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa378_y4;
  wire f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa377_y4;
  wire f_s_dadda_rca24_fa379_y0;
  wire f_s_dadda_rca24_fa379_y1;
  wire f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa282_y2;
  wire f_s_dadda_rca24_fa379_y2;
  wire f_s_dadda_rca24_fa379_y3;
  wire f_s_dadda_rca24_fa379_y4;
  wire f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa283_y2;
  wire f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa284_y2;
  wire f_s_dadda_rca24_fa380_y0;
  wire f_s_dadda_rca24_fa380_y1;
  wire f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa285_y2;
  wire f_s_dadda_rca24_fa380_y2;
  wire f_s_dadda_rca24_fa380_y3;
  wire f_s_dadda_rca24_fa380_y4;
  wire f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa380_y4;
  wire f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa379_y4;
  wire f_s_dadda_rca24_fa381_y0;
  wire f_s_dadda_rca24_fa381_y1;
  wire f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa290_y2;
  wire f_s_dadda_rca24_fa381_y2;
  wire f_s_dadda_rca24_fa381_y3;
  wire f_s_dadda_rca24_fa381_y4;
  wire f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa291_y2;
  wire f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa292_y2;
  wire f_s_dadda_rca24_fa382_y0;
  wire f_s_dadda_rca24_fa382_y1;
  wire f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa293_y2;
  wire f_s_dadda_rca24_fa382_y2;
  wire f_s_dadda_rca24_fa382_y3;
  wire f_s_dadda_rca24_fa382_y4;
  wire f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa382_y4;
  wire f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa381_y4;
  wire f_s_dadda_rca24_fa383_y0;
  wire f_s_dadda_rca24_fa383_y1;
  wire f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa297_y2;
  wire f_s_dadda_rca24_fa383_y2;
  wire f_s_dadda_rca24_fa383_y3;
  wire f_s_dadda_rca24_fa383_y4;
  wire f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa298_y2;
  wire f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa299_y2;
  wire f_s_dadda_rca24_fa384_y0;
  wire f_s_dadda_rca24_fa384_y1;
  wire f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa300_y2;
  wire f_s_dadda_rca24_fa384_y2;
  wire f_s_dadda_rca24_fa384_y3;
  wire f_s_dadda_rca24_fa384_y4;
  wire f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa384_y4;
  wire f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa383_y4;
  wire f_s_dadda_rca24_fa385_y0;
  wire f_s_dadda_rca24_fa385_y1;
  wire f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa303_y2;
  wire f_s_dadda_rca24_fa385_y2;
  wire f_s_dadda_rca24_fa385_y3;
  wire f_s_dadda_rca24_fa385_y4;
  wire f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa304_y2;
  wire f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa305_y2;
  wire f_s_dadda_rca24_fa386_y0;
  wire f_s_dadda_rca24_fa386_y1;
  wire f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa306_y2;
  wire f_s_dadda_rca24_fa386_y2;
  wire f_s_dadda_rca24_fa386_y3;
  wire f_s_dadda_rca24_fa386_y4;
  wire f_s_dadda_rca24_nand_14_23_a_14;
  wire f_s_dadda_rca24_nand_14_23_b_23;
  wire f_s_dadda_rca24_nand_14_23_y0;
  wire f_s_dadda_rca24_fa387_f_s_dadda_rca24_fa386_y4;
  wire f_s_dadda_rca24_fa387_f_s_dadda_rca24_fa385_y4;
  wire f_s_dadda_rca24_fa387_y0;
  wire f_s_dadda_rca24_fa387_y1;
  wire f_s_dadda_rca24_fa387_f_s_dadda_rca24_nand_14_23_y0;
  wire f_s_dadda_rca24_fa387_y2;
  wire f_s_dadda_rca24_fa387_y3;
  wire f_s_dadda_rca24_fa387_y4;
  wire f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa309_y2;
  wire f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa310_y2;
  wire f_s_dadda_rca24_fa388_y0;
  wire f_s_dadda_rca24_fa388_y1;
  wire f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa311_y2;
  wire f_s_dadda_rca24_fa388_y2;
  wire f_s_dadda_rca24_fa388_y3;
  wire f_s_dadda_rca24_fa388_y4;
  wire f_s_dadda_rca24_and_16_22_a_16;
  wire f_s_dadda_rca24_and_16_22_b_22;
  wire f_s_dadda_rca24_and_16_22_y0;
  wire f_s_dadda_rca24_fa389_f_s_dadda_rca24_fa388_y4;
  wire f_s_dadda_rca24_fa389_f_s_dadda_rca24_fa387_y4;
  wire f_s_dadda_rca24_fa389_y0;
  wire f_s_dadda_rca24_fa389_y1;
  wire f_s_dadda_rca24_fa389_f_s_dadda_rca24_and_16_22_y0;
  wire f_s_dadda_rca24_fa389_y2;
  wire f_s_dadda_rca24_fa389_y3;
  wire f_s_dadda_rca24_fa389_y4;
  wire f_s_dadda_rca24_nand_15_23_a_15;
  wire f_s_dadda_rca24_nand_15_23_b_23;
  wire f_s_dadda_rca24_nand_15_23_y0;
  wire f_s_dadda_rca24_fa390_f_s_dadda_rca24_nand_15_23_y0;
  wire f_s_dadda_rca24_fa390_f_s_dadda_rca24_fa314_y2;
  wire f_s_dadda_rca24_fa390_y0;
  wire f_s_dadda_rca24_fa390_y1;
  wire f_s_dadda_rca24_fa390_f_s_dadda_rca24_fa315_y2;
  wire f_s_dadda_rca24_fa390_y2;
  wire f_s_dadda_rca24_fa390_y3;
  wire f_s_dadda_rca24_fa390_y4;
  wire f_s_dadda_rca24_and_18_21_a_18;
  wire f_s_dadda_rca24_and_18_21_b_21;
  wire f_s_dadda_rca24_and_18_21_y0;
  wire f_s_dadda_rca24_fa391_f_s_dadda_rca24_fa390_y4;
  wire f_s_dadda_rca24_fa391_f_s_dadda_rca24_fa389_y4;
  wire f_s_dadda_rca24_fa391_y0;
  wire f_s_dadda_rca24_fa391_y1;
  wire f_s_dadda_rca24_fa391_f_s_dadda_rca24_and_18_21_y0;
  wire f_s_dadda_rca24_fa391_y2;
  wire f_s_dadda_rca24_fa391_y3;
  wire f_s_dadda_rca24_fa391_y4;
  wire f_s_dadda_rca24_and_17_22_a_17;
  wire f_s_dadda_rca24_and_17_22_b_22;
  wire f_s_dadda_rca24_and_17_22_y0;
  wire f_s_dadda_rca24_nand_16_23_a_16;
  wire f_s_dadda_rca24_nand_16_23_b_23;
  wire f_s_dadda_rca24_nand_16_23_y0;
  wire f_s_dadda_rca24_fa392_f_s_dadda_rca24_and_17_22_y0;
  wire f_s_dadda_rca24_fa392_f_s_dadda_rca24_nand_16_23_y0;
  wire f_s_dadda_rca24_fa392_y0;
  wire f_s_dadda_rca24_fa392_y1;
  wire f_s_dadda_rca24_fa392_f_s_dadda_rca24_fa318_y2;
  wire f_s_dadda_rca24_fa392_y2;
  wire f_s_dadda_rca24_fa392_y3;
  wire f_s_dadda_rca24_fa392_y4;
  wire f_s_dadda_rca24_and_20_20_a_20;
  wire f_s_dadda_rca24_and_20_20_b_20;
  wire f_s_dadda_rca24_and_20_20_y0;
  wire f_s_dadda_rca24_fa393_f_s_dadda_rca24_fa392_y4;
  wire f_s_dadda_rca24_fa393_f_s_dadda_rca24_fa391_y4;
  wire f_s_dadda_rca24_fa393_y0;
  wire f_s_dadda_rca24_fa393_y1;
  wire f_s_dadda_rca24_fa393_f_s_dadda_rca24_and_20_20_y0;
  wire f_s_dadda_rca24_fa393_y2;
  wire f_s_dadda_rca24_fa393_y3;
  wire f_s_dadda_rca24_fa393_y4;
  wire f_s_dadda_rca24_and_19_21_a_19;
  wire f_s_dadda_rca24_and_19_21_b_21;
  wire f_s_dadda_rca24_and_19_21_y0;
  wire f_s_dadda_rca24_and_18_22_a_18;
  wire f_s_dadda_rca24_and_18_22_b_22;
  wire f_s_dadda_rca24_and_18_22_y0;
  wire f_s_dadda_rca24_nand_17_23_a_17;
  wire f_s_dadda_rca24_nand_17_23_b_23;
  wire f_s_dadda_rca24_nand_17_23_y0;
  wire f_s_dadda_rca24_fa394_f_s_dadda_rca24_and_19_21_y0;
  wire f_s_dadda_rca24_fa394_f_s_dadda_rca24_and_18_22_y0;
  wire f_s_dadda_rca24_fa394_y0;
  wire f_s_dadda_rca24_fa394_y1;
  wire f_s_dadda_rca24_fa394_f_s_dadda_rca24_nand_17_23_y0;
  wire f_s_dadda_rca24_fa394_y2;
  wire f_s_dadda_rca24_fa394_y3;
  wire f_s_dadda_rca24_fa394_y4;
  wire f_s_dadda_rca24_and_22_19_a_22;
  wire f_s_dadda_rca24_and_22_19_b_19;
  wire f_s_dadda_rca24_and_22_19_y0;
  wire f_s_dadda_rca24_fa395_f_s_dadda_rca24_fa394_y4;
  wire f_s_dadda_rca24_fa395_f_s_dadda_rca24_fa393_y4;
  wire f_s_dadda_rca24_fa395_y0;
  wire f_s_dadda_rca24_fa395_y1;
  wire f_s_dadda_rca24_fa395_f_s_dadda_rca24_and_22_19_y0;
  wire f_s_dadda_rca24_fa395_y2;
  wire f_s_dadda_rca24_fa395_y3;
  wire f_s_dadda_rca24_fa395_y4;
  wire f_s_dadda_rca24_and_21_20_a_21;
  wire f_s_dadda_rca24_and_21_20_b_20;
  wire f_s_dadda_rca24_and_21_20_y0;
  wire f_s_dadda_rca24_and_20_21_a_20;
  wire f_s_dadda_rca24_and_20_21_b_21;
  wire f_s_dadda_rca24_and_20_21_y0;
  wire f_s_dadda_rca24_and_19_22_a_19;
  wire f_s_dadda_rca24_and_19_22_b_22;
  wire f_s_dadda_rca24_and_19_22_y0;
  wire f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_21_20_y0;
  wire f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_20_21_y0;
  wire f_s_dadda_rca24_fa396_y0;
  wire f_s_dadda_rca24_fa396_y1;
  wire f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_19_22_y0;
  wire f_s_dadda_rca24_fa396_y2;
  wire f_s_dadda_rca24_fa396_y3;
  wire f_s_dadda_rca24_fa396_y4;
  wire f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa396_y4;
  wire f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa395_y4;
  wire f_s_dadda_rca24_fa397_y0;
  wire f_s_dadda_rca24_fa397_y1;
  wire f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa323_y4;
  wire f_s_dadda_rca24_fa397_y2;
  wire f_s_dadda_rca24_fa397_y3;
  wire f_s_dadda_rca24_fa397_y4;
  wire f_s_dadda_rca24_nand_23_19_a_23;
  wire f_s_dadda_rca24_nand_23_19_b_19;
  wire f_s_dadda_rca24_nand_23_19_y0;
  wire f_s_dadda_rca24_and_22_20_a_22;
  wire f_s_dadda_rca24_and_22_20_b_20;
  wire f_s_dadda_rca24_and_22_20_y0;
  wire f_s_dadda_rca24_and_21_21_a_21;
  wire f_s_dadda_rca24_and_21_21_b_21;
  wire f_s_dadda_rca24_and_21_21_y0;
  wire f_s_dadda_rca24_fa398_f_s_dadda_rca24_nand_23_19_y0;
  wire f_s_dadda_rca24_fa398_f_s_dadda_rca24_and_22_20_y0;
  wire f_s_dadda_rca24_fa398_y0;
  wire f_s_dadda_rca24_fa398_y1;
  wire f_s_dadda_rca24_fa398_f_s_dadda_rca24_and_21_21_y0;
  wire f_s_dadda_rca24_fa398_y2;
  wire f_s_dadda_rca24_fa398_y3;
  wire f_s_dadda_rca24_fa398_y4;
  wire f_s_dadda_rca24_nand_23_20_a_23;
  wire f_s_dadda_rca24_nand_23_20_b_20;
  wire f_s_dadda_rca24_nand_23_20_y0;
  wire f_s_dadda_rca24_fa399_f_s_dadda_rca24_fa398_y4;
  wire f_s_dadda_rca24_fa399_f_s_dadda_rca24_fa397_y4;
  wire f_s_dadda_rca24_fa399_y0;
  wire f_s_dadda_rca24_fa399_y1;
  wire f_s_dadda_rca24_fa399_f_s_dadda_rca24_nand_23_20_y0;
  wire f_s_dadda_rca24_fa399_y2;
  wire f_s_dadda_rca24_fa399_y3;
  wire f_s_dadda_rca24_fa399_y4;
  wire f_s_dadda_rca24_and_3_0_a_3;
  wire f_s_dadda_rca24_and_3_0_b_0;
  wire f_s_dadda_rca24_and_3_0_y0;
  wire f_s_dadda_rca24_and_2_1_a_2;
  wire f_s_dadda_rca24_and_2_1_b_1;
  wire f_s_dadda_rca24_and_2_1_y0;
  wire f_s_dadda_rca24_ha20_f_s_dadda_rca24_and_3_0_y0;
  wire f_s_dadda_rca24_ha20_f_s_dadda_rca24_and_2_1_y0;
  wire f_s_dadda_rca24_ha20_y0;
  wire f_s_dadda_rca24_ha20_y1;
  wire f_s_dadda_rca24_and_2_2_a_2;
  wire f_s_dadda_rca24_and_2_2_b_2;
  wire f_s_dadda_rca24_and_2_2_y0;
  wire f_s_dadda_rca24_and_1_3_a_1;
  wire f_s_dadda_rca24_and_1_3_b_3;
  wire f_s_dadda_rca24_and_1_3_y0;
  wire f_s_dadda_rca24_fa400_f_s_dadda_rca24_ha20_y1;
  wire f_s_dadda_rca24_fa400_f_s_dadda_rca24_and_2_2_y0;
  wire f_s_dadda_rca24_fa400_y0;
  wire f_s_dadda_rca24_fa400_y1;
  wire f_s_dadda_rca24_fa400_f_s_dadda_rca24_and_1_3_y0;
  wire f_s_dadda_rca24_fa400_y2;
  wire f_s_dadda_rca24_fa400_y3;
  wire f_s_dadda_rca24_fa400_y4;
  wire f_s_dadda_rca24_and_1_4_a_1;
  wire f_s_dadda_rca24_and_1_4_b_4;
  wire f_s_dadda_rca24_and_1_4_y0;
  wire f_s_dadda_rca24_and_0_5_a_0;
  wire f_s_dadda_rca24_and_0_5_b_5;
  wire f_s_dadda_rca24_and_0_5_y0;
  wire f_s_dadda_rca24_fa401_f_s_dadda_rca24_fa400_y4;
  wire f_s_dadda_rca24_fa401_f_s_dadda_rca24_and_1_4_y0;
  wire f_s_dadda_rca24_fa401_y0;
  wire f_s_dadda_rca24_fa401_y1;
  wire f_s_dadda_rca24_fa401_f_s_dadda_rca24_and_0_5_y0;
  wire f_s_dadda_rca24_fa401_y2;
  wire f_s_dadda_rca24_fa401_y3;
  wire f_s_dadda_rca24_fa401_y4;
  wire f_s_dadda_rca24_and_0_6_a_0;
  wire f_s_dadda_rca24_and_0_6_b_6;
  wire f_s_dadda_rca24_and_0_6_y0;
  wire f_s_dadda_rca24_fa402_f_s_dadda_rca24_fa401_y4;
  wire f_s_dadda_rca24_fa402_f_s_dadda_rca24_and_0_6_y0;
  wire f_s_dadda_rca24_fa402_y0;
  wire f_s_dadda_rca24_fa402_y1;
  wire f_s_dadda_rca24_fa402_f_s_dadda_rca24_ha5_y0;
  wire f_s_dadda_rca24_fa402_y2;
  wire f_s_dadda_rca24_fa402_y3;
  wire f_s_dadda_rca24_fa402_y4;
  wire f_s_dadda_rca24_fa403_f_s_dadda_rca24_fa402_y4;
  wire f_s_dadda_rca24_fa403_f_s_dadda_rca24_fa25_y2;
  wire f_s_dadda_rca24_fa403_y0;
  wire f_s_dadda_rca24_fa403_y1;
  wire f_s_dadda_rca24_fa403_f_s_dadda_rca24_ha6_y0;
  wire f_s_dadda_rca24_fa403_y2;
  wire f_s_dadda_rca24_fa403_y3;
  wire f_s_dadda_rca24_fa403_y4;
  wire f_s_dadda_rca24_fa404_f_s_dadda_rca24_fa403_y4;
  wire f_s_dadda_rca24_fa404_f_s_dadda_rca24_fa27_y2;
  wire f_s_dadda_rca24_fa404_y0;
  wire f_s_dadda_rca24_fa404_y1;
  wire f_s_dadda_rca24_fa404_f_s_dadda_rca24_ha7_y0;
  wire f_s_dadda_rca24_fa404_y2;
  wire f_s_dadda_rca24_fa404_y3;
  wire f_s_dadda_rca24_fa404_y4;
  wire f_s_dadda_rca24_fa405_f_s_dadda_rca24_fa404_y4;
  wire f_s_dadda_rca24_fa405_f_s_dadda_rca24_fa30_y2;
  wire f_s_dadda_rca24_fa405_y0;
  wire f_s_dadda_rca24_fa405_y1;
  wire f_s_dadda_rca24_fa405_f_s_dadda_rca24_ha8_y0;
  wire f_s_dadda_rca24_fa405_y2;
  wire f_s_dadda_rca24_fa405_y3;
  wire f_s_dadda_rca24_fa405_y4;
  wire f_s_dadda_rca24_fa406_f_s_dadda_rca24_fa405_y4;
  wire f_s_dadda_rca24_fa406_f_s_dadda_rca24_fa34_y2;
  wire f_s_dadda_rca24_fa406_y0;
  wire f_s_dadda_rca24_fa406_y1;
  wire f_s_dadda_rca24_fa406_f_s_dadda_rca24_ha9_y0;
  wire f_s_dadda_rca24_fa406_y2;
  wire f_s_dadda_rca24_fa406_y3;
  wire f_s_dadda_rca24_fa406_y4;
  wire f_s_dadda_rca24_fa407_f_s_dadda_rca24_fa406_y4;
  wire f_s_dadda_rca24_fa407_f_s_dadda_rca24_fa39_y2;
  wire f_s_dadda_rca24_fa407_y0;
  wire f_s_dadda_rca24_fa407_y1;
  wire f_s_dadda_rca24_fa407_f_s_dadda_rca24_ha10_y0;
  wire f_s_dadda_rca24_fa407_y2;
  wire f_s_dadda_rca24_fa407_y3;
  wire f_s_dadda_rca24_fa407_y4;
  wire f_s_dadda_rca24_fa408_f_s_dadda_rca24_fa407_y4;
  wire f_s_dadda_rca24_fa408_f_s_dadda_rca24_fa45_y2;
  wire f_s_dadda_rca24_fa408_y0;
  wire f_s_dadda_rca24_fa408_y1;
  wire f_s_dadda_rca24_fa408_f_s_dadda_rca24_ha11_y0;
  wire f_s_dadda_rca24_fa408_y2;
  wire f_s_dadda_rca24_fa408_y3;
  wire f_s_dadda_rca24_fa408_y4;
  wire f_s_dadda_rca24_fa409_f_s_dadda_rca24_fa408_y4;
  wire f_s_dadda_rca24_fa409_f_s_dadda_rca24_fa52_y2;
  wire f_s_dadda_rca24_fa409_y0;
  wire f_s_dadda_rca24_fa409_y1;
  wire f_s_dadda_rca24_fa409_f_s_dadda_rca24_ha12_y0;
  wire f_s_dadda_rca24_fa409_y2;
  wire f_s_dadda_rca24_fa409_y3;
  wire f_s_dadda_rca24_fa409_y4;
  wire f_s_dadda_rca24_fa410_f_s_dadda_rca24_fa409_y4;
  wire f_s_dadda_rca24_fa410_f_s_dadda_rca24_fa60_y2;
  wire f_s_dadda_rca24_fa410_y0;
  wire f_s_dadda_rca24_fa410_y1;
  wire f_s_dadda_rca24_fa410_f_s_dadda_rca24_ha13_y0;
  wire f_s_dadda_rca24_fa410_y2;
  wire f_s_dadda_rca24_fa410_y3;
  wire f_s_dadda_rca24_fa410_y4;
  wire f_s_dadda_rca24_fa411_f_s_dadda_rca24_fa410_y4;
  wire f_s_dadda_rca24_fa411_f_s_dadda_rca24_fa69_y2;
  wire f_s_dadda_rca24_fa411_y0;
  wire f_s_dadda_rca24_fa411_y1;
  wire f_s_dadda_rca24_fa411_f_s_dadda_rca24_ha14_y0;
  wire f_s_dadda_rca24_fa411_y2;
  wire f_s_dadda_rca24_fa411_y3;
  wire f_s_dadda_rca24_fa411_y4;
  wire f_s_dadda_rca24_fa412_f_s_dadda_rca24_fa411_y4;
  wire f_s_dadda_rca24_fa412_f_s_dadda_rca24_fa79_y2;
  wire f_s_dadda_rca24_fa412_y0;
  wire f_s_dadda_rca24_fa412_y1;
  wire f_s_dadda_rca24_fa412_f_s_dadda_rca24_ha15_y0;
  wire f_s_dadda_rca24_fa412_y2;
  wire f_s_dadda_rca24_fa412_y3;
  wire f_s_dadda_rca24_fa412_y4;
  wire f_s_dadda_rca24_fa413_f_s_dadda_rca24_fa412_y4;
  wire f_s_dadda_rca24_fa413_f_s_dadda_rca24_fa90_y2;
  wire f_s_dadda_rca24_fa413_y0;
  wire f_s_dadda_rca24_fa413_y1;
  wire f_s_dadda_rca24_fa413_f_s_dadda_rca24_ha16_y0;
  wire f_s_dadda_rca24_fa413_y2;
  wire f_s_dadda_rca24_fa413_y3;
  wire f_s_dadda_rca24_fa413_y4;
  wire f_s_dadda_rca24_fa414_f_s_dadda_rca24_fa413_y4;
  wire f_s_dadda_rca24_fa414_f_s_dadda_rca24_fa102_y2;
  wire f_s_dadda_rca24_fa414_y0;
  wire f_s_dadda_rca24_fa414_y1;
  wire f_s_dadda_rca24_fa414_f_s_dadda_rca24_ha17_y0;
  wire f_s_dadda_rca24_fa414_y2;
  wire f_s_dadda_rca24_fa414_y3;
  wire f_s_dadda_rca24_fa414_y4;
  wire f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa414_y4;
  wire f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa114_y2;
  wire f_s_dadda_rca24_fa415_y0;
  wire f_s_dadda_rca24_fa415_y1;
  wire f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa115_y2;
  wire f_s_dadda_rca24_fa415_y2;
  wire f_s_dadda_rca24_fa415_y3;
  wire f_s_dadda_rca24_fa415_y4;
  wire f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa415_y4;
  wire f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa127_y2;
  wire f_s_dadda_rca24_fa416_y0;
  wire f_s_dadda_rca24_fa416_y1;
  wire f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa128_y2;
  wire f_s_dadda_rca24_fa416_y2;
  wire f_s_dadda_rca24_fa416_y3;
  wire f_s_dadda_rca24_fa416_y4;
  wire f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa416_y4;
  wire f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa140_y2;
  wire f_s_dadda_rca24_fa417_y0;
  wire f_s_dadda_rca24_fa417_y1;
  wire f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa141_y2;
  wire f_s_dadda_rca24_fa417_y2;
  wire f_s_dadda_rca24_fa417_y3;
  wire f_s_dadda_rca24_fa417_y4;
  wire f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa417_y4;
  wire f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa153_y2;
  wire f_s_dadda_rca24_fa418_y0;
  wire f_s_dadda_rca24_fa418_y1;
  wire f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa154_y2;
  wire f_s_dadda_rca24_fa418_y2;
  wire f_s_dadda_rca24_fa418_y3;
  wire f_s_dadda_rca24_fa418_y4;
  wire f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa418_y4;
  wire f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa166_y2;
  wire f_s_dadda_rca24_fa419_y0;
  wire f_s_dadda_rca24_fa419_y1;
  wire f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa167_y2;
  wire f_s_dadda_rca24_fa419_y2;
  wire f_s_dadda_rca24_fa419_y3;
  wire f_s_dadda_rca24_fa419_y4;
  wire f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa419_y4;
  wire f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa179_y2;
  wire f_s_dadda_rca24_fa420_y0;
  wire f_s_dadda_rca24_fa420_y1;
  wire f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa180_y2;
  wire f_s_dadda_rca24_fa420_y2;
  wire f_s_dadda_rca24_fa420_y3;
  wire f_s_dadda_rca24_fa420_y4;
  wire f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa420_y4;
  wire f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa192_y2;
  wire f_s_dadda_rca24_fa421_y0;
  wire f_s_dadda_rca24_fa421_y1;
  wire f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa193_y2;
  wire f_s_dadda_rca24_fa421_y2;
  wire f_s_dadda_rca24_fa421_y3;
  wire f_s_dadda_rca24_fa421_y4;
  wire f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa421_y4;
  wire f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa205_y2;
  wire f_s_dadda_rca24_fa422_y0;
  wire f_s_dadda_rca24_fa422_y1;
  wire f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa206_y2;
  wire f_s_dadda_rca24_fa422_y2;
  wire f_s_dadda_rca24_fa422_y3;
  wire f_s_dadda_rca24_fa422_y4;
  wire f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa422_y4;
  wire f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa218_y2;
  wire f_s_dadda_rca24_fa423_y0;
  wire f_s_dadda_rca24_fa423_y1;
  wire f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa219_y2;
  wire f_s_dadda_rca24_fa423_y2;
  wire f_s_dadda_rca24_fa423_y3;
  wire f_s_dadda_rca24_fa423_y4;
  wire f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa423_y4;
  wire f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa231_y2;
  wire f_s_dadda_rca24_fa424_y0;
  wire f_s_dadda_rca24_fa424_y1;
  wire f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa232_y2;
  wire f_s_dadda_rca24_fa424_y2;
  wire f_s_dadda_rca24_fa424_y3;
  wire f_s_dadda_rca24_fa424_y4;
  wire f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa424_y4;
  wire f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa244_y2;
  wire f_s_dadda_rca24_fa425_y0;
  wire f_s_dadda_rca24_fa425_y1;
  wire f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa245_y2;
  wire f_s_dadda_rca24_fa425_y2;
  wire f_s_dadda_rca24_fa425_y3;
  wire f_s_dadda_rca24_fa425_y4;
  wire f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa425_y4;
  wire f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa256_y2;
  wire f_s_dadda_rca24_fa426_y0;
  wire f_s_dadda_rca24_fa426_y1;
  wire f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa257_y2;
  wire f_s_dadda_rca24_fa426_y2;
  wire f_s_dadda_rca24_fa426_y3;
  wire f_s_dadda_rca24_fa426_y4;
  wire f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa426_y4;
  wire f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa267_y2;
  wire f_s_dadda_rca24_fa427_y0;
  wire f_s_dadda_rca24_fa427_y1;
  wire f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa268_y2;
  wire f_s_dadda_rca24_fa427_y2;
  wire f_s_dadda_rca24_fa427_y3;
  wire f_s_dadda_rca24_fa427_y4;
  wire f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa427_y4;
  wire f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa277_y2;
  wire f_s_dadda_rca24_fa428_y0;
  wire f_s_dadda_rca24_fa428_y1;
  wire f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa278_y2;
  wire f_s_dadda_rca24_fa428_y2;
  wire f_s_dadda_rca24_fa428_y3;
  wire f_s_dadda_rca24_fa428_y4;
  wire f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa428_y4;
  wire f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa286_y2;
  wire f_s_dadda_rca24_fa429_y0;
  wire f_s_dadda_rca24_fa429_y1;
  wire f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa287_y2;
  wire f_s_dadda_rca24_fa429_y2;
  wire f_s_dadda_rca24_fa429_y3;
  wire f_s_dadda_rca24_fa429_y4;
  wire f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa429_y4;
  wire f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa294_y2;
  wire f_s_dadda_rca24_fa430_y0;
  wire f_s_dadda_rca24_fa430_y1;
  wire f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa295_y2;
  wire f_s_dadda_rca24_fa430_y2;
  wire f_s_dadda_rca24_fa430_y3;
  wire f_s_dadda_rca24_fa430_y4;
  wire f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa430_y4;
  wire f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa301_y2;
  wire f_s_dadda_rca24_fa431_y0;
  wire f_s_dadda_rca24_fa431_y1;
  wire f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa302_y2;
  wire f_s_dadda_rca24_fa431_y2;
  wire f_s_dadda_rca24_fa431_y3;
  wire f_s_dadda_rca24_fa431_y4;
  wire f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa431_y4;
  wire f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa307_y2;
  wire f_s_dadda_rca24_fa432_y0;
  wire f_s_dadda_rca24_fa432_y1;
  wire f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa308_y2;
  wire f_s_dadda_rca24_fa432_y2;
  wire f_s_dadda_rca24_fa432_y3;
  wire f_s_dadda_rca24_fa432_y4;
  wire f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa432_y4;
  wire f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa312_y2;
  wire f_s_dadda_rca24_fa433_y0;
  wire f_s_dadda_rca24_fa433_y1;
  wire f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa313_y2;
  wire f_s_dadda_rca24_fa433_y2;
  wire f_s_dadda_rca24_fa433_y3;
  wire f_s_dadda_rca24_fa433_y4;
  wire f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa433_y4;
  wire f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa316_y2;
  wire f_s_dadda_rca24_fa434_y0;
  wire f_s_dadda_rca24_fa434_y1;
  wire f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa317_y2;
  wire f_s_dadda_rca24_fa434_y2;
  wire f_s_dadda_rca24_fa434_y3;
  wire f_s_dadda_rca24_fa434_y4;
  wire f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa434_y4;
  wire f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa319_y2;
  wire f_s_dadda_rca24_fa435_y0;
  wire f_s_dadda_rca24_fa435_y1;
  wire f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa320_y2;
  wire f_s_dadda_rca24_fa435_y2;
  wire f_s_dadda_rca24_fa435_y3;
  wire f_s_dadda_rca24_fa435_y4;
  wire f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa435_y4;
  wire f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa321_y2;
  wire f_s_dadda_rca24_fa436_y0;
  wire f_s_dadda_rca24_fa436_y1;
  wire f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa322_y2;
  wire f_s_dadda_rca24_fa436_y2;
  wire f_s_dadda_rca24_fa436_y3;
  wire f_s_dadda_rca24_fa436_y4;
  wire f_s_dadda_rca24_nand_18_23_a_18;
  wire f_s_dadda_rca24_nand_18_23_b_23;
  wire f_s_dadda_rca24_nand_18_23_y0;
  wire f_s_dadda_rca24_fa437_f_s_dadda_rca24_fa436_y4;
  wire f_s_dadda_rca24_fa437_f_s_dadda_rca24_nand_18_23_y0;
  wire f_s_dadda_rca24_fa437_y0;
  wire f_s_dadda_rca24_fa437_y1;
  wire f_s_dadda_rca24_fa437_f_s_dadda_rca24_fa323_y2;
  wire f_s_dadda_rca24_fa437_y2;
  wire f_s_dadda_rca24_fa437_y3;
  wire f_s_dadda_rca24_fa437_y4;
  wire f_s_dadda_rca24_and_20_22_a_20;
  wire f_s_dadda_rca24_and_20_22_b_22;
  wire f_s_dadda_rca24_and_20_22_y0;
  wire f_s_dadda_rca24_nand_19_23_a_19;
  wire f_s_dadda_rca24_nand_19_23_b_23;
  wire f_s_dadda_rca24_nand_19_23_y0;
  wire f_s_dadda_rca24_fa438_f_s_dadda_rca24_fa437_y4;
  wire f_s_dadda_rca24_fa438_f_s_dadda_rca24_and_20_22_y0;
  wire f_s_dadda_rca24_fa438_y0;
  wire f_s_dadda_rca24_fa438_y1;
  wire f_s_dadda_rca24_fa438_f_s_dadda_rca24_nand_19_23_y0;
  wire f_s_dadda_rca24_fa438_y2;
  wire f_s_dadda_rca24_fa438_y3;
  wire f_s_dadda_rca24_fa438_y4;
  wire f_s_dadda_rca24_and_22_21_a_22;
  wire f_s_dadda_rca24_and_22_21_b_21;
  wire f_s_dadda_rca24_and_22_21_y0;
  wire f_s_dadda_rca24_and_21_22_a_21;
  wire f_s_dadda_rca24_and_21_22_b_22;
  wire f_s_dadda_rca24_and_21_22_y0;
  wire f_s_dadda_rca24_fa439_f_s_dadda_rca24_fa438_y4;
  wire f_s_dadda_rca24_fa439_f_s_dadda_rca24_and_22_21_y0;
  wire f_s_dadda_rca24_fa439_y0;
  wire f_s_dadda_rca24_fa439_y1;
  wire f_s_dadda_rca24_fa439_f_s_dadda_rca24_and_21_22_y0;
  wire f_s_dadda_rca24_fa439_y2;
  wire f_s_dadda_rca24_fa439_y3;
  wire f_s_dadda_rca24_fa439_y4;
  wire f_s_dadda_rca24_nand_23_21_a_23;
  wire f_s_dadda_rca24_nand_23_21_b_21;
  wire f_s_dadda_rca24_nand_23_21_y0;
  wire f_s_dadda_rca24_fa440_f_s_dadda_rca24_fa439_y4;
  wire f_s_dadda_rca24_fa440_f_s_dadda_rca24_fa399_y4;
  wire f_s_dadda_rca24_fa440_y0;
  wire f_s_dadda_rca24_fa440_y1;
  wire f_s_dadda_rca24_fa440_f_s_dadda_rca24_nand_23_21_y0;
  wire f_s_dadda_rca24_fa440_y2;
  wire f_s_dadda_rca24_fa440_y3;
  wire f_s_dadda_rca24_fa440_y4;
  wire f_s_dadda_rca24_and_2_0_a_2;
  wire f_s_dadda_rca24_and_2_0_b_0;
  wire f_s_dadda_rca24_and_2_0_y0;
  wire f_s_dadda_rca24_and_1_1_a_1;
  wire f_s_dadda_rca24_and_1_1_b_1;
  wire f_s_dadda_rca24_and_1_1_y0;
  wire f_s_dadda_rca24_ha21_f_s_dadda_rca24_and_2_0_y0;
  wire f_s_dadda_rca24_ha21_f_s_dadda_rca24_and_1_1_y0;
  wire f_s_dadda_rca24_ha21_y0;
  wire f_s_dadda_rca24_ha21_y1;
  wire f_s_dadda_rca24_and_1_2_a_1;
  wire f_s_dadda_rca24_and_1_2_b_2;
  wire f_s_dadda_rca24_and_1_2_y0;
  wire f_s_dadda_rca24_and_0_3_a_0;
  wire f_s_dadda_rca24_and_0_3_b_3;
  wire f_s_dadda_rca24_and_0_3_y0;
  wire f_s_dadda_rca24_fa441_f_s_dadda_rca24_ha21_y1;
  wire f_s_dadda_rca24_fa441_f_s_dadda_rca24_and_1_2_y0;
  wire f_s_dadda_rca24_fa441_y0;
  wire f_s_dadda_rca24_fa441_y1;
  wire f_s_dadda_rca24_fa441_f_s_dadda_rca24_and_0_3_y0;
  wire f_s_dadda_rca24_fa441_y2;
  wire f_s_dadda_rca24_fa441_y3;
  wire f_s_dadda_rca24_fa441_y4;
  wire f_s_dadda_rca24_and_0_4_a_0;
  wire f_s_dadda_rca24_and_0_4_b_4;
  wire f_s_dadda_rca24_and_0_4_y0;
  wire f_s_dadda_rca24_fa442_f_s_dadda_rca24_fa441_y4;
  wire f_s_dadda_rca24_fa442_f_s_dadda_rca24_and_0_4_y0;
  wire f_s_dadda_rca24_fa442_y0;
  wire f_s_dadda_rca24_fa442_y1;
  wire f_s_dadda_rca24_fa442_f_s_dadda_rca24_ha18_y0;
  wire f_s_dadda_rca24_fa442_y2;
  wire f_s_dadda_rca24_fa442_y3;
  wire f_s_dadda_rca24_fa442_y4;
  wire f_s_dadda_rca24_fa443_f_s_dadda_rca24_fa442_y4;
  wire f_s_dadda_rca24_fa443_f_s_dadda_rca24_fa324_y2;
  wire f_s_dadda_rca24_fa443_y0;
  wire f_s_dadda_rca24_fa443_y1;
  wire f_s_dadda_rca24_fa443_f_s_dadda_rca24_ha19_y0;
  wire f_s_dadda_rca24_fa443_y2;
  wire f_s_dadda_rca24_fa443_y3;
  wire f_s_dadda_rca24_fa443_y4;
  wire f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa443_y4;
  wire f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa325_y2;
  wire f_s_dadda_rca24_fa444_y0;
  wire f_s_dadda_rca24_fa444_y1;
  wire f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa326_y2;
  wire f_s_dadda_rca24_fa444_y2;
  wire f_s_dadda_rca24_fa444_y3;
  wire f_s_dadda_rca24_fa444_y4;
  wire f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa444_y4;
  wire f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa327_y2;
  wire f_s_dadda_rca24_fa445_y0;
  wire f_s_dadda_rca24_fa445_y1;
  wire f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa328_y2;
  wire f_s_dadda_rca24_fa445_y2;
  wire f_s_dadda_rca24_fa445_y3;
  wire f_s_dadda_rca24_fa445_y4;
  wire f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa445_y4;
  wire f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa329_y2;
  wire f_s_dadda_rca24_fa446_y0;
  wire f_s_dadda_rca24_fa446_y1;
  wire f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa330_y2;
  wire f_s_dadda_rca24_fa446_y2;
  wire f_s_dadda_rca24_fa446_y3;
  wire f_s_dadda_rca24_fa446_y4;
  wire f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa446_y4;
  wire f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa331_y2;
  wire f_s_dadda_rca24_fa447_y0;
  wire f_s_dadda_rca24_fa447_y1;
  wire f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa332_y2;
  wire f_s_dadda_rca24_fa447_y2;
  wire f_s_dadda_rca24_fa447_y3;
  wire f_s_dadda_rca24_fa447_y4;
  wire f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa447_y4;
  wire f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa333_y2;
  wire f_s_dadda_rca24_fa448_y0;
  wire f_s_dadda_rca24_fa448_y1;
  wire f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa334_y2;
  wire f_s_dadda_rca24_fa448_y2;
  wire f_s_dadda_rca24_fa448_y3;
  wire f_s_dadda_rca24_fa448_y4;
  wire f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa448_y4;
  wire f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa335_y2;
  wire f_s_dadda_rca24_fa449_y0;
  wire f_s_dadda_rca24_fa449_y1;
  wire f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa336_y2;
  wire f_s_dadda_rca24_fa449_y2;
  wire f_s_dadda_rca24_fa449_y3;
  wire f_s_dadda_rca24_fa449_y4;
  wire f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa449_y4;
  wire f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa337_y2;
  wire f_s_dadda_rca24_fa450_y0;
  wire f_s_dadda_rca24_fa450_y1;
  wire f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa338_y2;
  wire f_s_dadda_rca24_fa450_y2;
  wire f_s_dadda_rca24_fa450_y3;
  wire f_s_dadda_rca24_fa450_y4;
  wire f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa450_y4;
  wire f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa339_y2;
  wire f_s_dadda_rca24_fa451_y0;
  wire f_s_dadda_rca24_fa451_y1;
  wire f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa340_y2;
  wire f_s_dadda_rca24_fa451_y2;
  wire f_s_dadda_rca24_fa451_y3;
  wire f_s_dadda_rca24_fa451_y4;
  wire f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa451_y4;
  wire f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa341_y2;
  wire f_s_dadda_rca24_fa452_y0;
  wire f_s_dadda_rca24_fa452_y1;
  wire f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa342_y2;
  wire f_s_dadda_rca24_fa452_y2;
  wire f_s_dadda_rca24_fa452_y3;
  wire f_s_dadda_rca24_fa452_y4;
  wire f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa452_y4;
  wire f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa343_y2;
  wire f_s_dadda_rca24_fa453_y0;
  wire f_s_dadda_rca24_fa453_y1;
  wire f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa344_y2;
  wire f_s_dadda_rca24_fa453_y2;
  wire f_s_dadda_rca24_fa453_y3;
  wire f_s_dadda_rca24_fa453_y4;
  wire f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa453_y4;
  wire f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa345_y2;
  wire f_s_dadda_rca24_fa454_y0;
  wire f_s_dadda_rca24_fa454_y1;
  wire f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa346_y2;
  wire f_s_dadda_rca24_fa454_y2;
  wire f_s_dadda_rca24_fa454_y3;
  wire f_s_dadda_rca24_fa454_y4;
  wire f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa454_y4;
  wire f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa347_y2;
  wire f_s_dadda_rca24_fa455_y0;
  wire f_s_dadda_rca24_fa455_y1;
  wire f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa348_y2;
  wire f_s_dadda_rca24_fa455_y2;
  wire f_s_dadda_rca24_fa455_y3;
  wire f_s_dadda_rca24_fa455_y4;
  wire f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa455_y4;
  wire f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa349_y2;
  wire f_s_dadda_rca24_fa456_y0;
  wire f_s_dadda_rca24_fa456_y1;
  wire f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa350_y2;
  wire f_s_dadda_rca24_fa456_y2;
  wire f_s_dadda_rca24_fa456_y3;
  wire f_s_dadda_rca24_fa456_y4;
  wire f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa456_y4;
  wire f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa351_y2;
  wire f_s_dadda_rca24_fa457_y0;
  wire f_s_dadda_rca24_fa457_y1;
  wire f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa352_y2;
  wire f_s_dadda_rca24_fa457_y2;
  wire f_s_dadda_rca24_fa457_y3;
  wire f_s_dadda_rca24_fa457_y4;
  wire f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa457_y4;
  wire f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa353_y2;
  wire f_s_dadda_rca24_fa458_y0;
  wire f_s_dadda_rca24_fa458_y1;
  wire f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa354_y2;
  wire f_s_dadda_rca24_fa458_y2;
  wire f_s_dadda_rca24_fa458_y3;
  wire f_s_dadda_rca24_fa458_y4;
  wire f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa458_y4;
  wire f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa355_y2;
  wire f_s_dadda_rca24_fa459_y0;
  wire f_s_dadda_rca24_fa459_y1;
  wire f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa356_y2;
  wire f_s_dadda_rca24_fa459_y2;
  wire f_s_dadda_rca24_fa459_y3;
  wire f_s_dadda_rca24_fa459_y4;
  wire f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa459_y4;
  wire f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa357_y2;
  wire f_s_dadda_rca24_fa460_y0;
  wire f_s_dadda_rca24_fa460_y1;
  wire f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa358_y2;
  wire f_s_dadda_rca24_fa460_y2;
  wire f_s_dadda_rca24_fa460_y3;
  wire f_s_dadda_rca24_fa460_y4;
  wire f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa460_y4;
  wire f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa359_y2;
  wire f_s_dadda_rca24_fa461_y0;
  wire f_s_dadda_rca24_fa461_y1;
  wire f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa360_y2;
  wire f_s_dadda_rca24_fa461_y2;
  wire f_s_dadda_rca24_fa461_y3;
  wire f_s_dadda_rca24_fa461_y4;
  wire f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa461_y4;
  wire f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa361_y2;
  wire f_s_dadda_rca24_fa462_y0;
  wire f_s_dadda_rca24_fa462_y1;
  wire f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa362_y2;
  wire f_s_dadda_rca24_fa462_y2;
  wire f_s_dadda_rca24_fa462_y3;
  wire f_s_dadda_rca24_fa462_y4;
  wire f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa462_y4;
  wire f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa363_y2;
  wire f_s_dadda_rca24_fa463_y0;
  wire f_s_dadda_rca24_fa463_y1;
  wire f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa364_y2;
  wire f_s_dadda_rca24_fa463_y2;
  wire f_s_dadda_rca24_fa463_y3;
  wire f_s_dadda_rca24_fa463_y4;
  wire f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa463_y4;
  wire f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa365_y2;
  wire f_s_dadda_rca24_fa464_y0;
  wire f_s_dadda_rca24_fa464_y1;
  wire f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa366_y2;
  wire f_s_dadda_rca24_fa464_y2;
  wire f_s_dadda_rca24_fa464_y3;
  wire f_s_dadda_rca24_fa464_y4;
  wire f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa464_y4;
  wire f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa367_y2;
  wire f_s_dadda_rca24_fa465_y0;
  wire f_s_dadda_rca24_fa465_y1;
  wire f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa368_y2;
  wire f_s_dadda_rca24_fa465_y2;
  wire f_s_dadda_rca24_fa465_y3;
  wire f_s_dadda_rca24_fa465_y4;
  wire f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa465_y4;
  wire f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa369_y2;
  wire f_s_dadda_rca24_fa466_y0;
  wire f_s_dadda_rca24_fa466_y1;
  wire f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa370_y2;
  wire f_s_dadda_rca24_fa466_y2;
  wire f_s_dadda_rca24_fa466_y3;
  wire f_s_dadda_rca24_fa466_y4;
  wire f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa466_y4;
  wire f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa371_y2;
  wire f_s_dadda_rca24_fa467_y0;
  wire f_s_dadda_rca24_fa467_y1;
  wire f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa372_y2;
  wire f_s_dadda_rca24_fa467_y2;
  wire f_s_dadda_rca24_fa467_y3;
  wire f_s_dadda_rca24_fa467_y4;
  wire f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa467_y4;
  wire f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa373_y2;
  wire f_s_dadda_rca24_fa468_y0;
  wire f_s_dadda_rca24_fa468_y1;
  wire f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa374_y2;
  wire f_s_dadda_rca24_fa468_y2;
  wire f_s_dadda_rca24_fa468_y3;
  wire f_s_dadda_rca24_fa468_y4;
  wire f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa468_y4;
  wire f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa375_y2;
  wire f_s_dadda_rca24_fa469_y0;
  wire f_s_dadda_rca24_fa469_y1;
  wire f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa376_y2;
  wire f_s_dadda_rca24_fa469_y2;
  wire f_s_dadda_rca24_fa469_y3;
  wire f_s_dadda_rca24_fa469_y4;
  wire f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa469_y4;
  wire f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa377_y2;
  wire f_s_dadda_rca24_fa470_y0;
  wire f_s_dadda_rca24_fa470_y1;
  wire f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa378_y2;
  wire f_s_dadda_rca24_fa470_y2;
  wire f_s_dadda_rca24_fa470_y3;
  wire f_s_dadda_rca24_fa470_y4;
  wire f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa470_y4;
  wire f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa379_y2;
  wire f_s_dadda_rca24_fa471_y0;
  wire f_s_dadda_rca24_fa471_y1;
  wire f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa380_y2;
  wire f_s_dadda_rca24_fa471_y2;
  wire f_s_dadda_rca24_fa471_y3;
  wire f_s_dadda_rca24_fa471_y4;
  wire f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa471_y4;
  wire f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa381_y2;
  wire f_s_dadda_rca24_fa472_y0;
  wire f_s_dadda_rca24_fa472_y1;
  wire f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa382_y2;
  wire f_s_dadda_rca24_fa472_y2;
  wire f_s_dadda_rca24_fa472_y3;
  wire f_s_dadda_rca24_fa472_y4;
  wire f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa472_y4;
  wire f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa383_y2;
  wire f_s_dadda_rca24_fa473_y0;
  wire f_s_dadda_rca24_fa473_y1;
  wire f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa384_y2;
  wire f_s_dadda_rca24_fa473_y2;
  wire f_s_dadda_rca24_fa473_y3;
  wire f_s_dadda_rca24_fa473_y4;
  wire f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa473_y4;
  wire f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa385_y2;
  wire f_s_dadda_rca24_fa474_y0;
  wire f_s_dadda_rca24_fa474_y1;
  wire f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa386_y2;
  wire f_s_dadda_rca24_fa474_y2;
  wire f_s_dadda_rca24_fa474_y3;
  wire f_s_dadda_rca24_fa474_y4;
  wire f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa474_y4;
  wire f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa387_y2;
  wire f_s_dadda_rca24_fa475_y0;
  wire f_s_dadda_rca24_fa475_y1;
  wire f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa388_y2;
  wire f_s_dadda_rca24_fa475_y2;
  wire f_s_dadda_rca24_fa475_y3;
  wire f_s_dadda_rca24_fa475_y4;
  wire f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa475_y4;
  wire f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa389_y2;
  wire f_s_dadda_rca24_fa476_y0;
  wire f_s_dadda_rca24_fa476_y1;
  wire f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa390_y2;
  wire f_s_dadda_rca24_fa476_y2;
  wire f_s_dadda_rca24_fa476_y3;
  wire f_s_dadda_rca24_fa476_y4;
  wire f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa476_y4;
  wire f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa391_y2;
  wire f_s_dadda_rca24_fa477_y0;
  wire f_s_dadda_rca24_fa477_y1;
  wire f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa392_y2;
  wire f_s_dadda_rca24_fa477_y2;
  wire f_s_dadda_rca24_fa477_y3;
  wire f_s_dadda_rca24_fa477_y4;
  wire f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa477_y4;
  wire f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa393_y2;
  wire f_s_dadda_rca24_fa478_y0;
  wire f_s_dadda_rca24_fa478_y1;
  wire f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa394_y2;
  wire f_s_dadda_rca24_fa478_y2;
  wire f_s_dadda_rca24_fa478_y3;
  wire f_s_dadda_rca24_fa478_y4;
  wire f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa478_y4;
  wire f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa395_y2;
  wire f_s_dadda_rca24_fa479_y0;
  wire f_s_dadda_rca24_fa479_y1;
  wire f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa396_y2;
  wire f_s_dadda_rca24_fa479_y2;
  wire f_s_dadda_rca24_fa479_y3;
  wire f_s_dadda_rca24_fa479_y4;
  wire f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa479_y4;
  wire f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa397_y2;
  wire f_s_dadda_rca24_fa480_y0;
  wire f_s_dadda_rca24_fa480_y1;
  wire f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa398_y2;
  wire f_s_dadda_rca24_fa480_y2;
  wire f_s_dadda_rca24_fa480_y3;
  wire f_s_dadda_rca24_fa480_y4;
  wire f_s_dadda_rca24_nand_20_23_a_20;
  wire f_s_dadda_rca24_nand_20_23_b_23;
  wire f_s_dadda_rca24_nand_20_23_y0;
  wire f_s_dadda_rca24_fa481_f_s_dadda_rca24_fa480_y4;
  wire f_s_dadda_rca24_fa481_f_s_dadda_rca24_nand_20_23_y0;
  wire f_s_dadda_rca24_fa481_y0;
  wire f_s_dadda_rca24_fa481_y1;
  wire f_s_dadda_rca24_fa481_f_s_dadda_rca24_fa399_y2;
  wire f_s_dadda_rca24_fa481_y2;
  wire f_s_dadda_rca24_fa481_y3;
  wire f_s_dadda_rca24_fa481_y4;
  wire f_s_dadda_rca24_and_22_22_a_22;
  wire f_s_dadda_rca24_and_22_22_b_22;
  wire f_s_dadda_rca24_and_22_22_y0;
  wire f_s_dadda_rca24_nand_21_23_a_21;
  wire f_s_dadda_rca24_nand_21_23_b_23;
  wire f_s_dadda_rca24_nand_21_23_y0;
  wire f_s_dadda_rca24_fa482_f_s_dadda_rca24_fa481_y4;
  wire f_s_dadda_rca24_fa482_f_s_dadda_rca24_and_22_22_y0;
  wire f_s_dadda_rca24_fa482_y0;
  wire f_s_dadda_rca24_fa482_y1;
  wire f_s_dadda_rca24_fa482_f_s_dadda_rca24_nand_21_23_y0;
  wire f_s_dadda_rca24_fa482_y2;
  wire f_s_dadda_rca24_fa482_y3;
  wire f_s_dadda_rca24_fa482_y4;
  wire f_s_dadda_rca24_nand_23_22_a_23;
  wire f_s_dadda_rca24_nand_23_22_b_22;
  wire f_s_dadda_rca24_nand_23_22_y0;
  wire f_s_dadda_rca24_fa483_f_s_dadda_rca24_fa482_y4;
  wire f_s_dadda_rca24_fa483_f_s_dadda_rca24_fa440_y4;
  wire f_s_dadda_rca24_fa483_y0;
  wire f_s_dadda_rca24_fa483_y1;
  wire f_s_dadda_rca24_fa483_f_s_dadda_rca24_nand_23_22_y0;
  wire f_s_dadda_rca24_fa483_y2;
  wire f_s_dadda_rca24_fa483_y3;
  wire f_s_dadda_rca24_fa483_y4;
  wire f_s_dadda_rca24_and_0_0_a_0;
  wire f_s_dadda_rca24_and_0_0_b_0;
  wire f_s_dadda_rca24_and_0_0_y0;
  wire f_s_dadda_rca24_and_1_0_a_1;
  wire f_s_dadda_rca24_and_1_0_b_0;
  wire f_s_dadda_rca24_and_1_0_y0;
  wire f_s_dadda_rca24_and_0_2_a_0;
  wire f_s_dadda_rca24_and_0_2_b_2;
  wire f_s_dadda_rca24_and_0_2_y0;
  wire f_s_dadda_rca24_nand_22_23_a_22;
  wire f_s_dadda_rca24_nand_22_23_b_23;
  wire f_s_dadda_rca24_nand_22_23_y0;
  wire f_s_dadda_rca24_and_0_1_a_0;
  wire f_s_dadda_rca24_and_0_1_b_1;
  wire f_s_dadda_rca24_and_0_1_y0;
  wire f_s_dadda_rca24_and_23_23_a_23;
  wire f_s_dadda_rca24_and_23_23_b_23;
  wire f_s_dadda_rca24_and_23_23_y0;
  wire f_s_dadda_rca24_u_rca_ha_f_s_dadda_rca24_and_1_0_y0;
  wire f_s_dadda_rca24_u_rca_ha_f_s_dadda_rca24_and_0_1_y0;
  wire f_s_dadda_rca24_u_rca_ha_y0;
  wire f_s_dadda_rca24_u_rca_ha_y1;
  wire f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_and_0_2_y0;
  wire f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_ha21_y0;
  wire f_s_dadda_rca24_u_rca_fa1_y0;
  wire f_s_dadda_rca24_u_rca_fa1_y1;
  wire f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_u_rca_ha_y1;
  wire f_s_dadda_rca24_u_rca_fa1_y2;
  wire f_s_dadda_rca24_u_rca_fa1_y3;
  wire f_s_dadda_rca24_u_rca_fa1_y4;
  wire f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_ha20_y0;
  wire f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_fa441_y2;
  wire f_s_dadda_rca24_u_rca_fa2_y0;
  wire f_s_dadda_rca24_u_rca_fa2_y1;
  wire f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_u_rca_fa1_y4;
  wire f_s_dadda_rca24_u_rca_fa2_y2;
  wire f_s_dadda_rca24_u_rca_fa2_y3;
  wire f_s_dadda_rca24_u_rca_fa2_y4;
  wire f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_fa400_y2;
  wire f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_fa442_y2;
  wire f_s_dadda_rca24_u_rca_fa3_y0;
  wire f_s_dadda_rca24_u_rca_fa3_y1;
  wire f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_u_rca_fa2_y4;
  wire f_s_dadda_rca24_u_rca_fa3_y2;
  wire f_s_dadda_rca24_u_rca_fa3_y3;
  wire f_s_dadda_rca24_u_rca_fa3_y4;
  wire f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_fa401_y2;
  wire f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_fa443_y2;
  wire f_s_dadda_rca24_u_rca_fa4_y0;
  wire f_s_dadda_rca24_u_rca_fa4_y1;
  wire f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_u_rca_fa3_y4;
  wire f_s_dadda_rca24_u_rca_fa4_y2;
  wire f_s_dadda_rca24_u_rca_fa4_y3;
  wire f_s_dadda_rca24_u_rca_fa4_y4;
  wire f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_fa402_y2;
  wire f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_fa444_y2;
  wire f_s_dadda_rca24_u_rca_fa5_y0;
  wire f_s_dadda_rca24_u_rca_fa5_y1;
  wire f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_u_rca_fa4_y4;
  wire f_s_dadda_rca24_u_rca_fa5_y2;
  wire f_s_dadda_rca24_u_rca_fa5_y3;
  wire f_s_dadda_rca24_u_rca_fa5_y4;
  wire f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_fa403_y2;
  wire f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_fa445_y2;
  wire f_s_dadda_rca24_u_rca_fa6_y0;
  wire f_s_dadda_rca24_u_rca_fa6_y1;
  wire f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_u_rca_fa5_y4;
  wire f_s_dadda_rca24_u_rca_fa6_y2;
  wire f_s_dadda_rca24_u_rca_fa6_y3;
  wire f_s_dadda_rca24_u_rca_fa6_y4;
  wire f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_fa404_y2;
  wire f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_fa446_y2;
  wire f_s_dadda_rca24_u_rca_fa7_y0;
  wire f_s_dadda_rca24_u_rca_fa7_y1;
  wire f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_u_rca_fa6_y4;
  wire f_s_dadda_rca24_u_rca_fa7_y2;
  wire f_s_dadda_rca24_u_rca_fa7_y3;
  wire f_s_dadda_rca24_u_rca_fa7_y4;
  wire f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_fa405_y2;
  wire f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_fa447_y2;
  wire f_s_dadda_rca24_u_rca_fa8_y0;
  wire f_s_dadda_rca24_u_rca_fa8_y1;
  wire f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_u_rca_fa7_y4;
  wire f_s_dadda_rca24_u_rca_fa8_y2;
  wire f_s_dadda_rca24_u_rca_fa8_y3;
  wire f_s_dadda_rca24_u_rca_fa8_y4;
  wire f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_fa406_y2;
  wire f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_fa448_y2;
  wire f_s_dadda_rca24_u_rca_fa9_y0;
  wire f_s_dadda_rca24_u_rca_fa9_y1;
  wire f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_u_rca_fa8_y4;
  wire f_s_dadda_rca24_u_rca_fa9_y2;
  wire f_s_dadda_rca24_u_rca_fa9_y3;
  wire f_s_dadda_rca24_u_rca_fa9_y4;
  wire f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_fa407_y2;
  wire f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_fa449_y2;
  wire f_s_dadda_rca24_u_rca_fa10_y0;
  wire f_s_dadda_rca24_u_rca_fa10_y1;
  wire f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_u_rca_fa9_y4;
  wire f_s_dadda_rca24_u_rca_fa10_y2;
  wire f_s_dadda_rca24_u_rca_fa10_y3;
  wire f_s_dadda_rca24_u_rca_fa10_y4;
  wire f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_fa408_y2;
  wire f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_fa450_y2;
  wire f_s_dadda_rca24_u_rca_fa11_y0;
  wire f_s_dadda_rca24_u_rca_fa11_y1;
  wire f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_u_rca_fa10_y4;
  wire f_s_dadda_rca24_u_rca_fa11_y2;
  wire f_s_dadda_rca24_u_rca_fa11_y3;
  wire f_s_dadda_rca24_u_rca_fa11_y4;
  wire f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_fa409_y2;
  wire f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_fa451_y2;
  wire f_s_dadda_rca24_u_rca_fa12_y0;
  wire f_s_dadda_rca24_u_rca_fa12_y1;
  wire f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_u_rca_fa11_y4;
  wire f_s_dadda_rca24_u_rca_fa12_y2;
  wire f_s_dadda_rca24_u_rca_fa12_y3;
  wire f_s_dadda_rca24_u_rca_fa12_y4;
  wire f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_fa410_y2;
  wire f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_fa452_y2;
  wire f_s_dadda_rca24_u_rca_fa13_y0;
  wire f_s_dadda_rca24_u_rca_fa13_y1;
  wire f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_u_rca_fa12_y4;
  wire f_s_dadda_rca24_u_rca_fa13_y2;
  wire f_s_dadda_rca24_u_rca_fa13_y3;
  wire f_s_dadda_rca24_u_rca_fa13_y4;
  wire f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_fa411_y2;
  wire f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_fa453_y2;
  wire f_s_dadda_rca24_u_rca_fa14_y0;
  wire f_s_dadda_rca24_u_rca_fa14_y1;
  wire f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_u_rca_fa13_y4;
  wire f_s_dadda_rca24_u_rca_fa14_y2;
  wire f_s_dadda_rca24_u_rca_fa14_y3;
  wire f_s_dadda_rca24_u_rca_fa14_y4;
  wire f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_fa412_y2;
  wire f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_fa454_y2;
  wire f_s_dadda_rca24_u_rca_fa15_y0;
  wire f_s_dadda_rca24_u_rca_fa15_y1;
  wire f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_u_rca_fa14_y4;
  wire f_s_dadda_rca24_u_rca_fa15_y2;
  wire f_s_dadda_rca24_u_rca_fa15_y3;
  wire f_s_dadda_rca24_u_rca_fa15_y4;
  wire f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_fa413_y2;
  wire f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_fa455_y2;
  wire f_s_dadda_rca24_u_rca_fa16_y0;
  wire f_s_dadda_rca24_u_rca_fa16_y1;
  wire f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_u_rca_fa15_y4;
  wire f_s_dadda_rca24_u_rca_fa16_y2;
  wire f_s_dadda_rca24_u_rca_fa16_y3;
  wire f_s_dadda_rca24_u_rca_fa16_y4;
  wire f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_fa414_y2;
  wire f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_fa456_y2;
  wire f_s_dadda_rca24_u_rca_fa17_y0;
  wire f_s_dadda_rca24_u_rca_fa17_y1;
  wire f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_u_rca_fa16_y4;
  wire f_s_dadda_rca24_u_rca_fa17_y2;
  wire f_s_dadda_rca24_u_rca_fa17_y3;
  wire f_s_dadda_rca24_u_rca_fa17_y4;
  wire f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_fa415_y2;
  wire f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_fa457_y2;
  wire f_s_dadda_rca24_u_rca_fa18_y0;
  wire f_s_dadda_rca24_u_rca_fa18_y1;
  wire f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_u_rca_fa17_y4;
  wire f_s_dadda_rca24_u_rca_fa18_y2;
  wire f_s_dadda_rca24_u_rca_fa18_y3;
  wire f_s_dadda_rca24_u_rca_fa18_y4;
  wire f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_fa416_y2;
  wire f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_fa458_y2;
  wire f_s_dadda_rca24_u_rca_fa19_y0;
  wire f_s_dadda_rca24_u_rca_fa19_y1;
  wire f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_u_rca_fa18_y4;
  wire f_s_dadda_rca24_u_rca_fa19_y2;
  wire f_s_dadda_rca24_u_rca_fa19_y3;
  wire f_s_dadda_rca24_u_rca_fa19_y4;
  wire f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_fa417_y2;
  wire f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_fa459_y2;
  wire f_s_dadda_rca24_u_rca_fa20_y0;
  wire f_s_dadda_rca24_u_rca_fa20_y1;
  wire f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_u_rca_fa19_y4;
  wire f_s_dadda_rca24_u_rca_fa20_y2;
  wire f_s_dadda_rca24_u_rca_fa20_y3;
  wire f_s_dadda_rca24_u_rca_fa20_y4;
  wire f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_fa418_y2;
  wire f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_fa460_y2;
  wire f_s_dadda_rca24_u_rca_fa21_y0;
  wire f_s_dadda_rca24_u_rca_fa21_y1;
  wire f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_u_rca_fa20_y4;
  wire f_s_dadda_rca24_u_rca_fa21_y2;
  wire f_s_dadda_rca24_u_rca_fa21_y3;
  wire f_s_dadda_rca24_u_rca_fa21_y4;
  wire f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_fa419_y2;
  wire f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_fa461_y2;
  wire f_s_dadda_rca24_u_rca_fa22_y0;
  wire f_s_dadda_rca24_u_rca_fa22_y1;
  wire f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_u_rca_fa21_y4;
  wire f_s_dadda_rca24_u_rca_fa22_y2;
  wire f_s_dadda_rca24_u_rca_fa22_y3;
  wire f_s_dadda_rca24_u_rca_fa22_y4;
  wire f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_fa420_y2;
  wire f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_fa462_y2;
  wire f_s_dadda_rca24_u_rca_fa23_y0;
  wire f_s_dadda_rca24_u_rca_fa23_y1;
  wire f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_u_rca_fa22_y4;
  wire f_s_dadda_rca24_u_rca_fa23_y2;
  wire f_s_dadda_rca24_u_rca_fa23_y3;
  wire f_s_dadda_rca24_u_rca_fa23_y4;
  wire f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_fa421_y2;
  wire f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_fa463_y2;
  wire f_s_dadda_rca24_u_rca_fa24_y0;
  wire f_s_dadda_rca24_u_rca_fa24_y1;
  wire f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_u_rca_fa23_y4;
  wire f_s_dadda_rca24_u_rca_fa24_y2;
  wire f_s_dadda_rca24_u_rca_fa24_y3;
  wire f_s_dadda_rca24_u_rca_fa24_y4;
  wire f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_fa422_y2;
  wire f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_fa464_y2;
  wire f_s_dadda_rca24_u_rca_fa25_y0;
  wire f_s_dadda_rca24_u_rca_fa25_y1;
  wire f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_u_rca_fa24_y4;
  wire f_s_dadda_rca24_u_rca_fa25_y2;
  wire f_s_dadda_rca24_u_rca_fa25_y3;
  wire f_s_dadda_rca24_u_rca_fa25_y4;
  wire f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_fa423_y2;
  wire f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_fa465_y2;
  wire f_s_dadda_rca24_u_rca_fa26_y0;
  wire f_s_dadda_rca24_u_rca_fa26_y1;
  wire f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_u_rca_fa25_y4;
  wire f_s_dadda_rca24_u_rca_fa26_y2;
  wire f_s_dadda_rca24_u_rca_fa26_y3;
  wire f_s_dadda_rca24_u_rca_fa26_y4;
  wire f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_fa424_y2;
  wire f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_fa466_y2;
  wire f_s_dadda_rca24_u_rca_fa27_y0;
  wire f_s_dadda_rca24_u_rca_fa27_y1;
  wire f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_u_rca_fa26_y4;
  wire f_s_dadda_rca24_u_rca_fa27_y2;
  wire f_s_dadda_rca24_u_rca_fa27_y3;
  wire f_s_dadda_rca24_u_rca_fa27_y4;
  wire f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_fa425_y2;
  wire f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_fa467_y2;
  wire f_s_dadda_rca24_u_rca_fa28_y0;
  wire f_s_dadda_rca24_u_rca_fa28_y1;
  wire f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_u_rca_fa27_y4;
  wire f_s_dadda_rca24_u_rca_fa28_y2;
  wire f_s_dadda_rca24_u_rca_fa28_y3;
  wire f_s_dadda_rca24_u_rca_fa28_y4;
  wire f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_fa426_y2;
  wire f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_fa468_y2;
  wire f_s_dadda_rca24_u_rca_fa29_y0;
  wire f_s_dadda_rca24_u_rca_fa29_y1;
  wire f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_u_rca_fa28_y4;
  wire f_s_dadda_rca24_u_rca_fa29_y2;
  wire f_s_dadda_rca24_u_rca_fa29_y3;
  wire f_s_dadda_rca24_u_rca_fa29_y4;
  wire f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_fa427_y2;
  wire f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_fa469_y2;
  wire f_s_dadda_rca24_u_rca_fa30_y0;
  wire f_s_dadda_rca24_u_rca_fa30_y1;
  wire f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_u_rca_fa29_y4;
  wire f_s_dadda_rca24_u_rca_fa30_y2;
  wire f_s_dadda_rca24_u_rca_fa30_y3;
  wire f_s_dadda_rca24_u_rca_fa30_y4;
  wire f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_fa428_y2;
  wire f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_fa470_y2;
  wire f_s_dadda_rca24_u_rca_fa31_y0;
  wire f_s_dadda_rca24_u_rca_fa31_y1;
  wire f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_u_rca_fa30_y4;
  wire f_s_dadda_rca24_u_rca_fa31_y2;
  wire f_s_dadda_rca24_u_rca_fa31_y3;
  wire f_s_dadda_rca24_u_rca_fa31_y4;
  wire f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_fa429_y2;
  wire f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_fa471_y2;
  wire f_s_dadda_rca24_u_rca_fa32_y0;
  wire f_s_dadda_rca24_u_rca_fa32_y1;
  wire f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_u_rca_fa31_y4;
  wire f_s_dadda_rca24_u_rca_fa32_y2;
  wire f_s_dadda_rca24_u_rca_fa32_y3;
  wire f_s_dadda_rca24_u_rca_fa32_y4;
  wire f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_fa430_y2;
  wire f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_fa472_y2;
  wire f_s_dadda_rca24_u_rca_fa33_y0;
  wire f_s_dadda_rca24_u_rca_fa33_y1;
  wire f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_u_rca_fa32_y4;
  wire f_s_dadda_rca24_u_rca_fa33_y2;
  wire f_s_dadda_rca24_u_rca_fa33_y3;
  wire f_s_dadda_rca24_u_rca_fa33_y4;
  wire f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_fa431_y2;
  wire f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_fa473_y2;
  wire f_s_dadda_rca24_u_rca_fa34_y0;
  wire f_s_dadda_rca24_u_rca_fa34_y1;
  wire f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_u_rca_fa33_y4;
  wire f_s_dadda_rca24_u_rca_fa34_y2;
  wire f_s_dadda_rca24_u_rca_fa34_y3;
  wire f_s_dadda_rca24_u_rca_fa34_y4;
  wire f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_fa432_y2;
  wire f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_fa474_y2;
  wire f_s_dadda_rca24_u_rca_fa35_y0;
  wire f_s_dadda_rca24_u_rca_fa35_y1;
  wire f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_u_rca_fa34_y4;
  wire f_s_dadda_rca24_u_rca_fa35_y2;
  wire f_s_dadda_rca24_u_rca_fa35_y3;
  wire f_s_dadda_rca24_u_rca_fa35_y4;
  wire f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_fa433_y2;
  wire f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_fa475_y2;
  wire f_s_dadda_rca24_u_rca_fa36_y0;
  wire f_s_dadda_rca24_u_rca_fa36_y1;
  wire f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_u_rca_fa35_y4;
  wire f_s_dadda_rca24_u_rca_fa36_y2;
  wire f_s_dadda_rca24_u_rca_fa36_y3;
  wire f_s_dadda_rca24_u_rca_fa36_y4;
  wire f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_fa434_y2;
  wire f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_fa476_y2;
  wire f_s_dadda_rca24_u_rca_fa37_y0;
  wire f_s_dadda_rca24_u_rca_fa37_y1;
  wire f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_u_rca_fa36_y4;
  wire f_s_dadda_rca24_u_rca_fa37_y2;
  wire f_s_dadda_rca24_u_rca_fa37_y3;
  wire f_s_dadda_rca24_u_rca_fa37_y4;
  wire f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_fa435_y2;
  wire f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_fa477_y2;
  wire f_s_dadda_rca24_u_rca_fa38_y0;
  wire f_s_dadda_rca24_u_rca_fa38_y1;
  wire f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_u_rca_fa37_y4;
  wire f_s_dadda_rca24_u_rca_fa38_y2;
  wire f_s_dadda_rca24_u_rca_fa38_y3;
  wire f_s_dadda_rca24_u_rca_fa38_y4;
  wire f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_fa436_y2;
  wire f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_fa478_y2;
  wire f_s_dadda_rca24_u_rca_fa39_y0;
  wire f_s_dadda_rca24_u_rca_fa39_y1;
  wire f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_u_rca_fa38_y4;
  wire f_s_dadda_rca24_u_rca_fa39_y2;
  wire f_s_dadda_rca24_u_rca_fa39_y3;
  wire f_s_dadda_rca24_u_rca_fa39_y4;
  wire f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_fa437_y2;
  wire f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_fa479_y2;
  wire f_s_dadda_rca24_u_rca_fa40_y0;
  wire f_s_dadda_rca24_u_rca_fa40_y1;
  wire f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_u_rca_fa39_y4;
  wire f_s_dadda_rca24_u_rca_fa40_y2;
  wire f_s_dadda_rca24_u_rca_fa40_y3;
  wire f_s_dadda_rca24_u_rca_fa40_y4;
  wire f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_fa438_y2;
  wire f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_fa480_y2;
  wire f_s_dadda_rca24_u_rca_fa41_y0;
  wire f_s_dadda_rca24_u_rca_fa41_y1;
  wire f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_u_rca_fa40_y4;
  wire f_s_dadda_rca24_u_rca_fa41_y2;
  wire f_s_dadda_rca24_u_rca_fa41_y3;
  wire f_s_dadda_rca24_u_rca_fa41_y4;
  wire f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_fa439_y2;
  wire f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_fa481_y2;
  wire f_s_dadda_rca24_u_rca_fa42_y0;
  wire f_s_dadda_rca24_u_rca_fa42_y1;
  wire f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_u_rca_fa41_y4;
  wire f_s_dadda_rca24_u_rca_fa42_y2;
  wire f_s_dadda_rca24_u_rca_fa42_y3;
  wire f_s_dadda_rca24_u_rca_fa42_y4;
  wire f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_fa440_y2;
  wire f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_fa482_y2;
  wire f_s_dadda_rca24_u_rca_fa43_y0;
  wire f_s_dadda_rca24_u_rca_fa43_y1;
  wire f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_u_rca_fa42_y4;
  wire f_s_dadda_rca24_u_rca_fa43_y2;
  wire f_s_dadda_rca24_u_rca_fa43_y3;
  wire f_s_dadda_rca24_u_rca_fa43_y4;
  wire f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_nand_22_23_y0;
  wire f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_fa483_y2;
  wire f_s_dadda_rca24_u_rca_fa44_y0;
  wire f_s_dadda_rca24_u_rca_fa44_y1;
  wire f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_u_rca_fa43_y4;
  wire f_s_dadda_rca24_u_rca_fa44_y2;
  wire f_s_dadda_rca24_u_rca_fa44_y3;
  wire f_s_dadda_rca24_u_rca_fa44_y4;
  wire f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_fa483_y4;
  wire f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_and_23_23_y0;
  wire f_s_dadda_rca24_u_rca_fa45_y0;
  wire f_s_dadda_rca24_u_rca_fa45_y1;
  wire f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_u_rca_fa44_y4;
  wire f_s_dadda_rca24_u_rca_fa45_y2;
  wire f_s_dadda_rca24_u_rca_fa45_y3;
  wire f_s_dadda_rca24_u_rca_fa45_y4;
  wire f_s_dadda_rca24_xor0_constant_wire_1;
  wire f_s_dadda_rca24_xor0_f_s_dadda_rca24_u_rca_fa45_y4;
  wire f_s_dadda_rca24_xor0_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign a_16 = a[16];
  assign a_17 = a[17];
  assign a_18 = a[18];
  assign a_19 = a[19];
  assign a_20 = a[20];
  assign a_21 = a[21];
  assign a_22 = a[22];
  assign a_23 = a[23];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign b_16 = b[16];
  assign b_17 = b[17];
  assign b_18 = b[18];
  assign b_19 = b[19];
  assign b_20 = b[20];
  assign b_21 = b[21];
  assign b_22 = b[22];
  assign b_23 = b[23];
  assign constant_wire_value_1_a_0 = a_0;
  assign constant_wire_value_1_b_0 = b_0;
  assign constant_wire_value_1_y0 = constant_wire_value_1_a_0 ^ constant_wire_value_1_b_0;
  assign constant_wire_value_1_y1 = ~(constant_wire_value_1_a_0 ^ constant_wire_value_1_b_0);
  assign constant_wire_1 = constant_wire_value_1_y0 | constant_wire_value_1_y1;
  assign f_s_dadda_rca24_and_19_0_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_19_0_y0 = f_s_dadda_rca24_and_19_0_a_19 & f_s_dadda_rca24_and_19_0_b_0;
  assign f_s_dadda_rca24_and_18_1_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_18_1_y0 = f_s_dadda_rca24_and_18_1_a_18 & f_s_dadda_rca24_and_18_1_b_1;
  assign f_s_dadda_rca24_ha0_f_s_dadda_rca24_and_19_0_y0 = f_s_dadda_rca24_and_19_0_y0;
  assign f_s_dadda_rca24_ha0_f_s_dadda_rca24_and_18_1_y0 = f_s_dadda_rca24_and_18_1_y0;
  assign f_s_dadda_rca24_ha0_y0 = f_s_dadda_rca24_ha0_f_s_dadda_rca24_and_19_0_y0 ^ f_s_dadda_rca24_ha0_f_s_dadda_rca24_and_18_1_y0;
  assign f_s_dadda_rca24_ha0_y1 = f_s_dadda_rca24_ha0_f_s_dadda_rca24_and_19_0_y0 & f_s_dadda_rca24_ha0_f_s_dadda_rca24_and_18_1_y0;
  assign f_s_dadda_rca24_and_20_0_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_20_0_y0 = f_s_dadda_rca24_and_20_0_a_20 & f_s_dadda_rca24_and_20_0_b_0;
  assign f_s_dadda_rca24_and_19_1_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_19_1_y0 = f_s_dadda_rca24_and_19_1_a_19 & f_s_dadda_rca24_and_19_1_b_1;
  assign f_s_dadda_rca24_fa0_f_s_dadda_rca24_ha0_y1 = f_s_dadda_rca24_ha0_y1;
  assign f_s_dadda_rca24_fa0_f_s_dadda_rca24_and_20_0_y0 = f_s_dadda_rca24_and_20_0_y0;
  assign f_s_dadda_rca24_fa0_f_s_dadda_rca24_and_19_1_y0 = f_s_dadda_rca24_and_19_1_y0;
  assign f_s_dadda_rca24_fa0_y0 = f_s_dadda_rca24_fa0_f_s_dadda_rca24_ha0_y1 ^ f_s_dadda_rca24_fa0_f_s_dadda_rca24_and_20_0_y0;
  assign f_s_dadda_rca24_fa0_y1 = f_s_dadda_rca24_fa0_f_s_dadda_rca24_ha0_y1 & f_s_dadda_rca24_fa0_f_s_dadda_rca24_and_20_0_y0;
  assign f_s_dadda_rca24_fa0_y2 = f_s_dadda_rca24_fa0_y0 ^ f_s_dadda_rca24_fa0_f_s_dadda_rca24_and_19_1_y0;
  assign f_s_dadda_rca24_fa0_y3 = f_s_dadda_rca24_fa0_y0 & f_s_dadda_rca24_fa0_f_s_dadda_rca24_and_19_1_y0;
  assign f_s_dadda_rca24_fa0_y4 = f_s_dadda_rca24_fa0_y1 | f_s_dadda_rca24_fa0_y3;
  assign f_s_dadda_rca24_and_18_2_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_18_2_y0 = f_s_dadda_rca24_and_18_2_a_18 & f_s_dadda_rca24_and_18_2_b_2;
  assign f_s_dadda_rca24_and_17_3_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_17_3_y0 = f_s_dadda_rca24_and_17_3_a_17 & f_s_dadda_rca24_and_17_3_b_3;
  assign f_s_dadda_rca24_ha1_f_s_dadda_rca24_and_18_2_y0 = f_s_dadda_rca24_and_18_2_y0;
  assign f_s_dadda_rca24_ha1_f_s_dadda_rca24_and_17_3_y0 = f_s_dadda_rca24_and_17_3_y0;
  assign f_s_dadda_rca24_ha1_y0 = f_s_dadda_rca24_ha1_f_s_dadda_rca24_and_18_2_y0 ^ f_s_dadda_rca24_ha1_f_s_dadda_rca24_and_17_3_y0;
  assign f_s_dadda_rca24_ha1_y1 = f_s_dadda_rca24_ha1_f_s_dadda_rca24_and_18_2_y0 & f_s_dadda_rca24_ha1_f_s_dadda_rca24_and_17_3_y0;
  assign f_s_dadda_rca24_and_21_0_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_21_0_y0 = f_s_dadda_rca24_and_21_0_a_21 & f_s_dadda_rca24_and_21_0_b_0;
  assign f_s_dadda_rca24_fa1_f_s_dadda_rca24_ha1_y1 = f_s_dadda_rca24_ha1_y1;
  assign f_s_dadda_rca24_fa1_f_s_dadda_rca24_fa0_y4 = f_s_dadda_rca24_fa0_y4;
  assign f_s_dadda_rca24_fa1_f_s_dadda_rca24_and_21_0_y0 = f_s_dadda_rca24_and_21_0_y0;
  assign f_s_dadda_rca24_fa1_y0 = f_s_dadda_rca24_fa1_f_s_dadda_rca24_ha1_y1 ^ f_s_dadda_rca24_fa1_f_s_dadda_rca24_fa0_y4;
  assign f_s_dadda_rca24_fa1_y1 = f_s_dadda_rca24_fa1_f_s_dadda_rca24_ha1_y1 & f_s_dadda_rca24_fa1_f_s_dadda_rca24_fa0_y4;
  assign f_s_dadda_rca24_fa1_y2 = f_s_dadda_rca24_fa1_y0 ^ f_s_dadda_rca24_fa1_f_s_dadda_rca24_and_21_0_y0;
  assign f_s_dadda_rca24_fa1_y3 = f_s_dadda_rca24_fa1_y0 & f_s_dadda_rca24_fa1_f_s_dadda_rca24_and_21_0_y0;
  assign f_s_dadda_rca24_fa1_y4 = f_s_dadda_rca24_fa1_y1 | f_s_dadda_rca24_fa1_y3;
  assign f_s_dadda_rca24_and_20_1_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_20_1_y0 = f_s_dadda_rca24_and_20_1_a_20 & f_s_dadda_rca24_and_20_1_b_1;
  assign f_s_dadda_rca24_and_19_2_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_19_2_y0 = f_s_dadda_rca24_and_19_2_a_19 & f_s_dadda_rca24_and_19_2_b_2;
  assign f_s_dadda_rca24_and_18_3_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_18_3_y0 = f_s_dadda_rca24_and_18_3_a_18 & f_s_dadda_rca24_and_18_3_b_3;
  assign f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_20_1_y0 = f_s_dadda_rca24_and_20_1_y0;
  assign f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_19_2_y0 = f_s_dadda_rca24_and_19_2_y0;
  assign f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_18_3_y0 = f_s_dadda_rca24_and_18_3_y0;
  assign f_s_dadda_rca24_fa2_y0 = f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_20_1_y0 ^ f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_19_2_y0;
  assign f_s_dadda_rca24_fa2_y1 = f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_20_1_y0 & f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_19_2_y0;
  assign f_s_dadda_rca24_fa2_y2 = f_s_dadda_rca24_fa2_y0 ^ f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_18_3_y0;
  assign f_s_dadda_rca24_fa2_y3 = f_s_dadda_rca24_fa2_y0 & f_s_dadda_rca24_fa2_f_s_dadda_rca24_and_18_3_y0;
  assign f_s_dadda_rca24_fa2_y4 = f_s_dadda_rca24_fa2_y1 | f_s_dadda_rca24_fa2_y3;
  assign f_s_dadda_rca24_and_17_4_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_17_4_y0 = f_s_dadda_rca24_and_17_4_a_17 & f_s_dadda_rca24_and_17_4_b_4;
  assign f_s_dadda_rca24_and_16_5_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_16_5_y0 = f_s_dadda_rca24_and_16_5_a_16 & f_s_dadda_rca24_and_16_5_b_5;
  assign f_s_dadda_rca24_ha2_f_s_dadda_rca24_and_17_4_y0 = f_s_dadda_rca24_and_17_4_y0;
  assign f_s_dadda_rca24_ha2_f_s_dadda_rca24_and_16_5_y0 = f_s_dadda_rca24_and_16_5_y0;
  assign f_s_dadda_rca24_ha2_y0 = f_s_dadda_rca24_ha2_f_s_dadda_rca24_and_17_4_y0 ^ f_s_dadda_rca24_ha2_f_s_dadda_rca24_and_16_5_y0;
  assign f_s_dadda_rca24_ha2_y1 = f_s_dadda_rca24_ha2_f_s_dadda_rca24_and_17_4_y0 & f_s_dadda_rca24_ha2_f_s_dadda_rca24_and_16_5_y0;
  assign f_s_dadda_rca24_fa3_f_s_dadda_rca24_ha2_y1 = f_s_dadda_rca24_ha2_y1;
  assign f_s_dadda_rca24_fa3_f_s_dadda_rca24_fa2_y4 = f_s_dadda_rca24_fa2_y4;
  assign f_s_dadda_rca24_fa3_f_s_dadda_rca24_fa1_y4 = f_s_dadda_rca24_fa1_y4;
  assign f_s_dadda_rca24_fa3_y0 = f_s_dadda_rca24_fa3_f_s_dadda_rca24_ha2_y1 ^ f_s_dadda_rca24_fa3_f_s_dadda_rca24_fa2_y4;
  assign f_s_dadda_rca24_fa3_y1 = f_s_dadda_rca24_fa3_f_s_dadda_rca24_ha2_y1 & f_s_dadda_rca24_fa3_f_s_dadda_rca24_fa2_y4;
  assign f_s_dadda_rca24_fa3_y2 = f_s_dadda_rca24_fa3_y0 ^ f_s_dadda_rca24_fa3_f_s_dadda_rca24_fa1_y4;
  assign f_s_dadda_rca24_fa3_y3 = f_s_dadda_rca24_fa3_y0 & f_s_dadda_rca24_fa3_f_s_dadda_rca24_fa1_y4;
  assign f_s_dadda_rca24_fa3_y4 = f_s_dadda_rca24_fa3_y1 | f_s_dadda_rca24_fa3_y3;
  assign f_s_dadda_rca24_and_22_0_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_22_0_y0 = f_s_dadda_rca24_and_22_0_a_22 & f_s_dadda_rca24_and_22_0_b_0;
  assign f_s_dadda_rca24_and_21_1_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_21_1_y0 = f_s_dadda_rca24_and_21_1_a_21 & f_s_dadda_rca24_and_21_1_b_1;
  assign f_s_dadda_rca24_and_20_2_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_20_2_y0 = f_s_dadda_rca24_and_20_2_a_20 & f_s_dadda_rca24_and_20_2_b_2;
  assign f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_22_0_y0 = f_s_dadda_rca24_and_22_0_y0;
  assign f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_21_1_y0 = f_s_dadda_rca24_and_21_1_y0;
  assign f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_20_2_y0 = f_s_dadda_rca24_and_20_2_y0;
  assign f_s_dadda_rca24_fa4_y0 = f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_22_0_y0 ^ f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_21_1_y0;
  assign f_s_dadda_rca24_fa4_y1 = f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_22_0_y0 & f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_21_1_y0;
  assign f_s_dadda_rca24_fa4_y2 = f_s_dadda_rca24_fa4_y0 ^ f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_20_2_y0;
  assign f_s_dadda_rca24_fa4_y3 = f_s_dadda_rca24_fa4_y0 & f_s_dadda_rca24_fa4_f_s_dadda_rca24_and_20_2_y0;
  assign f_s_dadda_rca24_fa4_y4 = f_s_dadda_rca24_fa4_y1 | f_s_dadda_rca24_fa4_y3;
  assign f_s_dadda_rca24_and_19_3_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_19_3_y0 = f_s_dadda_rca24_and_19_3_a_19 & f_s_dadda_rca24_and_19_3_b_3;
  assign f_s_dadda_rca24_and_18_4_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_18_4_y0 = f_s_dadda_rca24_and_18_4_a_18 & f_s_dadda_rca24_and_18_4_b_4;
  assign f_s_dadda_rca24_and_17_5_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_17_5_y0 = f_s_dadda_rca24_and_17_5_a_17 & f_s_dadda_rca24_and_17_5_b_5;
  assign f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_19_3_y0 = f_s_dadda_rca24_and_19_3_y0;
  assign f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_18_4_y0 = f_s_dadda_rca24_and_18_4_y0;
  assign f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_17_5_y0 = f_s_dadda_rca24_and_17_5_y0;
  assign f_s_dadda_rca24_fa5_y0 = f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_19_3_y0 ^ f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_18_4_y0;
  assign f_s_dadda_rca24_fa5_y1 = f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_19_3_y0 & f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_18_4_y0;
  assign f_s_dadda_rca24_fa5_y2 = f_s_dadda_rca24_fa5_y0 ^ f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_17_5_y0;
  assign f_s_dadda_rca24_fa5_y3 = f_s_dadda_rca24_fa5_y0 & f_s_dadda_rca24_fa5_f_s_dadda_rca24_and_17_5_y0;
  assign f_s_dadda_rca24_fa5_y4 = f_s_dadda_rca24_fa5_y1 | f_s_dadda_rca24_fa5_y3;
  assign f_s_dadda_rca24_and_16_6_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_16_6_y0 = f_s_dadda_rca24_and_16_6_a_16 & f_s_dadda_rca24_and_16_6_b_6;
  assign f_s_dadda_rca24_and_15_7_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_15_7_y0 = f_s_dadda_rca24_and_15_7_a_15 & f_s_dadda_rca24_and_15_7_b_7;
  assign f_s_dadda_rca24_ha3_f_s_dadda_rca24_and_16_6_y0 = f_s_dadda_rca24_and_16_6_y0;
  assign f_s_dadda_rca24_ha3_f_s_dadda_rca24_and_15_7_y0 = f_s_dadda_rca24_and_15_7_y0;
  assign f_s_dadda_rca24_ha3_y0 = f_s_dadda_rca24_ha3_f_s_dadda_rca24_and_16_6_y0 ^ f_s_dadda_rca24_ha3_f_s_dadda_rca24_and_15_7_y0;
  assign f_s_dadda_rca24_ha3_y1 = f_s_dadda_rca24_ha3_f_s_dadda_rca24_and_16_6_y0 & f_s_dadda_rca24_ha3_f_s_dadda_rca24_and_15_7_y0;
  assign f_s_dadda_rca24_fa6_f_s_dadda_rca24_ha3_y1 = f_s_dadda_rca24_ha3_y1;
  assign f_s_dadda_rca24_fa6_f_s_dadda_rca24_fa5_y4 = f_s_dadda_rca24_fa5_y4;
  assign f_s_dadda_rca24_fa6_f_s_dadda_rca24_fa4_y4 = f_s_dadda_rca24_fa4_y4;
  assign f_s_dadda_rca24_fa6_y0 = f_s_dadda_rca24_fa6_f_s_dadda_rca24_ha3_y1 ^ f_s_dadda_rca24_fa6_f_s_dadda_rca24_fa5_y4;
  assign f_s_dadda_rca24_fa6_y1 = f_s_dadda_rca24_fa6_f_s_dadda_rca24_ha3_y1 & f_s_dadda_rca24_fa6_f_s_dadda_rca24_fa5_y4;
  assign f_s_dadda_rca24_fa6_y2 = f_s_dadda_rca24_fa6_y0 ^ f_s_dadda_rca24_fa6_f_s_dadda_rca24_fa4_y4;
  assign f_s_dadda_rca24_fa6_y3 = f_s_dadda_rca24_fa6_y0 & f_s_dadda_rca24_fa6_f_s_dadda_rca24_fa4_y4;
  assign f_s_dadda_rca24_fa6_y4 = f_s_dadda_rca24_fa6_y1 | f_s_dadda_rca24_fa6_y3;
  assign f_s_dadda_rca24_nand_23_0_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_0_b_0 = b_0;
  assign f_s_dadda_rca24_nand_23_0_y0 = ~(f_s_dadda_rca24_nand_23_0_a_23 & f_s_dadda_rca24_nand_23_0_b_0);
  assign f_s_dadda_rca24_and_22_1_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_22_1_y0 = f_s_dadda_rca24_and_22_1_a_22 & f_s_dadda_rca24_and_22_1_b_1;
  assign f_s_dadda_rca24_fa7_f_s_dadda_rca24_fa3_y4 = f_s_dadda_rca24_fa3_y4;
  assign f_s_dadda_rca24_fa7_f_s_dadda_rca24_nand_23_0_y0 = f_s_dadda_rca24_nand_23_0_y0;
  assign f_s_dadda_rca24_fa7_f_s_dadda_rca24_and_22_1_y0 = f_s_dadda_rca24_and_22_1_y0;
  assign f_s_dadda_rca24_fa7_y0 = f_s_dadda_rca24_fa7_f_s_dadda_rca24_fa3_y4 ^ f_s_dadda_rca24_fa7_f_s_dadda_rca24_nand_23_0_y0;
  assign f_s_dadda_rca24_fa7_y1 = f_s_dadda_rca24_fa7_f_s_dadda_rca24_fa3_y4 & f_s_dadda_rca24_fa7_f_s_dadda_rca24_nand_23_0_y0;
  assign f_s_dadda_rca24_fa7_y2 = f_s_dadda_rca24_fa7_y0 ^ f_s_dadda_rca24_fa7_f_s_dadda_rca24_and_22_1_y0;
  assign f_s_dadda_rca24_fa7_y3 = f_s_dadda_rca24_fa7_y0 & f_s_dadda_rca24_fa7_f_s_dadda_rca24_and_22_1_y0;
  assign f_s_dadda_rca24_fa7_y4 = f_s_dadda_rca24_fa7_y1 | f_s_dadda_rca24_fa7_y3;
  assign f_s_dadda_rca24_and_21_2_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_21_2_y0 = f_s_dadda_rca24_and_21_2_a_21 & f_s_dadda_rca24_and_21_2_b_2;
  assign f_s_dadda_rca24_and_20_3_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_20_3_y0 = f_s_dadda_rca24_and_20_3_a_20 & f_s_dadda_rca24_and_20_3_b_3;
  assign f_s_dadda_rca24_and_19_4_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_19_4_y0 = f_s_dadda_rca24_and_19_4_a_19 & f_s_dadda_rca24_and_19_4_b_4;
  assign f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_21_2_y0 = f_s_dadda_rca24_and_21_2_y0;
  assign f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_20_3_y0 = f_s_dadda_rca24_and_20_3_y0;
  assign f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_19_4_y0 = f_s_dadda_rca24_and_19_4_y0;
  assign f_s_dadda_rca24_fa8_y0 = f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_21_2_y0 ^ f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_20_3_y0;
  assign f_s_dadda_rca24_fa8_y1 = f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_21_2_y0 & f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_20_3_y0;
  assign f_s_dadda_rca24_fa8_y2 = f_s_dadda_rca24_fa8_y0 ^ f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_19_4_y0;
  assign f_s_dadda_rca24_fa8_y3 = f_s_dadda_rca24_fa8_y0 & f_s_dadda_rca24_fa8_f_s_dadda_rca24_and_19_4_y0;
  assign f_s_dadda_rca24_fa8_y4 = f_s_dadda_rca24_fa8_y1 | f_s_dadda_rca24_fa8_y3;
  assign f_s_dadda_rca24_and_18_5_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_18_5_y0 = f_s_dadda_rca24_and_18_5_a_18 & f_s_dadda_rca24_and_18_5_b_5;
  assign f_s_dadda_rca24_and_17_6_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_17_6_y0 = f_s_dadda_rca24_and_17_6_a_17 & f_s_dadda_rca24_and_17_6_b_6;
  assign f_s_dadda_rca24_and_16_7_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_16_7_y0 = f_s_dadda_rca24_and_16_7_a_16 & f_s_dadda_rca24_and_16_7_b_7;
  assign f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_18_5_y0 = f_s_dadda_rca24_and_18_5_y0;
  assign f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_17_6_y0 = f_s_dadda_rca24_and_17_6_y0;
  assign f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_16_7_y0 = f_s_dadda_rca24_and_16_7_y0;
  assign f_s_dadda_rca24_fa9_y0 = f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_18_5_y0 ^ f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_17_6_y0;
  assign f_s_dadda_rca24_fa9_y1 = f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_18_5_y0 & f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_17_6_y0;
  assign f_s_dadda_rca24_fa9_y2 = f_s_dadda_rca24_fa9_y0 ^ f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_16_7_y0;
  assign f_s_dadda_rca24_fa9_y3 = f_s_dadda_rca24_fa9_y0 & f_s_dadda_rca24_fa9_f_s_dadda_rca24_and_16_7_y0;
  assign f_s_dadda_rca24_fa9_y4 = f_s_dadda_rca24_fa9_y1 | f_s_dadda_rca24_fa9_y3;
  assign f_s_dadda_rca24_and_15_8_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_15_8_y0 = f_s_dadda_rca24_and_15_8_a_15 & f_s_dadda_rca24_and_15_8_b_8;
  assign f_s_dadda_rca24_and_14_9_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_14_9_y0 = f_s_dadda_rca24_and_14_9_a_14 & f_s_dadda_rca24_and_14_9_b_9;
  assign f_s_dadda_rca24_ha4_f_s_dadda_rca24_and_15_8_y0 = f_s_dadda_rca24_and_15_8_y0;
  assign f_s_dadda_rca24_ha4_f_s_dadda_rca24_and_14_9_y0 = f_s_dadda_rca24_and_14_9_y0;
  assign f_s_dadda_rca24_ha4_y0 = f_s_dadda_rca24_ha4_f_s_dadda_rca24_and_15_8_y0 ^ f_s_dadda_rca24_ha4_f_s_dadda_rca24_and_14_9_y0;
  assign f_s_dadda_rca24_ha4_y1 = f_s_dadda_rca24_ha4_f_s_dadda_rca24_and_15_8_y0 & f_s_dadda_rca24_ha4_f_s_dadda_rca24_and_14_9_y0;
  assign f_s_dadda_rca24_fa10_f_s_dadda_rca24_ha4_y1 = f_s_dadda_rca24_ha4_y1;
  assign f_s_dadda_rca24_fa10_f_s_dadda_rca24_fa9_y4 = f_s_dadda_rca24_fa9_y4;
  assign f_s_dadda_rca24_fa10_f_s_dadda_rca24_fa8_y4 = f_s_dadda_rca24_fa8_y4;
  assign f_s_dadda_rca24_fa10_y0 = f_s_dadda_rca24_fa10_f_s_dadda_rca24_ha4_y1 ^ f_s_dadda_rca24_fa10_f_s_dadda_rca24_fa9_y4;
  assign f_s_dadda_rca24_fa10_y1 = f_s_dadda_rca24_fa10_f_s_dadda_rca24_ha4_y1 & f_s_dadda_rca24_fa10_f_s_dadda_rca24_fa9_y4;
  assign f_s_dadda_rca24_fa10_y2 = f_s_dadda_rca24_fa10_y0 ^ f_s_dadda_rca24_fa10_f_s_dadda_rca24_fa8_y4;
  assign f_s_dadda_rca24_fa10_y3 = f_s_dadda_rca24_fa10_y0 & f_s_dadda_rca24_fa10_f_s_dadda_rca24_fa8_y4;
  assign f_s_dadda_rca24_fa10_y4 = f_s_dadda_rca24_fa10_y1 | f_s_dadda_rca24_fa10_y3;
  assign f_s_dadda_rca24_fa11_f_s_dadda_rca24_fa7_y4 = f_s_dadda_rca24_fa7_y4;
  assign f_s_dadda_rca24_fa11_f_s_dadda_rca24_fa6_y4 = f_s_dadda_rca24_fa6_y4;
  assign f_s_dadda_rca24_fa11_constant_wire_1 = constant_wire_1;
  assign f_s_dadda_rca24_fa11_y0 = f_s_dadda_rca24_fa11_f_s_dadda_rca24_fa7_y4 ^ f_s_dadda_rca24_fa11_f_s_dadda_rca24_fa6_y4;
  assign f_s_dadda_rca24_fa11_y1 = f_s_dadda_rca24_fa11_f_s_dadda_rca24_fa7_y4 & f_s_dadda_rca24_fa11_f_s_dadda_rca24_fa6_y4;
  assign f_s_dadda_rca24_fa11_y2 = f_s_dadda_rca24_fa11_y0 ^ f_s_dadda_rca24_fa11_constant_wire_1;
  assign f_s_dadda_rca24_fa11_y3 = f_s_dadda_rca24_fa11_y0 & f_s_dadda_rca24_fa11_constant_wire_1;
  assign f_s_dadda_rca24_fa11_y4 = f_s_dadda_rca24_fa11_y1 | f_s_dadda_rca24_fa11_y3;
  assign f_s_dadda_rca24_nand_23_1_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_1_b_1 = b_1;
  assign f_s_dadda_rca24_nand_23_1_y0 = ~(f_s_dadda_rca24_nand_23_1_a_23 & f_s_dadda_rca24_nand_23_1_b_1);
  assign f_s_dadda_rca24_and_22_2_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_22_2_y0 = f_s_dadda_rca24_and_22_2_a_22 & f_s_dadda_rca24_and_22_2_b_2;
  assign f_s_dadda_rca24_and_21_3_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_21_3_y0 = f_s_dadda_rca24_and_21_3_a_21 & f_s_dadda_rca24_and_21_3_b_3;
  assign f_s_dadda_rca24_fa12_f_s_dadda_rca24_nand_23_1_y0 = f_s_dadda_rca24_nand_23_1_y0;
  assign f_s_dadda_rca24_fa12_f_s_dadda_rca24_and_22_2_y0 = f_s_dadda_rca24_and_22_2_y0;
  assign f_s_dadda_rca24_fa12_f_s_dadda_rca24_and_21_3_y0 = f_s_dadda_rca24_and_21_3_y0;
  assign f_s_dadda_rca24_fa12_y0 = f_s_dadda_rca24_fa12_f_s_dadda_rca24_nand_23_1_y0 ^ f_s_dadda_rca24_fa12_f_s_dadda_rca24_and_22_2_y0;
  assign f_s_dadda_rca24_fa12_y1 = f_s_dadda_rca24_fa12_f_s_dadda_rca24_nand_23_1_y0 & f_s_dadda_rca24_fa12_f_s_dadda_rca24_and_22_2_y0;
  assign f_s_dadda_rca24_fa12_y2 = f_s_dadda_rca24_fa12_y0 ^ f_s_dadda_rca24_fa12_f_s_dadda_rca24_and_21_3_y0;
  assign f_s_dadda_rca24_fa12_y3 = f_s_dadda_rca24_fa12_y0 & f_s_dadda_rca24_fa12_f_s_dadda_rca24_and_21_3_y0;
  assign f_s_dadda_rca24_fa12_y4 = f_s_dadda_rca24_fa12_y1 | f_s_dadda_rca24_fa12_y3;
  assign f_s_dadda_rca24_and_20_4_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_20_4_y0 = f_s_dadda_rca24_and_20_4_a_20 & f_s_dadda_rca24_and_20_4_b_4;
  assign f_s_dadda_rca24_and_19_5_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_19_5_y0 = f_s_dadda_rca24_and_19_5_a_19 & f_s_dadda_rca24_and_19_5_b_5;
  assign f_s_dadda_rca24_and_18_6_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_18_6_y0 = f_s_dadda_rca24_and_18_6_a_18 & f_s_dadda_rca24_and_18_6_b_6;
  assign f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_20_4_y0 = f_s_dadda_rca24_and_20_4_y0;
  assign f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_19_5_y0 = f_s_dadda_rca24_and_19_5_y0;
  assign f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_18_6_y0 = f_s_dadda_rca24_and_18_6_y0;
  assign f_s_dadda_rca24_fa13_y0 = f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_20_4_y0 ^ f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_19_5_y0;
  assign f_s_dadda_rca24_fa13_y1 = f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_20_4_y0 & f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_19_5_y0;
  assign f_s_dadda_rca24_fa13_y2 = f_s_dadda_rca24_fa13_y0 ^ f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_18_6_y0;
  assign f_s_dadda_rca24_fa13_y3 = f_s_dadda_rca24_fa13_y0 & f_s_dadda_rca24_fa13_f_s_dadda_rca24_and_18_6_y0;
  assign f_s_dadda_rca24_fa13_y4 = f_s_dadda_rca24_fa13_y1 | f_s_dadda_rca24_fa13_y3;
  assign f_s_dadda_rca24_and_17_7_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_17_7_y0 = f_s_dadda_rca24_and_17_7_a_17 & f_s_dadda_rca24_and_17_7_b_7;
  assign f_s_dadda_rca24_and_16_8_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_16_8_y0 = f_s_dadda_rca24_and_16_8_a_16 & f_s_dadda_rca24_and_16_8_b_8;
  assign f_s_dadda_rca24_and_15_9_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_15_9_y0 = f_s_dadda_rca24_and_15_9_a_15 & f_s_dadda_rca24_and_15_9_b_9;
  assign f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_17_7_y0 = f_s_dadda_rca24_and_17_7_y0;
  assign f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_16_8_y0 = f_s_dadda_rca24_and_16_8_y0;
  assign f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_15_9_y0 = f_s_dadda_rca24_and_15_9_y0;
  assign f_s_dadda_rca24_fa14_y0 = f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_17_7_y0 ^ f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_16_8_y0;
  assign f_s_dadda_rca24_fa14_y1 = f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_17_7_y0 & f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_16_8_y0;
  assign f_s_dadda_rca24_fa14_y2 = f_s_dadda_rca24_fa14_y0 ^ f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_15_9_y0;
  assign f_s_dadda_rca24_fa14_y3 = f_s_dadda_rca24_fa14_y0 & f_s_dadda_rca24_fa14_f_s_dadda_rca24_and_15_9_y0;
  assign f_s_dadda_rca24_fa14_y4 = f_s_dadda_rca24_fa14_y1 | f_s_dadda_rca24_fa14_y3;
  assign f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa14_y4 = f_s_dadda_rca24_fa14_y4;
  assign f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa13_y4 = f_s_dadda_rca24_fa13_y4;
  assign f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa12_y4 = f_s_dadda_rca24_fa12_y4;
  assign f_s_dadda_rca24_fa15_y0 = f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa14_y4 ^ f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa13_y4;
  assign f_s_dadda_rca24_fa15_y1 = f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa14_y4 & f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa13_y4;
  assign f_s_dadda_rca24_fa15_y2 = f_s_dadda_rca24_fa15_y0 ^ f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa12_y4;
  assign f_s_dadda_rca24_fa15_y3 = f_s_dadda_rca24_fa15_y0 & f_s_dadda_rca24_fa15_f_s_dadda_rca24_fa12_y4;
  assign f_s_dadda_rca24_fa15_y4 = f_s_dadda_rca24_fa15_y1 | f_s_dadda_rca24_fa15_y3;
  assign f_s_dadda_rca24_nand_23_2_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_2_b_2 = b_2;
  assign f_s_dadda_rca24_nand_23_2_y0 = ~(f_s_dadda_rca24_nand_23_2_a_23 & f_s_dadda_rca24_nand_23_2_b_2);
  assign f_s_dadda_rca24_fa16_f_s_dadda_rca24_fa11_y4 = f_s_dadda_rca24_fa11_y4;
  assign f_s_dadda_rca24_fa16_f_s_dadda_rca24_fa10_y4 = f_s_dadda_rca24_fa10_y4;
  assign f_s_dadda_rca24_fa16_f_s_dadda_rca24_nand_23_2_y0 = f_s_dadda_rca24_nand_23_2_y0;
  assign f_s_dadda_rca24_fa16_y0 = f_s_dadda_rca24_fa16_f_s_dadda_rca24_fa11_y4 ^ f_s_dadda_rca24_fa16_f_s_dadda_rca24_fa10_y4;
  assign f_s_dadda_rca24_fa16_y1 = f_s_dadda_rca24_fa16_f_s_dadda_rca24_fa11_y4 & f_s_dadda_rca24_fa16_f_s_dadda_rca24_fa10_y4;
  assign f_s_dadda_rca24_fa16_y2 = f_s_dadda_rca24_fa16_y0 ^ f_s_dadda_rca24_fa16_f_s_dadda_rca24_nand_23_2_y0;
  assign f_s_dadda_rca24_fa16_y3 = f_s_dadda_rca24_fa16_y0 & f_s_dadda_rca24_fa16_f_s_dadda_rca24_nand_23_2_y0;
  assign f_s_dadda_rca24_fa16_y4 = f_s_dadda_rca24_fa16_y1 | f_s_dadda_rca24_fa16_y3;
  assign f_s_dadda_rca24_and_22_3_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_22_3_y0 = f_s_dadda_rca24_and_22_3_a_22 & f_s_dadda_rca24_and_22_3_b_3;
  assign f_s_dadda_rca24_and_21_4_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_21_4_y0 = f_s_dadda_rca24_and_21_4_a_21 & f_s_dadda_rca24_and_21_4_b_4;
  assign f_s_dadda_rca24_and_20_5_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_20_5_y0 = f_s_dadda_rca24_and_20_5_a_20 & f_s_dadda_rca24_and_20_5_b_5;
  assign f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_22_3_y0 = f_s_dadda_rca24_and_22_3_y0;
  assign f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_21_4_y0 = f_s_dadda_rca24_and_21_4_y0;
  assign f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_20_5_y0 = f_s_dadda_rca24_and_20_5_y0;
  assign f_s_dadda_rca24_fa17_y0 = f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_22_3_y0 ^ f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_21_4_y0;
  assign f_s_dadda_rca24_fa17_y1 = f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_22_3_y0 & f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_21_4_y0;
  assign f_s_dadda_rca24_fa17_y2 = f_s_dadda_rca24_fa17_y0 ^ f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_20_5_y0;
  assign f_s_dadda_rca24_fa17_y3 = f_s_dadda_rca24_fa17_y0 & f_s_dadda_rca24_fa17_f_s_dadda_rca24_and_20_5_y0;
  assign f_s_dadda_rca24_fa17_y4 = f_s_dadda_rca24_fa17_y1 | f_s_dadda_rca24_fa17_y3;
  assign f_s_dadda_rca24_and_19_6_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_19_6_y0 = f_s_dadda_rca24_and_19_6_a_19 & f_s_dadda_rca24_and_19_6_b_6;
  assign f_s_dadda_rca24_and_18_7_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_18_7_y0 = f_s_dadda_rca24_and_18_7_a_18 & f_s_dadda_rca24_and_18_7_b_7;
  assign f_s_dadda_rca24_and_17_8_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_17_8_y0 = f_s_dadda_rca24_and_17_8_a_17 & f_s_dadda_rca24_and_17_8_b_8;
  assign f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_19_6_y0 = f_s_dadda_rca24_and_19_6_y0;
  assign f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_18_7_y0 = f_s_dadda_rca24_and_18_7_y0;
  assign f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_17_8_y0 = f_s_dadda_rca24_and_17_8_y0;
  assign f_s_dadda_rca24_fa18_y0 = f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_19_6_y0 ^ f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_18_7_y0;
  assign f_s_dadda_rca24_fa18_y1 = f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_19_6_y0 & f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_18_7_y0;
  assign f_s_dadda_rca24_fa18_y2 = f_s_dadda_rca24_fa18_y0 ^ f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_17_8_y0;
  assign f_s_dadda_rca24_fa18_y3 = f_s_dadda_rca24_fa18_y0 & f_s_dadda_rca24_fa18_f_s_dadda_rca24_and_17_8_y0;
  assign f_s_dadda_rca24_fa18_y4 = f_s_dadda_rca24_fa18_y1 | f_s_dadda_rca24_fa18_y3;
  assign f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa18_y4 = f_s_dadda_rca24_fa18_y4;
  assign f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa17_y4 = f_s_dadda_rca24_fa17_y4;
  assign f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa16_y4 = f_s_dadda_rca24_fa16_y4;
  assign f_s_dadda_rca24_fa19_y0 = f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa18_y4 ^ f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa17_y4;
  assign f_s_dadda_rca24_fa19_y1 = f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa18_y4 & f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa17_y4;
  assign f_s_dadda_rca24_fa19_y2 = f_s_dadda_rca24_fa19_y0 ^ f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa16_y4;
  assign f_s_dadda_rca24_fa19_y3 = f_s_dadda_rca24_fa19_y0 & f_s_dadda_rca24_fa19_f_s_dadda_rca24_fa16_y4;
  assign f_s_dadda_rca24_fa19_y4 = f_s_dadda_rca24_fa19_y1 | f_s_dadda_rca24_fa19_y3;
  assign f_s_dadda_rca24_nand_23_3_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_3_b_3 = b_3;
  assign f_s_dadda_rca24_nand_23_3_y0 = ~(f_s_dadda_rca24_nand_23_3_a_23 & f_s_dadda_rca24_nand_23_3_b_3);
  assign f_s_dadda_rca24_and_22_4_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_22_4_y0 = f_s_dadda_rca24_and_22_4_a_22 & f_s_dadda_rca24_and_22_4_b_4;
  assign f_s_dadda_rca24_fa20_f_s_dadda_rca24_fa15_y4 = f_s_dadda_rca24_fa15_y4;
  assign f_s_dadda_rca24_fa20_f_s_dadda_rca24_nand_23_3_y0 = f_s_dadda_rca24_nand_23_3_y0;
  assign f_s_dadda_rca24_fa20_f_s_dadda_rca24_and_22_4_y0 = f_s_dadda_rca24_and_22_4_y0;
  assign f_s_dadda_rca24_fa20_y0 = f_s_dadda_rca24_fa20_f_s_dadda_rca24_fa15_y4 ^ f_s_dadda_rca24_fa20_f_s_dadda_rca24_nand_23_3_y0;
  assign f_s_dadda_rca24_fa20_y1 = f_s_dadda_rca24_fa20_f_s_dadda_rca24_fa15_y4 & f_s_dadda_rca24_fa20_f_s_dadda_rca24_nand_23_3_y0;
  assign f_s_dadda_rca24_fa20_y2 = f_s_dadda_rca24_fa20_y0 ^ f_s_dadda_rca24_fa20_f_s_dadda_rca24_and_22_4_y0;
  assign f_s_dadda_rca24_fa20_y3 = f_s_dadda_rca24_fa20_y0 & f_s_dadda_rca24_fa20_f_s_dadda_rca24_and_22_4_y0;
  assign f_s_dadda_rca24_fa20_y4 = f_s_dadda_rca24_fa20_y1 | f_s_dadda_rca24_fa20_y3;
  assign f_s_dadda_rca24_and_21_5_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_21_5_y0 = f_s_dadda_rca24_and_21_5_a_21 & f_s_dadda_rca24_and_21_5_b_5;
  assign f_s_dadda_rca24_and_20_6_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_20_6_y0 = f_s_dadda_rca24_and_20_6_a_20 & f_s_dadda_rca24_and_20_6_b_6;
  assign f_s_dadda_rca24_and_19_7_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_19_7_y0 = f_s_dadda_rca24_and_19_7_a_19 & f_s_dadda_rca24_and_19_7_b_7;
  assign f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_21_5_y0 = f_s_dadda_rca24_and_21_5_y0;
  assign f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_20_6_y0 = f_s_dadda_rca24_and_20_6_y0;
  assign f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_19_7_y0 = f_s_dadda_rca24_and_19_7_y0;
  assign f_s_dadda_rca24_fa21_y0 = f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_21_5_y0 ^ f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_20_6_y0;
  assign f_s_dadda_rca24_fa21_y1 = f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_21_5_y0 & f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_20_6_y0;
  assign f_s_dadda_rca24_fa21_y2 = f_s_dadda_rca24_fa21_y0 ^ f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_19_7_y0;
  assign f_s_dadda_rca24_fa21_y3 = f_s_dadda_rca24_fa21_y0 & f_s_dadda_rca24_fa21_f_s_dadda_rca24_and_19_7_y0;
  assign f_s_dadda_rca24_fa21_y4 = f_s_dadda_rca24_fa21_y1 | f_s_dadda_rca24_fa21_y3;
  assign f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa21_y4 = f_s_dadda_rca24_fa21_y4;
  assign f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa20_y4 = f_s_dadda_rca24_fa20_y4;
  assign f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa19_y4 = f_s_dadda_rca24_fa19_y4;
  assign f_s_dadda_rca24_fa22_y0 = f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa21_y4 ^ f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa20_y4;
  assign f_s_dadda_rca24_fa22_y1 = f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa21_y4 & f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa20_y4;
  assign f_s_dadda_rca24_fa22_y2 = f_s_dadda_rca24_fa22_y0 ^ f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa19_y4;
  assign f_s_dadda_rca24_fa22_y3 = f_s_dadda_rca24_fa22_y0 & f_s_dadda_rca24_fa22_f_s_dadda_rca24_fa19_y4;
  assign f_s_dadda_rca24_fa22_y4 = f_s_dadda_rca24_fa22_y1 | f_s_dadda_rca24_fa22_y3;
  assign f_s_dadda_rca24_nand_23_4_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_4_b_4 = b_4;
  assign f_s_dadda_rca24_nand_23_4_y0 = ~(f_s_dadda_rca24_nand_23_4_a_23 & f_s_dadda_rca24_nand_23_4_b_4);
  assign f_s_dadda_rca24_and_22_5_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_22_5_y0 = f_s_dadda_rca24_and_22_5_a_22 & f_s_dadda_rca24_and_22_5_b_5;
  assign f_s_dadda_rca24_and_21_6_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_21_6_y0 = f_s_dadda_rca24_and_21_6_a_21 & f_s_dadda_rca24_and_21_6_b_6;
  assign f_s_dadda_rca24_fa23_f_s_dadda_rca24_nand_23_4_y0 = f_s_dadda_rca24_nand_23_4_y0;
  assign f_s_dadda_rca24_fa23_f_s_dadda_rca24_and_22_5_y0 = f_s_dadda_rca24_and_22_5_y0;
  assign f_s_dadda_rca24_fa23_f_s_dadda_rca24_and_21_6_y0 = f_s_dadda_rca24_and_21_6_y0;
  assign f_s_dadda_rca24_fa23_y0 = f_s_dadda_rca24_fa23_f_s_dadda_rca24_nand_23_4_y0 ^ f_s_dadda_rca24_fa23_f_s_dadda_rca24_and_22_5_y0;
  assign f_s_dadda_rca24_fa23_y1 = f_s_dadda_rca24_fa23_f_s_dadda_rca24_nand_23_4_y0 & f_s_dadda_rca24_fa23_f_s_dadda_rca24_and_22_5_y0;
  assign f_s_dadda_rca24_fa23_y2 = f_s_dadda_rca24_fa23_y0 ^ f_s_dadda_rca24_fa23_f_s_dadda_rca24_and_21_6_y0;
  assign f_s_dadda_rca24_fa23_y3 = f_s_dadda_rca24_fa23_y0 & f_s_dadda_rca24_fa23_f_s_dadda_rca24_and_21_6_y0;
  assign f_s_dadda_rca24_fa23_y4 = f_s_dadda_rca24_fa23_y1 | f_s_dadda_rca24_fa23_y3;
  assign f_s_dadda_rca24_nand_23_5_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_5_b_5 = b_5;
  assign f_s_dadda_rca24_nand_23_5_y0 = ~(f_s_dadda_rca24_nand_23_5_a_23 & f_s_dadda_rca24_nand_23_5_b_5);
  assign f_s_dadda_rca24_fa24_f_s_dadda_rca24_fa23_y4 = f_s_dadda_rca24_fa23_y4;
  assign f_s_dadda_rca24_fa24_f_s_dadda_rca24_fa22_y4 = f_s_dadda_rca24_fa22_y4;
  assign f_s_dadda_rca24_fa24_f_s_dadda_rca24_nand_23_5_y0 = f_s_dadda_rca24_nand_23_5_y0;
  assign f_s_dadda_rca24_fa24_y0 = f_s_dadda_rca24_fa24_f_s_dadda_rca24_fa23_y4 ^ f_s_dadda_rca24_fa24_f_s_dadda_rca24_fa22_y4;
  assign f_s_dadda_rca24_fa24_y1 = f_s_dadda_rca24_fa24_f_s_dadda_rca24_fa23_y4 & f_s_dadda_rca24_fa24_f_s_dadda_rca24_fa22_y4;
  assign f_s_dadda_rca24_fa24_y2 = f_s_dadda_rca24_fa24_y0 ^ f_s_dadda_rca24_fa24_f_s_dadda_rca24_nand_23_5_y0;
  assign f_s_dadda_rca24_fa24_y3 = f_s_dadda_rca24_fa24_y0 & f_s_dadda_rca24_fa24_f_s_dadda_rca24_nand_23_5_y0;
  assign f_s_dadda_rca24_fa24_y4 = f_s_dadda_rca24_fa24_y1 | f_s_dadda_rca24_fa24_y3;
  assign f_s_dadda_rca24_and_6_0_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_6_0_y0 = f_s_dadda_rca24_and_6_0_a_6 & f_s_dadda_rca24_and_6_0_b_0;
  assign f_s_dadda_rca24_and_5_1_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_5_1_y0 = f_s_dadda_rca24_and_5_1_a_5 & f_s_dadda_rca24_and_5_1_b_1;
  assign f_s_dadda_rca24_ha5_f_s_dadda_rca24_and_6_0_y0 = f_s_dadda_rca24_and_6_0_y0;
  assign f_s_dadda_rca24_ha5_f_s_dadda_rca24_and_5_1_y0 = f_s_dadda_rca24_and_5_1_y0;
  assign f_s_dadda_rca24_ha5_y0 = f_s_dadda_rca24_ha5_f_s_dadda_rca24_and_6_0_y0 ^ f_s_dadda_rca24_ha5_f_s_dadda_rca24_and_5_1_y0;
  assign f_s_dadda_rca24_ha5_y1 = f_s_dadda_rca24_ha5_f_s_dadda_rca24_and_6_0_y0 & f_s_dadda_rca24_ha5_f_s_dadda_rca24_and_5_1_y0;
  assign f_s_dadda_rca24_and_7_0_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_7_0_y0 = f_s_dadda_rca24_and_7_0_a_7 & f_s_dadda_rca24_and_7_0_b_0;
  assign f_s_dadda_rca24_and_6_1_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_6_1_y0 = f_s_dadda_rca24_and_6_1_a_6 & f_s_dadda_rca24_and_6_1_b_1;
  assign f_s_dadda_rca24_fa25_f_s_dadda_rca24_ha5_y1 = f_s_dadda_rca24_ha5_y1;
  assign f_s_dadda_rca24_fa25_f_s_dadda_rca24_and_7_0_y0 = f_s_dadda_rca24_and_7_0_y0;
  assign f_s_dadda_rca24_fa25_f_s_dadda_rca24_and_6_1_y0 = f_s_dadda_rca24_and_6_1_y0;
  assign f_s_dadda_rca24_fa25_y0 = f_s_dadda_rca24_fa25_f_s_dadda_rca24_ha5_y1 ^ f_s_dadda_rca24_fa25_f_s_dadda_rca24_and_7_0_y0;
  assign f_s_dadda_rca24_fa25_y1 = f_s_dadda_rca24_fa25_f_s_dadda_rca24_ha5_y1 & f_s_dadda_rca24_fa25_f_s_dadda_rca24_and_7_0_y0;
  assign f_s_dadda_rca24_fa25_y2 = f_s_dadda_rca24_fa25_y0 ^ f_s_dadda_rca24_fa25_f_s_dadda_rca24_and_6_1_y0;
  assign f_s_dadda_rca24_fa25_y3 = f_s_dadda_rca24_fa25_y0 & f_s_dadda_rca24_fa25_f_s_dadda_rca24_and_6_1_y0;
  assign f_s_dadda_rca24_fa25_y4 = f_s_dadda_rca24_fa25_y1 | f_s_dadda_rca24_fa25_y3;
  assign f_s_dadda_rca24_and_5_2_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_5_2_y0 = f_s_dadda_rca24_and_5_2_a_5 & f_s_dadda_rca24_and_5_2_b_2;
  assign f_s_dadda_rca24_and_4_3_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_4_3_y0 = f_s_dadda_rca24_and_4_3_a_4 & f_s_dadda_rca24_and_4_3_b_3;
  assign f_s_dadda_rca24_ha6_f_s_dadda_rca24_and_5_2_y0 = f_s_dadda_rca24_and_5_2_y0;
  assign f_s_dadda_rca24_ha6_f_s_dadda_rca24_and_4_3_y0 = f_s_dadda_rca24_and_4_3_y0;
  assign f_s_dadda_rca24_ha6_y0 = f_s_dadda_rca24_ha6_f_s_dadda_rca24_and_5_2_y0 ^ f_s_dadda_rca24_ha6_f_s_dadda_rca24_and_4_3_y0;
  assign f_s_dadda_rca24_ha6_y1 = f_s_dadda_rca24_ha6_f_s_dadda_rca24_and_5_2_y0 & f_s_dadda_rca24_ha6_f_s_dadda_rca24_and_4_3_y0;
  assign f_s_dadda_rca24_and_8_0_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_8_0_y0 = f_s_dadda_rca24_and_8_0_a_8 & f_s_dadda_rca24_and_8_0_b_0;
  assign f_s_dadda_rca24_fa26_f_s_dadda_rca24_ha6_y1 = f_s_dadda_rca24_ha6_y1;
  assign f_s_dadda_rca24_fa26_f_s_dadda_rca24_fa25_y4 = f_s_dadda_rca24_fa25_y4;
  assign f_s_dadda_rca24_fa26_f_s_dadda_rca24_and_8_0_y0 = f_s_dadda_rca24_and_8_0_y0;
  assign f_s_dadda_rca24_fa26_y0 = f_s_dadda_rca24_fa26_f_s_dadda_rca24_ha6_y1 ^ f_s_dadda_rca24_fa26_f_s_dadda_rca24_fa25_y4;
  assign f_s_dadda_rca24_fa26_y1 = f_s_dadda_rca24_fa26_f_s_dadda_rca24_ha6_y1 & f_s_dadda_rca24_fa26_f_s_dadda_rca24_fa25_y4;
  assign f_s_dadda_rca24_fa26_y2 = f_s_dadda_rca24_fa26_y0 ^ f_s_dadda_rca24_fa26_f_s_dadda_rca24_and_8_0_y0;
  assign f_s_dadda_rca24_fa26_y3 = f_s_dadda_rca24_fa26_y0 & f_s_dadda_rca24_fa26_f_s_dadda_rca24_and_8_0_y0;
  assign f_s_dadda_rca24_fa26_y4 = f_s_dadda_rca24_fa26_y1 | f_s_dadda_rca24_fa26_y3;
  assign f_s_dadda_rca24_and_7_1_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_7_1_y0 = f_s_dadda_rca24_and_7_1_a_7 & f_s_dadda_rca24_and_7_1_b_1;
  assign f_s_dadda_rca24_and_6_2_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_6_2_y0 = f_s_dadda_rca24_and_6_2_a_6 & f_s_dadda_rca24_and_6_2_b_2;
  assign f_s_dadda_rca24_and_5_3_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_5_3_y0 = f_s_dadda_rca24_and_5_3_a_5 & f_s_dadda_rca24_and_5_3_b_3;
  assign f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_7_1_y0 = f_s_dadda_rca24_and_7_1_y0;
  assign f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_6_2_y0 = f_s_dadda_rca24_and_6_2_y0;
  assign f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_5_3_y0 = f_s_dadda_rca24_and_5_3_y0;
  assign f_s_dadda_rca24_fa27_y0 = f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_7_1_y0 ^ f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_6_2_y0;
  assign f_s_dadda_rca24_fa27_y1 = f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_7_1_y0 & f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_6_2_y0;
  assign f_s_dadda_rca24_fa27_y2 = f_s_dadda_rca24_fa27_y0 ^ f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_5_3_y0;
  assign f_s_dadda_rca24_fa27_y3 = f_s_dadda_rca24_fa27_y0 & f_s_dadda_rca24_fa27_f_s_dadda_rca24_and_5_3_y0;
  assign f_s_dadda_rca24_fa27_y4 = f_s_dadda_rca24_fa27_y1 | f_s_dadda_rca24_fa27_y3;
  assign f_s_dadda_rca24_and_4_4_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_4_4_y0 = f_s_dadda_rca24_and_4_4_a_4 & f_s_dadda_rca24_and_4_4_b_4;
  assign f_s_dadda_rca24_and_3_5_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_3_5_y0 = f_s_dadda_rca24_and_3_5_a_3 & f_s_dadda_rca24_and_3_5_b_5;
  assign f_s_dadda_rca24_ha7_f_s_dadda_rca24_and_4_4_y0 = f_s_dadda_rca24_and_4_4_y0;
  assign f_s_dadda_rca24_ha7_f_s_dadda_rca24_and_3_5_y0 = f_s_dadda_rca24_and_3_5_y0;
  assign f_s_dadda_rca24_ha7_y0 = f_s_dadda_rca24_ha7_f_s_dadda_rca24_and_4_4_y0 ^ f_s_dadda_rca24_ha7_f_s_dadda_rca24_and_3_5_y0;
  assign f_s_dadda_rca24_ha7_y1 = f_s_dadda_rca24_ha7_f_s_dadda_rca24_and_4_4_y0 & f_s_dadda_rca24_ha7_f_s_dadda_rca24_and_3_5_y0;
  assign f_s_dadda_rca24_fa28_f_s_dadda_rca24_ha7_y1 = f_s_dadda_rca24_ha7_y1;
  assign f_s_dadda_rca24_fa28_f_s_dadda_rca24_fa27_y4 = f_s_dadda_rca24_fa27_y4;
  assign f_s_dadda_rca24_fa28_f_s_dadda_rca24_fa26_y4 = f_s_dadda_rca24_fa26_y4;
  assign f_s_dadda_rca24_fa28_y0 = f_s_dadda_rca24_fa28_f_s_dadda_rca24_ha7_y1 ^ f_s_dadda_rca24_fa28_f_s_dadda_rca24_fa27_y4;
  assign f_s_dadda_rca24_fa28_y1 = f_s_dadda_rca24_fa28_f_s_dadda_rca24_ha7_y1 & f_s_dadda_rca24_fa28_f_s_dadda_rca24_fa27_y4;
  assign f_s_dadda_rca24_fa28_y2 = f_s_dadda_rca24_fa28_y0 ^ f_s_dadda_rca24_fa28_f_s_dadda_rca24_fa26_y4;
  assign f_s_dadda_rca24_fa28_y3 = f_s_dadda_rca24_fa28_y0 & f_s_dadda_rca24_fa28_f_s_dadda_rca24_fa26_y4;
  assign f_s_dadda_rca24_fa28_y4 = f_s_dadda_rca24_fa28_y1 | f_s_dadda_rca24_fa28_y3;
  assign f_s_dadda_rca24_and_9_0_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_9_0_y0 = f_s_dadda_rca24_and_9_0_a_9 & f_s_dadda_rca24_and_9_0_b_0;
  assign f_s_dadda_rca24_and_8_1_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_8_1_y0 = f_s_dadda_rca24_and_8_1_a_8 & f_s_dadda_rca24_and_8_1_b_1;
  assign f_s_dadda_rca24_and_7_2_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_7_2_y0 = f_s_dadda_rca24_and_7_2_a_7 & f_s_dadda_rca24_and_7_2_b_2;
  assign f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_9_0_y0 = f_s_dadda_rca24_and_9_0_y0;
  assign f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_8_1_y0 = f_s_dadda_rca24_and_8_1_y0;
  assign f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_7_2_y0 = f_s_dadda_rca24_and_7_2_y0;
  assign f_s_dadda_rca24_fa29_y0 = f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_9_0_y0 ^ f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_8_1_y0;
  assign f_s_dadda_rca24_fa29_y1 = f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_9_0_y0 & f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_8_1_y0;
  assign f_s_dadda_rca24_fa29_y2 = f_s_dadda_rca24_fa29_y0 ^ f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_7_2_y0;
  assign f_s_dadda_rca24_fa29_y3 = f_s_dadda_rca24_fa29_y0 & f_s_dadda_rca24_fa29_f_s_dadda_rca24_and_7_2_y0;
  assign f_s_dadda_rca24_fa29_y4 = f_s_dadda_rca24_fa29_y1 | f_s_dadda_rca24_fa29_y3;
  assign f_s_dadda_rca24_and_6_3_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_6_3_y0 = f_s_dadda_rca24_and_6_3_a_6 & f_s_dadda_rca24_and_6_3_b_3;
  assign f_s_dadda_rca24_and_5_4_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_5_4_y0 = f_s_dadda_rca24_and_5_4_a_5 & f_s_dadda_rca24_and_5_4_b_4;
  assign f_s_dadda_rca24_and_4_5_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_4_5_y0 = f_s_dadda_rca24_and_4_5_a_4 & f_s_dadda_rca24_and_4_5_b_5;
  assign f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_6_3_y0 = f_s_dadda_rca24_and_6_3_y0;
  assign f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_5_4_y0 = f_s_dadda_rca24_and_5_4_y0;
  assign f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_4_5_y0 = f_s_dadda_rca24_and_4_5_y0;
  assign f_s_dadda_rca24_fa30_y0 = f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_6_3_y0 ^ f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_5_4_y0;
  assign f_s_dadda_rca24_fa30_y1 = f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_6_3_y0 & f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_5_4_y0;
  assign f_s_dadda_rca24_fa30_y2 = f_s_dadda_rca24_fa30_y0 ^ f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_4_5_y0;
  assign f_s_dadda_rca24_fa30_y3 = f_s_dadda_rca24_fa30_y0 & f_s_dadda_rca24_fa30_f_s_dadda_rca24_and_4_5_y0;
  assign f_s_dadda_rca24_fa30_y4 = f_s_dadda_rca24_fa30_y1 | f_s_dadda_rca24_fa30_y3;
  assign f_s_dadda_rca24_and_3_6_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_3_6_y0 = f_s_dadda_rca24_and_3_6_a_3 & f_s_dadda_rca24_and_3_6_b_6;
  assign f_s_dadda_rca24_and_2_7_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_2_7_y0 = f_s_dadda_rca24_and_2_7_a_2 & f_s_dadda_rca24_and_2_7_b_7;
  assign f_s_dadda_rca24_ha8_f_s_dadda_rca24_and_3_6_y0 = f_s_dadda_rca24_and_3_6_y0;
  assign f_s_dadda_rca24_ha8_f_s_dadda_rca24_and_2_7_y0 = f_s_dadda_rca24_and_2_7_y0;
  assign f_s_dadda_rca24_ha8_y0 = f_s_dadda_rca24_ha8_f_s_dadda_rca24_and_3_6_y0 ^ f_s_dadda_rca24_ha8_f_s_dadda_rca24_and_2_7_y0;
  assign f_s_dadda_rca24_ha8_y1 = f_s_dadda_rca24_ha8_f_s_dadda_rca24_and_3_6_y0 & f_s_dadda_rca24_ha8_f_s_dadda_rca24_and_2_7_y0;
  assign f_s_dadda_rca24_fa31_f_s_dadda_rca24_ha8_y1 = f_s_dadda_rca24_ha8_y1;
  assign f_s_dadda_rca24_fa31_f_s_dadda_rca24_fa30_y4 = f_s_dadda_rca24_fa30_y4;
  assign f_s_dadda_rca24_fa31_f_s_dadda_rca24_fa29_y4 = f_s_dadda_rca24_fa29_y4;
  assign f_s_dadda_rca24_fa31_y0 = f_s_dadda_rca24_fa31_f_s_dadda_rca24_ha8_y1 ^ f_s_dadda_rca24_fa31_f_s_dadda_rca24_fa30_y4;
  assign f_s_dadda_rca24_fa31_y1 = f_s_dadda_rca24_fa31_f_s_dadda_rca24_ha8_y1 & f_s_dadda_rca24_fa31_f_s_dadda_rca24_fa30_y4;
  assign f_s_dadda_rca24_fa31_y2 = f_s_dadda_rca24_fa31_y0 ^ f_s_dadda_rca24_fa31_f_s_dadda_rca24_fa29_y4;
  assign f_s_dadda_rca24_fa31_y3 = f_s_dadda_rca24_fa31_y0 & f_s_dadda_rca24_fa31_f_s_dadda_rca24_fa29_y4;
  assign f_s_dadda_rca24_fa31_y4 = f_s_dadda_rca24_fa31_y1 | f_s_dadda_rca24_fa31_y3;
  assign f_s_dadda_rca24_and_10_0_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_10_0_y0 = f_s_dadda_rca24_and_10_0_a_10 & f_s_dadda_rca24_and_10_0_b_0;
  assign f_s_dadda_rca24_and_9_1_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_9_1_y0 = f_s_dadda_rca24_and_9_1_a_9 & f_s_dadda_rca24_and_9_1_b_1;
  assign f_s_dadda_rca24_fa32_f_s_dadda_rca24_fa28_y4 = f_s_dadda_rca24_fa28_y4;
  assign f_s_dadda_rca24_fa32_f_s_dadda_rca24_and_10_0_y0 = f_s_dadda_rca24_and_10_0_y0;
  assign f_s_dadda_rca24_fa32_f_s_dadda_rca24_and_9_1_y0 = f_s_dadda_rca24_and_9_1_y0;
  assign f_s_dadda_rca24_fa32_y0 = f_s_dadda_rca24_fa32_f_s_dadda_rca24_fa28_y4 ^ f_s_dadda_rca24_fa32_f_s_dadda_rca24_and_10_0_y0;
  assign f_s_dadda_rca24_fa32_y1 = f_s_dadda_rca24_fa32_f_s_dadda_rca24_fa28_y4 & f_s_dadda_rca24_fa32_f_s_dadda_rca24_and_10_0_y0;
  assign f_s_dadda_rca24_fa32_y2 = f_s_dadda_rca24_fa32_y0 ^ f_s_dadda_rca24_fa32_f_s_dadda_rca24_and_9_1_y0;
  assign f_s_dadda_rca24_fa32_y3 = f_s_dadda_rca24_fa32_y0 & f_s_dadda_rca24_fa32_f_s_dadda_rca24_and_9_1_y0;
  assign f_s_dadda_rca24_fa32_y4 = f_s_dadda_rca24_fa32_y1 | f_s_dadda_rca24_fa32_y3;
  assign f_s_dadda_rca24_and_8_2_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_8_2_y0 = f_s_dadda_rca24_and_8_2_a_8 & f_s_dadda_rca24_and_8_2_b_2;
  assign f_s_dadda_rca24_and_7_3_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_7_3_y0 = f_s_dadda_rca24_and_7_3_a_7 & f_s_dadda_rca24_and_7_3_b_3;
  assign f_s_dadda_rca24_and_6_4_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_6_4_y0 = f_s_dadda_rca24_and_6_4_a_6 & f_s_dadda_rca24_and_6_4_b_4;
  assign f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_8_2_y0 = f_s_dadda_rca24_and_8_2_y0;
  assign f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_7_3_y0 = f_s_dadda_rca24_and_7_3_y0;
  assign f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_6_4_y0 = f_s_dadda_rca24_and_6_4_y0;
  assign f_s_dadda_rca24_fa33_y0 = f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_8_2_y0 ^ f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_7_3_y0;
  assign f_s_dadda_rca24_fa33_y1 = f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_8_2_y0 & f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_7_3_y0;
  assign f_s_dadda_rca24_fa33_y2 = f_s_dadda_rca24_fa33_y0 ^ f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_6_4_y0;
  assign f_s_dadda_rca24_fa33_y3 = f_s_dadda_rca24_fa33_y0 & f_s_dadda_rca24_fa33_f_s_dadda_rca24_and_6_4_y0;
  assign f_s_dadda_rca24_fa33_y4 = f_s_dadda_rca24_fa33_y1 | f_s_dadda_rca24_fa33_y3;
  assign f_s_dadda_rca24_and_5_5_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_5_5_y0 = f_s_dadda_rca24_and_5_5_a_5 & f_s_dadda_rca24_and_5_5_b_5;
  assign f_s_dadda_rca24_and_4_6_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_4_6_y0 = f_s_dadda_rca24_and_4_6_a_4 & f_s_dadda_rca24_and_4_6_b_6;
  assign f_s_dadda_rca24_and_3_7_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_3_7_y0 = f_s_dadda_rca24_and_3_7_a_3 & f_s_dadda_rca24_and_3_7_b_7;
  assign f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_5_5_y0 = f_s_dadda_rca24_and_5_5_y0;
  assign f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_4_6_y0 = f_s_dadda_rca24_and_4_6_y0;
  assign f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_3_7_y0 = f_s_dadda_rca24_and_3_7_y0;
  assign f_s_dadda_rca24_fa34_y0 = f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_5_5_y0 ^ f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_4_6_y0;
  assign f_s_dadda_rca24_fa34_y1 = f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_5_5_y0 & f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_4_6_y0;
  assign f_s_dadda_rca24_fa34_y2 = f_s_dadda_rca24_fa34_y0 ^ f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_3_7_y0;
  assign f_s_dadda_rca24_fa34_y3 = f_s_dadda_rca24_fa34_y0 & f_s_dadda_rca24_fa34_f_s_dadda_rca24_and_3_7_y0;
  assign f_s_dadda_rca24_fa34_y4 = f_s_dadda_rca24_fa34_y1 | f_s_dadda_rca24_fa34_y3;
  assign f_s_dadda_rca24_and_2_8_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_2_8_y0 = f_s_dadda_rca24_and_2_8_a_2 & f_s_dadda_rca24_and_2_8_b_8;
  assign f_s_dadda_rca24_and_1_9_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_1_9_y0 = f_s_dadda_rca24_and_1_9_a_1 & f_s_dadda_rca24_and_1_9_b_9;
  assign f_s_dadda_rca24_ha9_f_s_dadda_rca24_and_2_8_y0 = f_s_dadda_rca24_and_2_8_y0;
  assign f_s_dadda_rca24_ha9_f_s_dadda_rca24_and_1_9_y0 = f_s_dadda_rca24_and_1_9_y0;
  assign f_s_dadda_rca24_ha9_y0 = f_s_dadda_rca24_ha9_f_s_dadda_rca24_and_2_8_y0 ^ f_s_dadda_rca24_ha9_f_s_dadda_rca24_and_1_9_y0;
  assign f_s_dadda_rca24_ha9_y1 = f_s_dadda_rca24_ha9_f_s_dadda_rca24_and_2_8_y0 & f_s_dadda_rca24_ha9_f_s_dadda_rca24_and_1_9_y0;
  assign f_s_dadda_rca24_fa35_f_s_dadda_rca24_ha9_y1 = f_s_dadda_rca24_ha9_y1;
  assign f_s_dadda_rca24_fa35_f_s_dadda_rca24_fa34_y4 = f_s_dadda_rca24_fa34_y4;
  assign f_s_dadda_rca24_fa35_f_s_dadda_rca24_fa33_y4 = f_s_dadda_rca24_fa33_y4;
  assign f_s_dadda_rca24_fa35_y0 = f_s_dadda_rca24_fa35_f_s_dadda_rca24_ha9_y1 ^ f_s_dadda_rca24_fa35_f_s_dadda_rca24_fa34_y4;
  assign f_s_dadda_rca24_fa35_y1 = f_s_dadda_rca24_fa35_f_s_dadda_rca24_ha9_y1 & f_s_dadda_rca24_fa35_f_s_dadda_rca24_fa34_y4;
  assign f_s_dadda_rca24_fa35_y2 = f_s_dadda_rca24_fa35_y0 ^ f_s_dadda_rca24_fa35_f_s_dadda_rca24_fa33_y4;
  assign f_s_dadda_rca24_fa35_y3 = f_s_dadda_rca24_fa35_y0 & f_s_dadda_rca24_fa35_f_s_dadda_rca24_fa33_y4;
  assign f_s_dadda_rca24_fa35_y4 = f_s_dadda_rca24_fa35_y1 | f_s_dadda_rca24_fa35_y3;
  assign f_s_dadda_rca24_and_11_0_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_11_0_y0 = f_s_dadda_rca24_and_11_0_a_11 & f_s_dadda_rca24_and_11_0_b_0;
  assign f_s_dadda_rca24_fa36_f_s_dadda_rca24_fa32_y4 = f_s_dadda_rca24_fa32_y4;
  assign f_s_dadda_rca24_fa36_f_s_dadda_rca24_fa31_y4 = f_s_dadda_rca24_fa31_y4;
  assign f_s_dadda_rca24_fa36_f_s_dadda_rca24_and_11_0_y0 = f_s_dadda_rca24_and_11_0_y0;
  assign f_s_dadda_rca24_fa36_y0 = f_s_dadda_rca24_fa36_f_s_dadda_rca24_fa32_y4 ^ f_s_dadda_rca24_fa36_f_s_dadda_rca24_fa31_y4;
  assign f_s_dadda_rca24_fa36_y1 = f_s_dadda_rca24_fa36_f_s_dadda_rca24_fa32_y4 & f_s_dadda_rca24_fa36_f_s_dadda_rca24_fa31_y4;
  assign f_s_dadda_rca24_fa36_y2 = f_s_dadda_rca24_fa36_y0 ^ f_s_dadda_rca24_fa36_f_s_dadda_rca24_and_11_0_y0;
  assign f_s_dadda_rca24_fa36_y3 = f_s_dadda_rca24_fa36_y0 & f_s_dadda_rca24_fa36_f_s_dadda_rca24_and_11_0_y0;
  assign f_s_dadda_rca24_fa36_y4 = f_s_dadda_rca24_fa36_y1 | f_s_dadda_rca24_fa36_y3;
  assign f_s_dadda_rca24_and_10_1_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_10_1_y0 = f_s_dadda_rca24_and_10_1_a_10 & f_s_dadda_rca24_and_10_1_b_1;
  assign f_s_dadda_rca24_and_9_2_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_9_2_y0 = f_s_dadda_rca24_and_9_2_a_9 & f_s_dadda_rca24_and_9_2_b_2;
  assign f_s_dadda_rca24_and_8_3_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_8_3_y0 = f_s_dadda_rca24_and_8_3_a_8 & f_s_dadda_rca24_and_8_3_b_3;
  assign f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_10_1_y0 = f_s_dadda_rca24_and_10_1_y0;
  assign f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_9_2_y0 = f_s_dadda_rca24_and_9_2_y0;
  assign f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_8_3_y0 = f_s_dadda_rca24_and_8_3_y0;
  assign f_s_dadda_rca24_fa37_y0 = f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_10_1_y0 ^ f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_9_2_y0;
  assign f_s_dadda_rca24_fa37_y1 = f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_10_1_y0 & f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_9_2_y0;
  assign f_s_dadda_rca24_fa37_y2 = f_s_dadda_rca24_fa37_y0 ^ f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_8_3_y0;
  assign f_s_dadda_rca24_fa37_y3 = f_s_dadda_rca24_fa37_y0 & f_s_dadda_rca24_fa37_f_s_dadda_rca24_and_8_3_y0;
  assign f_s_dadda_rca24_fa37_y4 = f_s_dadda_rca24_fa37_y1 | f_s_dadda_rca24_fa37_y3;
  assign f_s_dadda_rca24_and_7_4_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_7_4_y0 = f_s_dadda_rca24_and_7_4_a_7 & f_s_dadda_rca24_and_7_4_b_4;
  assign f_s_dadda_rca24_and_6_5_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_6_5_y0 = f_s_dadda_rca24_and_6_5_a_6 & f_s_dadda_rca24_and_6_5_b_5;
  assign f_s_dadda_rca24_and_5_6_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_5_6_y0 = f_s_dadda_rca24_and_5_6_a_5 & f_s_dadda_rca24_and_5_6_b_6;
  assign f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_7_4_y0 = f_s_dadda_rca24_and_7_4_y0;
  assign f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_6_5_y0 = f_s_dadda_rca24_and_6_5_y0;
  assign f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_5_6_y0 = f_s_dadda_rca24_and_5_6_y0;
  assign f_s_dadda_rca24_fa38_y0 = f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_7_4_y0 ^ f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_6_5_y0;
  assign f_s_dadda_rca24_fa38_y1 = f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_7_4_y0 & f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_6_5_y0;
  assign f_s_dadda_rca24_fa38_y2 = f_s_dadda_rca24_fa38_y0 ^ f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_5_6_y0;
  assign f_s_dadda_rca24_fa38_y3 = f_s_dadda_rca24_fa38_y0 & f_s_dadda_rca24_fa38_f_s_dadda_rca24_and_5_6_y0;
  assign f_s_dadda_rca24_fa38_y4 = f_s_dadda_rca24_fa38_y1 | f_s_dadda_rca24_fa38_y3;
  assign f_s_dadda_rca24_and_4_7_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_4_7_y0 = f_s_dadda_rca24_and_4_7_a_4 & f_s_dadda_rca24_and_4_7_b_7;
  assign f_s_dadda_rca24_and_3_8_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_3_8_y0 = f_s_dadda_rca24_and_3_8_a_3 & f_s_dadda_rca24_and_3_8_b_8;
  assign f_s_dadda_rca24_and_2_9_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_2_9_y0 = f_s_dadda_rca24_and_2_9_a_2 & f_s_dadda_rca24_and_2_9_b_9;
  assign f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_4_7_y0 = f_s_dadda_rca24_and_4_7_y0;
  assign f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_3_8_y0 = f_s_dadda_rca24_and_3_8_y0;
  assign f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_2_9_y0 = f_s_dadda_rca24_and_2_9_y0;
  assign f_s_dadda_rca24_fa39_y0 = f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_4_7_y0 ^ f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_3_8_y0;
  assign f_s_dadda_rca24_fa39_y1 = f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_4_7_y0 & f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_3_8_y0;
  assign f_s_dadda_rca24_fa39_y2 = f_s_dadda_rca24_fa39_y0 ^ f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_2_9_y0;
  assign f_s_dadda_rca24_fa39_y3 = f_s_dadda_rca24_fa39_y0 & f_s_dadda_rca24_fa39_f_s_dadda_rca24_and_2_9_y0;
  assign f_s_dadda_rca24_fa39_y4 = f_s_dadda_rca24_fa39_y1 | f_s_dadda_rca24_fa39_y3;
  assign f_s_dadda_rca24_and_1_10_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_1_10_y0 = f_s_dadda_rca24_and_1_10_a_1 & f_s_dadda_rca24_and_1_10_b_10;
  assign f_s_dadda_rca24_and_0_11_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_0_11_y0 = f_s_dadda_rca24_and_0_11_a_0 & f_s_dadda_rca24_and_0_11_b_11;
  assign f_s_dadda_rca24_ha10_f_s_dadda_rca24_and_1_10_y0 = f_s_dadda_rca24_and_1_10_y0;
  assign f_s_dadda_rca24_ha10_f_s_dadda_rca24_and_0_11_y0 = f_s_dadda_rca24_and_0_11_y0;
  assign f_s_dadda_rca24_ha10_y0 = f_s_dadda_rca24_ha10_f_s_dadda_rca24_and_1_10_y0 ^ f_s_dadda_rca24_ha10_f_s_dadda_rca24_and_0_11_y0;
  assign f_s_dadda_rca24_ha10_y1 = f_s_dadda_rca24_ha10_f_s_dadda_rca24_and_1_10_y0 & f_s_dadda_rca24_ha10_f_s_dadda_rca24_and_0_11_y0;
  assign f_s_dadda_rca24_fa40_f_s_dadda_rca24_ha10_y1 = f_s_dadda_rca24_ha10_y1;
  assign f_s_dadda_rca24_fa40_f_s_dadda_rca24_fa39_y4 = f_s_dadda_rca24_fa39_y4;
  assign f_s_dadda_rca24_fa40_f_s_dadda_rca24_fa38_y4 = f_s_dadda_rca24_fa38_y4;
  assign f_s_dadda_rca24_fa40_y0 = f_s_dadda_rca24_fa40_f_s_dadda_rca24_ha10_y1 ^ f_s_dadda_rca24_fa40_f_s_dadda_rca24_fa39_y4;
  assign f_s_dadda_rca24_fa40_y1 = f_s_dadda_rca24_fa40_f_s_dadda_rca24_ha10_y1 & f_s_dadda_rca24_fa40_f_s_dadda_rca24_fa39_y4;
  assign f_s_dadda_rca24_fa40_y2 = f_s_dadda_rca24_fa40_y0 ^ f_s_dadda_rca24_fa40_f_s_dadda_rca24_fa38_y4;
  assign f_s_dadda_rca24_fa40_y3 = f_s_dadda_rca24_fa40_y0 & f_s_dadda_rca24_fa40_f_s_dadda_rca24_fa38_y4;
  assign f_s_dadda_rca24_fa40_y4 = f_s_dadda_rca24_fa40_y1 | f_s_dadda_rca24_fa40_y3;
  assign f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa37_y4 = f_s_dadda_rca24_fa37_y4;
  assign f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa36_y4 = f_s_dadda_rca24_fa36_y4;
  assign f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa35_y4 = f_s_dadda_rca24_fa35_y4;
  assign f_s_dadda_rca24_fa41_y0 = f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa37_y4 ^ f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa36_y4;
  assign f_s_dadda_rca24_fa41_y1 = f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa37_y4 & f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa36_y4;
  assign f_s_dadda_rca24_fa41_y2 = f_s_dadda_rca24_fa41_y0 ^ f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa35_y4;
  assign f_s_dadda_rca24_fa41_y3 = f_s_dadda_rca24_fa41_y0 & f_s_dadda_rca24_fa41_f_s_dadda_rca24_fa35_y4;
  assign f_s_dadda_rca24_fa41_y4 = f_s_dadda_rca24_fa41_y1 | f_s_dadda_rca24_fa41_y3;
  assign f_s_dadda_rca24_and_12_0_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_12_0_y0 = f_s_dadda_rca24_and_12_0_a_12 & f_s_dadda_rca24_and_12_0_b_0;
  assign f_s_dadda_rca24_and_11_1_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_11_1_y0 = f_s_dadda_rca24_and_11_1_a_11 & f_s_dadda_rca24_and_11_1_b_1;
  assign f_s_dadda_rca24_and_10_2_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_10_2_y0 = f_s_dadda_rca24_and_10_2_a_10 & f_s_dadda_rca24_and_10_2_b_2;
  assign f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_12_0_y0 = f_s_dadda_rca24_and_12_0_y0;
  assign f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_11_1_y0 = f_s_dadda_rca24_and_11_1_y0;
  assign f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_10_2_y0 = f_s_dadda_rca24_and_10_2_y0;
  assign f_s_dadda_rca24_fa42_y0 = f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_12_0_y0 ^ f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_11_1_y0;
  assign f_s_dadda_rca24_fa42_y1 = f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_12_0_y0 & f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_11_1_y0;
  assign f_s_dadda_rca24_fa42_y2 = f_s_dadda_rca24_fa42_y0 ^ f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_10_2_y0;
  assign f_s_dadda_rca24_fa42_y3 = f_s_dadda_rca24_fa42_y0 & f_s_dadda_rca24_fa42_f_s_dadda_rca24_and_10_2_y0;
  assign f_s_dadda_rca24_fa42_y4 = f_s_dadda_rca24_fa42_y1 | f_s_dadda_rca24_fa42_y3;
  assign f_s_dadda_rca24_and_9_3_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_9_3_y0 = f_s_dadda_rca24_and_9_3_a_9 & f_s_dadda_rca24_and_9_3_b_3;
  assign f_s_dadda_rca24_and_8_4_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_8_4_y0 = f_s_dadda_rca24_and_8_4_a_8 & f_s_dadda_rca24_and_8_4_b_4;
  assign f_s_dadda_rca24_and_7_5_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_7_5_y0 = f_s_dadda_rca24_and_7_5_a_7 & f_s_dadda_rca24_and_7_5_b_5;
  assign f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_9_3_y0 = f_s_dadda_rca24_and_9_3_y0;
  assign f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_8_4_y0 = f_s_dadda_rca24_and_8_4_y0;
  assign f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_7_5_y0 = f_s_dadda_rca24_and_7_5_y0;
  assign f_s_dadda_rca24_fa43_y0 = f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_9_3_y0 ^ f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_8_4_y0;
  assign f_s_dadda_rca24_fa43_y1 = f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_9_3_y0 & f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_8_4_y0;
  assign f_s_dadda_rca24_fa43_y2 = f_s_dadda_rca24_fa43_y0 ^ f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_7_5_y0;
  assign f_s_dadda_rca24_fa43_y3 = f_s_dadda_rca24_fa43_y0 & f_s_dadda_rca24_fa43_f_s_dadda_rca24_and_7_5_y0;
  assign f_s_dadda_rca24_fa43_y4 = f_s_dadda_rca24_fa43_y1 | f_s_dadda_rca24_fa43_y3;
  assign f_s_dadda_rca24_and_6_6_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_6_6_y0 = f_s_dadda_rca24_and_6_6_a_6 & f_s_dadda_rca24_and_6_6_b_6;
  assign f_s_dadda_rca24_and_5_7_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_5_7_y0 = f_s_dadda_rca24_and_5_7_a_5 & f_s_dadda_rca24_and_5_7_b_7;
  assign f_s_dadda_rca24_and_4_8_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_4_8_y0 = f_s_dadda_rca24_and_4_8_a_4 & f_s_dadda_rca24_and_4_8_b_8;
  assign f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_6_6_y0 = f_s_dadda_rca24_and_6_6_y0;
  assign f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_5_7_y0 = f_s_dadda_rca24_and_5_7_y0;
  assign f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_4_8_y0 = f_s_dadda_rca24_and_4_8_y0;
  assign f_s_dadda_rca24_fa44_y0 = f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_6_6_y0 ^ f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_5_7_y0;
  assign f_s_dadda_rca24_fa44_y1 = f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_6_6_y0 & f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_5_7_y0;
  assign f_s_dadda_rca24_fa44_y2 = f_s_dadda_rca24_fa44_y0 ^ f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_4_8_y0;
  assign f_s_dadda_rca24_fa44_y3 = f_s_dadda_rca24_fa44_y0 & f_s_dadda_rca24_fa44_f_s_dadda_rca24_and_4_8_y0;
  assign f_s_dadda_rca24_fa44_y4 = f_s_dadda_rca24_fa44_y1 | f_s_dadda_rca24_fa44_y3;
  assign f_s_dadda_rca24_and_3_9_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_3_9_y0 = f_s_dadda_rca24_and_3_9_a_3 & f_s_dadda_rca24_and_3_9_b_9;
  assign f_s_dadda_rca24_and_2_10_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_2_10_y0 = f_s_dadda_rca24_and_2_10_a_2 & f_s_dadda_rca24_and_2_10_b_10;
  assign f_s_dadda_rca24_and_1_11_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_1_11_y0 = f_s_dadda_rca24_and_1_11_a_1 & f_s_dadda_rca24_and_1_11_b_11;
  assign f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_3_9_y0 = f_s_dadda_rca24_and_3_9_y0;
  assign f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_2_10_y0 = f_s_dadda_rca24_and_2_10_y0;
  assign f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_1_11_y0 = f_s_dadda_rca24_and_1_11_y0;
  assign f_s_dadda_rca24_fa45_y0 = f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_3_9_y0 ^ f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_2_10_y0;
  assign f_s_dadda_rca24_fa45_y1 = f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_3_9_y0 & f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_2_10_y0;
  assign f_s_dadda_rca24_fa45_y2 = f_s_dadda_rca24_fa45_y0 ^ f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_1_11_y0;
  assign f_s_dadda_rca24_fa45_y3 = f_s_dadda_rca24_fa45_y0 & f_s_dadda_rca24_fa45_f_s_dadda_rca24_and_1_11_y0;
  assign f_s_dadda_rca24_fa45_y4 = f_s_dadda_rca24_fa45_y1 | f_s_dadda_rca24_fa45_y3;
  assign f_s_dadda_rca24_and_0_12_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_0_12_y0 = f_s_dadda_rca24_and_0_12_a_0 & f_s_dadda_rca24_and_0_12_b_12;
  assign f_s_dadda_rca24_ha11_f_s_dadda_rca24_and_0_12_y0 = f_s_dadda_rca24_and_0_12_y0;
  assign f_s_dadda_rca24_ha11_f_s_dadda_rca24_fa40_y2 = f_s_dadda_rca24_fa40_y2;
  assign f_s_dadda_rca24_ha11_y0 = f_s_dadda_rca24_ha11_f_s_dadda_rca24_and_0_12_y0 ^ f_s_dadda_rca24_ha11_f_s_dadda_rca24_fa40_y2;
  assign f_s_dadda_rca24_ha11_y1 = f_s_dadda_rca24_ha11_f_s_dadda_rca24_and_0_12_y0 & f_s_dadda_rca24_ha11_f_s_dadda_rca24_fa40_y2;
  assign f_s_dadda_rca24_fa46_f_s_dadda_rca24_ha11_y1 = f_s_dadda_rca24_ha11_y1;
  assign f_s_dadda_rca24_fa46_f_s_dadda_rca24_fa45_y4 = f_s_dadda_rca24_fa45_y4;
  assign f_s_dadda_rca24_fa46_f_s_dadda_rca24_fa44_y4 = f_s_dadda_rca24_fa44_y4;
  assign f_s_dadda_rca24_fa46_y0 = f_s_dadda_rca24_fa46_f_s_dadda_rca24_ha11_y1 ^ f_s_dadda_rca24_fa46_f_s_dadda_rca24_fa45_y4;
  assign f_s_dadda_rca24_fa46_y1 = f_s_dadda_rca24_fa46_f_s_dadda_rca24_ha11_y1 & f_s_dadda_rca24_fa46_f_s_dadda_rca24_fa45_y4;
  assign f_s_dadda_rca24_fa46_y2 = f_s_dadda_rca24_fa46_y0 ^ f_s_dadda_rca24_fa46_f_s_dadda_rca24_fa44_y4;
  assign f_s_dadda_rca24_fa46_y3 = f_s_dadda_rca24_fa46_y0 & f_s_dadda_rca24_fa46_f_s_dadda_rca24_fa44_y4;
  assign f_s_dadda_rca24_fa46_y4 = f_s_dadda_rca24_fa46_y1 | f_s_dadda_rca24_fa46_y3;
  assign f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa43_y4 = f_s_dadda_rca24_fa43_y4;
  assign f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa42_y4 = f_s_dadda_rca24_fa42_y4;
  assign f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa41_y4 = f_s_dadda_rca24_fa41_y4;
  assign f_s_dadda_rca24_fa47_y0 = f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa43_y4 ^ f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa42_y4;
  assign f_s_dadda_rca24_fa47_y1 = f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa43_y4 & f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa42_y4;
  assign f_s_dadda_rca24_fa47_y2 = f_s_dadda_rca24_fa47_y0 ^ f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa41_y4;
  assign f_s_dadda_rca24_fa47_y3 = f_s_dadda_rca24_fa47_y0 & f_s_dadda_rca24_fa47_f_s_dadda_rca24_fa41_y4;
  assign f_s_dadda_rca24_fa47_y4 = f_s_dadda_rca24_fa47_y1 | f_s_dadda_rca24_fa47_y3;
  assign f_s_dadda_rca24_and_13_0_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_13_0_y0 = f_s_dadda_rca24_and_13_0_a_13 & f_s_dadda_rca24_and_13_0_b_0;
  assign f_s_dadda_rca24_and_12_1_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_12_1_y0 = f_s_dadda_rca24_and_12_1_a_12 & f_s_dadda_rca24_and_12_1_b_1;
  assign f_s_dadda_rca24_fa48_f_s_dadda_rca24_fa40_y4 = f_s_dadda_rca24_fa40_y4;
  assign f_s_dadda_rca24_fa48_f_s_dadda_rca24_and_13_0_y0 = f_s_dadda_rca24_and_13_0_y0;
  assign f_s_dadda_rca24_fa48_f_s_dadda_rca24_and_12_1_y0 = f_s_dadda_rca24_and_12_1_y0;
  assign f_s_dadda_rca24_fa48_y0 = f_s_dadda_rca24_fa48_f_s_dadda_rca24_fa40_y4 ^ f_s_dadda_rca24_fa48_f_s_dadda_rca24_and_13_0_y0;
  assign f_s_dadda_rca24_fa48_y1 = f_s_dadda_rca24_fa48_f_s_dadda_rca24_fa40_y4 & f_s_dadda_rca24_fa48_f_s_dadda_rca24_and_13_0_y0;
  assign f_s_dadda_rca24_fa48_y2 = f_s_dadda_rca24_fa48_y0 ^ f_s_dadda_rca24_fa48_f_s_dadda_rca24_and_12_1_y0;
  assign f_s_dadda_rca24_fa48_y3 = f_s_dadda_rca24_fa48_y0 & f_s_dadda_rca24_fa48_f_s_dadda_rca24_and_12_1_y0;
  assign f_s_dadda_rca24_fa48_y4 = f_s_dadda_rca24_fa48_y1 | f_s_dadda_rca24_fa48_y3;
  assign f_s_dadda_rca24_and_11_2_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_11_2_y0 = f_s_dadda_rca24_and_11_2_a_11 & f_s_dadda_rca24_and_11_2_b_2;
  assign f_s_dadda_rca24_and_10_3_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_10_3_y0 = f_s_dadda_rca24_and_10_3_a_10 & f_s_dadda_rca24_and_10_3_b_3;
  assign f_s_dadda_rca24_and_9_4_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_9_4_y0 = f_s_dadda_rca24_and_9_4_a_9 & f_s_dadda_rca24_and_9_4_b_4;
  assign f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_11_2_y0 = f_s_dadda_rca24_and_11_2_y0;
  assign f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_10_3_y0 = f_s_dadda_rca24_and_10_3_y0;
  assign f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_9_4_y0 = f_s_dadda_rca24_and_9_4_y0;
  assign f_s_dadda_rca24_fa49_y0 = f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_11_2_y0 ^ f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_10_3_y0;
  assign f_s_dadda_rca24_fa49_y1 = f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_11_2_y0 & f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_10_3_y0;
  assign f_s_dadda_rca24_fa49_y2 = f_s_dadda_rca24_fa49_y0 ^ f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_9_4_y0;
  assign f_s_dadda_rca24_fa49_y3 = f_s_dadda_rca24_fa49_y0 & f_s_dadda_rca24_fa49_f_s_dadda_rca24_and_9_4_y0;
  assign f_s_dadda_rca24_fa49_y4 = f_s_dadda_rca24_fa49_y1 | f_s_dadda_rca24_fa49_y3;
  assign f_s_dadda_rca24_and_8_5_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_8_5_y0 = f_s_dadda_rca24_and_8_5_a_8 & f_s_dadda_rca24_and_8_5_b_5;
  assign f_s_dadda_rca24_and_7_6_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_7_6_y0 = f_s_dadda_rca24_and_7_6_a_7 & f_s_dadda_rca24_and_7_6_b_6;
  assign f_s_dadda_rca24_and_6_7_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_6_7_y0 = f_s_dadda_rca24_and_6_7_a_6 & f_s_dadda_rca24_and_6_7_b_7;
  assign f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_8_5_y0 = f_s_dadda_rca24_and_8_5_y0;
  assign f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_7_6_y0 = f_s_dadda_rca24_and_7_6_y0;
  assign f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_6_7_y0 = f_s_dadda_rca24_and_6_7_y0;
  assign f_s_dadda_rca24_fa50_y0 = f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_8_5_y0 ^ f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_7_6_y0;
  assign f_s_dadda_rca24_fa50_y1 = f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_8_5_y0 & f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_7_6_y0;
  assign f_s_dadda_rca24_fa50_y2 = f_s_dadda_rca24_fa50_y0 ^ f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_6_7_y0;
  assign f_s_dadda_rca24_fa50_y3 = f_s_dadda_rca24_fa50_y0 & f_s_dadda_rca24_fa50_f_s_dadda_rca24_and_6_7_y0;
  assign f_s_dadda_rca24_fa50_y4 = f_s_dadda_rca24_fa50_y1 | f_s_dadda_rca24_fa50_y3;
  assign f_s_dadda_rca24_and_5_8_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_5_8_y0 = f_s_dadda_rca24_and_5_8_a_5 & f_s_dadda_rca24_and_5_8_b_8;
  assign f_s_dadda_rca24_and_4_9_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_4_9_y0 = f_s_dadda_rca24_and_4_9_a_4 & f_s_dadda_rca24_and_4_9_b_9;
  assign f_s_dadda_rca24_and_3_10_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_3_10_y0 = f_s_dadda_rca24_and_3_10_a_3 & f_s_dadda_rca24_and_3_10_b_10;
  assign f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_5_8_y0 = f_s_dadda_rca24_and_5_8_y0;
  assign f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_4_9_y0 = f_s_dadda_rca24_and_4_9_y0;
  assign f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_3_10_y0 = f_s_dadda_rca24_and_3_10_y0;
  assign f_s_dadda_rca24_fa51_y0 = f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_5_8_y0 ^ f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_4_9_y0;
  assign f_s_dadda_rca24_fa51_y1 = f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_5_8_y0 & f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_4_9_y0;
  assign f_s_dadda_rca24_fa51_y2 = f_s_dadda_rca24_fa51_y0 ^ f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_3_10_y0;
  assign f_s_dadda_rca24_fa51_y3 = f_s_dadda_rca24_fa51_y0 & f_s_dadda_rca24_fa51_f_s_dadda_rca24_and_3_10_y0;
  assign f_s_dadda_rca24_fa51_y4 = f_s_dadda_rca24_fa51_y1 | f_s_dadda_rca24_fa51_y3;
  assign f_s_dadda_rca24_and_2_11_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_2_11_y0 = f_s_dadda_rca24_and_2_11_a_2 & f_s_dadda_rca24_and_2_11_b_11;
  assign f_s_dadda_rca24_and_1_12_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_1_12_y0 = f_s_dadda_rca24_and_1_12_a_1 & f_s_dadda_rca24_and_1_12_b_12;
  assign f_s_dadda_rca24_and_0_13_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_0_13_y0 = f_s_dadda_rca24_and_0_13_a_0 & f_s_dadda_rca24_and_0_13_b_13;
  assign f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_2_11_y0 = f_s_dadda_rca24_and_2_11_y0;
  assign f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_1_12_y0 = f_s_dadda_rca24_and_1_12_y0;
  assign f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_0_13_y0 = f_s_dadda_rca24_and_0_13_y0;
  assign f_s_dadda_rca24_fa52_y0 = f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_2_11_y0 ^ f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_1_12_y0;
  assign f_s_dadda_rca24_fa52_y1 = f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_2_11_y0 & f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_1_12_y0;
  assign f_s_dadda_rca24_fa52_y2 = f_s_dadda_rca24_fa52_y0 ^ f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_0_13_y0;
  assign f_s_dadda_rca24_fa52_y3 = f_s_dadda_rca24_fa52_y0 & f_s_dadda_rca24_fa52_f_s_dadda_rca24_and_0_13_y0;
  assign f_s_dadda_rca24_fa52_y4 = f_s_dadda_rca24_fa52_y1 | f_s_dadda_rca24_fa52_y3;
  assign f_s_dadda_rca24_ha12_f_s_dadda_rca24_fa46_y2 = f_s_dadda_rca24_fa46_y2;
  assign f_s_dadda_rca24_ha12_f_s_dadda_rca24_fa47_y2 = f_s_dadda_rca24_fa47_y2;
  assign f_s_dadda_rca24_ha12_y0 = f_s_dadda_rca24_ha12_f_s_dadda_rca24_fa46_y2 ^ f_s_dadda_rca24_ha12_f_s_dadda_rca24_fa47_y2;
  assign f_s_dadda_rca24_ha12_y1 = f_s_dadda_rca24_ha12_f_s_dadda_rca24_fa46_y2 & f_s_dadda_rca24_ha12_f_s_dadda_rca24_fa47_y2;
  assign f_s_dadda_rca24_fa53_f_s_dadda_rca24_ha12_y1 = f_s_dadda_rca24_ha12_y1;
  assign f_s_dadda_rca24_fa53_f_s_dadda_rca24_fa52_y4 = f_s_dadda_rca24_fa52_y4;
  assign f_s_dadda_rca24_fa53_f_s_dadda_rca24_fa51_y4 = f_s_dadda_rca24_fa51_y4;
  assign f_s_dadda_rca24_fa53_y0 = f_s_dadda_rca24_fa53_f_s_dadda_rca24_ha12_y1 ^ f_s_dadda_rca24_fa53_f_s_dadda_rca24_fa52_y4;
  assign f_s_dadda_rca24_fa53_y1 = f_s_dadda_rca24_fa53_f_s_dadda_rca24_ha12_y1 & f_s_dadda_rca24_fa53_f_s_dadda_rca24_fa52_y4;
  assign f_s_dadda_rca24_fa53_y2 = f_s_dadda_rca24_fa53_y0 ^ f_s_dadda_rca24_fa53_f_s_dadda_rca24_fa51_y4;
  assign f_s_dadda_rca24_fa53_y3 = f_s_dadda_rca24_fa53_y0 & f_s_dadda_rca24_fa53_f_s_dadda_rca24_fa51_y4;
  assign f_s_dadda_rca24_fa53_y4 = f_s_dadda_rca24_fa53_y1 | f_s_dadda_rca24_fa53_y3;
  assign f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa50_y4 = f_s_dadda_rca24_fa50_y4;
  assign f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa49_y4 = f_s_dadda_rca24_fa49_y4;
  assign f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa48_y4 = f_s_dadda_rca24_fa48_y4;
  assign f_s_dadda_rca24_fa54_y0 = f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa50_y4 ^ f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa49_y4;
  assign f_s_dadda_rca24_fa54_y1 = f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa50_y4 & f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa49_y4;
  assign f_s_dadda_rca24_fa54_y2 = f_s_dadda_rca24_fa54_y0 ^ f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa48_y4;
  assign f_s_dadda_rca24_fa54_y3 = f_s_dadda_rca24_fa54_y0 & f_s_dadda_rca24_fa54_f_s_dadda_rca24_fa48_y4;
  assign f_s_dadda_rca24_fa54_y4 = f_s_dadda_rca24_fa54_y1 | f_s_dadda_rca24_fa54_y3;
  assign f_s_dadda_rca24_and_14_0_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_14_0_y0 = f_s_dadda_rca24_and_14_0_a_14 & f_s_dadda_rca24_and_14_0_b_0;
  assign f_s_dadda_rca24_fa55_f_s_dadda_rca24_fa47_y4 = f_s_dadda_rca24_fa47_y4;
  assign f_s_dadda_rca24_fa55_f_s_dadda_rca24_fa46_y4 = f_s_dadda_rca24_fa46_y4;
  assign f_s_dadda_rca24_fa55_f_s_dadda_rca24_and_14_0_y0 = f_s_dadda_rca24_and_14_0_y0;
  assign f_s_dadda_rca24_fa55_y0 = f_s_dadda_rca24_fa55_f_s_dadda_rca24_fa47_y4 ^ f_s_dadda_rca24_fa55_f_s_dadda_rca24_fa46_y4;
  assign f_s_dadda_rca24_fa55_y1 = f_s_dadda_rca24_fa55_f_s_dadda_rca24_fa47_y4 & f_s_dadda_rca24_fa55_f_s_dadda_rca24_fa46_y4;
  assign f_s_dadda_rca24_fa55_y2 = f_s_dadda_rca24_fa55_y0 ^ f_s_dadda_rca24_fa55_f_s_dadda_rca24_and_14_0_y0;
  assign f_s_dadda_rca24_fa55_y3 = f_s_dadda_rca24_fa55_y0 & f_s_dadda_rca24_fa55_f_s_dadda_rca24_and_14_0_y0;
  assign f_s_dadda_rca24_fa55_y4 = f_s_dadda_rca24_fa55_y1 | f_s_dadda_rca24_fa55_y3;
  assign f_s_dadda_rca24_and_13_1_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_13_1_y0 = f_s_dadda_rca24_and_13_1_a_13 & f_s_dadda_rca24_and_13_1_b_1;
  assign f_s_dadda_rca24_and_12_2_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_12_2_y0 = f_s_dadda_rca24_and_12_2_a_12 & f_s_dadda_rca24_and_12_2_b_2;
  assign f_s_dadda_rca24_and_11_3_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_11_3_y0 = f_s_dadda_rca24_and_11_3_a_11 & f_s_dadda_rca24_and_11_3_b_3;
  assign f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_13_1_y0 = f_s_dadda_rca24_and_13_1_y0;
  assign f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_12_2_y0 = f_s_dadda_rca24_and_12_2_y0;
  assign f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_11_3_y0 = f_s_dadda_rca24_and_11_3_y0;
  assign f_s_dadda_rca24_fa56_y0 = f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_13_1_y0 ^ f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_12_2_y0;
  assign f_s_dadda_rca24_fa56_y1 = f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_13_1_y0 & f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_12_2_y0;
  assign f_s_dadda_rca24_fa56_y2 = f_s_dadda_rca24_fa56_y0 ^ f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_11_3_y0;
  assign f_s_dadda_rca24_fa56_y3 = f_s_dadda_rca24_fa56_y0 & f_s_dadda_rca24_fa56_f_s_dadda_rca24_and_11_3_y0;
  assign f_s_dadda_rca24_fa56_y4 = f_s_dadda_rca24_fa56_y1 | f_s_dadda_rca24_fa56_y3;
  assign f_s_dadda_rca24_and_10_4_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_10_4_y0 = f_s_dadda_rca24_and_10_4_a_10 & f_s_dadda_rca24_and_10_4_b_4;
  assign f_s_dadda_rca24_and_9_5_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_9_5_y0 = f_s_dadda_rca24_and_9_5_a_9 & f_s_dadda_rca24_and_9_5_b_5;
  assign f_s_dadda_rca24_and_8_6_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_8_6_y0 = f_s_dadda_rca24_and_8_6_a_8 & f_s_dadda_rca24_and_8_6_b_6;
  assign f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_10_4_y0 = f_s_dadda_rca24_and_10_4_y0;
  assign f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_9_5_y0 = f_s_dadda_rca24_and_9_5_y0;
  assign f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_8_6_y0 = f_s_dadda_rca24_and_8_6_y0;
  assign f_s_dadda_rca24_fa57_y0 = f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_10_4_y0 ^ f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_9_5_y0;
  assign f_s_dadda_rca24_fa57_y1 = f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_10_4_y0 & f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_9_5_y0;
  assign f_s_dadda_rca24_fa57_y2 = f_s_dadda_rca24_fa57_y0 ^ f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_8_6_y0;
  assign f_s_dadda_rca24_fa57_y3 = f_s_dadda_rca24_fa57_y0 & f_s_dadda_rca24_fa57_f_s_dadda_rca24_and_8_6_y0;
  assign f_s_dadda_rca24_fa57_y4 = f_s_dadda_rca24_fa57_y1 | f_s_dadda_rca24_fa57_y3;
  assign f_s_dadda_rca24_and_7_7_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_7_7_y0 = f_s_dadda_rca24_and_7_7_a_7 & f_s_dadda_rca24_and_7_7_b_7;
  assign f_s_dadda_rca24_and_6_8_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_6_8_y0 = f_s_dadda_rca24_and_6_8_a_6 & f_s_dadda_rca24_and_6_8_b_8;
  assign f_s_dadda_rca24_and_5_9_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_5_9_y0 = f_s_dadda_rca24_and_5_9_a_5 & f_s_dadda_rca24_and_5_9_b_9;
  assign f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_7_7_y0 = f_s_dadda_rca24_and_7_7_y0;
  assign f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_6_8_y0 = f_s_dadda_rca24_and_6_8_y0;
  assign f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_5_9_y0 = f_s_dadda_rca24_and_5_9_y0;
  assign f_s_dadda_rca24_fa58_y0 = f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_7_7_y0 ^ f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_6_8_y0;
  assign f_s_dadda_rca24_fa58_y1 = f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_7_7_y0 & f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_6_8_y0;
  assign f_s_dadda_rca24_fa58_y2 = f_s_dadda_rca24_fa58_y0 ^ f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_5_9_y0;
  assign f_s_dadda_rca24_fa58_y3 = f_s_dadda_rca24_fa58_y0 & f_s_dadda_rca24_fa58_f_s_dadda_rca24_and_5_9_y0;
  assign f_s_dadda_rca24_fa58_y4 = f_s_dadda_rca24_fa58_y1 | f_s_dadda_rca24_fa58_y3;
  assign f_s_dadda_rca24_and_4_10_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_4_10_y0 = f_s_dadda_rca24_and_4_10_a_4 & f_s_dadda_rca24_and_4_10_b_10;
  assign f_s_dadda_rca24_and_3_11_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_3_11_y0 = f_s_dadda_rca24_and_3_11_a_3 & f_s_dadda_rca24_and_3_11_b_11;
  assign f_s_dadda_rca24_and_2_12_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_2_12_y0 = f_s_dadda_rca24_and_2_12_a_2 & f_s_dadda_rca24_and_2_12_b_12;
  assign f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_4_10_y0 = f_s_dadda_rca24_and_4_10_y0;
  assign f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_3_11_y0 = f_s_dadda_rca24_and_3_11_y0;
  assign f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_2_12_y0 = f_s_dadda_rca24_and_2_12_y0;
  assign f_s_dadda_rca24_fa59_y0 = f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_4_10_y0 ^ f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_3_11_y0;
  assign f_s_dadda_rca24_fa59_y1 = f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_4_10_y0 & f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_3_11_y0;
  assign f_s_dadda_rca24_fa59_y2 = f_s_dadda_rca24_fa59_y0 ^ f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_2_12_y0;
  assign f_s_dadda_rca24_fa59_y3 = f_s_dadda_rca24_fa59_y0 & f_s_dadda_rca24_fa59_f_s_dadda_rca24_and_2_12_y0;
  assign f_s_dadda_rca24_fa59_y4 = f_s_dadda_rca24_fa59_y1 | f_s_dadda_rca24_fa59_y3;
  assign f_s_dadda_rca24_and_1_13_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_1_13_y0 = f_s_dadda_rca24_and_1_13_a_1 & f_s_dadda_rca24_and_1_13_b_13;
  assign f_s_dadda_rca24_and_0_14_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_0_14_y0 = f_s_dadda_rca24_and_0_14_a_0 & f_s_dadda_rca24_and_0_14_b_14;
  assign f_s_dadda_rca24_fa60_f_s_dadda_rca24_and_1_13_y0 = f_s_dadda_rca24_and_1_13_y0;
  assign f_s_dadda_rca24_fa60_f_s_dadda_rca24_and_0_14_y0 = f_s_dadda_rca24_and_0_14_y0;
  assign f_s_dadda_rca24_fa60_f_s_dadda_rca24_fa53_y2 = f_s_dadda_rca24_fa53_y2;
  assign f_s_dadda_rca24_fa60_y0 = f_s_dadda_rca24_fa60_f_s_dadda_rca24_and_1_13_y0 ^ f_s_dadda_rca24_fa60_f_s_dadda_rca24_and_0_14_y0;
  assign f_s_dadda_rca24_fa60_y1 = f_s_dadda_rca24_fa60_f_s_dadda_rca24_and_1_13_y0 & f_s_dadda_rca24_fa60_f_s_dadda_rca24_and_0_14_y0;
  assign f_s_dadda_rca24_fa60_y2 = f_s_dadda_rca24_fa60_y0 ^ f_s_dadda_rca24_fa60_f_s_dadda_rca24_fa53_y2;
  assign f_s_dadda_rca24_fa60_y3 = f_s_dadda_rca24_fa60_y0 & f_s_dadda_rca24_fa60_f_s_dadda_rca24_fa53_y2;
  assign f_s_dadda_rca24_fa60_y4 = f_s_dadda_rca24_fa60_y1 | f_s_dadda_rca24_fa60_y3;
  assign f_s_dadda_rca24_ha13_f_s_dadda_rca24_fa54_y2 = f_s_dadda_rca24_fa54_y2;
  assign f_s_dadda_rca24_ha13_f_s_dadda_rca24_fa55_y2 = f_s_dadda_rca24_fa55_y2;
  assign f_s_dadda_rca24_ha13_y0 = f_s_dadda_rca24_ha13_f_s_dadda_rca24_fa54_y2 ^ f_s_dadda_rca24_ha13_f_s_dadda_rca24_fa55_y2;
  assign f_s_dadda_rca24_ha13_y1 = f_s_dadda_rca24_ha13_f_s_dadda_rca24_fa54_y2 & f_s_dadda_rca24_ha13_f_s_dadda_rca24_fa55_y2;
  assign f_s_dadda_rca24_fa61_f_s_dadda_rca24_ha13_y1 = f_s_dadda_rca24_ha13_y1;
  assign f_s_dadda_rca24_fa61_f_s_dadda_rca24_fa60_y4 = f_s_dadda_rca24_fa60_y4;
  assign f_s_dadda_rca24_fa61_f_s_dadda_rca24_fa59_y4 = f_s_dadda_rca24_fa59_y4;
  assign f_s_dadda_rca24_fa61_y0 = f_s_dadda_rca24_fa61_f_s_dadda_rca24_ha13_y1 ^ f_s_dadda_rca24_fa61_f_s_dadda_rca24_fa60_y4;
  assign f_s_dadda_rca24_fa61_y1 = f_s_dadda_rca24_fa61_f_s_dadda_rca24_ha13_y1 & f_s_dadda_rca24_fa61_f_s_dadda_rca24_fa60_y4;
  assign f_s_dadda_rca24_fa61_y2 = f_s_dadda_rca24_fa61_y0 ^ f_s_dadda_rca24_fa61_f_s_dadda_rca24_fa59_y4;
  assign f_s_dadda_rca24_fa61_y3 = f_s_dadda_rca24_fa61_y0 & f_s_dadda_rca24_fa61_f_s_dadda_rca24_fa59_y4;
  assign f_s_dadda_rca24_fa61_y4 = f_s_dadda_rca24_fa61_y1 | f_s_dadda_rca24_fa61_y3;
  assign f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa58_y4 = f_s_dadda_rca24_fa58_y4;
  assign f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa57_y4 = f_s_dadda_rca24_fa57_y4;
  assign f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa56_y4 = f_s_dadda_rca24_fa56_y4;
  assign f_s_dadda_rca24_fa62_y0 = f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa58_y4 ^ f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa57_y4;
  assign f_s_dadda_rca24_fa62_y1 = f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa58_y4 & f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa57_y4;
  assign f_s_dadda_rca24_fa62_y2 = f_s_dadda_rca24_fa62_y0 ^ f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa56_y4;
  assign f_s_dadda_rca24_fa62_y3 = f_s_dadda_rca24_fa62_y0 & f_s_dadda_rca24_fa62_f_s_dadda_rca24_fa56_y4;
  assign f_s_dadda_rca24_fa62_y4 = f_s_dadda_rca24_fa62_y1 | f_s_dadda_rca24_fa62_y3;
  assign f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa55_y4 = f_s_dadda_rca24_fa55_y4;
  assign f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa54_y4 = f_s_dadda_rca24_fa54_y4;
  assign f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa53_y4 = f_s_dadda_rca24_fa53_y4;
  assign f_s_dadda_rca24_fa63_y0 = f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa55_y4 ^ f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa54_y4;
  assign f_s_dadda_rca24_fa63_y1 = f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa55_y4 & f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa54_y4;
  assign f_s_dadda_rca24_fa63_y2 = f_s_dadda_rca24_fa63_y0 ^ f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa53_y4;
  assign f_s_dadda_rca24_fa63_y3 = f_s_dadda_rca24_fa63_y0 & f_s_dadda_rca24_fa63_f_s_dadda_rca24_fa53_y4;
  assign f_s_dadda_rca24_fa63_y4 = f_s_dadda_rca24_fa63_y1 | f_s_dadda_rca24_fa63_y3;
  assign f_s_dadda_rca24_and_15_0_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_15_0_y0 = f_s_dadda_rca24_and_15_0_a_15 & f_s_dadda_rca24_and_15_0_b_0;
  assign f_s_dadda_rca24_and_14_1_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_14_1_y0 = f_s_dadda_rca24_and_14_1_a_14 & f_s_dadda_rca24_and_14_1_b_1;
  assign f_s_dadda_rca24_and_13_2_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_13_2_y0 = f_s_dadda_rca24_and_13_2_a_13 & f_s_dadda_rca24_and_13_2_b_2;
  assign f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_15_0_y0 = f_s_dadda_rca24_and_15_0_y0;
  assign f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_14_1_y0 = f_s_dadda_rca24_and_14_1_y0;
  assign f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_13_2_y0 = f_s_dadda_rca24_and_13_2_y0;
  assign f_s_dadda_rca24_fa64_y0 = f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_15_0_y0 ^ f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_14_1_y0;
  assign f_s_dadda_rca24_fa64_y1 = f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_15_0_y0 & f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_14_1_y0;
  assign f_s_dadda_rca24_fa64_y2 = f_s_dadda_rca24_fa64_y0 ^ f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_13_2_y0;
  assign f_s_dadda_rca24_fa64_y3 = f_s_dadda_rca24_fa64_y0 & f_s_dadda_rca24_fa64_f_s_dadda_rca24_and_13_2_y0;
  assign f_s_dadda_rca24_fa64_y4 = f_s_dadda_rca24_fa64_y1 | f_s_dadda_rca24_fa64_y3;
  assign f_s_dadda_rca24_and_12_3_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_12_3_y0 = f_s_dadda_rca24_and_12_3_a_12 & f_s_dadda_rca24_and_12_3_b_3;
  assign f_s_dadda_rca24_and_11_4_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_11_4_y0 = f_s_dadda_rca24_and_11_4_a_11 & f_s_dadda_rca24_and_11_4_b_4;
  assign f_s_dadda_rca24_and_10_5_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_10_5_y0 = f_s_dadda_rca24_and_10_5_a_10 & f_s_dadda_rca24_and_10_5_b_5;
  assign f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_12_3_y0 = f_s_dadda_rca24_and_12_3_y0;
  assign f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_11_4_y0 = f_s_dadda_rca24_and_11_4_y0;
  assign f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_10_5_y0 = f_s_dadda_rca24_and_10_5_y0;
  assign f_s_dadda_rca24_fa65_y0 = f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_12_3_y0 ^ f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_11_4_y0;
  assign f_s_dadda_rca24_fa65_y1 = f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_12_3_y0 & f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_11_4_y0;
  assign f_s_dadda_rca24_fa65_y2 = f_s_dadda_rca24_fa65_y0 ^ f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_10_5_y0;
  assign f_s_dadda_rca24_fa65_y3 = f_s_dadda_rca24_fa65_y0 & f_s_dadda_rca24_fa65_f_s_dadda_rca24_and_10_5_y0;
  assign f_s_dadda_rca24_fa65_y4 = f_s_dadda_rca24_fa65_y1 | f_s_dadda_rca24_fa65_y3;
  assign f_s_dadda_rca24_and_9_6_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_9_6_y0 = f_s_dadda_rca24_and_9_6_a_9 & f_s_dadda_rca24_and_9_6_b_6;
  assign f_s_dadda_rca24_and_8_7_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_8_7_y0 = f_s_dadda_rca24_and_8_7_a_8 & f_s_dadda_rca24_and_8_7_b_7;
  assign f_s_dadda_rca24_and_7_8_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_7_8_y0 = f_s_dadda_rca24_and_7_8_a_7 & f_s_dadda_rca24_and_7_8_b_8;
  assign f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_9_6_y0 = f_s_dadda_rca24_and_9_6_y0;
  assign f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_8_7_y0 = f_s_dadda_rca24_and_8_7_y0;
  assign f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_7_8_y0 = f_s_dadda_rca24_and_7_8_y0;
  assign f_s_dadda_rca24_fa66_y0 = f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_9_6_y0 ^ f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_8_7_y0;
  assign f_s_dadda_rca24_fa66_y1 = f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_9_6_y0 & f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_8_7_y0;
  assign f_s_dadda_rca24_fa66_y2 = f_s_dadda_rca24_fa66_y0 ^ f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_7_8_y0;
  assign f_s_dadda_rca24_fa66_y3 = f_s_dadda_rca24_fa66_y0 & f_s_dadda_rca24_fa66_f_s_dadda_rca24_and_7_8_y0;
  assign f_s_dadda_rca24_fa66_y4 = f_s_dadda_rca24_fa66_y1 | f_s_dadda_rca24_fa66_y3;
  assign f_s_dadda_rca24_and_6_9_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_6_9_y0 = f_s_dadda_rca24_and_6_9_a_6 & f_s_dadda_rca24_and_6_9_b_9;
  assign f_s_dadda_rca24_and_5_10_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_5_10_y0 = f_s_dadda_rca24_and_5_10_a_5 & f_s_dadda_rca24_and_5_10_b_10;
  assign f_s_dadda_rca24_and_4_11_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_4_11_y0 = f_s_dadda_rca24_and_4_11_a_4 & f_s_dadda_rca24_and_4_11_b_11;
  assign f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_6_9_y0 = f_s_dadda_rca24_and_6_9_y0;
  assign f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_5_10_y0 = f_s_dadda_rca24_and_5_10_y0;
  assign f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_4_11_y0 = f_s_dadda_rca24_and_4_11_y0;
  assign f_s_dadda_rca24_fa67_y0 = f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_6_9_y0 ^ f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_5_10_y0;
  assign f_s_dadda_rca24_fa67_y1 = f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_6_9_y0 & f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_5_10_y0;
  assign f_s_dadda_rca24_fa67_y2 = f_s_dadda_rca24_fa67_y0 ^ f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_4_11_y0;
  assign f_s_dadda_rca24_fa67_y3 = f_s_dadda_rca24_fa67_y0 & f_s_dadda_rca24_fa67_f_s_dadda_rca24_and_4_11_y0;
  assign f_s_dadda_rca24_fa67_y4 = f_s_dadda_rca24_fa67_y1 | f_s_dadda_rca24_fa67_y3;
  assign f_s_dadda_rca24_and_3_12_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_3_12_y0 = f_s_dadda_rca24_and_3_12_a_3 & f_s_dadda_rca24_and_3_12_b_12;
  assign f_s_dadda_rca24_and_2_13_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_2_13_y0 = f_s_dadda_rca24_and_2_13_a_2 & f_s_dadda_rca24_and_2_13_b_13;
  assign f_s_dadda_rca24_and_1_14_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_1_14_y0 = f_s_dadda_rca24_and_1_14_a_1 & f_s_dadda_rca24_and_1_14_b_14;
  assign f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_3_12_y0 = f_s_dadda_rca24_and_3_12_y0;
  assign f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_2_13_y0 = f_s_dadda_rca24_and_2_13_y0;
  assign f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_1_14_y0 = f_s_dadda_rca24_and_1_14_y0;
  assign f_s_dadda_rca24_fa68_y0 = f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_3_12_y0 ^ f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_2_13_y0;
  assign f_s_dadda_rca24_fa68_y1 = f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_3_12_y0 & f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_2_13_y0;
  assign f_s_dadda_rca24_fa68_y2 = f_s_dadda_rca24_fa68_y0 ^ f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_1_14_y0;
  assign f_s_dadda_rca24_fa68_y3 = f_s_dadda_rca24_fa68_y0 & f_s_dadda_rca24_fa68_f_s_dadda_rca24_and_1_14_y0;
  assign f_s_dadda_rca24_fa68_y4 = f_s_dadda_rca24_fa68_y1 | f_s_dadda_rca24_fa68_y3;
  assign f_s_dadda_rca24_and_0_15_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_0_15_y0 = f_s_dadda_rca24_and_0_15_a_0 & f_s_dadda_rca24_and_0_15_b_15;
  assign f_s_dadda_rca24_fa69_f_s_dadda_rca24_and_0_15_y0 = f_s_dadda_rca24_and_0_15_y0;
  assign f_s_dadda_rca24_fa69_f_s_dadda_rca24_fa61_y2 = f_s_dadda_rca24_fa61_y2;
  assign f_s_dadda_rca24_fa69_f_s_dadda_rca24_fa62_y2 = f_s_dadda_rca24_fa62_y2;
  assign f_s_dadda_rca24_fa69_y0 = f_s_dadda_rca24_fa69_f_s_dadda_rca24_and_0_15_y0 ^ f_s_dadda_rca24_fa69_f_s_dadda_rca24_fa61_y2;
  assign f_s_dadda_rca24_fa69_y1 = f_s_dadda_rca24_fa69_f_s_dadda_rca24_and_0_15_y0 & f_s_dadda_rca24_fa69_f_s_dadda_rca24_fa61_y2;
  assign f_s_dadda_rca24_fa69_y2 = f_s_dadda_rca24_fa69_y0 ^ f_s_dadda_rca24_fa69_f_s_dadda_rca24_fa62_y2;
  assign f_s_dadda_rca24_fa69_y3 = f_s_dadda_rca24_fa69_y0 & f_s_dadda_rca24_fa69_f_s_dadda_rca24_fa62_y2;
  assign f_s_dadda_rca24_fa69_y4 = f_s_dadda_rca24_fa69_y1 | f_s_dadda_rca24_fa69_y3;
  assign f_s_dadda_rca24_ha14_f_s_dadda_rca24_fa63_y2 = f_s_dadda_rca24_fa63_y2;
  assign f_s_dadda_rca24_ha14_f_s_dadda_rca24_fa64_y2 = f_s_dadda_rca24_fa64_y2;
  assign f_s_dadda_rca24_ha14_y0 = f_s_dadda_rca24_ha14_f_s_dadda_rca24_fa63_y2 ^ f_s_dadda_rca24_ha14_f_s_dadda_rca24_fa64_y2;
  assign f_s_dadda_rca24_ha14_y1 = f_s_dadda_rca24_ha14_f_s_dadda_rca24_fa63_y2 & f_s_dadda_rca24_ha14_f_s_dadda_rca24_fa64_y2;
  assign f_s_dadda_rca24_fa70_f_s_dadda_rca24_ha14_y1 = f_s_dadda_rca24_ha14_y1;
  assign f_s_dadda_rca24_fa70_f_s_dadda_rca24_fa69_y4 = f_s_dadda_rca24_fa69_y4;
  assign f_s_dadda_rca24_fa70_f_s_dadda_rca24_fa68_y4 = f_s_dadda_rca24_fa68_y4;
  assign f_s_dadda_rca24_fa70_y0 = f_s_dadda_rca24_fa70_f_s_dadda_rca24_ha14_y1 ^ f_s_dadda_rca24_fa70_f_s_dadda_rca24_fa69_y4;
  assign f_s_dadda_rca24_fa70_y1 = f_s_dadda_rca24_fa70_f_s_dadda_rca24_ha14_y1 & f_s_dadda_rca24_fa70_f_s_dadda_rca24_fa69_y4;
  assign f_s_dadda_rca24_fa70_y2 = f_s_dadda_rca24_fa70_y0 ^ f_s_dadda_rca24_fa70_f_s_dadda_rca24_fa68_y4;
  assign f_s_dadda_rca24_fa70_y3 = f_s_dadda_rca24_fa70_y0 & f_s_dadda_rca24_fa70_f_s_dadda_rca24_fa68_y4;
  assign f_s_dadda_rca24_fa70_y4 = f_s_dadda_rca24_fa70_y1 | f_s_dadda_rca24_fa70_y3;
  assign f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa67_y4 = f_s_dadda_rca24_fa67_y4;
  assign f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa66_y4 = f_s_dadda_rca24_fa66_y4;
  assign f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa65_y4 = f_s_dadda_rca24_fa65_y4;
  assign f_s_dadda_rca24_fa71_y0 = f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa67_y4 ^ f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa66_y4;
  assign f_s_dadda_rca24_fa71_y1 = f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa67_y4 & f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa66_y4;
  assign f_s_dadda_rca24_fa71_y2 = f_s_dadda_rca24_fa71_y0 ^ f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa65_y4;
  assign f_s_dadda_rca24_fa71_y3 = f_s_dadda_rca24_fa71_y0 & f_s_dadda_rca24_fa71_f_s_dadda_rca24_fa65_y4;
  assign f_s_dadda_rca24_fa71_y4 = f_s_dadda_rca24_fa71_y1 | f_s_dadda_rca24_fa71_y3;
  assign f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa64_y4 = f_s_dadda_rca24_fa64_y4;
  assign f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa63_y4 = f_s_dadda_rca24_fa63_y4;
  assign f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa62_y4 = f_s_dadda_rca24_fa62_y4;
  assign f_s_dadda_rca24_fa72_y0 = f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa64_y4 ^ f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa63_y4;
  assign f_s_dadda_rca24_fa72_y1 = f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa64_y4 & f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa63_y4;
  assign f_s_dadda_rca24_fa72_y2 = f_s_dadda_rca24_fa72_y0 ^ f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa62_y4;
  assign f_s_dadda_rca24_fa72_y3 = f_s_dadda_rca24_fa72_y0 & f_s_dadda_rca24_fa72_f_s_dadda_rca24_fa62_y4;
  assign f_s_dadda_rca24_fa72_y4 = f_s_dadda_rca24_fa72_y1 | f_s_dadda_rca24_fa72_y3;
  assign f_s_dadda_rca24_and_16_0_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_16_0_y0 = f_s_dadda_rca24_and_16_0_a_16 & f_s_dadda_rca24_and_16_0_b_0;
  assign f_s_dadda_rca24_and_15_1_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_15_1_y0 = f_s_dadda_rca24_and_15_1_a_15 & f_s_dadda_rca24_and_15_1_b_1;
  assign f_s_dadda_rca24_fa73_f_s_dadda_rca24_fa61_y4 = f_s_dadda_rca24_fa61_y4;
  assign f_s_dadda_rca24_fa73_f_s_dadda_rca24_and_16_0_y0 = f_s_dadda_rca24_and_16_0_y0;
  assign f_s_dadda_rca24_fa73_f_s_dadda_rca24_and_15_1_y0 = f_s_dadda_rca24_and_15_1_y0;
  assign f_s_dadda_rca24_fa73_y0 = f_s_dadda_rca24_fa73_f_s_dadda_rca24_fa61_y4 ^ f_s_dadda_rca24_fa73_f_s_dadda_rca24_and_16_0_y0;
  assign f_s_dadda_rca24_fa73_y1 = f_s_dadda_rca24_fa73_f_s_dadda_rca24_fa61_y4 & f_s_dadda_rca24_fa73_f_s_dadda_rca24_and_16_0_y0;
  assign f_s_dadda_rca24_fa73_y2 = f_s_dadda_rca24_fa73_y0 ^ f_s_dadda_rca24_fa73_f_s_dadda_rca24_and_15_1_y0;
  assign f_s_dadda_rca24_fa73_y3 = f_s_dadda_rca24_fa73_y0 & f_s_dadda_rca24_fa73_f_s_dadda_rca24_and_15_1_y0;
  assign f_s_dadda_rca24_fa73_y4 = f_s_dadda_rca24_fa73_y1 | f_s_dadda_rca24_fa73_y3;
  assign f_s_dadda_rca24_and_14_2_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_14_2_y0 = f_s_dadda_rca24_and_14_2_a_14 & f_s_dadda_rca24_and_14_2_b_2;
  assign f_s_dadda_rca24_and_13_3_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_13_3_y0 = f_s_dadda_rca24_and_13_3_a_13 & f_s_dadda_rca24_and_13_3_b_3;
  assign f_s_dadda_rca24_and_12_4_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_12_4_y0 = f_s_dadda_rca24_and_12_4_a_12 & f_s_dadda_rca24_and_12_4_b_4;
  assign f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_14_2_y0 = f_s_dadda_rca24_and_14_2_y0;
  assign f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_13_3_y0 = f_s_dadda_rca24_and_13_3_y0;
  assign f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_12_4_y0 = f_s_dadda_rca24_and_12_4_y0;
  assign f_s_dadda_rca24_fa74_y0 = f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_14_2_y0 ^ f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_13_3_y0;
  assign f_s_dadda_rca24_fa74_y1 = f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_14_2_y0 & f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_13_3_y0;
  assign f_s_dadda_rca24_fa74_y2 = f_s_dadda_rca24_fa74_y0 ^ f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_12_4_y0;
  assign f_s_dadda_rca24_fa74_y3 = f_s_dadda_rca24_fa74_y0 & f_s_dadda_rca24_fa74_f_s_dadda_rca24_and_12_4_y0;
  assign f_s_dadda_rca24_fa74_y4 = f_s_dadda_rca24_fa74_y1 | f_s_dadda_rca24_fa74_y3;
  assign f_s_dadda_rca24_and_11_5_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_11_5_y0 = f_s_dadda_rca24_and_11_5_a_11 & f_s_dadda_rca24_and_11_5_b_5;
  assign f_s_dadda_rca24_and_10_6_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_10_6_y0 = f_s_dadda_rca24_and_10_6_a_10 & f_s_dadda_rca24_and_10_6_b_6;
  assign f_s_dadda_rca24_and_9_7_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_9_7_y0 = f_s_dadda_rca24_and_9_7_a_9 & f_s_dadda_rca24_and_9_7_b_7;
  assign f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_11_5_y0 = f_s_dadda_rca24_and_11_5_y0;
  assign f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_10_6_y0 = f_s_dadda_rca24_and_10_6_y0;
  assign f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_9_7_y0 = f_s_dadda_rca24_and_9_7_y0;
  assign f_s_dadda_rca24_fa75_y0 = f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_11_5_y0 ^ f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_10_6_y0;
  assign f_s_dadda_rca24_fa75_y1 = f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_11_5_y0 & f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_10_6_y0;
  assign f_s_dadda_rca24_fa75_y2 = f_s_dadda_rca24_fa75_y0 ^ f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_9_7_y0;
  assign f_s_dadda_rca24_fa75_y3 = f_s_dadda_rca24_fa75_y0 & f_s_dadda_rca24_fa75_f_s_dadda_rca24_and_9_7_y0;
  assign f_s_dadda_rca24_fa75_y4 = f_s_dadda_rca24_fa75_y1 | f_s_dadda_rca24_fa75_y3;
  assign f_s_dadda_rca24_and_8_8_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_8_8_y0 = f_s_dadda_rca24_and_8_8_a_8 & f_s_dadda_rca24_and_8_8_b_8;
  assign f_s_dadda_rca24_and_7_9_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_7_9_y0 = f_s_dadda_rca24_and_7_9_a_7 & f_s_dadda_rca24_and_7_9_b_9;
  assign f_s_dadda_rca24_and_6_10_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_6_10_y0 = f_s_dadda_rca24_and_6_10_a_6 & f_s_dadda_rca24_and_6_10_b_10;
  assign f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_8_8_y0 = f_s_dadda_rca24_and_8_8_y0;
  assign f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_7_9_y0 = f_s_dadda_rca24_and_7_9_y0;
  assign f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_6_10_y0 = f_s_dadda_rca24_and_6_10_y0;
  assign f_s_dadda_rca24_fa76_y0 = f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_8_8_y0 ^ f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_7_9_y0;
  assign f_s_dadda_rca24_fa76_y1 = f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_8_8_y0 & f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_7_9_y0;
  assign f_s_dadda_rca24_fa76_y2 = f_s_dadda_rca24_fa76_y0 ^ f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_6_10_y0;
  assign f_s_dadda_rca24_fa76_y3 = f_s_dadda_rca24_fa76_y0 & f_s_dadda_rca24_fa76_f_s_dadda_rca24_and_6_10_y0;
  assign f_s_dadda_rca24_fa76_y4 = f_s_dadda_rca24_fa76_y1 | f_s_dadda_rca24_fa76_y3;
  assign f_s_dadda_rca24_and_5_11_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_5_11_y0 = f_s_dadda_rca24_and_5_11_a_5 & f_s_dadda_rca24_and_5_11_b_11;
  assign f_s_dadda_rca24_and_4_12_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_4_12_y0 = f_s_dadda_rca24_and_4_12_a_4 & f_s_dadda_rca24_and_4_12_b_12;
  assign f_s_dadda_rca24_and_3_13_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_3_13_y0 = f_s_dadda_rca24_and_3_13_a_3 & f_s_dadda_rca24_and_3_13_b_13;
  assign f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_5_11_y0 = f_s_dadda_rca24_and_5_11_y0;
  assign f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_4_12_y0 = f_s_dadda_rca24_and_4_12_y0;
  assign f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_3_13_y0 = f_s_dadda_rca24_and_3_13_y0;
  assign f_s_dadda_rca24_fa77_y0 = f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_5_11_y0 ^ f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_4_12_y0;
  assign f_s_dadda_rca24_fa77_y1 = f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_5_11_y0 & f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_4_12_y0;
  assign f_s_dadda_rca24_fa77_y2 = f_s_dadda_rca24_fa77_y0 ^ f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_3_13_y0;
  assign f_s_dadda_rca24_fa77_y3 = f_s_dadda_rca24_fa77_y0 & f_s_dadda_rca24_fa77_f_s_dadda_rca24_and_3_13_y0;
  assign f_s_dadda_rca24_fa77_y4 = f_s_dadda_rca24_fa77_y1 | f_s_dadda_rca24_fa77_y3;
  assign f_s_dadda_rca24_and_2_14_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_2_14_y0 = f_s_dadda_rca24_and_2_14_a_2 & f_s_dadda_rca24_and_2_14_b_14;
  assign f_s_dadda_rca24_and_1_15_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_1_15_y0 = f_s_dadda_rca24_and_1_15_a_1 & f_s_dadda_rca24_and_1_15_b_15;
  assign f_s_dadda_rca24_and_0_16_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_0_16_y0 = f_s_dadda_rca24_and_0_16_a_0 & f_s_dadda_rca24_and_0_16_b_16;
  assign f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_2_14_y0 = f_s_dadda_rca24_and_2_14_y0;
  assign f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_1_15_y0 = f_s_dadda_rca24_and_1_15_y0;
  assign f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_0_16_y0 = f_s_dadda_rca24_and_0_16_y0;
  assign f_s_dadda_rca24_fa78_y0 = f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_2_14_y0 ^ f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_1_15_y0;
  assign f_s_dadda_rca24_fa78_y1 = f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_2_14_y0 & f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_1_15_y0;
  assign f_s_dadda_rca24_fa78_y2 = f_s_dadda_rca24_fa78_y0 ^ f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_0_16_y0;
  assign f_s_dadda_rca24_fa78_y3 = f_s_dadda_rca24_fa78_y0 & f_s_dadda_rca24_fa78_f_s_dadda_rca24_and_0_16_y0;
  assign f_s_dadda_rca24_fa78_y4 = f_s_dadda_rca24_fa78_y1 | f_s_dadda_rca24_fa78_y3;
  assign f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa70_y2 = f_s_dadda_rca24_fa70_y2;
  assign f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa71_y2 = f_s_dadda_rca24_fa71_y2;
  assign f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa72_y2 = f_s_dadda_rca24_fa72_y2;
  assign f_s_dadda_rca24_fa79_y0 = f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa70_y2 ^ f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa71_y2;
  assign f_s_dadda_rca24_fa79_y1 = f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa70_y2 & f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa71_y2;
  assign f_s_dadda_rca24_fa79_y2 = f_s_dadda_rca24_fa79_y0 ^ f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa72_y2;
  assign f_s_dadda_rca24_fa79_y3 = f_s_dadda_rca24_fa79_y0 & f_s_dadda_rca24_fa79_f_s_dadda_rca24_fa72_y2;
  assign f_s_dadda_rca24_fa79_y4 = f_s_dadda_rca24_fa79_y1 | f_s_dadda_rca24_fa79_y3;
  assign f_s_dadda_rca24_ha15_f_s_dadda_rca24_fa73_y2 = f_s_dadda_rca24_fa73_y2;
  assign f_s_dadda_rca24_ha15_f_s_dadda_rca24_fa74_y2 = f_s_dadda_rca24_fa74_y2;
  assign f_s_dadda_rca24_ha15_y0 = f_s_dadda_rca24_ha15_f_s_dadda_rca24_fa73_y2 ^ f_s_dadda_rca24_ha15_f_s_dadda_rca24_fa74_y2;
  assign f_s_dadda_rca24_ha15_y1 = f_s_dadda_rca24_ha15_f_s_dadda_rca24_fa73_y2 & f_s_dadda_rca24_ha15_f_s_dadda_rca24_fa74_y2;
  assign f_s_dadda_rca24_fa80_f_s_dadda_rca24_ha15_y1 = f_s_dadda_rca24_ha15_y1;
  assign f_s_dadda_rca24_fa80_f_s_dadda_rca24_fa79_y4 = f_s_dadda_rca24_fa79_y4;
  assign f_s_dadda_rca24_fa80_f_s_dadda_rca24_fa78_y4 = f_s_dadda_rca24_fa78_y4;
  assign f_s_dadda_rca24_fa80_y0 = f_s_dadda_rca24_fa80_f_s_dadda_rca24_ha15_y1 ^ f_s_dadda_rca24_fa80_f_s_dadda_rca24_fa79_y4;
  assign f_s_dadda_rca24_fa80_y1 = f_s_dadda_rca24_fa80_f_s_dadda_rca24_ha15_y1 & f_s_dadda_rca24_fa80_f_s_dadda_rca24_fa79_y4;
  assign f_s_dadda_rca24_fa80_y2 = f_s_dadda_rca24_fa80_y0 ^ f_s_dadda_rca24_fa80_f_s_dadda_rca24_fa78_y4;
  assign f_s_dadda_rca24_fa80_y3 = f_s_dadda_rca24_fa80_y0 & f_s_dadda_rca24_fa80_f_s_dadda_rca24_fa78_y4;
  assign f_s_dadda_rca24_fa80_y4 = f_s_dadda_rca24_fa80_y1 | f_s_dadda_rca24_fa80_y3;
  assign f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa77_y4 = f_s_dadda_rca24_fa77_y4;
  assign f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa76_y4 = f_s_dadda_rca24_fa76_y4;
  assign f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa75_y4 = f_s_dadda_rca24_fa75_y4;
  assign f_s_dadda_rca24_fa81_y0 = f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa77_y4 ^ f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa76_y4;
  assign f_s_dadda_rca24_fa81_y1 = f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa77_y4 & f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa76_y4;
  assign f_s_dadda_rca24_fa81_y2 = f_s_dadda_rca24_fa81_y0 ^ f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa75_y4;
  assign f_s_dadda_rca24_fa81_y3 = f_s_dadda_rca24_fa81_y0 & f_s_dadda_rca24_fa81_f_s_dadda_rca24_fa75_y4;
  assign f_s_dadda_rca24_fa81_y4 = f_s_dadda_rca24_fa81_y1 | f_s_dadda_rca24_fa81_y3;
  assign f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa74_y4 = f_s_dadda_rca24_fa74_y4;
  assign f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa73_y4 = f_s_dadda_rca24_fa73_y4;
  assign f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa72_y4 = f_s_dadda_rca24_fa72_y4;
  assign f_s_dadda_rca24_fa82_y0 = f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa74_y4 ^ f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa73_y4;
  assign f_s_dadda_rca24_fa82_y1 = f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa74_y4 & f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa73_y4;
  assign f_s_dadda_rca24_fa82_y2 = f_s_dadda_rca24_fa82_y0 ^ f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa72_y4;
  assign f_s_dadda_rca24_fa82_y3 = f_s_dadda_rca24_fa82_y0 & f_s_dadda_rca24_fa82_f_s_dadda_rca24_fa72_y4;
  assign f_s_dadda_rca24_fa82_y4 = f_s_dadda_rca24_fa82_y1 | f_s_dadda_rca24_fa82_y3;
  assign f_s_dadda_rca24_and_17_0_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_17_0_y0 = f_s_dadda_rca24_and_17_0_a_17 & f_s_dadda_rca24_and_17_0_b_0;
  assign f_s_dadda_rca24_fa83_f_s_dadda_rca24_fa71_y4 = f_s_dadda_rca24_fa71_y4;
  assign f_s_dadda_rca24_fa83_f_s_dadda_rca24_fa70_y4 = f_s_dadda_rca24_fa70_y4;
  assign f_s_dadda_rca24_fa83_f_s_dadda_rca24_and_17_0_y0 = f_s_dadda_rca24_and_17_0_y0;
  assign f_s_dadda_rca24_fa83_y0 = f_s_dadda_rca24_fa83_f_s_dadda_rca24_fa71_y4 ^ f_s_dadda_rca24_fa83_f_s_dadda_rca24_fa70_y4;
  assign f_s_dadda_rca24_fa83_y1 = f_s_dadda_rca24_fa83_f_s_dadda_rca24_fa71_y4 & f_s_dadda_rca24_fa83_f_s_dadda_rca24_fa70_y4;
  assign f_s_dadda_rca24_fa83_y2 = f_s_dadda_rca24_fa83_y0 ^ f_s_dadda_rca24_fa83_f_s_dadda_rca24_and_17_0_y0;
  assign f_s_dadda_rca24_fa83_y3 = f_s_dadda_rca24_fa83_y0 & f_s_dadda_rca24_fa83_f_s_dadda_rca24_and_17_0_y0;
  assign f_s_dadda_rca24_fa83_y4 = f_s_dadda_rca24_fa83_y1 | f_s_dadda_rca24_fa83_y3;
  assign f_s_dadda_rca24_and_16_1_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_16_1_y0 = f_s_dadda_rca24_and_16_1_a_16 & f_s_dadda_rca24_and_16_1_b_1;
  assign f_s_dadda_rca24_and_15_2_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_15_2_y0 = f_s_dadda_rca24_and_15_2_a_15 & f_s_dadda_rca24_and_15_2_b_2;
  assign f_s_dadda_rca24_and_14_3_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_14_3_y0 = f_s_dadda_rca24_and_14_3_a_14 & f_s_dadda_rca24_and_14_3_b_3;
  assign f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_16_1_y0 = f_s_dadda_rca24_and_16_1_y0;
  assign f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_15_2_y0 = f_s_dadda_rca24_and_15_2_y0;
  assign f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_14_3_y0 = f_s_dadda_rca24_and_14_3_y0;
  assign f_s_dadda_rca24_fa84_y0 = f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_16_1_y0 ^ f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_15_2_y0;
  assign f_s_dadda_rca24_fa84_y1 = f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_16_1_y0 & f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_15_2_y0;
  assign f_s_dadda_rca24_fa84_y2 = f_s_dadda_rca24_fa84_y0 ^ f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_14_3_y0;
  assign f_s_dadda_rca24_fa84_y3 = f_s_dadda_rca24_fa84_y0 & f_s_dadda_rca24_fa84_f_s_dadda_rca24_and_14_3_y0;
  assign f_s_dadda_rca24_fa84_y4 = f_s_dadda_rca24_fa84_y1 | f_s_dadda_rca24_fa84_y3;
  assign f_s_dadda_rca24_and_13_4_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_13_4_y0 = f_s_dadda_rca24_and_13_4_a_13 & f_s_dadda_rca24_and_13_4_b_4;
  assign f_s_dadda_rca24_and_12_5_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_12_5_y0 = f_s_dadda_rca24_and_12_5_a_12 & f_s_dadda_rca24_and_12_5_b_5;
  assign f_s_dadda_rca24_and_11_6_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_11_6_y0 = f_s_dadda_rca24_and_11_6_a_11 & f_s_dadda_rca24_and_11_6_b_6;
  assign f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_13_4_y0 = f_s_dadda_rca24_and_13_4_y0;
  assign f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_12_5_y0 = f_s_dadda_rca24_and_12_5_y0;
  assign f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_11_6_y0 = f_s_dadda_rca24_and_11_6_y0;
  assign f_s_dadda_rca24_fa85_y0 = f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_13_4_y0 ^ f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_12_5_y0;
  assign f_s_dadda_rca24_fa85_y1 = f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_13_4_y0 & f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_12_5_y0;
  assign f_s_dadda_rca24_fa85_y2 = f_s_dadda_rca24_fa85_y0 ^ f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_11_6_y0;
  assign f_s_dadda_rca24_fa85_y3 = f_s_dadda_rca24_fa85_y0 & f_s_dadda_rca24_fa85_f_s_dadda_rca24_and_11_6_y0;
  assign f_s_dadda_rca24_fa85_y4 = f_s_dadda_rca24_fa85_y1 | f_s_dadda_rca24_fa85_y3;
  assign f_s_dadda_rca24_and_10_7_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_10_7_y0 = f_s_dadda_rca24_and_10_7_a_10 & f_s_dadda_rca24_and_10_7_b_7;
  assign f_s_dadda_rca24_and_9_8_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_9_8_y0 = f_s_dadda_rca24_and_9_8_a_9 & f_s_dadda_rca24_and_9_8_b_8;
  assign f_s_dadda_rca24_and_8_9_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_8_9_y0 = f_s_dadda_rca24_and_8_9_a_8 & f_s_dadda_rca24_and_8_9_b_9;
  assign f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_10_7_y0 = f_s_dadda_rca24_and_10_7_y0;
  assign f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_9_8_y0 = f_s_dadda_rca24_and_9_8_y0;
  assign f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_8_9_y0 = f_s_dadda_rca24_and_8_9_y0;
  assign f_s_dadda_rca24_fa86_y0 = f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_10_7_y0 ^ f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_9_8_y0;
  assign f_s_dadda_rca24_fa86_y1 = f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_10_7_y0 & f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_9_8_y0;
  assign f_s_dadda_rca24_fa86_y2 = f_s_dadda_rca24_fa86_y0 ^ f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_8_9_y0;
  assign f_s_dadda_rca24_fa86_y3 = f_s_dadda_rca24_fa86_y0 & f_s_dadda_rca24_fa86_f_s_dadda_rca24_and_8_9_y0;
  assign f_s_dadda_rca24_fa86_y4 = f_s_dadda_rca24_fa86_y1 | f_s_dadda_rca24_fa86_y3;
  assign f_s_dadda_rca24_and_7_10_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_7_10_y0 = f_s_dadda_rca24_and_7_10_a_7 & f_s_dadda_rca24_and_7_10_b_10;
  assign f_s_dadda_rca24_and_6_11_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_6_11_y0 = f_s_dadda_rca24_and_6_11_a_6 & f_s_dadda_rca24_and_6_11_b_11;
  assign f_s_dadda_rca24_and_5_12_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_5_12_y0 = f_s_dadda_rca24_and_5_12_a_5 & f_s_dadda_rca24_and_5_12_b_12;
  assign f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_7_10_y0 = f_s_dadda_rca24_and_7_10_y0;
  assign f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_6_11_y0 = f_s_dadda_rca24_and_6_11_y0;
  assign f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_5_12_y0 = f_s_dadda_rca24_and_5_12_y0;
  assign f_s_dadda_rca24_fa87_y0 = f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_7_10_y0 ^ f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_6_11_y0;
  assign f_s_dadda_rca24_fa87_y1 = f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_7_10_y0 & f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_6_11_y0;
  assign f_s_dadda_rca24_fa87_y2 = f_s_dadda_rca24_fa87_y0 ^ f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_5_12_y0;
  assign f_s_dadda_rca24_fa87_y3 = f_s_dadda_rca24_fa87_y0 & f_s_dadda_rca24_fa87_f_s_dadda_rca24_and_5_12_y0;
  assign f_s_dadda_rca24_fa87_y4 = f_s_dadda_rca24_fa87_y1 | f_s_dadda_rca24_fa87_y3;
  assign f_s_dadda_rca24_and_4_13_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_4_13_y0 = f_s_dadda_rca24_and_4_13_a_4 & f_s_dadda_rca24_and_4_13_b_13;
  assign f_s_dadda_rca24_and_3_14_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_3_14_y0 = f_s_dadda_rca24_and_3_14_a_3 & f_s_dadda_rca24_and_3_14_b_14;
  assign f_s_dadda_rca24_and_2_15_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_2_15_y0 = f_s_dadda_rca24_and_2_15_a_2 & f_s_dadda_rca24_and_2_15_b_15;
  assign f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_4_13_y0 = f_s_dadda_rca24_and_4_13_y0;
  assign f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_3_14_y0 = f_s_dadda_rca24_and_3_14_y0;
  assign f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_2_15_y0 = f_s_dadda_rca24_and_2_15_y0;
  assign f_s_dadda_rca24_fa88_y0 = f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_4_13_y0 ^ f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_3_14_y0;
  assign f_s_dadda_rca24_fa88_y1 = f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_4_13_y0 & f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_3_14_y0;
  assign f_s_dadda_rca24_fa88_y2 = f_s_dadda_rca24_fa88_y0 ^ f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_2_15_y0;
  assign f_s_dadda_rca24_fa88_y3 = f_s_dadda_rca24_fa88_y0 & f_s_dadda_rca24_fa88_f_s_dadda_rca24_and_2_15_y0;
  assign f_s_dadda_rca24_fa88_y4 = f_s_dadda_rca24_fa88_y1 | f_s_dadda_rca24_fa88_y3;
  assign f_s_dadda_rca24_and_1_16_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_1_16_y0 = f_s_dadda_rca24_and_1_16_a_1 & f_s_dadda_rca24_and_1_16_b_16;
  assign f_s_dadda_rca24_and_0_17_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_0_17_y0 = f_s_dadda_rca24_and_0_17_a_0 & f_s_dadda_rca24_and_0_17_b_17;
  assign f_s_dadda_rca24_fa89_f_s_dadda_rca24_and_1_16_y0 = f_s_dadda_rca24_and_1_16_y0;
  assign f_s_dadda_rca24_fa89_f_s_dadda_rca24_and_0_17_y0 = f_s_dadda_rca24_and_0_17_y0;
  assign f_s_dadda_rca24_fa89_f_s_dadda_rca24_fa80_y2 = f_s_dadda_rca24_fa80_y2;
  assign f_s_dadda_rca24_fa89_y0 = f_s_dadda_rca24_fa89_f_s_dadda_rca24_and_1_16_y0 ^ f_s_dadda_rca24_fa89_f_s_dadda_rca24_and_0_17_y0;
  assign f_s_dadda_rca24_fa89_y1 = f_s_dadda_rca24_fa89_f_s_dadda_rca24_and_1_16_y0 & f_s_dadda_rca24_fa89_f_s_dadda_rca24_and_0_17_y0;
  assign f_s_dadda_rca24_fa89_y2 = f_s_dadda_rca24_fa89_y0 ^ f_s_dadda_rca24_fa89_f_s_dadda_rca24_fa80_y2;
  assign f_s_dadda_rca24_fa89_y3 = f_s_dadda_rca24_fa89_y0 & f_s_dadda_rca24_fa89_f_s_dadda_rca24_fa80_y2;
  assign f_s_dadda_rca24_fa89_y4 = f_s_dadda_rca24_fa89_y1 | f_s_dadda_rca24_fa89_y3;
  assign f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa81_y2 = f_s_dadda_rca24_fa81_y2;
  assign f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa82_y2 = f_s_dadda_rca24_fa82_y2;
  assign f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa83_y2 = f_s_dadda_rca24_fa83_y2;
  assign f_s_dadda_rca24_fa90_y0 = f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa81_y2 ^ f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa82_y2;
  assign f_s_dadda_rca24_fa90_y1 = f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa81_y2 & f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa82_y2;
  assign f_s_dadda_rca24_fa90_y2 = f_s_dadda_rca24_fa90_y0 ^ f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa83_y2;
  assign f_s_dadda_rca24_fa90_y3 = f_s_dadda_rca24_fa90_y0 & f_s_dadda_rca24_fa90_f_s_dadda_rca24_fa83_y2;
  assign f_s_dadda_rca24_fa90_y4 = f_s_dadda_rca24_fa90_y1 | f_s_dadda_rca24_fa90_y3;
  assign f_s_dadda_rca24_ha16_f_s_dadda_rca24_fa84_y2 = f_s_dadda_rca24_fa84_y2;
  assign f_s_dadda_rca24_ha16_f_s_dadda_rca24_fa85_y2 = f_s_dadda_rca24_fa85_y2;
  assign f_s_dadda_rca24_ha16_y0 = f_s_dadda_rca24_ha16_f_s_dadda_rca24_fa84_y2 ^ f_s_dadda_rca24_ha16_f_s_dadda_rca24_fa85_y2;
  assign f_s_dadda_rca24_ha16_y1 = f_s_dadda_rca24_ha16_f_s_dadda_rca24_fa84_y2 & f_s_dadda_rca24_ha16_f_s_dadda_rca24_fa85_y2;
  assign f_s_dadda_rca24_fa91_f_s_dadda_rca24_ha16_y1 = f_s_dadda_rca24_ha16_y1;
  assign f_s_dadda_rca24_fa91_f_s_dadda_rca24_fa90_y4 = f_s_dadda_rca24_fa90_y4;
  assign f_s_dadda_rca24_fa91_f_s_dadda_rca24_fa89_y4 = f_s_dadda_rca24_fa89_y4;
  assign f_s_dadda_rca24_fa91_y0 = f_s_dadda_rca24_fa91_f_s_dadda_rca24_ha16_y1 ^ f_s_dadda_rca24_fa91_f_s_dadda_rca24_fa90_y4;
  assign f_s_dadda_rca24_fa91_y1 = f_s_dadda_rca24_fa91_f_s_dadda_rca24_ha16_y1 & f_s_dadda_rca24_fa91_f_s_dadda_rca24_fa90_y4;
  assign f_s_dadda_rca24_fa91_y2 = f_s_dadda_rca24_fa91_y0 ^ f_s_dadda_rca24_fa91_f_s_dadda_rca24_fa89_y4;
  assign f_s_dadda_rca24_fa91_y3 = f_s_dadda_rca24_fa91_y0 & f_s_dadda_rca24_fa91_f_s_dadda_rca24_fa89_y4;
  assign f_s_dadda_rca24_fa91_y4 = f_s_dadda_rca24_fa91_y1 | f_s_dadda_rca24_fa91_y3;
  assign f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa88_y4 = f_s_dadda_rca24_fa88_y4;
  assign f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa87_y4 = f_s_dadda_rca24_fa87_y4;
  assign f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa86_y4 = f_s_dadda_rca24_fa86_y4;
  assign f_s_dadda_rca24_fa92_y0 = f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa88_y4 ^ f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa87_y4;
  assign f_s_dadda_rca24_fa92_y1 = f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa88_y4 & f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa87_y4;
  assign f_s_dadda_rca24_fa92_y2 = f_s_dadda_rca24_fa92_y0 ^ f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa86_y4;
  assign f_s_dadda_rca24_fa92_y3 = f_s_dadda_rca24_fa92_y0 & f_s_dadda_rca24_fa92_f_s_dadda_rca24_fa86_y4;
  assign f_s_dadda_rca24_fa92_y4 = f_s_dadda_rca24_fa92_y1 | f_s_dadda_rca24_fa92_y3;
  assign f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa85_y4 = f_s_dadda_rca24_fa85_y4;
  assign f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa84_y4 = f_s_dadda_rca24_fa84_y4;
  assign f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa83_y4 = f_s_dadda_rca24_fa83_y4;
  assign f_s_dadda_rca24_fa93_y0 = f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa85_y4 ^ f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa84_y4;
  assign f_s_dadda_rca24_fa93_y1 = f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa85_y4 & f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa84_y4;
  assign f_s_dadda_rca24_fa93_y2 = f_s_dadda_rca24_fa93_y0 ^ f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa83_y4;
  assign f_s_dadda_rca24_fa93_y3 = f_s_dadda_rca24_fa93_y0 & f_s_dadda_rca24_fa93_f_s_dadda_rca24_fa83_y4;
  assign f_s_dadda_rca24_fa93_y4 = f_s_dadda_rca24_fa93_y1 | f_s_dadda_rca24_fa93_y3;
  assign f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa82_y4 = f_s_dadda_rca24_fa82_y4;
  assign f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa81_y4 = f_s_dadda_rca24_fa81_y4;
  assign f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa80_y4 = f_s_dadda_rca24_fa80_y4;
  assign f_s_dadda_rca24_fa94_y0 = f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa82_y4 ^ f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa81_y4;
  assign f_s_dadda_rca24_fa94_y1 = f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa82_y4 & f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa81_y4;
  assign f_s_dadda_rca24_fa94_y2 = f_s_dadda_rca24_fa94_y0 ^ f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa80_y4;
  assign f_s_dadda_rca24_fa94_y3 = f_s_dadda_rca24_fa94_y0 & f_s_dadda_rca24_fa94_f_s_dadda_rca24_fa80_y4;
  assign f_s_dadda_rca24_fa94_y4 = f_s_dadda_rca24_fa94_y1 | f_s_dadda_rca24_fa94_y3;
  assign f_s_dadda_rca24_and_18_0_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_18_0_y0 = f_s_dadda_rca24_and_18_0_a_18 & f_s_dadda_rca24_and_18_0_b_0;
  assign f_s_dadda_rca24_and_17_1_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_17_1_y0 = f_s_dadda_rca24_and_17_1_a_17 & f_s_dadda_rca24_and_17_1_b_1;
  assign f_s_dadda_rca24_and_16_2_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_16_2_y0 = f_s_dadda_rca24_and_16_2_a_16 & f_s_dadda_rca24_and_16_2_b_2;
  assign f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_18_0_y0 = f_s_dadda_rca24_and_18_0_y0;
  assign f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_17_1_y0 = f_s_dadda_rca24_and_17_1_y0;
  assign f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_16_2_y0 = f_s_dadda_rca24_and_16_2_y0;
  assign f_s_dadda_rca24_fa95_y0 = f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_18_0_y0 ^ f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_17_1_y0;
  assign f_s_dadda_rca24_fa95_y1 = f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_18_0_y0 & f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_17_1_y0;
  assign f_s_dadda_rca24_fa95_y2 = f_s_dadda_rca24_fa95_y0 ^ f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_16_2_y0;
  assign f_s_dadda_rca24_fa95_y3 = f_s_dadda_rca24_fa95_y0 & f_s_dadda_rca24_fa95_f_s_dadda_rca24_and_16_2_y0;
  assign f_s_dadda_rca24_fa95_y4 = f_s_dadda_rca24_fa95_y1 | f_s_dadda_rca24_fa95_y3;
  assign f_s_dadda_rca24_and_15_3_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_15_3_y0 = f_s_dadda_rca24_and_15_3_a_15 & f_s_dadda_rca24_and_15_3_b_3;
  assign f_s_dadda_rca24_and_14_4_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_14_4_y0 = f_s_dadda_rca24_and_14_4_a_14 & f_s_dadda_rca24_and_14_4_b_4;
  assign f_s_dadda_rca24_and_13_5_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_13_5_y0 = f_s_dadda_rca24_and_13_5_a_13 & f_s_dadda_rca24_and_13_5_b_5;
  assign f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_15_3_y0 = f_s_dadda_rca24_and_15_3_y0;
  assign f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_14_4_y0 = f_s_dadda_rca24_and_14_4_y0;
  assign f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_13_5_y0 = f_s_dadda_rca24_and_13_5_y0;
  assign f_s_dadda_rca24_fa96_y0 = f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_15_3_y0 ^ f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_14_4_y0;
  assign f_s_dadda_rca24_fa96_y1 = f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_15_3_y0 & f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_14_4_y0;
  assign f_s_dadda_rca24_fa96_y2 = f_s_dadda_rca24_fa96_y0 ^ f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_13_5_y0;
  assign f_s_dadda_rca24_fa96_y3 = f_s_dadda_rca24_fa96_y0 & f_s_dadda_rca24_fa96_f_s_dadda_rca24_and_13_5_y0;
  assign f_s_dadda_rca24_fa96_y4 = f_s_dadda_rca24_fa96_y1 | f_s_dadda_rca24_fa96_y3;
  assign f_s_dadda_rca24_and_12_6_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_12_6_y0 = f_s_dadda_rca24_and_12_6_a_12 & f_s_dadda_rca24_and_12_6_b_6;
  assign f_s_dadda_rca24_and_11_7_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_11_7_y0 = f_s_dadda_rca24_and_11_7_a_11 & f_s_dadda_rca24_and_11_7_b_7;
  assign f_s_dadda_rca24_and_10_8_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_10_8_y0 = f_s_dadda_rca24_and_10_8_a_10 & f_s_dadda_rca24_and_10_8_b_8;
  assign f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_12_6_y0 = f_s_dadda_rca24_and_12_6_y0;
  assign f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_11_7_y0 = f_s_dadda_rca24_and_11_7_y0;
  assign f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_10_8_y0 = f_s_dadda_rca24_and_10_8_y0;
  assign f_s_dadda_rca24_fa97_y0 = f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_12_6_y0 ^ f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_11_7_y0;
  assign f_s_dadda_rca24_fa97_y1 = f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_12_6_y0 & f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_11_7_y0;
  assign f_s_dadda_rca24_fa97_y2 = f_s_dadda_rca24_fa97_y0 ^ f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_10_8_y0;
  assign f_s_dadda_rca24_fa97_y3 = f_s_dadda_rca24_fa97_y0 & f_s_dadda_rca24_fa97_f_s_dadda_rca24_and_10_8_y0;
  assign f_s_dadda_rca24_fa97_y4 = f_s_dadda_rca24_fa97_y1 | f_s_dadda_rca24_fa97_y3;
  assign f_s_dadda_rca24_and_9_9_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_9_9_y0 = f_s_dadda_rca24_and_9_9_a_9 & f_s_dadda_rca24_and_9_9_b_9;
  assign f_s_dadda_rca24_and_8_10_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_8_10_y0 = f_s_dadda_rca24_and_8_10_a_8 & f_s_dadda_rca24_and_8_10_b_10;
  assign f_s_dadda_rca24_and_7_11_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_7_11_y0 = f_s_dadda_rca24_and_7_11_a_7 & f_s_dadda_rca24_and_7_11_b_11;
  assign f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_9_9_y0 = f_s_dadda_rca24_and_9_9_y0;
  assign f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_8_10_y0 = f_s_dadda_rca24_and_8_10_y0;
  assign f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_7_11_y0 = f_s_dadda_rca24_and_7_11_y0;
  assign f_s_dadda_rca24_fa98_y0 = f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_9_9_y0 ^ f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_8_10_y0;
  assign f_s_dadda_rca24_fa98_y1 = f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_9_9_y0 & f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_8_10_y0;
  assign f_s_dadda_rca24_fa98_y2 = f_s_dadda_rca24_fa98_y0 ^ f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_7_11_y0;
  assign f_s_dadda_rca24_fa98_y3 = f_s_dadda_rca24_fa98_y0 & f_s_dadda_rca24_fa98_f_s_dadda_rca24_and_7_11_y0;
  assign f_s_dadda_rca24_fa98_y4 = f_s_dadda_rca24_fa98_y1 | f_s_dadda_rca24_fa98_y3;
  assign f_s_dadda_rca24_and_6_12_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_6_12_y0 = f_s_dadda_rca24_and_6_12_a_6 & f_s_dadda_rca24_and_6_12_b_12;
  assign f_s_dadda_rca24_and_5_13_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_5_13_y0 = f_s_dadda_rca24_and_5_13_a_5 & f_s_dadda_rca24_and_5_13_b_13;
  assign f_s_dadda_rca24_and_4_14_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_4_14_y0 = f_s_dadda_rca24_and_4_14_a_4 & f_s_dadda_rca24_and_4_14_b_14;
  assign f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_6_12_y0 = f_s_dadda_rca24_and_6_12_y0;
  assign f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_5_13_y0 = f_s_dadda_rca24_and_5_13_y0;
  assign f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_4_14_y0 = f_s_dadda_rca24_and_4_14_y0;
  assign f_s_dadda_rca24_fa99_y0 = f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_6_12_y0 ^ f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_5_13_y0;
  assign f_s_dadda_rca24_fa99_y1 = f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_6_12_y0 & f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_5_13_y0;
  assign f_s_dadda_rca24_fa99_y2 = f_s_dadda_rca24_fa99_y0 ^ f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_4_14_y0;
  assign f_s_dadda_rca24_fa99_y3 = f_s_dadda_rca24_fa99_y0 & f_s_dadda_rca24_fa99_f_s_dadda_rca24_and_4_14_y0;
  assign f_s_dadda_rca24_fa99_y4 = f_s_dadda_rca24_fa99_y1 | f_s_dadda_rca24_fa99_y3;
  assign f_s_dadda_rca24_and_3_15_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_3_15_y0 = f_s_dadda_rca24_and_3_15_a_3 & f_s_dadda_rca24_and_3_15_b_15;
  assign f_s_dadda_rca24_and_2_16_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_2_16_y0 = f_s_dadda_rca24_and_2_16_a_2 & f_s_dadda_rca24_and_2_16_b_16;
  assign f_s_dadda_rca24_and_1_17_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_1_17_y0 = f_s_dadda_rca24_and_1_17_a_1 & f_s_dadda_rca24_and_1_17_b_17;
  assign f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_3_15_y0 = f_s_dadda_rca24_and_3_15_y0;
  assign f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_2_16_y0 = f_s_dadda_rca24_and_2_16_y0;
  assign f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_1_17_y0 = f_s_dadda_rca24_and_1_17_y0;
  assign f_s_dadda_rca24_fa100_y0 = f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_3_15_y0 ^ f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_2_16_y0;
  assign f_s_dadda_rca24_fa100_y1 = f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_3_15_y0 & f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_2_16_y0;
  assign f_s_dadda_rca24_fa100_y2 = f_s_dadda_rca24_fa100_y0 ^ f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_1_17_y0;
  assign f_s_dadda_rca24_fa100_y3 = f_s_dadda_rca24_fa100_y0 & f_s_dadda_rca24_fa100_f_s_dadda_rca24_and_1_17_y0;
  assign f_s_dadda_rca24_fa100_y4 = f_s_dadda_rca24_fa100_y1 | f_s_dadda_rca24_fa100_y3;
  assign f_s_dadda_rca24_and_0_18_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_0_18_y0 = f_s_dadda_rca24_and_0_18_a_0 & f_s_dadda_rca24_and_0_18_b_18;
  assign f_s_dadda_rca24_fa101_f_s_dadda_rca24_and_0_18_y0 = f_s_dadda_rca24_and_0_18_y0;
  assign f_s_dadda_rca24_fa101_f_s_dadda_rca24_fa91_y2 = f_s_dadda_rca24_fa91_y2;
  assign f_s_dadda_rca24_fa101_f_s_dadda_rca24_fa92_y2 = f_s_dadda_rca24_fa92_y2;
  assign f_s_dadda_rca24_fa101_y0 = f_s_dadda_rca24_fa101_f_s_dadda_rca24_and_0_18_y0 ^ f_s_dadda_rca24_fa101_f_s_dadda_rca24_fa91_y2;
  assign f_s_dadda_rca24_fa101_y1 = f_s_dadda_rca24_fa101_f_s_dadda_rca24_and_0_18_y0 & f_s_dadda_rca24_fa101_f_s_dadda_rca24_fa91_y2;
  assign f_s_dadda_rca24_fa101_y2 = f_s_dadda_rca24_fa101_y0 ^ f_s_dadda_rca24_fa101_f_s_dadda_rca24_fa92_y2;
  assign f_s_dadda_rca24_fa101_y3 = f_s_dadda_rca24_fa101_y0 & f_s_dadda_rca24_fa101_f_s_dadda_rca24_fa92_y2;
  assign f_s_dadda_rca24_fa101_y4 = f_s_dadda_rca24_fa101_y1 | f_s_dadda_rca24_fa101_y3;
  assign f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa93_y2 = f_s_dadda_rca24_fa93_y2;
  assign f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa94_y2 = f_s_dadda_rca24_fa94_y2;
  assign f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa95_y2 = f_s_dadda_rca24_fa95_y2;
  assign f_s_dadda_rca24_fa102_y0 = f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa93_y2 ^ f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa94_y2;
  assign f_s_dadda_rca24_fa102_y1 = f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa93_y2 & f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa94_y2;
  assign f_s_dadda_rca24_fa102_y2 = f_s_dadda_rca24_fa102_y0 ^ f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa95_y2;
  assign f_s_dadda_rca24_fa102_y3 = f_s_dadda_rca24_fa102_y0 & f_s_dadda_rca24_fa102_f_s_dadda_rca24_fa95_y2;
  assign f_s_dadda_rca24_fa102_y4 = f_s_dadda_rca24_fa102_y1 | f_s_dadda_rca24_fa102_y3;
  assign f_s_dadda_rca24_ha17_f_s_dadda_rca24_fa96_y2 = f_s_dadda_rca24_fa96_y2;
  assign f_s_dadda_rca24_ha17_f_s_dadda_rca24_fa97_y2 = f_s_dadda_rca24_fa97_y2;
  assign f_s_dadda_rca24_ha17_y0 = f_s_dadda_rca24_ha17_f_s_dadda_rca24_fa96_y2 ^ f_s_dadda_rca24_ha17_f_s_dadda_rca24_fa97_y2;
  assign f_s_dadda_rca24_ha17_y1 = f_s_dadda_rca24_ha17_f_s_dadda_rca24_fa96_y2 & f_s_dadda_rca24_ha17_f_s_dadda_rca24_fa97_y2;
  assign f_s_dadda_rca24_fa103_f_s_dadda_rca24_ha17_y1 = f_s_dadda_rca24_ha17_y1;
  assign f_s_dadda_rca24_fa103_f_s_dadda_rca24_fa102_y4 = f_s_dadda_rca24_fa102_y4;
  assign f_s_dadda_rca24_fa103_f_s_dadda_rca24_fa101_y4 = f_s_dadda_rca24_fa101_y4;
  assign f_s_dadda_rca24_fa103_y0 = f_s_dadda_rca24_fa103_f_s_dadda_rca24_ha17_y1 ^ f_s_dadda_rca24_fa103_f_s_dadda_rca24_fa102_y4;
  assign f_s_dadda_rca24_fa103_y1 = f_s_dadda_rca24_fa103_f_s_dadda_rca24_ha17_y1 & f_s_dadda_rca24_fa103_f_s_dadda_rca24_fa102_y4;
  assign f_s_dadda_rca24_fa103_y2 = f_s_dadda_rca24_fa103_y0 ^ f_s_dadda_rca24_fa103_f_s_dadda_rca24_fa101_y4;
  assign f_s_dadda_rca24_fa103_y3 = f_s_dadda_rca24_fa103_y0 & f_s_dadda_rca24_fa103_f_s_dadda_rca24_fa101_y4;
  assign f_s_dadda_rca24_fa103_y4 = f_s_dadda_rca24_fa103_y1 | f_s_dadda_rca24_fa103_y3;
  assign f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa100_y4 = f_s_dadda_rca24_fa100_y4;
  assign f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa99_y4 = f_s_dadda_rca24_fa99_y4;
  assign f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa98_y4 = f_s_dadda_rca24_fa98_y4;
  assign f_s_dadda_rca24_fa104_y0 = f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa100_y4 ^ f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa99_y4;
  assign f_s_dadda_rca24_fa104_y1 = f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa100_y4 & f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa99_y4;
  assign f_s_dadda_rca24_fa104_y2 = f_s_dadda_rca24_fa104_y0 ^ f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa98_y4;
  assign f_s_dadda_rca24_fa104_y3 = f_s_dadda_rca24_fa104_y0 & f_s_dadda_rca24_fa104_f_s_dadda_rca24_fa98_y4;
  assign f_s_dadda_rca24_fa104_y4 = f_s_dadda_rca24_fa104_y1 | f_s_dadda_rca24_fa104_y3;
  assign f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa97_y4 = f_s_dadda_rca24_fa97_y4;
  assign f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa96_y4 = f_s_dadda_rca24_fa96_y4;
  assign f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa95_y4 = f_s_dadda_rca24_fa95_y4;
  assign f_s_dadda_rca24_fa105_y0 = f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa97_y4 ^ f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa96_y4;
  assign f_s_dadda_rca24_fa105_y1 = f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa97_y4 & f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa96_y4;
  assign f_s_dadda_rca24_fa105_y2 = f_s_dadda_rca24_fa105_y0 ^ f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa95_y4;
  assign f_s_dadda_rca24_fa105_y3 = f_s_dadda_rca24_fa105_y0 & f_s_dadda_rca24_fa105_f_s_dadda_rca24_fa95_y4;
  assign f_s_dadda_rca24_fa105_y4 = f_s_dadda_rca24_fa105_y1 | f_s_dadda_rca24_fa105_y3;
  assign f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa94_y4 = f_s_dadda_rca24_fa94_y4;
  assign f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa93_y4 = f_s_dadda_rca24_fa93_y4;
  assign f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa92_y4 = f_s_dadda_rca24_fa92_y4;
  assign f_s_dadda_rca24_fa106_y0 = f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa94_y4 ^ f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa93_y4;
  assign f_s_dadda_rca24_fa106_y1 = f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa94_y4 & f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa93_y4;
  assign f_s_dadda_rca24_fa106_y2 = f_s_dadda_rca24_fa106_y0 ^ f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa92_y4;
  assign f_s_dadda_rca24_fa106_y3 = f_s_dadda_rca24_fa106_y0 & f_s_dadda_rca24_fa106_f_s_dadda_rca24_fa92_y4;
  assign f_s_dadda_rca24_fa106_y4 = f_s_dadda_rca24_fa106_y1 | f_s_dadda_rca24_fa106_y3;
  assign f_s_dadda_rca24_and_17_2_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_17_2_y0 = f_s_dadda_rca24_and_17_2_a_17 & f_s_dadda_rca24_and_17_2_b_2;
  assign f_s_dadda_rca24_and_16_3_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_16_3_y0 = f_s_dadda_rca24_and_16_3_a_16 & f_s_dadda_rca24_and_16_3_b_3;
  assign f_s_dadda_rca24_fa107_f_s_dadda_rca24_fa91_y4 = f_s_dadda_rca24_fa91_y4;
  assign f_s_dadda_rca24_fa107_f_s_dadda_rca24_and_17_2_y0 = f_s_dadda_rca24_and_17_2_y0;
  assign f_s_dadda_rca24_fa107_f_s_dadda_rca24_and_16_3_y0 = f_s_dadda_rca24_and_16_3_y0;
  assign f_s_dadda_rca24_fa107_y0 = f_s_dadda_rca24_fa107_f_s_dadda_rca24_fa91_y4 ^ f_s_dadda_rca24_fa107_f_s_dadda_rca24_and_17_2_y0;
  assign f_s_dadda_rca24_fa107_y1 = f_s_dadda_rca24_fa107_f_s_dadda_rca24_fa91_y4 & f_s_dadda_rca24_fa107_f_s_dadda_rca24_and_17_2_y0;
  assign f_s_dadda_rca24_fa107_y2 = f_s_dadda_rca24_fa107_y0 ^ f_s_dadda_rca24_fa107_f_s_dadda_rca24_and_16_3_y0;
  assign f_s_dadda_rca24_fa107_y3 = f_s_dadda_rca24_fa107_y0 & f_s_dadda_rca24_fa107_f_s_dadda_rca24_and_16_3_y0;
  assign f_s_dadda_rca24_fa107_y4 = f_s_dadda_rca24_fa107_y1 | f_s_dadda_rca24_fa107_y3;
  assign f_s_dadda_rca24_and_15_4_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_15_4_y0 = f_s_dadda_rca24_and_15_4_a_15 & f_s_dadda_rca24_and_15_4_b_4;
  assign f_s_dadda_rca24_and_14_5_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_14_5_y0 = f_s_dadda_rca24_and_14_5_a_14 & f_s_dadda_rca24_and_14_5_b_5;
  assign f_s_dadda_rca24_and_13_6_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_13_6_y0 = f_s_dadda_rca24_and_13_6_a_13 & f_s_dadda_rca24_and_13_6_b_6;
  assign f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_15_4_y0 = f_s_dadda_rca24_and_15_4_y0;
  assign f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_14_5_y0 = f_s_dadda_rca24_and_14_5_y0;
  assign f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_13_6_y0 = f_s_dadda_rca24_and_13_6_y0;
  assign f_s_dadda_rca24_fa108_y0 = f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_15_4_y0 ^ f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_14_5_y0;
  assign f_s_dadda_rca24_fa108_y1 = f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_15_4_y0 & f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_14_5_y0;
  assign f_s_dadda_rca24_fa108_y2 = f_s_dadda_rca24_fa108_y0 ^ f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_13_6_y0;
  assign f_s_dadda_rca24_fa108_y3 = f_s_dadda_rca24_fa108_y0 & f_s_dadda_rca24_fa108_f_s_dadda_rca24_and_13_6_y0;
  assign f_s_dadda_rca24_fa108_y4 = f_s_dadda_rca24_fa108_y1 | f_s_dadda_rca24_fa108_y3;
  assign f_s_dadda_rca24_and_12_7_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_12_7_y0 = f_s_dadda_rca24_and_12_7_a_12 & f_s_dadda_rca24_and_12_7_b_7;
  assign f_s_dadda_rca24_and_11_8_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_11_8_y0 = f_s_dadda_rca24_and_11_8_a_11 & f_s_dadda_rca24_and_11_8_b_8;
  assign f_s_dadda_rca24_and_10_9_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_10_9_y0 = f_s_dadda_rca24_and_10_9_a_10 & f_s_dadda_rca24_and_10_9_b_9;
  assign f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_12_7_y0 = f_s_dadda_rca24_and_12_7_y0;
  assign f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_11_8_y0 = f_s_dadda_rca24_and_11_8_y0;
  assign f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_10_9_y0 = f_s_dadda_rca24_and_10_9_y0;
  assign f_s_dadda_rca24_fa109_y0 = f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_12_7_y0 ^ f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_11_8_y0;
  assign f_s_dadda_rca24_fa109_y1 = f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_12_7_y0 & f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_11_8_y0;
  assign f_s_dadda_rca24_fa109_y2 = f_s_dadda_rca24_fa109_y0 ^ f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_10_9_y0;
  assign f_s_dadda_rca24_fa109_y3 = f_s_dadda_rca24_fa109_y0 & f_s_dadda_rca24_fa109_f_s_dadda_rca24_and_10_9_y0;
  assign f_s_dadda_rca24_fa109_y4 = f_s_dadda_rca24_fa109_y1 | f_s_dadda_rca24_fa109_y3;
  assign f_s_dadda_rca24_and_9_10_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_9_10_y0 = f_s_dadda_rca24_and_9_10_a_9 & f_s_dadda_rca24_and_9_10_b_10;
  assign f_s_dadda_rca24_and_8_11_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_8_11_y0 = f_s_dadda_rca24_and_8_11_a_8 & f_s_dadda_rca24_and_8_11_b_11;
  assign f_s_dadda_rca24_and_7_12_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_7_12_y0 = f_s_dadda_rca24_and_7_12_a_7 & f_s_dadda_rca24_and_7_12_b_12;
  assign f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_9_10_y0 = f_s_dadda_rca24_and_9_10_y0;
  assign f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_8_11_y0 = f_s_dadda_rca24_and_8_11_y0;
  assign f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_7_12_y0 = f_s_dadda_rca24_and_7_12_y0;
  assign f_s_dadda_rca24_fa110_y0 = f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_9_10_y0 ^ f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_8_11_y0;
  assign f_s_dadda_rca24_fa110_y1 = f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_9_10_y0 & f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_8_11_y0;
  assign f_s_dadda_rca24_fa110_y2 = f_s_dadda_rca24_fa110_y0 ^ f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_7_12_y0;
  assign f_s_dadda_rca24_fa110_y3 = f_s_dadda_rca24_fa110_y0 & f_s_dadda_rca24_fa110_f_s_dadda_rca24_and_7_12_y0;
  assign f_s_dadda_rca24_fa110_y4 = f_s_dadda_rca24_fa110_y1 | f_s_dadda_rca24_fa110_y3;
  assign f_s_dadda_rca24_and_6_13_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_6_13_y0 = f_s_dadda_rca24_and_6_13_a_6 & f_s_dadda_rca24_and_6_13_b_13;
  assign f_s_dadda_rca24_and_5_14_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_5_14_y0 = f_s_dadda_rca24_and_5_14_a_5 & f_s_dadda_rca24_and_5_14_b_14;
  assign f_s_dadda_rca24_and_4_15_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_4_15_y0 = f_s_dadda_rca24_and_4_15_a_4 & f_s_dadda_rca24_and_4_15_b_15;
  assign f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_6_13_y0 = f_s_dadda_rca24_and_6_13_y0;
  assign f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_5_14_y0 = f_s_dadda_rca24_and_5_14_y0;
  assign f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_4_15_y0 = f_s_dadda_rca24_and_4_15_y0;
  assign f_s_dadda_rca24_fa111_y0 = f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_6_13_y0 ^ f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_5_14_y0;
  assign f_s_dadda_rca24_fa111_y1 = f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_6_13_y0 & f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_5_14_y0;
  assign f_s_dadda_rca24_fa111_y2 = f_s_dadda_rca24_fa111_y0 ^ f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_4_15_y0;
  assign f_s_dadda_rca24_fa111_y3 = f_s_dadda_rca24_fa111_y0 & f_s_dadda_rca24_fa111_f_s_dadda_rca24_and_4_15_y0;
  assign f_s_dadda_rca24_fa111_y4 = f_s_dadda_rca24_fa111_y1 | f_s_dadda_rca24_fa111_y3;
  assign f_s_dadda_rca24_and_3_16_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_3_16_y0 = f_s_dadda_rca24_and_3_16_a_3 & f_s_dadda_rca24_and_3_16_b_16;
  assign f_s_dadda_rca24_and_2_17_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_2_17_y0 = f_s_dadda_rca24_and_2_17_a_2 & f_s_dadda_rca24_and_2_17_b_17;
  assign f_s_dadda_rca24_and_1_18_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_1_18_y0 = f_s_dadda_rca24_and_1_18_a_1 & f_s_dadda_rca24_and_1_18_b_18;
  assign f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_3_16_y0 = f_s_dadda_rca24_and_3_16_y0;
  assign f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_2_17_y0 = f_s_dadda_rca24_and_2_17_y0;
  assign f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_1_18_y0 = f_s_dadda_rca24_and_1_18_y0;
  assign f_s_dadda_rca24_fa112_y0 = f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_3_16_y0 ^ f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_2_17_y0;
  assign f_s_dadda_rca24_fa112_y1 = f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_3_16_y0 & f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_2_17_y0;
  assign f_s_dadda_rca24_fa112_y2 = f_s_dadda_rca24_fa112_y0 ^ f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_1_18_y0;
  assign f_s_dadda_rca24_fa112_y3 = f_s_dadda_rca24_fa112_y0 & f_s_dadda_rca24_fa112_f_s_dadda_rca24_and_1_18_y0;
  assign f_s_dadda_rca24_fa112_y4 = f_s_dadda_rca24_fa112_y1 | f_s_dadda_rca24_fa112_y3;
  assign f_s_dadda_rca24_and_0_19_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_0_19_y0 = f_s_dadda_rca24_and_0_19_a_0 & f_s_dadda_rca24_and_0_19_b_19;
  assign f_s_dadda_rca24_fa113_f_s_dadda_rca24_and_0_19_y0 = f_s_dadda_rca24_and_0_19_y0;
  assign f_s_dadda_rca24_fa113_f_s_dadda_rca24_ha0_y0 = f_s_dadda_rca24_ha0_y0;
  assign f_s_dadda_rca24_fa113_f_s_dadda_rca24_fa103_y2 = f_s_dadda_rca24_fa103_y2;
  assign f_s_dadda_rca24_fa113_y0 = f_s_dadda_rca24_fa113_f_s_dadda_rca24_and_0_19_y0 ^ f_s_dadda_rca24_fa113_f_s_dadda_rca24_ha0_y0;
  assign f_s_dadda_rca24_fa113_y1 = f_s_dadda_rca24_fa113_f_s_dadda_rca24_and_0_19_y0 & f_s_dadda_rca24_fa113_f_s_dadda_rca24_ha0_y0;
  assign f_s_dadda_rca24_fa113_y2 = f_s_dadda_rca24_fa113_y0 ^ f_s_dadda_rca24_fa113_f_s_dadda_rca24_fa103_y2;
  assign f_s_dadda_rca24_fa113_y3 = f_s_dadda_rca24_fa113_y0 & f_s_dadda_rca24_fa113_f_s_dadda_rca24_fa103_y2;
  assign f_s_dadda_rca24_fa113_y4 = f_s_dadda_rca24_fa113_y1 | f_s_dadda_rca24_fa113_y3;
  assign f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa104_y2 = f_s_dadda_rca24_fa104_y2;
  assign f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa105_y2 = f_s_dadda_rca24_fa105_y2;
  assign f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa106_y2 = f_s_dadda_rca24_fa106_y2;
  assign f_s_dadda_rca24_fa114_y0 = f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa104_y2 ^ f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa105_y2;
  assign f_s_dadda_rca24_fa114_y1 = f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa104_y2 & f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa105_y2;
  assign f_s_dadda_rca24_fa114_y2 = f_s_dadda_rca24_fa114_y0 ^ f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa106_y2;
  assign f_s_dadda_rca24_fa114_y3 = f_s_dadda_rca24_fa114_y0 & f_s_dadda_rca24_fa114_f_s_dadda_rca24_fa106_y2;
  assign f_s_dadda_rca24_fa114_y4 = f_s_dadda_rca24_fa114_y1 | f_s_dadda_rca24_fa114_y3;
  assign f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa107_y2 = f_s_dadda_rca24_fa107_y2;
  assign f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa108_y2 = f_s_dadda_rca24_fa108_y2;
  assign f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa109_y2 = f_s_dadda_rca24_fa109_y2;
  assign f_s_dadda_rca24_fa115_y0 = f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa107_y2 ^ f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa108_y2;
  assign f_s_dadda_rca24_fa115_y1 = f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa107_y2 & f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa108_y2;
  assign f_s_dadda_rca24_fa115_y2 = f_s_dadda_rca24_fa115_y0 ^ f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa109_y2;
  assign f_s_dadda_rca24_fa115_y3 = f_s_dadda_rca24_fa115_y0 & f_s_dadda_rca24_fa115_f_s_dadda_rca24_fa109_y2;
  assign f_s_dadda_rca24_fa115_y4 = f_s_dadda_rca24_fa115_y1 | f_s_dadda_rca24_fa115_y3;
  assign f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa115_y4 = f_s_dadda_rca24_fa115_y4;
  assign f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa114_y4 = f_s_dadda_rca24_fa114_y4;
  assign f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa113_y4 = f_s_dadda_rca24_fa113_y4;
  assign f_s_dadda_rca24_fa116_y0 = f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa115_y4 ^ f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa114_y4;
  assign f_s_dadda_rca24_fa116_y1 = f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa115_y4 & f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa114_y4;
  assign f_s_dadda_rca24_fa116_y2 = f_s_dadda_rca24_fa116_y0 ^ f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa113_y4;
  assign f_s_dadda_rca24_fa116_y3 = f_s_dadda_rca24_fa116_y0 & f_s_dadda_rca24_fa116_f_s_dadda_rca24_fa113_y4;
  assign f_s_dadda_rca24_fa116_y4 = f_s_dadda_rca24_fa116_y1 | f_s_dadda_rca24_fa116_y3;
  assign f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa112_y4 = f_s_dadda_rca24_fa112_y4;
  assign f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa111_y4 = f_s_dadda_rca24_fa111_y4;
  assign f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa110_y4 = f_s_dadda_rca24_fa110_y4;
  assign f_s_dadda_rca24_fa117_y0 = f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa112_y4 ^ f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa111_y4;
  assign f_s_dadda_rca24_fa117_y1 = f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa112_y4 & f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa111_y4;
  assign f_s_dadda_rca24_fa117_y2 = f_s_dadda_rca24_fa117_y0 ^ f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa110_y4;
  assign f_s_dadda_rca24_fa117_y3 = f_s_dadda_rca24_fa117_y0 & f_s_dadda_rca24_fa117_f_s_dadda_rca24_fa110_y4;
  assign f_s_dadda_rca24_fa117_y4 = f_s_dadda_rca24_fa117_y1 | f_s_dadda_rca24_fa117_y3;
  assign f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa109_y4 = f_s_dadda_rca24_fa109_y4;
  assign f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa108_y4 = f_s_dadda_rca24_fa108_y4;
  assign f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa107_y4 = f_s_dadda_rca24_fa107_y4;
  assign f_s_dadda_rca24_fa118_y0 = f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa109_y4 ^ f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa108_y4;
  assign f_s_dadda_rca24_fa118_y1 = f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa109_y4 & f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa108_y4;
  assign f_s_dadda_rca24_fa118_y2 = f_s_dadda_rca24_fa118_y0 ^ f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa107_y4;
  assign f_s_dadda_rca24_fa118_y3 = f_s_dadda_rca24_fa118_y0 & f_s_dadda_rca24_fa118_f_s_dadda_rca24_fa107_y4;
  assign f_s_dadda_rca24_fa118_y4 = f_s_dadda_rca24_fa118_y1 | f_s_dadda_rca24_fa118_y3;
  assign f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa106_y4 = f_s_dadda_rca24_fa106_y4;
  assign f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa105_y4 = f_s_dadda_rca24_fa105_y4;
  assign f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa104_y4 = f_s_dadda_rca24_fa104_y4;
  assign f_s_dadda_rca24_fa119_y0 = f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa106_y4 ^ f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa105_y4;
  assign f_s_dadda_rca24_fa119_y1 = f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa106_y4 & f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa105_y4;
  assign f_s_dadda_rca24_fa119_y2 = f_s_dadda_rca24_fa119_y0 ^ f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa104_y4;
  assign f_s_dadda_rca24_fa119_y3 = f_s_dadda_rca24_fa119_y0 & f_s_dadda_rca24_fa119_f_s_dadda_rca24_fa104_y4;
  assign f_s_dadda_rca24_fa119_y4 = f_s_dadda_rca24_fa119_y1 | f_s_dadda_rca24_fa119_y3;
  assign f_s_dadda_rca24_and_16_4_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_16_4_y0 = f_s_dadda_rca24_and_16_4_a_16 & f_s_dadda_rca24_and_16_4_b_4;
  assign f_s_dadda_rca24_and_15_5_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_15_5_y0 = f_s_dadda_rca24_and_15_5_a_15 & f_s_dadda_rca24_and_15_5_b_5;
  assign f_s_dadda_rca24_fa120_f_s_dadda_rca24_fa103_y4 = f_s_dadda_rca24_fa103_y4;
  assign f_s_dadda_rca24_fa120_f_s_dadda_rca24_and_16_4_y0 = f_s_dadda_rca24_and_16_4_y0;
  assign f_s_dadda_rca24_fa120_f_s_dadda_rca24_and_15_5_y0 = f_s_dadda_rca24_and_15_5_y0;
  assign f_s_dadda_rca24_fa120_y0 = f_s_dadda_rca24_fa120_f_s_dadda_rca24_fa103_y4 ^ f_s_dadda_rca24_fa120_f_s_dadda_rca24_and_16_4_y0;
  assign f_s_dadda_rca24_fa120_y1 = f_s_dadda_rca24_fa120_f_s_dadda_rca24_fa103_y4 & f_s_dadda_rca24_fa120_f_s_dadda_rca24_and_16_4_y0;
  assign f_s_dadda_rca24_fa120_y2 = f_s_dadda_rca24_fa120_y0 ^ f_s_dadda_rca24_fa120_f_s_dadda_rca24_and_15_5_y0;
  assign f_s_dadda_rca24_fa120_y3 = f_s_dadda_rca24_fa120_y0 & f_s_dadda_rca24_fa120_f_s_dadda_rca24_and_15_5_y0;
  assign f_s_dadda_rca24_fa120_y4 = f_s_dadda_rca24_fa120_y1 | f_s_dadda_rca24_fa120_y3;
  assign f_s_dadda_rca24_and_14_6_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_14_6_y0 = f_s_dadda_rca24_and_14_6_a_14 & f_s_dadda_rca24_and_14_6_b_6;
  assign f_s_dadda_rca24_and_13_7_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_13_7_y0 = f_s_dadda_rca24_and_13_7_a_13 & f_s_dadda_rca24_and_13_7_b_7;
  assign f_s_dadda_rca24_and_12_8_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_12_8_y0 = f_s_dadda_rca24_and_12_8_a_12 & f_s_dadda_rca24_and_12_8_b_8;
  assign f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_14_6_y0 = f_s_dadda_rca24_and_14_6_y0;
  assign f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_13_7_y0 = f_s_dadda_rca24_and_13_7_y0;
  assign f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_12_8_y0 = f_s_dadda_rca24_and_12_8_y0;
  assign f_s_dadda_rca24_fa121_y0 = f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_14_6_y0 ^ f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_13_7_y0;
  assign f_s_dadda_rca24_fa121_y1 = f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_14_6_y0 & f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_13_7_y0;
  assign f_s_dadda_rca24_fa121_y2 = f_s_dadda_rca24_fa121_y0 ^ f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_12_8_y0;
  assign f_s_dadda_rca24_fa121_y3 = f_s_dadda_rca24_fa121_y0 & f_s_dadda_rca24_fa121_f_s_dadda_rca24_and_12_8_y0;
  assign f_s_dadda_rca24_fa121_y4 = f_s_dadda_rca24_fa121_y1 | f_s_dadda_rca24_fa121_y3;
  assign f_s_dadda_rca24_and_11_9_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_11_9_y0 = f_s_dadda_rca24_and_11_9_a_11 & f_s_dadda_rca24_and_11_9_b_9;
  assign f_s_dadda_rca24_and_10_10_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_10_10_y0 = f_s_dadda_rca24_and_10_10_a_10 & f_s_dadda_rca24_and_10_10_b_10;
  assign f_s_dadda_rca24_and_9_11_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_9_11_y0 = f_s_dadda_rca24_and_9_11_a_9 & f_s_dadda_rca24_and_9_11_b_11;
  assign f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_11_9_y0 = f_s_dadda_rca24_and_11_9_y0;
  assign f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_10_10_y0 = f_s_dadda_rca24_and_10_10_y0;
  assign f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_9_11_y0 = f_s_dadda_rca24_and_9_11_y0;
  assign f_s_dadda_rca24_fa122_y0 = f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_11_9_y0 ^ f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_10_10_y0;
  assign f_s_dadda_rca24_fa122_y1 = f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_11_9_y0 & f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_10_10_y0;
  assign f_s_dadda_rca24_fa122_y2 = f_s_dadda_rca24_fa122_y0 ^ f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_9_11_y0;
  assign f_s_dadda_rca24_fa122_y3 = f_s_dadda_rca24_fa122_y0 & f_s_dadda_rca24_fa122_f_s_dadda_rca24_and_9_11_y0;
  assign f_s_dadda_rca24_fa122_y4 = f_s_dadda_rca24_fa122_y1 | f_s_dadda_rca24_fa122_y3;
  assign f_s_dadda_rca24_and_8_12_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_8_12_y0 = f_s_dadda_rca24_and_8_12_a_8 & f_s_dadda_rca24_and_8_12_b_12;
  assign f_s_dadda_rca24_and_7_13_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_7_13_y0 = f_s_dadda_rca24_and_7_13_a_7 & f_s_dadda_rca24_and_7_13_b_13;
  assign f_s_dadda_rca24_and_6_14_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_6_14_y0 = f_s_dadda_rca24_and_6_14_a_6 & f_s_dadda_rca24_and_6_14_b_14;
  assign f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_8_12_y0 = f_s_dadda_rca24_and_8_12_y0;
  assign f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_7_13_y0 = f_s_dadda_rca24_and_7_13_y0;
  assign f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_6_14_y0 = f_s_dadda_rca24_and_6_14_y0;
  assign f_s_dadda_rca24_fa123_y0 = f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_8_12_y0 ^ f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_7_13_y0;
  assign f_s_dadda_rca24_fa123_y1 = f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_8_12_y0 & f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_7_13_y0;
  assign f_s_dadda_rca24_fa123_y2 = f_s_dadda_rca24_fa123_y0 ^ f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_6_14_y0;
  assign f_s_dadda_rca24_fa123_y3 = f_s_dadda_rca24_fa123_y0 & f_s_dadda_rca24_fa123_f_s_dadda_rca24_and_6_14_y0;
  assign f_s_dadda_rca24_fa123_y4 = f_s_dadda_rca24_fa123_y1 | f_s_dadda_rca24_fa123_y3;
  assign f_s_dadda_rca24_and_5_15_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_5_15_y0 = f_s_dadda_rca24_and_5_15_a_5 & f_s_dadda_rca24_and_5_15_b_15;
  assign f_s_dadda_rca24_and_4_16_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_4_16_y0 = f_s_dadda_rca24_and_4_16_a_4 & f_s_dadda_rca24_and_4_16_b_16;
  assign f_s_dadda_rca24_and_3_17_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_3_17_y0 = f_s_dadda_rca24_and_3_17_a_3 & f_s_dadda_rca24_and_3_17_b_17;
  assign f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_5_15_y0 = f_s_dadda_rca24_and_5_15_y0;
  assign f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_4_16_y0 = f_s_dadda_rca24_and_4_16_y0;
  assign f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_3_17_y0 = f_s_dadda_rca24_and_3_17_y0;
  assign f_s_dadda_rca24_fa124_y0 = f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_5_15_y0 ^ f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_4_16_y0;
  assign f_s_dadda_rca24_fa124_y1 = f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_5_15_y0 & f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_4_16_y0;
  assign f_s_dadda_rca24_fa124_y2 = f_s_dadda_rca24_fa124_y0 ^ f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_3_17_y0;
  assign f_s_dadda_rca24_fa124_y3 = f_s_dadda_rca24_fa124_y0 & f_s_dadda_rca24_fa124_f_s_dadda_rca24_and_3_17_y0;
  assign f_s_dadda_rca24_fa124_y4 = f_s_dadda_rca24_fa124_y1 | f_s_dadda_rca24_fa124_y3;
  assign f_s_dadda_rca24_and_2_18_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_2_18_y0 = f_s_dadda_rca24_and_2_18_a_2 & f_s_dadda_rca24_and_2_18_b_18;
  assign f_s_dadda_rca24_and_1_19_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_1_19_y0 = f_s_dadda_rca24_and_1_19_a_1 & f_s_dadda_rca24_and_1_19_b_19;
  assign f_s_dadda_rca24_and_0_20_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_0_20_y0 = f_s_dadda_rca24_and_0_20_a_0 & f_s_dadda_rca24_and_0_20_b_20;
  assign f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_2_18_y0 = f_s_dadda_rca24_and_2_18_y0;
  assign f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_1_19_y0 = f_s_dadda_rca24_and_1_19_y0;
  assign f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_0_20_y0 = f_s_dadda_rca24_and_0_20_y0;
  assign f_s_dadda_rca24_fa125_y0 = f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_2_18_y0 ^ f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_1_19_y0;
  assign f_s_dadda_rca24_fa125_y1 = f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_2_18_y0 & f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_1_19_y0;
  assign f_s_dadda_rca24_fa125_y2 = f_s_dadda_rca24_fa125_y0 ^ f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_0_20_y0;
  assign f_s_dadda_rca24_fa125_y3 = f_s_dadda_rca24_fa125_y0 & f_s_dadda_rca24_fa125_f_s_dadda_rca24_and_0_20_y0;
  assign f_s_dadda_rca24_fa125_y4 = f_s_dadda_rca24_fa125_y1 | f_s_dadda_rca24_fa125_y3;
  assign f_s_dadda_rca24_fa126_f_s_dadda_rca24_fa0_y2 = f_s_dadda_rca24_fa0_y2;
  assign f_s_dadda_rca24_fa126_f_s_dadda_rca24_ha1_y0 = f_s_dadda_rca24_ha1_y0;
  assign f_s_dadda_rca24_fa126_f_s_dadda_rca24_fa116_y2 = f_s_dadda_rca24_fa116_y2;
  assign f_s_dadda_rca24_fa126_y0 = f_s_dadda_rca24_fa126_f_s_dadda_rca24_fa0_y2 ^ f_s_dadda_rca24_fa126_f_s_dadda_rca24_ha1_y0;
  assign f_s_dadda_rca24_fa126_y1 = f_s_dadda_rca24_fa126_f_s_dadda_rca24_fa0_y2 & f_s_dadda_rca24_fa126_f_s_dadda_rca24_ha1_y0;
  assign f_s_dadda_rca24_fa126_y2 = f_s_dadda_rca24_fa126_y0 ^ f_s_dadda_rca24_fa126_f_s_dadda_rca24_fa116_y2;
  assign f_s_dadda_rca24_fa126_y3 = f_s_dadda_rca24_fa126_y0 & f_s_dadda_rca24_fa126_f_s_dadda_rca24_fa116_y2;
  assign f_s_dadda_rca24_fa126_y4 = f_s_dadda_rca24_fa126_y1 | f_s_dadda_rca24_fa126_y3;
  assign f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa117_y2 = f_s_dadda_rca24_fa117_y2;
  assign f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa118_y2 = f_s_dadda_rca24_fa118_y2;
  assign f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa119_y2 = f_s_dadda_rca24_fa119_y2;
  assign f_s_dadda_rca24_fa127_y0 = f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa117_y2 ^ f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa118_y2;
  assign f_s_dadda_rca24_fa127_y1 = f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa117_y2 & f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa118_y2;
  assign f_s_dadda_rca24_fa127_y2 = f_s_dadda_rca24_fa127_y0 ^ f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa119_y2;
  assign f_s_dadda_rca24_fa127_y3 = f_s_dadda_rca24_fa127_y0 & f_s_dadda_rca24_fa127_f_s_dadda_rca24_fa119_y2;
  assign f_s_dadda_rca24_fa127_y4 = f_s_dadda_rca24_fa127_y1 | f_s_dadda_rca24_fa127_y3;
  assign f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa120_y2 = f_s_dadda_rca24_fa120_y2;
  assign f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa121_y2 = f_s_dadda_rca24_fa121_y2;
  assign f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa122_y2 = f_s_dadda_rca24_fa122_y2;
  assign f_s_dadda_rca24_fa128_y0 = f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa120_y2 ^ f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa121_y2;
  assign f_s_dadda_rca24_fa128_y1 = f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa120_y2 & f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa121_y2;
  assign f_s_dadda_rca24_fa128_y2 = f_s_dadda_rca24_fa128_y0 ^ f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa122_y2;
  assign f_s_dadda_rca24_fa128_y3 = f_s_dadda_rca24_fa128_y0 & f_s_dadda_rca24_fa128_f_s_dadda_rca24_fa122_y2;
  assign f_s_dadda_rca24_fa128_y4 = f_s_dadda_rca24_fa128_y1 | f_s_dadda_rca24_fa128_y3;
  assign f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa128_y4 = f_s_dadda_rca24_fa128_y4;
  assign f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa127_y4 = f_s_dadda_rca24_fa127_y4;
  assign f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa126_y4 = f_s_dadda_rca24_fa126_y4;
  assign f_s_dadda_rca24_fa129_y0 = f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa128_y4 ^ f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa127_y4;
  assign f_s_dadda_rca24_fa129_y1 = f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa128_y4 & f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa127_y4;
  assign f_s_dadda_rca24_fa129_y2 = f_s_dadda_rca24_fa129_y0 ^ f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa126_y4;
  assign f_s_dadda_rca24_fa129_y3 = f_s_dadda_rca24_fa129_y0 & f_s_dadda_rca24_fa129_f_s_dadda_rca24_fa126_y4;
  assign f_s_dadda_rca24_fa129_y4 = f_s_dadda_rca24_fa129_y1 | f_s_dadda_rca24_fa129_y3;
  assign f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa125_y4 = f_s_dadda_rca24_fa125_y4;
  assign f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa124_y4 = f_s_dadda_rca24_fa124_y4;
  assign f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa123_y4 = f_s_dadda_rca24_fa123_y4;
  assign f_s_dadda_rca24_fa130_y0 = f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa125_y4 ^ f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa124_y4;
  assign f_s_dadda_rca24_fa130_y1 = f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa125_y4 & f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa124_y4;
  assign f_s_dadda_rca24_fa130_y2 = f_s_dadda_rca24_fa130_y0 ^ f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa123_y4;
  assign f_s_dadda_rca24_fa130_y3 = f_s_dadda_rca24_fa130_y0 & f_s_dadda_rca24_fa130_f_s_dadda_rca24_fa123_y4;
  assign f_s_dadda_rca24_fa130_y4 = f_s_dadda_rca24_fa130_y1 | f_s_dadda_rca24_fa130_y3;
  assign f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa122_y4 = f_s_dadda_rca24_fa122_y4;
  assign f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa121_y4 = f_s_dadda_rca24_fa121_y4;
  assign f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa120_y4 = f_s_dadda_rca24_fa120_y4;
  assign f_s_dadda_rca24_fa131_y0 = f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa122_y4 ^ f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa121_y4;
  assign f_s_dadda_rca24_fa131_y1 = f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa122_y4 & f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa121_y4;
  assign f_s_dadda_rca24_fa131_y2 = f_s_dadda_rca24_fa131_y0 ^ f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa120_y4;
  assign f_s_dadda_rca24_fa131_y3 = f_s_dadda_rca24_fa131_y0 & f_s_dadda_rca24_fa131_f_s_dadda_rca24_fa120_y4;
  assign f_s_dadda_rca24_fa131_y4 = f_s_dadda_rca24_fa131_y1 | f_s_dadda_rca24_fa131_y3;
  assign f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa119_y4 = f_s_dadda_rca24_fa119_y4;
  assign f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa118_y4 = f_s_dadda_rca24_fa118_y4;
  assign f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa117_y4 = f_s_dadda_rca24_fa117_y4;
  assign f_s_dadda_rca24_fa132_y0 = f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa119_y4 ^ f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa118_y4;
  assign f_s_dadda_rca24_fa132_y1 = f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa119_y4 & f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa118_y4;
  assign f_s_dadda_rca24_fa132_y2 = f_s_dadda_rca24_fa132_y0 ^ f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa117_y4;
  assign f_s_dadda_rca24_fa132_y3 = f_s_dadda_rca24_fa132_y0 & f_s_dadda_rca24_fa132_f_s_dadda_rca24_fa117_y4;
  assign f_s_dadda_rca24_fa132_y4 = f_s_dadda_rca24_fa132_y1 | f_s_dadda_rca24_fa132_y3;
  assign f_s_dadda_rca24_and_15_6_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_15_6_y0 = f_s_dadda_rca24_and_15_6_a_15 & f_s_dadda_rca24_and_15_6_b_6;
  assign f_s_dadda_rca24_and_14_7_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_14_7_y0 = f_s_dadda_rca24_and_14_7_a_14 & f_s_dadda_rca24_and_14_7_b_7;
  assign f_s_dadda_rca24_fa133_f_s_dadda_rca24_fa116_y4 = f_s_dadda_rca24_fa116_y4;
  assign f_s_dadda_rca24_fa133_f_s_dadda_rca24_and_15_6_y0 = f_s_dadda_rca24_and_15_6_y0;
  assign f_s_dadda_rca24_fa133_f_s_dadda_rca24_and_14_7_y0 = f_s_dadda_rca24_and_14_7_y0;
  assign f_s_dadda_rca24_fa133_y0 = f_s_dadda_rca24_fa133_f_s_dadda_rca24_fa116_y4 ^ f_s_dadda_rca24_fa133_f_s_dadda_rca24_and_15_6_y0;
  assign f_s_dadda_rca24_fa133_y1 = f_s_dadda_rca24_fa133_f_s_dadda_rca24_fa116_y4 & f_s_dadda_rca24_fa133_f_s_dadda_rca24_and_15_6_y0;
  assign f_s_dadda_rca24_fa133_y2 = f_s_dadda_rca24_fa133_y0 ^ f_s_dadda_rca24_fa133_f_s_dadda_rca24_and_14_7_y0;
  assign f_s_dadda_rca24_fa133_y3 = f_s_dadda_rca24_fa133_y0 & f_s_dadda_rca24_fa133_f_s_dadda_rca24_and_14_7_y0;
  assign f_s_dadda_rca24_fa133_y4 = f_s_dadda_rca24_fa133_y1 | f_s_dadda_rca24_fa133_y3;
  assign f_s_dadda_rca24_and_13_8_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_13_8_y0 = f_s_dadda_rca24_and_13_8_a_13 & f_s_dadda_rca24_and_13_8_b_8;
  assign f_s_dadda_rca24_and_12_9_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_12_9_y0 = f_s_dadda_rca24_and_12_9_a_12 & f_s_dadda_rca24_and_12_9_b_9;
  assign f_s_dadda_rca24_and_11_10_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_11_10_y0 = f_s_dadda_rca24_and_11_10_a_11 & f_s_dadda_rca24_and_11_10_b_10;
  assign f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_13_8_y0 = f_s_dadda_rca24_and_13_8_y0;
  assign f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_12_9_y0 = f_s_dadda_rca24_and_12_9_y0;
  assign f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_11_10_y0 = f_s_dadda_rca24_and_11_10_y0;
  assign f_s_dadda_rca24_fa134_y0 = f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_13_8_y0 ^ f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_12_9_y0;
  assign f_s_dadda_rca24_fa134_y1 = f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_13_8_y0 & f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_12_9_y0;
  assign f_s_dadda_rca24_fa134_y2 = f_s_dadda_rca24_fa134_y0 ^ f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_11_10_y0;
  assign f_s_dadda_rca24_fa134_y3 = f_s_dadda_rca24_fa134_y0 & f_s_dadda_rca24_fa134_f_s_dadda_rca24_and_11_10_y0;
  assign f_s_dadda_rca24_fa134_y4 = f_s_dadda_rca24_fa134_y1 | f_s_dadda_rca24_fa134_y3;
  assign f_s_dadda_rca24_and_10_11_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_10_11_y0 = f_s_dadda_rca24_and_10_11_a_10 & f_s_dadda_rca24_and_10_11_b_11;
  assign f_s_dadda_rca24_and_9_12_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_9_12_y0 = f_s_dadda_rca24_and_9_12_a_9 & f_s_dadda_rca24_and_9_12_b_12;
  assign f_s_dadda_rca24_and_8_13_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_8_13_y0 = f_s_dadda_rca24_and_8_13_a_8 & f_s_dadda_rca24_and_8_13_b_13;
  assign f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_10_11_y0 = f_s_dadda_rca24_and_10_11_y0;
  assign f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_9_12_y0 = f_s_dadda_rca24_and_9_12_y0;
  assign f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_8_13_y0 = f_s_dadda_rca24_and_8_13_y0;
  assign f_s_dadda_rca24_fa135_y0 = f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_10_11_y0 ^ f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_9_12_y0;
  assign f_s_dadda_rca24_fa135_y1 = f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_10_11_y0 & f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_9_12_y0;
  assign f_s_dadda_rca24_fa135_y2 = f_s_dadda_rca24_fa135_y0 ^ f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_8_13_y0;
  assign f_s_dadda_rca24_fa135_y3 = f_s_dadda_rca24_fa135_y0 & f_s_dadda_rca24_fa135_f_s_dadda_rca24_and_8_13_y0;
  assign f_s_dadda_rca24_fa135_y4 = f_s_dadda_rca24_fa135_y1 | f_s_dadda_rca24_fa135_y3;
  assign f_s_dadda_rca24_and_7_14_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_7_14_y0 = f_s_dadda_rca24_and_7_14_a_7 & f_s_dadda_rca24_and_7_14_b_14;
  assign f_s_dadda_rca24_and_6_15_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_6_15_y0 = f_s_dadda_rca24_and_6_15_a_6 & f_s_dadda_rca24_and_6_15_b_15;
  assign f_s_dadda_rca24_and_5_16_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_5_16_y0 = f_s_dadda_rca24_and_5_16_a_5 & f_s_dadda_rca24_and_5_16_b_16;
  assign f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_7_14_y0 = f_s_dadda_rca24_and_7_14_y0;
  assign f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_6_15_y0 = f_s_dadda_rca24_and_6_15_y0;
  assign f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_5_16_y0 = f_s_dadda_rca24_and_5_16_y0;
  assign f_s_dadda_rca24_fa136_y0 = f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_7_14_y0 ^ f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_6_15_y0;
  assign f_s_dadda_rca24_fa136_y1 = f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_7_14_y0 & f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_6_15_y0;
  assign f_s_dadda_rca24_fa136_y2 = f_s_dadda_rca24_fa136_y0 ^ f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_5_16_y0;
  assign f_s_dadda_rca24_fa136_y3 = f_s_dadda_rca24_fa136_y0 & f_s_dadda_rca24_fa136_f_s_dadda_rca24_and_5_16_y0;
  assign f_s_dadda_rca24_fa136_y4 = f_s_dadda_rca24_fa136_y1 | f_s_dadda_rca24_fa136_y3;
  assign f_s_dadda_rca24_and_4_17_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_4_17_y0 = f_s_dadda_rca24_and_4_17_a_4 & f_s_dadda_rca24_and_4_17_b_17;
  assign f_s_dadda_rca24_and_3_18_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_3_18_y0 = f_s_dadda_rca24_and_3_18_a_3 & f_s_dadda_rca24_and_3_18_b_18;
  assign f_s_dadda_rca24_and_2_19_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_2_19_y0 = f_s_dadda_rca24_and_2_19_a_2 & f_s_dadda_rca24_and_2_19_b_19;
  assign f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_4_17_y0 = f_s_dadda_rca24_and_4_17_y0;
  assign f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_3_18_y0 = f_s_dadda_rca24_and_3_18_y0;
  assign f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_2_19_y0 = f_s_dadda_rca24_and_2_19_y0;
  assign f_s_dadda_rca24_fa137_y0 = f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_4_17_y0 ^ f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_3_18_y0;
  assign f_s_dadda_rca24_fa137_y1 = f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_4_17_y0 & f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_3_18_y0;
  assign f_s_dadda_rca24_fa137_y2 = f_s_dadda_rca24_fa137_y0 ^ f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_2_19_y0;
  assign f_s_dadda_rca24_fa137_y3 = f_s_dadda_rca24_fa137_y0 & f_s_dadda_rca24_fa137_f_s_dadda_rca24_and_2_19_y0;
  assign f_s_dadda_rca24_fa137_y4 = f_s_dadda_rca24_fa137_y1 | f_s_dadda_rca24_fa137_y3;
  assign f_s_dadda_rca24_and_1_20_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_1_20_y0 = f_s_dadda_rca24_and_1_20_a_1 & f_s_dadda_rca24_and_1_20_b_20;
  assign f_s_dadda_rca24_and_0_21_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_0_21_y0 = f_s_dadda_rca24_and_0_21_a_0 & f_s_dadda_rca24_and_0_21_b_21;
  assign f_s_dadda_rca24_fa138_f_s_dadda_rca24_and_1_20_y0 = f_s_dadda_rca24_and_1_20_y0;
  assign f_s_dadda_rca24_fa138_f_s_dadda_rca24_and_0_21_y0 = f_s_dadda_rca24_and_0_21_y0;
  assign f_s_dadda_rca24_fa138_f_s_dadda_rca24_fa1_y2 = f_s_dadda_rca24_fa1_y2;
  assign f_s_dadda_rca24_fa138_y0 = f_s_dadda_rca24_fa138_f_s_dadda_rca24_and_1_20_y0 ^ f_s_dadda_rca24_fa138_f_s_dadda_rca24_and_0_21_y0;
  assign f_s_dadda_rca24_fa138_y1 = f_s_dadda_rca24_fa138_f_s_dadda_rca24_and_1_20_y0 & f_s_dadda_rca24_fa138_f_s_dadda_rca24_and_0_21_y0;
  assign f_s_dadda_rca24_fa138_y2 = f_s_dadda_rca24_fa138_y0 ^ f_s_dadda_rca24_fa138_f_s_dadda_rca24_fa1_y2;
  assign f_s_dadda_rca24_fa138_y3 = f_s_dadda_rca24_fa138_y0 & f_s_dadda_rca24_fa138_f_s_dadda_rca24_fa1_y2;
  assign f_s_dadda_rca24_fa138_y4 = f_s_dadda_rca24_fa138_y1 | f_s_dadda_rca24_fa138_y3;
  assign f_s_dadda_rca24_fa139_f_s_dadda_rca24_fa2_y2 = f_s_dadda_rca24_fa2_y2;
  assign f_s_dadda_rca24_fa139_f_s_dadda_rca24_ha2_y0 = f_s_dadda_rca24_ha2_y0;
  assign f_s_dadda_rca24_fa139_f_s_dadda_rca24_fa129_y2 = f_s_dadda_rca24_fa129_y2;
  assign f_s_dadda_rca24_fa139_y0 = f_s_dadda_rca24_fa139_f_s_dadda_rca24_fa2_y2 ^ f_s_dadda_rca24_fa139_f_s_dadda_rca24_ha2_y0;
  assign f_s_dadda_rca24_fa139_y1 = f_s_dadda_rca24_fa139_f_s_dadda_rca24_fa2_y2 & f_s_dadda_rca24_fa139_f_s_dadda_rca24_ha2_y0;
  assign f_s_dadda_rca24_fa139_y2 = f_s_dadda_rca24_fa139_y0 ^ f_s_dadda_rca24_fa139_f_s_dadda_rca24_fa129_y2;
  assign f_s_dadda_rca24_fa139_y3 = f_s_dadda_rca24_fa139_y0 & f_s_dadda_rca24_fa139_f_s_dadda_rca24_fa129_y2;
  assign f_s_dadda_rca24_fa139_y4 = f_s_dadda_rca24_fa139_y1 | f_s_dadda_rca24_fa139_y3;
  assign f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa130_y2 = f_s_dadda_rca24_fa130_y2;
  assign f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa131_y2 = f_s_dadda_rca24_fa131_y2;
  assign f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa132_y2 = f_s_dadda_rca24_fa132_y2;
  assign f_s_dadda_rca24_fa140_y0 = f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa130_y2 ^ f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa131_y2;
  assign f_s_dadda_rca24_fa140_y1 = f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa130_y2 & f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa131_y2;
  assign f_s_dadda_rca24_fa140_y2 = f_s_dadda_rca24_fa140_y0 ^ f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa132_y2;
  assign f_s_dadda_rca24_fa140_y3 = f_s_dadda_rca24_fa140_y0 & f_s_dadda_rca24_fa140_f_s_dadda_rca24_fa132_y2;
  assign f_s_dadda_rca24_fa140_y4 = f_s_dadda_rca24_fa140_y1 | f_s_dadda_rca24_fa140_y3;
  assign f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa133_y2 = f_s_dadda_rca24_fa133_y2;
  assign f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa134_y2 = f_s_dadda_rca24_fa134_y2;
  assign f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa135_y2 = f_s_dadda_rca24_fa135_y2;
  assign f_s_dadda_rca24_fa141_y0 = f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa133_y2 ^ f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa134_y2;
  assign f_s_dadda_rca24_fa141_y1 = f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa133_y2 & f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa134_y2;
  assign f_s_dadda_rca24_fa141_y2 = f_s_dadda_rca24_fa141_y0 ^ f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa135_y2;
  assign f_s_dadda_rca24_fa141_y3 = f_s_dadda_rca24_fa141_y0 & f_s_dadda_rca24_fa141_f_s_dadda_rca24_fa135_y2;
  assign f_s_dadda_rca24_fa141_y4 = f_s_dadda_rca24_fa141_y1 | f_s_dadda_rca24_fa141_y3;
  assign f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa141_y4 = f_s_dadda_rca24_fa141_y4;
  assign f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa140_y4 = f_s_dadda_rca24_fa140_y4;
  assign f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa139_y4 = f_s_dadda_rca24_fa139_y4;
  assign f_s_dadda_rca24_fa142_y0 = f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa141_y4 ^ f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa140_y4;
  assign f_s_dadda_rca24_fa142_y1 = f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa141_y4 & f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa140_y4;
  assign f_s_dadda_rca24_fa142_y2 = f_s_dadda_rca24_fa142_y0 ^ f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa139_y4;
  assign f_s_dadda_rca24_fa142_y3 = f_s_dadda_rca24_fa142_y0 & f_s_dadda_rca24_fa142_f_s_dadda_rca24_fa139_y4;
  assign f_s_dadda_rca24_fa142_y4 = f_s_dadda_rca24_fa142_y1 | f_s_dadda_rca24_fa142_y3;
  assign f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa138_y4 = f_s_dadda_rca24_fa138_y4;
  assign f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa137_y4 = f_s_dadda_rca24_fa137_y4;
  assign f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa136_y4 = f_s_dadda_rca24_fa136_y4;
  assign f_s_dadda_rca24_fa143_y0 = f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa138_y4 ^ f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa137_y4;
  assign f_s_dadda_rca24_fa143_y1 = f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa138_y4 & f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa137_y4;
  assign f_s_dadda_rca24_fa143_y2 = f_s_dadda_rca24_fa143_y0 ^ f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa136_y4;
  assign f_s_dadda_rca24_fa143_y3 = f_s_dadda_rca24_fa143_y0 & f_s_dadda_rca24_fa143_f_s_dadda_rca24_fa136_y4;
  assign f_s_dadda_rca24_fa143_y4 = f_s_dadda_rca24_fa143_y1 | f_s_dadda_rca24_fa143_y3;
  assign f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa135_y4 = f_s_dadda_rca24_fa135_y4;
  assign f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa134_y4 = f_s_dadda_rca24_fa134_y4;
  assign f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa133_y4 = f_s_dadda_rca24_fa133_y4;
  assign f_s_dadda_rca24_fa144_y0 = f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa135_y4 ^ f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa134_y4;
  assign f_s_dadda_rca24_fa144_y1 = f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa135_y4 & f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa134_y4;
  assign f_s_dadda_rca24_fa144_y2 = f_s_dadda_rca24_fa144_y0 ^ f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa133_y4;
  assign f_s_dadda_rca24_fa144_y3 = f_s_dadda_rca24_fa144_y0 & f_s_dadda_rca24_fa144_f_s_dadda_rca24_fa133_y4;
  assign f_s_dadda_rca24_fa144_y4 = f_s_dadda_rca24_fa144_y1 | f_s_dadda_rca24_fa144_y3;
  assign f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa132_y4 = f_s_dadda_rca24_fa132_y4;
  assign f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa131_y4 = f_s_dadda_rca24_fa131_y4;
  assign f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa130_y4 = f_s_dadda_rca24_fa130_y4;
  assign f_s_dadda_rca24_fa145_y0 = f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa132_y4 ^ f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa131_y4;
  assign f_s_dadda_rca24_fa145_y1 = f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa132_y4 & f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa131_y4;
  assign f_s_dadda_rca24_fa145_y2 = f_s_dadda_rca24_fa145_y0 ^ f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa130_y4;
  assign f_s_dadda_rca24_fa145_y3 = f_s_dadda_rca24_fa145_y0 & f_s_dadda_rca24_fa145_f_s_dadda_rca24_fa130_y4;
  assign f_s_dadda_rca24_fa145_y4 = f_s_dadda_rca24_fa145_y1 | f_s_dadda_rca24_fa145_y3;
  assign f_s_dadda_rca24_and_14_8_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_14_8_y0 = f_s_dadda_rca24_and_14_8_a_14 & f_s_dadda_rca24_and_14_8_b_8;
  assign f_s_dadda_rca24_and_13_9_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_13_9_y0 = f_s_dadda_rca24_and_13_9_a_13 & f_s_dadda_rca24_and_13_9_b_9;
  assign f_s_dadda_rca24_fa146_f_s_dadda_rca24_fa129_y4 = f_s_dadda_rca24_fa129_y4;
  assign f_s_dadda_rca24_fa146_f_s_dadda_rca24_and_14_8_y0 = f_s_dadda_rca24_and_14_8_y0;
  assign f_s_dadda_rca24_fa146_f_s_dadda_rca24_and_13_9_y0 = f_s_dadda_rca24_and_13_9_y0;
  assign f_s_dadda_rca24_fa146_y0 = f_s_dadda_rca24_fa146_f_s_dadda_rca24_fa129_y4 ^ f_s_dadda_rca24_fa146_f_s_dadda_rca24_and_14_8_y0;
  assign f_s_dadda_rca24_fa146_y1 = f_s_dadda_rca24_fa146_f_s_dadda_rca24_fa129_y4 & f_s_dadda_rca24_fa146_f_s_dadda_rca24_and_14_8_y0;
  assign f_s_dadda_rca24_fa146_y2 = f_s_dadda_rca24_fa146_y0 ^ f_s_dadda_rca24_fa146_f_s_dadda_rca24_and_13_9_y0;
  assign f_s_dadda_rca24_fa146_y3 = f_s_dadda_rca24_fa146_y0 & f_s_dadda_rca24_fa146_f_s_dadda_rca24_and_13_9_y0;
  assign f_s_dadda_rca24_fa146_y4 = f_s_dadda_rca24_fa146_y1 | f_s_dadda_rca24_fa146_y3;
  assign f_s_dadda_rca24_and_12_10_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_12_10_y0 = f_s_dadda_rca24_and_12_10_a_12 & f_s_dadda_rca24_and_12_10_b_10;
  assign f_s_dadda_rca24_and_11_11_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_11_11_y0 = f_s_dadda_rca24_and_11_11_a_11 & f_s_dadda_rca24_and_11_11_b_11;
  assign f_s_dadda_rca24_and_10_12_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_10_12_y0 = f_s_dadda_rca24_and_10_12_a_10 & f_s_dadda_rca24_and_10_12_b_12;
  assign f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_12_10_y0 = f_s_dadda_rca24_and_12_10_y0;
  assign f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_11_11_y0 = f_s_dadda_rca24_and_11_11_y0;
  assign f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_10_12_y0 = f_s_dadda_rca24_and_10_12_y0;
  assign f_s_dadda_rca24_fa147_y0 = f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_12_10_y0 ^ f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_11_11_y0;
  assign f_s_dadda_rca24_fa147_y1 = f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_12_10_y0 & f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_11_11_y0;
  assign f_s_dadda_rca24_fa147_y2 = f_s_dadda_rca24_fa147_y0 ^ f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_10_12_y0;
  assign f_s_dadda_rca24_fa147_y3 = f_s_dadda_rca24_fa147_y0 & f_s_dadda_rca24_fa147_f_s_dadda_rca24_and_10_12_y0;
  assign f_s_dadda_rca24_fa147_y4 = f_s_dadda_rca24_fa147_y1 | f_s_dadda_rca24_fa147_y3;
  assign f_s_dadda_rca24_and_9_13_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_9_13_y0 = f_s_dadda_rca24_and_9_13_a_9 & f_s_dadda_rca24_and_9_13_b_13;
  assign f_s_dadda_rca24_and_8_14_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_8_14_y0 = f_s_dadda_rca24_and_8_14_a_8 & f_s_dadda_rca24_and_8_14_b_14;
  assign f_s_dadda_rca24_and_7_15_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_7_15_y0 = f_s_dadda_rca24_and_7_15_a_7 & f_s_dadda_rca24_and_7_15_b_15;
  assign f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_9_13_y0 = f_s_dadda_rca24_and_9_13_y0;
  assign f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_8_14_y0 = f_s_dadda_rca24_and_8_14_y0;
  assign f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_7_15_y0 = f_s_dadda_rca24_and_7_15_y0;
  assign f_s_dadda_rca24_fa148_y0 = f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_9_13_y0 ^ f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_8_14_y0;
  assign f_s_dadda_rca24_fa148_y1 = f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_9_13_y0 & f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_8_14_y0;
  assign f_s_dadda_rca24_fa148_y2 = f_s_dadda_rca24_fa148_y0 ^ f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_7_15_y0;
  assign f_s_dadda_rca24_fa148_y3 = f_s_dadda_rca24_fa148_y0 & f_s_dadda_rca24_fa148_f_s_dadda_rca24_and_7_15_y0;
  assign f_s_dadda_rca24_fa148_y4 = f_s_dadda_rca24_fa148_y1 | f_s_dadda_rca24_fa148_y3;
  assign f_s_dadda_rca24_and_6_16_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_6_16_y0 = f_s_dadda_rca24_and_6_16_a_6 & f_s_dadda_rca24_and_6_16_b_16;
  assign f_s_dadda_rca24_and_5_17_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_5_17_y0 = f_s_dadda_rca24_and_5_17_a_5 & f_s_dadda_rca24_and_5_17_b_17;
  assign f_s_dadda_rca24_and_4_18_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_4_18_y0 = f_s_dadda_rca24_and_4_18_a_4 & f_s_dadda_rca24_and_4_18_b_18;
  assign f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_6_16_y0 = f_s_dadda_rca24_and_6_16_y0;
  assign f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_5_17_y0 = f_s_dadda_rca24_and_5_17_y0;
  assign f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_4_18_y0 = f_s_dadda_rca24_and_4_18_y0;
  assign f_s_dadda_rca24_fa149_y0 = f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_6_16_y0 ^ f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_5_17_y0;
  assign f_s_dadda_rca24_fa149_y1 = f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_6_16_y0 & f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_5_17_y0;
  assign f_s_dadda_rca24_fa149_y2 = f_s_dadda_rca24_fa149_y0 ^ f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_4_18_y0;
  assign f_s_dadda_rca24_fa149_y3 = f_s_dadda_rca24_fa149_y0 & f_s_dadda_rca24_fa149_f_s_dadda_rca24_and_4_18_y0;
  assign f_s_dadda_rca24_fa149_y4 = f_s_dadda_rca24_fa149_y1 | f_s_dadda_rca24_fa149_y3;
  assign f_s_dadda_rca24_and_3_19_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_3_19_y0 = f_s_dadda_rca24_and_3_19_a_3 & f_s_dadda_rca24_and_3_19_b_19;
  assign f_s_dadda_rca24_and_2_20_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_2_20_y0 = f_s_dadda_rca24_and_2_20_a_2 & f_s_dadda_rca24_and_2_20_b_20;
  assign f_s_dadda_rca24_and_1_21_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_1_21_y0 = f_s_dadda_rca24_and_1_21_a_1 & f_s_dadda_rca24_and_1_21_b_21;
  assign f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_3_19_y0 = f_s_dadda_rca24_and_3_19_y0;
  assign f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_2_20_y0 = f_s_dadda_rca24_and_2_20_y0;
  assign f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_1_21_y0 = f_s_dadda_rca24_and_1_21_y0;
  assign f_s_dadda_rca24_fa150_y0 = f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_3_19_y0 ^ f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_2_20_y0;
  assign f_s_dadda_rca24_fa150_y1 = f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_3_19_y0 & f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_2_20_y0;
  assign f_s_dadda_rca24_fa150_y2 = f_s_dadda_rca24_fa150_y0 ^ f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_1_21_y0;
  assign f_s_dadda_rca24_fa150_y3 = f_s_dadda_rca24_fa150_y0 & f_s_dadda_rca24_fa150_f_s_dadda_rca24_and_1_21_y0;
  assign f_s_dadda_rca24_fa150_y4 = f_s_dadda_rca24_fa150_y1 | f_s_dadda_rca24_fa150_y3;
  assign f_s_dadda_rca24_and_0_22_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_0_22_y0 = f_s_dadda_rca24_and_0_22_a_0 & f_s_dadda_rca24_and_0_22_b_22;
  assign f_s_dadda_rca24_fa151_f_s_dadda_rca24_and_0_22_y0 = f_s_dadda_rca24_and_0_22_y0;
  assign f_s_dadda_rca24_fa151_f_s_dadda_rca24_fa3_y2 = f_s_dadda_rca24_fa3_y2;
  assign f_s_dadda_rca24_fa151_f_s_dadda_rca24_fa4_y2 = f_s_dadda_rca24_fa4_y2;
  assign f_s_dadda_rca24_fa151_y0 = f_s_dadda_rca24_fa151_f_s_dadda_rca24_and_0_22_y0 ^ f_s_dadda_rca24_fa151_f_s_dadda_rca24_fa3_y2;
  assign f_s_dadda_rca24_fa151_y1 = f_s_dadda_rca24_fa151_f_s_dadda_rca24_and_0_22_y0 & f_s_dadda_rca24_fa151_f_s_dadda_rca24_fa3_y2;
  assign f_s_dadda_rca24_fa151_y2 = f_s_dadda_rca24_fa151_y0 ^ f_s_dadda_rca24_fa151_f_s_dadda_rca24_fa4_y2;
  assign f_s_dadda_rca24_fa151_y3 = f_s_dadda_rca24_fa151_y0 & f_s_dadda_rca24_fa151_f_s_dadda_rca24_fa4_y2;
  assign f_s_dadda_rca24_fa151_y4 = f_s_dadda_rca24_fa151_y1 | f_s_dadda_rca24_fa151_y3;
  assign f_s_dadda_rca24_fa152_f_s_dadda_rca24_fa5_y2 = f_s_dadda_rca24_fa5_y2;
  assign f_s_dadda_rca24_fa152_f_s_dadda_rca24_ha3_y0 = f_s_dadda_rca24_ha3_y0;
  assign f_s_dadda_rca24_fa152_f_s_dadda_rca24_fa142_y2 = f_s_dadda_rca24_fa142_y2;
  assign f_s_dadda_rca24_fa152_y0 = f_s_dadda_rca24_fa152_f_s_dadda_rca24_fa5_y2 ^ f_s_dadda_rca24_fa152_f_s_dadda_rca24_ha3_y0;
  assign f_s_dadda_rca24_fa152_y1 = f_s_dadda_rca24_fa152_f_s_dadda_rca24_fa5_y2 & f_s_dadda_rca24_fa152_f_s_dadda_rca24_ha3_y0;
  assign f_s_dadda_rca24_fa152_y2 = f_s_dadda_rca24_fa152_y0 ^ f_s_dadda_rca24_fa152_f_s_dadda_rca24_fa142_y2;
  assign f_s_dadda_rca24_fa152_y3 = f_s_dadda_rca24_fa152_y0 & f_s_dadda_rca24_fa152_f_s_dadda_rca24_fa142_y2;
  assign f_s_dadda_rca24_fa152_y4 = f_s_dadda_rca24_fa152_y1 | f_s_dadda_rca24_fa152_y3;
  assign f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa143_y2 = f_s_dadda_rca24_fa143_y2;
  assign f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa144_y2 = f_s_dadda_rca24_fa144_y2;
  assign f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa145_y2 = f_s_dadda_rca24_fa145_y2;
  assign f_s_dadda_rca24_fa153_y0 = f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa143_y2 ^ f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa144_y2;
  assign f_s_dadda_rca24_fa153_y1 = f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa143_y2 & f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa144_y2;
  assign f_s_dadda_rca24_fa153_y2 = f_s_dadda_rca24_fa153_y0 ^ f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa145_y2;
  assign f_s_dadda_rca24_fa153_y3 = f_s_dadda_rca24_fa153_y0 & f_s_dadda_rca24_fa153_f_s_dadda_rca24_fa145_y2;
  assign f_s_dadda_rca24_fa153_y4 = f_s_dadda_rca24_fa153_y1 | f_s_dadda_rca24_fa153_y3;
  assign f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa146_y2 = f_s_dadda_rca24_fa146_y2;
  assign f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa147_y2 = f_s_dadda_rca24_fa147_y2;
  assign f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa148_y2 = f_s_dadda_rca24_fa148_y2;
  assign f_s_dadda_rca24_fa154_y0 = f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa146_y2 ^ f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa147_y2;
  assign f_s_dadda_rca24_fa154_y1 = f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa146_y2 & f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa147_y2;
  assign f_s_dadda_rca24_fa154_y2 = f_s_dadda_rca24_fa154_y0 ^ f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa148_y2;
  assign f_s_dadda_rca24_fa154_y3 = f_s_dadda_rca24_fa154_y0 & f_s_dadda_rca24_fa154_f_s_dadda_rca24_fa148_y2;
  assign f_s_dadda_rca24_fa154_y4 = f_s_dadda_rca24_fa154_y1 | f_s_dadda_rca24_fa154_y3;
  assign f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa154_y4 = f_s_dadda_rca24_fa154_y4;
  assign f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa153_y4 = f_s_dadda_rca24_fa153_y4;
  assign f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa152_y4 = f_s_dadda_rca24_fa152_y4;
  assign f_s_dadda_rca24_fa155_y0 = f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa154_y4 ^ f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa153_y4;
  assign f_s_dadda_rca24_fa155_y1 = f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa154_y4 & f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa153_y4;
  assign f_s_dadda_rca24_fa155_y2 = f_s_dadda_rca24_fa155_y0 ^ f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa152_y4;
  assign f_s_dadda_rca24_fa155_y3 = f_s_dadda_rca24_fa155_y0 & f_s_dadda_rca24_fa155_f_s_dadda_rca24_fa152_y4;
  assign f_s_dadda_rca24_fa155_y4 = f_s_dadda_rca24_fa155_y1 | f_s_dadda_rca24_fa155_y3;
  assign f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa151_y4 = f_s_dadda_rca24_fa151_y4;
  assign f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa150_y4 = f_s_dadda_rca24_fa150_y4;
  assign f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa149_y4 = f_s_dadda_rca24_fa149_y4;
  assign f_s_dadda_rca24_fa156_y0 = f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa151_y4 ^ f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa150_y4;
  assign f_s_dadda_rca24_fa156_y1 = f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa151_y4 & f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa150_y4;
  assign f_s_dadda_rca24_fa156_y2 = f_s_dadda_rca24_fa156_y0 ^ f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa149_y4;
  assign f_s_dadda_rca24_fa156_y3 = f_s_dadda_rca24_fa156_y0 & f_s_dadda_rca24_fa156_f_s_dadda_rca24_fa149_y4;
  assign f_s_dadda_rca24_fa156_y4 = f_s_dadda_rca24_fa156_y1 | f_s_dadda_rca24_fa156_y3;
  assign f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa148_y4 = f_s_dadda_rca24_fa148_y4;
  assign f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa147_y4 = f_s_dadda_rca24_fa147_y4;
  assign f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa146_y4 = f_s_dadda_rca24_fa146_y4;
  assign f_s_dadda_rca24_fa157_y0 = f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa148_y4 ^ f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa147_y4;
  assign f_s_dadda_rca24_fa157_y1 = f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa148_y4 & f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa147_y4;
  assign f_s_dadda_rca24_fa157_y2 = f_s_dadda_rca24_fa157_y0 ^ f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa146_y4;
  assign f_s_dadda_rca24_fa157_y3 = f_s_dadda_rca24_fa157_y0 & f_s_dadda_rca24_fa157_f_s_dadda_rca24_fa146_y4;
  assign f_s_dadda_rca24_fa157_y4 = f_s_dadda_rca24_fa157_y1 | f_s_dadda_rca24_fa157_y3;
  assign f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa145_y4 = f_s_dadda_rca24_fa145_y4;
  assign f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa144_y4 = f_s_dadda_rca24_fa144_y4;
  assign f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa143_y4 = f_s_dadda_rca24_fa143_y4;
  assign f_s_dadda_rca24_fa158_y0 = f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa145_y4 ^ f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa144_y4;
  assign f_s_dadda_rca24_fa158_y1 = f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa145_y4 & f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa144_y4;
  assign f_s_dadda_rca24_fa158_y2 = f_s_dadda_rca24_fa158_y0 ^ f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa143_y4;
  assign f_s_dadda_rca24_fa158_y3 = f_s_dadda_rca24_fa158_y0 & f_s_dadda_rca24_fa158_f_s_dadda_rca24_fa143_y4;
  assign f_s_dadda_rca24_fa158_y4 = f_s_dadda_rca24_fa158_y1 | f_s_dadda_rca24_fa158_y3;
  assign f_s_dadda_rca24_and_13_10_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_13_10_y0 = f_s_dadda_rca24_and_13_10_a_13 & f_s_dadda_rca24_and_13_10_b_10;
  assign f_s_dadda_rca24_and_12_11_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_12_11_y0 = f_s_dadda_rca24_and_12_11_a_12 & f_s_dadda_rca24_and_12_11_b_11;
  assign f_s_dadda_rca24_fa159_f_s_dadda_rca24_fa142_y4 = f_s_dadda_rca24_fa142_y4;
  assign f_s_dadda_rca24_fa159_f_s_dadda_rca24_and_13_10_y0 = f_s_dadda_rca24_and_13_10_y0;
  assign f_s_dadda_rca24_fa159_f_s_dadda_rca24_and_12_11_y0 = f_s_dadda_rca24_and_12_11_y0;
  assign f_s_dadda_rca24_fa159_y0 = f_s_dadda_rca24_fa159_f_s_dadda_rca24_fa142_y4 ^ f_s_dadda_rca24_fa159_f_s_dadda_rca24_and_13_10_y0;
  assign f_s_dadda_rca24_fa159_y1 = f_s_dadda_rca24_fa159_f_s_dadda_rca24_fa142_y4 & f_s_dadda_rca24_fa159_f_s_dadda_rca24_and_13_10_y0;
  assign f_s_dadda_rca24_fa159_y2 = f_s_dadda_rca24_fa159_y0 ^ f_s_dadda_rca24_fa159_f_s_dadda_rca24_and_12_11_y0;
  assign f_s_dadda_rca24_fa159_y3 = f_s_dadda_rca24_fa159_y0 & f_s_dadda_rca24_fa159_f_s_dadda_rca24_and_12_11_y0;
  assign f_s_dadda_rca24_fa159_y4 = f_s_dadda_rca24_fa159_y1 | f_s_dadda_rca24_fa159_y3;
  assign f_s_dadda_rca24_and_11_12_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_11_12_y0 = f_s_dadda_rca24_and_11_12_a_11 & f_s_dadda_rca24_and_11_12_b_12;
  assign f_s_dadda_rca24_and_10_13_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_10_13_y0 = f_s_dadda_rca24_and_10_13_a_10 & f_s_dadda_rca24_and_10_13_b_13;
  assign f_s_dadda_rca24_and_9_14_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_9_14_y0 = f_s_dadda_rca24_and_9_14_a_9 & f_s_dadda_rca24_and_9_14_b_14;
  assign f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_11_12_y0 = f_s_dadda_rca24_and_11_12_y0;
  assign f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_10_13_y0 = f_s_dadda_rca24_and_10_13_y0;
  assign f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_9_14_y0 = f_s_dadda_rca24_and_9_14_y0;
  assign f_s_dadda_rca24_fa160_y0 = f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_11_12_y0 ^ f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_10_13_y0;
  assign f_s_dadda_rca24_fa160_y1 = f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_11_12_y0 & f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_10_13_y0;
  assign f_s_dadda_rca24_fa160_y2 = f_s_dadda_rca24_fa160_y0 ^ f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_9_14_y0;
  assign f_s_dadda_rca24_fa160_y3 = f_s_dadda_rca24_fa160_y0 & f_s_dadda_rca24_fa160_f_s_dadda_rca24_and_9_14_y0;
  assign f_s_dadda_rca24_fa160_y4 = f_s_dadda_rca24_fa160_y1 | f_s_dadda_rca24_fa160_y3;
  assign f_s_dadda_rca24_and_8_15_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_8_15_y0 = f_s_dadda_rca24_and_8_15_a_8 & f_s_dadda_rca24_and_8_15_b_15;
  assign f_s_dadda_rca24_and_7_16_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_7_16_y0 = f_s_dadda_rca24_and_7_16_a_7 & f_s_dadda_rca24_and_7_16_b_16;
  assign f_s_dadda_rca24_and_6_17_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_6_17_y0 = f_s_dadda_rca24_and_6_17_a_6 & f_s_dadda_rca24_and_6_17_b_17;
  assign f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_8_15_y0 = f_s_dadda_rca24_and_8_15_y0;
  assign f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_7_16_y0 = f_s_dadda_rca24_and_7_16_y0;
  assign f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_6_17_y0 = f_s_dadda_rca24_and_6_17_y0;
  assign f_s_dadda_rca24_fa161_y0 = f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_8_15_y0 ^ f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_7_16_y0;
  assign f_s_dadda_rca24_fa161_y1 = f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_8_15_y0 & f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_7_16_y0;
  assign f_s_dadda_rca24_fa161_y2 = f_s_dadda_rca24_fa161_y0 ^ f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_6_17_y0;
  assign f_s_dadda_rca24_fa161_y3 = f_s_dadda_rca24_fa161_y0 & f_s_dadda_rca24_fa161_f_s_dadda_rca24_and_6_17_y0;
  assign f_s_dadda_rca24_fa161_y4 = f_s_dadda_rca24_fa161_y1 | f_s_dadda_rca24_fa161_y3;
  assign f_s_dadda_rca24_and_5_18_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_5_18_y0 = f_s_dadda_rca24_and_5_18_a_5 & f_s_dadda_rca24_and_5_18_b_18;
  assign f_s_dadda_rca24_and_4_19_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_4_19_y0 = f_s_dadda_rca24_and_4_19_a_4 & f_s_dadda_rca24_and_4_19_b_19;
  assign f_s_dadda_rca24_and_3_20_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_3_20_y0 = f_s_dadda_rca24_and_3_20_a_3 & f_s_dadda_rca24_and_3_20_b_20;
  assign f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_5_18_y0 = f_s_dadda_rca24_and_5_18_y0;
  assign f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_4_19_y0 = f_s_dadda_rca24_and_4_19_y0;
  assign f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_3_20_y0 = f_s_dadda_rca24_and_3_20_y0;
  assign f_s_dadda_rca24_fa162_y0 = f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_5_18_y0 ^ f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_4_19_y0;
  assign f_s_dadda_rca24_fa162_y1 = f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_5_18_y0 & f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_4_19_y0;
  assign f_s_dadda_rca24_fa162_y2 = f_s_dadda_rca24_fa162_y0 ^ f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_3_20_y0;
  assign f_s_dadda_rca24_fa162_y3 = f_s_dadda_rca24_fa162_y0 & f_s_dadda_rca24_fa162_f_s_dadda_rca24_and_3_20_y0;
  assign f_s_dadda_rca24_fa162_y4 = f_s_dadda_rca24_fa162_y1 | f_s_dadda_rca24_fa162_y3;
  assign f_s_dadda_rca24_and_2_21_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_2_21_y0 = f_s_dadda_rca24_and_2_21_a_2 & f_s_dadda_rca24_and_2_21_b_21;
  assign f_s_dadda_rca24_and_1_22_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_1_22_y0 = f_s_dadda_rca24_and_1_22_a_1 & f_s_dadda_rca24_and_1_22_b_22;
  assign f_s_dadda_rca24_nand_0_23_a_0 = a_0;
  assign f_s_dadda_rca24_nand_0_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_0_23_y0 = ~(f_s_dadda_rca24_nand_0_23_a_0 & f_s_dadda_rca24_nand_0_23_b_23);
  assign f_s_dadda_rca24_fa163_f_s_dadda_rca24_and_2_21_y0 = f_s_dadda_rca24_and_2_21_y0;
  assign f_s_dadda_rca24_fa163_f_s_dadda_rca24_and_1_22_y0 = f_s_dadda_rca24_and_1_22_y0;
  assign f_s_dadda_rca24_fa163_f_s_dadda_rca24_nand_0_23_y0 = f_s_dadda_rca24_nand_0_23_y0;
  assign f_s_dadda_rca24_fa163_y0 = f_s_dadda_rca24_fa163_f_s_dadda_rca24_and_2_21_y0 ^ f_s_dadda_rca24_fa163_f_s_dadda_rca24_and_1_22_y0;
  assign f_s_dadda_rca24_fa163_y1 = f_s_dadda_rca24_fa163_f_s_dadda_rca24_and_2_21_y0 & f_s_dadda_rca24_fa163_f_s_dadda_rca24_and_1_22_y0;
  assign f_s_dadda_rca24_fa163_y2 = f_s_dadda_rca24_fa163_y0 ^ f_s_dadda_rca24_fa163_f_s_dadda_rca24_nand_0_23_y0;
  assign f_s_dadda_rca24_fa163_y3 = f_s_dadda_rca24_fa163_y0 & f_s_dadda_rca24_fa163_f_s_dadda_rca24_nand_0_23_y0;
  assign f_s_dadda_rca24_fa163_y4 = f_s_dadda_rca24_fa163_y1 | f_s_dadda_rca24_fa163_y3;
  assign f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa6_y2 = f_s_dadda_rca24_fa6_y2;
  assign f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa7_y2 = f_s_dadda_rca24_fa7_y2;
  assign f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa8_y2 = f_s_dadda_rca24_fa8_y2;
  assign f_s_dadda_rca24_fa164_y0 = f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa6_y2 ^ f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa7_y2;
  assign f_s_dadda_rca24_fa164_y1 = f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa6_y2 & f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa7_y2;
  assign f_s_dadda_rca24_fa164_y2 = f_s_dadda_rca24_fa164_y0 ^ f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa8_y2;
  assign f_s_dadda_rca24_fa164_y3 = f_s_dadda_rca24_fa164_y0 & f_s_dadda_rca24_fa164_f_s_dadda_rca24_fa8_y2;
  assign f_s_dadda_rca24_fa164_y4 = f_s_dadda_rca24_fa164_y1 | f_s_dadda_rca24_fa164_y3;
  assign f_s_dadda_rca24_fa165_f_s_dadda_rca24_fa9_y2 = f_s_dadda_rca24_fa9_y2;
  assign f_s_dadda_rca24_fa165_f_s_dadda_rca24_ha4_y0 = f_s_dadda_rca24_ha4_y0;
  assign f_s_dadda_rca24_fa165_f_s_dadda_rca24_fa155_y2 = f_s_dadda_rca24_fa155_y2;
  assign f_s_dadda_rca24_fa165_y0 = f_s_dadda_rca24_fa165_f_s_dadda_rca24_fa9_y2 ^ f_s_dadda_rca24_fa165_f_s_dadda_rca24_ha4_y0;
  assign f_s_dadda_rca24_fa165_y1 = f_s_dadda_rca24_fa165_f_s_dadda_rca24_fa9_y2 & f_s_dadda_rca24_fa165_f_s_dadda_rca24_ha4_y0;
  assign f_s_dadda_rca24_fa165_y2 = f_s_dadda_rca24_fa165_y0 ^ f_s_dadda_rca24_fa165_f_s_dadda_rca24_fa155_y2;
  assign f_s_dadda_rca24_fa165_y3 = f_s_dadda_rca24_fa165_y0 & f_s_dadda_rca24_fa165_f_s_dadda_rca24_fa155_y2;
  assign f_s_dadda_rca24_fa165_y4 = f_s_dadda_rca24_fa165_y1 | f_s_dadda_rca24_fa165_y3;
  assign f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa156_y2 = f_s_dadda_rca24_fa156_y2;
  assign f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa157_y2 = f_s_dadda_rca24_fa157_y2;
  assign f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa158_y2 = f_s_dadda_rca24_fa158_y2;
  assign f_s_dadda_rca24_fa166_y0 = f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa156_y2 ^ f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa157_y2;
  assign f_s_dadda_rca24_fa166_y1 = f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa156_y2 & f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa157_y2;
  assign f_s_dadda_rca24_fa166_y2 = f_s_dadda_rca24_fa166_y0 ^ f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa158_y2;
  assign f_s_dadda_rca24_fa166_y3 = f_s_dadda_rca24_fa166_y0 & f_s_dadda_rca24_fa166_f_s_dadda_rca24_fa158_y2;
  assign f_s_dadda_rca24_fa166_y4 = f_s_dadda_rca24_fa166_y1 | f_s_dadda_rca24_fa166_y3;
  assign f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa159_y2 = f_s_dadda_rca24_fa159_y2;
  assign f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa160_y2 = f_s_dadda_rca24_fa160_y2;
  assign f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa161_y2 = f_s_dadda_rca24_fa161_y2;
  assign f_s_dadda_rca24_fa167_y0 = f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa159_y2 ^ f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa160_y2;
  assign f_s_dadda_rca24_fa167_y1 = f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa159_y2 & f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa160_y2;
  assign f_s_dadda_rca24_fa167_y2 = f_s_dadda_rca24_fa167_y0 ^ f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa161_y2;
  assign f_s_dadda_rca24_fa167_y3 = f_s_dadda_rca24_fa167_y0 & f_s_dadda_rca24_fa167_f_s_dadda_rca24_fa161_y2;
  assign f_s_dadda_rca24_fa167_y4 = f_s_dadda_rca24_fa167_y1 | f_s_dadda_rca24_fa167_y3;
  assign f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa167_y4 = f_s_dadda_rca24_fa167_y4;
  assign f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa166_y4 = f_s_dadda_rca24_fa166_y4;
  assign f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa165_y4 = f_s_dadda_rca24_fa165_y4;
  assign f_s_dadda_rca24_fa168_y0 = f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa167_y4 ^ f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa166_y4;
  assign f_s_dadda_rca24_fa168_y1 = f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa167_y4 & f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa166_y4;
  assign f_s_dadda_rca24_fa168_y2 = f_s_dadda_rca24_fa168_y0 ^ f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa165_y4;
  assign f_s_dadda_rca24_fa168_y3 = f_s_dadda_rca24_fa168_y0 & f_s_dadda_rca24_fa168_f_s_dadda_rca24_fa165_y4;
  assign f_s_dadda_rca24_fa168_y4 = f_s_dadda_rca24_fa168_y1 | f_s_dadda_rca24_fa168_y3;
  assign f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa164_y4 = f_s_dadda_rca24_fa164_y4;
  assign f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa163_y4 = f_s_dadda_rca24_fa163_y4;
  assign f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa162_y4 = f_s_dadda_rca24_fa162_y4;
  assign f_s_dadda_rca24_fa169_y0 = f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa164_y4 ^ f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa163_y4;
  assign f_s_dadda_rca24_fa169_y1 = f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa164_y4 & f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa163_y4;
  assign f_s_dadda_rca24_fa169_y2 = f_s_dadda_rca24_fa169_y0 ^ f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa162_y4;
  assign f_s_dadda_rca24_fa169_y3 = f_s_dadda_rca24_fa169_y0 & f_s_dadda_rca24_fa169_f_s_dadda_rca24_fa162_y4;
  assign f_s_dadda_rca24_fa169_y4 = f_s_dadda_rca24_fa169_y1 | f_s_dadda_rca24_fa169_y3;
  assign f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa161_y4 = f_s_dadda_rca24_fa161_y4;
  assign f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa160_y4 = f_s_dadda_rca24_fa160_y4;
  assign f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa159_y4 = f_s_dadda_rca24_fa159_y4;
  assign f_s_dadda_rca24_fa170_y0 = f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa161_y4 ^ f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa160_y4;
  assign f_s_dadda_rca24_fa170_y1 = f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa161_y4 & f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa160_y4;
  assign f_s_dadda_rca24_fa170_y2 = f_s_dadda_rca24_fa170_y0 ^ f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa159_y4;
  assign f_s_dadda_rca24_fa170_y3 = f_s_dadda_rca24_fa170_y0 & f_s_dadda_rca24_fa170_f_s_dadda_rca24_fa159_y4;
  assign f_s_dadda_rca24_fa170_y4 = f_s_dadda_rca24_fa170_y1 | f_s_dadda_rca24_fa170_y3;
  assign f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa158_y4 = f_s_dadda_rca24_fa158_y4;
  assign f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa157_y4 = f_s_dadda_rca24_fa157_y4;
  assign f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa156_y4 = f_s_dadda_rca24_fa156_y4;
  assign f_s_dadda_rca24_fa171_y0 = f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa158_y4 ^ f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa157_y4;
  assign f_s_dadda_rca24_fa171_y1 = f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa158_y4 & f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa157_y4;
  assign f_s_dadda_rca24_fa171_y2 = f_s_dadda_rca24_fa171_y0 ^ f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa156_y4;
  assign f_s_dadda_rca24_fa171_y3 = f_s_dadda_rca24_fa171_y0 & f_s_dadda_rca24_fa171_f_s_dadda_rca24_fa156_y4;
  assign f_s_dadda_rca24_fa171_y4 = f_s_dadda_rca24_fa171_y1 | f_s_dadda_rca24_fa171_y3;
  assign f_s_dadda_rca24_and_14_10_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_14_10_y0 = f_s_dadda_rca24_and_14_10_a_14 & f_s_dadda_rca24_and_14_10_b_10;
  assign f_s_dadda_rca24_and_13_11_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_13_11_y0 = f_s_dadda_rca24_and_13_11_a_13 & f_s_dadda_rca24_and_13_11_b_11;
  assign f_s_dadda_rca24_fa172_f_s_dadda_rca24_fa155_y4 = f_s_dadda_rca24_fa155_y4;
  assign f_s_dadda_rca24_fa172_f_s_dadda_rca24_and_14_10_y0 = f_s_dadda_rca24_and_14_10_y0;
  assign f_s_dadda_rca24_fa172_f_s_dadda_rca24_and_13_11_y0 = f_s_dadda_rca24_and_13_11_y0;
  assign f_s_dadda_rca24_fa172_y0 = f_s_dadda_rca24_fa172_f_s_dadda_rca24_fa155_y4 ^ f_s_dadda_rca24_fa172_f_s_dadda_rca24_and_14_10_y0;
  assign f_s_dadda_rca24_fa172_y1 = f_s_dadda_rca24_fa172_f_s_dadda_rca24_fa155_y4 & f_s_dadda_rca24_fa172_f_s_dadda_rca24_and_14_10_y0;
  assign f_s_dadda_rca24_fa172_y2 = f_s_dadda_rca24_fa172_y0 ^ f_s_dadda_rca24_fa172_f_s_dadda_rca24_and_13_11_y0;
  assign f_s_dadda_rca24_fa172_y3 = f_s_dadda_rca24_fa172_y0 & f_s_dadda_rca24_fa172_f_s_dadda_rca24_and_13_11_y0;
  assign f_s_dadda_rca24_fa172_y4 = f_s_dadda_rca24_fa172_y1 | f_s_dadda_rca24_fa172_y3;
  assign f_s_dadda_rca24_and_12_12_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_12_12_y0 = f_s_dadda_rca24_and_12_12_a_12 & f_s_dadda_rca24_and_12_12_b_12;
  assign f_s_dadda_rca24_and_11_13_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_11_13_y0 = f_s_dadda_rca24_and_11_13_a_11 & f_s_dadda_rca24_and_11_13_b_13;
  assign f_s_dadda_rca24_and_10_14_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_10_14_y0 = f_s_dadda_rca24_and_10_14_a_10 & f_s_dadda_rca24_and_10_14_b_14;
  assign f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_12_12_y0 = f_s_dadda_rca24_and_12_12_y0;
  assign f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_11_13_y0 = f_s_dadda_rca24_and_11_13_y0;
  assign f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_10_14_y0 = f_s_dadda_rca24_and_10_14_y0;
  assign f_s_dadda_rca24_fa173_y0 = f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_12_12_y0 ^ f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_11_13_y0;
  assign f_s_dadda_rca24_fa173_y1 = f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_12_12_y0 & f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_11_13_y0;
  assign f_s_dadda_rca24_fa173_y2 = f_s_dadda_rca24_fa173_y0 ^ f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_10_14_y0;
  assign f_s_dadda_rca24_fa173_y3 = f_s_dadda_rca24_fa173_y0 & f_s_dadda_rca24_fa173_f_s_dadda_rca24_and_10_14_y0;
  assign f_s_dadda_rca24_fa173_y4 = f_s_dadda_rca24_fa173_y1 | f_s_dadda_rca24_fa173_y3;
  assign f_s_dadda_rca24_and_9_15_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_9_15_y0 = f_s_dadda_rca24_and_9_15_a_9 & f_s_dadda_rca24_and_9_15_b_15;
  assign f_s_dadda_rca24_and_8_16_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_8_16_y0 = f_s_dadda_rca24_and_8_16_a_8 & f_s_dadda_rca24_and_8_16_b_16;
  assign f_s_dadda_rca24_and_7_17_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_7_17_y0 = f_s_dadda_rca24_and_7_17_a_7 & f_s_dadda_rca24_and_7_17_b_17;
  assign f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_9_15_y0 = f_s_dadda_rca24_and_9_15_y0;
  assign f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_8_16_y0 = f_s_dadda_rca24_and_8_16_y0;
  assign f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_7_17_y0 = f_s_dadda_rca24_and_7_17_y0;
  assign f_s_dadda_rca24_fa174_y0 = f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_9_15_y0 ^ f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_8_16_y0;
  assign f_s_dadda_rca24_fa174_y1 = f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_9_15_y0 & f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_8_16_y0;
  assign f_s_dadda_rca24_fa174_y2 = f_s_dadda_rca24_fa174_y0 ^ f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_7_17_y0;
  assign f_s_dadda_rca24_fa174_y3 = f_s_dadda_rca24_fa174_y0 & f_s_dadda_rca24_fa174_f_s_dadda_rca24_and_7_17_y0;
  assign f_s_dadda_rca24_fa174_y4 = f_s_dadda_rca24_fa174_y1 | f_s_dadda_rca24_fa174_y3;
  assign f_s_dadda_rca24_and_6_18_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_6_18_y0 = f_s_dadda_rca24_and_6_18_a_6 & f_s_dadda_rca24_and_6_18_b_18;
  assign f_s_dadda_rca24_and_5_19_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_5_19_y0 = f_s_dadda_rca24_and_5_19_a_5 & f_s_dadda_rca24_and_5_19_b_19;
  assign f_s_dadda_rca24_and_4_20_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_4_20_y0 = f_s_dadda_rca24_and_4_20_a_4 & f_s_dadda_rca24_and_4_20_b_20;
  assign f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_6_18_y0 = f_s_dadda_rca24_and_6_18_y0;
  assign f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_5_19_y0 = f_s_dadda_rca24_and_5_19_y0;
  assign f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_4_20_y0 = f_s_dadda_rca24_and_4_20_y0;
  assign f_s_dadda_rca24_fa175_y0 = f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_6_18_y0 ^ f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_5_19_y0;
  assign f_s_dadda_rca24_fa175_y1 = f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_6_18_y0 & f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_5_19_y0;
  assign f_s_dadda_rca24_fa175_y2 = f_s_dadda_rca24_fa175_y0 ^ f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_4_20_y0;
  assign f_s_dadda_rca24_fa175_y3 = f_s_dadda_rca24_fa175_y0 & f_s_dadda_rca24_fa175_f_s_dadda_rca24_and_4_20_y0;
  assign f_s_dadda_rca24_fa175_y4 = f_s_dadda_rca24_fa175_y1 | f_s_dadda_rca24_fa175_y3;
  assign f_s_dadda_rca24_and_3_21_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_3_21_y0 = f_s_dadda_rca24_and_3_21_a_3 & f_s_dadda_rca24_and_3_21_b_21;
  assign f_s_dadda_rca24_and_2_22_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_2_22_y0 = f_s_dadda_rca24_and_2_22_a_2 & f_s_dadda_rca24_and_2_22_b_22;
  assign f_s_dadda_rca24_nand_1_23_a_1 = a_1;
  assign f_s_dadda_rca24_nand_1_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_1_23_y0 = ~(f_s_dadda_rca24_nand_1_23_a_1 & f_s_dadda_rca24_nand_1_23_b_23);
  assign f_s_dadda_rca24_fa176_f_s_dadda_rca24_and_3_21_y0 = f_s_dadda_rca24_and_3_21_y0;
  assign f_s_dadda_rca24_fa176_f_s_dadda_rca24_and_2_22_y0 = f_s_dadda_rca24_and_2_22_y0;
  assign f_s_dadda_rca24_fa176_f_s_dadda_rca24_nand_1_23_y0 = f_s_dadda_rca24_nand_1_23_y0;
  assign f_s_dadda_rca24_fa176_y0 = f_s_dadda_rca24_fa176_f_s_dadda_rca24_and_3_21_y0 ^ f_s_dadda_rca24_fa176_f_s_dadda_rca24_and_2_22_y0;
  assign f_s_dadda_rca24_fa176_y1 = f_s_dadda_rca24_fa176_f_s_dadda_rca24_and_3_21_y0 & f_s_dadda_rca24_fa176_f_s_dadda_rca24_and_2_22_y0;
  assign f_s_dadda_rca24_fa176_y2 = f_s_dadda_rca24_fa176_y0 ^ f_s_dadda_rca24_fa176_f_s_dadda_rca24_nand_1_23_y0;
  assign f_s_dadda_rca24_fa176_y3 = f_s_dadda_rca24_fa176_y0 & f_s_dadda_rca24_fa176_f_s_dadda_rca24_nand_1_23_y0;
  assign f_s_dadda_rca24_fa176_y4 = f_s_dadda_rca24_fa176_y1 | f_s_dadda_rca24_fa176_y3;
  assign f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa10_y2 = f_s_dadda_rca24_fa10_y2;
  assign f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa11_y2 = f_s_dadda_rca24_fa11_y2;
  assign f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa12_y2 = f_s_dadda_rca24_fa12_y2;
  assign f_s_dadda_rca24_fa177_y0 = f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa10_y2 ^ f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa11_y2;
  assign f_s_dadda_rca24_fa177_y1 = f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa10_y2 & f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa11_y2;
  assign f_s_dadda_rca24_fa177_y2 = f_s_dadda_rca24_fa177_y0 ^ f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa12_y2;
  assign f_s_dadda_rca24_fa177_y3 = f_s_dadda_rca24_fa177_y0 & f_s_dadda_rca24_fa177_f_s_dadda_rca24_fa12_y2;
  assign f_s_dadda_rca24_fa177_y4 = f_s_dadda_rca24_fa177_y1 | f_s_dadda_rca24_fa177_y3;
  assign f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa13_y2 = f_s_dadda_rca24_fa13_y2;
  assign f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa14_y2 = f_s_dadda_rca24_fa14_y2;
  assign f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa168_y2 = f_s_dadda_rca24_fa168_y2;
  assign f_s_dadda_rca24_fa178_y0 = f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa13_y2 ^ f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa14_y2;
  assign f_s_dadda_rca24_fa178_y1 = f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa13_y2 & f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa14_y2;
  assign f_s_dadda_rca24_fa178_y2 = f_s_dadda_rca24_fa178_y0 ^ f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa168_y2;
  assign f_s_dadda_rca24_fa178_y3 = f_s_dadda_rca24_fa178_y0 & f_s_dadda_rca24_fa178_f_s_dadda_rca24_fa168_y2;
  assign f_s_dadda_rca24_fa178_y4 = f_s_dadda_rca24_fa178_y1 | f_s_dadda_rca24_fa178_y3;
  assign f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa169_y2 = f_s_dadda_rca24_fa169_y2;
  assign f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa170_y2 = f_s_dadda_rca24_fa170_y2;
  assign f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa171_y2 = f_s_dadda_rca24_fa171_y2;
  assign f_s_dadda_rca24_fa179_y0 = f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa169_y2 ^ f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa170_y2;
  assign f_s_dadda_rca24_fa179_y1 = f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa169_y2 & f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa170_y2;
  assign f_s_dadda_rca24_fa179_y2 = f_s_dadda_rca24_fa179_y0 ^ f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa171_y2;
  assign f_s_dadda_rca24_fa179_y3 = f_s_dadda_rca24_fa179_y0 & f_s_dadda_rca24_fa179_f_s_dadda_rca24_fa171_y2;
  assign f_s_dadda_rca24_fa179_y4 = f_s_dadda_rca24_fa179_y1 | f_s_dadda_rca24_fa179_y3;
  assign f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa172_y2 = f_s_dadda_rca24_fa172_y2;
  assign f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa173_y2 = f_s_dadda_rca24_fa173_y2;
  assign f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa174_y2 = f_s_dadda_rca24_fa174_y2;
  assign f_s_dadda_rca24_fa180_y0 = f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa172_y2 ^ f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa173_y2;
  assign f_s_dadda_rca24_fa180_y1 = f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa172_y2 & f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa173_y2;
  assign f_s_dadda_rca24_fa180_y2 = f_s_dadda_rca24_fa180_y0 ^ f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa174_y2;
  assign f_s_dadda_rca24_fa180_y3 = f_s_dadda_rca24_fa180_y0 & f_s_dadda_rca24_fa180_f_s_dadda_rca24_fa174_y2;
  assign f_s_dadda_rca24_fa180_y4 = f_s_dadda_rca24_fa180_y1 | f_s_dadda_rca24_fa180_y3;
  assign f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa180_y4 = f_s_dadda_rca24_fa180_y4;
  assign f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa179_y4 = f_s_dadda_rca24_fa179_y4;
  assign f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa178_y4 = f_s_dadda_rca24_fa178_y4;
  assign f_s_dadda_rca24_fa181_y0 = f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa180_y4 ^ f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa179_y4;
  assign f_s_dadda_rca24_fa181_y1 = f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa180_y4 & f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa179_y4;
  assign f_s_dadda_rca24_fa181_y2 = f_s_dadda_rca24_fa181_y0 ^ f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa178_y4;
  assign f_s_dadda_rca24_fa181_y3 = f_s_dadda_rca24_fa181_y0 & f_s_dadda_rca24_fa181_f_s_dadda_rca24_fa178_y4;
  assign f_s_dadda_rca24_fa181_y4 = f_s_dadda_rca24_fa181_y1 | f_s_dadda_rca24_fa181_y3;
  assign f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa177_y4 = f_s_dadda_rca24_fa177_y4;
  assign f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa176_y4 = f_s_dadda_rca24_fa176_y4;
  assign f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa175_y4 = f_s_dadda_rca24_fa175_y4;
  assign f_s_dadda_rca24_fa182_y0 = f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa177_y4 ^ f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa176_y4;
  assign f_s_dadda_rca24_fa182_y1 = f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa177_y4 & f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa176_y4;
  assign f_s_dadda_rca24_fa182_y2 = f_s_dadda_rca24_fa182_y0 ^ f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa175_y4;
  assign f_s_dadda_rca24_fa182_y3 = f_s_dadda_rca24_fa182_y0 & f_s_dadda_rca24_fa182_f_s_dadda_rca24_fa175_y4;
  assign f_s_dadda_rca24_fa182_y4 = f_s_dadda_rca24_fa182_y1 | f_s_dadda_rca24_fa182_y3;
  assign f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa174_y4 = f_s_dadda_rca24_fa174_y4;
  assign f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa173_y4 = f_s_dadda_rca24_fa173_y4;
  assign f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa172_y4 = f_s_dadda_rca24_fa172_y4;
  assign f_s_dadda_rca24_fa183_y0 = f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa174_y4 ^ f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa173_y4;
  assign f_s_dadda_rca24_fa183_y1 = f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa174_y4 & f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa173_y4;
  assign f_s_dadda_rca24_fa183_y2 = f_s_dadda_rca24_fa183_y0 ^ f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa172_y4;
  assign f_s_dadda_rca24_fa183_y3 = f_s_dadda_rca24_fa183_y0 & f_s_dadda_rca24_fa183_f_s_dadda_rca24_fa172_y4;
  assign f_s_dadda_rca24_fa183_y4 = f_s_dadda_rca24_fa183_y1 | f_s_dadda_rca24_fa183_y3;
  assign f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa171_y4 = f_s_dadda_rca24_fa171_y4;
  assign f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa170_y4 = f_s_dadda_rca24_fa170_y4;
  assign f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa169_y4 = f_s_dadda_rca24_fa169_y4;
  assign f_s_dadda_rca24_fa184_y0 = f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa171_y4 ^ f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa170_y4;
  assign f_s_dadda_rca24_fa184_y1 = f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa171_y4 & f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa170_y4;
  assign f_s_dadda_rca24_fa184_y2 = f_s_dadda_rca24_fa184_y0 ^ f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa169_y4;
  assign f_s_dadda_rca24_fa184_y3 = f_s_dadda_rca24_fa184_y0 & f_s_dadda_rca24_fa184_f_s_dadda_rca24_fa169_y4;
  assign f_s_dadda_rca24_fa184_y4 = f_s_dadda_rca24_fa184_y1 | f_s_dadda_rca24_fa184_y3;
  assign f_s_dadda_rca24_and_16_9_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_16_9_y0 = f_s_dadda_rca24_and_16_9_a_16 & f_s_dadda_rca24_and_16_9_b_9;
  assign f_s_dadda_rca24_and_15_10_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_15_10_y0 = f_s_dadda_rca24_and_15_10_a_15 & f_s_dadda_rca24_and_15_10_b_10;
  assign f_s_dadda_rca24_fa185_f_s_dadda_rca24_fa168_y4 = f_s_dadda_rca24_fa168_y4;
  assign f_s_dadda_rca24_fa185_f_s_dadda_rca24_and_16_9_y0 = f_s_dadda_rca24_and_16_9_y0;
  assign f_s_dadda_rca24_fa185_f_s_dadda_rca24_and_15_10_y0 = f_s_dadda_rca24_and_15_10_y0;
  assign f_s_dadda_rca24_fa185_y0 = f_s_dadda_rca24_fa185_f_s_dadda_rca24_fa168_y4 ^ f_s_dadda_rca24_fa185_f_s_dadda_rca24_and_16_9_y0;
  assign f_s_dadda_rca24_fa185_y1 = f_s_dadda_rca24_fa185_f_s_dadda_rca24_fa168_y4 & f_s_dadda_rca24_fa185_f_s_dadda_rca24_and_16_9_y0;
  assign f_s_dadda_rca24_fa185_y2 = f_s_dadda_rca24_fa185_y0 ^ f_s_dadda_rca24_fa185_f_s_dadda_rca24_and_15_10_y0;
  assign f_s_dadda_rca24_fa185_y3 = f_s_dadda_rca24_fa185_y0 & f_s_dadda_rca24_fa185_f_s_dadda_rca24_and_15_10_y0;
  assign f_s_dadda_rca24_fa185_y4 = f_s_dadda_rca24_fa185_y1 | f_s_dadda_rca24_fa185_y3;
  assign f_s_dadda_rca24_and_14_11_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_14_11_y0 = f_s_dadda_rca24_and_14_11_a_14 & f_s_dadda_rca24_and_14_11_b_11;
  assign f_s_dadda_rca24_and_13_12_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_13_12_y0 = f_s_dadda_rca24_and_13_12_a_13 & f_s_dadda_rca24_and_13_12_b_12;
  assign f_s_dadda_rca24_and_12_13_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_12_13_y0 = f_s_dadda_rca24_and_12_13_a_12 & f_s_dadda_rca24_and_12_13_b_13;
  assign f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_14_11_y0 = f_s_dadda_rca24_and_14_11_y0;
  assign f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_13_12_y0 = f_s_dadda_rca24_and_13_12_y0;
  assign f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_12_13_y0 = f_s_dadda_rca24_and_12_13_y0;
  assign f_s_dadda_rca24_fa186_y0 = f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_14_11_y0 ^ f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_13_12_y0;
  assign f_s_dadda_rca24_fa186_y1 = f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_14_11_y0 & f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_13_12_y0;
  assign f_s_dadda_rca24_fa186_y2 = f_s_dadda_rca24_fa186_y0 ^ f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_12_13_y0;
  assign f_s_dadda_rca24_fa186_y3 = f_s_dadda_rca24_fa186_y0 & f_s_dadda_rca24_fa186_f_s_dadda_rca24_and_12_13_y0;
  assign f_s_dadda_rca24_fa186_y4 = f_s_dadda_rca24_fa186_y1 | f_s_dadda_rca24_fa186_y3;
  assign f_s_dadda_rca24_and_11_14_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_11_14_y0 = f_s_dadda_rca24_and_11_14_a_11 & f_s_dadda_rca24_and_11_14_b_14;
  assign f_s_dadda_rca24_and_10_15_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_10_15_y0 = f_s_dadda_rca24_and_10_15_a_10 & f_s_dadda_rca24_and_10_15_b_15;
  assign f_s_dadda_rca24_and_9_16_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_9_16_y0 = f_s_dadda_rca24_and_9_16_a_9 & f_s_dadda_rca24_and_9_16_b_16;
  assign f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_11_14_y0 = f_s_dadda_rca24_and_11_14_y0;
  assign f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_10_15_y0 = f_s_dadda_rca24_and_10_15_y0;
  assign f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_9_16_y0 = f_s_dadda_rca24_and_9_16_y0;
  assign f_s_dadda_rca24_fa187_y0 = f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_11_14_y0 ^ f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_10_15_y0;
  assign f_s_dadda_rca24_fa187_y1 = f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_11_14_y0 & f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_10_15_y0;
  assign f_s_dadda_rca24_fa187_y2 = f_s_dadda_rca24_fa187_y0 ^ f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_9_16_y0;
  assign f_s_dadda_rca24_fa187_y3 = f_s_dadda_rca24_fa187_y0 & f_s_dadda_rca24_fa187_f_s_dadda_rca24_and_9_16_y0;
  assign f_s_dadda_rca24_fa187_y4 = f_s_dadda_rca24_fa187_y1 | f_s_dadda_rca24_fa187_y3;
  assign f_s_dadda_rca24_and_8_17_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_8_17_y0 = f_s_dadda_rca24_and_8_17_a_8 & f_s_dadda_rca24_and_8_17_b_17;
  assign f_s_dadda_rca24_and_7_18_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_7_18_y0 = f_s_dadda_rca24_and_7_18_a_7 & f_s_dadda_rca24_and_7_18_b_18;
  assign f_s_dadda_rca24_and_6_19_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_6_19_y0 = f_s_dadda_rca24_and_6_19_a_6 & f_s_dadda_rca24_and_6_19_b_19;
  assign f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_8_17_y0 = f_s_dadda_rca24_and_8_17_y0;
  assign f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_7_18_y0 = f_s_dadda_rca24_and_7_18_y0;
  assign f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_6_19_y0 = f_s_dadda_rca24_and_6_19_y0;
  assign f_s_dadda_rca24_fa188_y0 = f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_8_17_y0 ^ f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_7_18_y0;
  assign f_s_dadda_rca24_fa188_y1 = f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_8_17_y0 & f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_7_18_y0;
  assign f_s_dadda_rca24_fa188_y2 = f_s_dadda_rca24_fa188_y0 ^ f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_6_19_y0;
  assign f_s_dadda_rca24_fa188_y3 = f_s_dadda_rca24_fa188_y0 & f_s_dadda_rca24_fa188_f_s_dadda_rca24_and_6_19_y0;
  assign f_s_dadda_rca24_fa188_y4 = f_s_dadda_rca24_fa188_y1 | f_s_dadda_rca24_fa188_y3;
  assign f_s_dadda_rca24_and_5_20_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_5_20_y0 = f_s_dadda_rca24_and_5_20_a_5 & f_s_dadda_rca24_and_5_20_b_20;
  assign f_s_dadda_rca24_and_4_21_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_4_21_y0 = f_s_dadda_rca24_and_4_21_a_4 & f_s_dadda_rca24_and_4_21_b_21;
  assign f_s_dadda_rca24_and_3_22_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_3_22_y0 = f_s_dadda_rca24_and_3_22_a_3 & f_s_dadda_rca24_and_3_22_b_22;
  assign f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_5_20_y0 = f_s_dadda_rca24_and_5_20_y0;
  assign f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_4_21_y0 = f_s_dadda_rca24_and_4_21_y0;
  assign f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_3_22_y0 = f_s_dadda_rca24_and_3_22_y0;
  assign f_s_dadda_rca24_fa189_y0 = f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_5_20_y0 ^ f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_4_21_y0;
  assign f_s_dadda_rca24_fa189_y1 = f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_5_20_y0 & f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_4_21_y0;
  assign f_s_dadda_rca24_fa189_y2 = f_s_dadda_rca24_fa189_y0 ^ f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_3_22_y0;
  assign f_s_dadda_rca24_fa189_y3 = f_s_dadda_rca24_fa189_y0 & f_s_dadda_rca24_fa189_f_s_dadda_rca24_and_3_22_y0;
  assign f_s_dadda_rca24_fa189_y4 = f_s_dadda_rca24_fa189_y1 | f_s_dadda_rca24_fa189_y3;
  assign f_s_dadda_rca24_nand_2_23_a_2 = a_2;
  assign f_s_dadda_rca24_nand_2_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_2_23_y0 = ~(f_s_dadda_rca24_nand_2_23_a_2 & f_s_dadda_rca24_nand_2_23_b_23);
  assign f_s_dadda_rca24_fa190_f_s_dadda_rca24_nand_2_23_y0 = f_s_dadda_rca24_nand_2_23_y0;
  assign f_s_dadda_rca24_fa190_f_s_dadda_rca24_fa15_y2 = f_s_dadda_rca24_fa15_y2;
  assign f_s_dadda_rca24_fa190_f_s_dadda_rca24_fa16_y2 = f_s_dadda_rca24_fa16_y2;
  assign f_s_dadda_rca24_fa190_y0 = f_s_dadda_rca24_fa190_f_s_dadda_rca24_nand_2_23_y0 ^ f_s_dadda_rca24_fa190_f_s_dadda_rca24_fa15_y2;
  assign f_s_dadda_rca24_fa190_y1 = f_s_dadda_rca24_fa190_f_s_dadda_rca24_nand_2_23_y0 & f_s_dadda_rca24_fa190_f_s_dadda_rca24_fa15_y2;
  assign f_s_dadda_rca24_fa190_y2 = f_s_dadda_rca24_fa190_y0 ^ f_s_dadda_rca24_fa190_f_s_dadda_rca24_fa16_y2;
  assign f_s_dadda_rca24_fa190_y3 = f_s_dadda_rca24_fa190_y0 & f_s_dadda_rca24_fa190_f_s_dadda_rca24_fa16_y2;
  assign f_s_dadda_rca24_fa190_y4 = f_s_dadda_rca24_fa190_y1 | f_s_dadda_rca24_fa190_y3;
  assign f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa17_y2 = f_s_dadda_rca24_fa17_y2;
  assign f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa18_y2 = f_s_dadda_rca24_fa18_y2;
  assign f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa181_y2 = f_s_dadda_rca24_fa181_y2;
  assign f_s_dadda_rca24_fa191_y0 = f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa17_y2 ^ f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa18_y2;
  assign f_s_dadda_rca24_fa191_y1 = f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa17_y2 & f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa18_y2;
  assign f_s_dadda_rca24_fa191_y2 = f_s_dadda_rca24_fa191_y0 ^ f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa181_y2;
  assign f_s_dadda_rca24_fa191_y3 = f_s_dadda_rca24_fa191_y0 & f_s_dadda_rca24_fa191_f_s_dadda_rca24_fa181_y2;
  assign f_s_dadda_rca24_fa191_y4 = f_s_dadda_rca24_fa191_y1 | f_s_dadda_rca24_fa191_y3;
  assign f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa182_y2 = f_s_dadda_rca24_fa182_y2;
  assign f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa183_y2 = f_s_dadda_rca24_fa183_y2;
  assign f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa184_y2 = f_s_dadda_rca24_fa184_y2;
  assign f_s_dadda_rca24_fa192_y0 = f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa182_y2 ^ f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa183_y2;
  assign f_s_dadda_rca24_fa192_y1 = f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa182_y2 & f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa183_y2;
  assign f_s_dadda_rca24_fa192_y2 = f_s_dadda_rca24_fa192_y0 ^ f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa184_y2;
  assign f_s_dadda_rca24_fa192_y3 = f_s_dadda_rca24_fa192_y0 & f_s_dadda_rca24_fa192_f_s_dadda_rca24_fa184_y2;
  assign f_s_dadda_rca24_fa192_y4 = f_s_dadda_rca24_fa192_y1 | f_s_dadda_rca24_fa192_y3;
  assign f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa185_y2 = f_s_dadda_rca24_fa185_y2;
  assign f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa186_y2 = f_s_dadda_rca24_fa186_y2;
  assign f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa187_y2 = f_s_dadda_rca24_fa187_y2;
  assign f_s_dadda_rca24_fa193_y0 = f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa185_y2 ^ f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa186_y2;
  assign f_s_dadda_rca24_fa193_y1 = f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa185_y2 & f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa186_y2;
  assign f_s_dadda_rca24_fa193_y2 = f_s_dadda_rca24_fa193_y0 ^ f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa187_y2;
  assign f_s_dadda_rca24_fa193_y3 = f_s_dadda_rca24_fa193_y0 & f_s_dadda_rca24_fa193_f_s_dadda_rca24_fa187_y2;
  assign f_s_dadda_rca24_fa193_y4 = f_s_dadda_rca24_fa193_y1 | f_s_dadda_rca24_fa193_y3;
  assign f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa193_y4 = f_s_dadda_rca24_fa193_y4;
  assign f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa192_y4 = f_s_dadda_rca24_fa192_y4;
  assign f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa191_y4 = f_s_dadda_rca24_fa191_y4;
  assign f_s_dadda_rca24_fa194_y0 = f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa193_y4 ^ f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa192_y4;
  assign f_s_dadda_rca24_fa194_y1 = f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa193_y4 & f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa192_y4;
  assign f_s_dadda_rca24_fa194_y2 = f_s_dadda_rca24_fa194_y0 ^ f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa191_y4;
  assign f_s_dadda_rca24_fa194_y3 = f_s_dadda_rca24_fa194_y0 & f_s_dadda_rca24_fa194_f_s_dadda_rca24_fa191_y4;
  assign f_s_dadda_rca24_fa194_y4 = f_s_dadda_rca24_fa194_y1 | f_s_dadda_rca24_fa194_y3;
  assign f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa190_y4 = f_s_dadda_rca24_fa190_y4;
  assign f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa189_y4 = f_s_dadda_rca24_fa189_y4;
  assign f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa188_y4 = f_s_dadda_rca24_fa188_y4;
  assign f_s_dadda_rca24_fa195_y0 = f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa190_y4 ^ f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa189_y4;
  assign f_s_dadda_rca24_fa195_y1 = f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa190_y4 & f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa189_y4;
  assign f_s_dadda_rca24_fa195_y2 = f_s_dadda_rca24_fa195_y0 ^ f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa188_y4;
  assign f_s_dadda_rca24_fa195_y3 = f_s_dadda_rca24_fa195_y0 & f_s_dadda_rca24_fa195_f_s_dadda_rca24_fa188_y4;
  assign f_s_dadda_rca24_fa195_y4 = f_s_dadda_rca24_fa195_y1 | f_s_dadda_rca24_fa195_y3;
  assign f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa187_y4 = f_s_dadda_rca24_fa187_y4;
  assign f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa186_y4 = f_s_dadda_rca24_fa186_y4;
  assign f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa185_y4 = f_s_dadda_rca24_fa185_y4;
  assign f_s_dadda_rca24_fa196_y0 = f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa187_y4 ^ f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa186_y4;
  assign f_s_dadda_rca24_fa196_y1 = f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa187_y4 & f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa186_y4;
  assign f_s_dadda_rca24_fa196_y2 = f_s_dadda_rca24_fa196_y0 ^ f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa185_y4;
  assign f_s_dadda_rca24_fa196_y3 = f_s_dadda_rca24_fa196_y0 & f_s_dadda_rca24_fa196_f_s_dadda_rca24_fa185_y4;
  assign f_s_dadda_rca24_fa196_y4 = f_s_dadda_rca24_fa196_y1 | f_s_dadda_rca24_fa196_y3;
  assign f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa184_y4 = f_s_dadda_rca24_fa184_y4;
  assign f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa183_y4 = f_s_dadda_rca24_fa183_y4;
  assign f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa182_y4 = f_s_dadda_rca24_fa182_y4;
  assign f_s_dadda_rca24_fa197_y0 = f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa184_y4 ^ f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa183_y4;
  assign f_s_dadda_rca24_fa197_y1 = f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa184_y4 & f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa183_y4;
  assign f_s_dadda_rca24_fa197_y2 = f_s_dadda_rca24_fa197_y0 ^ f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa182_y4;
  assign f_s_dadda_rca24_fa197_y3 = f_s_dadda_rca24_fa197_y0 & f_s_dadda_rca24_fa197_f_s_dadda_rca24_fa182_y4;
  assign f_s_dadda_rca24_fa197_y4 = f_s_dadda_rca24_fa197_y1 | f_s_dadda_rca24_fa197_y3;
  assign f_s_dadda_rca24_and_18_8_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_18_8_y0 = f_s_dadda_rca24_and_18_8_a_18 & f_s_dadda_rca24_and_18_8_b_8;
  assign f_s_dadda_rca24_and_17_9_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_17_9_y0 = f_s_dadda_rca24_and_17_9_a_17 & f_s_dadda_rca24_and_17_9_b_9;
  assign f_s_dadda_rca24_fa198_f_s_dadda_rca24_fa181_y4 = f_s_dadda_rca24_fa181_y4;
  assign f_s_dadda_rca24_fa198_f_s_dadda_rca24_and_18_8_y0 = f_s_dadda_rca24_and_18_8_y0;
  assign f_s_dadda_rca24_fa198_f_s_dadda_rca24_and_17_9_y0 = f_s_dadda_rca24_and_17_9_y0;
  assign f_s_dadda_rca24_fa198_y0 = f_s_dadda_rca24_fa198_f_s_dadda_rca24_fa181_y4 ^ f_s_dadda_rca24_fa198_f_s_dadda_rca24_and_18_8_y0;
  assign f_s_dadda_rca24_fa198_y1 = f_s_dadda_rca24_fa198_f_s_dadda_rca24_fa181_y4 & f_s_dadda_rca24_fa198_f_s_dadda_rca24_and_18_8_y0;
  assign f_s_dadda_rca24_fa198_y2 = f_s_dadda_rca24_fa198_y0 ^ f_s_dadda_rca24_fa198_f_s_dadda_rca24_and_17_9_y0;
  assign f_s_dadda_rca24_fa198_y3 = f_s_dadda_rca24_fa198_y0 & f_s_dadda_rca24_fa198_f_s_dadda_rca24_and_17_9_y0;
  assign f_s_dadda_rca24_fa198_y4 = f_s_dadda_rca24_fa198_y1 | f_s_dadda_rca24_fa198_y3;
  assign f_s_dadda_rca24_and_16_10_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_16_10_y0 = f_s_dadda_rca24_and_16_10_a_16 & f_s_dadda_rca24_and_16_10_b_10;
  assign f_s_dadda_rca24_and_15_11_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_15_11_y0 = f_s_dadda_rca24_and_15_11_a_15 & f_s_dadda_rca24_and_15_11_b_11;
  assign f_s_dadda_rca24_and_14_12_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_14_12_y0 = f_s_dadda_rca24_and_14_12_a_14 & f_s_dadda_rca24_and_14_12_b_12;
  assign f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_16_10_y0 = f_s_dadda_rca24_and_16_10_y0;
  assign f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_15_11_y0 = f_s_dadda_rca24_and_15_11_y0;
  assign f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_14_12_y0 = f_s_dadda_rca24_and_14_12_y0;
  assign f_s_dadda_rca24_fa199_y0 = f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_16_10_y0 ^ f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_15_11_y0;
  assign f_s_dadda_rca24_fa199_y1 = f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_16_10_y0 & f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_15_11_y0;
  assign f_s_dadda_rca24_fa199_y2 = f_s_dadda_rca24_fa199_y0 ^ f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_14_12_y0;
  assign f_s_dadda_rca24_fa199_y3 = f_s_dadda_rca24_fa199_y0 & f_s_dadda_rca24_fa199_f_s_dadda_rca24_and_14_12_y0;
  assign f_s_dadda_rca24_fa199_y4 = f_s_dadda_rca24_fa199_y1 | f_s_dadda_rca24_fa199_y3;
  assign f_s_dadda_rca24_and_13_13_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_13_13_y0 = f_s_dadda_rca24_and_13_13_a_13 & f_s_dadda_rca24_and_13_13_b_13;
  assign f_s_dadda_rca24_and_12_14_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_12_14_y0 = f_s_dadda_rca24_and_12_14_a_12 & f_s_dadda_rca24_and_12_14_b_14;
  assign f_s_dadda_rca24_and_11_15_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_11_15_y0 = f_s_dadda_rca24_and_11_15_a_11 & f_s_dadda_rca24_and_11_15_b_15;
  assign f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_13_13_y0 = f_s_dadda_rca24_and_13_13_y0;
  assign f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_12_14_y0 = f_s_dadda_rca24_and_12_14_y0;
  assign f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_11_15_y0 = f_s_dadda_rca24_and_11_15_y0;
  assign f_s_dadda_rca24_fa200_y0 = f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_13_13_y0 ^ f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_12_14_y0;
  assign f_s_dadda_rca24_fa200_y1 = f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_13_13_y0 & f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_12_14_y0;
  assign f_s_dadda_rca24_fa200_y2 = f_s_dadda_rca24_fa200_y0 ^ f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_11_15_y0;
  assign f_s_dadda_rca24_fa200_y3 = f_s_dadda_rca24_fa200_y0 & f_s_dadda_rca24_fa200_f_s_dadda_rca24_and_11_15_y0;
  assign f_s_dadda_rca24_fa200_y4 = f_s_dadda_rca24_fa200_y1 | f_s_dadda_rca24_fa200_y3;
  assign f_s_dadda_rca24_and_10_16_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_10_16_y0 = f_s_dadda_rca24_and_10_16_a_10 & f_s_dadda_rca24_and_10_16_b_16;
  assign f_s_dadda_rca24_and_9_17_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_9_17_y0 = f_s_dadda_rca24_and_9_17_a_9 & f_s_dadda_rca24_and_9_17_b_17;
  assign f_s_dadda_rca24_and_8_18_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_8_18_y0 = f_s_dadda_rca24_and_8_18_a_8 & f_s_dadda_rca24_and_8_18_b_18;
  assign f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_10_16_y0 = f_s_dadda_rca24_and_10_16_y0;
  assign f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_9_17_y0 = f_s_dadda_rca24_and_9_17_y0;
  assign f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_8_18_y0 = f_s_dadda_rca24_and_8_18_y0;
  assign f_s_dadda_rca24_fa201_y0 = f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_10_16_y0 ^ f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_9_17_y0;
  assign f_s_dadda_rca24_fa201_y1 = f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_10_16_y0 & f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_9_17_y0;
  assign f_s_dadda_rca24_fa201_y2 = f_s_dadda_rca24_fa201_y0 ^ f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_8_18_y0;
  assign f_s_dadda_rca24_fa201_y3 = f_s_dadda_rca24_fa201_y0 & f_s_dadda_rca24_fa201_f_s_dadda_rca24_and_8_18_y0;
  assign f_s_dadda_rca24_fa201_y4 = f_s_dadda_rca24_fa201_y1 | f_s_dadda_rca24_fa201_y3;
  assign f_s_dadda_rca24_and_7_19_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_7_19_y0 = f_s_dadda_rca24_and_7_19_a_7 & f_s_dadda_rca24_and_7_19_b_19;
  assign f_s_dadda_rca24_and_6_20_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_6_20_y0 = f_s_dadda_rca24_and_6_20_a_6 & f_s_dadda_rca24_and_6_20_b_20;
  assign f_s_dadda_rca24_and_5_21_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_5_21_y0 = f_s_dadda_rca24_and_5_21_a_5 & f_s_dadda_rca24_and_5_21_b_21;
  assign f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_7_19_y0 = f_s_dadda_rca24_and_7_19_y0;
  assign f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_6_20_y0 = f_s_dadda_rca24_and_6_20_y0;
  assign f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_5_21_y0 = f_s_dadda_rca24_and_5_21_y0;
  assign f_s_dadda_rca24_fa202_y0 = f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_7_19_y0 ^ f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_6_20_y0;
  assign f_s_dadda_rca24_fa202_y1 = f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_7_19_y0 & f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_6_20_y0;
  assign f_s_dadda_rca24_fa202_y2 = f_s_dadda_rca24_fa202_y0 ^ f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_5_21_y0;
  assign f_s_dadda_rca24_fa202_y3 = f_s_dadda_rca24_fa202_y0 & f_s_dadda_rca24_fa202_f_s_dadda_rca24_and_5_21_y0;
  assign f_s_dadda_rca24_fa202_y4 = f_s_dadda_rca24_fa202_y1 | f_s_dadda_rca24_fa202_y3;
  assign f_s_dadda_rca24_and_4_22_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_4_22_y0 = f_s_dadda_rca24_and_4_22_a_4 & f_s_dadda_rca24_and_4_22_b_22;
  assign f_s_dadda_rca24_nand_3_23_a_3 = a_3;
  assign f_s_dadda_rca24_nand_3_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_3_23_y0 = ~(f_s_dadda_rca24_nand_3_23_a_3 & f_s_dadda_rca24_nand_3_23_b_23);
  assign f_s_dadda_rca24_fa203_f_s_dadda_rca24_and_4_22_y0 = f_s_dadda_rca24_and_4_22_y0;
  assign f_s_dadda_rca24_fa203_f_s_dadda_rca24_nand_3_23_y0 = f_s_dadda_rca24_nand_3_23_y0;
  assign f_s_dadda_rca24_fa203_f_s_dadda_rca24_fa19_y2 = f_s_dadda_rca24_fa19_y2;
  assign f_s_dadda_rca24_fa203_y0 = f_s_dadda_rca24_fa203_f_s_dadda_rca24_and_4_22_y0 ^ f_s_dadda_rca24_fa203_f_s_dadda_rca24_nand_3_23_y0;
  assign f_s_dadda_rca24_fa203_y1 = f_s_dadda_rca24_fa203_f_s_dadda_rca24_and_4_22_y0 & f_s_dadda_rca24_fa203_f_s_dadda_rca24_nand_3_23_y0;
  assign f_s_dadda_rca24_fa203_y2 = f_s_dadda_rca24_fa203_y0 ^ f_s_dadda_rca24_fa203_f_s_dadda_rca24_fa19_y2;
  assign f_s_dadda_rca24_fa203_y3 = f_s_dadda_rca24_fa203_y0 & f_s_dadda_rca24_fa203_f_s_dadda_rca24_fa19_y2;
  assign f_s_dadda_rca24_fa203_y4 = f_s_dadda_rca24_fa203_y1 | f_s_dadda_rca24_fa203_y3;
  assign f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa20_y2 = f_s_dadda_rca24_fa20_y2;
  assign f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa21_y2 = f_s_dadda_rca24_fa21_y2;
  assign f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa194_y2 = f_s_dadda_rca24_fa194_y2;
  assign f_s_dadda_rca24_fa204_y0 = f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa20_y2 ^ f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa21_y2;
  assign f_s_dadda_rca24_fa204_y1 = f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa20_y2 & f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa21_y2;
  assign f_s_dadda_rca24_fa204_y2 = f_s_dadda_rca24_fa204_y0 ^ f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa194_y2;
  assign f_s_dadda_rca24_fa204_y3 = f_s_dadda_rca24_fa204_y0 & f_s_dadda_rca24_fa204_f_s_dadda_rca24_fa194_y2;
  assign f_s_dadda_rca24_fa204_y4 = f_s_dadda_rca24_fa204_y1 | f_s_dadda_rca24_fa204_y3;
  assign f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa195_y2 = f_s_dadda_rca24_fa195_y2;
  assign f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa196_y2 = f_s_dadda_rca24_fa196_y2;
  assign f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa197_y2 = f_s_dadda_rca24_fa197_y2;
  assign f_s_dadda_rca24_fa205_y0 = f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa195_y2 ^ f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa196_y2;
  assign f_s_dadda_rca24_fa205_y1 = f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa195_y2 & f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa196_y2;
  assign f_s_dadda_rca24_fa205_y2 = f_s_dadda_rca24_fa205_y0 ^ f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa197_y2;
  assign f_s_dadda_rca24_fa205_y3 = f_s_dadda_rca24_fa205_y0 & f_s_dadda_rca24_fa205_f_s_dadda_rca24_fa197_y2;
  assign f_s_dadda_rca24_fa205_y4 = f_s_dadda_rca24_fa205_y1 | f_s_dadda_rca24_fa205_y3;
  assign f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa198_y2 = f_s_dadda_rca24_fa198_y2;
  assign f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa199_y2 = f_s_dadda_rca24_fa199_y2;
  assign f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa200_y2 = f_s_dadda_rca24_fa200_y2;
  assign f_s_dadda_rca24_fa206_y0 = f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa198_y2 ^ f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa199_y2;
  assign f_s_dadda_rca24_fa206_y1 = f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa198_y2 & f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa199_y2;
  assign f_s_dadda_rca24_fa206_y2 = f_s_dadda_rca24_fa206_y0 ^ f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa200_y2;
  assign f_s_dadda_rca24_fa206_y3 = f_s_dadda_rca24_fa206_y0 & f_s_dadda_rca24_fa206_f_s_dadda_rca24_fa200_y2;
  assign f_s_dadda_rca24_fa206_y4 = f_s_dadda_rca24_fa206_y1 | f_s_dadda_rca24_fa206_y3;
  assign f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa206_y4 = f_s_dadda_rca24_fa206_y4;
  assign f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa205_y4 = f_s_dadda_rca24_fa205_y4;
  assign f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa204_y4 = f_s_dadda_rca24_fa204_y4;
  assign f_s_dadda_rca24_fa207_y0 = f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa206_y4 ^ f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa205_y4;
  assign f_s_dadda_rca24_fa207_y1 = f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa206_y4 & f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa205_y4;
  assign f_s_dadda_rca24_fa207_y2 = f_s_dadda_rca24_fa207_y0 ^ f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa204_y4;
  assign f_s_dadda_rca24_fa207_y3 = f_s_dadda_rca24_fa207_y0 & f_s_dadda_rca24_fa207_f_s_dadda_rca24_fa204_y4;
  assign f_s_dadda_rca24_fa207_y4 = f_s_dadda_rca24_fa207_y1 | f_s_dadda_rca24_fa207_y3;
  assign f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa203_y4 = f_s_dadda_rca24_fa203_y4;
  assign f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa202_y4 = f_s_dadda_rca24_fa202_y4;
  assign f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa201_y4 = f_s_dadda_rca24_fa201_y4;
  assign f_s_dadda_rca24_fa208_y0 = f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa203_y4 ^ f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa202_y4;
  assign f_s_dadda_rca24_fa208_y1 = f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa203_y4 & f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa202_y4;
  assign f_s_dadda_rca24_fa208_y2 = f_s_dadda_rca24_fa208_y0 ^ f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa201_y4;
  assign f_s_dadda_rca24_fa208_y3 = f_s_dadda_rca24_fa208_y0 & f_s_dadda_rca24_fa208_f_s_dadda_rca24_fa201_y4;
  assign f_s_dadda_rca24_fa208_y4 = f_s_dadda_rca24_fa208_y1 | f_s_dadda_rca24_fa208_y3;
  assign f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa200_y4 = f_s_dadda_rca24_fa200_y4;
  assign f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa199_y4 = f_s_dadda_rca24_fa199_y4;
  assign f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa198_y4 = f_s_dadda_rca24_fa198_y4;
  assign f_s_dadda_rca24_fa209_y0 = f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa200_y4 ^ f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa199_y4;
  assign f_s_dadda_rca24_fa209_y1 = f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa200_y4 & f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa199_y4;
  assign f_s_dadda_rca24_fa209_y2 = f_s_dadda_rca24_fa209_y0 ^ f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa198_y4;
  assign f_s_dadda_rca24_fa209_y3 = f_s_dadda_rca24_fa209_y0 & f_s_dadda_rca24_fa209_f_s_dadda_rca24_fa198_y4;
  assign f_s_dadda_rca24_fa209_y4 = f_s_dadda_rca24_fa209_y1 | f_s_dadda_rca24_fa209_y3;
  assign f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa197_y4 = f_s_dadda_rca24_fa197_y4;
  assign f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa196_y4 = f_s_dadda_rca24_fa196_y4;
  assign f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa195_y4 = f_s_dadda_rca24_fa195_y4;
  assign f_s_dadda_rca24_fa210_y0 = f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa197_y4 ^ f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa196_y4;
  assign f_s_dadda_rca24_fa210_y1 = f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa197_y4 & f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa196_y4;
  assign f_s_dadda_rca24_fa210_y2 = f_s_dadda_rca24_fa210_y0 ^ f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa195_y4;
  assign f_s_dadda_rca24_fa210_y3 = f_s_dadda_rca24_fa210_y0 & f_s_dadda_rca24_fa210_f_s_dadda_rca24_fa195_y4;
  assign f_s_dadda_rca24_fa210_y4 = f_s_dadda_rca24_fa210_y1 | f_s_dadda_rca24_fa210_y3;
  assign f_s_dadda_rca24_and_20_7_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_20_7_y0 = f_s_dadda_rca24_and_20_7_a_20 & f_s_dadda_rca24_and_20_7_b_7;
  assign f_s_dadda_rca24_and_19_8_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_19_8_y0 = f_s_dadda_rca24_and_19_8_a_19 & f_s_dadda_rca24_and_19_8_b_8;
  assign f_s_dadda_rca24_fa211_f_s_dadda_rca24_fa194_y4 = f_s_dadda_rca24_fa194_y4;
  assign f_s_dadda_rca24_fa211_f_s_dadda_rca24_and_20_7_y0 = f_s_dadda_rca24_and_20_7_y0;
  assign f_s_dadda_rca24_fa211_f_s_dadda_rca24_and_19_8_y0 = f_s_dadda_rca24_and_19_8_y0;
  assign f_s_dadda_rca24_fa211_y0 = f_s_dadda_rca24_fa211_f_s_dadda_rca24_fa194_y4 ^ f_s_dadda_rca24_fa211_f_s_dadda_rca24_and_20_7_y0;
  assign f_s_dadda_rca24_fa211_y1 = f_s_dadda_rca24_fa211_f_s_dadda_rca24_fa194_y4 & f_s_dadda_rca24_fa211_f_s_dadda_rca24_and_20_7_y0;
  assign f_s_dadda_rca24_fa211_y2 = f_s_dadda_rca24_fa211_y0 ^ f_s_dadda_rca24_fa211_f_s_dadda_rca24_and_19_8_y0;
  assign f_s_dadda_rca24_fa211_y3 = f_s_dadda_rca24_fa211_y0 & f_s_dadda_rca24_fa211_f_s_dadda_rca24_and_19_8_y0;
  assign f_s_dadda_rca24_fa211_y4 = f_s_dadda_rca24_fa211_y1 | f_s_dadda_rca24_fa211_y3;
  assign f_s_dadda_rca24_and_18_9_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_18_9_y0 = f_s_dadda_rca24_and_18_9_a_18 & f_s_dadda_rca24_and_18_9_b_9;
  assign f_s_dadda_rca24_and_17_10_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_17_10_y0 = f_s_dadda_rca24_and_17_10_a_17 & f_s_dadda_rca24_and_17_10_b_10;
  assign f_s_dadda_rca24_and_16_11_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_16_11_y0 = f_s_dadda_rca24_and_16_11_a_16 & f_s_dadda_rca24_and_16_11_b_11;
  assign f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_18_9_y0 = f_s_dadda_rca24_and_18_9_y0;
  assign f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_17_10_y0 = f_s_dadda_rca24_and_17_10_y0;
  assign f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_16_11_y0 = f_s_dadda_rca24_and_16_11_y0;
  assign f_s_dadda_rca24_fa212_y0 = f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_18_9_y0 ^ f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_17_10_y0;
  assign f_s_dadda_rca24_fa212_y1 = f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_18_9_y0 & f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_17_10_y0;
  assign f_s_dadda_rca24_fa212_y2 = f_s_dadda_rca24_fa212_y0 ^ f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_16_11_y0;
  assign f_s_dadda_rca24_fa212_y3 = f_s_dadda_rca24_fa212_y0 & f_s_dadda_rca24_fa212_f_s_dadda_rca24_and_16_11_y0;
  assign f_s_dadda_rca24_fa212_y4 = f_s_dadda_rca24_fa212_y1 | f_s_dadda_rca24_fa212_y3;
  assign f_s_dadda_rca24_and_15_12_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_15_12_y0 = f_s_dadda_rca24_and_15_12_a_15 & f_s_dadda_rca24_and_15_12_b_12;
  assign f_s_dadda_rca24_and_14_13_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_14_13_y0 = f_s_dadda_rca24_and_14_13_a_14 & f_s_dadda_rca24_and_14_13_b_13;
  assign f_s_dadda_rca24_and_13_14_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_13_14_y0 = f_s_dadda_rca24_and_13_14_a_13 & f_s_dadda_rca24_and_13_14_b_14;
  assign f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_15_12_y0 = f_s_dadda_rca24_and_15_12_y0;
  assign f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_14_13_y0 = f_s_dadda_rca24_and_14_13_y0;
  assign f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_13_14_y0 = f_s_dadda_rca24_and_13_14_y0;
  assign f_s_dadda_rca24_fa213_y0 = f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_15_12_y0 ^ f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_14_13_y0;
  assign f_s_dadda_rca24_fa213_y1 = f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_15_12_y0 & f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_14_13_y0;
  assign f_s_dadda_rca24_fa213_y2 = f_s_dadda_rca24_fa213_y0 ^ f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_13_14_y0;
  assign f_s_dadda_rca24_fa213_y3 = f_s_dadda_rca24_fa213_y0 & f_s_dadda_rca24_fa213_f_s_dadda_rca24_and_13_14_y0;
  assign f_s_dadda_rca24_fa213_y4 = f_s_dadda_rca24_fa213_y1 | f_s_dadda_rca24_fa213_y3;
  assign f_s_dadda_rca24_and_12_15_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_12_15_y0 = f_s_dadda_rca24_and_12_15_a_12 & f_s_dadda_rca24_and_12_15_b_15;
  assign f_s_dadda_rca24_and_11_16_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_11_16_y0 = f_s_dadda_rca24_and_11_16_a_11 & f_s_dadda_rca24_and_11_16_b_16;
  assign f_s_dadda_rca24_and_10_17_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_10_17_y0 = f_s_dadda_rca24_and_10_17_a_10 & f_s_dadda_rca24_and_10_17_b_17;
  assign f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_12_15_y0 = f_s_dadda_rca24_and_12_15_y0;
  assign f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_11_16_y0 = f_s_dadda_rca24_and_11_16_y0;
  assign f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_10_17_y0 = f_s_dadda_rca24_and_10_17_y0;
  assign f_s_dadda_rca24_fa214_y0 = f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_12_15_y0 ^ f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_11_16_y0;
  assign f_s_dadda_rca24_fa214_y1 = f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_12_15_y0 & f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_11_16_y0;
  assign f_s_dadda_rca24_fa214_y2 = f_s_dadda_rca24_fa214_y0 ^ f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_10_17_y0;
  assign f_s_dadda_rca24_fa214_y3 = f_s_dadda_rca24_fa214_y0 & f_s_dadda_rca24_fa214_f_s_dadda_rca24_and_10_17_y0;
  assign f_s_dadda_rca24_fa214_y4 = f_s_dadda_rca24_fa214_y1 | f_s_dadda_rca24_fa214_y3;
  assign f_s_dadda_rca24_and_9_18_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_9_18_y0 = f_s_dadda_rca24_and_9_18_a_9 & f_s_dadda_rca24_and_9_18_b_18;
  assign f_s_dadda_rca24_and_8_19_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_8_19_y0 = f_s_dadda_rca24_and_8_19_a_8 & f_s_dadda_rca24_and_8_19_b_19;
  assign f_s_dadda_rca24_and_7_20_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_7_20_y0 = f_s_dadda_rca24_and_7_20_a_7 & f_s_dadda_rca24_and_7_20_b_20;
  assign f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_9_18_y0 = f_s_dadda_rca24_and_9_18_y0;
  assign f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_8_19_y0 = f_s_dadda_rca24_and_8_19_y0;
  assign f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_7_20_y0 = f_s_dadda_rca24_and_7_20_y0;
  assign f_s_dadda_rca24_fa215_y0 = f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_9_18_y0 ^ f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_8_19_y0;
  assign f_s_dadda_rca24_fa215_y1 = f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_9_18_y0 & f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_8_19_y0;
  assign f_s_dadda_rca24_fa215_y2 = f_s_dadda_rca24_fa215_y0 ^ f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_7_20_y0;
  assign f_s_dadda_rca24_fa215_y3 = f_s_dadda_rca24_fa215_y0 & f_s_dadda_rca24_fa215_f_s_dadda_rca24_and_7_20_y0;
  assign f_s_dadda_rca24_fa215_y4 = f_s_dadda_rca24_fa215_y1 | f_s_dadda_rca24_fa215_y3;
  assign f_s_dadda_rca24_and_6_21_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_6_21_y0 = f_s_dadda_rca24_and_6_21_a_6 & f_s_dadda_rca24_and_6_21_b_21;
  assign f_s_dadda_rca24_and_5_22_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_5_22_y0 = f_s_dadda_rca24_and_5_22_a_5 & f_s_dadda_rca24_and_5_22_b_22;
  assign f_s_dadda_rca24_nand_4_23_a_4 = a_4;
  assign f_s_dadda_rca24_nand_4_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_4_23_y0 = ~(f_s_dadda_rca24_nand_4_23_a_4 & f_s_dadda_rca24_nand_4_23_b_23);
  assign f_s_dadda_rca24_fa216_f_s_dadda_rca24_and_6_21_y0 = f_s_dadda_rca24_and_6_21_y0;
  assign f_s_dadda_rca24_fa216_f_s_dadda_rca24_and_5_22_y0 = f_s_dadda_rca24_and_5_22_y0;
  assign f_s_dadda_rca24_fa216_f_s_dadda_rca24_nand_4_23_y0 = f_s_dadda_rca24_nand_4_23_y0;
  assign f_s_dadda_rca24_fa216_y0 = f_s_dadda_rca24_fa216_f_s_dadda_rca24_and_6_21_y0 ^ f_s_dadda_rca24_fa216_f_s_dadda_rca24_and_5_22_y0;
  assign f_s_dadda_rca24_fa216_y1 = f_s_dadda_rca24_fa216_f_s_dadda_rca24_and_6_21_y0 & f_s_dadda_rca24_fa216_f_s_dadda_rca24_and_5_22_y0;
  assign f_s_dadda_rca24_fa216_y2 = f_s_dadda_rca24_fa216_y0 ^ f_s_dadda_rca24_fa216_f_s_dadda_rca24_nand_4_23_y0;
  assign f_s_dadda_rca24_fa216_y3 = f_s_dadda_rca24_fa216_y0 & f_s_dadda_rca24_fa216_f_s_dadda_rca24_nand_4_23_y0;
  assign f_s_dadda_rca24_fa216_y4 = f_s_dadda_rca24_fa216_y1 | f_s_dadda_rca24_fa216_y3;
  assign f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa22_y2 = f_s_dadda_rca24_fa22_y2;
  assign f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa23_y2 = f_s_dadda_rca24_fa23_y2;
  assign f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa207_y2 = f_s_dadda_rca24_fa207_y2;
  assign f_s_dadda_rca24_fa217_y0 = f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa22_y2 ^ f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa23_y2;
  assign f_s_dadda_rca24_fa217_y1 = f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa22_y2 & f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa23_y2;
  assign f_s_dadda_rca24_fa217_y2 = f_s_dadda_rca24_fa217_y0 ^ f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa207_y2;
  assign f_s_dadda_rca24_fa217_y3 = f_s_dadda_rca24_fa217_y0 & f_s_dadda_rca24_fa217_f_s_dadda_rca24_fa207_y2;
  assign f_s_dadda_rca24_fa217_y4 = f_s_dadda_rca24_fa217_y1 | f_s_dadda_rca24_fa217_y3;
  assign f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa208_y2 = f_s_dadda_rca24_fa208_y2;
  assign f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa209_y2 = f_s_dadda_rca24_fa209_y2;
  assign f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa210_y2 = f_s_dadda_rca24_fa210_y2;
  assign f_s_dadda_rca24_fa218_y0 = f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa208_y2 ^ f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa209_y2;
  assign f_s_dadda_rca24_fa218_y1 = f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa208_y2 & f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa209_y2;
  assign f_s_dadda_rca24_fa218_y2 = f_s_dadda_rca24_fa218_y0 ^ f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa210_y2;
  assign f_s_dadda_rca24_fa218_y3 = f_s_dadda_rca24_fa218_y0 & f_s_dadda_rca24_fa218_f_s_dadda_rca24_fa210_y2;
  assign f_s_dadda_rca24_fa218_y4 = f_s_dadda_rca24_fa218_y1 | f_s_dadda_rca24_fa218_y3;
  assign f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa211_y2 = f_s_dadda_rca24_fa211_y2;
  assign f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa212_y2 = f_s_dadda_rca24_fa212_y2;
  assign f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa213_y2 = f_s_dadda_rca24_fa213_y2;
  assign f_s_dadda_rca24_fa219_y0 = f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa211_y2 ^ f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa212_y2;
  assign f_s_dadda_rca24_fa219_y1 = f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa211_y2 & f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa212_y2;
  assign f_s_dadda_rca24_fa219_y2 = f_s_dadda_rca24_fa219_y0 ^ f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa213_y2;
  assign f_s_dadda_rca24_fa219_y3 = f_s_dadda_rca24_fa219_y0 & f_s_dadda_rca24_fa219_f_s_dadda_rca24_fa213_y2;
  assign f_s_dadda_rca24_fa219_y4 = f_s_dadda_rca24_fa219_y1 | f_s_dadda_rca24_fa219_y3;
  assign f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa219_y4 = f_s_dadda_rca24_fa219_y4;
  assign f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa218_y4 = f_s_dadda_rca24_fa218_y4;
  assign f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa217_y4 = f_s_dadda_rca24_fa217_y4;
  assign f_s_dadda_rca24_fa220_y0 = f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa219_y4 ^ f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa218_y4;
  assign f_s_dadda_rca24_fa220_y1 = f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa219_y4 & f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa218_y4;
  assign f_s_dadda_rca24_fa220_y2 = f_s_dadda_rca24_fa220_y0 ^ f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa217_y4;
  assign f_s_dadda_rca24_fa220_y3 = f_s_dadda_rca24_fa220_y0 & f_s_dadda_rca24_fa220_f_s_dadda_rca24_fa217_y4;
  assign f_s_dadda_rca24_fa220_y4 = f_s_dadda_rca24_fa220_y1 | f_s_dadda_rca24_fa220_y3;
  assign f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa216_y4 = f_s_dadda_rca24_fa216_y4;
  assign f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa215_y4 = f_s_dadda_rca24_fa215_y4;
  assign f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa214_y4 = f_s_dadda_rca24_fa214_y4;
  assign f_s_dadda_rca24_fa221_y0 = f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa216_y4 ^ f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa215_y4;
  assign f_s_dadda_rca24_fa221_y1 = f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa216_y4 & f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa215_y4;
  assign f_s_dadda_rca24_fa221_y2 = f_s_dadda_rca24_fa221_y0 ^ f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa214_y4;
  assign f_s_dadda_rca24_fa221_y3 = f_s_dadda_rca24_fa221_y0 & f_s_dadda_rca24_fa221_f_s_dadda_rca24_fa214_y4;
  assign f_s_dadda_rca24_fa221_y4 = f_s_dadda_rca24_fa221_y1 | f_s_dadda_rca24_fa221_y3;
  assign f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa213_y4 = f_s_dadda_rca24_fa213_y4;
  assign f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa212_y4 = f_s_dadda_rca24_fa212_y4;
  assign f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa211_y4 = f_s_dadda_rca24_fa211_y4;
  assign f_s_dadda_rca24_fa222_y0 = f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa213_y4 ^ f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa212_y4;
  assign f_s_dadda_rca24_fa222_y1 = f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa213_y4 & f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa212_y4;
  assign f_s_dadda_rca24_fa222_y2 = f_s_dadda_rca24_fa222_y0 ^ f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa211_y4;
  assign f_s_dadda_rca24_fa222_y3 = f_s_dadda_rca24_fa222_y0 & f_s_dadda_rca24_fa222_f_s_dadda_rca24_fa211_y4;
  assign f_s_dadda_rca24_fa222_y4 = f_s_dadda_rca24_fa222_y1 | f_s_dadda_rca24_fa222_y3;
  assign f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa210_y4 = f_s_dadda_rca24_fa210_y4;
  assign f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa209_y4 = f_s_dadda_rca24_fa209_y4;
  assign f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa208_y4 = f_s_dadda_rca24_fa208_y4;
  assign f_s_dadda_rca24_fa223_y0 = f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa210_y4 ^ f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa209_y4;
  assign f_s_dadda_rca24_fa223_y1 = f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa210_y4 & f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa209_y4;
  assign f_s_dadda_rca24_fa223_y2 = f_s_dadda_rca24_fa223_y0 ^ f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa208_y4;
  assign f_s_dadda_rca24_fa223_y3 = f_s_dadda_rca24_fa223_y0 & f_s_dadda_rca24_fa223_f_s_dadda_rca24_fa208_y4;
  assign f_s_dadda_rca24_fa223_y4 = f_s_dadda_rca24_fa223_y1 | f_s_dadda_rca24_fa223_y3;
  assign f_s_dadda_rca24_and_22_6_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_22_6_y0 = f_s_dadda_rca24_and_22_6_a_22 & f_s_dadda_rca24_and_22_6_b_6;
  assign f_s_dadda_rca24_and_21_7_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_21_7_y0 = f_s_dadda_rca24_and_21_7_a_21 & f_s_dadda_rca24_and_21_7_b_7;
  assign f_s_dadda_rca24_fa224_f_s_dadda_rca24_fa207_y4 = f_s_dadda_rca24_fa207_y4;
  assign f_s_dadda_rca24_fa224_f_s_dadda_rca24_and_22_6_y0 = f_s_dadda_rca24_and_22_6_y0;
  assign f_s_dadda_rca24_fa224_f_s_dadda_rca24_and_21_7_y0 = f_s_dadda_rca24_and_21_7_y0;
  assign f_s_dadda_rca24_fa224_y0 = f_s_dadda_rca24_fa224_f_s_dadda_rca24_fa207_y4 ^ f_s_dadda_rca24_fa224_f_s_dadda_rca24_and_22_6_y0;
  assign f_s_dadda_rca24_fa224_y1 = f_s_dadda_rca24_fa224_f_s_dadda_rca24_fa207_y4 & f_s_dadda_rca24_fa224_f_s_dadda_rca24_and_22_6_y0;
  assign f_s_dadda_rca24_fa224_y2 = f_s_dadda_rca24_fa224_y0 ^ f_s_dadda_rca24_fa224_f_s_dadda_rca24_and_21_7_y0;
  assign f_s_dadda_rca24_fa224_y3 = f_s_dadda_rca24_fa224_y0 & f_s_dadda_rca24_fa224_f_s_dadda_rca24_and_21_7_y0;
  assign f_s_dadda_rca24_fa224_y4 = f_s_dadda_rca24_fa224_y1 | f_s_dadda_rca24_fa224_y3;
  assign f_s_dadda_rca24_and_20_8_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_20_8_y0 = f_s_dadda_rca24_and_20_8_a_20 & f_s_dadda_rca24_and_20_8_b_8;
  assign f_s_dadda_rca24_and_19_9_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_19_9_y0 = f_s_dadda_rca24_and_19_9_a_19 & f_s_dadda_rca24_and_19_9_b_9;
  assign f_s_dadda_rca24_and_18_10_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_18_10_y0 = f_s_dadda_rca24_and_18_10_a_18 & f_s_dadda_rca24_and_18_10_b_10;
  assign f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_20_8_y0 = f_s_dadda_rca24_and_20_8_y0;
  assign f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_19_9_y0 = f_s_dadda_rca24_and_19_9_y0;
  assign f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_18_10_y0 = f_s_dadda_rca24_and_18_10_y0;
  assign f_s_dadda_rca24_fa225_y0 = f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_20_8_y0 ^ f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_19_9_y0;
  assign f_s_dadda_rca24_fa225_y1 = f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_20_8_y0 & f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_19_9_y0;
  assign f_s_dadda_rca24_fa225_y2 = f_s_dadda_rca24_fa225_y0 ^ f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_18_10_y0;
  assign f_s_dadda_rca24_fa225_y3 = f_s_dadda_rca24_fa225_y0 & f_s_dadda_rca24_fa225_f_s_dadda_rca24_and_18_10_y0;
  assign f_s_dadda_rca24_fa225_y4 = f_s_dadda_rca24_fa225_y1 | f_s_dadda_rca24_fa225_y3;
  assign f_s_dadda_rca24_and_17_11_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_17_11_y0 = f_s_dadda_rca24_and_17_11_a_17 & f_s_dadda_rca24_and_17_11_b_11;
  assign f_s_dadda_rca24_and_16_12_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_16_12_y0 = f_s_dadda_rca24_and_16_12_a_16 & f_s_dadda_rca24_and_16_12_b_12;
  assign f_s_dadda_rca24_and_15_13_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_15_13_y0 = f_s_dadda_rca24_and_15_13_a_15 & f_s_dadda_rca24_and_15_13_b_13;
  assign f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_17_11_y0 = f_s_dadda_rca24_and_17_11_y0;
  assign f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_16_12_y0 = f_s_dadda_rca24_and_16_12_y0;
  assign f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_15_13_y0 = f_s_dadda_rca24_and_15_13_y0;
  assign f_s_dadda_rca24_fa226_y0 = f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_17_11_y0 ^ f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_16_12_y0;
  assign f_s_dadda_rca24_fa226_y1 = f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_17_11_y0 & f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_16_12_y0;
  assign f_s_dadda_rca24_fa226_y2 = f_s_dadda_rca24_fa226_y0 ^ f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_15_13_y0;
  assign f_s_dadda_rca24_fa226_y3 = f_s_dadda_rca24_fa226_y0 & f_s_dadda_rca24_fa226_f_s_dadda_rca24_and_15_13_y0;
  assign f_s_dadda_rca24_fa226_y4 = f_s_dadda_rca24_fa226_y1 | f_s_dadda_rca24_fa226_y3;
  assign f_s_dadda_rca24_and_14_14_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_14_14_y0 = f_s_dadda_rca24_and_14_14_a_14 & f_s_dadda_rca24_and_14_14_b_14;
  assign f_s_dadda_rca24_and_13_15_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_13_15_y0 = f_s_dadda_rca24_and_13_15_a_13 & f_s_dadda_rca24_and_13_15_b_15;
  assign f_s_dadda_rca24_and_12_16_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_12_16_y0 = f_s_dadda_rca24_and_12_16_a_12 & f_s_dadda_rca24_and_12_16_b_16;
  assign f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_14_14_y0 = f_s_dadda_rca24_and_14_14_y0;
  assign f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_13_15_y0 = f_s_dadda_rca24_and_13_15_y0;
  assign f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_12_16_y0 = f_s_dadda_rca24_and_12_16_y0;
  assign f_s_dadda_rca24_fa227_y0 = f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_14_14_y0 ^ f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_13_15_y0;
  assign f_s_dadda_rca24_fa227_y1 = f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_14_14_y0 & f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_13_15_y0;
  assign f_s_dadda_rca24_fa227_y2 = f_s_dadda_rca24_fa227_y0 ^ f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_12_16_y0;
  assign f_s_dadda_rca24_fa227_y3 = f_s_dadda_rca24_fa227_y0 & f_s_dadda_rca24_fa227_f_s_dadda_rca24_and_12_16_y0;
  assign f_s_dadda_rca24_fa227_y4 = f_s_dadda_rca24_fa227_y1 | f_s_dadda_rca24_fa227_y3;
  assign f_s_dadda_rca24_and_11_17_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_11_17_y0 = f_s_dadda_rca24_and_11_17_a_11 & f_s_dadda_rca24_and_11_17_b_17;
  assign f_s_dadda_rca24_and_10_18_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_10_18_y0 = f_s_dadda_rca24_and_10_18_a_10 & f_s_dadda_rca24_and_10_18_b_18;
  assign f_s_dadda_rca24_and_9_19_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_9_19_y0 = f_s_dadda_rca24_and_9_19_a_9 & f_s_dadda_rca24_and_9_19_b_19;
  assign f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_11_17_y0 = f_s_dadda_rca24_and_11_17_y0;
  assign f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_10_18_y0 = f_s_dadda_rca24_and_10_18_y0;
  assign f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_9_19_y0 = f_s_dadda_rca24_and_9_19_y0;
  assign f_s_dadda_rca24_fa228_y0 = f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_11_17_y0 ^ f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_10_18_y0;
  assign f_s_dadda_rca24_fa228_y1 = f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_11_17_y0 & f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_10_18_y0;
  assign f_s_dadda_rca24_fa228_y2 = f_s_dadda_rca24_fa228_y0 ^ f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_9_19_y0;
  assign f_s_dadda_rca24_fa228_y3 = f_s_dadda_rca24_fa228_y0 & f_s_dadda_rca24_fa228_f_s_dadda_rca24_and_9_19_y0;
  assign f_s_dadda_rca24_fa228_y4 = f_s_dadda_rca24_fa228_y1 | f_s_dadda_rca24_fa228_y3;
  assign f_s_dadda_rca24_and_8_20_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_8_20_y0 = f_s_dadda_rca24_and_8_20_a_8 & f_s_dadda_rca24_and_8_20_b_20;
  assign f_s_dadda_rca24_and_7_21_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_7_21_y0 = f_s_dadda_rca24_and_7_21_a_7 & f_s_dadda_rca24_and_7_21_b_21;
  assign f_s_dadda_rca24_and_6_22_a_6 = a_6;
  assign f_s_dadda_rca24_and_6_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_6_22_y0 = f_s_dadda_rca24_and_6_22_a_6 & f_s_dadda_rca24_and_6_22_b_22;
  assign f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_8_20_y0 = f_s_dadda_rca24_and_8_20_y0;
  assign f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_7_21_y0 = f_s_dadda_rca24_and_7_21_y0;
  assign f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_6_22_y0 = f_s_dadda_rca24_and_6_22_y0;
  assign f_s_dadda_rca24_fa229_y0 = f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_8_20_y0 ^ f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_7_21_y0;
  assign f_s_dadda_rca24_fa229_y1 = f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_8_20_y0 & f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_7_21_y0;
  assign f_s_dadda_rca24_fa229_y2 = f_s_dadda_rca24_fa229_y0 ^ f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_6_22_y0;
  assign f_s_dadda_rca24_fa229_y3 = f_s_dadda_rca24_fa229_y0 & f_s_dadda_rca24_fa229_f_s_dadda_rca24_and_6_22_y0;
  assign f_s_dadda_rca24_fa229_y4 = f_s_dadda_rca24_fa229_y1 | f_s_dadda_rca24_fa229_y3;
  assign f_s_dadda_rca24_nand_5_23_a_5 = a_5;
  assign f_s_dadda_rca24_nand_5_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_5_23_y0 = ~(f_s_dadda_rca24_nand_5_23_a_5 & f_s_dadda_rca24_nand_5_23_b_23);
  assign f_s_dadda_rca24_fa230_f_s_dadda_rca24_nand_5_23_y0 = f_s_dadda_rca24_nand_5_23_y0;
  assign f_s_dadda_rca24_fa230_f_s_dadda_rca24_fa24_y2 = f_s_dadda_rca24_fa24_y2;
  assign f_s_dadda_rca24_fa230_f_s_dadda_rca24_fa220_y2 = f_s_dadda_rca24_fa220_y2;
  assign f_s_dadda_rca24_fa230_y0 = f_s_dadda_rca24_fa230_f_s_dadda_rca24_nand_5_23_y0 ^ f_s_dadda_rca24_fa230_f_s_dadda_rca24_fa24_y2;
  assign f_s_dadda_rca24_fa230_y1 = f_s_dadda_rca24_fa230_f_s_dadda_rca24_nand_5_23_y0 & f_s_dadda_rca24_fa230_f_s_dadda_rca24_fa24_y2;
  assign f_s_dadda_rca24_fa230_y2 = f_s_dadda_rca24_fa230_y0 ^ f_s_dadda_rca24_fa230_f_s_dadda_rca24_fa220_y2;
  assign f_s_dadda_rca24_fa230_y3 = f_s_dadda_rca24_fa230_y0 & f_s_dadda_rca24_fa230_f_s_dadda_rca24_fa220_y2;
  assign f_s_dadda_rca24_fa230_y4 = f_s_dadda_rca24_fa230_y1 | f_s_dadda_rca24_fa230_y3;
  assign f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa221_y2 = f_s_dadda_rca24_fa221_y2;
  assign f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa222_y2 = f_s_dadda_rca24_fa222_y2;
  assign f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa223_y2 = f_s_dadda_rca24_fa223_y2;
  assign f_s_dadda_rca24_fa231_y0 = f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa221_y2 ^ f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa222_y2;
  assign f_s_dadda_rca24_fa231_y1 = f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa221_y2 & f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa222_y2;
  assign f_s_dadda_rca24_fa231_y2 = f_s_dadda_rca24_fa231_y0 ^ f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa223_y2;
  assign f_s_dadda_rca24_fa231_y3 = f_s_dadda_rca24_fa231_y0 & f_s_dadda_rca24_fa231_f_s_dadda_rca24_fa223_y2;
  assign f_s_dadda_rca24_fa231_y4 = f_s_dadda_rca24_fa231_y1 | f_s_dadda_rca24_fa231_y3;
  assign f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa224_y2 = f_s_dadda_rca24_fa224_y2;
  assign f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa225_y2 = f_s_dadda_rca24_fa225_y2;
  assign f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa226_y2 = f_s_dadda_rca24_fa226_y2;
  assign f_s_dadda_rca24_fa232_y0 = f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa224_y2 ^ f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa225_y2;
  assign f_s_dadda_rca24_fa232_y1 = f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa224_y2 & f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa225_y2;
  assign f_s_dadda_rca24_fa232_y2 = f_s_dadda_rca24_fa232_y0 ^ f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa226_y2;
  assign f_s_dadda_rca24_fa232_y3 = f_s_dadda_rca24_fa232_y0 & f_s_dadda_rca24_fa232_f_s_dadda_rca24_fa226_y2;
  assign f_s_dadda_rca24_fa232_y4 = f_s_dadda_rca24_fa232_y1 | f_s_dadda_rca24_fa232_y3;
  assign f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa232_y4 = f_s_dadda_rca24_fa232_y4;
  assign f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa231_y4 = f_s_dadda_rca24_fa231_y4;
  assign f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa230_y4 = f_s_dadda_rca24_fa230_y4;
  assign f_s_dadda_rca24_fa233_y0 = f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa232_y4 ^ f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa231_y4;
  assign f_s_dadda_rca24_fa233_y1 = f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa232_y4 & f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa231_y4;
  assign f_s_dadda_rca24_fa233_y2 = f_s_dadda_rca24_fa233_y0 ^ f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa230_y4;
  assign f_s_dadda_rca24_fa233_y3 = f_s_dadda_rca24_fa233_y0 & f_s_dadda_rca24_fa233_f_s_dadda_rca24_fa230_y4;
  assign f_s_dadda_rca24_fa233_y4 = f_s_dadda_rca24_fa233_y1 | f_s_dadda_rca24_fa233_y3;
  assign f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa229_y4 = f_s_dadda_rca24_fa229_y4;
  assign f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa228_y4 = f_s_dadda_rca24_fa228_y4;
  assign f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa227_y4 = f_s_dadda_rca24_fa227_y4;
  assign f_s_dadda_rca24_fa234_y0 = f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa229_y4 ^ f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa228_y4;
  assign f_s_dadda_rca24_fa234_y1 = f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa229_y4 & f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa228_y4;
  assign f_s_dadda_rca24_fa234_y2 = f_s_dadda_rca24_fa234_y0 ^ f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa227_y4;
  assign f_s_dadda_rca24_fa234_y3 = f_s_dadda_rca24_fa234_y0 & f_s_dadda_rca24_fa234_f_s_dadda_rca24_fa227_y4;
  assign f_s_dadda_rca24_fa234_y4 = f_s_dadda_rca24_fa234_y1 | f_s_dadda_rca24_fa234_y3;
  assign f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa226_y4 = f_s_dadda_rca24_fa226_y4;
  assign f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa225_y4 = f_s_dadda_rca24_fa225_y4;
  assign f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa224_y4 = f_s_dadda_rca24_fa224_y4;
  assign f_s_dadda_rca24_fa235_y0 = f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa226_y4 ^ f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa225_y4;
  assign f_s_dadda_rca24_fa235_y1 = f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa226_y4 & f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa225_y4;
  assign f_s_dadda_rca24_fa235_y2 = f_s_dadda_rca24_fa235_y0 ^ f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa224_y4;
  assign f_s_dadda_rca24_fa235_y3 = f_s_dadda_rca24_fa235_y0 & f_s_dadda_rca24_fa235_f_s_dadda_rca24_fa224_y4;
  assign f_s_dadda_rca24_fa235_y4 = f_s_dadda_rca24_fa235_y1 | f_s_dadda_rca24_fa235_y3;
  assign f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa223_y4 = f_s_dadda_rca24_fa223_y4;
  assign f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa222_y4 = f_s_dadda_rca24_fa222_y4;
  assign f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa221_y4 = f_s_dadda_rca24_fa221_y4;
  assign f_s_dadda_rca24_fa236_y0 = f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa223_y4 ^ f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa222_y4;
  assign f_s_dadda_rca24_fa236_y1 = f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa223_y4 & f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa222_y4;
  assign f_s_dadda_rca24_fa236_y2 = f_s_dadda_rca24_fa236_y0 ^ f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa221_y4;
  assign f_s_dadda_rca24_fa236_y3 = f_s_dadda_rca24_fa236_y0 & f_s_dadda_rca24_fa236_f_s_dadda_rca24_fa221_y4;
  assign f_s_dadda_rca24_fa236_y4 = f_s_dadda_rca24_fa236_y1 | f_s_dadda_rca24_fa236_y3;
  assign f_s_dadda_rca24_nand_23_6_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_6_b_6 = b_6;
  assign f_s_dadda_rca24_nand_23_6_y0 = ~(f_s_dadda_rca24_nand_23_6_a_23 & f_s_dadda_rca24_nand_23_6_b_6);
  assign f_s_dadda_rca24_fa237_f_s_dadda_rca24_fa220_y4 = f_s_dadda_rca24_fa220_y4;
  assign f_s_dadda_rca24_fa237_f_s_dadda_rca24_fa24_y4 = f_s_dadda_rca24_fa24_y4;
  assign f_s_dadda_rca24_fa237_f_s_dadda_rca24_nand_23_6_y0 = f_s_dadda_rca24_nand_23_6_y0;
  assign f_s_dadda_rca24_fa237_y0 = f_s_dadda_rca24_fa237_f_s_dadda_rca24_fa220_y4 ^ f_s_dadda_rca24_fa237_f_s_dadda_rca24_fa24_y4;
  assign f_s_dadda_rca24_fa237_y1 = f_s_dadda_rca24_fa237_f_s_dadda_rca24_fa220_y4 & f_s_dadda_rca24_fa237_f_s_dadda_rca24_fa24_y4;
  assign f_s_dadda_rca24_fa237_y2 = f_s_dadda_rca24_fa237_y0 ^ f_s_dadda_rca24_fa237_f_s_dadda_rca24_nand_23_6_y0;
  assign f_s_dadda_rca24_fa237_y3 = f_s_dadda_rca24_fa237_y0 & f_s_dadda_rca24_fa237_f_s_dadda_rca24_nand_23_6_y0;
  assign f_s_dadda_rca24_fa237_y4 = f_s_dadda_rca24_fa237_y1 | f_s_dadda_rca24_fa237_y3;
  assign f_s_dadda_rca24_and_22_7_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_22_7_y0 = f_s_dadda_rca24_and_22_7_a_22 & f_s_dadda_rca24_and_22_7_b_7;
  assign f_s_dadda_rca24_and_21_8_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_21_8_y0 = f_s_dadda_rca24_and_21_8_a_21 & f_s_dadda_rca24_and_21_8_b_8;
  assign f_s_dadda_rca24_and_20_9_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_20_9_y0 = f_s_dadda_rca24_and_20_9_a_20 & f_s_dadda_rca24_and_20_9_b_9;
  assign f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_22_7_y0 = f_s_dadda_rca24_and_22_7_y0;
  assign f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_21_8_y0 = f_s_dadda_rca24_and_21_8_y0;
  assign f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_20_9_y0 = f_s_dadda_rca24_and_20_9_y0;
  assign f_s_dadda_rca24_fa238_y0 = f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_22_7_y0 ^ f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_21_8_y0;
  assign f_s_dadda_rca24_fa238_y1 = f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_22_7_y0 & f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_21_8_y0;
  assign f_s_dadda_rca24_fa238_y2 = f_s_dadda_rca24_fa238_y0 ^ f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_20_9_y0;
  assign f_s_dadda_rca24_fa238_y3 = f_s_dadda_rca24_fa238_y0 & f_s_dadda_rca24_fa238_f_s_dadda_rca24_and_20_9_y0;
  assign f_s_dadda_rca24_fa238_y4 = f_s_dadda_rca24_fa238_y1 | f_s_dadda_rca24_fa238_y3;
  assign f_s_dadda_rca24_and_19_10_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_19_10_y0 = f_s_dadda_rca24_and_19_10_a_19 & f_s_dadda_rca24_and_19_10_b_10;
  assign f_s_dadda_rca24_and_18_11_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_18_11_y0 = f_s_dadda_rca24_and_18_11_a_18 & f_s_dadda_rca24_and_18_11_b_11;
  assign f_s_dadda_rca24_and_17_12_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_17_12_y0 = f_s_dadda_rca24_and_17_12_a_17 & f_s_dadda_rca24_and_17_12_b_12;
  assign f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_19_10_y0 = f_s_dadda_rca24_and_19_10_y0;
  assign f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_18_11_y0 = f_s_dadda_rca24_and_18_11_y0;
  assign f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_17_12_y0 = f_s_dadda_rca24_and_17_12_y0;
  assign f_s_dadda_rca24_fa239_y0 = f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_19_10_y0 ^ f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_18_11_y0;
  assign f_s_dadda_rca24_fa239_y1 = f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_19_10_y0 & f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_18_11_y0;
  assign f_s_dadda_rca24_fa239_y2 = f_s_dadda_rca24_fa239_y0 ^ f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_17_12_y0;
  assign f_s_dadda_rca24_fa239_y3 = f_s_dadda_rca24_fa239_y0 & f_s_dadda_rca24_fa239_f_s_dadda_rca24_and_17_12_y0;
  assign f_s_dadda_rca24_fa239_y4 = f_s_dadda_rca24_fa239_y1 | f_s_dadda_rca24_fa239_y3;
  assign f_s_dadda_rca24_and_16_13_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_16_13_y0 = f_s_dadda_rca24_and_16_13_a_16 & f_s_dadda_rca24_and_16_13_b_13;
  assign f_s_dadda_rca24_and_15_14_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_15_14_y0 = f_s_dadda_rca24_and_15_14_a_15 & f_s_dadda_rca24_and_15_14_b_14;
  assign f_s_dadda_rca24_and_14_15_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_14_15_y0 = f_s_dadda_rca24_and_14_15_a_14 & f_s_dadda_rca24_and_14_15_b_15;
  assign f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_16_13_y0 = f_s_dadda_rca24_and_16_13_y0;
  assign f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_15_14_y0 = f_s_dadda_rca24_and_15_14_y0;
  assign f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_14_15_y0 = f_s_dadda_rca24_and_14_15_y0;
  assign f_s_dadda_rca24_fa240_y0 = f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_16_13_y0 ^ f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_15_14_y0;
  assign f_s_dadda_rca24_fa240_y1 = f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_16_13_y0 & f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_15_14_y0;
  assign f_s_dadda_rca24_fa240_y2 = f_s_dadda_rca24_fa240_y0 ^ f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_14_15_y0;
  assign f_s_dadda_rca24_fa240_y3 = f_s_dadda_rca24_fa240_y0 & f_s_dadda_rca24_fa240_f_s_dadda_rca24_and_14_15_y0;
  assign f_s_dadda_rca24_fa240_y4 = f_s_dadda_rca24_fa240_y1 | f_s_dadda_rca24_fa240_y3;
  assign f_s_dadda_rca24_and_13_16_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_13_16_y0 = f_s_dadda_rca24_and_13_16_a_13 & f_s_dadda_rca24_and_13_16_b_16;
  assign f_s_dadda_rca24_and_12_17_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_12_17_y0 = f_s_dadda_rca24_and_12_17_a_12 & f_s_dadda_rca24_and_12_17_b_17;
  assign f_s_dadda_rca24_and_11_18_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_11_18_y0 = f_s_dadda_rca24_and_11_18_a_11 & f_s_dadda_rca24_and_11_18_b_18;
  assign f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_13_16_y0 = f_s_dadda_rca24_and_13_16_y0;
  assign f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_12_17_y0 = f_s_dadda_rca24_and_12_17_y0;
  assign f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_11_18_y0 = f_s_dadda_rca24_and_11_18_y0;
  assign f_s_dadda_rca24_fa241_y0 = f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_13_16_y0 ^ f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_12_17_y0;
  assign f_s_dadda_rca24_fa241_y1 = f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_13_16_y0 & f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_12_17_y0;
  assign f_s_dadda_rca24_fa241_y2 = f_s_dadda_rca24_fa241_y0 ^ f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_11_18_y0;
  assign f_s_dadda_rca24_fa241_y3 = f_s_dadda_rca24_fa241_y0 & f_s_dadda_rca24_fa241_f_s_dadda_rca24_and_11_18_y0;
  assign f_s_dadda_rca24_fa241_y4 = f_s_dadda_rca24_fa241_y1 | f_s_dadda_rca24_fa241_y3;
  assign f_s_dadda_rca24_and_10_19_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_10_19_y0 = f_s_dadda_rca24_and_10_19_a_10 & f_s_dadda_rca24_and_10_19_b_19;
  assign f_s_dadda_rca24_and_9_20_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_9_20_y0 = f_s_dadda_rca24_and_9_20_a_9 & f_s_dadda_rca24_and_9_20_b_20;
  assign f_s_dadda_rca24_and_8_21_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_8_21_y0 = f_s_dadda_rca24_and_8_21_a_8 & f_s_dadda_rca24_and_8_21_b_21;
  assign f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_10_19_y0 = f_s_dadda_rca24_and_10_19_y0;
  assign f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_9_20_y0 = f_s_dadda_rca24_and_9_20_y0;
  assign f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_8_21_y0 = f_s_dadda_rca24_and_8_21_y0;
  assign f_s_dadda_rca24_fa242_y0 = f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_10_19_y0 ^ f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_9_20_y0;
  assign f_s_dadda_rca24_fa242_y1 = f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_10_19_y0 & f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_9_20_y0;
  assign f_s_dadda_rca24_fa242_y2 = f_s_dadda_rca24_fa242_y0 ^ f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_8_21_y0;
  assign f_s_dadda_rca24_fa242_y3 = f_s_dadda_rca24_fa242_y0 & f_s_dadda_rca24_fa242_f_s_dadda_rca24_and_8_21_y0;
  assign f_s_dadda_rca24_fa242_y4 = f_s_dadda_rca24_fa242_y1 | f_s_dadda_rca24_fa242_y3;
  assign f_s_dadda_rca24_and_7_22_a_7 = a_7;
  assign f_s_dadda_rca24_and_7_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_7_22_y0 = f_s_dadda_rca24_and_7_22_a_7 & f_s_dadda_rca24_and_7_22_b_22;
  assign f_s_dadda_rca24_nand_6_23_a_6 = a_6;
  assign f_s_dadda_rca24_nand_6_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_6_23_y0 = ~(f_s_dadda_rca24_nand_6_23_a_6 & f_s_dadda_rca24_nand_6_23_b_23);
  assign f_s_dadda_rca24_fa243_f_s_dadda_rca24_and_7_22_y0 = f_s_dadda_rca24_and_7_22_y0;
  assign f_s_dadda_rca24_fa243_f_s_dadda_rca24_nand_6_23_y0 = f_s_dadda_rca24_nand_6_23_y0;
  assign f_s_dadda_rca24_fa243_f_s_dadda_rca24_fa233_y2 = f_s_dadda_rca24_fa233_y2;
  assign f_s_dadda_rca24_fa243_y0 = f_s_dadda_rca24_fa243_f_s_dadda_rca24_and_7_22_y0 ^ f_s_dadda_rca24_fa243_f_s_dadda_rca24_nand_6_23_y0;
  assign f_s_dadda_rca24_fa243_y1 = f_s_dadda_rca24_fa243_f_s_dadda_rca24_and_7_22_y0 & f_s_dadda_rca24_fa243_f_s_dadda_rca24_nand_6_23_y0;
  assign f_s_dadda_rca24_fa243_y2 = f_s_dadda_rca24_fa243_y0 ^ f_s_dadda_rca24_fa243_f_s_dadda_rca24_fa233_y2;
  assign f_s_dadda_rca24_fa243_y3 = f_s_dadda_rca24_fa243_y0 & f_s_dadda_rca24_fa243_f_s_dadda_rca24_fa233_y2;
  assign f_s_dadda_rca24_fa243_y4 = f_s_dadda_rca24_fa243_y1 | f_s_dadda_rca24_fa243_y3;
  assign f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa234_y2 = f_s_dadda_rca24_fa234_y2;
  assign f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa235_y2 = f_s_dadda_rca24_fa235_y2;
  assign f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa236_y2 = f_s_dadda_rca24_fa236_y2;
  assign f_s_dadda_rca24_fa244_y0 = f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa234_y2 ^ f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa235_y2;
  assign f_s_dadda_rca24_fa244_y1 = f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa234_y2 & f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa235_y2;
  assign f_s_dadda_rca24_fa244_y2 = f_s_dadda_rca24_fa244_y0 ^ f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa236_y2;
  assign f_s_dadda_rca24_fa244_y3 = f_s_dadda_rca24_fa244_y0 & f_s_dadda_rca24_fa244_f_s_dadda_rca24_fa236_y2;
  assign f_s_dadda_rca24_fa244_y4 = f_s_dadda_rca24_fa244_y1 | f_s_dadda_rca24_fa244_y3;
  assign f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa237_y2 = f_s_dadda_rca24_fa237_y2;
  assign f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa238_y2 = f_s_dadda_rca24_fa238_y2;
  assign f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa239_y2 = f_s_dadda_rca24_fa239_y2;
  assign f_s_dadda_rca24_fa245_y0 = f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa237_y2 ^ f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa238_y2;
  assign f_s_dadda_rca24_fa245_y1 = f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa237_y2 & f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa238_y2;
  assign f_s_dadda_rca24_fa245_y2 = f_s_dadda_rca24_fa245_y0 ^ f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa239_y2;
  assign f_s_dadda_rca24_fa245_y3 = f_s_dadda_rca24_fa245_y0 & f_s_dadda_rca24_fa245_f_s_dadda_rca24_fa239_y2;
  assign f_s_dadda_rca24_fa245_y4 = f_s_dadda_rca24_fa245_y1 | f_s_dadda_rca24_fa245_y3;
  assign f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa245_y4 = f_s_dadda_rca24_fa245_y4;
  assign f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa244_y4 = f_s_dadda_rca24_fa244_y4;
  assign f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa243_y4 = f_s_dadda_rca24_fa243_y4;
  assign f_s_dadda_rca24_fa246_y0 = f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa245_y4 ^ f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa244_y4;
  assign f_s_dadda_rca24_fa246_y1 = f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa245_y4 & f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa244_y4;
  assign f_s_dadda_rca24_fa246_y2 = f_s_dadda_rca24_fa246_y0 ^ f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa243_y4;
  assign f_s_dadda_rca24_fa246_y3 = f_s_dadda_rca24_fa246_y0 & f_s_dadda_rca24_fa246_f_s_dadda_rca24_fa243_y4;
  assign f_s_dadda_rca24_fa246_y4 = f_s_dadda_rca24_fa246_y1 | f_s_dadda_rca24_fa246_y3;
  assign f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa242_y4 = f_s_dadda_rca24_fa242_y4;
  assign f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa241_y4 = f_s_dadda_rca24_fa241_y4;
  assign f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa240_y4 = f_s_dadda_rca24_fa240_y4;
  assign f_s_dadda_rca24_fa247_y0 = f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa242_y4 ^ f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa241_y4;
  assign f_s_dadda_rca24_fa247_y1 = f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa242_y4 & f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa241_y4;
  assign f_s_dadda_rca24_fa247_y2 = f_s_dadda_rca24_fa247_y0 ^ f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa240_y4;
  assign f_s_dadda_rca24_fa247_y3 = f_s_dadda_rca24_fa247_y0 & f_s_dadda_rca24_fa247_f_s_dadda_rca24_fa240_y4;
  assign f_s_dadda_rca24_fa247_y4 = f_s_dadda_rca24_fa247_y1 | f_s_dadda_rca24_fa247_y3;
  assign f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa239_y4 = f_s_dadda_rca24_fa239_y4;
  assign f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa238_y4 = f_s_dadda_rca24_fa238_y4;
  assign f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa237_y4 = f_s_dadda_rca24_fa237_y4;
  assign f_s_dadda_rca24_fa248_y0 = f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa239_y4 ^ f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa238_y4;
  assign f_s_dadda_rca24_fa248_y1 = f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa239_y4 & f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa238_y4;
  assign f_s_dadda_rca24_fa248_y2 = f_s_dadda_rca24_fa248_y0 ^ f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa237_y4;
  assign f_s_dadda_rca24_fa248_y3 = f_s_dadda_rca24_fa248_y0 & f_s_dadda_rca24_fa248_f_s_dadda_rca24_fa237_y4;
  assign f_s_dadda_rca24_fa248_y4 = f_s_dadda_rca24_fa248_y1 | f_s_dadda_rca24_fa248_y3;
  assign f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa236_y4 = f_s_dadda_rca24_fa236_y4;
  assign f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa235_y4 = f_s_dadda_rca24_fa235_y4;
  assign f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa234_y4 = f_s_dadda_rca24_fa234_y4;
  assign f_s_dadda_rca24_fa249_y0 = f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa236_y4 ^ f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa235_y4;
  assign f_s_dadda_rca24_fa249_y1 = f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa236_y4 & f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa235_y4;
  assign f_s_dadda_rca24_fa249_y2 = f_s_dadda_rca24_fa249_y0 ^ f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa234_y4;
  assign f_s_dadda_rca24_fa249_y3 = f_s_dadda_rca24_fa249_y0 & f_s_dadda_rca24_fa249_f_s_dadda_rca24_fa234_y4;
  assign f_s_dadda_rca24_fa249_y4 = f_s_dadda_rca24_fa249_y1 | f_s_dadda_rca24_fa249_y3;
  assign f_s_dadda_rca24_nand_23_7_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_7_b_7 = b_7;
  assign f_s_dadda_rca24_nand_23_7_y0 = ~(f_s_dadda_rca24_nand_23_7_a_23 & f_s_dadda_rca24_nand_23_7_b_7);
  assign f_s_dadda_rca24_and_22_8_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_22_8_y0 = f_s_dadda_rca24_and_22_8_a_22 & f_s_dadda_rca24_and_22_8_b_8;
  assign f_s_dadda_rca24_fa250_f_s_dadda_rca24_fa233_y4 = f_s_dadda_rca24_fa233_y4;
  assign f_s_dadda_rca24_fa250_f_s_dadda_rca24_nand_23_7_y0 = f_s_dadda_rca24_nand_23_7_y0;
  assign f_s_dadda_rca24_fa250_f_s_dadda_rca24_and_22_8_y0 = f_s_dadda_rca24_and_22_8_y0;
  assign f_s_dadda_rca24_fa250_y0 = f_s_dadda_rca24_fa250_f_s_dadda_rca24_fa233_y4 ^ f_s_dadda_rca24_fa250_f_s_dadda_rca24_nand_23_7_y0;
  assign f_s_dadda_rca24_fa250_y1 = f_s_dadda_rca24_fa250_f_s_dadda_rca24_fa233_y4 & f_s_dadda_rca24_fa250_f_s_dadda_rca24_nand_23_7_y0;
  assign f_s_dadda_rca24_fa250_y2 = f_s_dadda_rca24_fa250_y0 ^ f_s_dadda_rca24_fa250_f_s_dadda_rca24_and_22_8_y0;
  assign f_s_dadda_rca24_fa250_y3 = f_s_dadda_rca24_fa250_y0 & f_s_dadda_rca24_fa250_f_s_dadda_rca24_and_22_8_y0;
  assign f_s_dadda_rca24_fa250_y4 = f_s_dadda_rca24_fa250_y1 | f_s_dadda_rca24_fa250_y3;
  assign f_s_dadda_rca24_and_21_9_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_21_9_y0 = f_s_dadda_rca24_and_21_9_a_21 & f_s_dadda_rca24_and_21_9_b_9;
  assign f_s_dadda_rca24_and_20_10_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_20_10_y0 = f_s_dadda_rca24_and_20_10_a_20 & f_s_dadda_rca24_and_20_10_b_10;
  assign f_s_dadda_rca24_and_19_11_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_19_11_y0 = f_s_dadda_rca24_and_19_11_a_19 & f_s_dadda_rca24_and_19_11_b_11;
  assign f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_21_9_y0 = f_s_dadda_rca24_and_21_9_y0;
  assign f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_20_10_y0 = f_s_dadda_rca24_and_20_10_y0;
  assign f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_19_11_y0 = f_s_dadda_rca24_and_19_11_y0;
  assign f_s_dadda_rca24_fa251_y0 = f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_21_9_y0 ^ f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_20_10_y0;
  assign f_s_dadda_rca24_fa251_y1 = f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_21_9_y0 & f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_20_10_y0;
  assign f_s_dadda_rca24_fa251_y2 = f_s_dadda_rca24_fa251_y0 ^ f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_19_11_y0;
  assign f_s_dadda_rca24_fa251_y3 = f_s_dadda_rca24_fa251_y0 & f_s_dadda_rca24_fa251_f_s_dadda_rca24_and_19_11_y0;
  assign f_s_dadda_rca24_fa251_y4 = f_s_dadda_rca24_fa251_y1 | f_s_dadda_rca24_fa251_y3;
  assign f_s_dadda_rca24_and_18_12_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_18_12_y0 = f_s_dadda_rca24_and_18_12_a_18 & f_s_dadda_rca24_and_18_12_b_12;
  assign f_s_dadda_rca24_and_17_13_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_17_13_y0 = f_s_dadda_rca24_and_17_13_a_17 & f_s_dadda_rca24_and_17_13_b_13;
  assign f_s_dadda_rca24_and_16_14_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_16_14_y0 = f_s_dadda_rca24_and_16_14_a_16 & f_s_dadda_rca24_and_16_14_b_14;
  assign f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_18_12_y0 = f_s_dadda_rca24_and_18_12_y0;
  assign f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_17_13_y0 = f_s_dadda_rca24_and_17_13_y0;
  assign f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_16_14_y0 = f_s_dadda_rca24_and_16_14_y0;
  assign f_s_dadda_rca24_fa252_y0 = f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_18_12_y0 ^ f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_17_13_y0;
  assign f_s_dadda_rca24_fa252_y1 = f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_18_12_y0 & f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_17_13_y0;
  assign f_s_dadda_rca24_fa252_y2 = f_s_dadda_rca24_fa252_y0 ^ f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_16_14_y0;
  assign f_s_dadda_rca24_fa252_y3 = f_s_dadda_rca24_fa252_y0 & f_s_dadda_rca24_fa252_f_s_dadda_rca24_and_16_14_y0;
  assign f_s_dadda_rca24_fa252_y4 = f_s_dadda_rca24_fa252_y1 | f_s_dadda_rca24_fa252_y3;
  assign f_s_dadda_rca24_and_15_15_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_15_15_y0 = f_s_dadda_rca24_and_15_15_a_15 & f_s_dadda_rca24_and_15_15_b_15;
  assign f_s_dadda_rca24_and_14_16_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_14_16_y0 = f_s_dadda_rca24_and_14_16_a_14 & f_s_dadda_rca24_and_14_16_b_16;
  assign f_s_dadda_rca24_and_13_17_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_13_17_y0 = f_s_dadda_rca24_and_13_17_a_13 & f_s_dadda_rca24_and_13_17_b_17;
  assign f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_15_15_y0 = f_s_dadda_rca24_and_15_15_y0;
  assign f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_14_16_y0 = f_s_dadda_rca24_and_14_16_y0;
  assign f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_13_17_y0 = f_s_dadda_rca24_and_13_17_y0;
  assign f_s_dadda_rca24_fa253_y0 = f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_15_15_y0 ^ f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_14_16_y0;
  assign f_s_dadda_rca24_fa253_y1 = f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_15_15_y0 & f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_14_16_y0;
  assign f_s_dadda_rca24_fa253_y2 = f_s_dadda_rca24_fa253_y0 ^ f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_13_17_y0;
  assign f_s_dadda_rca24_fa253_y3 = f_s_dadda_rca24_fa253_y0 & f_s_dadda_rca24_fa253_f_s_dadda_rca24_and_13_17_y0;
  assign f_s_dadda_rca24_fa253_y4 = f_s_dadda_rca24_fa253_y1 | f_s_dadda_rca24_fa253_y3;
  assign f_s_dadda_rca24_and_12_18_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_12_18_y0 = f_s_dadda_rca24_and_12_18_a_12 & f_s_dadda_rca24_and_12_18_b_18;
  assign f_s_dadda_rca24_and_11_19_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_11_19_y0 = f_s_dadda_rca24_and_11_19_a_11 & f_s_dadda_rca24_and_11_19_b_19;
  assign f_s_dadda_rca24_and_10_20_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_10_20_y0 = f_s_dadda_rca24_and_10_20_a_10 & f_s_dadda_rca24_and_10_20_b_20;
  assign f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_12_18_y0 = f_s_dadda_rca24_and_12_18_y0;
  assign f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_11_19_y0 = f_s_dadda_rca24_and_11_19_y0;
  assign f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_10_20_y0 = f_s_dadda_rca24_and_10_20_y0;
  assign f_s_dadda_rca24_fa254_y0 = f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_12_18_y0 ^ f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_11_19_y0;
  assign f_s_dadda_rca24_fa254_y1 = f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_12_18_y0 & f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_11_19_y0;
  assign f_s_dadda_rca24_fa254_y2 = f_s_dadda_rca24_fa254_y0 ^ f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_10_20_y0;
  assign f_s_dadda_rca24_fa254_y3 = f_s_dadda_rca24_fa254_y0 & f_s_dadda_rca24_fa254_f_s_dadda_rca24_and_10_20_y0;
  assign f_s_dadda_rca24_fa254_y4 = f_s_dadda_rca24_fa254_y1 | f_s_dadda_rca24_fa254_y3;
  assign f_s_dadda_rca24_and_9_21_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_9_21_y0 = f_s_dadda_rca24_and_9_21_a_9 & f_s_dadda_rca24_and_9_21_b_21;
  assign f_s_dadda_rca24_and_8_22_a_8 = a_8;
  assign f_s_dadda_rca24_and_8_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_8_22_y0 = f_s_dadda_rca24_and_8_22_a_8 & f_s_dadda_rca24_and_8_22_b_22;
  assign f_s_dadda_rca24_nand_7_23_a_7 = a_7;
  assign f_s_dadda_rca24_nand_7_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_7_23_y0 = ~(f_s_dadda_rca24_nand_7_23_a_7 & f_s_dadda_rca24_nand_7_23_b_23);
  assign f_s_dadda_rca24_fa255_f_s_dadda_rca24_and_9_21_y0 = f_s_dadda_rca24_and_9_21_y0;
  assign f_s_dadda_rca24_fa255_f_s_dadda_rca24_and_8_22_y0 = f_s_dadda_rca24_and_8_22_y0;
  assign f_s_dadda_rca24_fa255_f_s_dadda_rca24_nand_7_23_y0 = f_s_dadda_rca24_nand_7_23_y0;
  assign f_s_dadda_rca24_fa255_y0 = f_s_dadda_rca24_fa255_f_s_dadda_rca24_and_9_21_y0 ^ f_s_dadda_rca24_fa255_f_s_dadda_rca24_and_8_22_y0;
  assign f_s_dadda_rca24_fa255_y1 = f_s_dadda_rca24_fa255_f_s_dadda_rca24_and_9_21_y0 & f_s_dadda_rca24_fa255_f_s_dadda_rca24_and_8_22_y0;
  assign f_s_dadda_rca24_fa255_y2 = f_s_dadda_rca24_fa255_y0 ^ f_s_dadda_rca24_fa255_f_s_dadda_rca24_nand_7_23_y0;
  assign f_s_dadda_rca24_fa255_y3 = f_s_dadda_rca24_fa255_y0 & f_s_dadda_rca24_fa255_f_s_dadda_rca24_nand_7_23_y0;
  assign f_s_dadda_rca24_fa255_y4 = f_s_dadda_rca24_fa255_y1 | f_s_dadda_rca24_fa255_y3;
  assign f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa246_y2 = f_s_dadda_rca24_fa246_y2;
  assign f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa247_y2 = f_s_dadda_rca24_fa247_y2;
  assign f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa248_y2 = f_s_dadda_rca24_fa248_y2;
  assign f_s_dadda_rca24_fa256_y0 = f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa246_y2 ^ f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa247_y2;
  assign f_s_dadda_rca24_fa256_y1 = f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa246_y2 & f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa247_y2;
  assign f_s_dadda_rca24_fa256_y2 = f_s_dadda_rca24_fa256_y0 ^ f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa248_y2;
  assign f_s_dadda_rca24_fa256_y3 = f_s_dadda_rca24_fa256_y0 & f_s_dadda_rca24_fa256_f_s_dadda_rca24_fa248_y2;
  assign f_s_dadda_rca24_fa256_y4 = f_s_dadda_rca24_fa256_y1 | f_s_dadda_rca24_fa256_y3;
  assign f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa249_y2 = f_s_dadda_rca24_fa249_y2;
  assign f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa250_y2 = f_s_dadda_rca24_fa250_y2;
  assign f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa251_y2 = f_s_dadda_rca24_fa251_y2;
  assign f_s_dadda_rca24_fa257_y0 = f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa249_y2 ^ f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa250_y2;
  assign f_s_dadda_rca24_fa257_y1 = f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa249_y2 & f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa250_y2;
  assign f_s_dadda_rca24_fa257_y2 = f_s_dadda_rca24_fa257_y0 ^ f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa251_y2;
  assign f_s_dadda_rca24_fa257_y3 = f_s_dadda_rca24_fa257_y0 & f_s_dadda_rca24_fa257_f_s_dadda_rca24_fa251_y2;
  assign f_s_dadda_rca24_fa257_y4 = f_s_dadda_rca24_fa257_y1 | f_s_dadda_rca24_fa257_y3;
  assign f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa257_y4 = f_s_dadda_rca24_fa257_y4;
  assign f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa256_y4 = f_s_dadda_rca24_fa256_y4;
  assign f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa255_y4 = f_s_dadda_rca24_fa255_y4;
  assign f_s_dadda_rca24_fa258_y0 = f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa257_y4 ^ f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa256_y4;
  assign f_s_dadda_rca24_fa258_y1 = f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa257_y4 & f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa256_y4;
  assign f_s_dadda_rca24_fa258_y2 = f_s_dadda_rca24_fa258_y0 ^ f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa255_y4;
  assign f_s_dadda_rca24_fa258_y3 = f_s_dadda_rca24_fa258_y0 & f_s_dadda_rca24_fa258_f_s_dadda_rca24_fa255_y4;
  assign f_s_dadda_rca24_fa258_y4 = f_s_dadda_rca24_fa258_y1 | f_s_dadda_rca24_fa258_y3;
  assign f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa254_y4 = f_s_dadda_rca24_fa254_y4;
  assign f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa253_y4 = f_s_dadda_rca24_fa253_y4;
  assign f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa252_y4 = f_s_dadda_rca24_fa252_y4;
  assign f_s_dadda_rca24_fa259_y0 = f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa254_y4 ^ f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa253_y4;
  assign f_s_dadda_rca24_fa259_y1 = f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa254_y4 & f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa253_y4;
  assign f_s_dadda_rca24_fa259_y2 = f_s_dadda_rca24_fa259_y0 ^ f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa252_y4;
  assign f_s_dadda_rca24_fa259_y3 = f_s_dadda_rca24_fa259_y0 & f_s_dadda_rca24_fa259_f_s_dadda_rca24_fa252_y4;
  assign f_s_dadda_rca24_fa259_y4 = f_s_dadda_rca24_fa259_y1 | f_s_dadda_rca24_fa259_y3;
  assign f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa251_y4 = f_s_dadda_rca24_fa251_y4;
  assign f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa250_y4 = f_s_dadda_rca24_fa250_y4;
  assign f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa249_y4 = f_s_dadda_rca24_fa249_y4;
  assign f_s_dadda_rca24_fa260_y0 = f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa251_y4 ^ f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa250_y4;
  assign f_s_dadda_rca24_fa260_y1 = f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa251_y4 & f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa250_y4;
  assign f_s_dadda_rca24_fa260_y2 = f_s_dadda_rca24_fa260_y0 ^ f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa249_y4;
  assign f_s_dadda_rca24_fa260_y3 = f_s_dadda_rca24_fa260_y0 & f_s_dadda_rca24_fa260_f_s_dadda_rca24_fa249_y4;
  assign f_s_dadda_rca24_fa260_y4 = f_s_dadda_rca24_fa260_y1 | f_s_dadda_rca24_fa260_y3;
  assign f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa248_y4 = f_s_dadda_rca24_fa248_y4;
  assign f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa247_y4 = f_s_dadda_rca24_fa247_y4;
  assign f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa246_y4 = f_s_dadda_rca24_fa246_y4;
  assign f_s_dadda_rca24_fa261_y0 = f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa248_y4 ^ f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa247_y4;
  assign f_s_dadda_rca24_fa261_y1 = f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa248_y4 & f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa247_y4;
  assign f_s_dadda_rca24_fa261_y2 = f_s_dadda_rca24_fa261_y0 ^ f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa246_y4;
  assign f_s_dadda_rca24_fa261_y3 = f_s_dadda_rca24_fa261_y0 & f_s_dadda_rca24_fa261_f_s_dadda_rca24_fa246_y4;
  assign f_s_dadda_rca24_fa261_y4 = f_s_dadda_rca24_fa261_y1 | f_s_dadda_rca24_fa261_y3;
  assign f_s_dadda_rca24_nand_23_8_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_8_b_8 = b_8;
  assign f_s_dadda_rca24_nand_23_8_y0 = ~(f_s_dadda_rca24_nand_23_8_a_23 & f_s_dadda_rca24_nand_23_8_b_8);
  assign f_s_dadda_rca24_and_22_9_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_22_9_y0 = f_s_dadda_rca24_and_22_9_a_22 & f_s_dadda_rca24_and_22_9_b_9;
  assign f_s_dadda_rca24_and_21_10_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_21_10_y0 = f_s_dadda_rca24_and_21_10_a_21 & f_s_dadda_rca24_and_21_10_b_10;
  assign f_s_dadda_rca24_fa262_f_s_dadda_rca24_nand_23_8_y0 = f_s_dadda_rca24_nand_23_8_y0;
  assign f_s_dadda_rca24_fa262_f_s_dadda_rca24_and_22_9_y0 = f_s_dadda_rca24_and_22_9_y0;
  assign f_s_dadda_rca24_fa262_f_s_dadda_rca24_and_21_10_y0 = f_s_dadda_rca24_and_21_10_y0;
  assign f_s_dadda_rca24_fa262_y0 = f_s_dadda_rca24_fa262_f_s_dadda_rca24_nand_23_8_y0 ^ f_s_dadda_rca24_fa262_f_s_dadda_rca24_and_22_9_y0;
  assign f_s_dadda_rca24_fa262_y1 = f_s_dadda_rca24_fa262_f_s_dadda_rca24_nand_23_8_y0 & f_s_dadda_rca24_fa262_f_s_dadda_rca24_and_22_9_y0;
  assign f_s_dadda_rca24_fa262_y2 = f_s_dadda_rca24_fa262_y0 ^ f_s_dadda_rca24_fa262_f_s_dadda_rca24_and_21_10_y0;
  assign f_s_dadda_rca24_fa262_y3 = f_s_dadda_rca24_fa262_y0 & f_s_dadda_rca24_fa262_f_s_dadda_rca24_and_21_10_y0;
  assign f_s_dadda_rca24_fa262_y4 = f_s_dadda_rca24_fa262_y1 | f_s_dadda_rca24_fa262_y3;
  assign f_s_dadda_rca24_and_20_11_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_20_11_y0 = f_s_dadda_rca24_and_20_11_a_20 & f_s_dadda_rca24_and_20_11_b_11;
  assign f_s_dadda_rca24_and_19_12_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_19_12_y0 = f_s_dadda_rca24_and_19_12_a_19 & f_s_dadda_rca24_and_19_12_b_12;
  assign f_s_dadda_rca24_and_18_13_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_18_13_y0 = f_s_dadda_rca24_and_18_13_a_18 & f_s_dadda_rca24_and_18_13_b_13;
  assign f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_20_11_y0 = f_s_dadda_rca24_and_20_11_y0;
  assign f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_19_12_y0 = f_s_dadda_rca24_and_19_12_y0;
  assign f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_18_13_y0 = f_s_dadda_rca24_and_18_13_y0;
  assign f_s_dadda_rca24_fa263_y0 = f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_20_11_y0 ^ f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_19_12_y0;
  assign f_s_dadda_rca24_fa263_y1 = f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_20_11_y0 & f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_19_12_y0;
  assign f_s_dadda_rca24_fa263_y2 = f_s_dadda_rca24_fa263_y0 ^ f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_18_13_y0;
  assign f_s_dadda_rca24_fa263_y3 = f_s_dadda_rca24_fa263_y0 & f_s_dadda_rca24_fa263_f_s_dadda_rca24_and_18_13_y0;
  assign f_s_dadda_rca24_fa263_y4 = f_s_dadda_rca24_fa263_y1 | f_s_dadda_rca24_fa263_y3;
  assign f_s_dadda_rca24_and_17_14_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_17_14_y0 = f_s_dadda_rca24_and_17_14_a_17 & f_s_dadda_rca24_and_17_14_b_14;
  assign f_s_dadda_rca24_and_16_15_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_16_15_y0 = f_s_dadda_rca24_and_16_15_a_16 & f_s_dadda_rca24_and_16_15_b_15;
  assign f_s_dadda_rca24_and_15_16_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_15_16_y0 = f_s_dadda_rca24_and_15_16_a_15 & f_s_dadda_rca24_and_15_16_b_16;
  assign f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_17_14_y0 = f_s_dadda_rca24_and_17_14_y0;
  assign f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_16_15_y0 = f_s_dadda_rca24_and_16_15_y0;
  assign f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_15_16_y0 = f_s_dadda_rca24_and_15_16_y0;
  assign f_s_dadda_rca24_fa264_y0 = f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_17_14_y0 ^ f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_16_15_y0;
  assign f_s_dadda_rca24_fa264_y1 = f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_17_14_y0 & f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_16_15_y0;
  assign f_s_dadda_rca24_fa264_y2 = f_s_dadda_rca24_fa264_y0 ^ f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_15_16_y0;
  assign f_s_dadda_rca24_fa264_y3 = f_s_dadda_rca24_fa264_y0 & f_s_dadda_rca24_fa264_f_s_dadda_rca24_and_15_16_y0;
  assign f_s_dadda_rca24_fa264_y4 = f_s_dadda_rca24_fa264_y1 | f_s_dadda_rca24_fa264_y3;
  assign f_s_dadda_rca24_and_14_17_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_14_17_y0 = f_s_dadda_rca24_and_14_17_a_14 & f_s_dadda_rca24_and_14_17_b_17;
  assign f_s_dadda_rca24_and_13_18_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_13_18_y0 = f_s_dadda_rca24_and_13_18_a_13 & f_s_dadda_rca24_and_13_18_b_18;
  assign f_s_dadda_rca24_and_12_19_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_12_19_y0 = f_s_dadda_rca24_and_12_19_a_12 & f_s_dadda_rca24_and_12_19_b_19;
  assign f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_14_17_y0 = f_s_dadda_rca24_and_14_17_y0;
  assign f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_13_18_y0 = f_s_dadda_rca24_and_13_18_y0;
  assign f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_12_19_y0 = f_s_dadda_rca24_and_12_19_y0;
  assign f_s_dadda_rca24_fa265_y0 = f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_14_17_y0 ^ f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_13_18_y0;
  assign f_s_dadda_rca24_fa265_y1 = f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_14_17_y0 & f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_13_18_y0;
  assign f_s_dadda_rca24_fa265_y2 = f_s_dadda_rca24_fa265_y0 ^ f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_12_19_y0;
  assign f_s_dadda_rca24_fa265_y3 = f_s_dadda_rca24_fa265_y0 & f_s_dadda_rca24_fa265_f_s_dadda_rca24_and_12_19_y0;
  assign f_s_dadda_rca24_fa265_y4 = f_s_dadda_rca24_fa265_y1 | f_s_dadda_rca24_fa265_y3;
  assign f_s_dadda_rca24_and_11_20_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_11_20_y0 = f_s_dadda_rca24_and_11_20_a_11 & f_s_dadda_rca24_and_11_20_b_20;
  assign f_s_dadda_rca24_and_10_21_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_10_21_y0 = f_s_dadda_rca24_and_10_21_a_10 & f_s_dadda_rca24_and_10_21_b_21;
  assign f_s_dadda_rca24_and_9_22_a_9 = a_9;
  assign f_s_dadda_rca24_and_9_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_9_22_y0 = f_s_dadda_rca24_and_9_22_a_9 & f_s_dadda_rca24_and_9_22_b_22;
  assign f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_11_20_y0 = f_s_dadda_rca24_and_11_20_y0;
  assign f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_10_21_y0 = f_s_dadda_rca24_and_10_21_y0;
  assign f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_9_22_y0 = f_s_dadda_rca24_and_9_22_y0;
  assign f_s_dadda_rca24_fa266_y0 = f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_11_20_y0 ^ f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_10_21_y0;
  assign f_s_dadda_rca24_fa266_y1 = f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_11_20_y0 & f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_10_21_y0;
  assign f_s_dadda_rca24_fa266_y2 = f_s_dadda_rca24_fa266_y0 ^ f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_9_22_y0;
  assign f_s_dadda_rca24_fa266_y3 = f_s_dadda_rca24_fa266_y0 & f_s_dadda_rca24_fa266_f_s_dadda_rca24_and_9_22_y0;
  assign f_s_dadda_rca24_fa266_y4 = f_s_dadda_rca24_fa266_y1 | f_s_dadda_rca24_fa266_y3;
  assign f_s_dadda_rca24_nand_8_23_a_8 = a_8;
  assign f_s_dadda_rca24_nand_8_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_8_23_y0 = ~(f_s_dadda_rca24_nand_8_23_a_8 & f_s_dadda_rca24_nand_8_23_b_23);
  assign f_s_dadda_rca24_fa267_f_s_dadda_rca24_nand_8_23_y0 = f_s_dadda_rca24_nand_8_23_y0;
  assign f_s_dadda_rca24_fa267_f_s_dadda_rca24_fa258_y2 = f_s_dadda_rca24_fa258_y2;
  assign f_s_dadda_rca24_fa267_f_s_dadda_rca24_fa259_y2 = f_s_dadda_rca24_fa259_y2;
  assign f_s_dadda_rca24_fa267_y0 = f_s_dadda_rca24_fa267_f_s_dadda_rca24_nand_8_23_y0 ^ f_s_dadda_rca24_fa267_f_s_dadda_rca24_fa258_y2;
  assign f_s_dadda_rca24_fa267_y1 = f_s_dadda_rca24_fa267_f_s_dadda_rca24_nand_8_23_y0 & f_s_dadda_rca24_fa267_f_s_dadda_rca24_fa258_y2;
  assign f_s_dadda_rca24_fa267_y2 = f_s_dadda_rca24_fa267_y0 ^ f_s_dadda_rca24_fa267_f_s_dadda_rca24_fa259_y2;
  assign f_s_dadda_rca24_fa267_y3 = f_s_dadda_rca24_fa267_y0 & f_s_dadda_rca24_fa267_f_s_dadda_rca24_fa259_y2;
  assign f_s_dadda_rca24_fa267_y4 = f_s_dadda_rca24_fa267_y1 | f_s_dadda_rca24_fa267_y3;
  assign f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa260_y2 = f_s_dadda_rca24_fa260_y2;
  assign f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa261_y2 = f_s_dadda_rca24_fa261_y2;
  assign f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa262_y2 = f_s_dadda_rca24_fa262_y2;
  assign f_s_dadda_rca24_fa268_y0 = f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa260_y2 ^ f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa261_y2;
  assign f_s_dadda_rca24_fa268_y1 = f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa260_y2 & f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa261_y2;
  assign f_s_dadda_rca24_fa268_y2 = f_s_dadda_rca24_fa268_y0 ^ f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa262_y2;
  assign f_s_dadda_rca24_fa268_y3 = f_s_dadda_rca24_fa268_y0 & f_s_dadda_rca24_fa268_f_s_dadda_rca24_fa262_y2;
  assign f_s_dadda_rca24_fa268_y4 = f_s_dadda_rca24_fa268_y1 | f_s_dadda_rca24_fa268_y3;
  assign f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa268_y4 = f_s_dadda_rca24_fa268_y4;
  assign f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa267_y4 = f_s_dadda_rca24_fa267_y4;
  assign f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa266_y4 = f_s_dadda_rca24_fa266_y4;
  assign f_s_dadda_rca24_fa269_y0 = f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa268_y4 ^ f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa267_y4;
  assign f_s_dadda_rca24_fa269_y1 = f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa268_y4 & f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa267_y4;
  assign f_s_dadda_rca24_fa269_y2 = f_s_dadda_rca24_fa269_y0 ^ f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa266_y4;
  assign f_s_dadda_rca24_fa269_y3 = f_s_dadda_rca24_fa269_y0 & f_s_dadda_rca24_fa269_f_s_dadda_rca24_fa266_y4;
  assign f_s_dadda_rca24_fa269_y4 = f_s_dadda_rca24_fa269_y1 | f_s_dadda_rca24_fa269_y3;
  assign f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa265_y4 = f_s_dadda_rca24_fa265_y4;
  assign f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa264_y4 = f_s_dadda_rca24_fa264_y4;
  assign f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa263_y4 = f_s_dadda_rca24_fa263_y4;
  assign f_s_dadda_rca24_fa270_y0 = f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa265_y4 ^ f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa264_y4;
  assign f_s_dadda_rca24_fa270_y1 = f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa265_y4 & f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa264_y4;
  assign f_s_dadda_rca24_fa270_y2 = f_s_dadda_rca24_fa270_y0 ^ f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa263_y4;
  assign f_s_dadda_rca24_fa270_y3 = f_s_dadda_rca24_fa270_y0 & f_s_dadda_rca24_fa270_f_s_dadda_rca24_fa263_y4;
  assign f_s_dadda_rca24_fa270_y4 = f_s_dadda_rca24_fa270_y1 | f_s_dadda_rca24_fa270_y3;
  assign f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa262_y4 = f_s_dadda_rca24_fa262_y4;
  assign f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa261_y4 = f_s_dadda_rca24_fa261_y4;
  assign f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa260_y4 = f_s_dadda_rca24_fa260_y4;
  assign f_s_dadda_rca24_fa271_y0 = f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa262_y4 ^ f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa261_y4;
  assign f_s_dadda_rca24_fa271_y1 = f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa262_y4 & f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa261_y4;
  assign f_s_dadda_rca24_fa271_y2 = f_s_dadda_rca24_fa271_y0 ^ f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa260_y4;
  assign f_s_dadda_rca24_fa271_y3 = f_s_dadda_rca24_fa271_y0 & f_s_dadda_rca24_fa271_f_s_dadda_rca24_fa260_y4;
  assign f_s_dadda_rca24_fa271_y4 = f_s_dadda_rca24_fa271_y1 | f_s_dadda_rca24_fa271_y3;
  assign f_s_dadda_rca24_nand_23_9_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_9_b_9 = b_9;
  assign f_s_dadda_rca24_nand_23_9_y0 = ~(f_s_dadda_rca24_nand_23_9_a_23 & f_s_dadda_rca24_nand_23_9_b_9);
  assign f_s_dadda_rca24_fa272_f_s_dadda_rca24_fa259_y4 = f_s_dadda_rca24_fa259_y4;
  assign f_s_dadda_rca24_fa272_f_s_dadda_rca24_fa258_y4 = f_s_dadda_rca24_fa258_y4;
  assign f_s_dadda_rca24_fa272_f_s_dadda_rca24_nand_23_9_y0 = f_s_dadda_rca24_nand_23_9_y0;
  assign f_s_dadda_rca24_fa272_y0 = f_s_dadda_rca24_fa272_f_s_dadda_rca24_fa259_y4 ^ f_s_dadda_rca24_fa272_f_s_dadda_rca24_fa258_y4;
  assign f_s_dadda_rca24_fa272_y1 = f_s_dadda_rca24_fa272_f_s_dadda_rca24_fa259_y4 & f_s_dadda_rca24_fa272_f_s_dadda_rca24_fa258_y4;
  assign f_s_dadda_rca24_fa272_y2 = f_s_dadda_rca24_fa272_y0 ^ f_s_dadda_rca24_fa272_f_s_dadda_rca24_nand_23_9_y0;
  assign f_s_dadda_rca24_fa272_y3 = f_s_dadda_rca24_fa272_y0 & f_s_dadda_rca24_fa272_f_s_dadda_rca24_nand_23_9_y0;
  assign f_s_dadda_rca24_fa272_y4 = f_s_dadda_rca24_fa272_y1 | f_s_dadda_rca24_fa272_y3;
  assign f_s_dadda_rca24_and_22_10_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_22_10_y0 = f_s_dadda_rca24_and_22_10_a_22 & f_s_dadda_rca24_and_22_10_b_10;
  assign f_s_dadda_rca24_and_21_11_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_21_11_y0 = f_s_dadda_rca24_and_21_11_a_21 & f_s_dadda_rca24_and_21_11_b_11;
  assign f_s_dadda_rca24_and_20_12_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_20_12_y0 = f_s_dadda_rca24_and_20_12_a_20 & f_s_dadda_rca24_and_20_12_b_12;
  assign f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_22_10_y0 = f_s_dadda_rca24_and_22_10_y0;
  assign f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_21_11_y0 = f_s_dadda_rca24_and_21_11_y0;
  assign f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_20_12_y0 = f_s_dadda_rca24_and_20_12_y0;
  assign f_s_dadda_rca24_fa273_y0 = f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_22_10_y0 ^ f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_21_11_y0;
  assign f_s_dadda_rca24_fa273_y1 = f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_22_10_y0 & f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_21_11_y0;
  assign f_s_dadda_rca24_fa273_y2 = f_s_dadda_rca24_fa273_y0 ^ f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_20_12_y0;
  assign f_s_dadda_rca24_fa273_y3 = f_s_dadda_rca24_fa273_y0 & f_s_dadda_rca24_fa273_f_s_dadda_rca24_and_20_12_y0;
  assign f_s_dadda_rca24_fa273_y4 = f_s_dadda_rca24_fa273_y1 | f_s_dadda_rca24_fa273_y3;
  assign f_s_dadda_rca24_and_19_13_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_19_13_y0 = f_s_dadda_rca24_and_19_13_a_19 & f_s_dadda_rca24_and_19_13_b_13;
  assign f_s_dadda_rca24_and_18_14_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_18_14_y0 = f_s_dadda_rca24_and_18_14_a_18 & f_s_dadda_rca24_and_18_14_b_14;
  assign f_s_dadda_rca24_and_17_15_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_17_15_y0 = f_s_dadda_rca24_and_17_15_a_17 & f_s_dadda_rca24_and_17_15_b_15;
  assign f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_19_13_y0 = f_s_dadda_rca24_and_19_13_y0;
  assign f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_18_14_y0 = f_s_dadda_rca24_and_18_14_y0;
  assign f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_17_15_y0 = f_s_dadda_rca24_and_17_15_y0;
  assign f_s_dadda_rca24_fa274_y0 = f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_19_13_y0 ^ f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_18_14_y0;
  assign f_s_dadda_rca24_fa274_y1 = f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_19_13_y0 & f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_18_14_y0;
  assign f_s_dadda_rca24_fa274_y2 = f_s_dadda_rca24_fa274_y0 ^ f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_17_15_y0;
  assign f_s_dadda_rca24_fa274_y3 = f_s_dadda_rca24_fa274_y0 & f_s_dadda_rca24_fa274_f_s_dadda_rca24_and_17_15_y0;
  assign f_s_dadda_rca24_fa274_y4 = f_s_dadda_rca24_fa274_y1 | f_s_dadda_rca24_fa274_y3;
  assign f_s_dadda_rca24_and_16_16_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_16_16_y0 = f_s_dadda_rca24_and_16_16_a_16 & f_s_dadda_rca24_and_16_16_b_16;
  assign f_s_dadda_rca24_and_15_17_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_15_17_y0 = f_s_dadda_rca24_and_15_17_a_15 & f_s_dadda_rca24_and_15_17_b_17;
  assign f_s_dadda_rca24_and_14_18_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_14_18_y0 = f_s_dadda_rca24_and_14_18_a_14 & f_s_dadda_rca24_and_14_18_b_18;
  assign f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_16_16_y0 = f_s_dadda_rca24_and_16_16_y0;
  assign f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_15_17_y0 = f_s_dadda_rca24_and_15_17_y0;
  assign f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_14_18_y0 = f_s_dadda_rca24_and_14_18_y0;
  assign f_s_dadda_rca24_fa275_y0 = f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_16_16_y0 ^ f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_15_17_y0;
  assign f_s_dadda_rca24_fa275_y1 = f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_16_16_y0 & f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_15_17_y0;
  assign f_s_dadda_rca24_fa275_y2 = f_s_dadda_rca24_fa275_y0 ^ f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_14_18_y0;
  assign f_s_dadda_rca24_fa275_y3 = f_s_dadda_rca24_fa275_y0 & f_s_dadda_rca24_fa275_f_s_dadda_rca24_and_14_18_y0;
  assign f_s_dadda_rca24_fa275_y4 = f_s_dadda_rca24_fa275_y1 | f_s_dadda_rca24_fa275_y3;
  assign f_s_dadda_rca24_and_13_19_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_13_19_y0 = f_s_dadda_rca24_and_13_19_a_13 & f_s_dadda_rca24_and_13_19_b_19;
  assign f_s_dadda_rca24_and_12_20_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_12_20_y0 = f_s_dadda_rca24_and_12_20_a_12 & f_s_dadda_rca24_and_12_20_b_20;
  assign f_s_dadda_rca24_and_11_21_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_11_21_y0 = f_s_dadda_rca24_and_11_21_a_11 & f_s_dadda_rca24_and_11_21_b_21;
  assign f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_13_19_y0 = f_s_dadda_rca24_and_13_19_y0;
  assign f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_12_20_y0 = f_s_dadda_rca24_and_12_20_y0;
  assign f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_11_21_y0 = f_s_dadda_rca24_and_11_21_y0;
  assign f_s_dadda_rca24_fa276_y0 = f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_13_19_y0 ^ f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_12_20_y0;
  assign f_s_dadda_rca24_fa276_y1 = f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_13_19_y0 & f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_12_20_y0;
  assign f_s_dadda_rca24_fa276_y2 = f_s_dadda_rca24_fa276_y0 ^ f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_11_21_y0;
  assign f_s_dadda_rca24_fa276_y3 = f_s_dadda_rca24_fa276_y0 & f_s_dadda_rca24_fa276_f_s_dadda_rca24_and_11_21_y0;
  assign f_s_dadda_rca24_fa276_y4 = f_s_dadda_rca24_fa276_y1 | f_s_dadda_rca24_fa276_y3;
  assign f_s_dadda_rca24_and_10_22_a_10 = a_10;
  assign f_s_dadda_rca24_and_10_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_10_22_y0 = f_s_dadda_rca24_and_10_22_a_10 & f_s_dadda_rca24_and_10_22_b_22;
  assign f_s_dadda_rca24_nand_9_23_a_9 = a_9;
  assign f_s_dadda_rca24_nand_9_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_9_23_y0 = ~(f_s_dadda_rca24_nand_9_23_a_9 & f_s_dadda_rca24_nand_9_23_b_23);
  assign f_s_dadda_rca24_fa277_f_s_dadda_rca24_and_10_22_y0 = f_s_dadda_rca24_and_10_22_y0;
  assign f_s_dadda_rca24_fa277_f_s_dadda_rca24_nand_9_23_y0 = f_s_dadda_rca24_nand_9_23_y0;
  assign f_s_dadda_rca24_fa277_f_s_dadda_rca24_fa269_y2 = f_s_dadda_rca24_fa269_y2;
  assign f_s_dadda_rca24_fa277_y0 = f_s_dadda_rca24_fa277_f_s_dadda_rca24_and_10_22_y0 ^ f_s_dadda_rca24_fa277_f_s_dadda_rca24_nand_9_23_y0;
  assign f_s_dadda_rca24_fa277_y1 = f_s_dadda_rca24_fa277_f_s_dadda_rca24_and_10_22_y0 & f_s_dadda_rca24_fa277_f_s_dadda_rca24_nand_9_23_y0;
  assign f_s_dadda_rca24_fa277_y2 = f_s_dadda_rca24_fa277_y0 ^ f_s_dadda_rca24_fa277_f_s_dadda_rca24_fa269_y2;
  assign f_s_dadda_rca24_fa277_y3 = f_s_dadda_rca24_fa277_y0 & f_s_dadda_rca24_fa277_f_s_dadda_rca24_fa269_y2;
  assign f_s_dadda_rca24_fa277_y4 = f_s_dadda_rca24_fa277_y1 | f_s_dadda_rca24_fa277_y3;
  assign f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa270_y2 = f_s_dadda_rca24_fa270_y2;
  assign f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa271_y2 = f_s_dadda_rca24_fa271_y2;
  assign f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa272_y2 = f_s_dadda_rca24_fa272_y2;
  assign f_s_dadda_rca24_fa278_y0 = f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa270_y2 ^ f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa271_y2;
  assign f_s_dadda_rca24_fa278_y1 = f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa270_y2 & f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa271_y2;
  assign f_s_dadda_rca24_fa278_y2 = f_s_dadda_rca24_fa278_y0 ^ f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa272_y2;
  assign f_s_dadda_rca24_fa278_y3 = f_s_dadda_rca24_fa278_y0 & f_s_dadda_rca24_fa278_f_s_dadda_rca24_fa272_y2;
  assign f_s_dadda_rca24_fa278_y4 = f_s_dadda_rca24_fa278_y1 | f_s_dadda_rca24_fa278_y3;
  assign f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa278_y4 = f_s_dadda_rca24_fa278_y4;
  assign f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa277_y4 = f_s_dadda_rca24_fa277_y4;
  assign f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa276_y4 = f_s_dadda_rca24_fa276_y4;
  assign f_s_dadda_rca24_fa279_y0 = f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa278_y4 ^ f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa277_y4;
  assign f_s_dadda_rca24_fa279_y1 = f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa278_y4 & f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa277_y4;
  assign f_s_dadda_rca24_fa279_y2 = f_s_dadda_rca24_fa279_y0 ^ f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa276_y4;
  assign f_s_dadda_rca24_fa279_y3 = f_s_dadda_rca24_fa279_y0 & f_s_dadda_rca24_fa279_f_s_dadda_rca24_fa276_y4;
  assign f_s_dadda_rca24_fa279_y4 = f_s_dadda_rca24_fa279_y1 | f_s_dadda_rca24_fa279_y3;
  assign f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa275_y4 = f_s_dadda_rca24_fa275_y4;
  assign f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa274_y4 = f_s_dadda_rca24_fa274_y4;
  assign f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa273_y4 = f_s_dadda_rca24_fa273_y4;
  assign f_s_dadda_rca24_fa280_y0 = f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa275_y4 ^ f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa274_y4;
  assign f_s_dadda_rca24_fa280_y1 = f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa275_y4 & f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa274_y4;
  assign f_s_dadda_rca24_fa280_y2 = f_s_dadda_rca24_fa280_y0 ^ f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa273_y4;
  assign f_s_dadda_rca24_fa280_y3 = f_s_dadda_rca24_fa280_y0 & f_s_dadda_rca24_fa280_f_s_dadda_rca24_fa273_y4;
  assign f_s_dadda_rca24_fa280_y4 = f_s_dadda_rca24_fa280_y1 | f_s_dadda_rca24_fa280_y3;
  assign f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa272_y4 = f_s_dadda_rca24_fa272_y4;
  assign f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa271_y4 = f_s_dadda_rca24_fa271_y4;
  assign f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa270_y4 = f_s_dadda_rca24_fa270_y4;
  assign f_s_dadda_rca24_fa281_y0 = f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa272_y4 ^ f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa271_y4;
  assign f_s_dadda_rca24_fa281_y1 = f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa272_y4 & f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa271_y4;
  assign f_s_dadda_rca24_fa281_y2 = f_s_dadda_rca24_fa281_y0 ^ f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa270_y4;
  assign f_s_dadda_rca24_fa281_y3 = f_s_dadda_rca24_fa281_y0 & f_s_dadda_rca24_fa281_f_s_dadda_rca24_fa270_y4;
  assign f_s_dadda_rca24_fa281_y4 = f_s_dadda_rca24_fa281_y1 | f_s_dadda_rca24_fa281_y3;
  assign f_s_dadda_rca24_nand_23_10_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_10_b_10 = b_10;
  assign f_s_dadda_rca24_nand_23_10_y0 = ~(f_s_dadda_rca24_nand_23_10_a_23 & f_s_dadda_rca24_nand_23_10_b_10);
  assign f_s_dadda_rca24_and_22_11_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_11_b_11 = b_11;
  assign f_s_dadda_rca24_and_22_11_y0 = f_s_dadda_rca24_and_22_11_a_22 & f_s_dadda_rca24_and_22_11_b_11;
  assign f_s_dadda_rca24_fa282_f_s_dadda_rca24_fa269_y4 = f_s_dadda_rca24_fa269_y4;
  assign f_s_dadda_rca24_fa282_f_s_dadda_rca24_nand_23_10_y0 = f_s_dadda_rca24_nand_23_10_y0;
  assign f_s_dadda_rca24_fa282_f_s_dadda_rca24_and_22_11_y0 = f_s_dadda_rca24_and_22_11_y0;
  assign f_s_dadda_rca24_fa282_y0 = f_s_dadda_rca24_fa282_f_s_dadda_rca24_fa269_y4 ^ f_s_dadda_rca24_fa282_f_s_dadda_rca24_nand_23_10_y0;
  assign f_s_dadda_rca24_fa282_y1 = f_s_dadda_rca24_fa282_f_s_dadda_rca24_fa269_y4 & f_s_dadda_rca24_fa282_f_s_dadda_rca24_nand_23_10_y0;
  assign f_s_dadda_rca24_fa282_y2 = f_s_dadda_rca24_fa282_y0 ^ f_s_dadda_rca24_fa282_f_s_dadda_rca24_and_22_11_y0;
  assign f_s_dadda_rca24_fa282_y3 = f_s_dadda_rca24_fa282_y0 & f_s_dadda_rca24_fa282_f_s_dadda_rca24_and_22_11_y0;
  assign f_s_dadda_rca24_fa282_y4 = f_s_dadda_rca24_fa282_y1 | f_s_dadda_rca24_fa282_y3;
  assign f_s_dadda_rca24_and_21_12_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_21_12_y0 = f_s_dadda_rca24_and_21_12_a_21 & f_s_dadda_rca24_and_21_12_b_12;
  assign f_s_dadda_rca24_and_20_13_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_20_13_y0 = f_s_dadda_rca24_and_20_13_a_20 & f_s_dadda_rca24_and_20_13_b_13;
  assign f_s_dadda_rca24_and_19_14_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_19_14_y0 = f_s_dadda_rca24_and_19_14_a_19 & f_s_dadda_rca24_and_19_14_b_14;
  assign f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_21_12_y0 = f_s_dadda_rca24_and_21_12_y0;
  assign f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_20_13_y0 = f_s_dadda_rca24_and_20_13_y0;
  assign f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_19_14_y0 = f_s_dadda_rca24_and_19_14_y0;
  assign f_s_dadda_rca24_fa283_y0 = f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_21_12_y0 ^ f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_20_13_y0;
  assign f_s_dadda_rca24_fa283_y1 = f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_21_12_y0 & f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_20_13_y0;
  assign f_s_dadda_rca24_fa283_y2 = f_s_dadda_rca24_fa283_y0 ^ f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_19_14_y0;
  assign f_s_dadda_rca24_fa283_y3 = f_s_dadda_rca24_fa283_y0 & f_s_dadda_rca24_fa283_f_s_dadda_rca24_and_19_14_y0;
  assign f_s_dadda_rca24_fa283_y4 = f_s_dadda_rca24_fa283_y1 | f_s_dadda_rca24_fa283_y3;
  assign f_s_dadda_rca24_and_18_15_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_18_15_y0 = f_s_dadda_rca24_and_18_15_a_18 & f_s_dadda_rca24_and_18_15_b_15;
  assign f_s_dadda_rca24_and_17_16_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_17_16_y0 = f_s_dadda_rca24_and_17_16_a_17 & f_s_dadda_rca24_and_17_16_b_16;
  assign f_s_dadda_rca24_and_16_17_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_16_17_y0 = f_s_dadda_rca24_and_16_17_a_16 & f_s_dadda_rca24_and_16_17_b_17;
  assign f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_18_15_y0 = f_s_dadda_rca24_and_18_15_y0;
  assign f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_17_16_y0 = f_s_dadda_rca24_and_17_16_y0;
  assign f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_16_17_y0 = f_s_dadda_rca24_and_16_17_y0;
  assign f_s_dadda_rca24_fa284_y0 = f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_18_15_y0 ^ f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_17_16_y0;
  assign f_s_dadda_rca24_fa284_y1 = f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_18_15_y0 & f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_17_16_y0;
  assign f_s_dadda_rca24_fa284_y2 = f_s_dadda_rca24_fa284_y0 ^ f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_16_17_y0;
  assign f_s_dadda_rca24_fa284_y3 = f_s_dadda_rca24_fa284_y0 & f_s_dadda_rca24_fa284_f_s_dadda_rca24_and_16_17_y0;
  assign f_s_dadda_rca24_fa284_y4 = f_s_dadda_rca24_fa284_y1 | f_s_dadda_rca24_fa284_y3;
  assign f_s_dadda_rca24_and_15_18_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_15_18_y0 = f_s_dadda_rca24_and_15_18_a_15 & f_s_dadda_rca24_and_15_18_b_18;
  assign f_s_dadda_rca24_and_14_19_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_14_19_y0 = f_s_dadda_rca24_and_14_19_a_14 & f_s_dadda_rca24_and_14_19_b_19;
  assign f_s_dadda_rca24_and_13_20_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_13_20_y0 = f_s_dadda_rca24_and_13_20_a_13 & f_s_dadda_rca24_and_13_20_b_20;
  assign f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_15_18_y0 = f_s_dadda_rca24_and_15_18_y0;
  assign f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_14_19_y0 = f_s_dadda_rca24_and_14_19_y0;
  assign f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_13_20_y0 = f_s_dadda_rca24_and_13_20_y0;
  assign f_s_dadda_rca24_fa285_y0 = f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_15_18_y0 ^ f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_14_19_y0;
  assign f_s_dadda_rca24_fa285_y1 = f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_15_18_y0 & f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_14_19_y0;
  assign f_s_dadda_rca24_fa285_y2 = f_s_dadda_rca24_fa285_y0 ^ f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_13_20_y0;
  assign f_s_dadda_rca24_fa285_y3 = f_s_dadda_rca24_fa285_y0 & f_s_dadda_rca24_fa285_f_s_dadda_rca24_and_13_20_y0;
  assign f_s_dadda_rca24_fa285_y4 = f_s_dadda_rca24_fa285_y1 | f_s_dadda_rca24_fa285_y3;
  assign f_s_dadda_rca24_and_12_21_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_12_21_y0 = f_s_dadda_rca24_and_12_21_a_12 & f_s_dadda_rca24_and_12_21_b_21;
  assign f_s_dadda_rca24_and_11_22_a_11 = a_11;
  assign f_s_dadda_rca24_and_11_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_11_22_y0 = f_s_dadda_rca24_and_11_22_a_11 & f_s_dadda_rca24_and_11_22_b_22;
  assign f_s_dadda_rca24_nand_10_23_a_10 = a_10;
  assign f_s_dadda_rca24_nand_10_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_10_23_y0 = ~(f_s_dadda_rca24_nand_10_23_a_10 & f_s_dadda_rca24_nand_10_23_b_23);
  assign f_s_dadda_rca24_fa286_f_s_dadda_rca24_and_12_21_y0 = f_s_dadda_rca24_and_12_21_y0;
  assign f_s_dadda_rca24_fa286_f_s_dadda_rca24_and_11_22_y0 = f_s_dadda_rca24_and_11_22_y0;
  assign f_s_dadda_rca24_fa286_f_s_dadda_rca24_nand_10_23_y0 = f_s_dadda_rca24_nand_10_23_y0;
  assign f_s_dadda_rca24_fa286_y0 = f_s_dadda_rca24_fa286_f_s_dadda_rca24_and_12_21_y0 ^ f_s_dadda_rca24_fa286_f_s_dadda_rca24_and_11_22_y0;
  assign f_s_dadda_rca24_fa286_y1 = f_s_dadda_rca24_fa286_f_s_dadda_rca24_and_12_21_y0 & f_s_dadda_rca24_fa286_f_s_dadda_rca24_and_11_22_y0;
  assign f_s_dadda_rca24_fa286_y2 = f_s_dadda_rca24_fa286_y0 ^ f_s_dadda_rca24_fa286_f_s_dadda_rca24_nand_10_23_y0;
  assign f_s_dadda_rca24_fa286_y3 = f_s_dadda_rca24_fa286_y0 & f_s_dadda_rca24_fa286_f_s_dadda_rca24_nand_10_23_y0;
  assign f_s_dadda_rca24_fa286_y4 = f_s_dadda_rca24_fa286_y1 | f_s_dadda_rca24_fa286_y3;
  assign f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa279_y2 = f_s_dadda_rca24_fa279_y2;
  assign f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa280_y2 = f_s_dadda_rca24_fa280_y2;
  assign f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa281_y2 = f_s_dadda_rca24_fa281_y2;
  assign f_s_dadda_rca24_fa287_y0 = f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa279_y2 ^ f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa280_y2;
  assign f_s_dadda_rca24_fa287_y1 = f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa279_y2 & f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa280_y2;
  assign f_s_dadda_rca24_fa287_y2 = f_s_dadda_rca24_fa287_y0 ^ f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa281_y2;
  assign f_s_dadda_rca24_fa287_y3 = f_s_dadda_rca24_fa287_y0 & f_s_dadda_rca24_fa287_f_s_dadda_rca24_fa281_y2;
  assign f_s_dadda_rca24_fa287_y4 = f_s_dadda_rca24_fa287_y1 | f_s_dadda_rca24_fa287_y3;
  assign f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa287_y4 = f_s_dadda_rca24_fa287_y4;
  assign f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa286_y4 = f_s_dadda_rca24_fa286_y4;
  assign f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa285_y4 = f_s_dadda_rca24_fa285_y4;
  assign f_s_dadda_rca24_fa288_y0 = f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa287_y4 ^ f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa286_y4;
  assign f_s_dadda_rca24_fa288_y1 = f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa287_y4 & f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa286_y4;
  assign f_s_dadda_rca24_fa288_y2 = f_s_dadda_rca24_fa288_y0 ^ f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa285_y4;
  assign f_s_dadda_rca24_fa288_y3 = f_s_dadda_rca24_fa288_y0 & f_s_dadda_rca24_fa288_f_s_dadda_rca24_fa285_y4;
  assign f_s_dadda_rca24_fa288_y4 = f_s_dadda_rca24_fa288_y1 | f_s_dadda_rca24_fa288_y3;
  assign f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa284_y4 = f_s_dadda_rca24_fa284_y4;
  assign f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa283_y4 = f_s_dadda_rca24_fa283_y4;
  assign f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa282_y4 = f_s_dadda_rca24_fa282_y4;
  assign f_s_dadda_rca24_fa289_y0 = f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa284_y4 ^ f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa283_y4;
  assign f_s_dadda_rca24_fa289_y1 = f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa284_y4 & f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa283_y4;
  assign f_s_dadda_rca24_fa289_y2 = f_s_dadda_rca24_fa289_y0 ^ f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa282_y4;
  assign f_s_dadda_rca24_fa289_y3 = f_s_dadda_rca24_fa289_y0 & f_s_dadda_rca24_fa289_f_s_dadda_rca24_fa282_y4;
  assign f_s_dadda_rca24_fa289_y4 = f_s_dadda_rca24_fa289_y1 | f_s_dadda_rca24_fa289_y3;
  assign f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa281_y4 = f_s_dadda_rca24_fa281_y4;
  assign f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa280_y4 = f_s_dadda_rca24_fa280_y4;
  assign f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa279_y4 = f_s_dadda_rca24_fa279_y4;
  assign f_s_dadda_rca24_fa290_y0 = f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa281_y4 ^ f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa280_y4;
  assign f_s_dadda_rca24_fa290_y1 = f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa281_y4 & f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa280_y4;
  assign f_s_dadda_rca24_fa290_y2 = f_s_dadda_rca24_fa290_y0 ^ f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa279_y4;
  assign f_s_dadda_rca24_fa290_y3 = f_s_dadda_rca24_fa290_y0 & f_s_dadda_rca24_fa290_f_s_dadda_rca24_fa279_y4;
  assign f_s_dadda_rca24_fa290_y4 = f_s_dadda_rca24_fa290_y1 | f_s_dadda_rca24_fa290_y3;
  assign f_s_dadda_rca24_nand_23_11_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_11_b_11 = b_11;
  assign f_s_dadda_rca24_nand_23_11_y0 = ~(f_s_dadda_rca24_nand_23_11_a_23 & f_s_dadda_rca24_nand_23_11_b_11);
  assign f_s_dadda_rca24_and_22_12_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_12_b_12 = b_12;
  assign f_s_dadda_rca24_and_22_12_y0 = f_s_dadda_rca24_and_22_12_a_22 & f_s_dadda_rca24_and_22_12_b_12;
  assign f_s_dadda_rca24_and_21_13_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_21_13_y0 = f_s_dadda_rca24_and_21_13_a_21 & f_s_dadda_rca24_and_21_13_b_13;
  assign f_s_dadda_rca24_fa291_f_s_dadda_rca24_nand_23_11_y0 = f_s_dadda_rca24_nand_23_11_y0;
  assign f_s_dadda_rca24_fa291_f_s_dadda_rca24_and_22_12_y0 = f_s_dadda_rca24_and_22_12_y0;
  assign f_s_dadda_rca24_fa291_f_s_dadda_rca24_and_21_13_y0 = f_s_dadda_rca24_and_21_13_y0;
  assign f_s_dadda_rca24_fa291_y0 = f_s_dadda_rca24_fa291_f_s_dadda_rca24_nand_23_11_y0 ^ f_s_dadda_rca24_fa291_f_s_dadda_rca24_and_22_12_y0;
  assign f_s_dadda_rca24_fa291_y1 = f_s_dadda_rca24_fa291_f_s_dadda_rca24_nand_23_11_y0 & f_s_dadda_rca24_fa291_f_s_dadda_rca24_and_22_12_y0;
  assign f_s_dadda_rca24_fa291_y2 = f_s_dadda_rca24_fa291_y0 ^ f_s_dadda_rca24_fa291_f_s_dadda_rca24_and_21_13_y0;
  assign f_s_dadda_rca24_fa291_y3 = f_s_dadda_rca24_fa291_y0 & f_s_dadda_rca24_fa291_f_s_dadda_rca24_and_21_13_y0;
  assign f_s_dadda_rca24_fa291_y4 = f_s_dadda_rca24_fa291_y1 | f_s_dadda_rca24_fa291_y3;
  assign f_s_dadda_rca24_and_20_14_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_20_14_y0 = f_s_dadda_rca24_and_20_14_a_20 & f_s_dadda_rca24_and_20_14_b_14;
  assign f_s_dadda_rca24_and_19_15_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_19_15_y0 = f_s_dadda_rca24_and_19_15_a_19 & f_s_dadda_rca24_and_19_15_b_15;
  assign f_s_dadda_rca24_and_18_16_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_18_16_y0 = f_s_dadda_rca24_and_18_16_a_18 & f_s_dadda_rca24_and_18_16_b_16;
  assign f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_20_14_y0 = f_s_dadda_rca24_and_20_14_y0;
  assign f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_19_15_y0 = f_s_dadda_rca24_and_19_15_y0;
  assign f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_18_16_y0 = f_s_dadda_rca24_and_18_16_y0;
  assign f_s_dadda_rca24_fa292_y0 = f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_20_14_y0 ^ f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_19_15_y0;
  assign f_s_dadda_rca24_fa292_y1 = f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_20_14_y0 & f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_19_15_y0;
  assign f_s_dadda_rca24_fa292_y2 = f_s_dadda_rca24_fa292_y0 ^ f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_18_16_y0;
  assign f_s_dadda_rca24_fa292_y3 = f_s_dadda_rca24_fa292_y0 & f_s_dadda_rca24_fa292_f_s_dadda_rca24_and_18_16_y0;
  assign f_s_dadda_rca24_fa292_y4 = f_s_dadda_rca24_fa292_y1 | f_s_dadda_rca24_fa292_y3;
  assign f_s_dadda_rca24_and_17_17_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_17_17_y0 = f_s_dadda_rca24_and_17_17_a_17 & f_s_dadda_rca24_and_17_17_b_17;
  assign f_s_dadda_rca24_and_16_18_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_16_18_y0 = f_s_dadda_rca24_and_16_18_a_16 & f_s_dadda_rca24_and_16_18_b_18;
  assign f_s_dadda_rca24_and_15_19_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_15_19_y0 = f_s_dadda_rca24_and_15_19_a_15 & f_s_dadda_rca24_and_15_19_b_19;
  assign f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_17_17_y0 = f_s_dadda_rca24_and_17_17_y0;
  assign f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_16_18_y0 = f_s_dadda_rca24_and_16_18_y0;
  assign f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_15_19_y0 = f_s_dadda_rca24_and_15_19_y0;
  assign f_s_dadda_rca24_fa293_y0 = f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_17_17_y0 ^ f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_16_18_y0;
  assign f_s_dadda_rca24_fa293_y1 = f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_17_17_y0 & f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_16_18_y0;
  assign f_s_dadda_rca24_fa293_y2 = f_s_dadda_rca24_fa293_y0 ^ f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_15_19_y0;
  assign f_s_dadda_rca24_fa293_y3 = f_s_dadda_rca24_fa293_y0 & f_s_dadda_rca24_fa293_f_s_dadda_rca24_and_15_19_y0;
  assign f_s_dadda_rca24_fa293_y4 = f_s_dadda_rca24_fa293_y1 | f_s_dadda_rca24_fa293_y3;
  assign f_s_dadda_rca24_and_14_20_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_14_20_y0 = f_s_dadda_rca24_and_14_20_a_14 & f_s_dadda_rca24_and_14_20_b_20;
  assign f_s_dadda_rca24_and_13_21_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_13_21_y0 = f_s_dadda_rca24_and_13_21_a_13 & f_s_dadda_rca24_and_13_21_b_21;
  assign f_s_dadda_rca24_and_12_22_a_12 = a_12;
  assign f_s_dadda_rca24_and_12_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_12_22_y0 = f_s_dadda_rca24_and_12_22_a_12 & f_s_dadda_rca24_and_12_22_b_22;
  assign f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_14_20_y0 = f_s_dadda_rca24_and_14_20_y0;
  assign f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_13_21_y0 = f_s_dadda_rca24_and_13_21_y0;
  assign f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_12_22_y0 = f_s_dadda_rca24_and_12_22_y0;
  assign f_s_dadda_rca24_fa294_y0 = f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_14_20_y0 ^ f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_13_21_y0;
  assign f_s_dadda_rca24_fa294_y1 = f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_14_20_y0 & f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_13_21_y0;
  assign f_s_dadda_rca24_fa294_y2 = f_s_dadda_rca24_fa294_y0 ^ f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_12_22_y0;
  assign f_s_dadda_rca24_fa294_y3 = f_s_dadda_rca24_fa294_y0 & f_s_dadda_rca24_fa294_f_s_dadda_rca24_and_12_22_y0;
  assign f_s_dadda_rca24_fa294_y4 = f_s_dadda_rca24_fa294_y1 | f_s_dadda_rca24_fa294_y3;
  assign f_s_dadda_rca24_nand_11_23_a_11 = a_11;
  assign f_s_dadda_rca24_nand_11_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_11_23_y0 = ~(f_s_dadda_rca24_nand_11_23_a_11 & f_s_dadda_rca24_nand_11_23_b_23);
  assign f_s_dadda_rca24_fa295_f_s_dadda_rca24_nand_11_23_y0 = f_s_dadda_rca24_nand_11_23_y0;
  assign f_s_dadda_rca24_fa295_f_s_dadda_rca24_fa288_y2 = f_s_dadda_rca24_fa288_y2;
  assign f_s_dadda_rca24_fa295_f_s_dadda_rca24_fa289_y2 = f_s_dadda_rca24_fa289_y2;
  assign f_s_dadda_rca24_fa295_y0 = f_s_dadda_rca24_fa295_f_s_dadda_rca24_nand_11_23_y0 ^ f_s_dadda_rca24_fa295_f_s_dadda_rca24_fa288_y2;
  assign f_s_dadda_rca24_fa295_y1 = f_s_dadda_rca24_fa295_f_s_dadda_rca24_nand_11_23_y0 & f_s_dadda_rca24_fa295_f_s_dadda_rca24_fa288_y2;
  assign f_s_dadda_rca24_fa295_y2 = f_s_dadda_rca24_fa295_y0 ^ f_s_dadda_rca24_fa295_f_s_dadda_rca24_fa289_y2;
  assign f_s_dadda_rca24_fa295_y3 = f_s_dadda_rca24_fa295_y0 & f_s_dadda_rca24_fa295_f_s_dadda_rca24_fa289_y2;
  assign f_s_dadda_rca24_fa295_y4 = f_s_dadda_rca24_fa295_y1 | f_s_dadda_rca24_fa295_y3;
  assign f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa295_y4 = f_s_dadda_rca24_fa295_y4;
  assign f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa294_y4 = f_s_dadda_rca24_fa294_y4;
  assign f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa293_y4 = f_s_dadda_rca24_fa293_y4;
  assign f_s_dadda_rca24_fa296_y0 = f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa295_y4 ^ f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa294_y4;
  assign f_s_dadda_rca24_fa296_y1 = f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa295_y4 & f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa294_y4;
  assign f_s_dadda_rca24_fa296_y2 = f_s_dadda_rca24_fa296_y0 ^ f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa293_y4;
  assign f_s_dadda_rca24_fa296_y3 = f_s_dadda_rca24_fa296_y0 & f_s_dadda_rca24_fa296_f_s_dadda_rca24_fa293_y4;
  assign f_s_dadda_rca24_fa296_y4 = f_s_dadda_rca24_fa296_y1 | f_s_dadda_rca24_fa296_y3;
  assign f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa292_y4 = f_s_dadda_rca24_fa292_y4;
  assign f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa291_y4 = f_s_dadda_rca24_fa291_y4;
  assign f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa290_y4 = f_s_dadda_rca24_fa290_y4;
  assign f_s_dadda_rca24_fa297_y0 = f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa292_y4 ^ f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa291_y4;
  assign f_s_dadda_rca24_fa297_y1 = f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa292_y4 & f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa291_y4;
  assign f_s_dadda_rca24_fa297_y2 = f_s_dadda_rca24_fa297_y0 ^ f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa290_y4;
  assign f_s_dadda_rca24_fa297_y3 = f_s_dadda_rca24_fa297_y0 & f_s_dadda_rca24_fa297_f_s_dadda_rca24_fa290_y4;
  assign f_s_dadda_rca24_fa297_y4 = f_s_dadda_rca24_fa297_y1 | f_s_dadda_rca24_fa297_y3;
  assign f_s_dadda_rca24_nand_23_12_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_12_b_12 = b_12;
  assign f_s_dadda_rca24_nand_23_12_y0 = ~(f_s_dadda_rca24_nand_23_12_a_23 & f_s_dadda_rca24_nand_23_12_b_12);
  assign f_s_dadda_rca24_fa298_f_s_dadda_rca24_fa289_y4 = f_s_dadda_rca24_fa289_y4;
  assign f_s_dadda_rca24_fa298_f_s_dadda_rca24_fa288_y4 = f_s_dadda_rca24_fa288_y4;
  assign f_s_dadda_rca24_fa298_f_s_dadda_rca24_nand_23_12_y0 = f_s_dadda_rca24_nand_23_12_y0;
  assign f_s_dadda_rca24_fa298_y0 = f_s_dadda_rca24_fa298_f_s_dadda_rca24_fa289_y4 ^ f_s_dadda_rca24_fa298_f_s_dadda_rca24_fa288_y4;
  assign f_s_dadda_rca24_fa298_y1 = f_s_dadda_rca24_fa298_f_s_dadda_rca24_fa289_y4 & f_s_dadda_rca24_fa298_f_s_dadda_rca24_fa288_y4;
  assign f_s_dadda_rca24_fa298_y2 = f_s_dadda_rca24_fa298_y0 ^ f_s_dadda_rca24_fa298_f_s_dadda_rca24_nand_23_12_y0;
  assign f_s_dadda_rca24_fa298_y3 = f_s_dadda_rca24_fa298_y0 & f_s_dadda_rca24_fa298_f_s_dadda_rca24_nand_23_12_y0;
  assign f_s_dadda_rca24_fa298_y4 = f_s_dadda_rca24_fa298_y1 | f_s_dadda_rca24_fa298_y3;
  assign f_s_dadda_rca24_and_22_13_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_13_b_13 = b_13;
  assign f_s_dadda_rca24_and_22_13_y0 = f_s_dadda_rca24_and_22_13_a_22 & f_s_dadda_rca24_and_22_13_b_13;
  assign f_s_dadda_rca24_and_21_14_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_21_14_y0 = f_s_dadda_rca24_and_21_14_a_21 & f_s_dadda_rca24_and_21_14_b_14;
  assign f_s_dadda_rca24_and_20_15_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_20_15_y0 = f_s_dadda_rca24_and_20_15_a_20 & f_s_dadda_rca24_and_20_15_b_15;
  assign f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_22_13_y0 = f_s_dadda_rca24_and_22_13_y0;
  assign f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_21_14_y0 = f_s_dadda_rca24_and_21_14_y0;
  assign f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_20_15_y0 = f_s_dadda_rca24_and_20_15_y0;
  assign f_s_dadda_rca24_fa299_y0 = f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_22_13_y0 ^ f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_21_14_y0;
  assign f_s_dadda_rca24_fa299_y1 = f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_22_13_y0 & f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_21_14_y0;
  assign f_s_dadda_rca24_fa299_y2 = f_s_dadda_rca24_fa299_y0 ^ f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_20_15_y0;
  assign f_s_dadda_rca24_fa299_y3 = f_s_dadda_rca24_fa299_y0 & f_s_dadda_rca24_fa299_f_s_dadda_rca24_and_20_15_y0;
  assign f_s_dadda_rca24_fa299_y4 = f_s_dadda_rca24_fa299_y1 | f_s_dadda_rca24_fa299_y3;
  assign f_s_dadda_rca24_and_19_16_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_19_16_y0 = f_s_dadda_rca24_and_19_16_a_19 & f_s_dadda_rca24_and_19_16_b_16;
  assign f_s_dadda_rca24_and_18_17_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_18_17_y0 = f_s_dadda_rca24_and_18_17_a_18 & f_s_dadda_rca24_and_18_17_b_17;
  assign f_s_dadda_rca24_and_17_18_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_17_18_y0 = f_s_dadda_rca24_and_17_18_a_17 & f_s_dadda_rca24_and_17_18_b_18;
  assign f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_19_16_y0 = f_s_dadda_rca24_and_19_16_y0;
  assign f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_18_17_y0 = f_s_dadda_rca24_and_18_17_y0;
  assign f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_17_18_y0 = f_s_dadda_rca24_and_17_18_y0;
  assign f_s_dadda_rca24_fa300_y0 = f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_19_16_y0 ^ f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_18_17_y0;
  assign f_s_dadda_rca24_fa300_y1 = f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_19_16_y0 & f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_18_17_y0;
  assign f_s_dadda_rca24_fa300_y2 = f_s_dadda_rca24_fa300_y0 ^ f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_17_18_y0;
  assign f_s_dadda_rca24_fa300_y3 = f_s_dadda_rca24_fa300_y0 & f_s_dadda_rca24_fa300_f_s_dadda_rca24_and_17_18_y0;
  assign f_s_dadda_rca24_fa300_y4 = f_s_dadda_rca24_fa300_y1 | f_s_dadda_rca24_fa300_y3;
  assign f_s_dadda_rca24_and_16_19_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_16_19_y0 = f_s_dadda_rca24_and_16_19_a_16 & f_s_dadda_rca24_and_16_19_b_19;
  assign f_s_dadda_rca24_and_15_20_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_15_20_y0 = f_s_dadda_rca24_and_15_20_a_15 & f_s_dadda_rca24_and_15_20_b_20;
  assign f_s_dadda_rca24_and_14_21_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_14_21_y0 = f_s_dadda_rca24_and_14_21_a_14 & f_s_dadda_rca24_and_14_21_b_21;
  assign f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_16_19_y0 = f_s_dadda_rca24_and_16_19_y0;
  assign f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_15_20_y0 = f_s_dadda_rca24_and_15_20_y0;
  assign f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_14_21_y0 = f_s_dadda_rca24_and_14_21_y0;
  assign f_s_dadda_rca24_fa301_y0 = f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_16_19_y0 ^ f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_15_20_y0;
  assign f_s_dadda_rca24_fa301_y1 = f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_16_19_y0 & f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_15_20_y0;
  assign f_s_dadda_rca24_fa301_y2 = f_s_dadda_rca24_fa301_y0 ^ f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_14_21_y0;
  assign f_s_dadda_rca24_fa301_y3 = f_s_dadda_rca24_fa301_y0 & f_s_dadda_rca24_fa301_f_s_dadda_rca24_and_14_21_y0;
  assign f_s_dadda_rca24_fa301_y4 = f_s_dadda_rca24_fa301_y1 | f_s_dadda_rca24_fa301_y3;
  assign f_s_dadda_rca24_and_13_22_a_13 = a_13;
  assign f_s_dadda_rca24_and_13_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_13_22_y0 = f_s_dadda_rca24_and_13_22_a_13 & f_s_dadda_rca24_and_13_22_b_22;
  assign f_s_dadda_rca24_nand_12_23_a_12 = a_12;
  assign f_s_dadda_rca24_nand_12_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_12_23_y0 = ~(f_s_dadda_rca24_nand_12_23_a_12 & f_s_dadda_rca24_nand_12_23_b_23);
  assign f_s_dadda_rca24_fa302_f_s_dadda_rca24_and_13_22_y0 = f_s_dadda_rca24_and_13_22_y0;
  assign f_s_dadda_rca24_fa302_f_s_dadda_rca24_nand_12_23_y0 = f_s_dadda_rca24_nand_12_23_y0;
  assign f_s_dadda_rca24_fa302_f_s_dadda_rca24_fa296_y2 = f_s_dadda_rca24_fa296_y2;
  assign f_s_dadda_rca24_fa302_y0 = f_s_dadda_rca24_fa302_f_s_dadda_rca24_and_13_22_y0 ^ f_s_dadda_rca24_fa302_f_s_dadda_rca24_nand_12_23_y0;
  assign f_s_dadda_rca24_fa302_y1 = f_s_dadda_rca24_fa302_f_s_dadda_rca24_and_13_22_y0 & f_s_dadda_rca24_fa302_f_s_dadda_rca24_nand_12_23_y0;
  assign f_s_dadda_rca24_fa302_y2 = f_s_dadda_rca24_fa302_y0 ^ f_s_dadda_rca24_fa302_f_s_dadda_rca24_fa296_y2;
  assign f_s_dadda_rca24_fa302_y3 = f_s_dadda_rca24_fa302_y0 & f_s_dadda_rca24_fa302_f_s_dadda_rca24_fa296_y2;
  assign f_s_dadda_rca24_fa302_y4 = f_s_dadda_rca24_fa302_y1 | f_s_dadda_rca24_fa302_y3;
  assign f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa302_y4 = f_s_dadda_rca24_fa302_y4;
  assign f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa301_y4 = f_s_dadda_rca24_fa301_y4;
  assign f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa300_y4 = f_s_dadda_rca24_fa300_y4;
  assign f_s_dadda_rca24_fa303_y0 = f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa302_y4 ^ f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa301_y4;
  assign f_s_dadda_rca24_fa303_y1 = f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa302_y4 & f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa301_y4;
  assign f_s_dadda_rca24_fa303_y2 = f_s_dadda_rca24_fa303_y0 ^ f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa300_y4;
  assign f_s_dadda_rca24_fa303_y3 = f_s_dadda_rca24_fa303_y0 & f_s_dadda_rca24_fa303_f_s_dadda_rca24_fa300_y4;
  assign f_s_dadda_rca24_fa303_y4 = f_s_dadda_rca24_fa303_y1 | f_s_dadda_rca24_fa303_y3;
  assign f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa299_y4 = f_s_dadda_rca24_fa299_y4;
  assign f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa298_y4 = f_s_dadda_rca24_fa298_y4;
  assign f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa297_y4 = f_s_dadda_rca24_fa297_y4;
  assign f_s_dadda_rca24_fa304_y0 = f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa299_y4 ^ f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa298_y4;
  assign f_s_dadda_rca24_fa304_y1 = f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa299_y4 & f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa298_y4;
  assign f_s_dadda_rca24_fa304_y2 = f_s_dadda_rca24_fa304_y0 ^ f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa297_y4;
  assign f_s_dadda_rca24_fa304_y3 = f_s_dadda_rca24_fa304_y0 & f_s_dadda_rca24_fa304_f_s_dadda_rca24_fa297_y4;
  assign f_s_dadda_rca24_fa304_y4 = f_s_dadda_rca24_fa304_y1 | f_s_dadda_rca24_fa304_y3;
  assign f_s_dadda_rca24_nand_23_13_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_13_b_13 = b_13;
  assign f_s_dadda_rca24_nand_23_13_y0 = ~(f_s_dadda_rca24_nand_23_13_a_23 & f_s_dadda_rca24_nand_23_13_b_13);
  assign f_s_dadda_rca24_and_22_14_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_14_b_14 = b_14;
  assign f_s_dadda_rca24_and_22_14_y0 = f_s_dadda_rca24_and_22_14_a_22 & f_s_dadda_rca24_and_22_14_b_14;
  assign f_s_dadda_rca24_fa305_f_s_dadda_rca24_fa296_y4 = f_s_dadda_rca24_fa296_y4;
  assign f_s_dadda_rca24_fa305_f_s_dadda_rca24_nand_23_13_y0 = f_s_dadda_rca24_nand_23_13_y0;
  assign f_s_dadda_rca24_fa305_f_s_dadda_rca24_and_22_14_y0 = f_s_dadda_rca24_and_22_14_y0;
  assign f_s_dadda_rca24_fa305_y0 = f_s_dadda_rca24_fa305_f_s_dadda_rca24_fa296_y4 ^ f_s_dadda_rca24_fa305_f_s_dadda_rca24_nand_23_13_y0;
  assign f_s_dadda_rca24_fa305_y1 = f_s_dadda_rca24_fa305_f_s_dadda_rca24_fa296_y4 & f_s_dadda_rca24_fa305_f_s_dadda_rca24_nand_23_13_y0;
  assign f_s_dadda_rca24_fa305_y2 = f_s_dadda_rca24_fa305_y0 ^ f_s_dadda_rca24_fa305_f_s_dadda_rca24_and_22_14_y0;
  assign f_s_dadda_rca24_fa305_y3 = f_s_dadda_rca24_fa305_y0 & f_s_dadda_rca24_fa305_f_s_dadda_rca24_and_22_14_y0;
  assign f_s_dadda_rca24_fa305_y4 = f_s_dadda_rca24_fa305_y1 | f_s_dadda_rca24_fa305_y3;
  assign f_s_dadda_rca24_and_21_15_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_21_15_y0 = f_s_dadda_rca24_and_21_15_a_21 & f_s_dadda_rca24_and_21_15_b_15;
  assign f_s_dadda_rca24_and_20_16_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_20_16_y0 = f_s_dadda_rca24_and_20_16_a_20 & f_s_dadda_rca24_and_20_16_b_16;
  assign f_s_dadda_rca24_and_19_17_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_19_17_y0 = f_s_dadda_rca24_and_19_17_a_19 & f_s_dadda_rca24_and_19_17_b_17;
  assign f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_21_15_y0 = f_s_dadda_rca24_and_21_15_y0;
  assign f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_20_16_y0 = f_s_dadda_rca24_and_20_16_y0;
  assign f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_19_17_y0 = f_s_dadda_rca24_and_19_17_y0;
  assign f_s_dadda_rca24_fa306_y0 = f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_21_15_y0 ^ f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_20_16_y0;
  assign f_s_dadda_rca24_fa306_y1 = f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_21_15_y0 & f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_20_16_y0;
  assign f_s_dadda_rca24_fa306_y2 = f_s_dadda_rca24_fa306_y0 ^ f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_19_17_y0;
  assign f_s_dadda_rca24_fa306_y3 = f_s_dadda_rca24_fa306_y0 & f_s_dadda_rca24_fa306_f_s_dadda_rca24_and_19_17_y0;
  assign f_s_dadda_rca24_fa306_y4 = f_s_dadda_rca24_fa306_y1 | f_s_dadda_rca24_fa306_y3;
  assign f_s_dadda_rca24_and_18_18_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_18_18_y0 = f_s_dadda_rca24_and_18_18_a_18 & f_s_dadda_rca24_and_18_18_b_18;
  assign f_s_dadda_rca24_and_17_19_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_17_19_y0 = f_s_dadda_rca24_and_17_19_a_17 & f_s_dadda_rca24_and_17_19_b_19;
  assign f_s_dadda_rca24_and_16_20_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_16_20_y0 = f_s_dadda_rca24_and_16_20_a_16 & f_s_dadda_rca24_and_16_20_b_20;
  assign f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_18_18_y0 = f_s_dadda_rca24_and_18_18_y0;
  assign f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_17_19_y0 = f_s_dadda_rca24_and_17_19_y0;
  assign f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_16_20_y0 = f_s_dadda_rca24_and_16_20_y0;
  assign f_s_dadda_rca24_fa307_y0 = f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_18_18_y0 ^ f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_17_19_y0;
  assign f_s_dadda_rca24_fa307_y1 = f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_18_18_y0 & f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_17_19_y0;
  assign f_s_dadda_rca24_fa307_y2 = f_s_dadda_rca24_fa307_y0 ^ f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_16_20_y0;
  assign f_s_dadda_rca24_fa307_y3 = f_s_dadda_rca24_fa307_y0 & f_s_dadda_rca24_fa307_f_s_dadda_rca24_and_16_20_y0;
  assign f_s_dadda_rca24_fa307_y4 = f_s_dadda_rca24_fa307_y1 | f_s_dadda_rca24_fa307_y3;
  assign f_s_dadda_rca24_and_15_21_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_15_21_y0 = f_s_dadda_rca24_and_15_21_a_15 & f_s_dadda_rca24_and_15_21_b_21;
  assign f_s_dadda_rca24_and_14_22_a_14 = a_14;
  assign f_s_dadda_rca24_and_14_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_14_22_y0 = f_s_dadda_rca24_and_14_22_a_14 & f_s_dadda_rca24_and_14_22_b_22;
  assign f_s_dadda_rca24_nand_13_23_a_13 = a_13;
  assign f_s_dadda_rca24_nand_13_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_13_23_y0 = ~(f_s_dadda_rca24_nand_13_23_a_13 & f_s_dadda_rca24_nand_13_23_b_23);
  assign f_s_dadda_rca24_fa308_f_s_dadda_rca24_and_15_21_y0 = f_s_dadda_rca24_and_15_21_y0;
  assign f_s_dadda_rca24_fa308_f_s_dadda_rca24_and_14_22_y0 = f_s_dadda_rca24_and_14_22_y0;
  assign f_s_dadda_rca24_fa308_f_s_dadda_rca24_nand_13_23_y0 = f_s_dadda_rca24_nand_13_23_y0;
  assign f_s_dadda_rca24_fa308_y0 = f_s_dadda_rca24_fa308_f_s_dadda_rca24_and_15_21_y0 ^ f_s_dadda_rca24_fa308_f_s_dadda_rca24_and_14_22_y0;
  assign f_s_dadda_rca24_fa308_y1 = f_s_dadda_rca24_fa308_f_s_dadda_rca24_and_15_21_y0 & f_s_dadda_rca24_fa308_f_s_dadda_rca24_and_14_22_y0;
  assign f_s_dadda_rca24_fa308_y2 = f_s_dadda_rca24_fa308_y0 ^ f_s_dadda_rca24_fa308_f_s_dadda_rca24_nand_13_23_y0;
  assign f_s_dadda_rca24_fa308_y3 = f_s_dadda_rca24_fa308_y0 & f_s_dadda_rca24_fa308_f_s_dadda_rca24_nand_13_23_y0;
  assign f_s_dadda_rca24_fa308_y4 = f_s_dadda_rca24_fa308_y1 | f_s_dadda_rca24_fa308_y3;
  assign f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa308_y4 = f_s_dadda_rca24_fa308_y4;
  assign f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa307_y4 = f_s_dadda_rca24_fa307_y4;
  assign f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa306_y4 = f_s_dadda_rca24_fa306_y4;
  assign f_s_dadda_rca24_fa309_y0 = f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa308_y4 ^ f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa307_y4;
  assign f_s_dadda_rca24_fa309_y1 = f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa308_y4 & f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa307_y4;
  assign f_s_dadda_rca24_fa309_y2 = f_s_dadda_rca24_fa309_y0 ^ f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa306_y4;
  assign f_s_dadda_rca24_fa309_y3 = f_s_dadda_rca24_fa309_y0 & f_s_dadda_rca24_fa309_f_s_dadda_rca24_fa306_y4;
  assign f_s_dadda_rca24_fa309_y4 = f_s_dadda_rca24_fa309_y1 | f_s_dadda_rca24_fa309_y3;
  assign f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa305_y4 = f_s_dadda_rca24_fa305_y4;
  assign f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa304_y4 = f_s_dadda_rca24_fa304_y4;
  assign f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa303_y4 = f_s_dadda_rca24_fa303_y4;
  assign f_s_dadda_rca24_fa310_y0 = f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa305_y4 ^ f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa304_y4;
  assign f_s_dadda_rca24_fa310_y1 = f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa305_y4 & f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa304_y4;
  assign f_s_dadda_rca24_fa310_y2 = f_s_dadda_rca24_fa310_y0 ^ f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa303_y4;
  assign f_s_dadda_rca24_fa310_y3 = f_s_dadda_rca24_fa310_y0 & f_s_dadda_rca24_fa310_f_s_dadda_rca24_fa303_y4;
  assign f_s_dadda_rca24_fa310_y4 = f_s_dadda_rca24_fa310_y1 | f_s_dadda_rca24_fa310_y3;
  assign f_s_dadda_rca24_nand_23_14_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_14_b_14 = b_14;
  assign f_s_dadda_rca24_nand_23_14_y0 = ~(f_s_dadda_rca24_nand_23_14_a_23 & f_s_dadda_rca24_nand_23_14_b_14);
  assign f_s_dadda_rca24_and_22_15_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_15_b_15 = b_15;
  assign f_s_dadda_rca24_and_22_15_y0 = f_s_dadda_rca24_and_22_15_a_22 & f_s_dadda_rca24_and_22_15_b_15;
  assign f_s_dadda_rca24_and_21_16_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_21_16_y0 = f_s_dadda_rca24_and_21_16_a_21 & f_s_dadda_rca24_and_21_16_b_16;
  assign f_s_dadda_rca24_fa311_f_s_dadda_rca24_nand_23_14_y0 = f_s_dadda_rca24_nand_23_14_y0;
  assign f_s_dadda_rca24_fa311_f_s_dadda_rca24_and_22_15_y0 = f_s_dadda_rca24_and_22_15_y0;
  assign f_s_dadda_rca24_fa311_f_s_dadda_rca24_and_21_16_y0 = f_s_dadda_rca24_and_21_16_y0;
  assign f_s_dadda_rca24_fa311_y0 = f_s_dadda_rca24_fa311_f_s_dadda_rca24_nand_23_14_y0 ^ f_s_dadda_rca24_fa311_f_s_dadda_rca24_and_22_15_y0;
  assign f_s_dadda_rca24_fa311_y1 = f_s_dadda_rca24_fa311_f_s_dadda_rca24_nand_23_14_y0 & f_s_dadda_rca24_fa311_f_s_dadda_rca24_and_22_15_y0;
  assign f_s_dadda_rca24_fa311_y2 = f_s_dadda_rca24_fa311_y0 ^ f_s_dadda_rca24_fa311_f_s_dadda_rca24_and_21_16_y0;
  assign f_s_dadda_rca24_fa311_y3 = f_s_dadda_rca24_fa311_y0 & f_s_dadda_rca24_fa311_f_s_dadda_rca24_and_21_16_y0;
  assign f_s_dadda_rca24_fa311_y4 = f_s_dadda_rca24_fa311_y1 | f_s_dadda_rca24_fa311_y3;
  assign f_s_dadda_rca24_and_20_17_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_20_17_y0 = f_s_dadda_rca24_and_20_17_a_20 & f_s_dadda_rca24_and_20_17_b_17;
  assign f_s_dadda_rca24_and_19_18_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_19_18_y0 = f_s_dadda_rca24_and_19_18_a_19 & f_s_dadda_rca24_and_19_18_b_18;
  assign f_s_dadda_rca24_and_18_19_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_18_19_y0 = f_s_dadda_rca24_and_18_19_a_18 & f_s_dadda_rca24_and_18_19_b_19;
  assign f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_20_17_y0 = f_s_dadda_rca24_and_20_17_y0;
  assign f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_19_18_y0 = f_s_dadda_rca24_and_19_18_y0;
  assign f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_18_19_y0 = f_s_dadda_rca24_and_18_19_y0;
  assign f_s_dadda_rca24_fa312_y0 = f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_20_17_y0 ^ f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_19_18_y0;
  assign f_s_dadda_rca24_fa312_y1 = f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_20_17_y0 & f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_19_18_y0;
  assign f_s_dadda_rca24_fa312_y2 = f_s_dadda_rca24_fa312_y0 ^ f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_18_19_y0;
  assign f_s_dadda_rca24_fa312_y3 = f_s_dadda_rca24_fa312_y0 & f_s_dadda_rca24_fa312_f_s_dadda_rca24_and_18_19_y0;
  assign f_s_dadda_rca24_fa312_y4 = f_s_dadda_rca24_fa312_y1 | f_s_dadda_rca24_fa312_y3;
  assign f_s_dadda_rca24_and_17_20_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_17_20_y0 = f_s_dadda_rca24_and_17_20_a_17 & f_s_dadda_rca24_and_17_20_b_20;
  assign f_s_dadda_rca24_and_16_21_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_16_21_y0 = f_s_dadda_rca24_and_16_21_a_16 & f_s_dadda_rca24_and_16_21_b_21;
  assign f_s_dadda_rca24_and_15_22_a_15 = a_15;
  assign f_s_dadda_rca24_and_15_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_15_22_y0 = f_s_dadda_rca24_and_15_22_a_15 & f_s_dadda_rca24_and_15_22_b_22;
  assign f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_17_20_y0 = f_s_dadda_rca24_and_17_20_y0;
  assign f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_16_21_y0 = f_s_dadda_rca24_and_16_21_y0;
  assign f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_15_22_y0 = f_s_dadda_rca24_and_15_22_y0;
  assign f_s_dadda_rca24_fa313_y0 = f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_17_20_y0 ^ f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_16_21_y0;
  assign f_s_dadda_rca24_fa313_y1 = f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_17_20_y0 & f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_16_21_y0;
  assign f_s_dadda_rca24_fa313_y2 = f_s_dadda_rca24_fa313_y0 ^ f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_15_22_y0;
  assign f_s_dadda_rca24_fa313_y3 = f_s_dadda_rca24_fa313_y0 & f_s_dadda_rca24_fa313_f_s_dadda_rca24_and_15_22_y0;
  assign f_s_dadda_rca24_fa313_y4 = f_s_dadda_rca24_fa313_y1 | f_s_dadda_rca24_fa313_y3;
  assign f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa313_y4 = f_s_dadda_rca24_fa313_y4;
  assign f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa312_y4 = f_s_dadda_rca24_fa312_y4;
  assign f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa311_y4 = f_s_dadda_rca24_fa311_y4;
  assign f_s_dadda_rca24_fa314_y0 = f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa313_y4 ^ f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa312_y4;
  assign f_s_dadda_rca24_fa314_y1 = f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa313_y4 & f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa312_y4;
  assign f_s_dadda_rca24_fa314_y2 = f_s_dadda_rca24_fa314_y0 ^ f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa311_y4;
  assign f_s_dadda_rca24_fa314_y3 = f_s_dadda_rca24_fa314_y0 & f_s_dadda_rca24_fa314_f_s_dadda_rca24_fa311_y4;
  assign f_s_dadda_rca24_fa314_y4 = f_s_dadda_rca24_fa314_y1 | f_s_dadda_rca24_fa314_y3;
  assign f_s_dadda_rca24_nand_23_15_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_15_b_15 = b_15;
  assign f_s_dadda_rca24_nand_23_15_y0 = ~(f_s_dadda_rca24_nand_23_15_a_23 & f_s_dadda_rca24_nand_23_15_b_15);
  assign f_s_dadda_rca24_fa315_f_s_dadda_rca24_fa310_y4 = f_s_dadda_rca24_fa310_y4;
  assign f_s_dadda_rca24_fa315_f_s_dadda_rca24_fa309_y4 = f_s_dadda_rca24_fa309_y4;
  assign f_s_dadda_rca24_fa315_f_s_dadda_rca24_nand_23_15_y0 = f_s_dadda_rca24_nand_23_15_y0;
  assign f_s_dadda_rca24_fa315_y0 = f_s_dadda_rca24_fa315_f_s_dadda_rca24_fa310_y4 ^ f_s_dadda_rca24_fa315_f_s_dadda_rca24_fa309_y4;
  assign f_s_dadda_rca24_fa315_y1 = f_s_dadda_rca24_fa315_f_s_dadda_rca24_fa310_y4 & f_s_dadda_rca24_fa315_f_s_dadda_rca24_fa309_y4;
  assign f_s_dadda_rca24_fa315_y2 = f_s_dadda_rca24_fa315_y0 ^ f_s_dadda_rca24_fa315_f_s_dadda_rca24_nand_23_15_y0;
  assign f_s_dadda_rca24_fa315_y3 = f_s_dadda_rca24_fa315_y0 & f_s_dadda_rca24_fa315_f_s_dadda_rca24_nand_23_15_y0;
  assign f_s_dadda_rca24_fa315_y4 = f_s_dadda_rca24_fa315_y1 | f_s_dadda_rca24_fa315_y3;
  assign f_s_dadda_rca24_and_22_16_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_16_b_16 = b_16;
  assign f_s_dadda_rca24_and_22_16_y0 = f_s_dadda_rca24_and_22_16_a_22 & f_s_dadda_rca24_and_22_16_b_16;
  assign f_s_dadda_rca24_and_21_17_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_21_17_y0 = f_s_dadda_rca24_and_21_17_a_21 & f_s_dadda_rca24_and_21_17_b_17;
  assign f_s_dadda_rca24_and_20_18_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_20_18_y0 = f_s_dadda_rca24_and_20_18_a_20 & f_s_dadda_rca24_and_20_18_b_18;
  assign f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_22_16_y0 = f_s_dadda_rca24_and_22_16_y0;
  assign f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_21_17_y0 = f_s_dadda_rca24_and_21_17_y0;
  assign f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_20_18_y0 = f_s_dadda_rca24_and_20_18_y0;
  assign f_s_dadda_rca24_fa316_y0 = f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_22_16_y0 ^ f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_21_17_y0;
  assign f_s_dadda_rca24_fa316_y1 = f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_22_16_y0 & f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_21_17_y0;
  assign f_s_dadda_rca24_fa316_y2 = f_s_dadda_rca24_fa316_y0 ^ f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_20_18_y0;
  assign f_s_dadda_rca24_fa316_y3 = f_s_dadda_rca24_fa316_y0 & f_s_dadda_rca24_fa316_f_s_dadda_rca24_and_20_18_y0;
  assign f_s_dadda_rca24_fa316_y4 = f_s_dadda_rca24_fa316_y1 | f_s_dadda_rca24_fa316_y3;
  assign f_s_dadda_rca24_and_19_19_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_19_19_y0 = f_s_dadda_rca24_and_19_19_a_19 & f_s_dadda_rca24_and_19_19_b_19;
  assign f_s_dadda_rca24_and_18_20_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_18_20_y0 = f_s_dadda_rca24_and_18_20_a_18 & f_s_dadda_rca24_and_18_20_b_20;
  assign f_s_dadda_rca24_and_17_21_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_17_21_y0 = f_s_dadda_rca24_and_17_21_a_17 & f_s_dadda_rca24_and_17_21_b_21;
  assign f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_19_19_y0 = f_s_dadda_rca24_and_19_19_y0;
  assign f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_18_20_y0 = f_s_dadda_rca24_and_18_20_y0;
  assign f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_17_21_y0 = f_s_dadda_rca24_and_17_21_y0;
  assign f_s_dadda_rca24_fa317_y0 = f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_19_19_y0 ^ f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_18_20_y0;
  assign f_s_dadda_rca24_fa317_y1 = f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_19_19_y0 & f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_18_20_y0;
  assign f_s_dadda_rca24_fa317_y2 = f_s_dadda_rca24_fa317_y0 ^ f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_17_21_y0;
  assign f_s_dadda_rca24_fa317_y3 = f_s_dadda_rca24_fa317_y0 & f_s_dadda_rca24_fa317_f_s_dadda_rca24_and_17_21_y0;
  assign f_s_dadda_rca24_fa317_y4 = f_s_dadda_rca24_fa317_y1 | f_s_dadda_rca24_fa317_y3;
  assign f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa317_y4 = f_s_dadda_rca24_fa317_y4;
  assign f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa316_y4 = f_s_dadda_rca24_fa316_y4;
  assign f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa315_y4 = f_s_dadda_rca24_fa315_y4;
  assign f_s_dadda_rca24_fa318_y0 = f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa317_y4 ^ f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa316_y4;
  assign f_s_dadda_rca24_fa318_y1 = f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa317_y4 & f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa316_y4;
  assign f_s_dadda_rca24_fa318_y2 = f_s_dadda_rca24_fa318_y0 ^ f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa315_y4;
  assign f_s_dadda_rca24_fa318_y3 = f_s_dadda_rca24_fa318_y0 & f_s_dadda_rca24_fa318_f_s_dadda_rca24_fa315_y4;
  assign f_s_dadda_rca24_fa318_y4 = f_s_dadda_rca24_fa318_y1 | f_s_dadda_rca24_fa318_y3;
  assign f_s_dadda_rca24_nand_23_16_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_16_b_16 = b_16;
  assign f_s_dadda_rca24_nand_23_16_y0 = ~(f_s_dadda_rca24_nand_23_16_a_23 & f_s_dadda_rca24_nand_23_16_b_16);
  assign f_s_dadda_rca24_and_22_17_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_17_b_17 = b_17;
  assign f_s_dadda_rca24_and_22_17_y0 = f_s_dadda_rca24_and_22_17_a_22 & f_s_dadda_rca24_and_22_17_b_17;
  assign f_s_dadda_rca24_fa319_f_s_dadda_rca24_fa314_y4 = f_s_dadda_rca24_fa314_y4;
  assign f_s_dadda_rca24_fa319_f_s_dadda_rca24_nand_23_16_y0 = f_s_dadda_rca24_nand_23_16_y0;
  assign f_s_dadda_rca24_fa319_f_s_dadda_rca24_and_22_17_y0 = f_s_dadda_rca24_and_22_17_y0;
  assign f_s_dadda_rca24_fa319_y0 = f_s_dadda_rca24_fa319_f_s_dadda_rca24_fa314_y4 ^ f_s_dadda_rca24_fa319_f_s_dadda_rca24_nand_23_16_y0;
  assign f_s_dadda_rca24_fa319_y1 = f_s_dadda_rca24_fa319_f_s_dadda_rca24_fa314_y4 & f_s_dadda_rca24_fa319_f_s_dadda_rca24_nand_23_16_y0;
  assign f_s_dadda_rca24_fa319_y2 = f_s_dadda_rca24_fa319_y0 ^ f_s_dadda_rca24_fa319_f_s_dadda_rca24_and_22_17_y0;
  assign f_s_dadda_rca24_fa319_y3 = f_s_dadda_rca24_fa319_y0 & f_s_dadda_rca24_fa319_f_s_dadda_rca24_and_22_17_y0;
  assign f_s_dadda_rca24_fa319_y4 = f_s_dadda_rca24_fa319_y1 | f_s_dadda_rca24_fa319_y3;
  assign f_s_dadda_rca24_and_21_18_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_21_18_y0 = f_s_dadda_rca24_and_21_18_a_21 & f_s_dadda_rca24_and_21_18_b_18;
  assign f_s_dadda_rca24_and_20_19_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_20_19_y0 = f_s_dadda_rca24_and_20_19_a_20 & f_s_dadda_rca24_and_20_19_b_19;
  assign f_s_dadda_rca24_and_19_20_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_19_20_y0 = f_s_dadda_rca24_and_19_20_a_19 & f_s_dadda_rca24_and_19_20_b_20;
  assign f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_21_18_y0 = f_s_dadda_rca24_and_21_18_y0;
  assign f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_20_19_y0 = f_s_dadda_rca24_and_20_19_y0;
  assign f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_19_20_y0 = f_s_dadda_rca24_and_19_20_y0;
  assign f_s_dadda_rca24_fa320_y0 = f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_21_18_y0 ^ f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_20_19_y0;
  assign f_s_dadda_rca24_fa320_y1 = f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_21_18_y0 & f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_20_19_y0;
  assign f_s_dadda_rca24_fa320_y2 = f_s_dadda_rca24_fa320_y0 ^ f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_19_20_y0;
  assign f_s_dadda_rca24_fa320_y3 = f_s_dadda_rca24_fa320_y0 & f_s_dadda_rca24_fa320_f_s_dadda_rca24_and_19_20_y0;
  assign f_s_dadda_rca24_fa320_y4 = f_s_dadda_rca24_fa320_y1 | f_s_dadda_rca24_fa320_y3;
  assign f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa320_y4 = f_s_dadda_rca24_fa320_y4;
  assign f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa319_y4 = f_s_dadda_rca24_fa319_y4;
  assign f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa318_y4 = f_s_dadda_rca24_fa318_y4;
  assign f_s_dadda_rca24_fa321_y0 = f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa320_y4 ^ f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa319_y4;
  assign f_s_dadda_rca24_fa321_y1 = f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa320_y4 & f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa319_y4;
  assign f_s_dadda_rca24_fa321_y2 = f_s_dadda_rca24_fa321_y0 ^ f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa318_y4;
  assign f_s_dadda_rca24_fa321_y3 = f_s_dadda_rca24_fa321_y0 & f_s_dadda_rca24_fa321_f_s_dadda_rca24_fa318_y4;
  assign f_s_dadda_rca24_fa321_y4 = f_s_dadda_rca24_fa321_y1 | f_s_dadda_rca24_fa321_y3;
  assign f_s_dadda_rca24_nand_23_17_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_17_b_17 = b_17;
  assign f_s_dadda_rca24_nand_23_17_y0 = ~(f_s_dadda_rca24_nand_23_17_a_23 & f_s_dadda_rca24_nand_23_17_b_17);
  assign f_s_dadda_rca24_and_22_18_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_18_b_18 = b_18;
  assign f_s_dadda_rca24_and_22_18_y0 = f_s_dadda_rca24_and_22_18_a_22 & f_s_dadda_rca24_and_22_18_b_18;
  assign f_s_dadda_rca24_and_21_19_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_21_19_y0 = f_s_dadda_rca24_and_21_19_a_21 & f_s_dadda_rca24_and_21_19_b_19;
  assign f_s_dadda_rca24_fa322_f_s_dadda_rca24_nand_23_17_y0 = f_s_dadda_rca24_nand_23_17_y0;
  assign f_s_dadda_rca24_fa322_f_s_dadda_rca24_and_22_18_y0 = f_s_dadda_rca24_and_22_18_y0;
  assign f_s_dadda_rca24_fa322_f_s_dadda_rca24_and_21_19_y0 = f_s_dadda_rca24_and_21_19_y0;
  assign f_s_dadda_rca24_fa322_y0 = f_s_dadda_rca24_fa322_f_s_dadda_rca24_nand_23_17_y0 ^ f_s_dadda_rca24_fa322_f_s_dadda_rca24_and_22_18_y0;
  assign f_s_dadda_rca24_fa322_y1 = f_s_dadda_rca24_fa322_f_s_dadda_rca24_nand_23_17_y0 & f_s_dadda_rca24_fa322_f_s_dadda_rca24_and_22_18_y0;
  assign f_s_dadda_rca24_fa322_y2 = f_s_dadda_rca24_fa322_y0 ^ f_s_dadda_rca24_fa322_f_s_dadda_rca24_and_21_19_y0;
  assign f_s_dadda_rca24_fa322_y3 = f_s_dadda_rca24_fa322_y0 & f_s_dadda_rca24_fa322_f_s_dadda_rca24_and_21_19_y0;
  assign f_s_dadda_rca24_fa322_y4 = f_s_dadda_rca24_fa322_y1 | f_s_dadda_rca24_fa322_y3;
  assign f_s_dadda_rca24_nand_23_18_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_18_b_18 = b_18;
  assign f_s_dadda_rca24_nand_23_18_y0 = ~(f_s_dadda_rca24_nand_23_18_a_23 & f_s_dadda_rca24_nand_23_18_b_18);
  assign f_s_dadda_rca24_fa323_f_s_dadda_rca24_fa322_y4 = f_s_dadda_rca24_fa322_y4;
  assign f_s_dadda_rca24_fa323_f_s_dadda_rca24_fa321_y4 = f_s_dadda_rca24_fa321_y4;
  assign f_s_dadda_rca24_fa323_f_s_dadda_rca24_nand_23_18_y0 = f_s_dadda_rca24_nand_23_18_y0;
  assign f_s_dadda_rca24_fa323_y0 = f_s_dadda_rca24_fa323_f_s_dadda_rca24_fa322_y4 ^ f_s_dadda_rca24_fa323_f_s_dadda_rca24_fa321_y4;
  assign f_s_dadda_rca24_fa323_y1 = f_s_dadda_rca24_fa323_f_s_dadda_rca24_fa322_y4 & f_s_dadda_rca24_fa323_f_s_dadda_rca24_fa321_y4;
  assign f_s_dadda_rca24_fa323_y2 = f_s_dadda_rca24_fa323_y0 ^ f_s_dadda_rca24_fa323_f_s_dadda_rca24_nand_23_18_y0;
  assign f_s_dadda_rca24_fa323_y3 = f_s_dadda_rca24_fa323_y0 & f_s_dadda_rca24_fa323_f_s_dadda_rca24_nand_23_18_y0;
  assign f_s_dadda_rca24_fa323_y4 = f_s_dadda_rca24_fa323_y1 | f_s_dadda_rca24_fa323_y3;
  assign f_s_dadda_rca24_and_4_0_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_4_0_y0 = f_s_dadda_rca24_and_4_0_a_4 & f_s_dadda_rca24_and_4_0_b_0;
  assign f_s_dadda_rca24_and_3_1_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_3_1_y0 = f_s_dadda_rca24_and_3_1_a_3 & f_s_dadda_rca24_and_3_1_b_1;
  assign f_s_dadda_rca24_ha18_f_s_dadda_rca24_and_4_0_y0 = f_s_dadda_rca24_and_4_0_y0;
  assign f_s_dadda_rca24_ha18_f_s_dadda_rca24_and_3_1_y0 = f_s_dadda_rca24_and_3_1_y0;
  assign f_s_dadda_rca24_ha18_y0 = f_s_dadda_rca24_ha18_f_s_dadda_rca24_and_4_0_y0 ^ f_s_dadda_rca24_ha18_f_s_dadda_rca24_and_3_1_y0;
  assign f_s_dadda_rca24_ha18_y1 = f_s_dadda_rca24_ha18_f_s_dadda_rca24_and_4_0_y0 & f_s_dadda_rca24_ha18_f_s_dadda_rca24_and_3_1_y0;
  assign f_s_dadda_rca24_and_5_0_a_5 = a_5;
  assign f_s_dadda_rca24_and_5_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_5_0_y0 = f_s_dadda_rca24_and_5_0_a_5 & f_s_dadda_rca24_and_5_0_b_0;
  assign f_s_dadda_rca24_and_4_1_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_4_1_y0 = f_s_dadda_rca24_and_4_1_a_4 & f_s_dadda_rca24_and_4_1_b_1;
  assign f_s_dadda_rca24_fa324_f_s_dadda_rca24_ha18_y1 = f_s_dadda_rca24_ha18_y1;
  assign f_s_dadda_rca24_fa324_f_s_dadda_rca24_and_5_0_y0 = f_s_dadda_rca24_and_5_0_y0;
  assign f_s_dadda_rca24_fa324_f_s_dadda_rca24_and_4_1_y0 = f_s_dadda_rca24_and_4_1_y0;
  assign f_s_dadda_rca24_fa324_y0 = f_s_dadda_rca24_fa324_f_s_dadda_rca24_ha18_y1 ^ f_s_dadda_rca24_fa324_f_s_dadda_rca24_and_5_0_y0;
  assign f_s_dadda_rca24_fa324_y1 = f_s_dadda_rca24_fa324_f_s_dadda_rca24_ha18_y1 & f_s_dadda_rca24_fa324_f_s_dadda_rca24_and_5_0_y0;
  assign f_s_dadda_rca24_fa324_y2 = f_s_dadda_rca24_fa324_y0 ^ f_s_dadda_rca24_fa324_f_s_dadda_rca24_and_4_1_y0;
  assign f_s_dadda_rca24_fa324_y3 = f_s_dadda_rca24_fa324_y0 & f_s_dadda_rca24_fa324_f_s_dadda_rca24_and_4_1_y0;
  assign f_s_dadda_rca24_fa324_y4 = f_s_dadda_rca24_fa324_y1 | f_s_dadda_rca24_fa324_y3;
  assign f_s_dadda_rca24_and_3_2_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_3_2_y0 = f_s_dadda_rca24_and_3_2_a_3 & f_s_dadda_rca24_and_3_2_b_2;
  assign f_s_dadda_rca24_and_2_3_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_2_3_y0 = f_s_dadda_rca24_and_2_3_a_2 & f_s_dadda_rca24_and_2_3_b_3;
  assign f_s_dadda_rca24_ha19_f_s_dadda_rca24_and_3_2_y0 = f_s_dadda_rca24_and_3_2_y0;
  assign f_s_dadda_rca24_ha19_f_s_dadda_rca24_and_2_3_y0 = f_s_dadda_rca24_and_2_3_y0;
  assign f_s_dadda_rca24_ha19_y0 = f_s_dadda_rca24_ha19_f_s_dadda_rca24_and_3_2_y0 ^ f_s_dadda_rca24_ha19_f_s_dadda_rca24_and_2_3_y0;
  assign f_s_dadda_rca24_ha19_y1 = f_s_dadda_rca24_ha19_f_s_dadda_rca24_and_3_2_y0 & f_s_dadda_rca24_ha19_f_s_dadda_rca24_and_2_3_y0;
  assign f_s_dadda_rca24_and_4_2_a_4 = a_4;
  assign f_s_dadda_rca24_and_4_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_4_2_y0 = f_s_dadda_rca24_and_4_2_a_4 & f_s_dadda_rca24_and_4_2_b_2;
  assign f_s_dadda_rca24_fa325_f_s_dadda_rca24_ha19_y1 = f_s_dadda_rca24_ha19_y1;
  assign f_s_dadda_rca24_fa325_f_s_dadda_rca24_fa324_y4 = f_s_dadda_rca24_fa324_y4;
  assign f_s_dadda_rca24_fa325_f_s_dadda_rca24_and_4_2_y0 = f_s_dadda_rca24_and_4_2_y0;
  assign f_s_dadda_rca24_fa325_y0 = f_s_dadda_rca24_fa325_f_s_dadda_rca24_ha19_y1 ^ f_s_dadda_rca24_fa325_f_s_dadda_rca24_fa324_y4;
  assign f_s_dadda_rca24_fa325_y1 = f_s_dadda_rca24_fa325_f_s_dadda_rca24_ha19_y1 & f_s_dadda_rca24_fa325_f_s_dadda_rca24_fa324_y4;
  assign f_s_dadda_rca24_fa325_y2 = f_s_dadda_rca24_fa325_y0 ^ f_s_dadda_rca24_fa325_f_s_dadda_rca24_and_4_2_y0;
  assign f_s_dadda_rca24_fa325_y3 = f_s_dadda_rca24_fa325_y0 & f_s_dadda_rca24_fa325_f_s_dadda_rca24_and_4_2_y0;
  assign f_s_dadda_rca24_fa325_y4 = f_s_dadda_rca24_fa325_y1 | f_s_dadda_rca24_fa325_y3;
  assign f_s_dadda_rca24_and_3_3_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_3_3_y0 = f_s_dadda_rca24_and_3_3_a_3 & f_s_dadda_rca24_and_3_3_b_3;
  assign f_s_dadda_rca24_and_2_4_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_2_4_y0 = f_s_dadda_rca24_and_2_4_a_2 & f_s_dadda_rca24_and_2_4_b_4;
  assign f_s_dadda_rca24_and_1_5_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_1_5_y0 = f_s_dadda_rca24_and_1_5_a_1 & f_s_dadda_rca24_and_1_5_b_5;
  assign f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_3_3_y0 = f_s_dadda_rca24_and_3_3_y0;
  assign f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_2_4_y0 = f_s_dadda_rca24_and_2_4_y0;
  assign f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_1_5_y0 = f_s_dadda_rca24_and_1_5_y0;
  assign f_s_dadda_rca24_fa326_y0 = f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_3_3_y0 ^ f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_2_4_y0;
  assign f_s_dadda_rca24_fa326_y1 = f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_3_3_y0 & f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_2_4_y0;
  assign f_s_dadda_rca24_fa326_y2 = f_s_dadda_rca24_fa326_y0 ^ f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_1_5_y0;
  assign f_s_dadda_rca24_fa326_y3 = f_s_dadda_rca24_fa326_y0 & f_s_dadda_rca24_fa326_f_s_dadda_rca24_and_1_5_y0;
  assign f_s_dadda_rca24_fa326_y4 = f_s_dadda_rca24_fa326_y1 | f_s_dadda_rca24_fa326_y3;
  assign f_s_dadda_rca24_and_3_4_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_3_4_y0 = f_s_dadda_rca24_and_3_4_a_3 & f_s_dadda_rca24_and_3_4_b_4;
  assign f_s_dadda_rca24_fa327_f_s_dadda_rca24_fa326_y4 = f_s_dadda_rca24_fa326_y4;
  assign f_s_dadda_rca24_fa327_f_s_dadda_rca24_fa325_y4 = f_s_dadda_rca24_fa325_y4;
  assign f_s_dadda_rca24_fa327_f_s_dadda_rca24_and_3_4_y0 = f_s_dadda_rca24_and_3_4_y0;
  assign f_s_dadda_rca24_fa327_y0 = f_s_dadda_rca24_fa327_f_s_dadda_rca24_fa326_y4 ^ f_s_dadda_rca24_fa327_f_s_dadda_rca24_fa325_y4;
  assign f_s_dadda_rca24_fa327_y1 = f_s_dadda_rca24_fa327_f_s_dadda_rca24_fa326_y4 & f_s_dadda_rca24_fa327_f_s_dadda_rca24_fa325_y4;
  assign f_s_dadda_rca24_fa327_y2 = f_s_dadda_rca24_fa327_y0 ^ f_s_dadda_rca24_fa327_f_s_dadda_rca24_and_3_4_y0;
  assign f_s_dadda_rca24_fa327_y3 = f_s_dadda_rca24_fa327_y0 & f_s_dadda_rca24_fa327_f_s_dadda_rca24_and_3_4_y0;
  assign f_s_dadda_rca24_fa327_y4 = f_s_dadda_rca24_fa327_y1 | f_s_dadda_rca24_fa327_y3;
  assign f_s_dadda_rca24_and_2_5_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_2_5_y0 = f_s_dadda_rca24_and_2_5_a_2 & f_s_dadda_rca24_and_2_5_b_5;
  assign f_s_dadda_rca24_and_1_6_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_1_6_y0 = f_s_dadda_rca24_and_1_6_a_1 & f_s_dadda_rca24_and_1_6_b_6;
  assign f_s_dadda_rca24_and_0_7_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_0_7_y0 = f_s_dadda_rca24_and_0_7_a_0 & f_s_dadda_rca24_and_0_7_b_7;
  assign f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_2_5_y0 = f_s_dadda_rca24_and_2_5_y0;
  assign f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_1_6_y0 = f_s_dadda_rca24_and_1_6_y0;
  assign f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_0_7_y0 = f_s_dadda_rca24_and_0_7_y0;
  assign f_s_dadda_rca24_fa328_y0 = f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_2_5_y0 ^ f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_1_6_y0;
  assign f_s_dadda_rca24_fa328_y1 = f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_2_5_y0 & f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_1_6_y0;
  assign f_s_dadda_rca24_fa328_y2 = f_s_dadda_rca24_fa328_y0 ^ f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_0_7_y0;
  assign f_s_dadda_rca24_fa328_y3 = f_s_dadda_rca24_fa328_y0 & f_s_dadda_rca24_fa328_f_s_dadda_rca24_and_0_7_y0;
  assign f_s_dadda_rca24_fa328_y4 = f_s_dadda_rca24_fa328_y1 | f_s_dadda_rca24_fa328_y3;
  assign f_s_dadda_rca24_and_2_6_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_2_6_y0 = f_s_dadda_rca24_and_2_6_a_2 & f_s_dadda_rca24_and_2_6_b_6;
  assign f_s_dadda_rca24_fa329_f_s_dadda_rca24_fa328_y4 = f_s_dadda_rca24_fa328_y4;
  assign f_s_dadda_rca24_fa329_f_s_dadda_rca24_fa327_y4 = f_s_dadda_rca24_fa327_y4;
  assign f_s_dadda_rca24_fa329_f_s_dadda_rca24_and_2_6_y0 = f_s_dadda_rca24_and_2_6_y0;
  assign f_s_dadda_rca24_fa329_y0 = f_s_dadda_rca24_fa329_f_s_dadda_rca24_fa328_y4 ^ f_s_dadda_rca24_fa329_f_s_dadda_rca24_fa327_y4;
  assign f_s_dadda_rca24_fa329_y1 = f_s_dadda_rca24_fa329_f_s_dadda_rca24_fa328_y4 & f_s_dadda_rca24_fa329_f_s_dadda_rca24_fa327_y4;
  assign f_s_dadda_rca24_fa329_y2 = f_s_dadda_rca24_fa329_y0 ^ f_s_dadda_rca24_fa329_f_s_dadda_rca24_and_2_6_y0;
  assign f_s_dadda_rca24_fa329_y3 = f_s_dadda_rca24_fa329_y0 & f_s_dadda_rca24_fa329_f_s_dadda_rca24_and_2_6_y0;
  assign f_s_dadda_rca24_fa329_y4 = f_s_dadda_rca24_fa329_y1 | f_s_dadda_rca24_fa329_y3;
  assign f_s_dadda_rca24_and_1_7_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_7_b_7 = b_7;
  assign f_s_dadda_rca24_and_1_7_y0 = f_s_dadda_rca24_and_1_7_a_1 & f_s_dadda_rca24_and_1_7_b_7;
  assign f_s_dadda_rca24_and_0_8_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_0_8_y0 = f_s_dadda_rca24_and_0_8_a_0 & f_s_dadda_rca24_and_0_8_b_8;
  assign f_s_dadda_rca24_fa330_f_s_dadda_rca24_and_1_7_y0 = f_s_dadda_rca24_and_1_7_y0;
  assign f_s_dadda_rca24_fa330_f_s_dadda_rca24_and_0_8_y0 = f_s_dadda_rca24_and_0_8_y0;
  assign f_s_dadda_rca24_fa330_f_s_dadda_rca24_fa26_y2 = f_s_dadda_rca24_fa26_y2;
  assign f_s_dadda_rca24_fa330_y0 = f_s_dadda_rca24_fa330_f_s_dadda_rca24_and_1_7_y0 ^ f_s_dadda_rca24_fa330_f_s_dadda_rca24_and_0_8_y0;
  assign f_s_dadda_rca24_fa330_y1 = f_s_dadda_rca24_fa330_f_s_dadda_rca24_and_1_7_y0 & f_s_dadda_rca24_fa330_f_s_dadda_rca24_and_0_8_y0;
  assign f_s_dadda_rca24_fa330_y2 = f_s_dadda_rca24_fa330_y0 ^ f_s_dadda_rca24_fa330_f_s_dadda_rca24_fa26_y2;
  assign f_s_dadda_rca24_fa330_y3 = f_s_dadda_rca24_fa330_y0 & f_s_dadda_rca24_fa330_f_s_dadda_rca24_fa26_y2;
  assign f_s_dadda_rca24_fa330_y4 = f_s_dadda_rca24_fa330_y1 | f_s_dadda_rca24_fa330_y3;
  assign f_s_dadda_rca24_and_1_8_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_8_b_8 = b_8;
  assign f_s_dadda_rca24_and_1_8_y0 = f_s_dadda_rca24_and_1_8_a_1 & f_s_dadda_rca24_and_1_8_b_8;
  assign f_s_dadda_rca24_fa331_f_s_dadda_rca24_fa330_y4 = f_s_dadda_rca24_fa330_y4;
  assign f_s_dadda_rca24_fa331_f_s_dadda_rca24_fa329_y4 = f_s_dadda_rca24_fa329_y4;
  assign f_s_dadda_rca24_fa331_f_s_dadda_rca24_and_1_8_y0 = f_s_dadda_rca24_and_1_8_y0;
  assign f_s_dadda_rca24_fa331_y0 = f_s_dadda_rca24_fa331_f_s_dadda_rca24_fa330_y4 ^ f_s_dadda_rca24_fa331_f_s_dadda_rca24_fa329_y4;
  assign f_s_dadda_rca24_fa331_y1 = f_s_dadda_rca24_fa331_f_s_dadda_rca24_fa330_y4 & f_s_dadda_rca24_fa331_f_s_dadda_rca24_fa329_y4;
  assign f_s_dadda_rca24_fa331_y2 = f_s_dadda_rca24_fa331_y0 ^ f_s_dadda_rca24_fa331_f_s_dadda_rca24_and_1_8_y0;
  assign f_s_dadda_rca24_fa331_y3 = f_s_dadda_rca24_fa331_y0 & f_s_dadda_rca24_fa331_f_s_dadda_rca24_and_1_8_y0;
  assign f_s_dadda_rca24_fa331_y4 = f_s_dadda_rca24_fa331_y1 | f_s_dadda_rca24_fa331_y3;
  assign f_s_dadda_rca24_and_0_9_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_9_b_9 = b_9;
  assign f_s_dadda_rca24_and_0_9_y0 = f_s_dadda_rca24_and_0_9_a_0 & f_s_dadda_rca24_and_0_9_b_9;
  assign f_s_dadda_rca24_fa332_f_s_dadda_rca24_and_0_9_y0 = f_s_dadda_rca24_and_0_9_y0;
  assign f_s_dadda_rca24_fa332_f_s_dadda_rca24_fa28_y2 = f_s_dadda_rca24_fa28_y2;
  assign f_s_dadda_rca24_fa332_f_s_dadda_rca24_fa29_y2 = f_s_dadda_rca24_fa29_y2;
  assign f_s_dadda_rca24_fa332_y0 = f_s_dadda_rca24_fa332_f_s_dadda_rca24_and_0_9_y0 ^ f_s_dadda_rca24_fa332_f_s_dadda_rca24_fa28_y2;
  assign f_s_dadda_rca24_fa332_y1 = f_s_dadda_rca24_fa332_f_s_dadda_rca24_and_0_9_y0 & f_s_dadda_rca24_fa332_f_s_dadda_rca24_fa28_y2;
  assign f_s_dadda_rca24_fa332_y2 = f_s_dadda_rca24_fa332_y0 ^ f_s_dadda_rca24_fa332_f_s_dadda_rca24_fa29_y2;
  assign f_s_dadda_rca24_fa332_y3 = f_s_dadda_rca24_fa332_y0 & f_s_dadda_rca24_fa332_f_s_dadda_rca24_fa29_y2;
  assign f_s_dadda_rca24_fa332_y4 = f_s_dadda_rca24_fa332_y1 | f_s_dadda_rca24_fa332_y3;
  assign f_s_dadda_rca24_and_0_10_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_10_b_10 = b_10;
  assign f_s_dadda_rca24_and_0_10_y0 = f_s_dadda_rca24_and_0_10_a_0 & f_s_dadda_rca24_and_0_10_b_10;
  assign f_s_dadda_rca24_fa333_f_s_dadda_rca24_fa332_y4 = f_s_dadda_rca24_fa332_y4;
  assign f_s_dadda_rca24_fa333_f_s_dadda_rca24_fa331_y4 = f_s_dadda_rca24_fa331_y4;
  assign f_s_dadda_rca24_fa333_f_s_dadda_rca24_and_0_10_y0 = f_s_dadda_rca24_and_0_10_y0;
  assign f_s_dadda_rca24_fa333_y0 = f_s_dadda_rca24_fa333_f_s_dadda_rca24_fa332_y4 ^ f_s_dadda_rca24_fa333_f_s_dadda_rca24_fa331_y4;
  assign f_s_dadda_rca24_fa333_y1 = f_s_dadda_rca24_fa333_f_s_dadda_rca24_fa332_y4 & f_s_dadda_rca24_fa333_f_s_dadda_rca24_fa331_y4;
  assign f_s_dadda_rca24_fa333_y2 = f_s_dadda_rca24_fa333_y0 ^ f_s_dadda_rca24_fa333_f_s_dadda_rca24_and_0_10_y0;
  assign f_s_dadda_rca24_fa333_y3 = f_s_dadda_rca24_fa333_y0 & f_s_dadda_rca24_fa333_f_s_dadda_rca24_and_0_10_y0;
  assign f_s_dadda_rca24_fa333_y4 = f_s_dadda_rca24_fa333_y1 | f_s_dadda_rca24_fa333_y3;
  assign f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa31_y2 = f_s_dadda_rca24_fa31_y2;
  assign f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa32_y2 = f_s_dadda_rca24_fa32_y2;
  assign f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa33_y2 = f_s_dadda_rca24_fa33_y2;
  assign f_s_dadda_rca24_fa334_y0 = f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa31_y2 ^ f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa32_y2;
  assign f_s_dadda_rca24_fa334_y1 = f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa31_y2 & f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa32_y2;
  assign f_s_dadda_rca24_fa334_y2 = f_s_dadda_rca24_fa334_y0 ^ f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa33_y2;
  assign f_s_dadda_rca24_fa334_y3 = f_s_dadda_rca24_fa334_y0 & f_s_dadda_rca24_fa334_f_s_dadda_rca24_fa33_y2;
  assign f_s_dadda_rca24_fa334_y4 = f_s_dadda_rca24_fa334_y1 | f_s_dadda_rca24_fa334_y3;
  assign f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa334_y4 = f_s_dadda_rca24_fa334_y4;
  assign f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa333_y4 = f_s_dadda_rca24_fa333_y4;
  assign f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa35_y2 = f_s_dadda_rca24_fa35_y2;
  assign f_s_dadda_rca24_fa335_y0 = f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa334_y4 ^ f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa333_y4;
  assign f_s_dadda_rca24_fa335_y1 = f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa334_y4 & f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa333_y4;
  assign f_s_dadda_rca24_fa335_y2 = f_s_dadda_rca24_fa335_y0 ^ f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa35_y2;
  assign f_s_dadda_rca24_fa335_y3 = f_s_dadda_rca24_fa335_y0 & f_s_dadda_rca24_fa335_f_s_dadda_rca24_fa35_y2;
  assign f_s_dadda_rca24_fa335_y4 = f_s_dadda_rca24_fa335_y1 | f_s_dadda_rca24_fa335_y3;
  assign f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa36_y2 = f_s_dadda_rca24_fa36_y2;
  assign f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa37_y2 = f_s_dadda_rca24_fa37_y2;
  assign f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa38_y2 = f_s_dadda_rca24_fa38_y2;
  assign f_s_dadda_rca24_fa336_y0 = f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa36_y2 ^ f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa37_y2;
  assign f_s_dadda_rca24_fa336_y1 = f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa36_y2 & f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa37_y2;
  assign f_s_dadda_rca24_fa336_y2 = f_s_dadda_rca24_fa336_y0 ^ f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa38_y2;
  assign f_s_dadda_rca24_fa336_y3 = f_s_dadda_rca24_fa336_y0 & f_s_dadda_rca24_fa336_f_s_dadda_rca24_fa38_y2;
  assign f_s_dadda_rca24_fa336_y4 = f_s_dadda_rca24_fa336_y1 | f_s_dadda_rca24_fa336_y3;
  assign f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa336_y4 = f_s_dadda_rca24_fa336_y4;
  assign f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa335_y4 = f_s_dadda_rca24_fa335_y4;
  assign f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa41_y2 = f_s_dadda_rca24_fa41_y2;
  assign f_s_dadda_rca24_fa337_y0 = f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa336_y4 ^ f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa335_y4;
  assign f_s_dadda_rca24_fa337_y1 = f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa336_y4 & f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa335_y4;
  assign f_s_dadda_rca24_fa337_y2 = f_s_dadda_rca24_fa337_y0 ^ f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa41_y2;
  assign f_s_dadda_rca24_fa337_y3 = f_s_dadda_rca24_fa337_y0 & f_s_dadda_rca24_fa337_f_s_dadda_rca24_fa41_y2;
  assign f_s_dadda_rca24_fa337_y4 = f_s_dadda_rca24_fa337_y1 | f_s_dadda_rca24_fa337_y3;
  assign f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa42_y2 = f_s_dadda_rca24_fa42_y2;
  assign f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa43_y2 = f_s_dadda_rca24_fa43_y2;
  assign f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa44_y2 = f_s_dadda_rca24_fa44_y2;
  assign f_s_dadda_rca24_fa338_y0 = f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa42_y2 ^ f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa43_y2;
  assign f_s_dadda_rca24_fa338_y1 = f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa42_y2 & f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa43_y2;
  assign f_s_dadda_rca24_fa338_y2 = f_s_dadda_rca24_fa338_y0 ^ f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa44_y2;
  assign f_s_dadda_rca24_fa338_y3 = f_s_dadda_rca24_fa338_y0 & f_s_dadda_rca24_fa338_f_s_dadda_rca24_fa44_y2;
  assign f_s_dadda_rca24_fa338_y4 = f_s_dadda_rca24_fa338_y1 | f_s_dadda_rca24_fa338_y3;
  assign f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa338_y4 = f_s_dadda_rca24_fa338_y4;
  assign f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa337_y4 = f_s_dadda_rca24_fa337_y4;
  assign f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa48_y2 = f_s_dadda_rca24_fa48_y2;
  assign f_s_dadda_rca24_fa339_y0 = f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa338_y4 ^ f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa337_y4;
  assign f_s_dadda_rca24_fa339_y1 = f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa338_y4 & f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa337_y4;
  assign f_s_dadda_rca24_fa339_y2 = f_s_dadda_rca24_fa339_y0 ^ f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa48_y2;
  assign f_s_dadda_rca24_fa339_y3 = f_s_dadda_rca24_fa339_y0 & f_s_dadda_rca24_fa339_f_s_dadda_rca24_fa48_y2;
  assign f_s_dadda_rca24_fa339_y4 = f_s_dadda_rca24_fa339_y1 | f_s_dadda_rca24_fa339_y3;
  assign f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa49_y2 = f_s_dadda_rca24_fa49_y2;
  assign f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa50_y2 = f_s_dadda_rca24_fa50_y2;
  assign f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa51_y2 = f_s_dadda_rca24_fa51_y2;
  assign f_s_dadda_rca24_fa340_y0 = f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa49_y2 ^ f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa50_y2;
  assign f_s_dadda_rca24_fa340_y1 = f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa49_y2 & f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa50_y2;
  assign f_s_dadda_rca24_fa340_y2 = f_s_dadda_rca24_fa340_y0 ^ f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa51_y2;
  assign f_s_dadda_rca24_fa340_y3 = f_s_dadda_rca24_fa340_y0 & f_s_dadda_rca24_fa340_f_s_dadda_rca24_fa51_y2;
  assign f_s_dadda_rca24_fa340_y4 = f_s_dadda_rca24_fa340_y1 | f_s_dadda_rca24_fa340_y3;
  assign f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa340_y4 = f_s_dadda_rca24_fa340_y4;
  assign f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa339_y4 = f_s_dadda_rca24_fa339_y4;
  assign f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa56_y2 = f_s_dadda_rca24_fa56_y2;
  assign f_s_dadda_rca24_fa341_y0 = f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa340_y4 ^ f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa339_y4;
  assign f_s_dadda_rca24_fa341_y1 = f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa340_y4 & f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa339_y4;
  assign f_s_dadda_rca24_fa341_y2 = f_s_dadda_rca24_fa341_y0 ^ f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa56_y2;
  assign f_s_dadda_rca24_fa341_y3 = f_s_dadda_rca24_fa341_y0 & f_s_dadda_rca24_fa341_f_s_dadda_rca24_fa56_y2;
  assign f_s_dadda_rca24_fa341_y4 = f_s_dadda_rca24_fa341_y1 | f_s_dadda_rca24_fa341_y3;
  assign f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa57_y2 = f_s_dadda_rca24_fa57_y2;
  assign f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa58_y2 = f_s_dadda_rca24_fa58_y2;
  assign f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa59_y2 = f_s_dadda_rca24_fa59_y2;
  assign f_s_dadda_rca24_fa342_y0 = f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa57_y2 ^ f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa58_y2;
  assign f_s_dadda_rca24_fa342_y1 = f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa57_y2 & f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa58_y2;
  assign f_s_dadda_rca24_fa342_y2 = f_s_dadda_rca24_fa342_y0 ^ f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa59_y2;
  assign f_s_dadda_rca24_fa342_y3 = f_s_dadda_rca24_fa342_y0 & f_s_dadda_rca24_fa342_f_s_dadda_rca24_fa59_y2;
  assign f_s_dadda_rca24_fa342_y4 = f_s_dadda_rca24_fa342_y1 | f_s_dadda_rca24_fa342_y3;
  assign f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa342_y4 = f_s_dadda_rca24_fa342_y4;
  assign f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa341_y4 = f_s_dadda_rca24_fa341_y4;
  assign f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa65_y2 = f_s_dadda_rca24_fa65_y2;
  assign f_s_dadda_rca24_fa343_y0 = f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa342_y4 ^ f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa341_y4;
  assign f_s_dadda_rca24_fa343_y1 = f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa342_y4 & f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa341_y4;
  assign f_s_dadda_rca24_fa343_y2 = f_s_dadda_rca24_fa343_y0 ^ f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa65_y2;
  assign f_s_dadda_rca24_fa343_y3 = f_s_dadda_rca24_fa343_y0 & f_s_dadda_rca24_fa343_f_s_dadda_rca24_fa65_y2;
  assign f_s_dadda_rca24_fa343_y4 = f_s_dadda_rca24_fa343_y1 | f_s_dadda_rca24_fa343_y3;
  assign f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa66_y2 = f_s_dadda_rca24_fa66_y2;
  assign f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa67_y2 = f_s_dadda_rca24_fa67_y2;
  assign f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa68_y2 = f_s_dadda_rca24_fa68_y2;
  assign f_s_dadda_rca24_fa344_y0 = f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa66_y2 ^ f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa67_y2;
  assign f_s_dadda_rca24_fa344_y1 = f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa66_y2 & f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa67_y2;
  assign f_s_dadda_rca24_fa344_y2 = f_s_dadda_rca24_fa344_y0 ^ f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa68_y2;
  assign f_s_dadda_rca24_fa344_y3 = f_s_dadda_rca24_fa344_y0 & f_s_dadda_rca24_fa344_f_s_dadda_rca24_fa68_y2;
  assign f_s_dadda_rca24_fa344_y4 = f_s_dadda_rca24_fa344_y1 | f_s_dadda_rca24_fa344_y3;
  assign f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa344_y4 = f_s_dadda_rca24_fa344_y4;
  assign f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa343_y4 = f_s_dadda_rca24_fa343_y4;
  assign f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa75_y2 = f_s_dadda_rca24_fa75_y2;
  assign f_s_dadda_rca24_fa345_y0 = f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa344_y4 ^ f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa343_y4;
  assign f_s_dadda_rca24_fa345_y1 = f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa344_y4 & f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa343_y4;
  assign f_s_dadda_rca24_fa345_y2 = f_s_dadda_rca24_fa345_y0 ^ f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa75_y2;
  assign f_s_dadda_rca24_fa345_y3 = f_s_dadda_rca24_fa345_y0 & f_s_dadda_rca24_fa345_f_s_dadda_rca24_fa75_y2;
  assign f_s_dadda_rca24_fa345_y4 = f_s_dadda_rca24_fa345_y1 | f_s_dadda_rca24_fa345_y3;
  assign f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa76_y2 = f_s_dadda_rca24_fa76_y2;
  assign f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa77_y2 = f_s_dadda_rca24_fa77_y2;
  assign f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa78_y2 = f_s_dadda_rca24_fa78_y2;
  assign f_s_dadda_rca24_fa346_y0 = f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa76_y2 ^ f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa77_y2;
  assign f_s_dadda_rca24_fa346_y1 = f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa76_y2 & f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa77_y2;
  assign f_s_dadda_rca24_fa346_y2 = f_s_dadda_rca24_fa346_y0 ^ f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa78_y2;
  assign f_s_dadda_rca24_fa346_y3 = f_s_dadda_rca24_fa346_y0 & f_s_dadda_rca24_fa346_f_s_dadda_rca24_fa78_y2;
  assign f_s_dadda_rca24_fa346_y4 = f_s_dadda_rca24_fa346_y1 | f_s_dadda_rca24_fa346_y3;
  assign f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa346_y4 = f_s_dadda_rca24_fa346_y4;
  assign f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa345_y4 = f_s_dadda_rca24_fa345_y4;
  assign f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa86_y2 = f_s_dadda_rca24_fa86_y2;
  assign f_s_dadda_rca24_fa347_y0 = f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa346_y4 ^ f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa345_y4;
  assign f_s_dadda_rca24_fa347_y1 = f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa346_y4 & f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa345_y4;
  assign f_s_dadda_rca24_fa347_y2 = f_s_dadda_rca24_fa347_y0 ^ f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa86_y2;
  assign f_s_dadda_rca24_fa347_y3 = f_s_dadda_rca24_fa347_y0 & f_s_dadda_rca24_fa347_f_s_dadda_rca24_fa86_y2;
  assign f_s_dadda_rca24_fa347_y4 = f_s_dadda_rca24_fa347_y1 | f_s_dadda_rca24_fa347_y3;
  assign f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa87_y2 = f_s_dadda_rca24_fa87_y2;
  assign f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa88_y2 = f_s_dadda_rca24_fa88_y2;
  assign f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa89_y2 = f_s_dadda_rca24_fa89_y2;
  assign f_s_dadda_rca24_fa348_y0 = f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa87_y2 ^ f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa88_y2;
  assign f_s_dadda_rca24_fa348_y1 = f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa87_y2 & f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa88_y2;
  assign f_s_dadda_rca24_fa348_y2 = f_s_dadda_rca24_fa348_y0 ^ f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa89_y2;
  assign f_s_dadda_rca24_fa348_y3 = f_s_dadda_rca24_fa348_y0 & f_s_dadda_rca24_fa348_f_s_dadda_rca24_fa89_y2;
  assign f_s_dadda_rca24_fa348_y4 = f_s_dadda_rca24_fa348_y1 | f_s_dadda_rca24_fa348_y3;
  assign f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa348_y4 = f_s_dadda_rca24_fa348_y4;
  assign f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa347_y4 = f_s_dadda_rca24_fa347_y4;
  assign f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa98_y2 = f_s_dadda_rca24_fa98_y2;
  assign f_s_dadda_rca24_fa349_y0 = f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa348_y4 ^ f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa347_y4;
  assign f_s_dadda_rca24_fa349_y1 = f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa348_y4 & f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa347_y4;
  assign f_s_dadda_rca24_fa349_y2 = f_s_dadda_rca24_fa349_y0 ^ f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa98_y2;
  assign f_s_dadda_rca24_fa349_y3 = f_s_dadda_rca24_fa349_y0 & f_s_dadda_rca24_fa349_f_s_dadda_rca24_fa98_y2;
  assign f_s_dadda_rca24_fa349_y4 = f_s_dadda_rca24_fa349_y1 | f_s_dadda_rca24_fa349_y3;
  assign f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa99_y2 = f_s_dadda_rca24_fa99_y2;
  assign f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa100_y2 = f_s_dadda_rca24_fa100_y2;
  assign f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa101_y2 = f_s_dadda_rca24_fa101_y2;
  assign f_s_dadda_rca24_fa350_y0 = f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa99_y2 ^ f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa100_y2;
  assign f_s_dadda_rca24_fa350_y1 = f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa99_y2 & f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa100_y2;
  assign f_s_dadda_rca24_fa350_y2 = f_s_dadda_rca24_fa350_y0 ^ f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa101_y2;
  assign f_s_dadda_rca24_fa350_y3 = f_s_dadda_rca24_fa350_y0 & f_s_dadda_rca24_fa350_f_s_dadda_rca24_fa101_y2;
  assign f_s_dadda_rca24_fa350_y4 = f_s_dadda_rca24_fa350_y1 | f_s_dadda_rca24_fa350_y3;
  assign f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa350_y4 = f_s_dadda_rca24_fa350_y4;
  assign f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa349_y4 = f_s_dadda_rca24_fa349_y4;
  assign f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa110_y2 = f_s_dadda_rca24_fa110_y2;
  assign f_s_dadda_rca24_fa351_y0 = f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa350_y4 ^ f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa349_y4;
  assign f_s_dadda_rca24_fa351_y1 = f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa350_y4 & f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa349_y4;
  assign f_s_dadda_rca24_fa351_y2 = f_s_dadda_rca24_fa351_y0 ^ f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa110_y2;
  assign f_s_dadda_rca24_fa351_y3 = f_s_dadda_rca24_fa351_y0 & f_s_dadda_rca24_fa351_f_s_dadda_rca24_fa110_y2;
  assign f_s_dadda_rca24_fa351_y4 = f_s_dadda_rca24_fa351_y1 | f_s_dadda_rca24_fa351_y3;
  assign f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa111_y2 = f_s_dadda_rca24_fa111_y2;
  assign f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa112_y2 = f_s_dadda_rca24_fa112_y2;
  assign f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa113_y2 = f_s_dadda_rca24_fa113_y2;
  assign f_s_dadda_rca24_fa352_y0 = f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa111_y2 ^ f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa112_y2;
  assign f_s_dadda_rca24_fa352_y1 = f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa111_y2 & f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa112_y2;
  assign f_s_dadda_rca24_fa352_y2 = f_s_dadda_rca24_fa352_y0 ^ f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa113_y2;
  assign f_s_dadda_rca24_fa352_y3 = f_s_dadda_rca24_fa352_y0 & f_s_dadda_rca24_fa352_f_s_dadda_rca24_fa113_y2;
  assign f_s_dadda_rca24_fa352_y4 = f_s_dadda_rca24_fa352_y1 | f_s_dadda_rca24_fa352_y3;
  assign f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa352_y4 = f_s_dadda_rca24_fa352_y4;
  assign f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa351_y4 = f_s_dadda_rca24_fa351_y4;
  assign f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa123_y2 = f_s_dadda_rca24_fa123_y2;
  assign f_s_dadda_rca24_fa353_y0 = f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa352_y4 ^ f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa351_y4;
  assign f_s_dadda_rca24_fa353_y1 = f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa352_y4 & f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa351_y4;
  assign f_s_dadda_rca24_fa353_y2 = f_s_dadda_rca24_fa353_y0 ^ f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa123_y2;
  assign f_s_dadda_rca24_fa353_y3 = f_s_dadda_rca24_fa353_y0 & f_s_dadda_rca24_fa353_f_s_dadda_rca24_fa123_y2;
  assign f_s_dadda_rca24_fa353_y4 = f_s_dadda_rca24_fa353_y1 | f_s_dadda_rca24_fa353_y3;
  assign f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa124_y2 = f_s_dadda_rca24_fa124_y2;
  assign f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa125_y2 = f_s_dadda_rca24_fa125_y2;
  assign f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa126_y2 = f_s_dadda_rca24_fa126_y2;
  assign f_s_dadda_rca24_fa354_y0 = f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa124_y2 ^ f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa125_y2;
  assign f_s_dadda_rca24_fa354_y1 = f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa124_y2 & f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa125_y2;
  assign f_s_dadda_rca24_fa354_y2 = f_s_dadda_rca24_fa354_y0 ^ f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa126_y2;
  assign f_s_dadda_rca24_fa354_y3 = f_s_dadda_rca24_fa354_y0 & f_s_dadda_rca24_fa354_f_s_dadda_rca24_fa126_y2;
  assign f_s_dadda_rca24_fa354_y4 = f_s_dadda_rca24_fa354_y1 | f_s_dadda_rca24_fa354_y3;
  assign f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa354_y4 = f_s_dadda_rca24_fa354_y4;
  assign f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa353_y4 = f_s_dadda_rca24_fa353_y4;
  assign f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa136_y2 = f_s_dadda_rca24_fa136_y2;
  assign f_s_dadda_rca24_fa355_y0 = f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa354_y4 ^ f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa353_y4;
  assign f_s_dadda_rca24_fa355_y1 = f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa354_y4 & f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa353_y4;
  assign f_s_dadda_rca24_fa355_y2 = f_s_dadda_rca24_fa355_y0 ^ f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa136_y2;
  assign f_s_dadda_rca24_fa355_y3 = f_s_dadda_rca24_fa355_y0 & f_s_dadda_rca24_fa355_f_s_dadda_rca24_fa136_y2;
  assign f_s_dadda_rca24_fa355_y4 = f_s_dadda_rca24_fa355_y1 | f_s_dadda_rca24_fa355_y3;
  assign f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa137_y2 = f_s_dadda_rca24_fa137_y2;
  assign f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa138_y2 = f_s_dadda_rca24_fa138_y2;
  assign f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa139_y2 = f_s_dadda_rca24_fa139_y2;
  assign f_s_dadda_rca24_fa356_y0 = f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa137_y2 ^ f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa138_y2;
  assign f_s_dadda_rca24_fa356_y1 = f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa137_y2 & f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa138_y2;
  assign f_s_dadda_rca24_fa356_y2 = f_s_dadda_rca24_fa356_y0 ^ f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa139_y2;
  assign f_s_dadda_rca24_fa356_y3 = f_s_dadda_rca24_fa356_y0 & f_s_dadda_rca24_fa356_f_s_dadda_rca24_fa139_y2;
  assign f_s_dadda_rca24_fa356_y4 = f_s_dadda_rca24_fa356_y1 | f_s_dadda_rca24_fa356_y3;
  assign f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa356_y4 = f_s_dadda_rca24_fa356_y4;
  assign f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa355_y4 = f_s_dadda_rca24_fa355_y4;
  assign f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa149_y2 = f_s_dadda_rca24_fa149_y2;
  assign f_s_dadda_rca24_fa357_y0 = f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa356_y4 ^ f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa355_y4;
  assign f_s_dadda_rca24_fa357_y1 = f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa356_y4 & f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa355_y4;
  assign f_s_dadda_rca24_fa357_y2 = f_s_dadda_rca24_fa357_y0 ^ f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa149_y2;
  assign f_s_dadda_rca24_fa357_y3 = f_s_dadda_rca24_fa357_y0 & f_s_dadda_rca24_fa357_f_s_dadda_rca24_fa149_y2;
  assign f_s_dadda_rca24_fa357_y4 = f_s_dadda_rca24_fa357_y1 | f_s_dadda_rca24_fa357_y3;
  assign f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa150_y2 = f_s_dadda_rca24_fa150_y2;
  assign f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa151_y2 = f_s_dadda_rca24_fa151_y2;
  assign f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa152_y2 = f_s_dadda_rca24_fa152_y2;
  assign f_s_dadda_rca24_fa358_y0 = f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa150_y2 ^ f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa151_y2;
  assign f_s_dadda_rca24_fa358_y1 = f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa150_y2 & f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa151_y2;
  assign f_s_dadda_rca24_fa358_y2 = f_s_dadda_rca24_fa358_y0 ^ f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa152_y2;
  assign f_s_dadda_rca24_fa358_y3 = f_s_dadda_rca24_fa358_y0 & f_s_dadda_rca24_fa358_f_s_dadda_rca24_fa152_y2;
  assign f_s_dadda_rca24_fa358_y4 = f_s_dadda_rca24_fa358_y1 | f_s_dadda_rca24_fa358_y3;
  assign f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa358_y4 = f_s_dadda_rca24_fa358_y4;
  assign f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa357_y4 = f_s_dadda_rca24_fa357_y4;
  assign f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa162_y2 = f_s_dadda_rca24_fa162_y2;
  assign f_s_dadda_rca24_fa359_y0 = f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa358_y4 ^ f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa357_y4;
  assign f_s_dadda_rca24_fa359_y1 = f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa358_y4 & f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa357_y4;
  assign f_s_dadda_rca24_fa359_y2 = f_s_dadda_rca24_fa359_y0 ^ f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa162_y2;
  assign f_s_dadda_rca24_fa359_y3 = f_s_dadda_rca24_fa359_y0 & f_s_dadda_rca24_fa359_f_s_dadda_rca24_fa162_y2;
  assign f_s_dadda_rca24_fa359_y4 = f_s_dadda_rca24_fa359_y1 | f_s_dadda_rca24_fa359_y3;
  assign f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa163_y2 = f_s_dadda_rca24_fa163_y2;
  assign f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa164_y2 = f_s_dadda_rca24_fa164_y2;
  assign f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa165_y2 = f_s_dadda_rca24_fa165_y2;
  assign f_s_dadda_rca24_fa360_y0 = f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa163_y2 ^ f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa164_y2;
  assign f_s_dadda_rca24_fa360_y1 = f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa163_y2 & f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa164_y2;
  assign f_s_dadda_rca24_fa360_y2 = f_s_dadda_rca24_fa360_y0 ^ f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa165_y2;
  assign f_s_dadda_rca24_fa360_y3 = f_s_dadda_rca24_fa360_y0 & f_s_dadda_rca24_fa360_f_s_dadda_rca24_fa165_y2;
  assign f_s_dadda_rca24_fa360_y4 = f_s_dadda_rca24_fa360_y1 | f_s_dadda_rca24_fa360_y3;
  assign f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa360_y4 = f_s_dadda_rca24_fa360_y4;
  assign f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa359_y4 = f_s_dadda_rca24_fa359_y4;
  assign f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa175_y2 = f_s_dadda_rca24_fa175_y2;
  assign f_s_dadda_rca24_fa361_y0 = f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa360_y4 ^ f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa359_y4;
  assign f_s_dadda_rca24_fa361_y1 = f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa360_y4 & f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa359_y4;
  assign f_s_dadda_rca24_fa361_y2 = f_s_dadda_rca24_fa361_y0 ^ f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa175_y2;
  assign f_s_dadda_rca24_fa361_y3 = f_s_dadda_rca24_fa361_y0 & f_s_dadda_rca24_fa361_f_s_dadda_rca24_fa175_y2;
  assign f_s_dadda_rca24_fa361_y4 = f_s_dadda_rca24_fa361_y1 | f_s_dadda_rca24_fa361_y3;
  assign f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa176_y2 = f_s_dadda_rca24_fa176_y2;
  assign f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa177_y2 = f_s_dadda_rca24_fa177_y2;
  assign f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa178_y2 = f_s_dadda_rca24_fa178_y2;
  assign f_s_dadda_rca24_fa362_y0 = f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa176_y2 ^ f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa177_y2;
  assign f_s_dadda_rca24_fa362_y1 = f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa176_y2 & f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa177_y2;
  assign f_s_dadda_rca24_fa362_y2 = f_s_dadda_rca24_fa362_y0 ^ f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa178_y2;
  assign f_s_dadda_rca24_fa362_y3 = f_s_dadda_rca24_fa362_y0 & f_s_dadda_rca24_fa362_f_s_dadda_rca24_fa178_y2;
  assign f_s_dadda_rca24_fa362_y4 = f_s_dadda_rca24_fa362_y1 | f_s_dadda_rca24_fa362_y3;
  assign f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa362_y4 = f_s_dadda_rca24_fa362_y4;
  assign f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa361_y4 = f_s_dadda_rca24_fa361_y4;
  assign f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa188_y2 = f_s_dadda_rca24_fa188_y2;
  assign f_s_dadda_rca24_fa363_y0 = f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa362_y4 ^ f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa361_y4;
  assign f_s_dadda_rca24_fa363_y1 = f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa362_y4 & f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa361_y4;
  assign f_s_dadda_rca24_fa363_y2 = f_s_dadda_rca24_fa363_y0 ^ f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa188_y2;
  assign f_s_dadda_rca24_fa363_y3 = f_s_dadda_rca24_fa363_y0 & f_s_dadda_rca24_fa363_f_s_dadda_rca24_fa188_y2;
  assign f_s_dadda_rca24_fa363_y4 = f_s_dadda_rca24_fa363_y1 | f_s_dadda_rca24_fa363_y3;
  assign f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa189_y2 = f_s_dadda_rca24_fa189_y2;
  assign f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa190_y2 = f_s_dadda_rca24_fa190_y2;
  assign f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa191_y2 = f_s_dadda_rca24_fa191_y2;
  assign f_s_dadda_rca24_fa364_y0 = f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa189_y2 ^ f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa190_y2;
  assign f_s_dadda_rca24_fa364_y1 = f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa189_y2 & f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa190_y2;
  assign f_s_dadda_rca24_fa364_y2 = f_s_dadda_rca24_fa364_y0 ^ f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa191_y2;
  assign f_s_dadda_rca24_fa364_y3 = f_s_dadda_rca24_fa364_y0 & f_s_dadda_rca24_fa364_f_s_dadda_rca24_fa191_y2;
  assign f_s_dadda_rca24_fa364_y4 = f_s_dadda_rca24_fa364_y1 | f_s_dadda_rca24_fa364_y3;
  assign f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa364_y4 = f_s_dadda_rca24_fa364_y4;
  assign f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa363_y4 = f_s_dadda_rca24_fa363_y4;
  assign f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa201_y2 = f_s_dadda_rca24_fa201_y2;
  assign f_s_dadda_rca24_fa365_y0 = f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa364_y4 ^ f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa363_y4;
  assign f_s_dadda_rca24_fa365_y1 = f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa364_y4 & f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa363_y4;
  assign f_s_dadda_rca24_fa365_y2 = f_s_dadda_rca24_fa365_y0 ^ f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa201_y2;
  assign f_s_dadda_rca24_fa365_y3 = f_s_dadda_rca24_fa365_y0 & f_s_dadda_rca24_fa365_f_s_dadda_rca24_fa201_y2;
  assign f_s_dadda_rca24_fa365_y4 = f_s_dadda_rca24_fa365_y1 | f_s_dadda_rca24_fa365_y3;
  assign f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa202_y2 = f_s_dadda_rca24_fa202_y2;
  assign f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa203_y2 = f_s_dadda_rca24_fa203_y2;
  assign f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa204_y2 = f_s_dadda_rca24_fa204_y2;
  assign f_s_dadda_rca24_fa366_y0 = f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa202_y2 ^ f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa203_y2;
  assign f_s_dadda_rca24_fa366_y1 = f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa202_y2 & f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa203_y2;
  assign f_s_dadda_rca24_fa366_y2 = f_s_dadda_rca24_fa366_y0 ^ f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa204_y2;
  assign f_s_dadda_rca24_fa366_y3 = f_s_dadda_rca24_fa366_y0 & f_s_dadda_rca24_fa366_f_s_dadda_rca24_fa204_y2;
  assign f_s_dadda_rca24_fa366_y4 = f_s_dadda_rca24_fa366_y1 | f_s_dadda_rca24_fa366_y3;
  assign f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa366_y4 = f_s_dadda_rca24_fa366_y4;
  assign f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa365_y4 = f_s_dadda_rca24_fa365_y4;
  assign f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa214_y2 = f_s_dadda_rca24_fa214_y2;
  assign f_s_dadda_rca24_fa367_y0 = f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa366_y4 ^ f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa365_y4;
  assign f_s_dadda_rca24_fa367_y1 = f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa366_y4 & f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa365_y4;
  assign f_s_dadda_rca24_fa367_y2 = f_s_dadda_rca24_fa367_y0 ^ f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa214_y2;
  assign f_s_dadda_rca24_fa367_y3 = f_s_dadda_rca24_fa367_y0 & f_s_dadda_rca24_fa367_f_s_dadda_rca24_fa214_y2;
  assign f_s_dadda_rca24_fa367_y4 = f_s_dadda_rca24_fa367_y1 | f_s_dadda_rca24_fa367_y3;
  assign f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa215_y2 = f_s_dadda_rca24_fa215_y2;
  assign f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa216_y2 = f_s_dadda_rca24_fa216_y2;
  assign f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa217_y2 = f_s_dadda_rca24_fa217_y2;
  assign f_s_dadda_rca24_fa368_y0 = f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa215_y2 ^ f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa216_y2;
  assign f_s_dadda_rca24_fa368_y1 = f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa215_y2 & f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa216_y2;
  assign f_s_dadda_rca24_fa368_y2 = f_s_dadda_rca24_fa368_y0 ^ f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa217_y2;
  assign f_s_dadda_rca24_fa368_y3 = f_s_dadda_rca24_fa368_y0 & f_s_dadda_rca24_fa368_f_s_dadda_rca24_fa217_y2;
  assign f_s_dadda_rca24_fa368_y4 = f_s_dadda_rca24_fa368_y1 | f_s_dadda_rca24_fa368_y3;
  assign f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa368_y4 = f_s_dadda_rca24_fa368_y4;
  assign f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa367_y4 = f_s_dadda_rca24_fa367_y4;
  assign f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa227_y2 = f_s_dadda_rca24_fa227_y2;
  assign f_s_dadda_rca24_fa369_y0 = f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa368_y4 ^ f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa367_y4;
  assign f_s_dadda_rca24_fa369_y1 = f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa368_y4 & f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa367_y4;
  assign f_s_dadda_rca24_fa369_y2 = f_s_dadda_rca24_fa369_y0 ^ f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa227_y2;
  assign f_s_dadda_rca24_fa369_y3 = f_s_dadda_rca24_fa369_y0 & f_s_dadda_rca24_fa369_f_s_dadda_rca24_fa227_y2;
  assign f_s_dadda_rca24_fa369_y4 = f_s_dadda_rca24_fa369_y1 | f_s_dadda_rca24_fa369_y3;
  assign f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa228_y2 = f_s_dadda_rca24_fa228_y2;
  assign f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa229_y2 = f_s_dadda_rca24_fa229_y2;
  assign f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa230_y2 = f_s_dadda_rca24_fa230_y2;
  assign f_s_dadda_rca24_fa370_y0 = f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa228_y2 ^ f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa229_y2;
  assign f_s_dadda_rca24_fa370_y1 = f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa228_y2 & f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa229_y2;
  assign f_s_dadda_rca24_fa370_y2 = f_s_dadda_rca24_fa370_y0 ^ f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa230_y2;
  assign f_s_dadda_rca24_fa370_y3 = f_s_dadda_rca24_fa370_y0 & f_s_dadda_rca24_fa370_f_s_dadda_rca24_fa230_y2;
  assign f_s_dadda_rca24_fa370_y4 = f_s_dadda_rca24_fa370_y1 | f_s_dadda_rca24_fa370_y3;
  assign f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa370_y4 = f_s_dadda_rca24_fa370_y4;
  assign f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa369_y4 = f_s_dadda_rca24_fa369_y4;
  assign f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa240_y2 = f_s_dadda_rca24_fa240_y2;
  assign f_s_dadda_rca24_fa371_y0 = f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa370_y4 ^ f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa369_y4;
  assign f_s_dadda_rca24_fa371_y1 = f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa370_y4 & f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa369_y4;
  assign f_s_dadda_rca24_fa371_y2 = f_s_dadda_rca24_fa371_y0 ^ f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa240_y2;
  assign f_s_dadda_rca24_fa371_y3 = f_s_dadda_rca24_fa371_y0 & f_s_dadda_rca24_fa371_f_s_dadda_rca24_fa240_y2;
  assign f_s_dadda_rca24_fa371_y4 = f_s_dadda_rca24_fa371_y1 | f_s_dadda_rca24_fa371_y3;
  assign f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa241_y2 = f_s_dadda_rca24_fa241_y2;
  assign f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa242_y2 = f_s_dadda_rca24_fa242_y2;
  assign f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa243_y2 = f_s_dadda_rca24_fa243_y2;
  assign f_s_dadda_rca24_fa372_y0 = f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa241_y2 ^ f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa242_y2;
  assign f_s_dadda_rca24_fa372_y1 = f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa241_y2 & f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa242_y2;
  assign f_s_dadda_rca24_fa372_y2 = f_s_dadda_rca24_fa372_y0 ^ f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa243_y2;
  assign f_s_dadda_rca24_fa372_y3 = f_s_dadda_rca24_fa372_y0 & f_s_dadda_rca24_fa372_f_s_dadda_rca24_fa243_y2;
  assign f_s_dadda_rca24_fa372_y4 = f_s_dadda_rca24_fa372_y1 | f_s_dadda_rca24_fa372_y3;
  assign f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa372_y4 = f_s_dadda_rca24_fa372_y4;
  assign f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa371_y4 = f_s_dadda_rca24_fa371_y4;
  assign f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa252_y2 = f_s_dadda_rca24_fa252_y2;
  assign f_s_dadda_rca24_fa373_y0 = f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa372_y4 ^ f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa371_y4;
  assign f_s_dadda_rca24_fa373_y1 = f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa372_y4 & f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa371_y4;
  assign f_s_dadda_rca24_fa373_y2 = f_s_dadda_rca24_fa373_y0 ^ f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa252_y2;
  assign f_s_dadda_rca24_fa373_y3 = f_s_dadda_rca24_fa373_y0 & f_s_dadda_rca24_fa373_f_s_dadda_rca24_fa252_y2;
  assign f_s_dadda_rca24_fa373_y4 = f_s_dadda_rca24_fa373_y1 | f_s_dadda_rca24_fa373_y3;
  assign f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa253_y2 = f_s_dadda_rca24_fa253_y2;
  assign f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa254_y2 = f_s_dadda_rca24_fa254_y2;
  assign f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa255_y2 = f_s_dadda_rca24_fa255_y2;
  assign f_s_dadda_rca24_fa374_y0 = f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa253_y2 ^ f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa254_y2;
  assign f_s_dadda_rca24_fa374_y1 = f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa253_y2 & f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa254_y2;
  assign f_s_dadda_rca24_fa374_y2 = f_s_dadda_rca24_fa374_y0 ^ f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa255_y2;
  assign f_s_dadda_rca24_fa374_y3 = f_s_dadda_rca24_fa374_y0 & f_s_dadda_rca24_fa374_f_s_dadda_rca24_fa255_y2;
  assign f_s_dadda_rca24_fa374_y4 = f_s_dadda_rca24_fa374_y1 | f_s_dadda_rca24_fa374_y3;
  assign f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa374_y4 = f_s_dadda_rca24_fa374_y4;
  assign f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa373_y4 = f_s_dadda_rca24_fa373_y4;
  assign f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa263_y2 = f_s_dadda_rca24_fa263_y2;
  assign f_s_dadda_rca24_fa375_y0 = f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa374_y4 ^ f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa373_y4;
  assign f_s_dadda_rca24_fa375_y1 = f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa374_y4 & f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa373_y4;
  assign f_s_dadda_rca24_fa375_y2 = f_s_dadda_rca24_fa375_y0 ^ f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa263_y2;
  assign f_s_dadda_rca24_fa375_y3 = f_s_dadda_rca24_fa375_y0 & f_s_dadda_rca24_fa375_f_s_dadda_rca24_fa263_y2;
  assign f_s_dadda_rca24_fa375_y4 = f_s_dadda_rca24_fa375_y1 | f_s_dadda_rca24_fa375_y3;
  assign f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa264_y2 = f_s_dadda_rca24_fa264_y2;
  assign f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa265_y2 = f_s_dadda_rca24_fa265_y2;
  assign f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa266_y2 = f_s_dadda_rca24_fa266_y2;
  assign f_s_dadda_rca24_fa376_y0 = f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa264_y2 ^ f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa265_y2;
  assign f_s_dadda_rca24_fa376_y1 = f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa264_y2 & f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa265_y2;
  assign f_s_dadda_rca24_fa376_y2 = f_s_dadda_rca24_fa376_y0 ^ f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa266_y2;
  assign f_s_dadda_rca24_fa376_y3 = f_s_dadda_rca24_fa376_y0 & f_s_dadda_rca24_fa376_f_s_dadda_rca24_fa266_y2;
  assign f_s_dadda_rca24_fa376_y4 = f_s_dadda_rca24_fa376_y1 | f_s_dadda_rca24_fa376_y3;
  assign f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa376_y4 = f_s_dadda_rca24_fa376_y4;
  assign f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa375_y4 = f_s_dadda_rca24_fa375_y4;
  assign f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa273_y2 = f_s_dadda_rca24_fa273_y2;
  assign f_s_dadda_rca24_fa377_y0 = f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa376_y4 ^ f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa375_y4;
  assign f_s_dadda_rca24_fa377_y1 = f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa376_y4 & f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa375_y4;
  assign f_s_dadda_rca24_fa377_y2 = f_s_dadda_rca24_fa377_y0 ^ f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa273_y2;
  assign f_s_dadda_rca24_fa377_y3 = f_s_dadda_rca24_fa377_y0 & f_s_dadda_rca24_fa377_f_s_dadda_rca24_fa273_y2;
  assign f_s_dadda_rca24_fa377_y4 = f_s_dadda_rca24_fa377_y1 | f_s_dadda_rca24_fa377_y3;
  assign f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa274_y2 = f_s_dadda_rca24_fa274_y2;
  assign f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa275_y2 = f_s_dadda_rca24_fa275_y2;
  assign f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa276_y2 = f_s_dadda_rca24_fa276_y2;
  assign f_s_dadda_rca24_fa378_y0 = f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa274_y2 ^ f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa275_y2;
  assign f_s_dadda_rca24_fa378_y1 = f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa274_y2 & f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa275_y2;
  assign f_s_dadda_rca24_fa378_y2 = f_s_dadda_rca24_fa378_y0 ^ f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa276_y2;
  assign f_s_dadda_rca24_fa378_y3 = f_s_dadda_rca24_fa378_y0 & f_s_dadda_rca24_fa378_f_s_dadda_rca24_fa276_y2;
  assign f_s_dadda_rca24_fa378_y4 = f_s_dadda_rca24_fa378_y1 | f_s_dadda_rca24_fa378_y3;
  assign f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa378_y4 = f_s_dadda_rca24_fa378_y4;
  assign f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa377_y4 = f_s_dadda_rca24_fa377_y4;
  assign f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa282_y2 = f_s_dadda_rca24_fa282_y2;
  assign f_s_dadda_rca24_fa379_y0 = f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa378_y4 ^ f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa377_y4;
  assign f_s_dadda_rca24_fa379_y1 = f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa378_y4 & f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa377_y4;
  assign f_s_dadda_rca24_fa379_y2 = f_s_dadda_rca24_fa379_y0 ^ f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa282_y2;
  assign f_s_dadda_rca24_fa379_y3 = f_s_dadda_rca24_fa379_y0 & f_s_dadda_rca24_fa379_f_s_dadda_rca24_fa282_y2;
  assign f_s_dadda_rca24_fa379_y4 = f_s_dadda_rca24_fa379_y1 | f_s_dadda_rca24_fa379_y3;
  assign f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa283_y2 = f_s_dadda_rca24_fa283_y2;
  assign f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa284_y2 = f_s_dadda_rca24_fa284_y2;
  assign f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa285_y2 = f_s_dadda_rca24_fa285_y2;
  assign f_s_dadda_rca24_fa380_y0 = f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa283_y2 ^ f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa284_y2;
  assign f_s_dadda_rca24_fa380_y1 = f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa283_y2 & f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa284_y2;
  assign f_s_dadda_rca24_fa380_y2 = f_s_dadda_rca24_fa380_y0 ^ f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa285_y2;
  assign f_s_dadda_rca24_fa380_y3 = f_s_dadda_rca24_fa380_y0 & f_s_dadda_rca24_fa380_f_s_dadda_rca24_fa285_y2;
  assign f_s_dadda_rca24_fa380_y4 = f_s_dadda_rca24_fa380_y1 | f_s_dadda_rca24_fa380_y3;
  assign f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa380_y4 = f_s_dadda_rca24_fa380_y4;
  assign f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa379_y4 = f_s_dadda_rca24_fa379_y4;
  assign f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa290_y2 = f_s_dadda_rca24_fa290_y2;
  assign f_s_dadda_rca24_fa381_y0 = f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa380_y4 ^ f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa379_y4;
  assign f_s_dadda_rca24_fa381_y1 = f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa380_y4 & f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa379_y4;
  assign f_s_dadda_rca24_fa381_y2 = f_s_dadda_rca24_fa381_y0 ^ f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa290_y2;
  assign f_s_dadda_rca24_fa381_y3 = f_s_dadda_rca24_fa381_y0 & f_s_dadda_rca24_fa381_f_s_dadda_rca24_fa290_y2;
  assign f_s_dadda_rca24_fa381_y4 = f_s_dadda_rca24_fa381_y1 | f_s_dadda_rca24_fa381_y3;
  assign f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa291_y2 = f_s_dadda_rca24_fa291_y2;
  assign f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa292_y2 = f_s_dadda_rca24_fa292_y2;
  assign f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa293_y2 = f_s_dadda_rca24_fa293_y2;
  assign f_s_dadda_rca24_fa382_y0 = f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa291_y2 ^ f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa292_y2;
  assign f_s_dadda_rca24_fa382_y1 = f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa291_y2 & f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa292_y2;
  assign f_s_dadda_rca24_fa382_y2 = f_s_dadda_rca24_fa382_y0 ^ f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa293_y2;
  assign f_s_dadda_rca24_fa382_y3 = f_s_dadda_rca24_fa382_y0 & f_s_dadda_rca24_fa382_f_s_dadda_rca24_fa293_y2;
  assign f_s_dadda_rca24_fa382_y4 = f_s_dadda_rca24_fa382_y1 | f_s_dadda_rca24_fa382_y3;
  assign f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa382_y4 = f_s_dadda_rca24_fa382_y4;
  assign f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa381_y4 = f_s_dadda_rca24_fa381_y4;
  assign f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa297_y2 = f_s_dadda_rca24_fa297_y2;
  assign f_s_dadda_rca24_fa383_y0 = f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa382_y4 ^ f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa381_y4;
  assign f_s_dadda_rca24_fa383_y1 = f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa382_y4 & f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa381_y4;
  assign f_s_dadda_rca24_fa383_y2 = f_s_dadda_rca24_fa383_y0 ^ f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa297_y2;
  assign f_s_dadda_rca24_fa383_y3 = f_s_dadda_rca24_fa383_y0 & f_s_dadda_rca24_fa383_f_s_dadda_rca24_fa297_y2;
  assign f_s_dadda_rca24_fa383_y4 = f_s_dadda_rca24_fa383_y1 | f_s_dadda_rca24_fa383_y3;
  assign f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa298_y2 = f_s_dadda_rca24_fa298_y2;
  assign f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa299_y2 = f_s_dadda_rca24_fa299_y2;
  assign f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa300_y2 = f_s_dadda_rca24_fa300_y2;
  assign f_s_dadda_rca24_fa384_y0 = f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa298_y2 ^ f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa299_y2;
  assign f_s_dadda_rca24_fa384_y1 = f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa298_y2 & f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa299_y2;
  assign f_s_dadda_rca24_fa384_y2 = f_s_dadda_rca24_fa384_y0 ^ f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa300_y2;
  assign f_s_dadda_rca24_fa384_y3 = f_s_dadda_rca24_fa384_y0 & f_s_dadda_rca24_fa384_f_s_dadda_rca24_fa300_y2;
  assign f_s_dadda_rca24_fa384_y4 = f_s_dadda_rca24_fa384_y1 | f_s_dadda_rca24_fa384_y3;
  assign f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa384_y4 = f_s_dadda_rca24_fa384_y4;
  assign f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa383_y4 = f_s_dadda_rca24_fa383_y4;
  assign f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa303_y2 = f_s_dadda_rca24_fa303_y2;
  assign f_s_dadda_rca24_fa385_y0 = f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa384_y4 ^ f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa383_y4;
  assign f_s_dadda_rca24_fa385_y1 = f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa384_y4 & f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa383_y4;
  assign f_s_dadda_rca24_fa385_y2 = f_s_dadda_rca24_fa385_y0 ^ f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa303_y2;
  assign f_s_dadda_rca24_fa385_y3 = f_s_dadda_rca24_fa385_y0 & f_s_dadda_rca24_fa385_f_s_dadda_rca24_fa303_y2;
  assign f_s_dadda_rca24_fa385_y4 = f_s_dadda_rca24_fa385_y1 | f_s_dadda_rca24_fa385_y3;
  assign f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa304_y2 = f_s_dadda_rca24_fa304_y2;
  assign f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa305_y2 = f_s_dadda_rca24_fa305_y2;
  assign f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa306_y2 = f_s_dadda_rca24_fa306_y2;
  assign f_s_dadda_rca24_fa386_y0 = f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa304_y2 ^ f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa305_y2;
  assign f_s_dadda_rca24_fa386_y1 = f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa304_y2 & f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa305_y2;
  assign f_s_dadda_rca24_fa386_y2 = f_s_dadda_rca24_fa386_y0 ^ f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa306_y2;
  assign f_s_dadda_rca24_fa386_y3 = f_s_dadda_rca24_fa386_y0 & f_s_dadda_rca24_fa386_f_s_dadda_rca24_fa306_y2;
  assign f_s_dadda_rca24_fa386_y4 = f_s_dadda_rca24_fa386_y1 | f_s_dadda_rca24_fa386_y3;
  assign f_s_dadda_rca24_nand_14_23_a_14 = a_14;
  assign f_s_dadda_rca24_nand_14_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_14_23_y0 = ~(f_s_dadda_rca24_nand_14_23_a_14 & f_s_dadda_rca24_nand_14_23_b_23);
  assign f_s_dadda_rca24_fa387_f_s_dadda_rca24_fa386_y4 = f_s_dadda_rca24_fa386_y4;
  assign f_s_dadda_rca24_fa387_f_s_dadda_rca24_fa385_y4 = f_s_dadda_rca24_fa385_y4;
  assign f_s_dadda_rca24_fa387_f_s_dadda_rca24_nand_14_23_y0 = f_s_dadda_rca24_nand_14_23_y0;
  assign f_s_dadda_rca24_fa387_y0 = f_s_dadda_rca24_fa387_f_s_dadda_rca24_fa386_y4 ^ f_s_dadda_rca24_fa387_f_s_dadda_rca24_fa385_y4;
  assign f_s_dadda_rca24_fa387_y1 = f_s_dadda_rca24_fa387_f_s_dadda_rca24_fa386_y4 & f_s_dadda_rca24_fa387_f_s_dadda_rca24_fa385_y4;
  assign f_s_dadda_rca24_fa387_y2 = f_s_dadda_rca24_fa387_y0 ^ f_s_dadda_rca24_fa387_f_s_dadda_rca24_nand_14_23_y0;
  assign f_s_dadda_rca24_fa387_y3 = f_s_dadda_rca24_fa387_y0 & f_s_dadda_rca24_fa387_f_s_dadda_rca24_nand_14_23_y0;
  assign f_s_dadda_rca24_fa387_y4 = f_s_dadda_rca24_fa387_y1 | f_s_dadda_rca24_fa387_y3;
  assign f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa309_y2 = f_s_dadda_rca24_fa309_y2;
  assign f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa310_y2 = f_s_dadda_rca24_fa310_y2;
  assign f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa311_y2 = f_s_dadda_rca24_fa311_y2;
  assign f_s_dadda_rca24_fa388_y0 = f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa309_y2 ^ f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa310_y2;
  assign f_s_dadda_rca24_fa388_y1 = f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa309_y2 & f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa310_y2;
  assign f_s_dadda_rca24_fa388_y2 = f_s_dadda_rca24_fa388_y0 ^ f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa311_y2;
  assign f_s_dadda_rca24_fa388_y3 = f_s_dadda_rca24_fa388_y0 & f_s_dadda_rca24_fa388_f_s_dadda_rca24_fa311_y2;
  assign f_s_dadda_rca24_fa388_y4 = f_s_dadda_rca24_fa388_y1 | f_s_dadda_rca24_fa388_y3;
  assign f_s_dadda_rca24_and_16_22_a_16 = a_16;
  assign f_s_dadda_rca24_and_16_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_16_22_y0 = f_s_dadda_rca24_and_16_22_a_16 & f_s_dadda_rca24_and_16_22_b_22;
  assign f_s_dadda_rca24_fa389_f_s_dadda_rca24_fa388_y4 = f_s_dadda_rca24_fa388_y4;
  assign f_s_dadda_rca24_fa389_f_s_dadda_rca24_fa387_y4 = f_s_dadda_rca24_fa387_y4;
  assign f_s_dadda_rca24_fa389_f_s_dadda_rca24_and_16_22_y0 = f_s_dadda_rca24_and_16_22_y0;
  assign f_s_dadda_rca24_fa389_y0 = f_s_dadda_rca24_fa389_f_s_dadda_rca24_fa388_y4 ^ f_s_dadda_rca24_fa389_f_s_dadda_rca24_fa387_y4;
  assign f_s_dadda_rca24_fa389_y1 = f_s_dadda_rca24_fa389_f_s_dadda_rca24_fa388_y4 & f_s_dadda_rca24_fa389_f_s_dadda_rca24_fa387_y4;
  assign f_s_dadda_rca24_fa389_y2 = f_s_dadda_rca24_fa389_y0 ^ f_s_dadda_rca24_fa389_f_s_dadda_rca24_and_16_22_y0;
  assign f_s_dadda_rca24_fa389_y3 = f_s_dadda_rca24_fa389_y0 & f_s_dadda_rca24_fa389_f_s_dadda_rca24_and_16_22_y0;
  assign f_s_dadda_rca24_fa389_y4 = f_s_dadda_rca24_fa389_y1 | f_s_dadda_rca24_fa389_y3;
  assign f_s_dadda_rca24_nand_15_23_a_15 = a_15;
  assign f_s_dadda_rca24_nand_15_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_15_23_y0 = ~(f_s_dadda_rca24_nand_15_23_a_15 & f_s_dadda_rca24_nand_15_23_b_23);
  assign f_s_dadda_rca24_fa390_f_s_dadda_rca24_nand_15_23_y0 = f_s_dadda_rca24_nand_15_23_y0;
  assign f_s_dadda_rca24_fa390_f_s_dadda_rca24_fa314_y2 = f_s_dadda_rca24_fa314_y2;
  assign f_s_dadda_rca24_fa390_f_s_dadda_rca24_fa315_y2 = f_s_dadda_rca24_fa315_y2;
  assign f_s_dadda_rca24_fa390_y0 = f_s_dadda_rca24_fa390_f_s_dadda_rca24_nand_15_23_y0 ^ f_s_dadda_rca24_fa390_f_s_dadda_rca24_fa314_y2;
  assign f_s_dadda_rca24_fa390_y1 = f_s_dadda_rca24_fa390_f_s_dadda_rca24_nand_15_23_y0 & f_s_dadda_rca24_fa390_f_s_dadda_rca24_fa314_y2;
  assign f_s_dadda_rca24_fa390_y2 = f_s_dadda_rca24_fa390_y0 ^ f_s_dadda_rca24_fa390_f_s_dadda_rca24_fa315_y2;
  assign f_s_dadda_rca24_fa390_y3 = f_s_dadda_rca24_fa390_y0 & f_s_dadda_rca24_fa390_f_s_dadda_rca24_fa315_y2;
  assign f_s_dadda_rca24_fa390_y4 = f_s_dadda_rca24_fa390_y1 | f_s_dadda_rca24_fa390_y3;
  assign f_s_dadda_rca24_and_18_21_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_18_21_y0 = f_s_dadda_rca24_and_18_21_a_18 & f_s_dadda_rca24_and_18_21_b_21;
  assign f_s_dadda_rca24_fa391_f_s_dadda_rca24_fa390_y4 = f_s_dadda_rca24_fa390_y4;
  assign f_s_dadda_rca24_fa391_f_s_dadda_rca24_fa389_y4 = f_s_dadda_rca24_fa389_y4;
  assign f_s_dadda_rca24_fa391_f_s_dadda_rca24_and_18_21_y0 = f_s_dadda_rca24_and_18_21_y0;
  assign f_s_dadda_rca24_fa391_y0 = f_s_dadda_rca24_fa391_f_s_dadda_rca24_fa390_y4 ^ f_s_dadda_rca24_fa391_f_s_dadda_rca24_fa389_y4;
  assign f_s_dadda_rca24_fa391_y1 = f_s_dadda_rca24_fa391_f_s_dadda_rca24_fa390_y4 & f_s_dadda_rca24_fa391_f_s_dadda_rca24_fa389_y4;
  assign f_s_dadda_rca24_fa391_y2 = f_s_dadda_rca24_fa391_y0 ^ f_s_dadda_rca24_fa391_f_s_dadda_rca24_and_18_21_y0;
  assign f_s_dadda_rca24_fa391_y3 = f_s_dadda_rca24_fa391_y0 & f_s_dadda_rca24_fa391_f_s_dadda_rca24_and_18_21_y0;
  assign f_s_dadda_rca24_fa391_y4 = f_s_dadda_rca24_fa391_y1 | f_s_dadda_rca24_fa391_y3;
  assign f_s_dadda_rca24_and_17_22_a_17 = a_17;
  assign f_s_dadda_rca24_and_17_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_17_22_y0 = f_s_dadda_rca24_and_17_22_a_17 & f_s_dadda_rca24_and_17_22_b_22;
  assign f_s_dadda_rca24_nand_16_23_a_16 = a_16;
  assign f_s_dadda_rca24_nand_16_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_16_23_y0 = ~(f_s_dadda_rca24_nand_16_23_a_16 & f_s_dadda_rca24_nand_16_23_b_23);
  assign f_s_dadda_rca24_fa392_f_s_dadda_rca24_and_17_22_y0 = f_s_dadda_rca24_and_17_22_y0;
  assign f_s_dadda_rca24_fa392_f_s_dadda_rca24_nand_16_23_y0 = f_s_dadda_rca24_nand_16_23_y0;
  assign f_s_dadda_rca24_fa392_f_s_dadda_rca24_fa318_y2 = f_s_dadda_rca24_fa318_y2;
  assign f_s_dadda_rca24_fa392_y0 = f_s_dadda_rca24_fa392_f_s_dadda_rca24_and_17_22_y0 ^ f_s_dadda_rca24_fa392_f_s_dadda_rca24_nand_16_23_y0;
  assign f_s_dadda_rca24_fa392_y1 = f_s_dadda_rca24_fa392_f_s_dadda_rca24_and_17_22_y0 & f_s_dadda_rca24_fa392_f_s_dadda_rca24_nand_16_23_y0;
  assign f_s_dadda_rca24_fa392_y2 = f_s_dadda_rca24_fa392_y0 ^ f_s_dadda_rca24_fa392_f_s_dadda_rca24_fa318_y2;
  assign f_s_dadda_rca24_fa392_y3 = f_s_dadda_rca24_fa392_y0 & f_s_dadda_rca24_fa392_f_s_dadda_rca24_fa318_y2;
  assign f_s_dadda_rca24_fa392_y4 = f_s_dadda_rca24_fa392_y1 | f_s_dadda_rca24_fa392_y3;
  assign f_s_dadda_rca24_and_20_20_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_20_20_y0 = f_s_dadda_rca24_and_20_20_a_20 & f_s_dadda_rca24_and_20_20_b_20;
  assign f_s_dadda_rca24_fa393_f_s_dadda_rca24_fa392_y4 = f_s_dadda_rca24_fa392_y4;
  assign f_s_dadda_rca24_fa393_f_s_dadda_rca24_fa391_y4 = f_s_dadda_rca24_fa391_y4;
  assign f_s_dadda_rca24_fa393_f_s_dadda_rca24_and_20_20_y0 = f_s_dadda_rca24_and_20_20_y0;
  assign f_s_dadda_rca24_fa393_y0 = f_s_dadda_rca24_fa393_f_s_dadda_rca24_fa392_y4 ^ f_s_dadda_rca24_fa393_f_s_dadda_rca24_fa391_y4;
  assign f_s_dadda_rca24_fa393_y1 = f_s_dadda_rca24_fa393_f_s_dadda_rca24_fa392_y4 & f_s_dadda_rca24_fa393_f_s_dadda_rca24_fa391_y4;
  assign f_s_dadda_rca24_fa393_y2 = f_s_dadda_rca24_fa393_y0 ^ f_s_dadda_rca24_fa393_f_s_dadda_rca24_and_20_20_y0;
  assign f_s_dadda_rca24_fa393_y3 = f_s_dadda_rca24_fa393_y0 & f_s_dadda_rca24_fa393_f_s_dadda_rca24_and_20_20_y0;
  assign f_s_dadda_rca24_fa393_y4 = f_s_dadda_rca24_fa393_y1 | f_s_dadda_rca24_fa393_y3;
  assign f_s_dadda_rca24_and_19_21_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_19_21_y0 = f_s_dadda_rca24_and_19_21_a_19 & f_s_dadda_rca24_and_19_21_b_21;
  assign f_s_dadda_rca24_and_18_22_a_18 = a_18;
  assign f_s_dadda_rca24_and_18_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_18_22_y0 = f_s_dadda_rca24_and_18_22_a_18 & f_s_dadda_rca24_and_18_22_b_22;
  assign f_s_dadda_rca24_nand_17_23_a_17 = a_17;
  assign f_s_dadda_rca24_nand_17_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_17_23_y0 = ~(f_s_dadda_rca24_nand_17_23_a_17 & f_s_dadda_rca24_nand_17_23_b_23);
  assign f_s_dadda_rca24_fa394_f_s_dadda_rca24_and_19_21_y0 = f_s_dadda_rca24_and_19_21_y0;
  assign f_s_dadda_rca24_fa394_f_s_dadda_rca24_and_18_22_y0 = f_s_dadda_rca24_and_18_22_y0;
  assign f_s_dadda_rca24_fa394_f_s_dadda_rca24_nand_17_23_y0 = f_s_dadda_rca24_nand_17_23_y0;
  assign f_s_dadda_rca24_fa394_y0 = f_s_dadda_rca24_fa394_f_s_dadda_rca24_and_19_21_y0 ^ f_s_dadda_rca24_fa394_f_s_dadda_rca24_and_18_22_y0;
  assign f_s_dadda_rca24_fa394_y1 = f_s_dadda_rca24_fa394_f_s_dadda_rca24_and_19_21_y0 & f_s_dadda_rca24_fa394_f_s_dadda_rca24_and_18_22_y0;
  assign f_s_dadda_rca24_fa394_y2 = f_s_dadda_rca24_fa394_y0 ^ f_s_dadda_rca24_fa394_f_s_dadda_rca24_nand_17_23_y0;
  assign f_s_dadda_rca24_fa394_y3 = f_s_dadda_rca24_fa394_y0 & f_s_dadda_rca24_fa394_f_s_dadda_rca24_nand_17_23_y0;
  assign f_s_dadda_rca24_fa394_y4 = f_s_dadda_rca24_fa394_y1 | f_s_dadda_rca24_fa394_y3;
  assign f_s_dadda_rca24_and_22_19_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_19_b_19 = b_19;
  assign f_s_dadda_rca24_and_22_19_y0 = f_s_dadda_rca24_and_22_19_a_22 & f_s_dadda_rca24_and_22_19_b_19;
  assign f_s_dadda_rca24_fa395_f_s_dadda_rca24_fa394_y4 = f_s_dadda_rca24_fa394_y4;
  assign f_s_dadda_rca24_fa395_f_s_dadda_rca24_fa393_y4 = f_s_dadda_rca24_fa393_y4;
  assign f_s_dadda_rca24_fa395_f_s_dadda_rca24_and_22_19_y0 = f_s_dadda_rca24_and_22_19_y0;
  assign f_s_dadda_rca24_fa395_y0 = f_s_dadda_rca24_fa395_f_s_dadda_rca24_fa394_y4 ^ f_s_dadda_rca24_fa395_f_s_dadda_rca24_fa393_y4;
  assign f_s_dadda_rca24_fa395_y1 = f_s_dadda_rca24_fa395_f_s_dadda_rca24_fa394_y4 & f_s_dadda_rca24_fa395_f_s_dadda_rca24_fa393_y4;
  assign f_s_dadda_rca24_fa395_y2 = f_s_dadda_rca24_fa395_y0 ^ f_s_dadda_rca24_fa395_f_s_dadda_rca24_and_22_19_y0;
  assign f_s_dadda_rca24_fa395_y3 = f_s_dadda_rca24_fa395_y0 & f_s_dadda_rca24_fa395_f_s_dadda_rca24_and_22_19_y0;
  assign f_s_dadda_rca24_fa395_y4 = f_s_dadda_rca24_fa395_y1 | f_s_dadda_rca24_fa395_y3;
  assign f_s_dadda_rca24_and_21_20_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_21_20_y0 = f_s_dadda_rca24_and_21_20_a_21 & f_s_dadda_rca24_and_21_20_b_20;
  assign f_s_dadda_rca24_and_20_21_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_20_21_y0 = f_s_dadda_rca24_and_20_21_a_20 & f_s_dadda_rca24_and_20_21_b_21;
  assign f_s_dadda_rca24_and_19_22_a_19 = a_19;
  assign f_s_dadda_rca24_and_19_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_19_22_y0 = f_s_dadda_rca24_and_19_22_a_19 & f_s_dadda_rca24_and_19_22_b_22;
  assign f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_21_20_y0 = f_s_dadda_rca24_and_21_20_y0;
  assign f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_20_21_y0 = f_s_dadda_rca24_and_20_21_y0;
  assign f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_19_22_y0 = f_s_dadda_rca24_and_19_22_y0;
  assign f_s_dadda_rca24_fa396_y0 = f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_21_20_y0 ^ f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_20_21_y0;
  assign f_s_dadda_rca24_fa396_y1 = f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_21_20_y0 & f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_20_21_y0;
  assign f_s_dadda_rca24_fa396_y2 = f_s_dadda_rca24_fa396_y0 ^ f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_19_22_y0;
  assign f_s_dadda_rca24_fa396_y3 = f_s_dadda_rca24_fa396_y0 & f_s_dadda_rca24_fa396_f_s_dadda_rca24_and_19_22_y0;
  assign f_s_dadda_rca24_fa396_y4 = f_s_dadda_rca24_fa396_y1 | f_s_dadda_rca24_fa396_y3;
  assign f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa396_y4 = f_s_dadda_rca24_fa396_y4;
  assign f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa395_y4 = f_s_dadda_rca24_fa395_y4;
  assign f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa323_y4 = f_s_dadda_rca24_fa323_y4;
  assign f_s_dadda_rca24_fa397_y0 = f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa396_y4 ^ f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa395_y4;
  assign f_s_dadda_rca24_fa397_y1 = f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa396_y4 & f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa395_y4;
  assign f_s_dadda_rca24_fa397_y2 = f_s_dadda_rca24_fa397_y0 ^ f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa323_y4;
  assign f_s_dadda_rca24_fa397_y3 = f_s_dadda_rca24_fa397_y0 & f_s_dadda_rca24_fa397_f_s_dadda_rca24_fa323_y4;
  assign f_s_dadda_rca24_fa397_y4 = f_s_dadda_rca24_fa397_y1 | f_s_dadda_rca24_fa397_y3;
  assign f_s_dadda_rca24_nand_23_19_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_19_b_19 = b_19;
  assign f_s_dadda_rca24_nand_23_19_y0 = ~(f_s_dadda_rca24_nand_23_19_a_23 & f_s_dadda_rca24_nand_23_19_b_19);
  assign f_s_dadda_rca24_and_22_20_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_20_b_20 = b_20;
  assign f_s_dadda_rca24_and_22_20_y0 = f_s_dadda_rca24_and_22_20_a_22 & f_s_dadda_rca24_and_22_20_b_20;
  assign f_s_dadda_rca24_and_21_21_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_21_21_y0 = f_s_dadda_rca24_and_21_21_a_21 & f_s_dadda_rca24_and_21_21_b_21;
  assign f_s_dadda_rca24_fa398_f_s_dadda_rca24_nand_23_19_y0 = f_s_dadda_rca24_nand_23_19_y0;
  assign f_s_dadda_rca24_fa398_f_s_dadda_rca24_and_22_20_y0 = f_s_dadda_rca24_and_22_20_y0;
  assign f_s_dadda_rca24_fa398_f_s_dadda_rca24_and_21_21_y0 = f_s_dadda_rca24_and_21_21_y0;
  assign f_s_dadda_rca24_fa398_y0 = f_s_dadda_rca24_fa398_f_s_dadda_rca24_nand_23_19_y0 ^ f_s_dadda_rca24_fa398_f_s_dadda_rca24_and_22_20_y0;
  assign f_s_dadda_rca24_fa398_y1 = f_s_dadda_rca24_fa398_f_s_dadda_rca24_nand_23_19_y0 & f_s_dadda_rca24_fa398_f_s_dadda_rca24_and_22_20_y0;
  assign f_s_dadda_rca24_fa398_y2 = f_s_dadda_rca24_fa398_y0 ^ f_s_dadda_rca24_fa398_f_s_dadda_rca24_and_21_21_y0;
  assign f_s_dadda_rca24_fa398_y3 = f_s_dadda_rca24_fa398_y0 & f_s_dadda_rca24_fa398_f_s_dadda_rca24_and_21_21_y0;
  assign f_s_dadda_rca24_fa398_y4 = f_s_dadda_rca24_fa398_y1 | f_s_dadda_rca24_fa398_y3;
  assign f_s_dadda_rca24_nand_23_20_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_20_b_20 = b_20;
  assign f_s_dadda_rca24_nand_23_20_y0 = ~(f_s_dadda_rca24_nand_23_20_a_23 & f_s_dadda_rca24_nand_23_20_b_20);
  assign f_s_dadda_rca24_fa399_f_s_dadda_rca24_fa398_y4 = f_s_dadda_rca24_fa398_y4;
  assign f_s_dadda_rca24_fa399_f_s_dadda_rca24_fa397_y4 = f_s_dadda_rca24_fa397_y4;
  assign f_s_dadda_rca24_fa399_f_s_dadda_rca24_nand_23_20_y0 = f_s_dadda_rca24_nand_23_20_y0;
  assign f_s_dadda_rca24_fa399_y0 = f_s_dadda_rca24_fa399_f_s_dadda_rca24_fa398_y4 ^ f_s_dadda_rca24_fa399_f_s_dadda_rca24_fa397_y4;
  assign f_s_dadda_rca24_fa399_y1 = f_s_dadda_rca24_fa399_f_s_dadda_rca24_fa398_y4 & f_s_dadda_rca24_fa399_f_s_dadda_rca24_fa397_y4;
  assign f_s_dadda_rca24_fa399_y2 = f_s_dadda_rca24_fa399_y0 ^ f_s_dadda_rca24_fa399_f_s_dadda_rca24_nand_23_20_y0;
  assign f_s_dadda_rca24_fa399_y3 = f_s_dadda_rca24_fa399_y0 & f_s_dadda_rca24_fa399_f_s_dadda_rca24_nand_23_20_y0;
  assign f_s_dadda_rca24_fa399_y4 = f_s_dadda_rca24_fa399_y1 | f_s_dadda_rca24_fa399_y3;
  assign f_s_dadda_rca24_and_3_0_a_3 = a_3;
  assign f_s_dadda_rca24_and_3_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_3_0_y0 = f_s_dadda_rca24_and_3_0_a_3 & f_s_dadda_rca24_and_3_0_b_0;
  assign f_s_dadda_rca24_and_2_1_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_2_1_y0 = f_s_dadda_rca24_and_2_1_a_2 & f_s_dadda_rca24_and_2_1_b_1;
  assign f_s_dadda_rca24_ha20_f_s_dadda_rca24_and_3_0_y0 = f_s_dadda_rca24_and_3_0_y0;
  assign f_s_dadda_rca24_ha20_f_s_dadda_rca24_and_2_1_y0 = f_s_dadda_rca24_and_2_1_y0;
  assign f_s_dadda_rca24_ha20_y0 = f_s_dadda_rca24_ha20_f_s_dadda_rca24_and_3_0_y0 ^ f_s_dadda_rca24_ha20_f_s_dadda_rca24_and_2_1_y0;
  assign f_s_dadda_rca24_ha20_y1 = f_s_dadda_rca24_ha20_f_s_dadda_rca24_and_3_0_y0 & f_s_dadda_rca24_ha20_f_s_dadda_rca24_and_2_1_y0;
  assign f_s_dadda_rca24_and_2_2_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_2_2_y0 = f_s_dadda_rca24_and_2_2_a_2 & f_s_dadda_rca24_and_2_2_b_2;
  assign f_s_dadda_rca24_and_1_3_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_1_3_y0 = f_s_dadda_rca24_and_1_3_a_1 & f_s_dadda_rca24_and_1_3_b_3;
  assign f_s_dadda_rca24_fa400_f_s_dadda_rca24_ha20_y1 = f_s_dadda_rca24_ha20_y1;
  assign f_s_dadda_rca24_fa400_f_s_dadda_rca24_and_2_2_y0 = f_s_dadda_rca24_and_2_2_y0;
  assign f_s_dadda_rca24_fa400_f_s_dadda_rca24_and_1_3_y0 = f_s_dadda_rca24_and_1_3_y0;
  assign f_s_dadda_rca24_fa400_y0 = f_s_dadda_rca24_fa400_f_s_dadda_rca24_ha20_y1 ^ f_s_dadda_rca24_fa400_f_s_dadda_rca24_and_2_2_y0;
  assign f_s_dadda_rca24_fa400_y1 = f_s_dadda_rca24_fa400_f_s_dadda_rca24_ha20_y1 & f_s_dadda_rca24_fa400_f_s_dadda_rca24_and_2_2_y0;
  assign f_s_dadda_rca24_fa400_y2 = f_s_dadda_rca24_fa400_y0 ^ f_s_dadda_rca24_fa400_f_s_dadda_rca24_and_1_3_y0;
  assign f_s_dadda_rca24_fa400_y3 = f_s_dadda_rca24_fa400_y0 & f_s_dadda_rca24_fa400_f_s_dadda_rca24_and_1_3_y0;
  assign f_s_dadda_rca24_fa400_y4 = f_s_dadda_rca24_fa400_y1 | f_s_dadda_rca24_fa400_y3;
  assign f_s_dadda_rca24_and_1_4_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_1_4_y0 = f_s_dadda_rca24_and_1_4_a_1 & f_s_dadda_rca24_and_1_4_b_4;
  assign f_s_dadda_rca24_and_0_5_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_5_b_5 = b_5;
  assign f_s_dadda_rca24_and_0_5_y0 = f_s_dadda_rca24_and_0_5_a_0 & f_s_dadda_rca24_and_0_5_b_5;
  assign f_s_dadda_rca24_fa401_f_s_dadda_rca24_fa400_y4 = f_s_dadda_rca24_fa400_y4;
  assign f_s_dadda_rca24_fa401_f_s_dadda_rca24_and_1_4_y0 = f_s_dadda_rca24_and_1_4_y0;
  assign f_s_dadda_rca24_fa401_f_s_dadda_rca24_and_0_5_y0 = f_s_dadda_rca24_and_0_5_y0;
  assign f_s_dadda_rca24_fa401_y0 = f_s_dadda_rca24_fa401_f_s_dadda_rca24_fa400_y4 ^ f_s_dadda_rca24_fa401_f_s_dadda_rca24_and_1_4_y0;
  assign f_s_dadda_rca24_fa401_y1 = f_s_dadda_rca24_fa401_f_s_dadda_rca24_fa400_y4 & f_s_dadda_rca24_fa401_f_s_dadda_rca24_and_1_4_y0;
  assign f_s_dadda_rca24_fa401_y2 = f_s_dadda_rca24_fa401_y0 ^ f_s_dadda_rca24_fa401_f_s_dadda_rca24_and_0_5_y0;
  assign f_s_dadda_rca24_fa401_y3 = f_s_dadda_rca24_fa401_y0 & f_s_dadda_rca24_fa401_f_s_dadda_rca24_and_0_5_y0;
  assign f_s_dadda_rca24_fa401_y4 = f_s_dadda_rca24_fa401_y1 | f_s_dadda_rca24_fa401_y3;
  assign f_s_dadda_rca24_and_0_6_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_6_b_6 = b_6;
  assign f_s_dadda_rca24_and_0_6_y0 = f_s_dadda_rca24_and_0_6_a_0 & f_s_dadda_rca24_and_0_6_b_6;
  assign f_s_dadda_rca24_fa402_f_s_dadda_rca24_fa401_y4 = f_s_dadda_rca24_fa401_y4;
  assign f_s_dadda_rca24_fa402_f_s_dadda_rca24_and_0_6_y0 = f_s_dadda_rca24_and_0_6_y0;
  assign f_s_dadda_rca24_fa402_f_s_dadda_rca24_ha5_y0 = f_s_dadda_rca24_ha5_y0;
  assign f_s_dadda_rca24_fa402_y0 = f_s_dadda_rca24_fa402_f_s_dadda_rca24_fa401_y4 ^ f_s_dadda_rca24_fa402_f_s_dadda_rca24_and_0_6_y0;
  assign f_s_dadda_rca24_fa402_y1 = f_s_dadda_rca24_fa402_f_s_dadda_rca24_fa401_y4 & f_s_dadda_rca24_fa402_f_s_dadda_rca24_and_0_6_y0;
  assign f_s_dadda_rca24_fa402_y2 = f_s_dadda_rca24_fa402_y0 ^ f_s_dadda_rca24_fa402_f_s_dadda_rca24_ha5_y0;
  assign f_s_dadda_rca24_fa402_y3 = f_s_dadda_rca24_fa402_y0 & f_s_dadda_rca24_fa402_f_s_dadda_rca24_ha5_y0;
  assign f_s_dadda_rca24_fa402_y4 = f_s_dadda_rca24_fa402_y1 | f_s_dadda_rca24_fa402_y3;
  assign f_s_dadda_rca24_fa403_f_s_dadda_rca24_fa402_y4 = f_s_dadda_rca24_fa402_y4;
  assign f_s_dadda_rca24_fa403_f_s_dadda_rca24_fa25_y2 = f_s_dadda_rca24_fa25_y2;
  assign f_s_dadda_rca24_fa403_f_s_dadda_rca24_ha6_y0 = f_s_dadda_rca24_ha6_y0;
  assign f_s_dadda_rca24_fa403_y0 = f_s_dadda_rca24_fa403_f_s_dadda_rca24_fa402_y4 ^ f_s_dadda_rca24_fa403_f_s_dadda_rca24_fa25_y2;
  assign f_s_dadda_rca24_fa403_y1 = f_s_dadda_rca24_fa403_f_s_dadda_rca24_fa402_y4 & f_s_dadda_rca24_fa403_f_s_dadda_rca24_fa25_y2;
  assign f_s_dadda_rca24_fa403_y2 = f_s_dadda_rca24_fa403_y0 ^ f_s_dadda_rca24_fa403_f_s_dadda_rca24_ha6_y0;
  assign f_s_dadda_rca24_fa403_y3 = f_s_dadda_rca24_fa403_y0 & f_s_dadda_rca24_fa403_f_s_dadda_rca24_ha6_y0;
  assign f_s_dadda_rca24_fa403_y4 = f_s_dadda_rca24_fa403_y1 | f_s_dadda_rca24_fa403_y3;
  assign f_s_dadda_rca24_fa404_f_s_dadda_rca24_fa403_y4 = f_s_dadda_rca24_fa403_y4;
  assign f_s_dadda_rca24_fa404_f_s_dadda_rca24_fa27_y2 = f_s_dadda_rca24_fa27_y2;
  assign f_s_dadda_rca24_fa404_f_s_dadda_rca24_ha7_y0 = f_s_dadda_rca24_ha7_y0;
  assign f_s_dadda_rca24_fa404_y0 = f_s_dadda_rca24_fa404_f_s_dadda_rca24_fa403_y4 ^ f_s_dadda_rca24_fa404_f_s_dadda_rca24_fa27_y2;
  assign f_s_dadda_rca24_fa404_y1 = f_s_dadda_rca24_fa404_f_s_dadda_rca24_fa403_y4 & f_s_dadda_rca24_fa404_f_s_dadda_rca24_fa27_y2;
  assign f_s_dadda_rca24_fa404_y2 = f_s_dadda_rca24_fa404_y0 ^ f_s_dadda_rca24_fa404_f_s_dadda_rca24_ha7_y0;
  assign f_s_dadda_rca24_fa404_y3 = f_s_dadda_rca24_fa404_y0 & f_s_dadda_rca24_fa404_f_s_dadda_rca24_ha7_y0;
  assign f_s_dadda_rca24_fa404_y4 = f_s_dadda_rca24_fa404_y1 | f_s_dadda_rca24_fa404_y3;
  assign f_s_dadda_rca24_fa405_f_s_dadda_rca24_fa404_y4 = f_s_dadda_rca24_fa404_y4;
  assign f_s_dadda_rca24_fa405_f_s_dadda_rca24_fa30_y2 = f_s_dadda_rca24_fa30_y2;
  assign f_s_dadda_rca24_fa405_f_s_dadda_rca24_ha8_y0 = f_s_dadda_rca24_ha8_y0;
  assign f_s_dadda_rca24_fa405_y0 = f_s_dadda_rca24_fa405_f_s_dadda_rca24_fa404_y4 ^ f_s_dadda_rca24_fa405_f_s_dadda_rca24_fa30_y2;
  assign f_s_dadda_rca24_fa405_y1 = f_s_dadda_rca24_fa405_f_s_dadda_rca24_fa404_y4 & f_s_dadda_rca24_fa405_f_s_dadda_rca24_fa30_y2;
  assign f_s_dadda_rca24_fa405_y2 = f_s_dadda_rca24_fa405_y0 ^ f_s_dadda_rca24_fa405_f_s_dadda_rca24_ha8_y0;
  assign f_s_dadda_rca24_fa405_y3 = f_s_dadda_rca24_fa405_y0 & f_s_dadda_rca24_fa405_f_s_dadda_rca24_ha8_y0;
  assign f_s_dadda_rca24_fa405_y4 = f_s_dadda_rca24_fa405_y1 | f_s_dadda_rca24_fa405_y3;
  assign f_s_dadda_rca24_fa406_f_s_dadda_rca24_fa405_y4 = f_s_dadda_rca24_fa405_y4;
  assign f_s_dadda_rca24_fa406_f_s_dadda_rca24_fa34_y2 = f_s_dadda_rca24_fa34_y2;
  assign f_s_dadda_rca24_fa406_f_s_dadda_rca24_ha9_y0 = f_s_dadda_rca24_ha9_y0;
  assign f_s_dadda_rca24_fa406_y0 = f_s_dadda_rca24_fa406_f_s_dadda_rca24_fa405_y4 ^ f_s_dadda_rca24_fa406_f_s_dadda_rca24_fa34_y2;
  assign f_s_dadda_rca24_fa406_y1 = f_s_dadda_rca24_fa406_f_s_dadda_rca24_fa405_y4 & f_s_dadda_rca24_fa406_f_s_dadda_rca24_fa34_y2;
  assign f_s_dadda_rca24_fa406_y2 = f_s_dadda_rca24_fa406_y0 ^ f_s_dadda_rca24_fa406_f_s_dadda_rca24_ha9_y0;
  assign f_s_dadda_rca24_fa406_y3 = f_s_dadda_rca24_fa406_y0 & f_s_dadda_rca24_fa406_f_s_dadda_rca24_ha9_y0;
  assign f_s_dadda_rca24_fa406_y4 = f_s_dadda_rca24_fa406_y1 | f_s_dadda_rca24_fa406_y3;
  assign f_s_dadda_rca24_fa407_f_s_dadda_rca24_fa406_y4 = f_s_dadda_rca24_fa406_y4;
  assign f_s_dadda_rca24_fa407_f_s_dadda_rca24_fa39_y2 = f_s_dadda_rca24_fa39_y2;
  assign f_s_dadda_rca24_fa407_f_s_dadda_rca24_ha10_y0 = f_s_dadda_rca24_ha10_y0;
  assign f_s_dadda_rca24_fa407_y0 = f_s_dadda_rca24_fa407_f_s_dadda_rca24_fa406_y4 ^ f_s_dadda_rca24_fa407_f_s_dadda_rca24_fa39_y2;
  assign f_s_dadda_rca24_fa407_y1 = f_s_dadda_rca24_fa407_f_s_dadda_rca24_fa406_y4 & f_s_dadda_rca24_fa407_f_s_dadda_rca24_fa39_y2;
  assign f_s_dadda_rca24_fa407_y2 = f_s_dadda_rca24_fa407_y0 ^ f_s_dadda_rca24_fa407_f_s_dadda_rca24_ha10_y0;
  assign f_s_dadda_rca24_fa407_y3 = f_s_dadda_rca24_fa407_y0 & f_s_dadda_rca24_fa407_f_s_dadda_rca24_ha10_y0;
  assign f_s_dadda_rca24_fa407_y4 = f_s_dadda_rca24_fa407_y1 | f_s_dadda_rca24_fa407_y3;
  assign f_s_dadda_rca24_fa408_f_s_dadda_rca24_fa407_y4 = f_s_dadda_rca24_fa407_y4;
  assign f_s_dadda_rca24_fa408_f_s_dadda_rca24_fa45_y2 = f_s_dadda_rca24_fa45_y2;
  assign f_s_dadda_rca24_fa408_f_s_dadda_rca24_ha11_y0 = f_s_dadda_rca24_ha11_y0;
  assign f_s_dadda_rca24_fa408_y0 = f_s_dadda_rca24_fa408_f_s_dadda_rca24_fa407_y4 ^ f_s_dadda_rca24_fa408_f_s_dadda_rca24_fa45_y2;
  assign f_s_dadda_rca24_fa408_y1 = f_s_dadda_rca24_fa408_f_s_dadda_rca24_fa407_y4 & f_s_dadda_rca24_fa408_f_s_dadda_rca24_fa45_y2;
  assign f_s_dadda_rca24_fa408_y2 = f_s_dadda_rca24_fa408_y0 ^ f_s_dadda_rca24_fa408_f_s_dadda_rca24_ha11_y0;
  assign f_s_dadda_rca24_fa408_y3 = f_s_dadda_rca24_fa408_y0 & f_s_dadda_rca24_fa408_f_s_dadda_rca24_ha11_y0;
  assign f_s_dadda_rca24_fa408_y4 = f_s_dadda_rca24_fa408_y1 | f_s_dadda_rca24_fa408_y3;
  assign f_s_dadda_rca24_fa409_f_s_dadda_rca24_fa408_y4 = f_s_dadda_rca24_fa408_y4;
  assign f_s_dadda_rca24_fa409_f_s_dadda_rca24_fa52_y2 = f_s_dadda_rca24_fa52_y2;
  assign f_s_dadda_rca24_fa409_f_s_dadda_rca24_ha12_y0 = f_s_dadda_rca24_ha12_y0;
  assign f_s_dadda_rca24_fa409_y0 = f_s_dadda_rca24_fa409_f_s_dadda_rca24_fa408_y4 ^ f_s_dadda_rca24_fa409_f_s_dadda_rca24_fa52_y2;
  assign f_s_dadda_rca24_fa409_y1 = f_s_dadda_rca24_fa409_f_s_dadda_rca24_fa408_y4 & f_s_dadda_rca24_fa409_f_s_dadda_rca24_fa52_y2;
  assign f_s_dadda_rca24_fa409_y2 = f_s_dadda_rca24_fa409_y0 ^ f_s_dadda_rca24_fa409_f_s_dadda_rca24_ha12_y0;
  assign f_s_dadda_rca24_fa409_y3 = f_s_dadda_rca24_fa409_y0 & f_s_dadda_rca24_fa409_f_s_dadda_rca24_ha12_y0;
  assign f_s_dadda_rca24_fa409_y4 = f_s_dadda_rca24_fa409_y1 | f_s_dadda_rca24_fa409_y3;
  assign f_s_dadda_rca24_fa410_f_s_dadda_rca24_fa409_y4 = f_s_dadda_rca24_fa409_y4;
  assign f_s_dadda_rca24_fa410_f_s_dadda_rca24_fa60_y2 = f_s_dadda_rca24_fa60_y2;
  assign f_s_dadda_rca24_fa410_f_s_dadda_rca24_ha13_y0 = f_s_dadda_rca24_ha13_y0;
  assign f_s_dadda_rca24_fa410_y0 = f_s_dadda_rca24_fa410_f_s_dadda_rca24_fa409_y4 ^ f_s_dadda_rca24_fa410_f_s_dadda_rca24_fa60_y2;
  assign f_s_dadda_rca24_fa410_y1 = f_s_dadda_rca24_fa410_f_s_dadda_rca24_fa409_y4 & f_s_dadda_rca24_fa410_f_s_dadda_rca24_fa60_y2;
  assign f_s_dadda_rca24_fa410_y2 = f_s_dadda_rca24_fa410_y0 ^ f_s_dadda_rca24_fa410_f_s_dadda_rca24_ha13_y0;
  assign f_s_dadda_rca24_fa410_y3 = f_s_dadda_rca24_fa410_y0 & f_s_dadda_rca24_fa410_f_s_dadda_rca24_ha13_y0;
  assign f_s_dadda_rca24_fa410_y4 = f_s_dadda_rca24_fa410_y1 | f_s_dadda_rca24_fa410_y3;
  assign f_s_dadda_rca24_fa411_f_s_dadda_rca24_fa410_y4 = f_s_dadda_rca24_fa410_y4;
  assign f_s_dadda_rca24_fa411_f_s_dadda_rca24_fa69_y2 = f_s_dadda_rca24_fa69_y2;
  assign f_s_dadda_rca24_fa411_f_s_dadda_rca24_ha14_y0 = f_s_dadda_rca24_ha14_y0;
  assign f_s_dadda_rca24_fa411_y0 = f_s_dadda_rca24_fa411_f_s_dadda_rca24_fa410_y4 ^ f_s_dadda_rca24_fa411_f_s_dadda_rca24_fa69_y2;
  assign f_s_dadda_rca24_fa411_y1 = f_s_dadda_rca24_fa411_f_s_dadda_rca24_fa410_y4 & f_s_dadda_rca24_fa411_f_s_dadda_rca24_fa69_y2;
  assign f_s_dadda_rca24_fa411_y2 = f_s_dadda_rca24_fa411_y0 ^ f_s_dadda_rca24_fa411_f_s_dadda_rca24_ha14_y0;
  assign f_s_dadda_rca24_fa411_y3 = f_s_dadda_rca24_fa411_y0 & f_s_dadda_rca24_fa411_f_s_dadda_rca24_ha14_y0;
  assign f_s_dadda_rca24_fa411_y4 = f_s_dadda_rca24_fa411_y1 | f_s_dadda_rca24_fa411_y3;
  assign f_s_dadda_rca24_fa412_f_s_dadda_rca24_fa411_y4 = f_s_dadda_rca24_fa411_y4;
  assign f_s_dadda_rca24_fa412_f_s_dadda_rca24_fa79_y2 = f_s_dadda_rca24_fa79_y2;
  assign f_s_dadda_rca24_fa412_f_s_dadda_rca24_ha15_y0 = f_s_dadda_rca24_ha15_y0;
  assign f_s_dadda_rca24_fa412_y0 = f_s_dadda_rca24_fa412_f_s_dadda_rca24_fa411_y4 ^ f_s_dadda_rca24_fa412_f_s_dadda_rca24_fa79_y2;
  assign f_s_dadda_rca24_fa412_y1 = f_s_dadda_rca24_fa412_f_s_dadda_rca24_fa411_y4 & f_s_dadda_rca24_fa412_f_s_dadda_rca24_fa79_y2;
  assign f_s_dadda_rca24_fa412_y2 = f_s_dadda_rca24_fa412_y0 ^ f_s_dadda_rca24_fa412_f_s_dadda_rca24_ha15_y0;
  assign f_s_dadda_rca24_fa412_y3 = f_s_dadda_rca24_fa412_y0 & f_s_dadda_rca24_fa412_f_s_dadda_rca24_ha15_y0;
  assign f_s_dadda_rca24_fa412_y4 = f_s_dadda_rca24_fa412_y1 | f_s_dadda_rca24_fa412_y3;
  assign f_s_dadda_rca24_fa413_f_s_dadda_rca24_fa412_y4 = f_s_dadda_rca24_fa412_y4;
  assign f_s_dadda_rca24_fa413_f_s_dadda_rca24_fa90_y2 = f_s_dadda_rca24_fa90_y2;
  assign f_s_dadda_rca24_fa413_f_s_dadda_rca24_ha16_y0 = f_s_dadda_rca24_ha16_y0;
  assign f_s_dadda_rca24_fa413_y0 = f_s_dadda_rca24_fa413_f_s_dadda_rca24_fa412_y4 ^ f_s_dadda_rca24_fa413_f_s_dadda_rca24_fa90_y2;
  assign f_s_dadda_rca24_fa413_y1 = f_s_dadda_rca24_fa413_f_s_dadda_rca24_fa412_y4 & f_s_dadda_rca24_fa413_f_s_dadda_rca24_fa90_y2;
  assign f_s_dadda_rca24_fa413_y2 = f_s_dadda_rca24_fa413_y0 ^ f_s_dadda_rca24_fa413_f_s_dadda_rca24_ha16_y0;
  assign f_s_dadda_rca24_fa413_y3 = f_s_dadda_rca24_fa413_y0 & f_s_dadda_rca24_fa413_f_s_dadda_rca24_ha16_y0;
  assign f_s_dadda_rca24_fa413_y4 = f_s_dadda_rca24_fa413_y1 | f_s_dadda_rca24_fa413_y3;
  assign f_s_dadda_rca24_fa414_f_s_dadda_rca24_fa413_y4 = f_s_dadda_rca24_fa413_y4;
  assign f_s_dadda_rca24_fa414_f_s_dadda_rca24_fa102_y2 = f_s_dadda_rca24_fa102_y2;
  assign f_s_dadda_rca24_fa414_f_s_dadda_rca24_ha17_y0 = f_s_dadda_rca24_ha17_y0;
  assign f_s_dadda_rca24_fa414_y0 = f_s_dadda_rca24_fa414_f_s_dadda_rca24_fa413_y4 ^ f_s_dadda_rca24_fa414_f_s_dadda_rca24_fa102_y2;
  assign f_s_dadda_rca24_fa414_y1 = f_s_dadda_rca24_fa414_f_s_dadda_rca24_fa413_y4 & f_s_dadda_rca24_fa414_f_s_dadda_rca24_fa102_y2;
  assign f_s_dadda_rca24_fa414_y2 = f_s_dadda_rca24_fa414_y0 ^ f_s_dadda_rca24_fa414_f_s_dadda_rca24_ha17_y0;
  assign f_s_dadda_rca24_fa414_y3 = f_s_dadda_rca24_fa414_y0 & f_s_dadda_rca24_fa414_f_s_dadda_rca24_ha17_y0;
  assign f_s_dadda_rca24_fa414_y4 = f_s_dadda_rca24_fa414_y1 | f_s_dadda_rca24_fa414_y3;
  assign f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa414_y4 = f_s_dadda_rca24_fa414_y4;
  assign f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa114_y2 = f_s_dadda_rca24_fa114_y2;
  assign f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa115_y2 = f_s_dadda_rca24_fa115_y2;
  assign f_s_dadda_rca24_fa415_y0 = f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa414_y4 ^ f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa114_y2;
  assign f_s_dadda_rca24_fa415_y1 = f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa414_y4 & f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa114_y2;
  assign f_s_dadda_rca24_fa415_y2 = f_s_dadda_rca24_fa415_y0 ^ f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa115_y2;
  assign f_s_dadda_rca24_fa415_y3 = f_s_dadda_rca24_fa415_y0 & f_s_dadda_rca24_fa415_f_s_dadda_rca24_fa115_y2;
  assign f_s_dadda_rca24_fa415_y4 = f_s_dadda_rca24_fa415_y1 | f_s_dadda_rca24_fa415_y3;
  assign f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa415_y4 = f_s_dadda_rca24_fa415_y4;
  assign f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa127_y2 = f_s_dadda_rca24_fa127_y2;
  assign f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa128_y2 = f_s_dadda_rca24_fa128_y2;
  assign f_s_dadda_rca24_fa416_y0 = f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa415_y4 ^ f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa127_y2;
  assign f_s_dadda_rca24_fa416_y1 = f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa415_y4 & f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa127_y2;
  assign f_s_dadda_rca24_fa416_y2 = f_s_dadda_rca24_fa416_y0 ^ f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa128_y2;
  assign f_s_dadda_rca24_fa416_y3 = f_s_dadda_rca24_fa416_y0 & f_s_dadda_rca24_fa416_f_s_dadda_rca24_fa128_y2;
  assign f_s_dadda_rca24_fa416_y4 = f_s_dadda_rca24_fa416_y1 | f_s_dadda_rca24_fa416_y3;
  assign f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa416_y4 = f_s_dadda_rca24_fa416_y4;
  assign f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa140_y2 = f_s_dadda_rca24_fa140_y2;
  assign f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa141_y2 = f_s_dadda_rca24_fa141_y2;
  assign f_s_dadda_rca24_fa417_y0 = f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa416_y4 ^ f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa140_y2;
  assign f_s_dadda_rca24_fa417_y1 = f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa416_y4 & f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa140_y2;
  assign f_s_dadda_rca24_fa417_y2 = f_s_dadda_rca24_fa417_y0 ^ f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa141_y2;
  assign f_s_dadda_rca24_fa417_y3 = f_s_dadda_rca24_fa417_y0 & f_s_dadda_rca24_fa417_f_s_dadda_rca24_fa141_y2;
  assign f_s_dadda_rca24_fa417_y4 = f_s_dadda_rca24_fa417_y1 | f_s_dadda_rca24_fa417_y3;
  assign f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa417_y4 = f_s_dadda_rca24_fa417_y4;
  assign f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa153_y2 = f_s_dadda_rca24_fa153_y2;
  assign f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa154_y2 = f_s_dadda_rca24_fa154_y2;
  assign f_s_dadda_rca24_fa418_y0 = f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa417_y4 ^ f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa153_y2;
  assign f_s_dadda_rca24_fa418_y1 = f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa417_y4 & f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa153_y2;
  assign f_s_dadda_rca24_fa418_y2 = f_s_dadda_rca24_fa418_y0 ^ f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa154_y2;
  assign f_s_dadda_rca24_fa418_y3 = f_s_dadda_rca24_fa418_y0 & f_s_dadda_rca24_fa418_f_s_dadda_rca24_fa154_y2;
  assign f_s_dadda_rca24_fa418_y4 = f_s_dadda_rca24_fa418_y1 | f_s_dadda_rca24_fa418_y3;
  assign f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa418_y4 = f_s_dadda_rca24_fa418_y4;
  assign f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa166_y2 = f_s_dadda_rca24_fa166_y2;
  assign f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa167_y2 = f_s_dadda_rca24_fa167_y2;
  assign f_s_dadda_rca24_fa419_y0 = f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa418_y4 ^ f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa166_y2;
  assign f_s_dadda_rca24_fa419_y1 = f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa418_y4 & f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa166_y2;
  assign f_s_dadda_rca24_fa419_y2 = f_s_dadda_rca24_fa419_y0 ^ f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa167_y2;
  assign f_s_dadda_rca24_fa419_y3 = f_s_dadda_rca24_fa419_y0 & f_s_dadda_rca24_fa419_f_s_dadda_rca24_fa167_y2;
  assign f_s_dadda_rca24_fa419_y4 = f_s_dadda_rca24_fa419_y1 | f_s_dadda_rca24_fa419_y3;
  assign f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa419_y4 = f_s_dadda_rca24_fa419_y4;
  assign f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa179_y2 = f_s_dadda_rca24_fa179_y2;
  assign f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa180_y2 = f_s_dadda_rca24_fa180_y2;
  assign f_s_dadda_rca24_fa420_y0 = f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa419_y4 ^ f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa179_y2;
  assign f_s_dadda_rca24_fa420_y1 = f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa419_y4 & f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa179_y2;
  assign f_s_dadda_rca24_fa420_y2 = f_s_dadda_rca24_fa420_y0 ^ f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa180_y2;
  assign f_s_dadda_rca24_fa420_y3 = f_s_dadda_rca24_fa420_y0 & f_s_dadda_rca24_fa420_f_s_dadda_rca24_fa180_y2;
  assign f_s_dadda_rca24_fa420_y4 = f_s_dadda_rca24_fa420_y1 | f_s_dadda_rca24_fa420_y3;
  assign f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa420_y4 = f_s_dadda_rca24_fa420_y4;
  assign f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa192_y2 = f_s_dadda_rca24_fa192_y2;
  assign f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa193_y2 = f_s_dadda_rca24_fa193_y2;
  assign f_s_dadda_rca24_fa421_y0 = f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa420_y4 ^ f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa192_y2;
  assign f_s_dadda_rca24_fa421_y1 = f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa420_y4 & f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa192_y2;
  assign f_s_dadda_rca24_fa421_y2 = f_s_dadda_rca24_fa421_y0 ^ f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa193_y2;
  assign f_s_dadda_rca24_fa421_y3 = f_s_dadda_rca24_fa421_y0 & f_s_dadda_rca24_fa421_f_s_dadda_rca24_fa193_y2;
  assign f_s_dadda_rca24_fa421_y4 = f_s_dadda_rca24_fa421_y1 | f_s_dadda_rca24_fa421_y3;
  assign f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa421_y4 = f_s_dadda_rca24_fa421_y4;
  assign f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa205_y2 = f_s_dadda_rca24_fa205_y2;
  assign f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa206_y2 = f_s_dadda_rca24_fa206_y2;
  assign f_s_dadda_rca24_fa422_y0 = f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa421_y4 ^ f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa205_y2;
  assign f_s_dadda_rca24_fa422_y1 = f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa421_y4 & f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa205_y2;
  assign f_s_dadda_rca24_fa422_y2 = f_s_dadda_rca24_fa422_y0 ^ f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa206_y2;
  assign f_s_dadda_rca24_fa422_y3 = f_s_dadda_rca24_fa422_y0 & f_s_dadda_rca24_fa422_f_s_dadda_rca24_fa206_y2;
  assign f_s_dadda_rca24_fa422_y4 = f_s_dadda_rca24_fa422_y1 | f_s_dadda_rca24_fa422_y3;
  assign f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa422_y4 = f_s_dadda_rca24_fa422_y4;
  assign f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa218_y2 = f_s_dadda_rca24_fa218_y2;
  assign f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa219_y2 = f_s_dadda_rca24_fa219_y2;
  assign f_s_dadda_rca24_fa423_y0 = f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa422_y4 ^ f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa218_y2;
  assign f_s_dadda_rca24_fa423_y1 = f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa422_y4 & f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa218_y2;
  assign f_s_dadda_rca24_fa423_y2 = f_s_dadda_rca24_fa423_y0 ^ f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa219_y2;
  assign f_s_dadda_rca24_fa423_y3 = f_s_dadda_rca24_fa423_y0 & f_s_dadda_rca24_fa423_f_s_dadda_rca24_fa219_y2;
  assign f_s_dadda_rca24_fa423_y4 = f_s_dadda_rca24_fa423_y1 | f_s_dadda_rca24_fa423_y3;
  assign f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa423_y4 = f_s_dadda_rca24_fa423_y4;
  assign f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa231_y2 = f_s_dadda_rca24_fa231_y2;
  assign f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa232_y2 = f_s_dadda_rca24_fa232_y2;
  assign f_s_dadda_rca24_fa424_y0 = f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa423_y4 ^ f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa231_y2;
  assign f_s_dadda_rca24_fa424_y1 = f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa423_y4 & f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa231_y2;
  assign f_s_dadda_rca24_fa424_y2 = f_s_dadda_rca24_fa424_y0 ^ f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa232_y2;
  assign f_s_dadda_rca24_fa424_y3 = f_s_dadda_rca24_fa424_y0 & f_s_dadda_rca24_fa424_f_s_dadda_rca24_fa232_y2;
  assign f_s_dadda_rca24_fa424_y4 = f_s_dadda_rca24_fa424_y1 | f_s_dadda_rca24_fa424_y3;
  assign f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa424_y4 = f_s_dadda_rca24_fa424_y4;
  assign f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa244_y2 = f_s_dadda_rca24_fa244_y2;
  assign f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa245_y2 = f_s_dadda_rca24_fa245_y2;
  assign f_s_dadda_rca24_fa425_y0 = f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa424_y4 ^ f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa244_y2;
  assign f_s_dadda_rca24_fa425_y1 = f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa424_y4 & f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa244_y2;
  assign f_s_dadda_rca24_fa425_y2 = f_s_dadda_rca24_fa425_y0 ^ f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa245_y2;
  assign f_s_dadda_rca24_fa425_y3 = f_s_dadda_rca24_fa425_y0 & f_s_dadda_rca24_fa425_f_s_dadda_rca24_fa245_y2;
  assign f_s_dadda_rca24_fa425_y4 = f_s_dadda_rca24_fa425_y1 | f_s_dadda_rca24_fa425_y3;
  assign f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa425_y4 = f_s_dadda_rca24_fa425_y4;
  assign f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa256_y2 = f_s_dadda_rca24_fa256_y2;
  assign f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa257_y2 = f_s_dadda_rca24_fa257_y2;
  assign f_s_dadda_rca24_fa426_y0 = f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa425_y4 ^ f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa256_y2;
  assign f_s_dadda_rca24_fa426_y1 = f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa425_y4 & f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa256_y2;
  assign f_s_dadda_rca24_fa426_y2 = f_s_dadda_rca24_fa426_y0 ^ f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa257_y2;
  assign f_s_dadda_rca24_fa426_y3 = f_s_dadda_rca24_fa426_y0 & f_s_dadda_rca24_fa426_f_s_dadda_rca24_fa257_y2;
  assign f_s_dadda_rca24_fa426_y4 = f_s_dadda_rca24_fa426_y1 | f_s_dadda_rca24_fa426_y3;
  assign f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa426_y4 = f_s_dadda_rca24_fa426_y4;
  assign f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa267_y2 = f_s_dadda_rca24_fa267_y2;
  assign f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa268_y2 = f_s_dadda_rca24_fa268_y2;
  assign f_s_dadda_rca24_fa427_y0 = f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa426_y4 ^ f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa267_y2;
  assign f_s_dadda_rca24_fa427_y1 = f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa426_y4 & f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa267_y2;
  assign f_s_dadda_rca24_fa427_y2 = f_s_dadda_rca24_fa427_y0 ^ f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa268_y2;
  assign f_s_dadda_rca24_fa427_y3 = f_s_dadda_rca24_fa427_y0 & f_s_dadda_rca24_fa427_f_s_dadda_rca24_fa268_y2;
  assign f_s_dadda_rca24_fa427_y4 = f_s_dadda_rca24_fa427_y1 | f_s_dadda_rca24_fa427_y3;
  assign f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa427_y4 = f_s_dadda_rca24_fa427_y4;
  assign f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa277_y2 = f_s_dadda_rca24_fa277_y2;
  assign f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa278_y2 = f_s_dadda_rca24_fa278_y2;
  assign f_s_dadda_rca24_fa428_y0 = f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa427_y4 ^ f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa277_y2;
  assign f_s_dadda_rca24_fa428_y1 = f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa427_y4 & f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa277_y2;
  assign f_s_dadda_rca24_fa428_y2 = f_s_dadda_rca24_fa428_y0 ^ f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa278_y2;
  assign f_s_dadda_rca24_fa428_y3 = f_s_dadda_rca24_fa428_y0 & f_s_dadda_rca24_fa428_f_s_dadda_rca24_fa278_y2;
  assign f_s_dadda_rca24_fa428_y4 = f_s_dadda_rca24_fa428_y1 | f_s_dadda_rca24_fa428_y3;
  assign f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa428_y4 = f_s_dadda_rca24_fa428_y4;
  assign f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa286_y2 = f_s_dadda_rca24_fa286_y2;
  assign f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa287_y2 = f_s_dadda_rca24_fa287_y2;
  assign f_s_dadda_rca24_fa429_y0 = f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa428_y4 ^ f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa286_y2;
  assign f_s_dadda_rca24_fa429_y1 = f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa428_y4 & f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa286_y2;
  assign f_s_dadda_rca24_fa429_y2 = f_s_dadda_rca24_fa429_y0 ^ f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa287_y2;
  assign f_s_dadda_rca24_fa429_y3 = f_s_dadda_rca24_fa429_y0 & f_s_dadda_rca24_fa429_f_s_dadda_rca24_fa287_y2;
  assign f_s_dadda_rca24_fa429_y4 = f_s_dadda_rca24_fa429_y1 | f_s_dadda_rca24_fa429_y3;
  assign f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa429_y4 = f_s_dadda_rca24_fa429_y4;
  assign f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa294_y2 = f_s_dadda_rca24_fa294_y2;
  assign f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa295_y2 = f_s_dadda_rca24_fa295_y2;
  assign f_s_dadda_rca24_fa430_y0 = f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa429_y4 ^ f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa294_y2;
  assign f_s_dadda_rca24_fa430_y1 = f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa429_y4 & f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa294_y2;
  assign f_s_dadda_rca24_fa430_y2 = f_s_dadda_rca24_fa430_y0 ^ f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa295_y2;
  assign f_s_dadda_rca24_fa430_y3 = f_s_dadda_rca24_fa430_y0 & f_s_dadda_rca24_fa430_f_s_dadda_rca24_fa295_y2;
  assign f_s_dadda_rca24_fa430_y4 = f_s_dadda_rca24_fa430_y1 | f_s_dadda_rca24_fa430_y3;
  assign f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa430_y4 = f_s_dadda_rca24_fa430_y4;
  assign f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa301_y2 = f_s_dadda_rca24_fa301_y2;
  assign f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa302_y2 = f_s_dadda_rca24_fa302_y2;
  assign f_s_dadda_rca24_fa431_y0 = f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa430_y4 ^ f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa301_y2;
  assign f_s_dadda_rca24_fa431_y1 = f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa430_y4 & f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa301_y2;
  assign f_s_dadda_rca24_fa431_y2 = f_s_dadda_rca24_fa431_y0 ^ f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa302_y2;
  assign f_s_dadda_rca24_fa431_y3 = f_s_dadda_rca24_fa431_y0 & f_s_dadda_rca24_fa431_f_s_dadda_rca24_fa302_y2;
  assign f_s_dadda_rca24_fa431_y4 = f_s_dadda_rca24_fa431_y1 | f_s_dadda_rca24_fa431_y3;
  assign f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa431_y4 = f_s_dadda_rca24_fa431_y4;
  assign f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa307_y2 = f_s_dadda_rca24_fa307_y2;
  assign f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa308_y2 = f_s_dadda_rca24_fa308_y2;
  assign f_s_dadda_rca24_fa432_y0 = f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa431_y4 ^ f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa307_y2;
  assign f_s_dadda_rca24_fa432_y1 = f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa431_y4 & f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa307_y2;
  assign f_s_dadda_rca24_fa432_y2 = f_s_dadda_rca24_fa432_y0 ^ f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa308_y2;
  assign f_s_dadda_rca24_fa432_y3 = f_s_dadda_rca24_fa432_y0 & f_s_dadda_rca24_fa432_f_s_dadda_rca24_fa308_y2;
  assign f_s_dadda_rca24_fa432_y4 = f_s_dadda_rca24_fa432_y1 | f_s_dadda_rca24_fa432_y3;
  assign f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa432_y4 = f_s_dadda_rca24_fa432_y4;
  assign f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa312_y2 = f_s_dadda_rca24_fa312_y2;
  assign f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa313_y2 = f_s_dadda_rca24_fa313_y2;
  assign f_s_dadda_rca24_fa433_y0 = f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa432_y4 ^ f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa312_y2;
  assign f_s_dadda_rca24_fa433_y1 = f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa432_y4 & f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa312_y2;
  assign f_s_dadda_rca24_fa433_y2 = f_s_dadda_rca24_fa433_y0 ^ f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa313_y2;
  assign f_s_dadda_rca24_fa433_y3 = f_s_dadda_rca24_fa433_y0 & f_s_dadda_rca24_fa433_f_s_dadda_rca24_fa313_y2;
  assign f_s_dadda_rca24_fa433_y4 = f_s_dadda_rca24_fa433_y1 | f_s_dadda_rca24_fa433_y3;
  assign f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa433_y4 = f_s_dadda_rca24_fa433_y4;
  assign f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa316_y2 = f_s_dadda_rca24_fa316_y2;
  assign f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa317_y2 = f_s_dadda_rca24_fa317_y2;
  assign f_s_dadda_rca24_fa434_y0 = f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa433_y4 ^ f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa316_y2;
  assign f_s_dadda_rca24_fa434_y1 = f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa433_y4 & f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa316_y2;
  assign f_s_dadda_rca24_fa434_y2 = f_s_dadda_rca24_fa434_y0 ^ f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa317_y2;
  assign f_s_dadda_rca24_fa434_y3 = f_s_dadda_rca24_fa434_y0 & f_s_dadda_rca24_fa434_f_s_dadda_rca24_fa317_y2;
  assign f_s_dadda_rca24_fa434_y4 = f_s_dadda_rca24_fa434_y1 | f_s_dadda_rca24_fa434_y3;
  assign f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa434_y4 = f_s_dadda_rca24_fa434_y4;
  assign f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa319_y2 = f_s_dadda_rca24_fa319_y2;
  assign f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa320_y2 = f_s_dadda_rca24_fa320_y2;
  assign f_s_dadda_rca24_fa435_y0 = f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa434_y4 ^ f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa319_y2;
  assign f_s_dadda_rca24_fa435_y1 = f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa434_y4 & f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa319_y2;
  assign f_s_dadda_rca24_fa435_y2 = f_s_dadda_rca24_fa435_y0 ^ f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa320_y2;
  assign f_s_dadda_rca24_fa435_y3 = f_s_dadda_rca24_fa435_y0 & f_s_dadda_rca24_fa435_f_s_dadda_rca24_fa320_y2;
  assign f_s_dadda_rca24_fa435_y4 = f_s_dadda_rca24_fa435_y1 | f_s_dadda_rca24_fa435_y3;
  assign f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa435_y4 = f_s_dadda_rca24_fa435_y4;
  assign f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa321_y2 = f_s_dadda_rca24_fa321_y2;
  assign f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa322_y2 = f_s_dadda_rca24_fa322_y2;
  assign f_s_dadda_rca24_fa436_y0 = f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa435_y4 ^ f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa321_y2;
  assign f_s_dadda_rca24_fa436_y1 = f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa435_y4 & f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa321_y2;
  assign f_s_dadda_rca24_fa436_y2 = f_s_dadda_rca24_fa436_y0 ^ f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa322_y2;
  assign f_s_dadda_rca24_fa436_y3 = f_s_dadda_rca24_fa436_y0 & f_s_dadda_rca24_fa436_f_s_dadda_rca24_fa322_y2;
  assign f_s_dadda_rca24_fa436_y4 = f_s_dadda_rca24_fa436_y1 | f_s_dadda_rca24_fa436_y3;
  assign f_s_dadda_rca24_nand_18_23_a_18 = a_18;
  assign f_s_dadda_rca24_nand_18_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_18_23_y0 = ~(f_s_dadda_rca24_nand_18_23_a_18 & f_s_dadda_rca24_nand_18_23_b_23);
  assign f_s_dadda_rca24_fa437_f_s_dadda_rca24_fa436_y4 = f_s_dadda_rca24_fa436_y4;
  assign f_s_dadda_rca24_fa437_f_s_dadda_rca24_nand_18_23_y0 = f_s_dadda_rca24_nand_18_23_y0;
  assign f_s_dadda_rca24_fa437_f_s_dadda_rca24_fa323_y2 = f_s_dadda_rca24_fa323_y2;
  assign f_s_dadda_rca24_fa437_y0 = f_s_dadda_rca24_fa437_f_s_dadda_rca24_fa436_y4 ^ f_s_dadda_rca24_fa437_f_s_dadda_rca24_nand_18_23_y0;
  assign f_s_dadda_rca24_fa437_y1 = f_s_dadda_rca24_fa437_f_s_dadda_rca24_fa436_y4 & f_s_dadda_rca24_fa437_f_s_dadda_rca24_nand_18_23_y0;
  assign f_s_dadda_rca24_fa437_y2 = f_s_dadda_rca24_fa437_y0 ^ f_s_dadda_rca24_fa437_f_s_dadda_rca24_fa323_y2;
  assign f_s_dadda_rca24_fa437_y3 = f_s_dadda_rca24_fa437_y0 & f_s_dadda_rca24_fa437_f_s_dadda_rca24_fa323_y2;
  assign f_s_dadda_rca24_fa437_y4 = f_s_dadda_rca24_fa437_y1 | f_s_dadda_rca24_fa437_y3;
  assign f_s_dadda_rca24_and_20_22_a_20 = a_20;
  assign f_s_dadda_rca24_and_20_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_20_22_y0 = f_s_dadda_rca24_and_20_22_a_20 & f_s_dadda_rca24_and_20_22_b_22;
  assign f_s_dadda_rca24_nand_19_23_a_19 = a_19;
  assign f_s_dadda_rca24_nand_19_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_19_23_y0 = ~(f_s_dadda_rca24_nand_19_23_a_19 & f_s_dadda_rca24_nand_19_23_b_23);
  assign f_s_dadda_rca24_fa438_f_s_dadda_rca24_fa437_y4 = f_s_dadda_rca24_fa437_y4;
  assign f_s_dadda_rca24_fa438_f_s_dadda_rca24_and_20_22_y0 = f_s_dadda_rca24_and_20_22_y0;
  assign f_s_dadda_rca24_fa438_f_s_dadda_rca24_nand_19_23_y0 = f_s_dadda_rca24_nand_19_23_y0;
  assign f_s_dadda_rca24_fa438_y0 = f_s_dadda_rca24_fa438_f_s_dadda_rca24_fa437_y4 ^ f_s_dadda_rca24_fa438_f_s_dadda_rca24_and_20_22_y0;
  assign f_s_dadda_rca24_fa438_y1 = f_s_dadda_rca24_fa438_f_s_dadda_rca24_fa437_y4 & f_s_dadda_rca24_fa438_f_s_dadda_rca24_and_20_22_y0;
  assign f_s_dadda_rca24_fa438_y2 = f_s_dadda_rca24_fa438_y0 ^ f_s_dadda_rca24_fa438_f_s_dadda_rca24_nand_19_23_y0;
  assign f_s_dadda_rca24_fa438_y3 = f_s_dadda_rca24_fa438_y0 & f_s_dadda_rca24_fa438_f_s_dadda_rca24_nand_19_23_y0;
  assign f_s_dadda_rca24_fa438_y4 = f_s_dadda_rca24_fa438_y1 | f_s_dadda_rca24_fa438_y3;
  assign f_s_dadda_rca24_and_22_21_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_21_b_21 = b_21;
  assign f_s_dadda_rca24_and_22_21_y0 = f_s_dadda_rca24_and_22_21_a_22 & f_s_dadda_rca24_and_22_21_b_21;
  assign f_s_dadda_rca24_and_21_22_a_21 = a_21;
  assign f_s_dadda_rca24_and_21_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_21_22_y0 = f_s_dadda_rca24_and_21_22_a_21 & f_s_dadda_rca24_and_21_22_b_22;
  assign f_s_dadda_rca24_fa439_f_s_dadda_rca24_fa438_y4 = f_s_dadda_rca24_fa438_y4;
  assign f_s_dadda_rca24_fa439_f_s_dadda_rca24_and_22_21_y0 = f_s_dadda_rca24_and_22_21_y0;
  assign f_s_dadda_rca24_fa439_f_s_dadda_rca24_and_21_22_y0 = f_s_dadda_rca24_and_21_22_y0;
  assign f_s_dadda_rca24_fa439_y0 = f_s_dadda_rca24_fa439_f_s_dadda_rca24_fa438_y4 ^ f_s_dadda_rca24_fa439_f_s_dadda_rca24_and_22_21_y0;
  assign f_s_dadda_rca24_fa439_y1 = f_s_dadda_rca24_fa439_f_s_dadda_rca24_fa438_y4 & f_s_dadda_rca24_fa439_f_s_dadda_rca24_and_22_21_y0;
  assign f_s_dadda_rca24_fa439_y2 = f_s_dadda_rca24_fa439_y0 ^ f_s_dadda_rca24_fa439_f_s_dadda_rca24_and_21_22_y0;
  assign f_s_dadda_rca24_fa439_y3 = f_s_dadda_rca24_fa439_y0 & f_s_dadda_rca24_fa439_f_s_dadda_rca24_and_21_22_y0;
  assign f_s_dadda_rca24_fa439_y4 = f_s_dadda_rca24_fa439_y1 | f_s_dadda_rca24_fa439_y3;
  assign f_s_dadda_rca24_nand_23_21_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_21_b_21 = b_21;
  assign f_s_dadda_rca24_nand_23_21_y0 = ~(f_s_dadda_rca24_nand_23_21_a_23 & f_s_dadda_rca24_nand_23_21_b_21);
  assign f_s_dadda_rca24_fa440_f_s_dadda_rca24_fa439_y4 = f_s_dadda_rca24_fa439_y4;
  assign f_s_dadda_rca24_fa440_f_s_dadda_rca24_fa399_y4 = f_s_dadda_rca24_fa399_y4;
  assign f_s_dadda_rca24_fa440_f_s_dadda_rca24_nand_23_21_y0 = f_s_dadda_rca24_nand_23_21_y0;
  assign f_s_dadda_rca24_fa440_y0 = f_s_dadda_rca24_fa440_f_s_dadda_rca24_fa439_y4 ^ f_s_dadda_rca24_fa440_f_s_dadda_rca24_fa399_y4;
  assign f_s_dadda_rca24_fa440_y1 = f_s_dadda_rca24_fa440_f_s_dadda_rca24_fa439_y4 & f_s_dadda_rca24_fa440_f_s_dadda_rca24_fa399_y4;
  assign f_s_dadda_rca24_fa440_y2 = f_s_dadda_rca24_fa440_y0 ^ f_s_dadda_rca24_fa440_f_s_dadda_rca24_nand_23_21_y0;
  assign f_s_dadda_rca24_fa440_y3 = f_s_dadda_rca24_fa440_y0 & f_s_dadda_rca24_fa440_f_s_dadda_rca24_nand_23_21_y0;
  assign f_s_dadda_rca24_fa440_y4 = f_s_dadda_rca24_fa440_y1 | f_s_dadda_rca24_fa440_y3;
  assign f_s_dadda_rca24_and_2_0_a_2 = a_2;
  assign f_s_dadda_rca24_and_2_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_2_0_y0 = f_s_dadda_rca24_and_2_0_a_2 & f_s_dadda_rca24_and_2_0_b_0;
  assign f_s_dadda_rca24_and_1_1_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_1_1_y0 = f_s_dadda_rca24_and_1_1_a_1 & f_s_dadda_rca24_and_1_1_b_1;
  assign f_s_dadda_rca24_ha21_f_s_dadda_rca24_and_2_0_y0 = f_s_dadda_rca24_and_2_0_y0;
  assign f_s_dadda_rca24_ha21_f_s_dadda_rca24_and_1_1_y0 = f_s_dadda_rca24_and_1_1_y0;
  assign f_s_dadda_rca24_ha21_y0 = f_s_dadda_rca24_ha21_f_s_dadda_rca24_and_2_0_y0 ^ f_s_dadda_rca24_ha21_f_s_dadda_rca24_and_1_1_y0;
  assign f_s_dadda_rca24_ha21_y1 = f_s_dadda_rca24_ha21_f_s_dadda_rca24_and_2_0_y0 & f_s_dadda_rca24_ha21_f_s_dadda_rca24_and_1_1_y0;
  assign f_s_dadda_rca24_and_1_2_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_1_2_y0 = f_s_dadda_rca24_and_1_2_a_1 & f_s_dadda_rca24_and_1_2_b_2;
  assign f_s_dadda_rca24_and_0_3_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_3_b_3 = b_3;
  assign f_s_dadda_rca24_and_0_3_y0 = f_s_dadda_rca24_and_0_3_a_0 & f_s_dadda_rca24_and_0_3_b_3;
  assign f_s_dadda_rca24_fa441_f_s_dadda_rca24_ha21_y1 = f_s_dadda_rca24_ha21_y1;
  assign f_s_dadda_rca24_fa441_f_s_dadda_rca24_and_1_2_y0 = f_s_dadda_rca24_and_1_2_y0;
  assign f_s_dadda_rca24_fa441_f_s_dadda_rca24_and_0_3_y0 = f_s_dadda_rca24_and_0_3_y0;
  assign f_s_dadda_rca24_fa441_y0 = f_s_dadda_rca24_fa441_f_s_dadda_rca24_ha21_y1 ^ f_s_dadda_rca24_fa441_f_s_dadda_rca24_and_1_2_y0;
  assign f_s_dadda_rca24_fa441_y1 = f_s_dadda_rca24_fa441_f_s_dadda_rca24_ha21_y1 & f_s_dadda_rca24_fa441_f_s_dadda_rca24_and_1_2_y0;
  assign f_s_dadda_rca24_fa441_y2 = f_s_dadda_rca24_fa441_y0 ^ f_s_dadda_rca24_fa441_f_s_dadda_rca24_and_0_3_y0;
  assign f_s_dadda_rca24_fa441_y3 = f_s_dadda_rca24_fa441_y0 & f_s_dadda_rca24_fa441_f_s_dadda_rca24_and_0_3_y0;
  assign f_s_dadda_rca24_fa441_y4 = f_s_dadda_rca24_fa441_y1 | f_s_dadda_rca24_fa441_y3;
  assign f_s_dadda_rca24_and_0_4_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_4_b_4 = b_4;
  assign f_s_dadda_rca24_and_0_4_y0 = f_s_dadda_rca24_and_0_4_a_0 & f_s_dadda_rca24_and_0_4_b_4;
  assign f_s_dadda_rca24_fa442_f_s_dadda_rca24_fa441_y4 = f_s_dadda_rca24_fa441_y4;
  assign f_s_dadda_rca24_fa442_f_s_dadda_rca24_and_0_4_y0 = f_s_dadda_rca24_and_0_4_y0;
  assign f_s_dadda_rca24_fa442_f_s_dadda_rca24_ha18_y0 = f_s_dadda_rca24_ha18_y0;
  assign f_s_dadda_rca24_fa442_y0 = f_s_dadda_rca24_fa442_f_s_dadda_rca24_fa441_y4 ^ f_s_dadda_rca24_fa442_f_s_dadda_rca24_and_0_4_y0;
  assign f_s_dadda_rca24_fa442_y1 = f_s_dadda_rca24_fa442_f_s_dadda_rca24_fa441_y4 & f_s_dadda_rca24_fa442_f_s_dadda_rca24_and_0_4_y0;
  assign f_s_dadda_rca24_fa442_y2 = f_s_dadda_rca24_fa442_y0 ^ f_s_dadda_rca24_fa442_f_s_dadda_rca24_ha18_y0;
  assign f_s_dadda_rca24_fa442_y3 = f_s_dadda_rca24_fa442_y0 & f_s_dadda_rca24_fa442_f_s_dadda_rca24_ha18_y0;
  assign f_s_dadda_rca24_fa442_y4 = f_s_dadda_rca24_fa442_y1 | f_s_dadda_rca24_fa442_y3;
  assign f_s_dadda_rca24_fa443_f_s_dadda_rca24_fa442_y4 = f_s_dadda_rca24_fa442_y4;
  assign f_s_dadda_rca24_fa443_f_s_dadda_rca24_fa324_y2 = f_s_dadda_rca24_fa324_y2;
  assign f_s_dadda_rca24_fa443_f_s_dadda_rca24_ha19_y0 = f_s_dadda_rca24_ha19_y0;
  assign f_s_dadda_rca24_fa443_y0 = f_s_dadda_rca24_fa443_f_s_dadda_rca24_fa442_y4 ^ f_s_dadda_rca24_fa443_f_s_dadda_rca24_fa324_y2;
  assign f_s_dadda_rca24_fa443_y1 = f_s_dadda_rca24_fa443_f_s_dadda_rca24_fa442_y4 & f_s_dadda_rca24_fa443_f_s_dadda_rca24_fa324_y2;
  assign f_s_dadda_rca24_fa443_y2 = f_s_dadda_rca24_fa443_y0 ^ f_s_dadda_rca24_fa443_f_s_dadda_rca24_ha19_y0;
  assign f_s_dadda_rca24_fa443_y3 = f_s_dadda_rca24_fa443_y0 & f_s_dadda_rca24_fa443_f_s_dadda_rca24_ha19_y0;
  assign f_s_dadda_rca24_fa443_y4 = f_s_dadda_rca24_fa443_y1 | f_s_dadda_rca24_fa443_y3;
  assign f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa443_y4 = f_s_dadda_rca24_fa443_y4;
  assign f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa325_y2 = f_s_dadda_rca24_fa325_y2;
  assign f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa326_y2 = f_s_dadda_rca24_fa326_y2;
  assign f_s_dadda_rca24_fa444_y0 = f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa443_y4 ^ f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa325_y2;
  assign f_s_dadda_rca24_fa444_y1 = f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa443_y4 & f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa325_y2;
  assign f_s_dadda_rca24_fa444_y2 = f_s_dadda_rca24_fa444_y0 ^ f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa326_y2;
  assign f_s_dadda_rca24_fa444_y3 = f_s_dadda_rca24_fa444_y0 & f_s_dadda_rca24_fa444_f_s_dadda_rca24_fa326_y2;
  assign f_s_dadda_rca24_fa444_y4 = f_s_dadda_rca24_fa444_y1 | f_s_dadda_rca24_fa444_y3;
  assign f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa444_y4 = f_s_dadda_rca24_fa444_y4;
  assign f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa327_y2 = f_s_dadda_rca24_fa327_y2;
  assign f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa328_y2 = f_s_dadda_rca24_fa328_y2;
  assign f_s_dadda_rca24_fa445_y0 = f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa444_y4 ^ f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa327_y2;
  assign f_s_dadda_rca24_fa445_y1 = f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa444_y4 & f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa327_y2;
  assign f_s_dadda_rca24_fa445_y2 = f_s_dadda_rca24_fa445_y0 ^ f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa328_y2;
  assign f_s_dadda_rca24_fa445_y3 = f_s_dadda_rca24_fa445_y0 & f_s_dadda_rca24_fa445_f_s_dadda_rca24_fa328_y2;
  assign f_s_dadda_rca24_fa445_y4 = f_s_dadda_rca24_fa445_y1 | f_s_dadda_rca24_fa445_y3;
  assign f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa445_y4 = f_s_dadda_rca24_fa445_y4;
  assign f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa329_y2 = f_s_dadda_rca24_fa329_y2;
  assign f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa330_y2 = f_s_dadda_rca24_fa330_y2;
  assign f_s_dadda_rca24_fa446_y0 = f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa445_y4 ^ f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa329_y2;
  assign f_s_dadda_rca24_fa446_y1 = f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa445_y4 & f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa329_y2;
  assign f_s_dadda_rca24_fa446_y2 = f_s_dadda_rca24_fa446_y0 ^ f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa330_y2;
  assign f_s_dadda_rca24_fa446_y3 = f_s_dadda_rca24_fa446_y0 & f_s_dadda_rca24_fa446_f_s_dadda_rca24_fa330_y2;
  assign f_s_dadda_rca24_fa446_y4 = f_s_dadda_rca24_fa446_y1 | f_s_dadda_rca24_fa446_y3;
  assign f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa446_y4 = f_s_dadda_rca24_fa446_y4;
  assign f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa331_y2 = f_s_dadda_rca24_fa331_y2;
  assign f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa332_y2 = f_s_dadda_rca24_fa332_y2;
  assign f_s_dadda_rca24_fa447_y0 = f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa446_y4 ^ f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa331_y2;
  assign f_s_dadda_rca24_fa447_y1 = f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa446_y4 & f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa331_y2;
  assign f_s_dadda_rca24_fa447_y2 = f_s_dadda_rca24_fa447_y0 ^ f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa332_y2;
  assign f_s_dadda_rca24_fa447_y3 = f_s_dadda_rca24_fa447_y0 & f_s_dadda_rca24_fa447_f_s_dadda_rca24_fa332_y2;
  assign f_s_dadda_rca24_fa447_y4 = f_s_dadda_rca24_fa447_y1 | f_s_dadda_rca24_fa447_y3;
  assign f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa447_y4 = f_s_dadda_rca24_fa447_y4;
  assign f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa333_y2 = f_s_dadda_rca24_fa333_y2;
  assign f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa334_y2 = f_s_dadda_rca24_fa334_y2;
  assign f_s_dadda_rca24_fa448_y0 = f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa447_y4 ^ f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa333_y2;
  assign f_s_dadda_rca24_fa448_y1 = f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa447_y4 & f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa333_y2;
  assign f_s_dadda_rca24_fa448_y2 = f_s_dadda_rca24_fa448_y0 ^ f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa334_y2;
  assign f_s_dadda_rca24_fa448_y3 = f_s_dadda_rca24_fa448_y0 & f_s_dadda_rca24_fa448_f_s_dadda_rca24_fa334_y2;
  assign f_s_dadda_rca24_fa448_y4 = f_s_dadda_rca24_fa448_y1 | f_s_dadda_rca24_fa448_y3;
  assign f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa448_y4 = f_s_dadda_rca24_fa448_y4;
  assign f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa335_y2 = f_s_dadda_rca24_fa335_y2;
  assign f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa336_y2 = f_s_dadda_rca24_fa336_y2;
  assign f_s_dadda_rca24_fa449_y0 = f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa448_y4 ^ f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa335_y2;
  assign f_s_dadda_rca24_fa449_y1 = f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa448_y4 & f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa335_y2;
  assign f_s_dadda_rca24_fa449_y2 = f_s_dadda_rca24_fa449_y0 ^ f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa336_y2;
  assign f_s_dadda_rca24_fa449_y3 = f_s_dadda_rca24_fa449_y0 & f_s_dadda_rca24_fa449_f_s_dadda_rca24_fa336_y2;
  assign f_s_dadda_rca24_fa449_y4 = f_s_dadda_rca24_fa449_y1 | f_s_dadda_rca24_fa449_y3;
  assign f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa449_y4 = f_s_dadda_rca24_fa449_y4;
  assign f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa337_y2 = f_s_dadda_rca24_fa337_y2;
  assign f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa338_y2 = f_s_dadda_rca24_fa338_y2;
  assign f_s_dadda_rca24_fa450_y0 = f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa449_y4 ^ f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa337_y2;
  assign f_s_dadda_rca24_fa450_y1 = f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa449_y4 & f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa337_y2;
  assign f_s_dadda_rca24_fa450_y2 = f_s_dadda_rca24_fa450_y0 ^ f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa338_y2;
  assign f_s_dadda_rca24_fa450_y3 = f_s_dadda_rca24_fa450_y0 & f_s_dadda_rca24_fa450_f_s_dadda_rca24_fa338_y2;
  assign f_s_dadda_rca24_fa450_y4 = f_s_dadda_rca24_fa450_y1 | f_s_dadda_rca24_fa450_y3;
  assign f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa450_y4 = f_s_dadda_rca24_fa450_y4;
  assign f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa339_y2 = f_s_dadda_rca24_fa339_y2;
  assign f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa340_y2 = f_s_dadda_rca24_fa340_y2;
  assign f_s_dadda_rca24_fa451_y0 = f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa450_y4 ^ f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa339_y2;
  assign f_s_dadda_rca24_fa451_y1 = f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa450_y4 & f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa339_y2;
  assign f_s_dadda_rca24_fa451_y2 = f_s_dadda_rca24_fa451_y0 ^ f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa340_y2;
  assign f_s_dadda_rca24_fa451_y3 = f_s_dadda_rca24_fa451_y0 & f_s_dadda_rca24_fa451_f_s_dadda_rca24_fa340_y2;
  assign f_s_dadda_rca24_fa451_y4 = f_s_dadda_rca24_fa451_y1 | f_s_dadda_rca24_fa451_y3;
  assign f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa451_y4 = f_s_dadda_rca24_fa451_y4;
  assign f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa341_y2 = f_s_dadda_rca24_fa341_y2;
  assign f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa342_y2 = f_s_dadda_rca24_fa342_y2;
  assign f_s_dadda_rca24_fa452_y0 = f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa451_y4 ^ f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa341_y2;
  assign f_s_dadda_rca24_fa452_y1 = f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa451_y4 & f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa341_y2;
  assign f_s_dadda_rca24_fa452_y2 = f_s_dadda_rca24_fa452_y0 ^ f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa342_y2;
  assign f_s_dadda_rca24_fa452_y3 = f_s_dadda_rca24_fa452_y0 & f_s_dadda_rca24_fa452_f_s_dadda_rca24_fa342_y2;
  assign f_s_dadda_rca24_fa452_y4 = f_s_dadda_rca24_fa452_y1 | f_s_dadda_rca24_fa452_y3;
  assign f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa452_y4 = f_s_dadda_rca24_fa452_y4;
  assign f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa343_y2 = f_s_dadda_rca24_fa343_y2;
  assign f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa344_y2 = f_s_dadda_rca24_fa344_y2;
  assign f_s_dadda_rca24_fa453_y0 = f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa452_y4 ^ f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa343_y2;
  assign f_s_dadda_rca24_fa453_y1 = f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa452_y4 & f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa343_y2;
  assign f_s_dadda_rca24_fa453_y2 = f_s_dadda_rca24_fa453_y0 ^ f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa344_y2;
  assign f_s_dadda_rca24_fa453_y3 = f_s_dadda_rca24_fa453_y0 & f_s_dadda_rca24_fa453_f_s_dadda_rca24_fa344_y2;
  assign f_s_dadda_rca24_fa453_y4 = f_s_dadda_rca24_fa453_y1 | f_s_dadda_rca24_fa453_y3;
  assign f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa453_y4 = f_s_dadda_rca24_fa453_y4;
  assign f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa345_y2 = f_s_dadda_rca24_fa345_y2;
  assign f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa346_y2 = f_s_dadda_rca24_fa346_y2;
  assign f_s_dadda_rca24_fa454_y0 = f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa453_y4 ^ f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa345_y2;
  assign f_s_dadda_rca24_fa454_y1 = f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa453_y4 & f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa345_y2;
  assign f_s_dadda_rca24_fa454_y2 = f_s_dadda_rca24_fa454_y0 ^ f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa346_y2;
  assign f_s_dadda_rca24_fa454_y3 = f_s_dadda_rca24_fa454_y0 & f_s_dadda_rca24_fa454_f_s_dadda_rca24_fa346_y2;
  assign f_s_dadda_rca24_fa454_y4 = f_s_dadda_rca24_fa454_y1 | f_s_dadda_rca24_fa454_y3;
  assign f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa454_y4 = f_s_dadda_rca24_fa454_y4;
  assign f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa347_y2 = f_s_dadda_rca24_fa347_y2;
  assign f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa348_y2 = f_s_dadda_rca24_fa348_y2;
  assign f_s_dadda_rca24_fa455_y0 = f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa454_y4 ^ f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa347_y2;
  assign f_s_dadda_rca24_fa455_y1 = f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa454_y4 & f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa347_y2;
  assign f_s_dadda_rca24_fa455_y2 = f_s_dadda_rca24_fa455_y0 ^ f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa348_y2;
  assign f_s_dadda_rca24_fa455_y3 = f_s_dadda_rca24_fa455_y0 & f_s_dadda_rca24_fa455_f_s_dadda_rca24_fa348_y2;
  assign f_s_dadda_rca24_fa455_y4 = f_s_dadda_rca24_fa455_y1 | f_s_dadda_rca24_fa455_y3;
  assign f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa455_y4 = f_s_dadda_rca24_fa455_y4;
  assign f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa349_y2 = f_s_dadda_rca24_fa349_y2;
  assign f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa350_y2 = f_s_dadda_rca24_fa350_y2;
  assign f_s_dadda_rca24_fa456_y0 = f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa455_y4 ^ f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa349_y2;
  assign f_s_dadda_rca24_fa456_y1 = f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa455_y4 & f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa349_y2;
  assign f_s_dadda_rca24_fa456_y2 = f_s_dadda_rca24_fa456_y0 ^ f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa350_y2;
  assign f_s_dadda_rca24_fa456_y3 = f_s_dadda_rca24_fa456_y0 & f_s_dadda_rca24_fa456_f_s_dadda_rca24_fa350_y2;
  assign f_s_dadda_rca24_fa456_y4 = f_s_dadda_rca24_fa456_y1 | f_s_dadda_rca24_fa456_y3;
  assign f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa456_y4 = f_s_dadda_rca24_fa456_y4;
  assign f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa351_y2 = f_s_dadda_rca24_fa351_y2;
  assign f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa352_y2 = f_s_dadda_rca24_fa352_y2;
  assign f_s_dadda_rca24_fa457_y0 = f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa456_y4 ^ f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa351_y2;
  assign f_s_dadda_rca24_fa457_y1 = f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa456_y4 & f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa351_y2;
  assign f_s_dadda_rca24_fa457_y2 = f_s_dadda_rca24_fa457_y0 ^ f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa352_y2;
  assign f_s_dadda_rca24_fa457_y3 = f_s_dadda_rca24_fa457_y0 & f_s_dadda_rca24_fa457_f_s_dadda_rca24_fa352_y2;
  assign f_s_dadda_rca24_fa457_y4 = f_s_dadda_rca24_fa457_y1 | f_s_dadda_rca24_fa457_y3;
  assign f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa457_y4 = f_s_dadda_rca24_fa457_y4;
  assign f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa353_y2 = f_s_dadda_rca24_fa353_y2;
  assign f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa354_y2 = f_s_dadda_rca24_fa354_y2;
  assign f_s_dadda_rca24_fa458_y0 = f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa457_y4 ^ f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa353_y2;
  assign f_s_dadda_rca24_fa458_y1 = f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa457_y4 & f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa353_y2;
  assign f_s_dadda_rca24_fa458_y2 = f_s_dadda_rca24_fa458_y0 ^ f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa354_y2;
  assign f_s_dadda_rca24_fa458_y3 = f_s_dadda_rca24_fa458_y0 & f_s_dadda_rca24_fa458_f_s_dadda_rca24_fa354_y2;
  assign f_s_dadda_rca24_fa458_y4 = f_s_dadda_rca24_fa458_y1 | f_s_dadda_rca24_fa458_y3;
  assign f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa458_y4 = f_s_dadda_rca24_fa458_y4;
  assign f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa355_y2 = f_s_dadda_rca24_fa355_y2;
  assign f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa356_y2 = f_s_dadda_rca24_fa356_y2;
  assign f_s_dadda_rca24_fa459_y0 = f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa458_y4 ^ f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa355_y2;
  assign f_s_dadda_rca24_fa459_y1 = f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa458_y4 & f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa355_y2;
  assign f_s_dadda_rca24_fa459_y2 = f_s_dadda_rca24_fa459_y0 ^ f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa356_y2;
  assign f_s_dadda_rca24_fa459_y3 = f_s_dadda_rca24_fa459_y0 & f_s_dadda_rca24_fa459_f_s_dadda_rca24_fa356_y2;
  assign f_s_dadda_rca24_fa459_y4 = f_s_dadda_rca24_fa459_y1 | f_s_dadda_rca24_fa459_y3;
  assign f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa459_y4 = f_s_dadda_rca24_fa459_y4;
  assign f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa357_y2 = f_s_dadda_rca24_fa357_y2;
  assign f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa358_y2 = f_s_dadda_rca24_fa358_y2;
  assign f_s_dadda_rca24_fa460_y0 = f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa459_y4 ^ f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa357_y2;
  assign f_s_dadda_rca24_fa460_y1 = f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa459_y4 & f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa357_y2;
  assign f_s_dadda_rca24_fa460_y2 = f_s_dadda_rca24_fa460_y0 ^ f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa358_y2;
  assign f_s_dadda_rca24_fa460_y3 = f_s_dadda_rca24_fa460_y0 & f_s_dadda_rca24_fa460_f_s_dadda_rca24_fa358_y2;
  assign f_s_dadda_rca24_fa460_y4 = f_s_dadda_rca24_fa460_y1 | f_s_dadda_rca24_fa460_y3;
  assign f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa460_y4 = f_s_dadda_rca24_fa460_y4;
  assign f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa359_y2 = f_s_dadda_rca24_fa359_y2;
  assign f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa360_y2 = f_s_dadda_rca24_fa360_y2;
  assign f_s_dadda_rca24_fa461_y0 = f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa460_y4 ^ f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa359_y2;
  assign f_s_dadda_rca24_fa461_y1 = f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa460_y4 & f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa359_y2;
  assign f_s_dadda_rca24_fa461_y2 = f_s_dadda_rca24_fa461_y0 ^ f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa360_y2;
  assign f_s_dadda_rca24_fa461_y3 = f_s_dadda_rca24_fa461_y0 & f_s_dadda_rca24_fa461_f_s_dadda_rca24_fa360_y2;
  assign f_s_dadda_rca24_fa461_y4 = f_s_dadda_rca24_fa461_y1 | f_s_dadda_rca24_fa461_y3;
  assign f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa461_y4 = f_s_dadda_rca24_fa461_y4;
  assign f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa361_y2 = f_s_dadda_rca24_fa361_y2;
  assign f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa362_y2 = f_s_dadda_rca24_fa362_y2;
  assign f_s_dadda_rca24_fa462_y0 = f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa461_y4 ^ f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa361_y2;
  assign f_s_dadda_rca24_fa462_y1 = f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa461_y4 & f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa361_y2;
  assign f_s_dadda_rca24_fa462_y2 = f_s_dadda_rca24_fa462_y0 ^ f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa362_y2;
  assign f_s_dadda_rca24_fa462_y3 = f_s_dadda_rca24_fa462_y0 & f_s_dadda_rca24_fa462_f_s_dadda_rca24_fa362_y2;
  assign f_s_dadda_rca24_fa462_y4 = f_s_dadda_rca24_fa462_y1 | f_s_dadda_rca24_fa462_y3;
  assign f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa462_y4 = f_s_dadda_rca24_fa462_y4;
  assign f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa363_y2 = f_s_dadda_rca24_fa363_y2;
  assign f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa364_y2 = f_s_dadda_rca24_fa364_y2;
  assign f_s_dadda_rca24_fa463_y0 = f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa462_y4 ^ f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa363_y2;
  assign f_s_dadda_rca24_fa463_y1 = f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa462_y4 & f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa363_y2;
  assign f_s_dadda_rca24_fa463_y2 = f_s_dadda_rca24_fa463_y0 ^ f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa364_y2;
  assign f_s_dadda_rca24_fa463_y3 = f_s_dadda_rca24_fa463_y0 & f_s_dadda_rca24_fa463_f_s_dadda_rca24_fa364_y2;
  assign f_s_dadda_rca24_fa463_y4 = f_s_dadda_rca24_fa463_y1 | f_s_dadda_rca24_fa463_y3;
  assign f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa463_y4 = f_s_dadda_rca24_fa463_y4;
  assign f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa365_y2 = f_s_dadda_rca24_fa365_y2;
  assign f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa366_y2 = f_s_dadda_rca24_fa366_y2;
  assign f_s_dadda_rca24_fa464_y0 = f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa463_y4 ^ f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa365_y2;
  assign f_s_dadda_rca24_fa464_y1 = f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa463_y4 & f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa365_y2;
  assign f_s_dadda_rca24_fa464_y2 = f_s_dadda_rca24_fa464_y0 ^ f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa366_y2;
  assign f_s_dadda_rca24_fa464_y3 = f_s_dadda_rca24_fa464_y0 & f_s_dadda_rca24_fa464_f_s_dadda_rca24_fa366_y2;
  assign f_s_dadda_rca24_fa464_y4 = f_s_dadda_rca24_fa464_y1 | f_s_dadda_rca24_fa464_y3;
  assign f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa464_y4 = f_s_dadda_rca24_fa464_y4;
  assign f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa367_y2 = f_s_dadda_rca24_fa367_y2;
  assign f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa368_y2 = f_s_dadda_rca24_fa368_y2;
  assign f_s_dadda_rca24_fa465_y0 = f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa464_y4 ^ f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa367_y2;
  assign f_s_dadda_rca24_fa465_y1 = f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa464_y4 & f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa367_y2;
  assign f_s_dadda_rca24_fa465_y2 = f_s_dadda_rca24_fa465_y0 ^ f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa368_y2;
  assign f_s_dadda_rca24_fa465_y3 = f_s_dadda_rca24_fa465_y0 & f_s_dadda_rca24_fa465_f_s_dadda_rca24_fa368_y2;
  assign f_s_dadda_rca24_fa465_y4 = f_s_dadda_rca24_fa465_y1 | f_s_dadda_rca24_fa465_y3;
  assign f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa465_y4 = f_s_dadda_rca24_fa465_y4;
  assign f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa369_y2 = f_s_dadda_rca24_fa369_y2;
  assign f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa370_y2 = f_s_dadda_rca24_fa370_y2;
  assign f_s_dadda_rca24_fa466_y0 = f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa465_y4 ^ f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa369_y2;
  assign f_s_dadda_rca24_fa466_y1 = f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa465_y4 & f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa369_y2;
  assign f_s_dadda_rca24_fa466_y2 = f_s_dadda_rca24_fa466_y0 ^ f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa370_y2;
  assign f_s_dadda_rca24_fa466_y3 = f_s_dadda_rca24_fa466_y0 & f_s_dadda_rca24_fa466_f_s_dadda_rca24_fa370_y2;
  assign f_s_dadda_rca24_fa466_y4 = f_s_dadda_rca24_fa466_y1 | f_s_dadda_rca24_fa466_y3;
  assign f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa466_y4 = f_s_dadda_rca24_fa466_y4;
  assign f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa371_y2 = f_s_dadda_rca24_fa371_y2;
  assign f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa372_y2 = f_s_dadda_rca24_fa372_y2;
  assign f_s_dadda_rca24_fa467_y0 = f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa466_y4 ^ f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa371_y2;
  assign f_s_dadda_rca24_fa467_y1 = f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa466_y4 & f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa371_y2;
  assign f_s_dadda_rca24_fa467_y2 = f_s_dadda_rca24_fa467_y0 ^ f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa372_y2;
  assign f_s_dadda_rca24_fa467_y3 = f_s_dadda_rca24_fa467_y0 & f_s_dadda_rca24_fa467_f_s_dadda_rca24_fa372_y2;
  assign f_s_dadda_rca24_fa467_y4 = f_s_dadda_rca24_fa467_y1 | f_s_dadda_rca24_fa467_y3;
  assign f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa467_y4 = f_s_dadda_rca24_fa467_y4;
  assign f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa373_y2 = f_s_dadda_rca24_fa373_y2;
  assign f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa374_y2 = f_s_dadda_rca24_fa374_y2;
  assign f_s_dadda_rca24_fa468_y0 = f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa467_y4 ^ f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa373_y2;
  assign f_s_dadda_rca24_fa468_y1 = f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa467_y4 & f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa373_y2;
  assign f_s_dadda_rca24_fa468_y2 = f_s_dadda_rca24_fa468_y0 ^ f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa374_y2;
  assign f_s_dadda_rca24_fa468_y3 = f_s_dadda_rca24_fa468_y0 & f_s_dadda_rca24_fa468_f_s_dadda_rca24_fa374_y2;
  assign f_s_dadda_rca24_fa468_y4 = f_s_dadda_rca24_fa468_y1 | f_s_dadda_rca24_fa468_y3;
  assign f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa468_y4 = f_s_dadda_rca24_fa468_y4;
  assign f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa375_y2 = f_s_dadda_rca24_fa375_y2;
  assign f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa376_y2 = f_s_dadda_rca24_fa376_y2;
  assign f_s_dadda_rca24_fa469_y0 = f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa468_y4 ^ f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa375_y2;
  assign f_s_dadda_rca24_fa469_y1 = f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa468_y4 & f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa375_y2;
  assign f_s_dadda_rca24_fa469_y2 = f_s_dadda_rca24_fa469_y0 ^ f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa376_y2;
  assign f_s_dadda_rca24_fa469_y3 = f_s_dadda_rca24_fa469_y0 & f_s_dadda_rca24_fa469_f_s_dadda_rca24_fa376_y2;
  assign f_s_dadda_rca24_fa469_y4 = f_s_dadda_rca24_fa469_y1 | f_s_dadda_rca24_fa469_y3;
  assign f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa469_y4 = f_s_dadda_rca24_fa469_y4;
  assign f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa377_y2 = f_s_dadda_rca24_fa377_y2;
  assign f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa378_y2 = f_s_dadda_rca24_fa378_y2;
  assign f_s_dadda_rca24_fa470_y0 = f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa469_y4 ^ f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa377_y2;
  assign f_s_dadda_rca24_fa470_y1 = f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa469_y4 & f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa377_y2;
  assign f_s_dadda_rca24_fa470_y2 = f_s_dadda_rca24_fa470_y0 ^ f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa378_y2;
  assign f_s_dadda_rca24_fa470_y3 = f_s_dadda_rca24_fa470_y0 & f_s_dadda_rca24_fa470_f_s_dadda_rca24_fa378_y2;
  assign f_s_dadda_rca24_fa470_y4 = f_s_dadda_rca24_fa470_y1 | f_s_dadda_rca24_fa470_y3;
  assign f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa470_y4 = f_s_dadda_rca24_fa470_y4;
  assign f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa379_y2 = f_s_dadda_rca24_fa379_y2;
  assign f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa380_y2 = f_s_dadda_rca24_fa380_y2;
  assign f_s_dadda_rca24_fa471_y0 = f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa470_y4 ^ f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa379_y2;
  assign f_s_dadda_rca24_fa471_y1 = f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa470_y4 & f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa379_y2;
  assign f_s_dadda_rca24_fa471_y2 = f_s_dadda_rca24_fa471_y0 ^ f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa380_y2;
  assign f_s_dadda_rca24_fa471_y3 = f_s_dadda_rca24_fa471_y0 & f_s_dadda_rca24_fa471_f_s_dadda_rca24_fa380_y2;
  assign f_s_dadda_rca24_fa471_y4 = f_s_dadda_rca24_fa471_y1 | f_s_dadda_rca24_fa471_y3;
  assign f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa471_y4 = f_s_dadda_rca24_fa471_y4;
  assign f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa381_y2 = f_s_dadda_rca24_fa381_y2;
  assign f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa382_y2 = f_s_dadda_rca24_fa382_y2;
  assign f_s_dadda_rca24_fa472_y0 = f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa471_y4 ^ f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa381_y2;
  assign f_s_dadda_rca24_fa472_y1 = f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa471_y4 & f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa381_y2;
  assign f_s_dadda_rca24_fa472_y2 = f_s_dadda_rca24_fa472_y0 ^ f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa382_y2;
  assign f_s_dadda_rca24_fa472_y3 = f_s_dadda_rca24_fa472_y0 & f_s_dadda_rca24_fa472_f_s_dadda_rca24_fa382_y2;
  assign f_s_dadda_rca24_fa472_y4 = f_s_dadda_rca24_fa472_y1 | f_s_dadda_rca24_fa472_y3;
  assign f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa472_y4 = f_s_dadda_rca24_fa472_y4;
  assign f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa383_y2 = f_s_dadda_rca24_fa383_y2;
  assign f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa384_y2 = f_s_dadda_rca24_fa384_y2;
  assign f_s_dadda_rca24_fa473_y0 = f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa472_y4 ^ f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa383_y2;
  assign f_s_dadda_rca24_fa473_y1 = f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa472_y4 & f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa383_y2;
  assign f_s_dadda_rca24_fa473_y2 = f_s_dadda_rca24_fa473_y0 ^ f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa384_y2;
  assign f_s_dadda_rca24_fa473_y3 = f_s_dadda_rca24_fa473_y0 & f_s_dadda_rca24_fa473_f_s_dadda_rca24_fa384_y2;
  assign f_s_dadda_rca24_fa473_y4 = f_s_dadda_rca24_fa473_y1 | f_s_dadda_rca24_fa473_y3;
  assign f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa473_y4 = f_s_dadda_rca24_fa473_y4;
  assign f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa385_y2 = f_s_dadda_rca24_fa385_y2;
  assign f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa386_y2 = f_s_dadda_rca24_fa386_y2;
  assign f_s_dadda_rca24_fa474_y0 = f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa473_y4 ^ f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa385_y2;
  assign f_s_dadda_rca24_fa474_y1 = f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa473_y4 & f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa385_y2;
  assign f_s_dadda_rca24_fa474_y2 = f_s_dadda_rca24_fa474_y0 ^ f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa386_y2;
  assign f_s_dadda_rca24_fa474_y3 = f_s_dadda_rca24_fa474_y0 & f_s_dadda_rca24_fa474_f_s_dadda_rca24_fa386_y2;
  assign f_s_dadda_rca24_fa474_y4 = f_s_dadda_rca24_fa474_y1 | f_s_dadda_rca24_fa474_y3;
  assign f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa474_y4 = f_s_dadda_rca24_fa474_y4;
  assign f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa387_y2 = f_s_dadda_rca24_fa387_y2;
  assign f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa388_y2 = f_s_dadda_rca24_fa388_y2;
  assign f_s_dadda_rca24_fa475_y0 = f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa474_y4 ^ f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa387_y2;
  assign f_s_dadda_rca24_fa475_y1 = f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa474_y4 & f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa387_y2;
  assign f_s_dadda_rca24_fa475_y2 = f_s_dadda_rca24_fa475_y0 ^ f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa388_y2;
  assign f_s_dadda_rca24_fa475_y3 = f_s_dadda_rca24_fa475_y0 & f_s_dadda_rca24_fa475_f_s_dadda_rca24_fa388_y2;
  assign f_s_dadda_rca24_fa475_y4 = f_s_dadda_rca24_fa475_y1 | f_s_dadda_rca24_fa475_y3;
  assign f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa475_y4 = f_s_dadda_rca24_fa475_y4;
  assign f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa389_y2 = f_s_dadda_rca24_fa389_y2;
  assign f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa390_y2 = f_s_dadda_rca24_fa390_y2;
  assign f_s_dadda_rca24_fa476_y0 = f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa475_y4 ^ f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa389_y2;
  assign f_s_dadda_rca24_fa476_y1 = f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa475_y4 & f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa389_y2;
  assign f_s_dadda_rca24_fa476_y2 = f_s_dadda_rca24_fa476_y0 ^ f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa390_y2;
  assign f_s_dadda_rca24_fa476_y3 = f_s_dadda_rca24_fa476_y0 & f_s_dadda_rca24_fa476_f_s_dadda_rca24_fa390_y2;
  assign f_s_dadda_rca24_fa476_y4 = f_s_dadda_rca24_fa476_y1 | f_s_dadda_rca24_fa476_y3;
  assign f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa476_y4 = f_s_dadda_rca24_fa476_y4;
  assign f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa391_y2 = f_s_dadda_rca24_fa391_y2;
  assign f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa392_y2 = f_s_dadda_rca24_fa392_y2;
  assign f_s_dadda_rca24_fa477_y0 = f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa476_y4 ^ f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa391_y2;
  assign f_s_dadda_rca24_fa477_y1 = f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa476_y4 & f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa391_y2;
  assign f_s_dadda_rca24_fa477_y2 = f_s_dadda_rca24_fa477_y0 ^ f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa392_y2;
  assign f_s_dadda_rca24_fa477_y3 = f_s_dadda_rca24_fa477_y0 & f_s_dadda_rca24_fa477_f_s_dadda_rca24_fa392_y2;
  assign f_s_dadda_rca24_fa477_y4 = f_s_dadda_rca24_fa477_y1 | f_s_dadda_rca24_fa477_y3;
  assign f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa477_y4 = f_s_dadda_rca24_fa477_y4;
  assign f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa393_y2 = f_s_dadda_rca24_fa393_y2;
  assign f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa394_y2 = f_s_dadda_rca24_fa394_y2;
  assign f_s_dadda_rca24_fa478_y0 = f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa477_y4 ^ f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa393_y2;
  assign f_s_dadda_rca24_fa478_y1 = f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa477_y4 & f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa393_y2;
  assign f_s_dadda_rca24_fa478_y2 = f_s_dadda_rca24_fa478_y0 ^ f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa394_y2;
  assign f_s_dadda_rca24_fa478_y3 = f_s_dadda_rca24_fa478_y0 & f_s_dadda_rca24_fa478_f_s_dadda_rca24_fa394_y2;
  assign f_s_dadda_rca24_fa478_y4 = f_s_dadda_rca24_fa478_y1 | f_s_dadda_rca24_fa478_y3;
  assign f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa478_y4 = f_s_dadda_rca24_fa478_y4;
  assign f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa395_y2 = f_s_dadda_rca24_fa395_y2;
  assign f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa396_y2 = f_s_dadda_rca24_fa396_y2;
  assign f_s_dadda_rca24_fa479_y0 = f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa478_y4 ^ f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa395_y2;
  assign f_s_dadda_rca24_fa479_y1 = f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa478_y4 & f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa395_y2;
  assign f_s_dadda_rca24_fa479_y2 = f_s_dadda_rca24_fa479_y0 ^ f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa396_y2;
  assign f_s_dadda_rca24_fa479_y3 = f_s_dadda_rca24_fa479_y0 & f_s_dadda_rca24_fa479_f_s_dadda_rca24_fa396_y2;
  assign f_s_dadda_rca24_fa479_y4 = f_s_dadda_rca24_fa479_y1 | f_s_dadda_rca24_fa479_y3;
  assign f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa479_y4 = f_s_dadda_rca24_fa479_y4;
  assign f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa397_y2 = f_s_dadda_rca24_fa397_y2;
  assign f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa398_y2 = f_s_dadda_rca24_fa398_y2;
  assign f_s_dadda_rca24_fa480_y0 = f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa479_y4 ^ f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa397_y2;
  assign f_s_dadda_rca24_fa480_y1 = f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa479_y4 & f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa397_y2;
  assign f_s_dadda_rca24_fa480_y2 = f_s_dadda_rca24_fa480_y0 ^ f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa398_y2;
  assign f_s_dadda_rca24_fa480_y3 = f_s_dadda_rca24_fa480_y0 & f_s_dadda_rca24_fa480_f_s_dadda_rca24_fa398_y2;
  assign f_s_dadda_rca24_fa480_y4 = f_s_dadda_rca24_fa480_y1 | f_s_dadda_rca24_fa480_y3;
  assign f_s_dadda_rca24_nand_20_23_a_20 = a_20;
  assign f_s_dadda_rca24_nand_20_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_20_23_y0 = ~(f_s_dadda_rca24_nand_20_23_a_20 & f_s_dadda_rca24_nand_20_23_b_23);
  assign f_s_dadda_rca24_fa481_f_s_dadda_rca24_fa480_y4 = f_s_dadda_rca24_fa480_y4;
  assign f_s_dadda_rca24_fa481_f_s_dadda_rca24_nand_20_23_y0 = f_s_dadda_rca24_nand_20_23_y0;
  assign f_s_dadda_rca24_fa481_f_s_dadda_rca24_fa399_y2 = f_s_dadda_rca24_fa399_y2;
  assign f_s_dadda_rca24_fa481_y0 = f_s_dadda_rca24_fa481_f_s_dadda_rca24_fa480_y4 ^ f_s_dadda_rca24_fa481_f_s_dadda_rca24_nand_20_23_y0;
  assign f_s_dadda_rca24_fa481_y1 = f_s_dadda_rca24_fa481_f_s_dadda_rca24_fa480_y4 & f_s_dadda_rca24_fa481_f_s_dadda_rca24_nand_20_23_y0;
  assign f_s_dadda_rca24_fa481_y2 = f_s_dadda_rca24_fa481_y0 ^ f_s_dadda_rca24_fa481_f_s_dadda_rca24_fa399_y2;
  assign f_s_dadda_rca24_fa481_y3 = f_s_dadda_rca24_fa481_y0 & f_s_dadda_rca24_fa481_f_s_dadda_rca24_fa399_y2;
  assign f_s_dadda_rca24_fa481_y4 = f_s_dadda_rca24_fa481_y1 | f_s_dadda_rca24_fa481_y3;
  assign f_s_dadda_rca24_and_22_22_a_22 = a_22;
  assign f_s_dadda_rca24_and_22_22_b_22 = b_22;
  assign f_s_dadda_rca24_and_22_22_y0 = f_s_dadda_rca24_and_22_22_a_22 & f_s_dadda_rca24_and_22_22_b_22;
  assign f_s_dadda_rca24_nand_21_23_a_21 = a_21;
  assign f_s_dadda_rca24_nand_21_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_21_23_y0 = ~(f_s_dadda_rca24_nand_21_23_a_21 & f_s_dadda_rca24_nand_21_23_b_23);
  assign f_s_dadda_rca24_fa482_f_s_dadda_rca24_fa481_y4 = f_s_dadda_rca24_fa481_y4;
  assign f_s_dadda_rca24_fa482_f_s_dadda_rca24_and_22_22_y0 = f_s_dadda_rca24_and_22_22_y0;
  assign f_s_dadda_rca24_fa482_f_s_dadda_rca24_nand_21_23_y0 = f_s_dadda_rca24_nand_21_23_y0;
  assign f_s_dadda_rca24_fa482_y0 = f_s_dadda_rca24_fa482_f_s_dadda_rca24_fa481_y4 ^ f_s_dadda_rca24_fa482_f_s_dadda_rca24_and_22_22_y0;
  assign f_s_dadda_rca24_fa482_y1 = f_s_dadda_rca24_fa482_f_s_dadda_rca24_fa481_y4 & f_s_dadda_rca24_fa482_f_s_dadda_rca24_and_22_22_y0;
  assign f_s_dadda_rca24_fa482_y2 = f_s_dadda_rca24_fa482_y0 ^ f_s_dadda_rca24_fa482_f_s_dadda_rca24_nand_21_23_y0;
  assign f_s_dadda_rca24_fa482_y3 = f_s_dadda_rca24_fa482_y0 & f_s_dadda_rca24_fa482_f_s_dadda_rca24_nand_21_23_y0;
  assign f_s_dadda_rca24_fa482_y4 = f_s_dadda_rca24_fa482_y1 | f_s_dadda_rca24_fa482_y3;
  assign f_s_dadda_rca24_nand_23_22_a_23 = a_23;
  assign f_s_dadda_rca24_nand_23_22_b_22 = b_22;
  assign f_s_dadda_rca24_nand_23_22_y0 = ~(f_s_dadda_rca24_nand_23_22_a_23 & f_s_dadda_rca24_nand_23_22_b_22);
  assign f_s_dadda_rca24_fa483_f_s_dadda_rca24_fa482_y4 = f_s_dadda_rca24_fa482_y4;
  assign f_s_dadda_rca24_fa483_f_s_dadda_rca24_fa440_y4 = f_s_dadda_rca24_fa440_y4;
  assign f_s_dadda_rca24_fa483_f_s_dadda_rca24_nand_23_22_y0 = f_s_dadda_rca24_nand_23_22_y0;
  assign f_s_dadda_rca24_fa483_y0 = f_s_dadda_rca24_fa483_f_s_dadda_rca24_fa482_y4 ^ f_s_dadda_rca24_fa483_f_s_dadda_rca24_fa440_y4;
  assign f_s_dadda_rca24_fa483_y1 = f_s_dadda_rca24_fa483_f_s_dadda_rca24_fa482_y4 & f_s_dadda_rca24_fa483_f_s_dadda_rca24_fa440_y4;
  assign f_s_dadda_rca24_fa483_y2 = f_s_dadda_rca24_fa483_y0 ^ f_s_dadda_rca24_fa483_f_s_dadda_rca24_nand_23_22_y0;
  assign f_s_dadda_rca24_fa483_y3 = f_s_dadda_rca24_fa483_y0 & f_s_dadda_rca24_fa483_f_s_dadda_rca24_nand_23_22_y0;
  assign f_s_dadda_rca24_fa483_y4 = f_s_dadda_rca24_fa483_y1 | f_s_dadda_rca24_fa483_y3;
  assign f_s_dadda_rca24_and_0_0_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_0_0_y0 = f_s_dadda_rca24_and_0_0_a_0 & f_s_dadda_rca24_and_0_0_b_0;
  assign f_s_dadda_rca24_and_1_0_a_1 = a_1;
  assign f_s_dadda_rca24_and_1_0_b_0 = b_0;
  assign f_s_dadda_rca24_and_1_0_y0 = f_s_dadda_rca24_and_1_0_a_1 & f_s_dadda_rca24_and_1_0_b_0;
  assign f_s_dadda_rca24_and_0_2_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_2_b_2 = b_2;
  assign f_s_dadda_rca24_and_0_2_y0 = f_s_dadda_rca24_and_0_2_a_0 & f_s_dadda_rca24_and_0_2_b_2;
  assign f_s_dadda_rca24_nand_22_23_a_22 = a_22;
  assign f_s_dadda_rca24_nand_22_23_b_23 = b_23;
  assign f_s_dadda_rca24_nand_22_23_y0 = ~(f_s_dadda_rca24_nand_22_23_a_22 & f_s_dadda_rca24_nand_22_23_b_23);
  assign f_s_dadda_rca24_and_0_1_a_0 = a_0;
  assign f_s_dadda_rca24_and_0_1_b_1 = b_1;
  assign f_s_dadda_rca24_and_0_1_y0 = f_s_dadda_rca24_and_0_1_a_0 & f_s_dadda_rca24_and_0_1_b_1;
  assign f_s_dadda_rca24_and_23_23_a_23 = a_23;
  assign f_s_dadda_rca24_and_23_23_b_23 = b_23;
  assign f_s_dadda_rca24_and_23_23_y0 = f_s_dadda_rca24_and_23_23_a_23 & f_s_dadda_rca24_and_23_23_b_23;
  assign f_s_dadda_rca24_u_rca_ha_f_s_dadda_rca24_and_1_0_y0 = f_s_dadda_rca24_and_1_0_y0;
  assign f_s_dadda_rca24_u_rca_ha_f_s_dadda_rca24_and_0_1_y0 = f_s_dadda_rca24_and_0_1_y0;
  assign f_s_dadda_rca24_u_rca_ha_y0 = f_s_dadda_rca24_u_rca_ha_f_s_dadda_rca24_and_1_0_y0 ^ f_s_dadda_rca24_u_rca_ha_f_s_dadda_rca24_and_0_1_y0;
  assign f_s_dadda_rca24_u_rca_ha_y1 = f_s_dadda_rca24_u_rca_ha_f_s_dadda_rca24_and_1_0_y0 & f_s_dadda_rca24_u_rca_ha_f_s_dadda_rca24_and_0_1_y0;
  assign f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_and_0_2_y0 = f_s_dadda_rca24_and_0_2_y0;
  assign f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_ha21_y0 = f_s_dadda_rca24_ha21_y0;
  assign f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_u_rca_ha_y1 = f_s_dadda_rca24_u_rca_ha_y1;
  assign f_s_dadda_rca24_u_rca_fa1_y0 = f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_and_0_2_y0 ^ f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_ha21_y0;
  assign f_s_dadda_rca24_u_rca_fa1_y1 = f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_and_0_2_y0 & f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_ha21_y0;
  assign f_s_dadda_rca24_u_rca_fa1_y2 = f_s_dadda_rca24_u_rca_fa1_y0 ^ f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_u_rca_ha_y1;
  assign f_s_dadda_rca24_u_rca_fa1_y3 = f_s_dadda_rca24_u_rca_fa1_y0 & f_s_dadda_rca24_u_rca_fa1_f_s_dadda_rca24_u_rca_ha_y1;
  assign f_s_dadda_rca24_u_rca_fa1_y4 = f_s_dadda_rca24_u_rca_fa1_y1 | f_s_dadda_rca24_u_rca_fa1_y3;
  assign f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_ha20_y0 = f_s_dadda_rca24_ha20_y0;
  assign f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_fa441_y2 = f_s_dadda_rca24_fa441_y2;
  assign f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_u_rca_fa1_y4 = f_s_dadda_rca24_u_rca_fa1_y4;
  assign f_s_dadda_rca24_u_rca_fa2_y0 = f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_ha20_y0 ^ f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_fa441_y2;
  assign f_s_dadda_rca24_u_rca_fa2_y1 = f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_ha20_y0 & f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_fa441_y2;
  assign f_s_dadda_rca24_u_rca_fa2_y2 = f_s_dadda_rca24_u_rca_fa2_y0 ^ f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_u_rca_fa1_y4;
  assign f_s_dadda_rca24_u_rca_fa2_y3 = f_s_dadda_rca24_u_rca_fa2_y0 & f_s_dadda_rca24_u_rca_fa2_f_s_dadda_rca24_u_rca_fa1_y4;
  assign f_s_dadda_rca24_u_rca_fa2_y4 = f_s_dadda_rca24_u_rca_fa2_y1 | f_s_dadda_rca24_u_rca_fa2_y3;
  assign f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_fa400_y2 = f_s_dadda_rca24_fa400_y2;
  assign f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_fa442_y2 = f_s_dadda_rca24_fa442_y2;
  assign f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_u_rca_fa2_y4 = f_s_dadda_rca24_u_rca_fa2_y4;
  assign f_s_dadda_rca24_u_rca_fa3_y0 = f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_fa400_y2 ^ f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_fa442_y2;
  assign f_s_dadda_rca24_u_rca_fa3_y1 = f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_fa400_y2 & f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_fa442_y2;
  assign f_s_dadda_rca24_u_rca_fa3_y2 = f_s_dadda_rca24_u_rca_fa3_y0 ^ f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_u_rca_fa2_y4;
  assign f_s_dadda_rca24_u_rca_fa3_y3 = f_s_dadda_rca24_u_rca_fa3_y0 & f_s_dadda_rca24_u_rca_fa3_f_s_dadda_rca24_u_rca_fa2_y4;
  assign f_s_dadda_rca24_u_rca_fa3_y4 = f_s_dadda_rca24_u_rca_fa3_y1 | f_s_dadda_rca24_u_rca_fa3_y3;
  assign f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_fa401_y2 = f_s_dadda_rca24_fa401_y2;
  assign f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_fa443_y2 = f_s_dadda_rca24_fa443_y2;
  assign f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_u_rca_fa3_y4 = f_s_dadda_rca24_u_rca_fa3_y4;
  assign f_s_dadda_rca24_u_rca_fa4_y0 = f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_fa401_y2 ^ f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_fa443_y2;
  assign f_s_dadda_rca24_u_rca_fa4_y1 = f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_fa401_y2 & f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_fa443_y2;
  assign f_s_dadda_rca24_u_rca_fa4_y2 = f_s_dadda_rca24_u_rca_fa4_y0 ^ f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_u_rca_fa3_y4;
  assign f_s_dadda_rca24_u_rca_fa4_y3 = f_s_dadda_rca24_u_rca_fa4_y0 & f_s_dadda_rca24_u_rca_fa4_f_s_dadda_rca24_u_rca_fa3_y4;
  assign f_s_dadda_rca24_u_rca_fa4_y4 = f_s_dadda_rca24_u_rca_fa4_y1 | f_s_dadda_rca24_u_rca_fa4_y3;
  assign f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_fa402_y2 = f_s_dadda_rca24_fa402_y2;
  assign f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_fa444_y2 = f_s_dadda_rca24_fa444_y2;
  assign f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_u_rca_fa4_y4 = f_s_dadda_rca24_u_rca_fa4_y4;
  assign f_s_dadda_rca24_u_rca_fa5_y0 = f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_fa402_y2 ^ f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_fa444_y2;
  assign f_s_dadda_rca24_u_rca_fa5_y1 = f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_fa402_y2 & f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_fa444_y2;
  assign f_s_dadda_rca24_u_rca_fa5_y2 = f_s_dadda_rca24_u_rca_fa5_y0 ^ f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_u_rca_fa4_y4;
  assign f_s_dadda_rca24_u_rca_fa5_y3 = f_s_dadda_rca24_u_rca_fa5_y0 & f_s_dadda_rca24_u_rca_fa5_f_s_dadda_rca24_u_rca_fa4_y4;
  assign f_s_dadda_rca24_u_rca_fa5_y4 = f_s_dadda_rca24_u_rca_fa5_y1 | f_s_dadda_rca24_u_rca_fa5_y3;
  assign f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_fa403_y2 = f_s_dadda_rca24_fa403_y2;
  assign f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_fa445_y2 = f_s_dadda_rca24_fa445_y2;
  assign f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_u_rca_fa5_y4 = f_s_dadda_rca24_u_rca_fa5_y4;
  assign f_s_dadda_rca24_u_rca_fa6_y0 = f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_fa403_y2 ^ f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_fa445_y2;
  assign f_s_dadda_rca24_u_rca_fa6_y1 = f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_fa403_y2 & f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_fa445_y2;
  assign f_s_dadda_rca24_u_rca_fa6_y2 = f_s_dadda_rca24_u_rca_fa6_y0 ^ f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_u_rca_fa5_y4;
  assign f_s_dadda_rca24_u_rca_fa6_y3 = f_s_dadda_rca24_u_rca_fa6_y0 & f_s_dadda_rca24_u_rca_fa6_f_s_dadda_rca24_u_rca_fa5_y4;
  assign f_s_dadda_rca24_u_rca_fa6_y4 = f_s_dadda_rca24_u_rca_fa6_y1 | f_s_dadda_rca24_u_rca_fa6_y3;
  assign f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_fa404_y2 = f_s_dadda_rca24_fa404_y2;
  assign f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_fa446_y2 = f_s_dadda_rca24_fa446_y2;
  assign f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_u_rca_fa6_y4 = f_s_dadda_rca24_u_rca_fa6_y4;
  assign f_s_dadda_rca24_u_rca_fa7_y0 = f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_fa404_y2 ^ f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_fa446_y2;
  assign f_s_dadda_rca24_u_rca_fa7_y1 = f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_fa404_y2 & f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_fa446_y2;
  assign f_s_dadda_rca24_u_rca_fa7_y2 = f_s_dadda_rca24_u_rca_fa7_y0 ^ f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_u_rca_fa6_y4;
  assign f_s_dadda_rca24_u_rca_fa7_y3 = f_s_dadda_rca24_u_rca_fa7_y0 & f_s_dadda_rca24_u_rca_fa7_f_s_dadda_rca24_u_rca_fa6_y4;
  assign f_s_dadda_rca24_u_rca_fa7_y4 = f_s_dadda_rca24_u_rca_fa7_y1 | f_s_dadda_rca24_u_rca_fa7_y3;
  assign f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_fa405_y2 = f_s_dadda_rca24_fa405_y2;
  assign f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_fa447_y2 = f_s_dadda_rca24_fa447_y2;
  assign f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_u_rca_fa7_y4 = f_s_dadda_rca24_u_rca_fa7_y4;
  assign f_s_dadda_rca24_u_rca_fa8_y0 = f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_fa405_y2 ^ f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_fa447_y2;
  assign f_s_dadda_rca24_u_rca_fa8_y1 = f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_fa405_y2 & f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_fa447_y2;
  assign f_s_dadda_rca24_u_rca_fa8_y2 = f_s_dadda_rca24_u_rca_fa8_y0 ^ f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_u_rca_fa7_y4;
  assign f_s_dadda_rca24_u_rca_fa8_y3 = f_s_dadda_rca24_u_rca_fa8_y0 & f_s_dadda_rca24_u_rca_fa8_f_s_dadda_rca24_u_rca_fa7_y4;
  assign f_s_dadda_rca24_u_rca_fa8_y4 = f_s_dadda_rca24_u_rca_fa8_y1 | f_s_dadda_rca24_u_rca_fa8_y3;
  assign f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_fa406_y2 = f_s_dadda_rca24_fa406_y2;
  assign f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_fa448_y2 = f_s_dadda_rca24_fa448_y2;
  assign f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_u_rca_fa8_y4 = f_s_dadda_rca24_u_rca_fa8_y4;
  assign f_s_dadda_rca24_u_rca_fa9_y0 = f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_fa406_y2 ^ f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_fa448_y2;
  assign f_s_dadda_rca24_u_rca_fa9_y1 = f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_fa406_y2 & f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_fa448_y2;
  assign f_s_dadda_rca24_u_rca_fa9_y2 = f_s_dadda_rca24_u_rca_fa9_y0 ^ f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_u_rca_fa8_y4;
  assign f_s_dadda_rca24_u_rca_fa9_y3 = f_s_dadda_rca24_u_rca_fa9_y0 & f_s_dadda_rca24_u_rca_fa9_f_s_dadda_rca24_u_rca_fa8_y4;
  assign f_s_dadda_rca24_u_rca_fa9_y4 = f_s_dadda_rca24_u_rca_fa9_y1 | f_s_dadda_rca24_u_rca_fa9_y3;
  assign f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_fa407_y2 = f_s_dadda_rca24_fa407_y2;
  assign f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_fa449_y2 = f_s_dadda_rca24_fa449_y2;
  assign f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_u_rca_fa9_y4 = f_s_dadda_rca24_u_rca_fa9_y4;
  assign f_s_dadda_rca24_u_rca_fa10_y0 = f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_fa407_y2 ^ f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_fa449_y2;
  assign f_s_dadda_rca24_u_rca_fa10_y1 = f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_fa407_y2 & f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_fa449_y2;
  assign f_s_dadda_rca24_u_rca_fa10_y2 = f_s_dadda_rca24_u_rca_fa10_y0 ^ f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_u_rca_fa9_y4;
  assign f_s_dadda_rca24_u_rca_fa10_y3 = f_s_dadda_rca24_u_rca_fa10_y0 & f_s_dadda_rca24_u_rca_fa10_f_s_dadda_rca24_u_rca_fa9_y4;
  assign f_s_dadda_rca24_u_rca_fa10_y4 = f_s_dadda_rca24_u_rca_fa10_y1 | f_s_dadda_rca24_u_rca_fa10_y3;
  assign f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_fa408_y2 = f_s_dadda_rca24_fa408_y2;
  assign f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_fa450_y2 = f_s_dadda_rca24_fa450_y2;
  assign f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_u_rca_fa10_y4 = f_s_dadda_rca24_u_rca_fa10_y4;
  assign f_s_dadda_rca24_u_rca_fa11_y0 = f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_fa408_y2 ^ f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_fa450_y2;
  assign f_s_dadda_rca24_u_rca_fa11_y1 = f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_fa408_y2 & f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_fa450_y2;
  assign f_s_dadda_rca24_u_rca_fa11_y2 = f_s_dadda_rca24_u_rca_fa11_y0 ^ f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_u_rca_fa10_y4;
  assign f_s_dadda_rca24_u_rca_fa11_y3 = f_s_dadda_rca24_u_rca_fa11_y0 & f_s_dadda_rca24_u_rca_fa11_f_s_dadda_rca24_u_rca_fa10_y4;
  assign f_s_dadda_rca24_u_rca_fa11_y4 = f_s_dadda_rca24_u_rca_fa11_y1 | f_s_dadda_rca24_u_rca_fa11_y3;
  assign f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_fa409_y2 = f_s_dadda_rca24_fa409_y2;
  assign f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_fa451_y2 = f_s_dadda_rca24_fa451_y2;
  assign f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_u_rca_fa11_y4 = f_s_dadda_rca24_u_rca_fa11_y4;
  assign f_s_dadda_rca24_u_rca_fa12_y0 = f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_fa409_y2 ^ f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_fa451_y2;
  assign f_s_dadda_rca24_u_rca_fa12_y1 = f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_fa409_y2 & f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_fa451_y2;
  assign f_s_dadda_rca24_u_rca_fa12_y2 = f_s_dadda_rca24_u_rca_fa12_y0 ^ f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_u_rca_fa11_y4;
  assign f_s_dadda_rca24_u_rca_fa12_y3 = f_s_dadda_rca24_u_rca_fa12_y0 & f_s_dadda_rca24_u_rca_fa12_f_s_dadda_rca24_u_rca_fa11_y4;
  assign f_s_dadda_rca24_u_rca_fa12_y4 = f_s_dadda_rca24_u_rca_fa12_y1 | f_s_dadda_rca24_u_rca_fa12_y3;
  assign f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_fa410_y2 = f_s_dadda_rca24_fa410_y2;
  assign f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_fa452_y2 = f_s_dadda_rca24_fa452_y2;
  assign f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_u_rca_fa12_y4 = f_s_dadda_rca24_u_rca_fa12_y4;
  assign f_s_dadda_rca24_u_rca_fa13_y0 = f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_fa410_y2 ^ f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_fa452_y2;
  assign f_s_dadda_rca24_u_rca_fa13_y1 = f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_fa410_y2 & f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_fa452_y2;
  assign f_s_dadda_rca24_u_rca_fa13_y2 = f_s_dadda_rca24_u_rca_fa13_y0 ^ f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_u_rca_fa12_y4;
  assign f_s_dadda_rca24_u_rca_fa13_y3 = f_s_dadda_rca24_u_rca_fa13_y0 & f_s_dadda_rca24_u_rca_fa13_f_s_dadda_rca24_u_rca_fa12_y4;
  assign f_s_dadda_rca24_u_rca_fa13_y4 = f_s_dadda_rca24_u_rca_fa13_y1 | f_s_dadda_rca24_u_rca_fa13_y3;
  assign f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_fa411_y2 = f_s_dadda_rca24_fa411_y2;
  assign f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_fa453_y2 = f_s_dadda_rca24_fa453_y2;
  assign f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_u_rca_fa13_y4 = f_s_dadda_rca24_u_rca_fa13_y4;
  assign f_s_dadda_rca24_u_rca_fa14_y0 = f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_fa411_y2 ^ f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_fa453_y2;
  assign f_s_dadda_rca24_u_rca_fa14_y1 = f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_fa411_y2 & f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_fa453_y2;
  assign f_s_dadda_rca24_u_rca_fa14_y2 = f_s_dadda_rca24_u_rca_fa14_y0 ^ f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_u_rca_fa13_y4;
  assign f_s_dadda_rca24_u_rca_fa14_y3 = f_s_dadda_rca24_u_rca_fa14_y0 & f_s_dadda_rca24_u_rca_fa14_f_s_dadda_rca24_u_rca_fa13_y4;
  assign f_s_dadda_rca24_u_rca_fa14_y4 = f_s_dadda_rca24_u_rca_fa14_y1 | f_s_dadda_rca24_u_rca_fa14_y3;
  assign f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_fa412_y2 = f_s_dadda_rca24_fa412_y2;
  assign f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_fa454_y2 = f_s_dadda_rca24_fa454_y2;
  assign f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_u_rca_fa14_y4 = f_s_dadda_rca24_u_rca_fa14_y4;
  assign f_s_dadda_rca24_u_rca_fa15_y0 = f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_fa412_y2 ^ f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_fa454_y2;
  assign f_s_dadda_rca24_u_rca_fa15_y1 = f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_fa412_y2 & f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_fa454_y2;
  assign f_s_dadda_rca24_u_rca_fa15_y2 = f_s_dadda_rca24_u_rca_fa15_y0 ^ f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_u_rca_fa14_y4;
  assign f_s_dadda_rca24_u_rca_fa15_y3 = f_s_dadda_rca24_u_rca_fa15_y0 & f_s_dadda_rca24_u_rca_fa15_f_s_dadda_rca24_u_rca_fa14_y4;
  assign f_s_dadda_rca24_u_rca_fa15_y4 = f_s_dadda_rca24_u_rca_fa15_y1 | f_s_dadda_rca24_u_rca_fa15_y3;
  assign f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_fa413_y2 = f_s_dadda_rca24_fa413_y2;
  assign f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_fa455_y2 = f_s_dadda_rca24_fa455_y2;
  assign f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_u_rca_fa15_y4 = f_s_dadda_rca24_u_rca_fa15_y4;
  assign f_s_dadda_rca24_u_rca_fa16_y0 = f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_fa413_y2 ^ f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_fa455_y2;
  assign f_s_dadda_rca24_u_rca_fa16_y1 = f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_fa413_y2 & f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_fa455_y2;
  assign f_s_dadda_rca24_u_rca_fa16_y2 = f_s_dadda_rca24_u_rca_fa16_y0 ^ f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_u_rca_fa15_y4;
  assign f_s_dadda_rca24_u_rca_fa16_y3 = f_s_dadda_rca24_u_rca_fa16_y0 & f_s_dadda_rca24_u_rca_fa16_f_s_dadda_rca24_u_rca_fa15_y4;
  assign f_s_dadda_rca24_u_rca_fa16_y4 = f_s_dadda_rca24_u_rca_fa16_y1 | f_s_dadda_rca24_u_rca_fa16_y3;
  assign f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_fa414_y2 = f_s_dadda_rca24_fa414_y2;
  assign f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_fa456_y2 = f_s_dadda_rca24_fa456_y2;
  assign f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_u_rca_fa16_y4 = f_s_dadda_rca24_u_rca_fa16_y4;
  assign f_s_dadda_rca24_u_rca_fa17_y0 = f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_fa414_y2 ^ f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_fa456_y2;
  assign f_s_dadda_rca24_u_rca_fa17_y1 = f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_fa414_y2 & f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_fa456_y2;
  assign f_s_dadda_rca24_u_rca_fa17_y2 = f_s_dadda_rca24_u_rca_fa17_y0 ^ f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_u_rca_fa16_y4;
  assign f_s_dadda_rca24_u_rca_fa17_y3 = f_s_dadda_rca24_u_rca_fa17_y0 & f_s_dadda_rca24_u_rca_fa17_f_s_dadda_rca24_u_rca_fa16_y4;
  assign f_s_dadda_rca24_u_rca_fa17_y4 = f_s_dadda_rca24_u_rca_fa17_y1 | f_s_dadda_rca24_u_rca_fa17_y3;
  assign f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_fa415_y2 = f_s_dadda_rca24_fa415_y2;
  assign f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_fa457_y2 = f_s_dadda_rca24_fa457_y2;
  assign f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_u_rca_fa17_y4 = f_s_dadda_rca24_u_rca_fa17_y4;
  assign f_s_dadda_rca24_u_rca_fa18_y0 = f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_fa415_y2 ^ f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_fa457_y2;
  assign f_s_dadda_rca24_u_rca_fa18_y1 = f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_fa415_y2 & f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_fa457_y2;
  assign f_s_dadda_rca24_u_rca_fa18_y2 = f_s_dadda_rca24_u_rca_fa18_y0 ^ f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_u_rca_fa17_y4;
  assign f_s_dadda_rca24_u_rca_fa18_y3 = f_s_dadda_rca24_u_rca_fa18_y0 & f_s_dadda_rca24_u_rca_fa18_f_s_dadda_rca24_u_rca_fa17_y4;
  assign f_s_dadda_rca24_u_rca_fa18_y4 = f_s_dadda_rca24_u_rca_fa18_y1 | f_s_dadda_rca24_u_rca_fa18_y3;
  assign f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_fa416_y2 = f_s_dadda_rca24_fa416_y2;
  assign f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_fa458_y2 = f_s_dadda_rca24_fa458_y2;
  assign f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_u_rca_fa18_y4 = f_s_dadda_rca24_u_rca_fa18_y4;
  assign f_s_dadda_rca24_u_rca_fa19_y0 = f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_fa416_y2 ^ f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_fa458_y2;
  assign f_s_dadda_rca24_u_rca_fa19_y1 = f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_fa416_y2 & f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_fa458_y2;
  assign f_s_dadda_rca24_u_rca_fa19_y2 = f_s_dadda_rca24_u_rca_fa19_y0 ^ f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_u_rca_fa18_y4;
  assign f_s_dadda_rca24_u_rca_fa19_y3 = f_s_dadda_rca24_u_rca_fa19_y0 & f_s_dadda_rca24_u_rca_fa19_f_s_dadda_rca24_u_rca_fa18_y4;
  assign f_s_dadda_rca24_u_rca_fa19_y4 = f_s_dadda_rca24_u_rca_fa19_y1 | f_s_dadda_rca24_u_rca_fa19_y3;
  assign f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_fa417_y2 = f_s_dadda_rca24_fa417_y2;
  assign f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_fa459_y2 = f_s_dadda_rca24_fa459_y2;
  assign f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_u_rca_fa19_y4 = f_s_dadda_rca24_u_rca_fa19_y4;
  assign f_s_dadda_rca24_u_rca_fa20_y0 = f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_fa417_y2 ^ f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_fa459_y2;
  assign f_s_dadda_rca24_u_rca_fa20_y1 = f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_fa417_y2 & f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_fa459_y2;
  assign f_s_dadda_rca24_u_rca_fa20_y2 = f_s_dadda_rca24_u_rca_fa20_y0 ^ f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_u_rca_fa19_y4;
  assign f_s_dadda_rca24_u_rca_fa20_y3 = f_s_dadda_rca24_u_rca_fa20_y0 & f_s_dadda_rca24_u_rca_fa20_f_s_dadda_rca24_u_rca_fa19_y4;
  assign f_s_dadda_rca24_u_rca_fa20_y4 = f_s_dadda_rca24_u_rca_fa20_y1 | f_s_dadda_rca24_u_rca_fa20_y3;
  assign f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_fa418_y2 = f_s_dadda_rca24_fa418_y2;
  assign f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_fa460_y2 = f_s_dadda_rca24_fa460_y2;
  assign f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_u_rca_fa20_y4 = f_s_dadda_rca24_u_rca_fa20_y4;
  assign f_s_dadda_rca24_u_rca_fa21_y0 = f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_fa418_y2 ^ f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_fa460_y2;
  assign f_s_dadda_rca24_u_rca_fa21_y1 = f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_fa418_y2 & f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_fa460_y2;
  assign f_s_dadda_rca24_u_rca_fa21_y2 = f_s_dadda_rca24_u_rca_fa21_y0 ^ f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_u_rca_fa20_y4;
  assign f_s_dadda_rca24_u_rca_fa21_y3 = f_s_dadda_rca24_u_rca_fa21_y0 & f_s_dadda_rca24_u_rca_fa21_f_s_dadda_rca24_u_rca_fa20_y4;
  assign f_s_dadda_rca24_u_rca_fa21_y4 = f_s_dadda_rca24_u_rca_fa21_y1 | f_s_dadda_rca24_u_rca_fa21_y3;
  assign f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_fa419_y2 = f_s_dadda_rca24_fa419_y2;
  assign f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_fa461_y2 = f_s_dadda_rca24_fa461_y2;
  assign f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_u_rca_fa21_y4 = f_s_dadda_rca24_u_rca_fa21_y4;
  assign f_s_dadda_rca24_u_rca_fa22_y0 = f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_fa419_y2 ^ f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_fa461_y2;
  assign f_s_dadda_rca24_u_rca_fa22_y1 = f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_fa419_y2 & f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_fa461_y2;
  assign f_s_dadda_rca24_u_rca_fa22_y2 = f_s_dadda_rca24_u_rca_fa22_y0 ^ f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_u_rca_fa21_y4;
  assign f_s_dadda_rca24_u_rca_fa22_y3 = f_s_dadda_rca24_u_rca_fa22_y0 & f_s_dadda_rca24_u_rca_fa22_f_s_dadda_rca24_u_rca_fa21_y4;
  assign f_s_dadda_rca24_u_rca_fa22_y4 = f_s_dadda_rca24_u_rca_fa22_y1 | f_s_dadda_rca24_u_rca_fa22_y3;
  assign f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_fa420_y2 = f_s_dadda_rca24_fa420_y2;
  assign f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_fa462_y2 = f_s_dadda_rca24_fa462_y2;
  assign f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_u_rca_fa22_y4 = f_s_dadda_rca24_u_rca_fa22_y4;
  assign f_s_dadda_rca24_u_rca_fa23_y0 = f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_fa420_y2 ^ f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_fa462_y2;
  assign f_s_dadda_rca24_u_rca_fa23_y1 = f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_fa420_y2 & f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_fa462_y2;
  assign f_s_dadda_rca24_u_rca_fa23_y2 = f_s_dadda_rca24_u_rca_fa23_y0 ^ f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_u_rca_fa22_y4;
  assign f_s_dadda_rca24_u_rca_fa23_y3 = f_s_dadda_rca24_u_rca_fa23_y0 & f_s_dadda_rca24_u_rca_fa23_f_s_dadda_rca24_u_rca_fa22_y4;
  assign f_s_dadda_rca24_u_rca_fa23_y4 = f_s_dadda_rca24_u_rca_fa23_y1 | f_s_dadda_rca24_u_rca_fa23_y3;
  assign f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_fa421_y2 = f_s_dadda_rca24_fa421_y2;
  assign f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_fa463_y2 = f_s_dadda_rca24_fa463_y2;
  assign f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_u_rca_fa23_y4 = f_s_dadda_rca24_u_rca_fa23_y4;
  assign f_s_dadda_rca24_u_rca_fa24_y0 = f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_fa421_y2 ^ f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_fa463_y2;
  assign f_s_dadda_rca24_u_rca_fa24_y1 = f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_fa421_y2 & f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_fa463_y2;
  assign f_s_dadda_rca24_u_rca_fa24_y2 = f_s_dadda_rca24_u_rca_fa24_y0 ^ f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_u_rca_fa23_y4;
  assign f_s_dadda_rca24_u_rca_fa24_y3 = f_s_dadda_rca24_u_rca_fa24_y0 & f_s_dadda_rca24_u_rca_fa24_f_s_dadda_rca24_u_rca_fa23_y4;
  assign f_s_dadda_rca24_u_rca_fa24_y4 = f_s_dadda_rca24_u_rca_fa24_y1 | f_s_dadda_rca24_u_rca_fa24_y3;
  assign f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_fa422_y2 = f_s_dadda_rca24_fa422_y2;
  assign f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_fa464_y2 = f_s_dadda_rca24_fa464_y2;
  assign f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_u_rca_fa24_y4 = f_s_dadda_rca24_u_rca_fa24_y4;
  assign f_s_dadda_rca24_u_rca_fa25_y0 = f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_fa422_y2 ^ f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_fa464_y2;
  assign f_s_dadda_rca24_u_rca_fa25_y1 = f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_fa422_y2 & f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_fa464_y2;
  assign f_s_dadda_rca24_u_rca_fa25_y2 = f_s_dadda_rca24_u_rca_fa25_y0 ^ f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_u_rca_fa24_y4;
  assign f_s_dadda_rca24_u_rca_fa25_y3 = f_s_dadda_rca24_u_rca_fa25_y0 & f_s_dadda_rca24_u_rca_fa25_f_s_dadda_rca24_u_rca_fa24_y4;
  assign f_s_dadda_rca24_u_rca_fa25_y4 = f_s_dadda_rca24_u_rca_fa25_y1 | f_s_dadda_rca24_u_rca_fa25_y3;
  assign f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_fa423_y2 = f_s_dadda_rca24_fa423_y2;
  assign f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_fa465_y2 = f_s_dadda_rca24_fa465_y2;
  assign f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_u_rca_fa25_y4 = f_s_dadda_rca24_u_rca_fa25_y4;
  assign f_s_dadda_rca24_u_rca_fa26_y0 = f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_fa423_y2 ^ f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_fa465_y2;
  assign f_s_dadda_rca24_u_rca_fa26_y1 = f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_fa423_y2 & f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_fa465_y2;
  assign f_s_dadda_rca24_u_rca_fa26_y2 = f_s_dadda_rca24_u_rca_fa26_y0 ^ f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_u_rca_fa25_y4;
  assign f_s_dadda_rca24_u_rca_fa26_y3 = f_s_dadda_rca24_u_rca_fa26_y0 & f_s_dadda_rca24_u_rca_fa26_f_s_dadda_rca24_u_rca_fa25_y4;
  assign f_s_dadda_rca24_u_rca_fa26_y4 = f_s_dadda_rca24_u_rca_fa26_y1 | f_s_dadda_rca24_u_rca_fa26_y3;
  assign f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_fa424_y2 = f_s_dadda_rca24_fa424_y2;
  assign f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_fa466_y2 = f_s_dadda_rca24_fa466_y2;
  assign f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_u_rca_fa26_y4 = f_s_dadda_rca24_u_rca_fa26_y4;
  assign f_s_dadda_rca24_u_rca_fa27_y0 = f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_fa424_y2 ^ f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_fa466_y2;
  assign f_s_dadda_rca24_u_rca_fa27_y1 = f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_fa424_y2 & f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_fa466_y2;
  assign f_s_dadda_rca24_u_rca_fa27_y2 = f_s_dadda_rca24_u_rca_fa27_y0 ^ f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_u_rca_fa26_y4;
  assign f_s_dadda_rca24_u_rca_fa27_y3 = f_s_dadda_rca24_u_rca_fa27_y0 & f_s_dadda_rca24_u_rca_fa27_f_s_dadda_rca24_u_rca_fa26_y4;
  assign f_s_dadda_rca24_u_rca_fa27_y4 = f_s_dadda_rca24_u_rca_fa27_y1 | f_s_dadda_rca24_u_rca_fa27_y3;
  assign f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_fa425_y2 = f_s_dadda_rca24_fa425_y2;
  assign f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_fa467_y2 = f_s_dadda_rca24_fa467_y2;
  assign f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_u_rca_fa27_y4 = f_s_dadda_rca24_u_rca_fa27_y4;
  assign f_s_dadda_rca24_u_rca_fa28_y0 = f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_fa425_y2 ^ f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_fa467_y2;
  assign f_s_dadda_rca24_u_rca_fa28_y1 = f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_fa425_y2 & f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_fa467_y2;
  assign f_s_dadda_rca24_u_rca_fa28_y2 = f_s_dadda_rca24_u_rca_fa28_y0 ^ f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_u_rca_fa27_y4;
  assign f_s_dadda_rca24_u_rca_fa28_y3 = f_s_dadda_rca24_u_rca_fa28_y0 & f_s_dadda_rca24_u_rca_fa28_f_s_dadda_rca24_u_rca_fa27_y4;
  assign f_s_dadda_rca24_u_rca_fa28_y4 = f_s_dadda_rca24_u_rca_fa28_y1 | f_s_dadda_rca24_u_rca_fa28_y3;
  assign f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_fa426_y2 = f_s_dadda_rca24_fa426_y2;
  assign f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_fa468_y2 = f_s_dadda_rca24_fa468_y2;
  assign f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_u_rca_fa28_y4 = f_s_dadda_rca24_u_rca_fa28_y4;
  assign f_s_dadda_rca24_u_rca_fa29_y0 = f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_fa426_y2 ^ f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_fa468_y2;
  assign f_s_dadda_rca24_u_rca_fa29_y1 = f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_fa426_y2 & f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_fa468_y2;
  assign f_s_dadda_rca24_u_rca_fa29_y2 = f_s_dadda_rca24_u_rca_fa29_y0 ^ f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_u_rca_fa28_y4;
  assign f_s_dadda_rca24_u_rca_fa29_y3 = f_s_dadda_rca24_u_rca_fa29_y0 & f_s_dadda_rca24_u_rca_fa29_f_s_dadda_rca24_u_rca_fa28_y4;
  assign f_s_dadda_rca24_u_rca_fa29_y4 = f_s_dadda_rca24_u_rca_fa29_y1 | f_s_dadda_rca24_u_rca_fa29_y3;
  assign f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_fa427_y2 = f_s_dadda_rca24_fa427_y2;
  assign f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_fa469_y2 = f_s_dadda_rca24_fa469_y2;
  assign f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_u_rca_fa29_y4 = f_s_dadda_rca24_u_rca_fa29_y4;
  assign f_s_dadda_rca24_u_rca_fa30_y0 = f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_fa427_y2 ^ f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_fa469_y2;
  assign f_s_dadda_rca24_u_rca_fa30_y1 = f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_fa427_y2 & f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_fa469_y2;
  assign f_s_dadda_rca24_u_rca_fa30_y2 = f_s_dadda_rca24_u_rca_fa30_y0 ^ f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_u_rca_fa29_y4;
  assign f_s_dadda_rca24_u_rca_fa30_y3 = f_s_dadda_rca24_u_rca_fa30_y0 & f_s_dadda_rca24_u_rca_fa30_f_s_dadda_rca24_u_rca_fa29_y4;
  assign f_s_dadda_rca24_u_rca_fa30_y4 = f_s_dadda_rca24_u_rca_fa30_y1 | f_s_dadda_rca24_u_rca_fa30_y3;
  assign f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_fa428_y2 = f_s_dadda_rca24_fa428_y2;
  assign f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_fa470_y2 = f_s_dadda_rca24_fa470_y2;
  assign f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_u_rca_fa30_y4 = f_s_dadda_rca24_u_rca_fa30_y4;
  assign f_s_dadda_rca24_u_rca_fa31_y0 = f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_fa428_y2 ^ f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_fa470_y2;
  assign f_s_dadda_rca24_u_rca_fa31_y1 = f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_fa428_y2 & f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_fa470_y2;
  assign f_s_dadda_rca24_u_rca_fa31_y2 = f_s_dadda_rca24_u_rca_fa31_y0 ^ f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_u_rca_fa30_y4;
  assign f_s_dadda_rca24_u_rca_fa31_y3 = f_s_dadda_rca24_u_rca_fa31_y0 & f_s_dadda_rca24_u_rca_fa31_f_s_dadda_rca24_u_rca_fa30_y4;
  assign f_s_dadda_rca24_u_rca_fa31_y4 = f_s_dadda_rca24_u_rca_fa31_y1 | f_s_dadda_rca24_u_rca_fa31_y3;
  assign f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_fa429_y2 = f_s_dadda_rca24_fa429_y2;
  assign f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_fa471_y2 = f_s_dadda_rca24_fa471_y2;
  assign f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_u_rca_fa31_y4 = f_s_dadda_rca24_u_rca_fa31_y4;
  assign f_s_dadda_rca24_u_rca_fa32_y0 = f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_fa429_y2 ^ f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_fa471_y2;
  assign f_s_dadda_rca24_u_rca_fa32_y1 = f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_fa429_y2 & f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_fa471_y2;
  assign f_s_dadda_rca24_u_rca_fa32_y2 = f_s_dadda_rca24_u_rca_fa32_y0 ^ f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_u_rca_fa31_y4;
  assign f_s_dadda_rca24_u_rca_fa32_y3 = f_s_dadda_rca24_u_rca_fa32_y0 & f_s_dadda_rca24_u_rca_fa32_f_s_dadda_rca24_u_rca_fa31_y4;
  assign f_s_dadda_rca24_u_rca_fa32_y4 = f_s_dadda_rca24_u_rca_fa32_y1 | f_s_dadda_rca24_u_rca_fa32_y3;
  assign f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_fa430_y2 = f_s_dadda_rca24_fa430_y2;
  assign f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_fa472_y2 = f_s_dadda_rca24_fa472_y2;
  assign f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_u_rca_fa32_y4 = f_s_dadda_rca24_u_rca_fa32_y4;
  assign f_s_dadda_rca24_u_rca_fa33_y0 = f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_fa430_y2 ^ f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_fa472_y2;
  assign f_s_dadda_rca24_u_rca_fa33_y1 = f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_fa430_y2 & f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_fa472_y2;
  assign f_s_dadda_rca24_u_rca_fa33_y2 = f_s_dadda_rca24_u_rca_fa33_y0 ^ f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_u_rca_fa32_y4;
  assign f_s_dadda_rca24_u_rca_fa33_y3 = f_s_dadda_rca24_u_rca_fa33_y0 & f_s_dadda_rca24_u_rca_fa33_f_s_dadda_rca24_u_rca_fa32_y4;
  assign f_s_dadda_rca24_u_rca_fa33_y4 = f_s_dadda_rca24_u_rca_fa33_y1 | f_s_dadda_rca24_u_rca_fa33_y3;
  assign f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_fa431_y2 = f_s_dadda_rca24_fa431_y2;
  assign f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_fa473_y2 = f_s_dadda_rca24_fa473_y2;
  assign f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_u_rca_fa33_y4 = f_s_dadda_rca24_u_rca_fa33_y4;
  assign f_s_dadda_rca24_u_rca_fa34_y0 = f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_fa431_y2 ^ f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_fa473_y2;
  assign f_s_dadda_rca24_u_rca_fa34_y1 = f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_fa431_y2 & f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_fa473_y2;
  assign f_s_dadda_rca24_u_rca_fa34_y2 = f_s_dadda_rca24_u_rca_fa34_y0 ^ f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_u_rca_fa33_y4;
  assign f_s_dadda_rca24_u_rca_fa34_y3 = f_s_dadda_rca24_u_rca_fa34_y0 & f_s_dadda_rca24_u_rca_fa34_f_s_dadda_rca24_u_rca_fa33_y4;
  assign f_s_dadda_rca24_u_rca_fa34_y4 = f_s_dadda_rca24_u_rca_fa34_y1 | f_s_dadda_rca24_u_rca_fa34_y3;
  assign f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_fa432_y2 = f_s_dadda_rca24_fa432_y2;
  assign f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_fa474_y2 = f_s_dadda_rca24_fa474_y2;
  assign f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_u_rca_fa34_y4 = f_s_dadda_rca24_u_rca_fa34_y4;
  assign f_s_dadda_rca24_u_rca_fa35_y0 = f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_fa432_y2 ^ f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_fa474_y2;
  assign f_s_dadda_rca24_u_rca_fa35_y1 = f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_fa432_y2 & f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_fa474_y2;
  assign f_s_dadda_rca24_u_rca_fa35_y2 = f_s_dadda_rca24_u_rca_fa35_y0 ^ f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_u_rca_fa34_y4;
  assign f_s_dadda_rca24_u_rca_fa35_y3 = f_s_dadda_rca24_u_rca_fa35_y0 & f_s_dadda_rca24_u_rca_fa35_f_s_dadda_rca24_u_rca_fa34_y4;
  assign f_s_dadda_rca24_u_rca_fa35_y4 = f_s_dadda_rca24_u_rca_fa35_y1 | f_s_dadda_rca24_u_rca_fa35_y3;
  assign f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_fa433_y2 = f_s_dadda_rca24_fa433_y2;
  assign f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_fa475_y2 = f_s_dadda_rca24_fa475_y2;
  assign f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_u_rca_fa35_y4 = f_s_dadda_rca24_u_rca_fa35_y4;
  assign f_s_dadda_rca24_u_rca_fa36_y0 = f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_fa433_y2 ^ f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_fa475_y2;
  assign f_s_dadda_rca24_u_rca_fa36_y1 = f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_fa433_y2 & f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_fa475_y2;
  assign f_s_dadda_rca24_u_rca_fa36_y2 = f_s_dadda_rca24_u_rca_fa36_y0 ^ f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_u_rca_fa35_y4;
  assign f_s_dadda_rca24_u_rca_fa36_y3 = f_s_dadda_rca24_u_rca_fa36_y0 & f_s_dadda_rca24_u_rca_fa36_f_s_dadda_rca24_u_rca_fa35_y4;
  assign f_s_dadda_rca24_u_rca_fa36_y4 = f_s_dadda_rca24_u_rca_fa36_y1 | f_s_dadda_rca24_u_rca_fa36_y3;
  assign f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_fa434_y2 = f_s_dadda_rca24_fa434_y2;
  assign f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_fa476_y2 = f_s_dadda_rca24_fa476_y2;
  assign f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_u_rca_fa36_y4 = f_s_dadda_rca24_u_rca_fa36_y4;
  assign f_s_dadda_rca24_u_rca_fa37_y0 = f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_fa434_y2 ^ f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_fa476_y2;
  assign f_s_dadda_rca24_u_rca_fa37_y1 = f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_fa434_y2 & f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_fa476_y2;
  assign f_s_dadda_rca24_u_rca_fa37_y2 = f_s_dadda_rca24_u_rca_fa37_y0 ^ f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_u_rca_fa36_y4;
  assign f_s_dadda_rca24_u_rca_fa37_y3 = f_s_dadda_rca24_u_rca_fa37_y0 & f_s_dadda_rca24_u_rca_fa37_f_s_dadda_rca24_u_rca_fa36_y4;
  assign f_s_dadda_rca24_u_rca_fa37_y4 = f_s_dadda_rca24_u_rca_fa37_y1 | f_s_dadda_rca24_u_rca_fa37_y3;
  assign f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_fa435_y2 = f_s_dadda_rca24_fa435_y2;
  assign f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_fa477_y2 = f_s_dadda_rca24_fa477_y2;
  assign f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_u_rca_fa37_y4 = f_s_dadda_rca24_u_rca_fa37_y4;
  assign f_s_dadda_rca24_u_rca_fa38_y0 = f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_fa435_y2 ^ f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_fa477_y2;
  assign f_s_dadda_rca24_u_rca_fa38_y1 = f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_fa435_y2 & f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_fa477_y2;
  assign f_s_dadda_rca24_u_rca_fa38_y2 = f_s_dadda_rca24_u_rca_fa38_y0 ^ f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_u_rca_fa37_y4;
  assign f_s_dadda_rca24_u_rca_fa38_y3 = f_s_dadda_rca24_u_rca_fa38_y0 & f_s_dadda_rca24_u_rca_fa38_f_s_dadda_rca24_u_rca_fa37_y4;
  assign f_s_dadda_rca24_u_rca_fa38_y4 = f_s_dadda_rca24_u_rca_fa38_y1 | f_s_dadda_rca24_u_rca_fa38_y3;
  assign f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_fa436_y2 = f_s_dadda_rca24_fa436_y2;
  assign f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_fa478_y2 = f_s_dadda_rca24_fa478_y2;
  assign f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_u_rca_fa38_y4 = f_s_dadda_rca24_u_rca_fa38_y4;
  assign f_s_dadda_rca24_u_rca_fa39_y0 = f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_fa436_y2 ^ f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_fa478_y2;
  assign f_s_dadda_rca24_u_rca_fa39_y1 = f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_fa436_y2 & f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_fa478_y2;
  assign f_s_dadda_rca24_u_rca_fa39_y2 = f_s_dadda_rca24_u_rca_fa39_y0 ^ f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_u_rca_fa38_y4;
  assign f_s_dadda_rca24_u_rca_fa39_y3 = f_s_dadda_rca24_u_rca_fa39_y0 & f_s_dadda_rca24_u_rca_fa39_f_s_dadda_rca24_u_rca_fa38_y4;
  assign f_s_dadda_rca24_u_rca_fa39_y4 = f_s_dadda_rca24_u_rca_fa39_y1 | f_s_dadda_rca24_u_rca_fa39_y3;
  assign f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_fa437_y2 = f_s_dadda_rca24_fa437_y2;
  assign f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_fa479_y2 = f_s_dadda_rca24_fa479_y2;
  assign f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_u_rca_fa39_y4 = f_s_dadda_rca24_u_rca_fa39_y4;
  assign f_s_dadda_rca24_u_rca_fa40_y0 = f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_fa437_y2 ^ f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_fa479_y2;
  assign f_s_dadda_rca24_u_rca_fa40_y1 = f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_fa437_y2 & f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_fa479_y2;
  assign f_s_dadda_rca24_u_rca_fa40_y2 = f_s_dadda_rca24_u_rca_fa40_y0 ^ f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_u_rca_fa39_y4;
  assign f_s_dadda_rca24_u_rca_fa40_y3 = f_s_dadda_rca24_u_rca_fa40_y0 & f_s_dadda_rca24_u_rca_fa40_f_s_dadda_rca24_u_rca_fa39_y4;
  assign f_s_dadda_rca24_u_rca_fa40_y4 = f_s_dadda_rca24_u_rca_fa40_y1 | f_s_dadda_rca24_u_rca_fa40_y3;
  assign f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_fa438_y2 = f_s_dadda_rca24_fa438_y2;
  assign f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_fa480_y2 = f_s_dadda_rca24_fa480_y2;
  assign f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_u_rca_fa40_y4 = f_s_dadda_rca24_u_rca_fa40_y4;
  assign f_s_dadda_rca24_u_rca_fa41_y0 = f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_fa438_y2 ^ f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_fa480_y2;
  assign f_s_dadda_rca24_u_rca_fa41_y1 = f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_fa438_y2 & f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_fa480_y2;
  assign f_s_dadda_rca24_u_rca_fa41_y2 = f_s_dadda_rca24_u_rca_fa41_y0 ^ f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_u_rca_fa40_y4;
  assign f_s_dadda_rca24_u_rca_fa41_y3 = f_s_dadda_rca24_u_rca_fa41_y0 & f_s_dadda_rca24_u_rca_fa41_f_s_dadda_rca24_u_rca_fa40_y4;
  assign f_s_dadda_rca24_u_rca_fa41_y4 = f_s_dadda_rca24_u_rca_fa41_y1 | f_s_dadda_rca24_u_rca_fa41_y3;
  assign f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_fa439_y2 = f_s_dadda_rca24_fa439_y2;
  assign f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_fa481_y2 = f_s_dadda_rca24_fa481_y2;
  assign f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_u_rca_fa41_y4 = f_s_dadda_rca24_u_rca_fa41_y4;
  assign f_s_dadda_rca24_u_rca_fa42_y0 = f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_fa439_y2 ^ f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_fa481_y2;
  assign f_s_dadda_rca24_u_rca_fa42_y1 = f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_fa439_y2 & f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_fa481_y2;
  assign f_s_dadda_rca24_u_rca_fa42_y2 = f_s_dadda_rca24_u_rca_fa42_y0 ^ f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_u_rca_fa41_y4;
  assign f_s_dadda_rca24_u_rca_fa42_y3 = f_s_dadda_rca24_u_rca_fa42_y0 & f_s_dadda_rca24_u_rca_fa42_f_s_dadda_rca24_u_rca_fa41_y4;
  assign f_s_dadda_rca24_u_rca_fa42_y4 = f_s_dadda_rca24_u_rca_fa42_y1 | f_s_dadda_rca24_u_rca_fa42_y3;
  assign f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_fa440_y2 = f_s_dadda_rca24_fa440_y2;
  assign f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_fa482_y2 = f_s_dadda_rca24_fa482_y2;
  assign f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_u_rca_fa42_y4 = f_s_dadda_rca24_u_rca_fa42_y4;
  assign f_s_dadda_rca24_u_rca_fa43_y0 = f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_fa440_y2 ^ f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_fa482_y2;
  assign f_s_dadda_rca24_u_rca_fa43_y1 = f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_fa440_y2 & f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_fa482_y2;
  assign f_s_dadda_rca24_u_rca_fa43_y2 = f_s_dadda_rca24_u_rca_fa43_y0 ^ f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_u_rca_fa42_y4;
  assign f_s_dadda_rca24_u_rca_fa43_y3 = f_s_dadda_rca24_u_rca_fa43_y0 & f_s_dadda_rca24_u_rca_fa43_f_s_dadda_rca24_u_rca_fa42_y4;
  assign f_s_dadda_rca24_u_rca_fa43_y4 = f_s_dadda_rca24_u_rca_fa43_y1 | f_s_dadda_rca24_u_rca_fa43_y3;
  assign f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_nand_22_23_y0 = f_s_dadda_rca24_nand_22_23_y0;
  assign f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_fa483_y2 = f_s_dadda_rca24_fa483_y2;
  assign f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_u_rca_fa43_y4 = f_s_dadda_rca24_u_rca_fa43_y4;
  assign f_s_dadda_rca24_u_rca_fa44_y0 = f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_nand_22_23_y0 ^ f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_fa483_y2;
  assign f_s_dadda_rca24_u_rca_fa44_y1 = f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_nand_22_23_y0 & f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_fa483_y2;
  assign f_s_dadda_rca24_u_rca_fa44_y2 = f_s_dadda_rca24_u_rca_fa44_y0 ^ f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_u_rca_fa43_y4;
  assign f_s_dadda_rca24_u_rca_fa44_y3 = f_s_dadda_rca24_u_rca_fa44_y0 & f_s_dadda_rca24_u_rca_fa44_f_s_dadda_rca24_u_rca_fa43_y4;
  assign f_s_dadda_rca24_u_rca_fa44_y4 = f_s_dadda_rca24_u_rca_fa44_y1 | f_s_dadda_rca24_u_rca_fa44_y3;
  assign f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_fa483_y4 = f_s_dadda_rca24_fa483_y4;
  assign f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_and_23_23_y0 = f_s_dadda_rca24_and_23_23_y0;
  assign f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_u_rca_fa44_y4 = f_s_dadda_rca24_u_rca_fa44_y4;
  assign f_s_dadda_rca24_u_rca_fa45_y0 = f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_fa483_y4 ^ f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_and_23_23_y0;
  assign f_s_dadda_rca24_u_rca_fa45_y1 = f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_fa483_y4 & f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_and_23_23_y0;
  assign f_s_dadda_rca24_u_rca_fa45_y2 = f_s_dadda_rca24_u_rca_fa45_y0 ^ f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_u_rca_fa44_y4;
  assign f_s_dadda_rca24_u_rca_fa45_y3 = f_s_dadda_rca24_u_rca_fa45_y0 & f_s_dadda_rca24_u_rca_fa45_f_s_dadda_rca24_u_rca_fa44_y4;
  assign f_s_dadda_rca24_u_rca_fa45_y4 = f_s_dadda_rca24_u_rca_fa45_y1 | f_s_dadda_rca24_u_rca_fa45_y3;
  assign f_s_dadda_rca24_xor0_constant_wire_1 = constant_wire_1;
  assign f_s_dadda_rca24_xor0_f_s_dadda_rca24_u_rca_fa45_y4 = f_s_dadda_rca24_u_rca_fa45_y4;
  assign f_s_dadda_rca24_xor0_y0 = f_s_dadda_rca24_xor0_constant_wire_1 ^ f_s_dadda_rca24_xor0_f_s_dadda_rca24_u_rca_fa45_y4;

  assign out[0] = f_s_dadda_rca24_and_0_0_y0;
  assign out[1] = f_s_dadda_rca24_u_rca_ha_y0;
  assign out[2] = f_s_dadda_rca24_u_rca_fa1_y2;
  assign out[3] = f_s_dadda_rca24_u_rca_fa2_y2;
  assign out[4] = f_s_dadda_rca24_u_rca_fa3_y2;
  assign out[5] = f_s_dadda_rca24_u_rca_fa4_y2;
  assign out[6] = f_s_dadda_rca24_u_rca_fa5_y2;
  assign out[7] = f_s_dadda_rca24_u_rca_fa6_y2;
  assign out[8] = f_s_dadda_rca24_u_rca_fa7_y2;
  assign out[9] = f_s_dadda_rca24_u_rca_fa8_y2;
  assign out[10] = f_s_dadda_rca24_u_rca_fa9_y2;
  assign out[11] = f_s_dadda_rca24_u_rca_fa10_y2;
  assign out[12] = f_s_dadda_rca24_u_rca_fa11_y2;
  assign out[13] = f_s_dadda_rca24_u_rca_fa12_y2;
  assign out[14] = f_s_dadda_rca24_u_rca_fa13_y2;
  assign out[15] = f_s_dadda_rca24_u_rca_fa14_y2;
  assign out[16] = f_s_dadda_rca24_u_rca_fa15_y2;
  assign out[17] = f_s_dadda_rca24_u_rca_fa16_y2;
  assign out[18] = f_s_dadda_rca24_u_rca_fa17_y2;
  assign out[19] = f_s_dadda_rca24_u_rca_fa18_y2;
  assign out[20] = f_s_dadda_rca24_u_rca_fa19_y2;
  assign out[21] = f_s_dadda_rca24_u_rca_fa20_y2;
  assign out[22] = f_s_dadda_rca24_u_rca_fa21_y2;
  assign out[23] = f_s_dadda_rca24_u_rca_fa22_y2;
  assign out[24] = f_s_dadda_rca24_u_rca_fa23_y2;
  assign out[25] = f_s_dadda_rca24_u_rca_fa24_y2;
  assign out[26] = f_s_dadda_rca24_u_rca_fa25_y2;
  assign out[27] = f_s_dadda_rca24_u_rca_fa26_y2;
  assign out[28] = f_s_dadda_rca24_u_rca_fa27_y2;
  assign out[29] = f_s_dadda_rca24_u_rca_fa28_y2;
  assign out[30] = f_s_dadda_rca24_u_rca_fa29_y2;
  assign out[31] = f_s_dadda_rca24_u_rca_fa30_y2;
  assign out[32] = f_s_dadda_rca24_u_rca_fa31_y2;
  assign out[33] = f_s_dadda_rca24_u_rca_fa32_y2;
  assign out[34] = f_s_dadda_rca24_u_rca_fa33_y2;
  assign out[35] = f_s_dadda_rca24_u_rca_fa34_y2;
  assign out[36] = f_s_dadda_rca24_u_rca_fa35_y2;
  assign out[37] = f_s_dadda_rca24_u_rca_fa36_y2;
  assign out[38] = f_s_dadda_rca24_u_rca_fa37_y2;
  assign out[39] = f_s_dadda_rca24_u_rca_fa38_y2;
  assign out[40] = f_s_dadda_rca24_u_rca_fa39_y2;
  assign out[41] = f_s_dadda_rca24_u_rca_fa40_y2;
  assign out[42] = f_s_dadda_rca24_u_rca_fa41_y2;
  assign out[43] = f_s_dadda_rca24_u_rca_fa42_y2;
  assign out[44] = f_s_dadda_rca24_u_rca_fa43_y2;
  assign out[45] = f_s_dadda_rca24_u_rca_fa44_y2;
  assign out[46] = f_s_dadda_rca24_u_rca_fa45_y2;
  assign out[47] = f_s_dadda_rca24_xor0_y0;
endmodule