module xor_gate(input _a, input _b, output _y0);
  assign _y0 = _a ^ _b;
endmodule

module xnor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a ^ _b);
endmodule

module nor_gate(input _a, input _b, output _y0);
  assign _y0 = ~(_a | _b);
endmodule

module or_gate(input _a, input _b, output _y0);
  assign _y0 = _a | _b;
endmodule

module and_gate(input _a, input _b, output _y0);
  assign _y0 = _a & _b;
endmodule

module constant_wire_value_0(input a, input b, output constant_wire_0);
  wire constant_wire_value_0_a;
  wire constant_wire_value_0_b;

  assign constant_wire_value_0_a = a;
  assign constant_wire_value_0_b = b;

  xor_gate xor_gate_constant_wire_value_0_y0(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y0);
  xnor_gate xnor_gate_constant_wire_value_0_y1(constant_wire_value_0_a, constant_wire_value_0_b, constant_wire_value_0_y1);
  nor_gate nor_gate_constant_wire_0(constant_wire_value_0_y0, constant_wire_value_0_y1, constant_wire_0);
endmodule

module pg_logic(input a, input b, output pg_logic_y0, output pg_logic_y1, output pg_logic_y2);
  wire pg_logic_a;
  wire pg_logic_b;

  assign pg_logic_a = a;
  assign pg_logic_b = b;

  or_gate or_gate_pg_logic_y0(pg_logic_a, pg_logic_b, pg_logic_y0);
  and_gate and_gate_pg_logic_y1(pg_logic_a, pg_logic_b, pg_logic_y1);
  xor_gate xor_gate_pg_logic_y2(pg_logic_a, pg_logic_b, pg_logic_y2);
endmodule

module h_s_cla16(input [15:0] a, input [15:0] b, output [16:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire constant_wire_0;
  wire h_s_cla16_pg_logic0_y0;
  wire h_s_cla16_pg_logic0_y1;
  wire h_s_cla16_pg_logic0_y2;
  wire h_s_cla16_xor0_y0;
  wire h_s_cla16_and0_y0;
  wire h_s_cla16_or0_y0;
  wire h_s_cla16_pg_logic1_y0;
  wire h_s_cla16_pg_logic1_y1;
  wire h_s_cla16_pg_logic1_y2;
  wire h_s_cla16_xor1_y0;
  wire h_s_cla16_and1_y0;
  wire h_s_cla16_and2_y0;
  wire h_s_cla16_and3_y0;
  wire h_s_cla16_and4_y0;
  wire h_s_cla16_or1_y0;
  wire h_s_cla16_or2_y0;
  wire h_s_cla16_pg_logic2_y0;
  wire h_s_cla16_pg_logic2_y1;
  wire h_s_cla16_pg_logic2_y2;
  wire h_s_cla16_xor2_y0;
  wire h_s_cla16_and5_y0;
  wire h_s_cla16_and6_y0;
  wire h_s_cla16_and7_y0;
  wire h_s_cla16_and8_y0;
  wire h_s_cla16_and9_y0;
  wire h_s_cla16_and10_y0;
  wire h_s_cla16_and11_y0;
  wire h_s_cla16_and12_y0;
  wire h_s_cla16_and13_y0;
  wire h_s_cla16_or3_y0;
  wire h_s_cla16_or4_y0;
  wire h_s_cla16_or5_y0;
  wire h_s_cla16_pg_logic3_y0;
  wire h_s_cla16_pg_logic3_y1;
  wire h_s_cla16_pg_logic3_y2;
  wire h_s_cla16_xor3_y0;
  wire h_s_cla16_and14_y0;
  wire h_s_cla16_and15_y0;
  wire h_s_cla16_and16_y0;
  wire h_s_cla16_and17_y0;
  wire h_s_cla16_and18_y0;
  wire h_s_cla16_and19_y0;
  wire h_s_cla16_and20_y0;
  wire h_s_cla16_and21_y0;
  wire h_s_cla16_and22_y0;
  wire h_s_cla16_and23_y0;
  wire h_s_cla16_and24_y0;
  wire h_s_cla16_and25_y0;
  wire h_s_cla16_and26_y0;
  wire h_s_cla16_and27_y0;
  wire h_s_cla16_and28_y0;
  wire h_s_cla16_and29_y0;
  wire h_s_cla16_or6_y0;
  wire h_s_cla16_or7_y0;
  wire h_s_cla16_or8_y0;
  wire h_s_cla16_or9_y0;
  wire h_s_cla16_pg_logic4_y0;
  wire h_s_cla16_pg_logic4_y1;
  wire h_s_cla16_pg_logic4_y2;
  wire h_s_cla16_xor4_y0;
  wire h_s_cla16_and30_y0;
  wire h_s_cla16_and31_y0;
  wire h_s_cla16_and32_y0;
  wire h_s_cla16_and33_y0;
  wire h_s_cla16_and34_y0;
  wire h_s_cla16_and35_y0;
  wire h_s_cla16_and36_y0;
  wire h_s_cla16_and37_y0;
  wire h_s_cla16_and38_y0;
  wire h_s_cla16_and39_y0;
  wire h_s_cla16_and40_y0;
  wire h_s_cla16_and41_y0;
  wire h_s_cla16_and42_y0;
  wire h_s_cla16_and43_y0;
  wire h_s_cla16_and44_y0;
  wire h_s_cla16_and45_y0;
  wire h_s_cla16_and46_y0;
  wire h_s_cla16_and47_y0;
  wire h_s_cla16_and48_y0;
  wire h_s_cla16_and49_y0;
  wire h_s_cla16_and50_y0;
  wire h_s_cla16_and51_y0;
  wire h_s_cla16_and52_y0;
  wire h_s_cla16_and53_y0;
  wire h_s_cla16_and54_y0;
  wire h_s_cla16_or10_y0;
  wire h_s_cla16_or11_y0;
  wire h_s_cla16_or12_y0;
  wire h_s_cla16_or13_y0;
  wire h_s_cla16_or14_y0;
  wire h_s_cla16_pg_logic5_y0;
  wire h_s_cla16_pg_logic5_y1;
  wire h_s_cla16_pg_logic5_y2;
  wire h_s_cla16_xor5_y0;
  wire h_s_cla16_and55_y0;
  wire h_s_cla16_and56_y0;
  wire h_s_cla16_and57_y0;
  wire h_s_cla16_and58_y0;
  wire h_s_cla16_and59_y0;
  wire h_s_cla16_and60_y0;
  wire h_s_cla16_and61_y0;
  wire h_s_cla16_and62_y0;
  wire h_s_cla16_and63_y0;
  wire h_s_cla16_and64_y0;
  wire h_s_cla16_and65_y0;
  wire h_s_cla16_and66_y0;
  wire h_s_cla16_and67_y0;
  wire h_s_cla16_and68_y0;
  wire h_s_cla16_and69_y0;
  wire h_s_cla16_and70_y0;
  wire h_s_cla16_and71_y0;
  wire h_s_cla16_and72_y0;
  wire h_s_cla16_and73_y0;
  wire h_s_cla16_and74_y0;
  wire h_s_cla16_and75_y0;
  wire h_s_cla16_and76_y0;
  wire h_s_cla16_and77_y0;
  wire h_s_cla16_and78_y0;
  wire h_s_cla16_and79_y0;
  wire h_s_cla16_and80_y0;
  wire h_s_cla16_and81_y0;
  wire h_s_cla16_and82_y0;
  wire h_s_cla16_and83_y0;
  wire h_s_cla16_and84_y0;
  wire h_s_cla16_and85_y0;
  wire h_s_cla16_and86_y0;
  wire h_s_cla16_and87_y0;
  wire h_s_cla16_and88_y0;
  wire h_s_cla16_and89_y0;
  wire h_s_cla16_and90_y0;
  wire h_s_cla16_or15_y0;
  wire h_s_cla16_or16_y0;
  wire h_s_cla16_or17_y0;
  wire h_s_cla16_or18_y0;
  wire h_s_cla16_or19_y0;
  wire h_s_cla16_or20_y0;
  wire h_s_cla16_pg_logic6_y0;
  wire h_s_cla16_pg_logic6_y1;
  wire h_s_cla16_pg_logic6_y2;
  wire h_s_cla16_xor6_y0;
  wire h_s_cla16_and91_y0;
  wire h_s_cla16_and92_y0;
  wire h_s_cla16_and93_y0;
  wire h_s_cla16_and94_y0;
  wire h_s_cla16_and95_y0;
  wire h_s_cla16_and96_y0;
  wire h_s_cla16_and97_y0;
  wire h_s_cla16_and98_y0;
  wire h_s_cla16_and99_y0;
  wire h_s_cla16_and100_y0;
  wire h_s_cla16_and101_y0;
  wire h_s_cla16_and102_y0;
  wire h_s_cla16_and103_y0;
  wire h_s_cla16_and104_y0;
  wire h_s_cla16_and105_y0;
  wire h_s_cla16_and106_y0;
  wire h_s_cla16_and107_y0;
  wire h_s_cla16_and108_y0;
  wire h_s_cla16_and109_y0;
  wire h_s_cla16_and110_y0;
  wire h_s_cla16_and111_y0;
  wire h_s_cla16_and112_y0;
  wire h_s_cla16_and113_y0;
  wire h_s_cla16_and114_y0;
  wire h_s_cla16_and115_y0;
  wire h_s_cla16_and116_y0;
  wire h_s_cla16_and117_y0;
  wire h_s_cla16_and118_y0;
  wire h_s_cla16_and119_y0;
  wire h_s_cla16_and120_y0;
  wire h_s_cla16_and121_y0;
  wire h_s_cla16_and122_y0;
  wire h_s_cla16_and123_y0;
  wire h_s_cla16_and124_y0;
  wire h_s_cla16_and125_y0;
  wire h_s_cla16_and126_y0;
  wire h_s_cla16_and127_y0;
  wire h_s_cla16_and128_y0;
  wire h_s_cla16_and129_y0;
  wire h_s_cla16_and130_y0;
  wire h_s_cla16_and131_y0;
  wire h_s_cla16_and132_y0;
  wire h_s_cla16_and133_y0;
  wire h_s_cla16_and134_y0;
  wire h_s_cla16_and135_y0;
  wire h_s_cla16_and136_y0;
  wire h_s_cla16_and137_y0;
  wire h_s_cla16_and138_y0;
  wire h_s_cla16_and139_y0;
  wire h_s_cla16_or21_y0;
  wire h_s_cla16_or22_y0;
  wire h_s_cla16_or23_y0;
  wire h_s_cla16_or24_y0;
  wire h_s_cla16_or25_y0;
  wire h_s_cla16_or26_y0;
  wire h_s_cla16_or27_y0;
  wire h_s_cla16_pg_logic7_y0;
  wire h_s_cla16_pg_logic7_y1;
  wire h_s_cla16_pg_logic7_y2;
  wire h_s_cla16_xor7_y0;
  wire h_s_cla16_and140_y0;
  wire h_s_cla16_and141_y0;
  wire h_s_cla16_and142_y0;
  wire h_s_cla16_and143_y0;
  wire h_s_cla16_and144_y0;
  wire h_s_cla16_and145_y0;
  wire h_s_cla16_and146_y0;
  wire h_s_cla16_and147_y0;
  wire h_s_cla16_and148_y0;
  wire h_s_cla16_and149_y0;
  wire h_s_cla16_and150_y0;
  wire h_s_cla16_and151_y0;
  wire h_s_cla16_and152_y0;
  wire h_s_cla16_and153_y0;
  wire h_s_cla16_and154_y0;
  wire h_s_cla16_and155_y0;
  wire h_s_cla16_and156_y0;
  wire h_s_cla16_and157_y0;
  wire h_s_cla16_and158_y0;
  wire h_s_cla16_and159_y0;
  wire h_s_cla16_and160_y0;
  wire h_s_cla16_and161_y0;
  wire h_s_cla16_and162_y0;
  wire h_s_cla16_and163_y0;
  wire h_s_cla16_and164_y0;
  wire h_s_cla16_and165_y0;
  wire h_s_cla16_and166_y0;
  wire h_s_cla16_and167_y0;
  wire h_s_cla16_and168_y0;
  wire h_s_cla16_and169_y0;
  wire h_s_cla16_and170_y0;
  wire h_s_cla16_and171_y0;
  wire h_s_cla16_and172_y0;
  wire h_s_cla16_and173_y0;
  wire h_s_cla16_and174_y0;
  wire h_s_cla16_and175_y0;
  wire h_s_cla16_and176_y0;
  wire h_s_cla16_and177_y0;
  wire h_s_cla16_and178_y0;
  wire h_s_cla16_and179_y0;
  wire h_s_cla16_and180_y0;
  wire h_s_cla16_and181_y0;
  wire h_s_cla16_and182_y0;
  wire h_s_cla16_and183_y0;
  wire h_s_cla16_and184_y0;
  wire h_s_cla16_and185_y0;
  wire h_s_cla16_and186_y0;
  wire h_s_cla16_and187_y0;
  wire h_s_cla16_and188_y0;
  wire h_s_cla16_and189_y0;
  wire h_s_cla16_and190_y0;
  wire h_s_cla16_and191_y0;
  wire h_s_cla16_and192_y0;
  wire h_s_cla16_and193_y0;
  wire h_s_cla16_and194_y0;
  wire h_s_cla16_and195_y0;
  wire h_s_cla16_and196_y0;
  wire h_s_cla16_and197_y0;
  wire h_s_cla16_and198_y0;
  wire h_s_cla16_and199_y0;
  wire h_s_cla16_and200_y0;
  wire h_s_cla16_and201_y0;
  wire h_s_cla16_and202_y0;
  wire h_s_cla16_and203_y0;
  wire h_s_cla16_or28_y0;
  wire h_s_cla16_or29_y0;
  wire h_s_cla16_or30_y0;
  wire h_s_cla16_or31_y0;
  wire h_s_cla16_or32_y0;
  wire h_s_cla16_or33_y0;
  wire h_s_cla16_or34_y0;
  wire h_s_cla16_or35_y0;
  wire h_s_cla16_pg_logic8_y0;
  wire h_s_cla16_pg_logic8_y1;
  wire h_s_cla16_pg_logic8_y2;
  wire h_s_cla16_xor8_y0;
  wire h_s_cla16_and204_y0;
  wire h_s_cla16_and205_y0;
  wire h_s_cla16_and206_y0;
  wire h_s_cla16_and207_y0;
  wire h_s_cla16_and208_y0;
  wire h_s_cla16_and209_y0;
  wire h_s_cla16_and210_y0;
  wire h_s_cla16_and211_y0;
  wire h_s_cla16_and212_y0;
  wire h_s_cla16_and213_y0;
  wire h_s_cla16_and214_y0;
  wire h_s_cla16_and215_y0;
  wire h_s_cla16_and216_y0;
  wire h_s_cla16_and217_y0;
  wire h_s_cla16_and218_y0;
  wire h_s_cla16_and219_y0;
  wire h_s_cla16_and220_y0;
  wire h_s_cla16_and221_y0;
  wire h_s_cla16_and222_y0;
  wire h_s_cla16_and223_y0;
  wire h_s_cla16_and224_y0;
  wire h_s_cla16_and225_y0;
  wire h_s_cla16_and226_y0;
  wire h_s_cla16_and227_y0;
  wire h_s_cla16_and228_y0;
  wire h_s_cla16_and229_y0;
  wire h_s_cla16_and230_y0;
  wire h_s_cla16_and231_y0;
  wire h_s_cla16_and232_y0;
  wire h_s_cla16_and233_y0;
  wire h_s_cla16_and234_y0;
  wire h_s_cla16_and235_y0;
  wire h_s_cla16_and236_y0;
  wire h_s_cla16_and237_y0;
  wire h_s_cla16_and238_y0;
  wire h_s_cla16_and239_y0;
  wire h_s_cla16_and240_y0;
  wire h_s_cla16_and241_y0;
  wire h_s_cla16_and242_y0;
  wire h_s_cla16_and243_y0;
  wire h_s_cla16_and244_y0;
  wire h_s_cla16_and245_y0;
  wire h_s_cla16_and246_y0;
  wire h_s_cla16_and247_y0;
  wire h_s_cla16_and248_y0;
  wire h_s_cla16_and249_y0;
  wire h_s_cla16_and250_y0;
  wire h_s_cla16_and251_y0;
  wire h_s_cla16_and252_y0;
  wire h_s_cla16_and253_y0;
  wire h_s_cla16_and254_y0;
  wire h_s_cla16_and255_y0;
  wire h_s_cla16_and256_y0;
  wire h_s_cla16_and257_y0;
  wire h_s_cla16_and258_y0;
  wire h_s_cla16_and259_y0;
  wire h_s_cla16_and260_y0;
  wire h_s_cla16_and261_y0;
  wire h_s_cla16_and262_y0;
  wire h_s_cla16_and263_y0;
  wire h_s_cla16_and264_y0;
  wire h_s_cla16_and265_y0;
  wire h_s_cla16_and266_y0;
  wire h_s_cla16_and267_y0;
  wire h_s_cla16_and268_y0;
  wire h_s_cla16_and269_y0;
  wire h_s_cla16_and270_y0;
  wire h_s_cla16_and271_y0;
  wire h_s_cla16_and272_y0;
  wire h_s_cla16_and273_y0;
  wire h_s_cla16_and274_y0;
  wire h_s_cla16_and275_y0;
  wire h_s_cla16_and276_y0;
  wire h_s_cla16_and277_y0;
  wire h_s_cla16_and278_y0;
  wire h_s_cla16_and279_y0;
  wire h_s_cla16_and280_y0;
  wire h_s_cla16_and281_y0;
  wire h_s_cla16_and282_y0;
  wire h_s_cla16_and283_y0;
  wire h_s_cla16_and284_y0;
  wire h_s_cla16_or36_y0;
  wire h_s_cla16_or37_y0;
  wire h_s_cla16_or38_y0;
  wire h_s_cla16_or39_y0;
  wire h_s_cla16_or40_y0;
  wire h_s_cla16_or41_y0;
  wire h_s_cla16_or42_y0;
  wire h_s_cla16_or43_y0;
  wire h_s_cla16_or44_y0;
  wire h_s_cla16_pg_logic9_y0;
  wire h_s_cla16_pg_logic9_y1;
  wire h_s_cla16_pg_logic9_y2;
  wire h_s_cla16_xor9_y0;
  wire h_s_cla16_and285_y0;
  wire h_s_cla16_and286_y0;
  wire h_s_cla16_and287_y0;
  wire h_s_cla16_and288_y0;
  wire h_s_cla16_and289_y0;
  wire h_s_cla16_and290_y0;
  wire h_s_cla16_and291_y0;
  wire h_s_cla16_and292_y0;
  wire h_s_cla16_and293_y0;
  wire h_s_cla16_and294_y0;
  wire h_s_cla16_and295_y0;
  wire h_s_cla16_and296_y0;
  wire h_s_cla16_and297_y0;
  wire h_s_cla16_and298_y0;
  wire h_s_cla16_and299_y0;
  wire h_s_cla16_and300_y0;
  wire h_s_cla16_and301_y0;
  wire h_s_cla16_and302_y0;
  wire h_s_cla16_and303_y0;
  wire h_s_cla16_and304_y0;
  wire h_s_cla16_and305_y0;
  wire h_s_cla16_and306_y0;
  wire h_s_cla16_and307_y0;
  wire h_s_cla16_and308_y0;
  wire h_s_cla16_and309_y0;
  wire h_s_cla16_and310_y0;
  wire h_s_cla16_and311_y0;
  wire h_s_cla16_and312_y0;
  wire h_s_cla16_and313_y0;
  wire h_s_cla16_and314_y0;
  wire h_s_cla16_and315_y0;
  wire h_s_cla16_and316_y0;
  wire h_s_cla16_and317_y0;
  wire h_s_cla16_and318_y0;
  wire h_s_cla16_and319_y0;
  wire h_s_cla16_and320_y0;
  wire h_s_cla16_and321_y0;
  wire h_s_cla16_and322_y0;
  wire h_s_cla16_and323_y0;
  wire h_s_cla16_and324_y0;
  wire h_s_cla16_and325_y0;
  wire h_s_cla16_and326_y0;
  wire h_s_cla16_and327_y0;
  wire h_s_cla16_and328_y0;
  wire h_s_cla16_and329_y0;
  wire h_s_cla16_and330_y0;
  wire h_s_cla16_and331_y0;
  wire h_s_cla16_and332_y0;
  wire h_s_cla16_and333_y0;
  wire h_s_cla16_and334_y0;
  wire h_s_cla16_and335_y0;
  wire h_s_cla16_and336_y0;
  wire h_s_cla16_and337_y0;
  wire h_s_cla16_and338_y0;
  wire h_s_cla16_and339_y0;
  wire h_s_cla16_and340_y0;
  wire h_s_cla16_and341_y0;
  wire h_s_cla16_and342_y0;
  wire h_s_cla16_and343_y0;
  wire h_s_cla16_and344_y0;
  wire h_s_cla16_and345_y0;
  wire h_s_cla16_and346_y0;
  wire h_s_cla16_and347_y0;
  wire h_s_cla16_and348_y0;
  wire h_s_cla16_and349_y0;
  wire h_s_cla16_and350_y0;
  wire h_s_cla16_and351_y0;
  wire h_s_cla16_and352_y0;
  wire h_s_cla16_and353_y0;
  wire h_s_cla16_and354_y0;
  wire h_s_cla16_and355_y0;
  wire h_s_cla16_and356_y0;
  wire h_s_cla16_and357_y0;
  wire h_s_cla16_and358_y0;
  wire h_s_cla16_and359_y0;
  wire h_s_cla16_and360_y0;
  wire h_s_cla16_and361_y0;
  wire h_s_cla16_and362_y0;
  wire h_s_cla16_and363_y0;
  wire h_s_cla16_and364_y0;
  wire h_s_cla16_and365_y0;
  wire h_s_cla16_and366_y0;
  wire h_s_cla16_and367_y0;
  wire h_s_cla16_and368_y0;
  wire h_s_cla16_and369_y0;
  wire h_s_cla16_and370_y0;
  wire h_s_cla16_and371_y0;
  wire h_s_cla16_and372_y0;
  wire h_s_cla16_and373_y0;
  wire h_s_cla16_and374_y0;
  wire h_s_cla16_and375_y0;
  wire h_s_cla16_and376_y0;
  wire h_s_cla16_and377_y0;
  wire h_s_cla16_and378_y0;
  wire h_s_cla16_and379_y0;
  wire h_s_cla16_and380_y0;
  wire h_s_cla16_and381_y0;
  wire h_s_cla16_and382_y0;
  wire h_s_cla16_and383_y0;
  wire h_s_cla16_and384_y0;
  wire h_s_cla16_or45_y0;
  wire h_s_cla16_or46_y0;
  wire h_s_cla16_or47_y0;
  wire h_s_cla16_or48_y0;
  wire h_s_cla16_or49_y0;
  wire h_s_cla16_or50_y0;
  wire h_s_cla16_or51_y0;
  wire h_s_cla16_or52_y0;
  wire h_s_cla16_or53_y0;
  wire h_s_cla16_or54_y0;
  wire h_s_cla16_pg_logic10_y0;
  wire h_s_cla16_pg_logic10_y1;
  wire h_s_cla16_pg_logic10_y2;
  wire h_s_cla16_xor10_y0;
  wire h_s_cla16_and385_y0;
  wire h_s_cla16_and386_y0;
  wire h_s_cla16_and387_y0;
  wire h_s_cla16_and388_y0;
  wire h_s_cla16_and389_y0;
  wire h_s_cla16_and390_y0;
  wire h_s_cla16_and391_y0;
  wire h_s_cla16_and392_y0;
  wire h_s_cla16_and393_y0;
  wire h_s_cla16_and394_y0;
  wire h_s_cla16_and395_y0;
  wire h_s_cla16_and396_y0;
  wire h_s_cla16_and397_y0;
  wire h_s_cla16_and398_y0;
  wire h_s_cla16_and399_y0;
  wire h_s_cla16_and400_y0;
  wire h_s_cla16_and401_y0;
  wire h_s_cla16_and402_y0;
  wire h_s_cla16_and403_y0;
  wire h_s_cla16_and404_y0;
  wire h_s_cla16_and405_y0;
  wire h_s_cla16_and406_y0;
  wire h_s_cla16_and407_y0;
  wire h_s_cla16_and408_y0;
  wire h_s_cla16_and409_y0;
  wire h_s_cla16_and410_y0;
  wire h_s_cla16_and411_y0;
  wire h_s_cla16_and412_y0;
  wire h_s_cla16_and413_y0;
  wire h_s_cla16_and414_y0;
  wire h_s_cla16_and415_y0;
  wire h_s_cla16_and416_y0;
  wire h_s_cla16_and417_y0;
  wire h_s_cla16_and418_y0;
  wire h_s_cla16_and419_y0;
  wire h_s_cla16_and420_y0;
  wire h_s_cla16_and421_y0;
  wire h_s_cla16_and422_y0;
  wire h_s_cla16_and423_y0;
  wire h_s_cla16_and424_y0;
  wire h_s_cla16_and425_y0;
  wire h_s_cla16_and426_y0;
  wire h_s_cla16_and427_y0;
  wire h_s_cla16_and428_y0;
  wire h_s_cla16_and429_y0;
  wire h_s_cla16_and430_y0;
  wire h_s_cla16_and431_y0;
  wire h_s_cla16_and432_y0;
  wire h_s_cla16_and433_y0;
  wire h_s_cla16_and434_y0;
  wire h_s_cla16_and435_y0;
  wire h_s_cla16_and436_y0;
  wire h_s_cla16_and437_y0;
  wire h_s_cla16_and438_y0;
  wire h_s_cla16_and439_y0;
  wire h_s_cla16_and440_y0;
  wire h_s_cla16_and441_y0;
  wire h_s_cla16_and442_y0;
  wire h_s_cla16_and443_y0;
  wire h_s_cla16_and444_y0;
  wire h_s_cla16_and445_y0;
  wire h_s_cla16_and446_y0;
  wire h_s_cla16_and447_y0;
  wire h_s_cla16_and448_y0;
  wire h_s_cla16_and449_y0;
  wire h_s_cla16_and450_y0;
  wire h_s_cla16_and451_y0;
  wire h_s_cla16_and452_y0;
  wire h_s_cla16_and453_y0;
  wire h_s_cla16_and454_y0;
  wire h_s_cla16_and455_y0;
  wire h_s_cla16_and456_y0;
  wire h_s_cla16_and457_y0;
  wire h_s_cla16_and458_y0;
  wire h_s_cla16_and459_y0;
  wire h_s_cla16_and460_y0;
  wire h_s_cla16_and461_y0;
  wire h_s_cla16_and462_y0;
  wire h_s_cla16_and463_y0;
  wire h_s_cla16_and464_y0;
  wire h_s_cla16_and465_y0;
  wire h_s_cla16_and466_y0;
  wire h_s_cla16_and467_y0;
  wire h_s_cla16_and468_y0;
  wire h_s_cla16_and469_y0;
  wire h_s_cla16_and470_y0;
  wire h_s_cla16_and471_y0;
  wire h_s_cla16_and472_y0;
  wire h_s_cla16_and473_y0;
  wire h_s_cla16_and474_y0;
  wire h_s_cla16_and475_y0;
  wire h_s_cla16_and476_y0;
  wire h_s_cla16_and477_y0;
  wire h_s_cla16_and478_y0;
  wire h_s_cla16_and479_y0;
  wire h_s_cla16_and480_y0;
  wire h_s_cla16_and481_y0;
  wire h_s_cla16_and482_y0;
  wire h_s_cla16_and483_y0;
  wire h_s_cla16_and484_y0;
  wire h_s_cla16_and485_y0;
  wire h_s_cla16_and486_y0;
  wire h_s_cla16_and487_y0;
  wire h_s_cla16_and488_y0;
  wire h_s_cla16_and489_y0;
  wire h_s_cla16_and490_y0;
  wire h_s_cla16_and491_y0;
  wire h_s_cla16_and492_y0;
  wire h_s_cla16_and493_y0;
  wire h_s_cla16_and494_y0;
  wire h_s_cla16_and495_y0;
  wire h_s_cla16_and496_y0;
  wire h_s_cla16_and497_y0;
  wire h_s_cla16_and498_y0;
  wire h_s_cla16_and499_y0;
  wire h_s_cla16_and500_y0;
  wire h_s_cla16_and501_y0;
  wire h_s_cla16_and502_y0;
  wire h_s_cla16_and503_y0;
  wire h_s_cla16_and504_y0;
  wire h_s_cla16_and505_y0;
  wire h_s_cla16_or55_y0;
  wire h_s_cla16_or56_y0;
  wire h_s_cla16_or57_y0;
  wire h_s_cla16_or58_y0;
  wire h_s_cla16_or59_y0;
  wire h_s_cla16_or60_y0;
  wire h_s_cla16_or61_y0;
  wire h_s_cla16_or62_y0;
  wire h_s_cla16_or63_y0;
  wire h_s_cla16_or64_y0;
  wire h_s_cla16_or65_y0;
  wire h_s_cla16_pg_logic11_y0;
  wire h_s_cla16_pg_logic11_y1;
  wire h_s_cla16_pg_logic11_y2;
  wire h_s_cla16_xor11_y0;
  wire h_s_cla16_and506_y0;
  wire h_s_cla16_and507_y0;
  wire h_s_cla16_and508_y0;
  wire h_s_cla16_and509_y0;
  wire h_s_cla16_and510_y0;
  wire h_s_cla16_and511_y0;
  wire h_s_cla16_and512_y0;
  wire h_s_cla16_and513_y0;
  wire h_s_cla16_and514_y0;
  wire h_s_cla16_and515_y0;
  wire h_s_cla16_and516_y0;
  wire h_s_cla16_and517_y0;
  wire h_s_cla16_and518_y0;
  wire h_s_cla16_and519_y0;
  wire h_s_cla16_and520_y0;
  wire h_s_cla16_and521_y0;
  wire h_s_cla16_and522_y0;
  wire h_s_cla16_and523_y0;
  wire h_s_cla16_and524_y0;
  wire h_s_cla16_and525_y0;
  wire h_s_cla16_and526_y0;
  wire h_s_cla16_and527_y0;
  wire h_s_cla16_and528_y0;
  wire h_s_cla16_and529_y0;
  wire h_s_cla16_and530_y0;
  wire h_s_cla16_and531_y0;
  wire h_s_cla16_and532_y0;
  wire h_s_cla16_and533_y0;
  wire h_s_cla16_and534_y0;
  wire h_s_cla16_and535_y0;
  wire h_s_cla16_and536_y0;
  wire h_s_cla16_and537_y0;
  wire h_s_cla16_and538_y0;
  wire h_s_cla16_and539_y0;
  wire h_s_cla16_and540_y0;
  wire h_s_cla16_and541_y0;
  wire h_s_cla16_and542_y0;
  wire h_s_cla16_and543_y0;
  wire h_s_cla16_and544_y0;
  wire h_s_cla16_and545_y0;
  wire h_s_cla16_and546_y0;
  wire h_s_cla16_and547_y0;
  wire h_s_cla16_and548_y0;
  wire h_s_cla16_and549_y0;
  wire h_s_cla16_and550_y0;
  wire h_s_cla16_and551_y0;
  wire h_s_cla16_and552_y0;
  wire h_s_cla16_and553_y0;
  wire h_s_cla16_and554_y0;
  wire h_s_cla16_and555_y0;
  wire h_s_cla16_and556_y0;
  wire h_s_cla16_and557_y0;
  wire h_s_cla16_and558_y0;
  wire h_s_cla16_and559_y0;
  wire h_s_cla16_and560_y0;
  wire h_s_cla16_and561_y0;
  wire h_s_cla16_and562_y0;
  wire h_s_cla16_and563_y0;
  wire h_s_cla16_and564_y0;
  wire h_s_cla16_and565_y0;
  wire h_s_cla16_and566_y0;
  wire h_s_cla16_and567_y0;
  wire h_s_cla16_and568_y0;
  wire h_s_cla16_and569_y0;
  wire h_s_cla16_and570_y0;
  wire h_s_cla16_and571_y0;
  wire h_s_cla16_and572_y0;
  wire h_s_cla16_and573_y0;
  wire h_s_cla16_and574_y0;
  wire h_s_cla16_and575_y0;
  wire h_s_cla16_and576_y0;
  wire h_s_cla16_and577_y0;
  wire h_s_cla16_and578_y0;
  wire h_s_cla16_and579_y0;
  wire h_s_cla16_and580_y0;
  wire h_s_cla16_and581_y0;
  wire h_s_cla16_and582_y0;
  wire h_s_cla16_and583_y0;
  wire h_s_cla16_and584_y0;
  wire h_s_cla16_and585_y0;
  wire h_s_cla16_and586_y0;
  wire h_s_cla16_and587_y0;
  wire h_s_cla16_and588_y0;
  wire h_s_cla16_and589_y0;
  wire h_s_cla16_and590_y0;
  wire h_s_cla16_and591_y0;
  wire h_s_cla16_and592_y0;
  wire h_s_cla16_and593_y0;
  wire h_s_cla16_and594_y0;
  wire h_s_cla16_and595_y0;
  wire h_s_cla16_and596_y0;
  wire h_s_cla16_and597_y0;
  wire h_s_cla16_and598_y0;
  wire h_s_cla16_and599_y0;
  wire h_s_cla16_and600_y0;
  wire h_s_cla16_and601_y0;
  wire h_s_cla16_and602_y0;
  wire h_s_cla16_and603_y0;
  wire h_s_cla16_and604_y0;
  wire h_s_cla16_and605_y0;
  wire h_s_cla16_and606_y0;
  wire h_s_cla16_and607_y0;
  wire h_s_cla16_and608_y0;
  wire h_s_cla16_and609_y0;
  wire h_s_cla16_and610_y0;
  wire h_s_cla16_and611_y0;
  wire h_s_cla16_and612_y0;
  wire h_s_cla16_and613_y0;
  wire h_s_cla16_and614_y0;
  wire h_s_cla16_and615_y0;
  wire h_s_cla16_and616_y0;
  wire h_s_cla16_and617_y0;
  wire h_s_cla16_and618_y0;
  wire h_s_cla16_and619_y0;
  wire h_s_cla16_and620_y0;
  wire h_s_cla16_and621_y0;
  wire h_s_cla16_and622_y0;
  wire h_s_cla16_and623_y0;
  wire h_s_cla16_and624_y0;
  wire h_s_cla16_and625_y0;
  wire h_s_cla16_and626_y0;
  wire h_s_cla16_and627_y0;
  wire h_s_cla16_and628_y0;
  wire h_s_cla16_and629_y0;
  wire h_s_cla16_and630_y0;
  wire h_s_cla16_and631_y0;
  wire h_s_cla16_and632_y0;
  wire h_s_cla16_and633_y0;
  wire h_s_cla16_and634_y0;
  wire h_s_cla16_and635_y0;
  wire h_s_cla16_and636_y0;
  wire h_s_cla16_and637_y0;
  wire h_s_cla16_and638_y0;
  wire h_s_cla16_and639_y0;
  wire h_s_cla16_and640_y0;
  wire h_s_cla16_and641_y0;
  wire h_s_cla16_and642_y0;
  wire h_s_cla16_and643_y0;
  wire h_s_cla16_and644_y0;
  wire h_s_cla16_and645_y0;
  wire h_s_cla16_and646_y0;
  wire h_s_cla16_and647_y0;
  wire h_s_cla16_and648_y0;
  wire h_s_cla16_and649_y0;
  wire h_s_cla16_or66_y0;
  wire h_s_cla16_or67_y0;
  wire h_s_cla16_or68_y0;
  wire h_s_cla16_or69_y0;
  wire h_s_cla16_or70_y0;
  wire h_s_cla16_or71_y0;
  wire h_s_cla16_or72_y0;
  wire h_s_cla16_or73_y0;
  wire h_s_cla16_or74_y0;
  wire h_s_cla16_or75_y0;
  wire h_s_cla16_or76_y0;
  wire h_s_cla16_or77_y0;
  wire h_s_cla16_pg_logic12_y0;
  wire h_s_cla16_pg_logic12_y1;
  wire h_s_cla16_pg_logic12_y2;
  wire h_s_cla16_xor12_y0;
  wire h_s_cla16_and650_y0;
  wire h_s_cla16_and651_y0;
  wire h_s_cla16_and652_y0;
  wire h_s_cla16_and653_y0;
  wire h_s_cla16_and654_y0;
  wire h_s_cla16_and655_y0;
  wire h_s_cla16_and656_y0;
  wire h_s_cla16_and657_y0;
  wire h_s_cla16_and658_y0;
  wire h_s_cla16_and659_y0;
  wire h_s_cla16_and660_y0;
  wire h_s_cla16_and661_y0;
  wire h_s_cla16_and662_y0;
  wire h_s_cla16_and663_y0;
  wire h_s_cla16_and664_y0;
  wire h_s_cla16_and665_y0;
  wire h_s_cla16_and666_y0;
  wire h_s_cla16_and667_y0;
  wire h_s_cla16_and668_y0;
  wire h_s_cla16_and669_y0;
  wire h_s_cla16_and670_y0;
  wire h_s_cla16_and671_y0;
  wire h_s_cla16_and672_y0;
  wire h_s_cla16_and673_y0;
  wire h_s_cla16_and674_y0;
  wire h_s_cla16_and675_y0;
  wire h_s_cla16_and676_y0;
  wire h_s_cla16_and677_y0;
  wire h_s_cla16_and678_y0;
  wire h_s_cla16_and679_y0;
  wire h_s_cla16_and680_y0;
  wire h_s_cla16_and681_y0;
  wire h_s_cla16_and682_y0;
  wire h_s_cla16_and683_y0;
  wire h_s_cla16_and684_y0;
  wire h_s_cla16_and685_y0;
  wire h_s_cla16_and686_y0;
  wire h_s_cla16_and687_y0;
  wire h_s_cla16_and688_y0;
  wire h_s_cla16_and689_y0;
  wire h_s_cla16_and690_y0;
  wire h_s_cla16_and691_y0;
  wire h_s_cla16_and692_y0;
  wire h_s_cla16_and693_y0;
  wire h_s_cla16_and694_y0;
  wire h_s_cla16_and695_y0;
  wire h_s_cla16_and696_y0;
  wire h_s_cla16_and697_y0;
  wire h_s_cla16_and698_y0;
  wire h_s_cla16_and699_y0;
  wire h_s_cla16_and700_y0;
  wire h_s_cla16_and701_y0;
  wire h_s_cla16_and702_y0;
  wire h_s_cla16_and703_y0;
  wire h_s_cla16_and704_y0;
  wire h_s_cla16_and705_y0;
  wire h_s_cla16_and706_y0;
  wire h_s_cla16_and707_y0;
  wire h_s_cla16_and708_y0;
  wire h_s_cla16_and709_y0;
  wire h_s_cla16_and710_y0;
  wire h_s_cla16_and711_y0;
  wire h_s_cla16_and712_y0;
  wire h_s_cla16_and713_y0;
  wire h_s_cla16_and714_y0;
  wire h_s_cla16_and715_y0;
  wire h_s_cla16_and716_y0;
  wire h_s_cla16_and717_y0;
  wire h_s_cla16_and718_y0;
  wire h_s_cla16_and719_y0;
  wire h_s_cla16_and720_y0;
  wire h_s_cla16_and721_y0;
  wire h_s_cla16_and722_y0;
  wire h_s_cla16_and723_y0;
  wire h_s_cla16_and724_y0;
  wire h_s_cla16_and725_y0;
  wire h_s_cla16_and726_y0;
  wire h_s_cla16_and727_y0;
  wire h_s_cla16_and728_y0;
  wire h_s_cla16_and729_y0;
  wire h_s_cla16_and730_y0;
  wire h_s_cla16_and731_y0;
  wire h_s_cla16_and732_y0;
  wire h_s_cla16_and733_y0;
  wire h_s_cla16_and734_y0;
  wire h_s_cla16_and735_y0;
  wire h_s_cla16_and736_y0;
  wire h_s_cla16_and737_y0;
  wire h_s_cla16_and738_y0;
  wire h_s_cla16_and739_y0;
  wire h_s_cla16_and740_y0;
  wire h_s_cla16_and741_y0;
  wire h_s_cla16_and742_y0;
  wire h_s_cla16_and743_y0;
  wire h_s_cla16_and744_y0;
  wire h_s_cla16_and745_y0;
  wire h_s_cla16_and746_y0;
  wire h_s_cla16_and747_y0;
  wire h_s_cla16_and748_y0;
  wire h_s_cla16_and749_y0;
  wire h_s_cla16_and750_y0;
  wire h_s_cla16_and751_y0;
  wire h_s_cla16_and752_y0;
  wire h_s_cla16_and753_y0;
  wire h_s_cla16_and754_y0;
  wire h_s_cla16_and755_y0;
  wire h_s_cla16_and756_y0;
  wire h_s_cla16_and757_y0;
  wire h_s_cla16_and758_y0;
  wire h_s_cla16_and759_y0;
  wire h_s_cla16_and760_y0;
  wire h_s_cla16_and761_y0;
  wire h_s_cla16_and762_y0;
  wire h_s_cla16_and763_y0;
  wire h_s_cla16_and764_y0;
  wire h_s_cla16_and765_y0;
  wire h_s_cla16_and766_y0;
  wire h_s_cla16_and767_y0;
  wire h_s_cla16_and768_y0;
  wire h_s_cla16_and769_y0;
  wire h_s_cla16_and770_y0;
  wire h_s_cla16_and771_y0;
  wire h_s_cla16_and772_y0;
  wire h_s_cla16_and773_y0;
  wire h_s_cla16_and774_y0;
  wire h_s_cla16_and775_y0;
  wire h_s_cla16_and776_y0;
  wire h_s_cla16_and777_y0;
  wire h_s_cla16_and778_y0;
  wire h_s_cla16_and779_y0;
  wire h_s_cla16_and780_y0;
  wire h_s_cla16_and781_y0;
  wire h_s_cla16_and782_y0;
  wire h_s_cla16_and783_y0;
  wire h_s_cla16_and784_y0;
  wire h_s_cla16_and785_y0;
  wire h_s_cla16_and786_y0;
  wire h_s_cla16_and787_y0;
  wire h_s_cla16_and788_y0;
  wire h_s_cla16_and789_y0;
  wire h_s_cla16_and790_y0;
  wire h_s_cla16_and791_y0;
  wire h_s_cla16_and792_y0;
  wire h_s_cla16_and793_y0;
  wire h_s_cla16_and794_y0;
  wire h_s_cla16_and795_y0;
  wire h_s_cla16_and796_y0;
  wire h_s_cla16_and797_y0;
  wire h_s_cla16_and798_y0;
  wire h_s_cla16_and799_y0;
  wire h_s_cla16_and800_y0;
  wire h_s_cla16_and801_y0;
  wire h_s_cla16_and802_y0;
  wire h_s_cla16_and803_y0;
  wire h_s_cla16_and804_y0;
  wire h_s_cla16_and805_y0;
  wire h_s_cla16_and806_y0;
  wire h_s_cla16_and807_y0;
  wire h_s_cla16_and808_y0;
  wire h_s_cla16_and809_y0;
  wire h_s_cla16_and810_y0;
  wire h_s_cla16_and811_y0;
  wire h_s_cla16_and812_y0;
  wire h_s_cla16_and813_y0;
  wire h_s_cla16_and814_y0;
  wire h_s_cla16_and815_y0;
  wire h_s_cla16_and816_y0;
  wire h_s_cla16_and817_y0;
  wire h_s_cla16_and818_y0;
  wire h_s_cla16_or78_y0;
  wire h_s_cla16_or79_y0;
  wire h_s_cla16_or80_y0;
  wire h_s_cla16_or81_y0;
  wire h_s_cla16_or82_y0;
  wire h_s_cla16_or83_y0;
  wire h_s_cla16_or84_y0;
  wire h_s_cla16_or85_y0;
  wire h_s_cla16_or86_y0;
  wire h_s_cla16_or87_y0;
  wire h_s_cla16_or88_y0;
  wire h_s_cla16_or89_y0;
  wire h_s_cla16_or90_y0;
  wire h_s_cla16_pg_logic13_y0;
  wire h_s_cla16_pg_logic13_y1;
  wire h_s_cla16_pg_logic13_y2;
  wire h_s_cla16_xor13_y0;
  wire h_s_cla16_and819_y0;
  wire h_s_cla16_and820_y0;
  wire h_s_cla16_and821_y0;
  wire h_s_cla16_and822_y0;
  wire h_s_cla16_and823_y0;
  wire h_s_cla16_and824_y0;
  wire h_s_cla16_and825_y0;
  wire h_s_cla16_and826_y0;
  wire h_s_cla16_and827_y0;
  wire h_s_cla16_and828_y0;
  wire h_s_cla16_and829_y0;
  wire h_s_cla16_and830_y0;
  wire h_s_cla16_and831_y0;
  wire h_s_cla16_and832_y0;
  wire h_s_cla16_and833_y0;
  wire h_s_cla16_and834_y0;
  wire h_s_cla16_and835_y0;
  wire h_s_cla16_and836_y0;
  wire h_s_cla16_and837_y0;
  wire h_s_cla16_and838_y0;
  wire h_s_cla16_and839_y0;
  wire h_s_cla16_and840_y0;
  wire h_s_cla16_and841_y0;
  wire h_s_cla16_and842_y0;
  wire h_s_cla16_and843_y0;
  wire h_s_cla16_and844_y0;
  wire h_s_cla16_and845_y0;
  wire h_s_cla16_and846_y0;
  wire h_s_cla16_and847_y0;
  wire h_s_cla16_and848_y0;
  wire h_s_cla16_and849_y0;
  wire h_s_cla16_and850_y0;
  wire h_s_cla16_and851_y0;
  wire h_s_cla16_and852_y0;
  wire h_s_cla16_and853_y0;
  wire h_s_cla16_and854_y0;
  wire h_s_cla16_and855_y0;
  wire h_s_cla16_and856_y0;
  wire h_s_cla16_and857_y0;
  wire h_s_cla16_and858_y0;
  wire h_s_cla16_and859_y0;
  wire h_s_cla16_and860_y0;
  wire h_s_cla16_and861_y0;
  wire h_s_cla16_and862_y0;
  wire h_s_cla16_and863_y0;
  wire h_s_cla16_and864_y0;
  wire h_s_cla16_and865_y0;
  wire h_s_cla16_and866_y0;
  wire h_s_cla16_and867_y0;
  wire h_s_cla16_and868_y0;
  wire h_s_cla16_and869_y0;
  wire h_s_cla16_and870_y0;
  wire h_s_cla16_and871_y0;
  wire h_s_cla16_and872_y0;
  wire h_s_cla16_and873_y0;
  wire h_s_cla16_and874_y0;
  wire h_s_cla16_and875_y0;
  wire h_s_cla16_and876_y0;
  wire h_s_cla16_and877_y0;
  wire h_s_cla16_and878_y0;
  wire h_s_cla16_and879_y0;
  wire h_s_cla16_and880_y0;
  wire h_s_cla16_and881_y0;
  wire h_s_cla16_and882_y0;
  wire h_s_cla16_and883_y0;
  wire h_s_cla16_and884_y0;
  wire h_s_cla16_and885_y0;
  wire h_s_cla16_and886_y0;
  wire h_s_cla16_and887_y0;
  wire h_s_cla16_and888_y0;
  wire h_s_cla16_and889_y0;
  wire h_s_cla16_and890_y0;
  wire h_s_cla16_and891_y0;
  wire h_s_cla16_and892_y0;
  wire h_s_cla16_and893_y0;
  wire h_s_cla16_and894_y0;
  wire h_s_cla16_and895_y0;
  wire h_s_cla16_and896_y0;
  wire h_s_cla16_and897_y0;
  wire h_s_cla16_and898_y0;
  wire h_s_cla16_and899_y0;
  wire h_s_cla16_and900_y0;
  wire h_s_cla16_and901_y0;
  wire h_s_cla16_and902_y0;
  wire h_s_cla16_and903_y0;
  wire h_s_cla16_and904_y0;
  wire h_s_cla16_and905_y0;
  wire h_s_cla16_and906_y0;
  wire h_s_cla16_and907_y0;
  wire h_s_cla16_and908_y0;
  wire h_s_cla16_and909_y0;
  wire h_s_cla16_and910_y0;
  wire h_s_cla16_and911_y0;
  wire h_s_cla16_and912_y0;
  wire h_s_cla16_and913_y0;
  wire h_s_cla16_and914_y0;
  wire h_s_cla16_and915_y0;
  wire h_s_cla16_and916_y0;
  wire h_s_cla16_and917_y0;
  wire h_s_cla16_and918_y0;
  wire h_s_cla16_and919_y0;
  wire h_s_cla16_and920_y0;
  wire h_s_cla16_and921_y0;
  wire h_s_cla16_and922_y0;
  wire h_s_cla16_and923_y0;
  wire h_s_cla16_and924_y0;
  wire h_s_cla16_and925_y0;
  wire h_s_cla16_and926_y0;
  wire h_s_cla16_and927_y0;
  wire h_s_cla16_and928_y0;
  wire h_s_cla16_and929_y0;
  wire h_s_cla16_and930_y0;
  wire h_s_cla16_and931_y0;
  wire h_s_cla16_and932_y0;
  wire h_s_cla16_and933_y0;
  wire h_s_cla16_and934_y0;
  wire h_s_cla16_and935_y0;
  wire h_s_cla16_and936_y0;
  wire h_s_cla16_and937_y0;
  wire h_s_cla16_and938_y0;
  wire h_s_cla16_and939_y0;
  wire h_s_cla16_and940_y0;
  wire h_s_cla16_and941_y0;
  wire h_s_cla16_and942_y0;
  wire h_s_cla16_and943_y0;
  wire h_s_cla16_and944_y0;
  wire h_s_cla16_and945_y0;
  wire h_s_cla16_and946_y0;
  wire h_s_cla16_and947_y0;
  wire h_s_cla16_and948_y0;
  wire h_s_cla16_and949_y0;
  wire h_s_cla16_and950_y0;
  wire h_s_cla16_and951_y0;
  wire h_s_cla16_and952_y0;
  wire h_s_cla16_and953_y0;
  wire h_s_cla16_and954_y0;
  wire h_s_cla16_and955_y0;
  wire h_s_cla16_and956_y0;
  wire h_s_cla16_and957_y0;
  wire h_s_cla16_and958_y0;
  wire h_s_cla16_and959_y0;
  wire h_s_cla16_and960_y0;
  wire h_s_cla16_and961_y0;
  wire h_s_cla16_and962_y0;
  wire h_s_cla16_and963_y0;
  wire h_s_cla16_and964_y0;
  wire h_s_cla16_and965_y0;
  wire h_s_cla16_and966_y0;
  wire h_s_cla16_and967_y0;
  wire h_s_cla16_and968_y0;
  wire h_s_cla16_and969_y0;
  wire h_s_cla16_and970_y0;
  wire h_s_cla16_and971_y0;
  wire h_s_cla16_and972_y0;
  wire h_s_cla16_and973_y0;
  wire h_s_cla16_and974_y0;
  wire h_s_cla16_and975_y0;
  wire h_s_cla16_and976_y0;
  wire h_s_cla16_and977_y0;
  wire h_s_cla16_and978_y0;
  wire h_s_cla16_and979_y0;
  wire h_s_cla16_and980_y0;
  wire h_s_cla16_and981_y0;
  wire h_s_cla16_and982_y0;
  wire h_s_cla16_and983_y0;
  wire h_s_cla16_and984_y0;
  wire h_s_cla16_and985_y0;
  wire h_s_cla16_and986_y0;
  wire h_s_cla16_and987_y0;
  wire h_s_cla16_and988_y0;
  wire h_s_cla16_and989_y0;
  wire h_s_cla16_and990_y0;
  wire h_s_cla16_and991_y0;
  wire h_s_cla16_and992_y0;
  wire h_s_cla16_and993_y0;
  wire h_s_cla16_and994_y0;
  wire h_s_cla16_and995_y0;
  wire h_s_cla16_and996_y0;
  wire h_s_cla16_and997_y0;
  wire h_s_cla16_and998_y0;
  wire h_s_cla16_and999_y0;
  wire h_s_cla16_and1000_y0;
  wire h_s_cla16_and1001_y0;
  wire h_s_cla16_and1002_y0;
  wire h_s_cla16_and1003_y0;
  wire h_s_cla16_and1004_y0;
  wire h_s_cla16_and1005_y0;
  wire h_s_cla16_and1006_y0;
  wire h_s_cla16_and1007_y0;
  wire h_s_cla16_and1008_y0;
  wire h_s_cla16_and1009_y0;
  wire h_s_cla16_and1010_y0;
  wire h_s_cla16_and1011_y0;
  wire h_s_cla16_and1012_y0;
  wire h_s_cla16_and1013_y0;
  wire h_s_cla16_and1014_y0;
  wire h_s_cla16_or91_y0;
  wire h_s_cla16_or92_y0;
  wire h_s_cla16_or93_y0;
  wire h_s_cla16_or94_y0;
  wire h_s_cla16_or95_y0;
  wire h_s_cla16_or96_y0;
  wire h_s_cla16_or97_y0;
  wire h_s_cla16_or98_y0;
  wire h_s_cla16_or99_y0;
  wire h_s_cla16_or100_y0;
  wire h_s_cla16_or101_y0;
  wire h_s_cla16_or102_y0;
  wire h_s_cla16_or103_y0;
  wire h_s_cla16_or104_y0;
  wire h_s_cla16_pg_logic14_y0;
  wire h_s_cla16_pg_logic14_y1;
  wire h_s_cla16_pg_logic14_y2;
  wire h_s_cla16_xor14_y0;
  wire h_s_cla16_and1015_y0;
  wire h_s_cla16_and1016_y0;
  wire h_s_cla16_and1017_y0;
  wire h_s_cla16_and1018_y0;
  wire h_s_cla16_and1019_y0;
  wire h_s_cla16_and1020_y0;
  wire h_s_cla16_and1021_y0;
  wire h_s_cla16_and1022_y0;
  wire h_s_cla16_and1023_y0;
  wire h_s_cla16_and1024_y0;
  wire h_s_cla16_and1025_y0;
  wire h_s_cla16_and1026_y0;
  wire h_s_cla16_and1027_y0;
  wire h_s_cla16_and1028_y0;
  wire h_s_cla16_and1029_y0;
  wire h_s_cla16_and1030_y0;
  wire h_s_cla16_and1031_y0;
  wire h_s_cla16_and1032_y0;
  wire h_s_cla16_and1033_y0;
  wire h_s_cla16_and1034_y0;
  wire h_s_cla16_and1035_y0;
  wire h_s_cla16_and1036_y0;
  wire h_s_cla16_and1037_y0;
  wire h_s_cla16_and1038_y0;
  wire h_s_cla16_and1039_y0;
  wire h_s_cla16_and1040_y0;
  wire h_s_cla16_and1041_y0;
  wire h_s_cla16_and1042_y0;
  wire h_s_cla16_and1043_y0;
  wire h_s_cla16_and1044_y0;
  wire h_s_cla16_and1045_y0;
  wire h_s_cla16_and1046_y0;
  wire h_s_cla16_and1047_y0;
  wire h_s_cla16_and1048_y0;
  wire h_s_cla16_and1049_y0;
  wire h_s_cla16_and1050_y0;
  wire h_s_cla16_and1051_y0;
  wire h_s_cla16_and1052_y0;
  wire h_s_cla16_and1053_y0;
  wire h_s_cla16_and1054_y0;
  wire h_s_cla16_and1055_y0;
  wire h_s_cla16_and1056_y0;
  wire h_s_cla16_and1057_y0;
  wire h_s_cla16_and1058_y0;
  wire h_s_cla16_and1059_y0;
  wire h_s_cla16_and1060_y0;
  wire h_s_cla16_and1061_y0;
  wire h_s_cla16_and1062_y0;
  wire h_s_cla16_and1063_y0;
  wire h_s_cla16_and1064_y0;
  wire h_s_cla16_and1065_y0;
  wire h_s_cla16_and1066_y0;
  wire h_s_cla16_and1067_y0;
  wire h_s_cla16_and1068_y0;
  wire h_s_cla16_and1069_y0;
  wire h_s_cla16_and1070_y0;
  wire h_s_cla16_and1071_y0;
  wire h_s_cla16_and1072_y0;
  wire h_s_cla16_and1073_y0;
  wire h_s_cla16_and1074_y0;
  wire h_s_cla16_and1075_y0;
  wire h_s_cla16_and1076_y0;
  wire h_s_cla16_and1077_y0;
  wire h_s_cla16_and1078_y0;
  wire h_s_cla16_and1079_y0;
  wire h_s_cla16_and1080_y0;
  wire h_s_cla16_and1081_y0;
  wire h_s_cla16_and1082_y0;
  wire h_s_cla16_and1083_y0;
  wire h_s_cla16_and1084_y0;
  wire h_s_cla16_and1085_y0;
  wire h_s_cla16_and1086_y0;
  wire h_s_cla16_and1087_y0;
  wire h_s_cla16_and1088_y0;
  wire h_s_cla16_and1089_y0;
  wire h_s_cla16_and1090_y0;
  wire h_s_cla16_and1091_y0;
  wire h_s_cla16_and1092_y0;
  wire h_s_cla16_and1093_y0;
  wire h_s_cla16_and1094_y0;
  wire h_s_cla16_and1095_y0;
  wire h_s_cla16_and1096_y0;
  wire h_s_cla16_and1097_y0;
  wire h_s_cla16_and1098_y0;
  wire h_s_cla16_and1099_y0;
  wire h_s_cla16_and1100_y0;
  wire h_s_cla16_and1101_y0;
  wire h_s_cla16_and1102_y0;
  wire h_s_cla16_and1103_y0;
  wire h_s_cla16_and1104_y0;
  wire h_s_cla16_and1105_y0;
  wire h_s_cla16_and1106_y0;
  wire h_s_cla16_and1107_y0;
  wire h_s_cla16_and1108_y0;
  wire h_s_cla16_and1109_y0;
  wire h_s_cla16_and1110_y0;
  wire h_s_cla16_and1111_y0;
  wire h_s_cla16_and1112_y0;
  wire h_s_cla16_and1113_y0;
  wire h_s_cla16_and1114_y0;
  wire h_s_cla16_and1115_y0;
  wire h_s_cla16_and1116_y0;
  wire h_s_cla16_and1117_y0;
  wire h_s_cla16_and1118_y0;
  wire h_s_cla16_and1119_y0;
  wire h_s_cla16_and1120_y0;
  wire h_s_cla16_and1121_y0;
  wire h_s_cla16_and1122_y0;
  wire h_s_cla16_and1123_y0;
  wire h_s_cla16_and1124_y0;
  wire h_s_cla16_and1125_y0;
  wire h_s_cla16_and1126_y0;
  wire h_s_cla16_and1127_y0;
  wire h_s_cla16_and1128_y0;
  wire h_s_cla16_and1129_y0;
  wire h_s_cla16_and1130_y0;
  wire h_s_cla16_and1131_y0;
  wire h_s_cla16_and1132_y0;
  wire h_s_cla16_and1133_y0;
  wire h_s_cla16_and1134_y0;
  wire h_s_cla16_and1135_y0;
  wire h_s_cla16_and1136_y0;
  wire h_s_cla16_and1137_y0;
  wire h_s_cla16_and1138_y0;
  wire h_s_cla16_and1139_y0;
  wire h_s_cla16_and1140_y0;
  wire h_s_cla16_and1141_y0;
  wire h_s_cla16_and1142_y0;
  wire h_s_cla16_and1143_y0;
  wire h_s_cla16_and1144_y0;
  wire h_s_cla16_and1145_y0;
  wire h_s_cla16_and1146_y0;
  wire h_s_cla16_and1147_y0;
  wire h_s_cla16_and1148_y0;
  wire h_s_cla16_and1149_y0;
  wire h_s_cla16_and1150_y0;
  wire h_s_cla16_and1151_y0;
  wire h_s_cla16_and1152_y0;
  wire h_s_cla16_and1153_y0;
  wire h_s_cla16_and1154_y0;
  wire h_s_cla16_and1155_y0;
  wire h_s_cla16_and1156_y0;
  wire h_s_cla16_and1157_y0;
  wire h_s_cla16_and1158_y0;
  wire h_s_cla16_and1159_y0;
  wire h_s_cla16_and1160_y0;
  wire h_s_cla16_and1161_y0;
  wire h_s_cla16_and1162_y0;
  wire h_s_cla16_and1163_y0;
  wire h_s_cla16_and1164_y0;
  wire h_s_cla16_and1165_y0;
  wire h_s_cla16_and1166_y0;
  wire h_s_cla16_and1167_y0;
  wire h_s_cla16_and1168_y0;
  wire h_s_cla16_and1169_y0;
  wire h_s_cla16_and1170_y0;
  wire h_s_cla16_and1171_y0;
  wire h_s_cla16_and1172_y0;
  wire h_s_cla16_and1173_y0;
  wire h_s_cla16_and1174_y0;
  wire h_s_cla16_and1175_y0;
  wire h_s_cla16_and1176_y0;
  wire h_s_cla16_and1177_y0;
  wire h_s_cla16_and1178_y0;
  wire h_s_cla16_and1179_y0;
  wire h_s_cla16_and1180_y0;
  wire h_s_cla16_and1181_y0;
  wire h_s_cla16_and1182_y0;
  wire h_s_cla16_and1183_y0;
  wire h_s_cla16_and1184_y0;
  wire h_s_cla16_and1185_y0;
  wire h_s_cla16_and1186_y0;
  wire h_s_cla16_and1187_y0;
  wire h_s_cla16_and1188_y0;
  wire h_s_cla16_and1189_y0;
  wire h_s_cla16_and1190_y0;
  wire h_s_cla16_and1191_y0;
  wire h_s_cla16_and1192_y0;
  wire h_s_cla16_and1193_y0;
  wire h_s_cla16_and1194_y0;
  wire h_s_cla16_and1195_y0;
  wire h_s_cla16_and1196_y0;
  wire h_s_cla16_and1197_y0;
  wire h_s_cla16_and1198_y0;
  wire h_s_cla16_and1199_y0;
  wire h_s_cla16_and1200_y0;
  wire h_s_cla16_and1201_y0;
  wire h_s_cla16_and1202_y0;
  wire h_s_cla16_and1203_y0;
  wire h_s_cla16_and1204_y0;
  wire h_s_cla16_and1205_y0;
  wire h_s_cla16_and1206_y0;
  wire h_s_cla16_and1207_y0;
  wire h_s_cla16_and1208_y0;
  wire h_s_cla16_and1209_y0;
  wire h_s_cla16_and1210_y0;
  wire h_s_cla16_and1211_y0;
  wire h_s_cla16_and1212_y0;
  wire h_s_cla16_and1213_y0;
  wire h_s_cla16_and1214_y0;
  wire h_s_cla16_and1215_y0;
  wire h_s_cla16_and1216_y0;
  wire h_s_cla16_and1217_y0;
  wire h_s_cla16_and1218_y0;
  wire h_s_cla16_and1219_y0;
  wire h_s_cla16_and1220_y0;
  wire h_s_cla16_and1221_y0;
  wire h_s_cla16_and1222_y0;
  wire h_s_cla16_and1223_y0;
  wire h_s_cla16_and1224_y0;
  wire h_s_cla16_and1225_y0;
  wire h_s_cla16_and1226_y0;
  wire h_s_cla16_and1227_y0;
  wire h_s_cla16_and1228_y0;
  wire h_s_cla16_and1229_y0;
  wire h_s_cla16_and1230_y0;
  wire h_s_cla16_and1231_y0;
  wire h_s_cla16_and1232_y0;
  wire h_s_cla16_and1233_y0;
  wire h_s_cla16_and1234_y0;
  wire h_s_cla16_and1235_y0;
  wire h_s_cla16_and1236_y0;
  wire h_s_cla16_and1237_y0;
  wire h_s_cla16_and1238_y0;
  wire h_s_cla16_and1239_y0;
  wire h_s_cla16_or105_y0;
  wire h_s_cla16_or106_y0;
  wire h_s_cla16_or107_y0;
  wire h_s_cla16_or108_y0;
  wire h_s_cla16_or109_y0;
  wire h_s_cla16_or110_y0;
  wire h_s_cla16_or111_y0;
  wire h_s_cla16_or112_y0;
  wire h_s_cla16_or113_y0;
  wire h_s_cla16_or114_y0;
  wire h_s_cla16_or115_y0;
  wire h_s_cla16_or116_y0;
  wire h_s_cla16_or117_y0;
  wire h_s_cla16_or118_y0;
  wire h_s_cla16_or119_y0;
  wire h_s_cla16_pg_logic15_y0;
  wire h_s_cla16_pg_logic15_y1;
  wire h_s_cla16_pg_logic15_y2;
  wire h_s_cla16_xor15_y0;
  wire h_s_cla16_and1240_y0;
  wire h_s_cla16_and1241_y0;
  wire h_s_cla16_and1242_y0;
  wire h_s_cla16_and1243_y0;
  wire h_s_cla16_and1244_y0;
  wire h_s_cla16_and1245_y0;
  wire h_s_cla16_and1246_y0;
  wire h_s_cla16_and1247_y0;
  wire h_s_cla16_and1248_y0;
  wire h_s_cla16_and1249_y0;
  wire h_s_cla16_and1250_y0;
  wire h_s_cla16_and1251_y0;
  wire h_s_cla16_and1252_y0;
  wire h_s_cla16_and1253_y0;
  wire h_s_cla16_and1254_y0;
  wire h_s_cla16_and1255_y0;
  wire h_s_cla16_and1256_y0;
  wire h_s_cla16_and1257_y0;
  wire h_s_cla16_and1258_y0;
  wire h_s_cla16_and1259_y0;
  wire h_s_cla16_and1260_y0;
  wire h_s_cla16_and1261_y0;
  wire h_s_cla16_and1262_y0;
  wire h_s_cla16_and1263_y0;
  wire h_s_cla16_and1264_y0;
  wire h_s_cla16_and1265_y0;
  wire h_s_cla16_and1266_y0;
  wire h_s_cla16_and1267_y0;
  wire h_s_cla16_and1268_y0;
  wire h_s_cla16_and1269_y0;
  wire h_s_cla16_and1270_y0;
  wire h_s_cla16_and1271_y0;
  wire h_s_cla16_and1272_y0;
  wire h_s_cla16_and1273_y0;
  wire h_s_cla16_and1274_y0;
  wire h_s_cla16_and1275_y0;
  wire h_s_cla16_and1276_y0;
  wire h_s_cla16_and1277_y0;
  wire h_s_cla16_and1278_y0;
  wire h_s_cla16_and1279_y0;
  wire h_s_cla16_and1280_y0;
  wire h_s_cla16_and1281_y0;
  wire h_s_cla16_and1282_y0;
  wire h_s_cla16_and1283_y0;
  wire h_s_cla16_and1284_y0;
  wire h_s_cla16_and1285_y0;
  wire h_s_cla16_and1286_y0;
  wire h_s_cla16_and1287_y0;
  wire h_s_cla16_and1288_y0;
  wire h_s_cla16_and1289_y0;
  wire h_s_cla16_and1290_y0;
  wire h_s_cla16_and1291_y0;
  wire h_s_cla16_and1292_y0;
  wire h_s_cla16_and1293_y0;
  wire h_s_cla16_and1294_y0;
  wire h_s_cla16_and1295_y0;
  wire h_s_cla16_and1296_y0;
  wire h_s_cla16_and1297_y0;
  wire h_s_cla16_and1298_y0;
  wire h_s_cla16_and1299_y0;
  wire h_s_cla16_and1300_y0;
  wire h_s_cla16_and1301_y0;
  wire h_s_cla16_and1302_y0;
  wire h_s_cla16_and1303_y0;
  wire h_s_cla16_and1304_y0;
  wire h_s_cla16_and1305_y0;
  wire h_s_cla16_and1306_y0;
  wire h_s_cla16_and1307_y0;
  wire h_s_cla16_and1308_y0;
  wire h_s_cla16_and1309_y0;
  wire h_s_cla16_and1310_y0;
  wire h_s_cla16_and1311_y0;
  wire h_s_cla16_and1312_y0;
  wire h_s_cla16_and1313_y0;
  wire h_s_cla16_and1314_y0;
  wire h_s_cla16_and1315_y0;
  wire h_s_cla16_and1316_y0;
  wire h_s_cla16_and1317_y0;
  wire h_s_cla16_and1318_y0;
  wire h_s_cla16_and1319_y0;
  wire h_s_cla16_and1320_y0;
  wire h_s_cla16_and1321_y0;
  wire h_s_cla16_and1322_y0;
  wire h_s_cla16_and1323_y0;
  wire h_s_cla16_and1324_y0;
  wire h_s_cla16_and1325_y0;
  wire h_s_cla16_and1326_y0;
  wire h_s_cla16_and1327_y0;
  wire h_s_cla16_and1328_y0;
  wire h_s_cla16_and1329_y0;
  wire h_s_cla16_and1330_y0;
  wire h_s_cla16_and1331_y0;
  wire h_s_cla16_and1332_y0;
  wire h_s_cla16_and1333_y0;
  wire h_s_cla16_and1334_y0;
  wire h_s_cla16_and1335_y0;
  wire h_s_cla16_and1336_y0;
  wire h_s_cla16_and1337_y0;
  wire h_s_cla16_and1338_y0;
  wire h_s_cla16_and1339_y0;
  wire h_s_cla16_and1340_y0;
  wire h_s_cla16_and1341_y0;
  wire h_s_cla16_and1342_y0;
  wire h_s_cla16_and1343_y0;
  wire h_s_cla16_and1344_y0;
  wire h_s_cla16_and1345_y0;
  wire h_s_cla16_and1346_y0;
  wire h_s_cla16_and1347_y0;
  wire h_s_cla16_and1348_y0;
  wire h_s_cla16_and1349_y0;
  wire h_s_cla16_and1350_y0;
  wire h_s_cla16_and1351_y0;
  wire h_s_cla16_and1352_y0;
  wire h_s_cla16_and1353_y0;
  wire h_s_cla16_and1354_y0;
  wire h_s_cla16_and1355_y0;
  wire h_s_cla16_and1356_y0;
  wire h_s_cla16_and1357_y0;
  wire h_s_cla16_and1358_y0;
  wire h_s_cla16_and1359_y0;
  wire h_s_cla16_and1360_y0;
  wire h_s_cla16_and1361_y0;
  wire h_s_cla16_and1362_y0;
  wire h_s_cla16_and1363_y0;
  wire h_s_cla16_and1364_y0;
  wire h_s_cla16_and1365_y0;
  wire h_s_cla16_and1366_y0;
  wire h_s_cla16_and1367_y0;
  wire h_s_cla16_and1368_y0;
  wire h_s_cla16_and1369_y0;
  wire h_s_cla16_and1370_y0;
  wire h_s_cla16_and1371_y0;
  wire h_s_cla16_and1372_y0;
  wire h_s_cla16_and1373_y0;
  wire h_s_cla16_and1374_y0;
  wire h_s_cla16_and1375_y0;
  wire h_s_cla16_and1376_y0;
  wire h_s_cla16_and1377_y0;
  wire h_s_cla16_and1378_y0;
  wire h_s_cla16_and1379_y0;
  wire h_s_cla16_and1380_y0;
  wire h_s_cla16_and1381_y0;
  wire h_s_cla16_and1382_y0;
  wire h_s_cla16_and1383_y0;
  wire h_s_cla16_and1384_y0;
  wire h_s_cla16_and1385_y0;
  wire h_s_cla16_and1386_y0;
  wire h_s_cla16_and1387_y0;
  wire h_s_cla16_and1388_y0;
  wire h_s_cla16_and1389_y0;
  wire h_s_cla16_and1390_y0;
  wire h_s_cla16_and1391_y0;
  wire h_s_cla16_and1392_y0;
  wire h_s_cla16_and1393_y0;
  wire h_s_cla16_and1394_y0;
  wire h_s_cla16_and1395_y0;
  wire h_s_cla16_and1396_y0;
  wire h_s_cla16_and1397_y0;
  wire h_s_cla16_and1398_y0;
  wire h_s_cla16_and1399_y0;
  wire h_s_cla16_and1400_y0;
  wire h_s_cla16_and1401_y0;
  wire h_s_cla16_and1402_y0;
  wire h_s_cla16_and1403_y0;
  wire h_s_cla16_and1404_y0;
  wire h_s_cla16_and1405_y0;
  wire h_s_cla16_and1406_y0;
  wire h_s_cla16_and1407_y0;
  wire h_s_cla16_and1408_y0;
  wire h_s_cla16_and1409_y0;
  wire h_s_cla16_and1410_y0;
  wire h_s_cla16_and1411_y0;
  wire h_s_cla16_and1412_y0;
  wire h_s_cla16_and1413_y0;
  wire h_s_cla16_and1414_y0;
  wire h_s_cla16_and1415_y0;
  wire h_s_cla16_and1416_y0;
  wire h_s_cla16_and1417_y0;
  wire h_s_cla16_and1418_y0;
  wire h_s_cla16_and1419_y0;
  wire h_s_cla16_and1420_y0;
  wire h_s_cla16_and1421_y0;
  wire h_s_cla16_and1422_y0;
  wire h_s_cla16_and1423_y0;
  wire h_s_cla16_and1424_y0;
  wire h_s_cla16_and1425_y0;
  wire h_s_cla16_and1426_y0;
  wire h_s_cla16_and1427_y0;
  wire h_s_cla16_and1428_y0;
  wire h_s_cla16_and1429_y0;
  wire h_s_cla16_and1430_y0;
  wire h_s_cla16_and1431_y0;
  wire h_s_cla16_and1432_y0;
  wire h_s_cla16_and1433_y0;
  wire h_s_cla16_and1434_y0;
  wire h_s_cla16_and1435_y0;
  wire h_s_cla16_and1436_y0;
  wire h_s_cla16_and1437_y0;
  wire h_s_cla16_and1438_y0;
  wire h_s_cla16_and1439_y0;
  wire h_s_cla16_and1440_y0;
  wire h_s_cla16_and1441_y0;
  wire h_s_cla16_and1442_y0;
  wire h_s_cla16_and1443_y0;
  wire h_s_cla16_and1444_y0;
  wire h_s_cla16_and1445_y0;
  wire h_s_cla16_and1446_y0;
  wire h_s_cla16_and1447_y0;
  wire h_s_cla16_and1448_y0;
  wire h_s_cla16_and1449_y0;
  wire h_s_cla16_and1450_y0;
  wire h_s_cla16_and1451_y0;
  wire h_s_cla16_and1452_y0;
  wire h_s_cla16_and1453_y0;
  wire h_s_cla16_and1454_y0;
  wire h_s_cla16_and1455_y0;
  wire h_s_cla16_and1456_y0;
  wire h_s_cla16_and1457_y0;
  wire h_s_cla16_and1458_y0;
  wire h_s_cla16_and1459_y0;
  wire h_s_cla16_and1460_y0;
  wire h_s_cla16_and1461_y0;
  wire h_s_cla16_and1462_y0;
  wire h_s_cla16_and1463_y0;
  wire h_s_cla16_and1464_y0;
  wire h_s_cla16_and1465_y0;
  wire h_s_cla16_and1466_y0;
  wire h_s_cla16_and1467_y0;
  wire h_s_cla16_and1468_y0;
  wire h_s_cla16_and1469_y0;
  wire h_s_cla16_and1470_y0;
  wire h_s_cla16_and1471_y0;
  wire h_s_cla16_and1472_y0;
  wire h_s_cla16_and1473_y0;
  wire h_s_cla16_and1474_y0;
  wire h_s_cla16_and1475_y0;
  wire h_s_cla16_and1476_y0;
  wire h_s_cla16_and1477_y0;
  wire h_s_cla16_and1478_y0;
  wire h_s_cla16_and1479_y0;
  wire h_s_cla16_and1480_y0;
  wire h_s_cla16_and1481_y0;
  wire h_s_cla16_and1482_y0;
  wire h_s_cla16_and1483_y0;
  wire h_s_cla16_and1484_y0;
  wire h_s_cla16_and1485_y0;
  wire h_s_cla16_and1486_y0;
  wire h_s_cla16_and1487_y0;
  wire h_s_cla16_and1488_y0;
  wire h_s_cla16_and1489_y0;
  wire h_s_cla16_and1490_y0;
  wire h_s_cla16_and1491_y0;
  wire h_s_cla16_and1492_y0;
  wire h_s_cla16_and1493_y0;
  wire h_s_cla16_and1494_y0;
  wire h_s_cla16_and1495_y0;
  wire h_s_cla16_or120_y0;
  wire h_s_cla16_or121_y0;
  wire h_s_cla16_or122_y0;
  wire h_s_cla16_or123_y0;
  wire h_s_cla16_or124_y0;
  wire h_s_cla16_or125_y0;
  wire h_s_cla16_or126_y0;
  wire h_s_cla16_or127_y0;
  wire h_s_cla16_or128_y0;
  wire h_s_cla16_or129_y0;
  wire h_s_cla16_or130_y0;
  wire h_s_cla16_or131_y0;
  wire h_s_cla16_or132_y0;
  wire h_s_cla16_or133_y0;
  wire h_s_cla16_or134_y0;
  wire h_s_cla16_or135_y0;
  wire h_s_cla16_xor16_y0;
  wire h_s_cla16_xor17_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  constant_wire_value_0 constant_wire_value_0_constant_wire_0(a_0, b_0, constant_wire_0);
  pg_logic pg_logic_h_s_cla16_pg_logic0_y0(a_0, b_0, h_s_cla16_pg_logic0_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_pg_logic0_y2);
  xor_gate xor_gate_h_s_cla16_xor0_y0(h_s_cla16_pg_logic0_y2, constant_wire_0, h_s_cla16_xor0_y0);
  and_gate and_gate_h_s_cla16_and0_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and0_y0);
  or_gate or_gate_h_s_cla16_or0_y0(h_s_cla16_pg_logic0_y1, h_s_cla16_and0_y0, h_s_cla16_or0_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic1_y0(a_1, b_1, h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_pg_logic1_y2);
  xor_gate xor_gate_h_s_cla16_xor1_y0(h_s_cla16_pg_logic1_y2, h_s_cla16_or0_y0, h_s_cla16_xor1_y0);
  and_gate and_gate_h_s_cla16_and1_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and1_y0);
  and_gate and_gate_h_s_cla16_and2_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and2_y0);
  and_gate and_gate_h_s_cla16_and3_y0(h_s_cla16_and2_y0, h_s_cla16_and1_y0, h_s_cla16_and3_y0);
  and_gate and_gate_h_s_cla16_and4_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and4_y0);
  or_gate or_gate_h_s_cla16_or1_y0(h_s_cla16_and4_y0, h_s_cla16_and3_y0, h_s_cla16_or1_y0);
  or_gate or_gate_h_s_cla16_or2_y0(h_s_cla16_pg_logic1_y1, h_s_cla16_or1_y0, h_s_cla16_or2_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic2_y0(a_2, b_2, h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_pg_logic2_y2);
  xor_gate xor_gate_h_s_cla16_xor2_y0(h_s_cla16_pg_logic2_y2, h_s_cla16_or2_y0, h_s_cla16_xor2_y0);
  and_gate and_gate_h_s_cla16_and5_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and5_y0);
  and_gate and_gate_h_s_cla16_and6_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and6_y0);
  and_gate and_gate_h_s_cla16_and7_y0(h_s_cla16_and6_y0, h_s_cla16_and5_y0, h_s_cla16_and7_y0);
  and_gate and_gate_h_s_cla16_and8_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and8_y0);
  and_gate and_gate_h_s_cla16_and9_y0(h_s_cla16_and8_y0, h_s_cla16_and7_y0, h_s_cla16_and9_y0);
  and_gate and_gate_h_s_cla16_and10_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and10_y0);
  and_gate and_gate_h_s_cla16_and11_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and11_y0);
  and_gate and_gate_h_s_cla16_and12_y0(h_s_cla16_and11_y0, h_s_cla16_and10_y0, h_s_cla16_and12_y0);
  and_gate and_gate_h_s_cla16_and13_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and13_y0);
  or_gate or_gate_h_s_cla16_or3_y0(h_s_cla16_and13_y0, h_s_cla16_and9_y0, h_s_cla16_or3_y0);
  or_gate or_gate_h_s_cla16_or4_y0(h_s_cla16_or3_y0, h_s_cla16_and12_y0, h_s_cla16_or4_y0);
  or_gate or_gate_h_s_cla16_or5_y0(h_s_cla16_pg_logic2_y1, h_s_cla16_or4_y0, h_s_cla16_or5_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic3_y0(a_3, b_3, h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_pg_logic3_y2);
  xor_gate xor_gate_h_s_cla16_xor3_y0(h_s_cla16_pg_logic3_y2, h_s_cla16_or5_y0, h_s_cla16_xor3_y0);
  and_gate and_gate_h_s_cla16_and14_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and14_y0);
  and_gate and_gate_h_s_cla16_and15_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and15_y0);
  and_gate and_gate_h_s_cla16_and16_y0(h_s_cla16_and15_y0, h_s_cla16_and14_y0, h_s_cla16_and16_y0);
  and_gate and_gate_h_s_cla16_and17_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and17_y0);
  and_gate and_gate_h_s_cla16_and18_y0(h_s_cla16_and17_y0, h_s_cla16_and16_y0, h_s_cla16_and18_y0);
  and_gate and_gate_h_s_cla16_and19_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and19_y0);
  and_gate and_gate_h_s_cla16_and20_y0(h_s_cla16_and19_y0, h_s_cla16_and18_y0, h_s_cla16_and20_y0);
  and_gate and_gate_h_s_cla16_and21_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and21_y0);
  and_gate and_gate_h_s_cla16_and22_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and22_y0);
  and_gate and_gate_h_s_cla16_and23_y0(h_s_cla16_and22_y0, h_s_cla16_and21_y0, h_s_cla16_and23_y0);
  and_gate and_gate_h_s_cla16_and24_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and24_y0);
  and_gate and_gate_h_s_cla16_and25_y0(h_s_cla16_and24_y0, h_s_cla16_and23_y0, h_s_cla16_and25_y0);
  and_gate and_gate_h_s_cla16_and26_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and26_y0);
  and_gate and_gate_h_s_cla16_and27_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and27_y0);
  and_gate and_gate_h_s_cla16_and28_y0(h_s_cla16_and27_y0, h_s_cla16_and26_y0, h_s_cla16_and28_y0);
  and_gate and_gate_h_s_cla16_and29_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and29_y0);
  or_gate or_gate_h_s_cla16_or6_y0(h_s_cla16_and29_y0, h_s_cla16_and20_y0, h_s_cla16_or6_y0);
  or_gate or_gate_h_s_cla16_or7_y0(h_s_cla16_or6_y0, h_s_cla16_and25_y0, h_s_cla16_or7_y0);
  or_gate or_gate_h_s_cla16_or8_y0(h_s_cla16_or7_y0, h_s_cla16_and28_y0, h_s_cla16_or8_y0);
  or_gate or_gate_h_s_cla16_or9_y0(h_s_cla16_pg_logic3_y1, h_s_cla16_or8_y0, h_s_cla16_or9_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic4_y0(a_4, b_4, h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_pg_logic4_y2);
  xor_gate xor_gate_h_s_cla16_xor4_y0(h_s_cla16_pg_logic4_y2, h_s_cla16_or9_y0, h_s_cla16_xor4_y0);
  and_gate and_gate_h_s_cla16_and30_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and30_y0);
  and_gate and_gate_h_s_cla16_and31_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and31_y0);
  and_gate and_gate_h_s_cla16_and32_y0(h_s_cla16_and31_y0, h_s_cla16_and30_y0, h_s_cla16_and32_y0);
  and_gate and_gate_h_s_cla16_and33_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and33_y0);
  and_gate and_gate_h_s_cla16_and34_y0(h_s_cla16_and33_y0, h_s_cla16_and32_y0, h_s_cla16_and34_y0);
  and_gate and_gate_h_s_cla16_and35_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and35_y0);
  and_gate and_gate_h_s_cla16_and36_y0(h_s_cla16_and35_y0, h_s_cla16_and34_y0, h_s_cla16_and36_y0);
  and_gate and_gate_h_s_cla16_and37_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and37_y0);
  and_gate and_gate_h_s_cla16_and38_y0(h_s_cla16_and37_y0, h_s_cla16_and36_y0, h_s_cla16_and38_y0);
  and_gate and_gate_h_s_cla16_and39_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and39_y0);
  and_gate and_gate_h_s_cla16_and40_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and40_y0);
  and_gate and_gate_h_s_cla16_and41_y0(h_s_cla16_and40_y0, h_s_cla16_and39_y0, h_s_cla16_and41_y0);
  and_gate and_gate_h_s_cla16_and42_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and42_y0);
  and_gate and_gate_h_s_cla16_and43_y0(h_s_cla16_and42_y0, h_s_cla16_and41_y0, h_s_cla16_and43_y0);
  and_gate and_gate_h_s_cla16_and44_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and44_y0);
  and_gate and_gate_h_s_cla16_and45_y0(h_s_cla16_and44_y0, h_s_cla16_and43_y0, h_s_cla16_and45_y0);
  and_gate and_gate_h_s_cla16_and46_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and46_y0);
  and_gate and_gate_h_s_cla16_and47_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and47_y0);
  and_gate and_gate_h_s_cla16_and48_y0(h_s_cla16_and47_y0, h_s_cla16_and46_y0, h_s_cla16_and48_y0);
  and_gate and_gate_h_s_cla16_and49_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and49_y0);
  and_gate and_gate_h_s_cla16_and50_y0(h_s_cla16_and49_y0, h_s_cla16_and48_y0, h_s_cla16_and50_y0);
  and_gate and_gate_h_s_cla16_and51_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and51_y0);
  and_gate and_gate_h_s_cla16_and52_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and52_y0);
  and_gate and_gate_h_s_cla16_and53_y0(h_s_cla16_and52_y0, h_s_cla16_and51_y0, h_s_cla16_and53_y0);
  and_gate and_gate_h_s_cla16_and54_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and54_y0);
  or_gate or_gate_h_s_cla16_or10_y0(h_s_cla16_and54_y0, h_s_cla16_and38_y0, h_s_cla16_or10_y0);
  or_gate or_gate_h_s_cla16_or11_y0(h_s_cla16_or10_y0, h_s_cla16_and45_y0, h_s_cla16_or11_y0);
  or_gate or_gate_h_s_cla16_or12_y0(h_s_cla16_or11_y0, h_s_cla16_and50_y0, h_s_cla16_or12_y0);
  or_gate or_gate_h_s_cla16_or13_y0(h_s_cla16_or12_y0, h_s_cla16_and53_y0, h_s_cla16_or13_y0);
  or_gate or_gate_h_s_cla16_or14_y0(h_s_cla16_pg_logic4_y1, h_s_cla16_or13_y0, h_s_cla16_or14_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic5_y0(a_5, b_5, h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_pg_logic5_y2);
  xor_gate xor_gate_h_s_cla16_xor5_y0(h_s_cla16_pg_logic5_y2, h_s_cla16_or14_y0, h_s_cla16_xor5_y0);
  and_gate and_gate_h_s_cla16_and55_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and55_y0);
  and_gate and_gate_h_s_cla16_and56_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and56_y0);
  and_gate and_gate_h_s_cla16_and57_y0(h_s_cla16_and56_y0, h_s_cla16_and55_y0, h_s_cla16_and57_y0);
  and_gate and_gate_h_s_cla16_and58_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and58_y0);
  and_gate and_gate_h_s_cla16_and59_y0(h_s_cla16_and58_y0, h_s_cla16_and57_y0, h_s_cla16_and59_y0);
  and_gate and_gate_h_s_cla16_and60_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and60_y0);
  and_gate and_gate_h_s_cla16_and61_y0(h_s_cla16_and60_y0, h_s_cla16_and59_y0, h_s_cla16_and61_y0);
  and_gate and_gate_h_s_cla16_and62_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and62_y0);
  and_gate and_gate_h_s_cla16_and63_y0(h_s_cla16_and62_y0, h_s_cla16_and61_y0, h_s_cla16_and63_y0);
  and_gate and_gate_h_s_cla16_and64_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and64_y0);
  and_gate and_gate_h_s_cla16_and65_y0(h_s_cla16_and64_y0, h_s_cla16_and63_y0, h_s_cla16_and65_y0);
  and_gate and_gate_h_s_cla16_and66_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and66_y0);
  and_gate and_gate_h_s_cla16_and67_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and67_y0);
  and_gate and_gate_h_s_cla16_and68_y0(h_s_cla16_and67_y0, h_s_cla16_and66_y0, h_s_cla16_and68_y0);
  and_gate and_gate_h_s_cla16_and69_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and69_y0);
  and_gate and_gate_h_s_cla16_and70_y0(h_s_cla16_and69_y0, h_s_cla16_and68_y0, h_s_cla16_and70_y0);
  and_gate and_gate_h_s_cla16_and71_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and71_y0);
  and_gate and_gate_h_s_cla16_and72_y0(h_s_cla16_and71_y0, h_s_cla16_and70_y0, h_s_cla16_and72_y0);
  and_gate and_gate_h_s_cla16_and73_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and73_y0);
  and_gate and_gate_h_s_cla16_and74_y0(h_s_cla16_and73_y0, h_s_cla16_and72_y0, h_s_cla16_and74_y0);
  and_gate and_gate_h_s_cla16_and75_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and75_y0);
  and_gate and_gate_h_s_cla16_and76_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and76_y0);
  and_gate and_gate_h_s_cla16_and77_y0(h_s_cla16_and76_y0, h_s_cla16_and75_y0, h_s_cla16_and77_y0);
  and_gate and_gate_h_s_cla16_and78_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and78_y0);
  and_gate and_gate_h_s_cla16_and79_y0(h_s_cla16_and78_y0, h_s_cla16_and77_y0, h_s_cla16_and79_y0);
  and_gate and_gate_h_s_cla16_and80_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and80_y0);
  and_gate and_gate_h_s_cla16_and81_y0(h_s_cla16_and80_y0, h_s_cla16_and79_y0, h_s_cla16_and81_y0);
  and_gate and_gate_h_s_cla16_and82_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and82_y0);
  and_gate and_gate_h_s_cla16_and83_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and83_y0);
  and_gate and_gate_h_s_cla16_and84_y0(h_s_cla16_and83_y0, h_s_cla16_and82_y0, h_s_cla16_and84_y0);
  and_gate and_gate_h_s_cla16_and85_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and85_y0);
  and_gate and_gate_h_s_cla16_and86_y0(h_s_cla16_and85_y0, h_s_cla16_and84_y0, h_s_cla16_and86_y0);
  and_gate and_gate_h_s_cla16_and87_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and87_y0);
  and_gate and_gate_h_s_cla16_and88_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and88_y0);
  and_gate and_gate_h_s_cla16_and89_y0(h_s_cla16_and88_y0, h_s_cla16_and87_y0, h_s_cla16_and89_y0);
  and_gate and_gate_h_s_cla16_and90_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and90_y0);
  or_gate or_gate_h_s_cla16_or15_y0(h_s_cla16_and90_y0, h_s_cla16_and65_y0, h_s_cla16_or15_y0);
  or_gate or_gate_h_s_cla16_or16_y0(h_s_cla16_or15_y0, h_s_cla16_and74_y0, h_s_cla16_or16_y0);
  or_gate or_gate_h_s_cla16_or17_y0(h_s_cla16_or16_y0, h_s_cla16_and81_y0, h_s_cla16_or17_y0);
  or_gate or_gate_h_s_cla16_or18_y0(h_s_cla16_or17_y0, h_s_cla16_and86_y0, h_s_cla16_or18_y0);
  or_gate or_gate_h_s_cla16_or19_y0(h_s_cla16_or18_y0, h_s_cla16_and89_y0, h_s_cla16_or19_y0);
  or_gate or_gate_h_s_cla16_or20_y0(h_s_cla16_pg_logic5_y1, h_s_cla16_or19_y0, h_s_cla16_or20_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic6_y0(a_6, b_6, h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_pg_logic6_y2);
  xor_gate xor_gate_h_s_cla16_xor6_y0(h_s_cla16_pg_logic6_y2, h_s_cla16_or20_y0, h_s_cla16_xor6_y0);
  and_gate and_gate_h_s_cla16_and91_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and91_y0);
  and_gate and_gate_h_s_cla16_and92_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and92_y0);
  and_gate and_gate_h_s_cla16_and93_y0(h_s_cla16_and92_y0, h_s_cla16_and91_y0, h_s_cla16_and93_y0);
  and_gate and_gate_h_s_cla16_and94_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and94_y0);
  and_gate and_gate_h_s_cla16_and95_y0(h_s_cla16_and94_y0, h_s_cla16_and93_y0, h_s_cla16_and95_y0);
  and_gate and_gate_h_s_cla16_and96_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and96_y0);
  and_gate and_gate_h_s_cla16_and97_y0(h_s_cla16_and96_y0, h_s_cla16_and95_y0, h_s_cla16_and97_y0);
  and_gate and_gate_h_s_cla16_and98_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and98_y0);
  and_gate and_gate_h_s_cla16_and99_y0(h_s_cla16_and98_y0, h_s_cla16_and97_y0, h_s_cla16_and99_y0);
  and_gate and_gate_h_s_cla16_and100_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and100_y0);
  and_gate and_gate_h_s_cla16_and101_y0(h_s_cla16_and100_y0, h_s_cla16_and99_y0, h_s_cla16_and101_y0);
  and_gate and_gate_h_s_cla16_and102_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and102_y0);
  and_gate and_gate_h_s_cla16_and103_y0(h_s_cla16_and102_y0, h_s_cla16_and101_y0, h_s_cla16_and103_y0);
  and_gate and_gate_h_s_cla16_and104_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and104_y0);
  and_gate and_gate_h_s_cla16_and105_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and105_y0);
  and_gate and_gate_h_s_cla16_and106_y0(h_s_cla16_and105_y0, h_s_cla16_and104_y0, h_s_cla16_and106_y0);
  and_gate and_gate_h_s_cla16_and107_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and107_y0);
  and_gate and_gate_h_s_cla16_and108_y0(h_s_cla16_and107_y0, h_s_cla16_and106_y0, h_s_cla16_and108_y0);
  and_gate and_gate_h_s_cla16_and109_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and109_y0);
  and_gate and_gate_h_s_cla16_and110_y0(h_s_cla16_and109_y0, h_s_cla16_and108_y0, h_s_cla16_and110_y0);
  and_gate and_gate_h_s_cla16_and111_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and111_y0);
  and_gate and_gate_h_s_cla16_and112_y0(h_s_cla16_and111_y0, h_s_cla16_and110_y0, h_s_cla16_and112_y0);
  and_gate and_gate_h_s_cla16_and113_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and113_y0);
  and_gate and_gate_h_s_cla16_and114_y0(h_s_cla16_and113_y0, h_s_cla16_and112_y0, h_s_cla16_and114_y0);
  and_gate and_gate_h_s_cla16_and115_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and115_y0);
  and_gate and_gate_h_s_cla16_and116_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and116_y0);
  and_gate and_gate_h_s_cla16_and117_y0(h_s_cla16_and116_y0, h_s_cla16_and115_y0, h_s_cla16_and117_y0);
  and_gate and_gate_h_s_cla16_and118_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and118_y0);
  and_gate and_gate_h_s_cla16_and119_y0(h_s_cla16_and118_y0, h_s_cla16_and117_y0, h_s_cla16_and119_y0);
  and_gate and_gate_h_s_cla16_and120_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and120_y0);
  and_gate and_gate_h_s_cla16_and121_y0(h_s_cla16_and120_y0, h_s_cla16_and119_y0, h_s_cla16_and121_y0);
  and_gate and_gate_h_s_cla16_and122_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and122_y0);
  and_gate and_gate_h_s_cla16_and123_y0(h_s_cla16_and122_y0, h_s_cla16_and121_y0, h_s_cla16_and123_y0);
  and_gate and_gate_h_s_cla16_and124_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and124_y0);
  and_gate and_gate_h_s_cla16_and125_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and125_y0);
  and_gate and_gate_h_s_cla16_and126_y0(h_s_cla16_and125_y0, h_s_cla16_and124_y0, h_s_cla16_and126_y0);
  and_gate and_gate_h_s_cla16_and127_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and127_y0);
  and_gate and_gate_h_s_cla16_and128_y0(h_s_cla16_and127_y0, h_s_cla16_and126_y0, h_s_cla16_and128_y0);
  and_gate and_gate_h_s_cla16_and129_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and129_y0);
  and_gate and_gate_h_s_cla16_and130_y0(h_s_cla16_and129_y0, h_s_cla16_and128_y0, h_s_cla16_and130_y0);
  and_gate and_gate_h_s_cla16_and131_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and131_y0);
  and_gate and_gate_h_s_cla16_and132_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and132_y0);
  and_gate and_gate_h_s_cla16_and133_y0(h_s_cla16_and132_y0, h_s_cla16_and131_y0, h_s_cla16_and133_y0);
  and_gate and_gate_h_s_cla16_and134_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and134_y0);
  and_gate and_gate_h_s_cla16_and135_y0(h_s_cla16_and134_y0, h_s_cla16_and133_y0, h_s_cla16_and135_y0);
  and_gate and_gate_h_s_cla16_and136_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and136_y0);
  and_gate and_gate_h_s_cla16_and137_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and137_y0);
  and_gate and_gate_h_s_cla16_and138_y0(h_s_cla16_and137_y0, h_s_cla16_and136_y0, h_s_cla16_and138_y0);
  and_gate and_gate_h_s_cla16_and139_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and139_y0);
  or_gate or_gate_h_s_cla16_or21_y0(h_s_cla16_and139_y0, h_s_cla16_and103_y0, h_s_cla16_or21_y0);
  or_gate or_gate_h_s_cla16_or22_y0(h_s_cla16_or21_y0, h_s_cla16_and114_y0, h_s_cla16_or22_y0);
  or_gate or_gate_h_s_cla16_or23_y0(h_s_cla16_or22_y0, h_s_cla16_and123_y0, h_s_cla16_or23_y0);
  or_gate or_gate_h_s_cla16_or24_y0(h_s_cla16_or23_y0, h_s_cla16_and130_y0, h_s_cla16_or24_y0);
  or_gate or_gate_h_s_cla16_or25_y0(h_s_cla16_or24_y0, h_s_cla16_and135_y0, h_s_cla16_or25_y0);
  or_gate or_gate_h_s_cla16_or26_y0(h_s_cla16_or25_y0, h_s_cla16_and138_y0, h_s_cla16_or26_y0);
  or_gate or_gate_h_s_cla16_or27_y0(h_s_cla16_pg_logic6_y1, h_s_cla16_or26_y0, h_s_cla16_or27_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic7_y0(a_7, b_7, h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_pg_logic7_y2);
  xor_gate xor_gate_h_s_cla16_xor7_y0(h_s_cla16_pg_logic7_y2, h_s_cla16_or27_y0, h_s_cla16_xor7_y0);
  and_gate and_gate_h_s_cla16_and140_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and140_y0);
  and_gate and_gate_h_s_cla16_and141_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and141_y0);
  and_gate and_gate_h_s_cla16_and142_y0(h_s_cla16_and141_y0, h_s_cla16_and140_y0, h_s_cla16_and142_y0);
  and_gate and_gate_h_s_cla16_and143_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and143_y0);
  and_gate and_gate_h_s_cla16_and144_y0(h_s_cla16_and143_y0, h_s_cla16_and142_y0, h_s_cla16_and144_y0);
  and_gate and_gate_h_s_cla16_and145_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and145_y0);
  and_gate and_gate_h_s_cla16_and146_y0(h_s_cla16_and145_y0, h_s_cla16_and144_y0, h_s_cla16_and146_y0);
  and_gate and_gate_h_s_cla16_and147_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and147_y0);
  and_gate and_gate_h_s_cla16_and148_y0(h_s_cla16_and147_y0, h_s_cla16_and146_y0, h_s_cla16_and148_y0);
  and_gate and_gate_h_s_cla16_and149_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and149_y0);
  and_gate and_gate_h_s_cla16_and150_y0(h_s_cla16_and149_y0, h_s_cla16_and148_y0, h_s_cla16_and150_y0);
  and_gate and_gate_h_s_cla16_and151_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and151_y0);
  and_gate and_gate_h_s_cla16_and152_y0(h_s_cla16_and151_y0, h_s_cla16_and150_y0, h_s_cla16_and152_y0);
  and_gate and_gate_h_s_cla16_and153_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and153_y0);
  and_gate and_gate_h_s_cla16_and154_y0(h_s_cla16_and153_y0, h_s_cla16_and152_y0, h_s_cla16_and154_y0);
  and_gate and_gate_h_s_cla16_and155_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and155_y0);
  and_gate and_gate_h_s_cla16_and156_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and156_y0);
  and_gate and_gate_h_s_cla16_and157_y0(h_s_cla16_and156_y0, h_s_cla16_and155_y0, h_s_cla16_and157_y0);
  and_gate and_gate_h_s_cla16_and158_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and158_y0);
  and_gate and_gate_h_s_cla16_and159_y0(h_s_cla16_and158_y0, h_s_cla16_and157_y0, h_s_cla16_and159_y0);
  and_gate and_gate_h_s_cla16_and160_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and160_y0);
  and_gate and_gate_h_s_cla16_and161_y0(h_s_cla16_and160_y0, h_s_cla16_and159_y0, h_s_cla16_and161_y0);
  and_gate and_gate_h_s_cla16_and162_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and162_y0);
  and_gate and_gate_h_s_cla16_and163_y0(h_s_cla16_and162_y0, h_s_cla16_and161_y0, h_s_cla16_and163_y0);
  and_gate and_gate_h_s_cla16_and164_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and164_y0);
  and_gate and_gate_h_s_cla16_and165_y0(h_s_cla16_and164_y0, h_s_cla16_and163_y0, h_s_cla16_and165_y0);
  and_gate and_gate_h_s_cla16_and166_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and166_y0);
  and_gate and_gate_h_s_cla16_and167_y0(h_s_cla16_and166_y0, h_s_cla16_and165_y0, h_s_cla16_and167_y0);
  and_gate and_gate_h_s_cla16_and168_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and168_y0);
  and_gate and_gate_h_s_cla16_and169_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and169_y0);
  and_gate and_gate_h_s_cla16_and170_y0(h_s_cla16_and169_y0, h_s_cla16_and168_y0, h_s_cla16_and170_y0);
  and_gate and_gate_h_s_cla16_and171_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and171_y0);
  and_gate and_gate_h_s_cla16_and172_y0(h_s_cla16_and171_y0, h_s_cla16_and170_y0, h_s_cla16_and172_y0);
  and_gate and_gate_h_s_cla16_and173_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and173_y0);
  and_gate and_gate_h_s_cla16_and174_y0(h_s_cla16_and173_y0, h_s_cla16_and172_y0, h_s_cla16_and174_y0);
  and_gate and_gate_h_s_cla16_and175_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and175_y0);
  and_gate and_gate_h_s_cla16_and176_y0(h_s_cla16_and175_y0, h_s_cla16_and174_y0, h_s_cla16_and176_y0);
  and_gate and_gate_h_s_cla16_and177_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and177_y0);
  and_gate and_gate_h_s_cla16_and178_y0(h_s_cla16_and177_y0, h_s_cla16_and176_y0, h_s_cla16_and178_y0);
  and_gate and_gate_h_s_cla16_and179_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and179_y0);
  and_gate and_gate_h_s_cla16_and180_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and180_y0);
  and_gate and_gate_h_s_cla16_and181_y0(h_s_cla16_and180_y0, h_s_cla16_and179_y0, h_s_cla16_and181_y0);
  and_gate and_gate_h_s_cla16_and182_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and182_y0);
  and_gate and_gate_h_s_cla16_and183_y0(h_s_cla16_and182_y0, h_s_cla16_and181_y0, h_s_cla16_and183_y0);
  and_gate and_gate_h_s_cla16_and184_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and184_y0);
  and_gate and_gate_h_s_cla16_and185_y0(h_s_cla16_and184_y0, h_s_cla16_and183_y0, h_s_cla16_and185_y0);
  and_gate and_gate_h_s_cla16_and186_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and186_y0);
  and_gate and_gate_h_s_cla16_and187_y0(h_s_cla16_and186_y0, h_s_cla16_and185_y0, h_s_cla16_and187_y0);
  and_gate and_gate_h_s_cla16_and188_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and188_y0);
  and_gate and_gate_h_s_cla16_and189_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and189_y0);
  and_gate and_gate_h_s_cla16_and190_y0(h_s_cla16_and189_y0, h_s_cla16_and188_y0, h_s_cla16_and190_y0);
  and_gate and_gate_h_s_cla16_and191_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and191_y0);
  and_gate and_gate_h_s_cla16_and192_y0(h_s_cla16_and191_y0, h_s_cla16_and190_y0, h_s_cla16_and192_y0);
  and_gate and_gate_h_s_cla16_and193_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and193_y0);
  and_gate and_gate_h_s_cla16_and194_y0(h_s_cla16_and193_y0, h_s_cla16_and192_y0, h_s_cla16_and194_y0);
  and_gate and_gate_h_s_cla16_and195_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and195_y0);
  and_gate and_gate_h_s_cla16_and196_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and196_y0);
  and_gate and_gate_h_s_cla16_and197_y0(h_s_cla16_and196_y0, h_s_cla16_and195_y0, h_s_cla16_and197_y0);
  and_gate and_gate_h_s_cla16_and198_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and198_y0);
  and_gate and_gate_h_s_cla16_and199_y0(h_s_cla16_and198_y0, h_s_cla16_and197_y0, h_s_cla16_and199_y0);
  and_gate and_gate_h_s_cla16_and200_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and200_y0);
  and_gate and_gate_h_s_cla16_and201_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and201_y0);
  and_gate and_gate_h_s_cla16_and202_y0(h_s_cla16_and201_y0, h_s_cla16_and200_y0, h_s_cla16_and202_y0);
  and_gate and_gate_h_s_cla16_and203_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and203_y0);
  or_gate or_gate_h_s_cla16_or28_y0(h_s_cla16_and203_y0, h_s_cla16_and154_y0, h_s_cla16_or28_y0);
  or_gate or_gate_h_s_cla16_or29_y0(h_s_cla16_or28_y0, h_s_cla16_and167_y0, h_s_cla16_or29_y0);
  or_gate or_gate_h_s_cla16_or30_y0(h_s_cla16_or29_y0, h_s_cla16_and178_y0, h_s_cla16_or30_y0);
  or_gate or_gate_h_s_cla16_or31_y0(h_s_cla16_or30_y0, h_s_cla16_and187_y0, h_s_cla16_or31_y0);
  or_gate or_gate_h_s_cla16_or32_y0(h_s_cla16_or31_y0, h_s_cla16_and194_y0, h_s_cla16_or32_y0);
  or_gate or_gate_h_s_cla16_or33_y0(h_s_cla16_or32_y0, h_s_cla16_and199_y0, h_s_cla16_or33_y0);
  or_gate or_gate_h_s_cla16_or34_y0(h_s_cla16_or33_y0, h_s_cla16_and202_y0, h_s_cla16_or34_y0);
  or_gate or_gate_h_s_cla16_or35_y0(h_s_cla16_pg_logic7_y1, h_s_cla16_or34_y0, h_s_cla16_or35_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic8_y0(a_8, b_8, h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_pg_logic8_y2);
  xor_gate xor_gate_h_s_cla16_xor8_y0(h_s_cla16_pg_logic8_y2, h_s_cla16_or35_y0, h_s_cla16_xor8_y0);
  and_gate and_gate_h_s_cla16_and204_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and204_y0);
  and_gate and_gate_h_s_cla16_and205_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and205_y0);
  and_gate and_gate_h_s_cla16_and206_y0(h_s_cla16_and205_y0, h_s_cla16_and204_y0, h_s_cla16_and206_y0);
  and_gate and_gate_h_s_cla16_and207_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and207_y0);
  and_gate and_gate_h_s_cla16_and208_y0(h_s_cla16_and207_y0, h_s_cla16_and206_y0, h_s_cla16_and208_y0);
  and_gate and_gate_h_s_cla16_and209_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and209_y0);
  and_gate and_gate_h_s_cla16_and210_y0(h_s_cla16_and209_y0, h_s_cla16_and208_y0, h_s_cla16_and210_y0);
  and_gate and_gate_h_s_cla16_and211_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and211_y0);
  and_gate and_gate_h_s_cla16_and212_y0(h_s_cla16_and211_y0, h_s_cla16_and210_y0, h_s_cla16_and212_y0);
  and_gate and_gate_h_s_cla16_and213_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and213_y0);
  and_gate and_gate_h_s_cla16_and214_y0(h_s_cla16_and213_y0, h_s_cla16_and212_y0, h_s_cla16_and214_y0);
  and_gate and_gate_h_s_cla16_and215_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and215_y0);
  and_gate and_gate_h_s_cla16_and216_y0(h_s_cla16_and215_y0, h_s_cla16_and214_y0, h_s_cla16_and216_y0);
  and_gate and_gate_h_s_cla16_and217_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and217_y0);
  and_gate and_gate_h_s_cla16_and218_y0(h_s_cla16_and217_y0, h_s_cla16_and216_y0, h_s_cla16_and218_y0);
  and_gate and_gate_h_s_cla16_and219_y0(h_s_cla16_pg_logic8_y0, constant_wire_0, h_s_cla16_and219_y0);
  and_gate and_gate_h_s_cla16_and220_y0(h_s_cla16_and219_y0, h_s_cla16_and218_y0, h_s_cla16_and220_y0);
  and_gate and_gate_h_s_cla16_and221_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and221_y0);
  and_gate and_gate_h_s_cla16_and222_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and222_y0);
  and_gate and_gate_h_s_cla16_and223_y0(h_s_cla16_and222_y0, h_s_cla16_and221_y0, h_s_cla16_and223_y0);
  and_gate and_gate_h_s_cla16_and224_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and224_y0);
  and_gate and_gate_h_s_cla16_and225_y0(h_s_cla16_and224_y0, h_s_cla16_and223_y0, h_s_cla16_and225_y0);
  and_gate and_gate_h_s_cla16_and226_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and226_y0);
  and_gate and_gate_h_s_cla16_and227_y0(h_s_cla16_and226_y0, h_s_cla16_and225_y0, h_s_cla16_and227_y0);
  and_gate and_gate_h_s_cla16_and228_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and228_y0);
  and_gate and_gate_h_s_cla16_and229_y0(h_s_cla16_and228_y0, h_s_cla16_and227_y0, h_s_cla16_and229_y0);
  and_gate and_gate_h_s_cla16_and230_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and230_y0);
  and_gate and_gate_h_s_cla16_and231_y0(h_s_cla16_and230_y0, h_s_cla16_and229_y0, h_s_cla16_and231_y0);
  and_gate and_gate_h_s_cla16_and232_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and232_y0);
  and_gate and_gate_h_s_cla16_and233_y0(h_s_cla16_and232_y0, h_s_cla16_and231_y0, h_s_cla16_and233_y0);
  and_gate and_gate_h_s_cla16_and234_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and234_y0);
  and_gate and_gate_h_s_cla16_and235_y0(h_s_cla16_and234_y0, h_s_cla16_and233_y0, h_s_cla16_and235_y0);
  and_gate and_gate_h_s_cla16_and236_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and236_y0);
  and_gate and_gate_h_s_cla16_and237_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and237_y0);
  and_gate and_gate_h_s_cla16_and238_y0(h_s_cla16_and237_y0, h_s_cla16_and236_y0, h_s_cla16_and238_y0);
  and_gate and_gate_h_s_cla16_and239_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and239_y0);
  and_gate and_gate_h_s_cla16_and240_y0(h_s_cla16_and239_y0, h_s_cla16_and238_y0, h_s_cla16_and240_y0);
  and_gate and_gate_h_s_cla16_and241_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and241_y0);
  and_gate and_gate_h_s_cla16_and242_y0(h_s_cla16_and241_y0, h_s_cla16_and240_y0, h_s_cla16_and242_y0);
  and_gate and_gate_h_s_cla16_and243_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and243_y0);
  and_gate and_gate_h_s_cla16_and244_y0(h_s_cla16_and243_y0, h_s_cla16_and242_y0, h_s_cla16_and244_y0);
  and_gate and_gate_h_s_cla16_and245_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and245_y0);
  and_gate and_gate_h_s_cla16_and246_y0(h_s_cla16_and245_y0, h_s_cla16_and244_y0, h_s_cla16_and246_y0);
  and_gate and_gate_h_s_cla16_and247_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and247_y0);
  and_gate and_gate_h_s_cla16_and248_y0(h_s_cla16_and247_y0, h_s_cla16_and246_y0, h_s_cla16_and248_y0);
  and_gate and_gate_h_s_cla16_and249_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and249_y0);
  and_gate and_gate_h_s_cla16_and250_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and250_y0);
  and_gate and_gate_h_s_cla16_and251_y0(h_s_cla16_and250_y0, h_s_cla16_and249_y0, h_s_cla16_and251_y0);
  and_gate and_gate_h_s_cla16_and252_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and252_y0);
  and_gate and_gate_h_s_cla16_and253_y0(h_s_cla16_and252_y0, h_s_cla16_and251_y0, h_s_cla16_and253_y0);
  and_gate and_gate_h_s_cla16_and254_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and254_y0);
  and_gate and_gate_h_s_cla16_and255_y0(h_s_cla16_and254_y0, h_s_cla16_and253_y0, h_s_cla16_and255_y0);
  and_gate and_gate_h_s_cla16_and256_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and256_y0);
  and_gate and_gate_h_s_cla16_and257_y0(h_s_cla16_and256_y0, h_s_cla16_and255_y0, h_s_cla16_and257_y0);
  and_gate and_gate_h_s_cla16_and258_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and258_y0);
  and_gate and_gate_h_s_cla16_and259_y0(h_s_cla16_and258_y0, h_s_cla16_and257_y0, h_s_cla16_and259_y0);
  and_gate and_gate_h_s_cla16_and260_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and260_y0);
  and_gate and_gate_h_s_cla16_and261_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and261_y0);
  and_gate and_gate_h_s_cla16_and262_y0(h_s_cla16_and261_y0, h_s_cla16_and260_y0, h_s_cla16_and262_y0);
  and_gate and_gate_h_s_cla16_and263_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and263_y0);
  and_gate and_gate_h_s_cla16_and264_y0(h_s_cla16_and263_y0, h_s_cla16_and262_y0, h_s_cla16_and264_y0);
  and_gate and_gate_h_s_cla16_and265_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and265_y0);
  and_gate and_gate_h_s_cla16_and266_y0(h_s_cla16_and265_y0, h_s_cla16_and264_y0, h_s_cla16_and266_y0);
  and_gate and_gate_h_s_cla16_and267_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and267_y0);
  and_gate and_gate_h_s_cla16_and268_y0(h_s_cla16_and267_y0, h_s_cla16_and266_y0, h_s_cla16_and268_y0);
  and_gate and_gate_h_s_cla16_and269_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and269_y0);
  and_gate and_gate_h_s_cla16_and270_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and270_y0);
  and_gate and_gate_h_s_cla16_and271_y0(h_s_cla16_and270_y0, h_s_cla16_and269_y0, h_s_cla16_and271_y0);
  and_gate and_gate_h_s_cla16_and272_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and272_y0);
  and_gate and_gate_h_s_cla16_and273_y0(h_s_cla16_and272_y0, h_s_cla16_and271_y0, h_s_cla16_and273_y0);
  and_gate and_gate_h_s_cla16_and274_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and274_y0);
  and_gate and_gate_h_s_cla16_and275_y0(h_s_cla16_and274_y0, h_s_cla16_and273_y0, h_s_cla16_and275_y0);
  and_gate and_gate_h_s_cla16_and276_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and276_y0);
  and_gate and_gate_h_s_cla16_and277_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and277_y0);
  and_gate and_gate_h_s_cla16_and278_y0(h_s_cla16_and277_y0, h_s_cla16_and276_y0, h_s_cla16_and278_y0);
  and_gate and_gate_h_s_cla16_and279_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and279_y0);
  and_gate and_gate_h_s_cla16_and280_y0(h_s_cla16_and279_y0, h_s_cla16_and278_y0, h_s_cla16_and280_y0);
  and_gate and_gate_h_s_cla16_and281_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and281_y0);
  and_gate and_gate_h_s_cla16_and282_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and282_y0);
  and_gate and_gate_h_s_cla16_and283_y0(h_s_cla16_and282_y0, h_s_cla16_and281_y0, h_s_cla16_and283_y0);
  and_gate and_gate_h_s_cla16_and284_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and284_y0);
  or_gate or_gate_h_s_cla16_or36_y0(h_s_cla16_and284_y0, h_s_cla16_and220_y0, h_s_cla16_or36_y0);
  or_gate or_gate_h_s_cla16_or37_y0(h_s_cla16_or36_y0, h_s_cla16_and235_y0, h_s_cla16_or37_y0);
  or_gate or_gate_h_s_cla16_or38_y0(h_s_cla16_or37_y0, h_s_cla16_and248_y0, h_s_cla16_or38_y0);
  or_gate or_gate_h_s_cla16_or39_y0(h_s_cla16_or38_y0, h_s_cla16_and259_y0, h_s_cla16_or39_y0);
  or_gate or_gate_h_s_cla16_or40_y0(h_s_cla16_or39_y0, h_s_cla16_and268_y0, h_s_cla16_or40_y0);
  or_gate or_gate_h_s_cla16_or41_y0(h_s_cla16_or40_y0, h_s_cla16_and275_y0, h_s_cla16_or41_y0);
  or_gate or_gate_h_s_cla16_or42_y0(h_s_cla16_or41_y0, h_s_cla16_and280_y0, h_s_cla16_or42_y0);
  or_gate or_gate_h_s_cla16_or43_y0(h_s_cla16_or42_y0, h_s_cla16_and283_y0, h_s_cla16_or43_y0);
  or_gate or_gate_h_s_cla16_or44_y0(h_s_cla16_pg_logic8_y1, h_s_cla16_or43_y0, h_s_cla16_or44_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic9_y0(a_9, b_9, h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_pg_logic9_y2);
  xor_gate xor_gate_h_s_cla16_xor9_y0(h_s_cla16_pg_logic9_y2, h_s_cla16_or44_y0, h_s_cla16_xor9_y0);
  and_gate and_gate_h_s_cla16_and285_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and285_y0);
  and_gate and_gate_h_s_cla16_and286_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and286_y0);
  and_gate and_gate_h_s_cla16_and287_y0(h_s_cla16_and286_y0, h_s_cla16_and285_y0, h_s_cla16_and287_y0);
  and_gate and_gate_h_s_cla16_and288_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and288_y0);
  and_gate and_gate_h_s_cla16_and289_y0(h_s_cla16_and288_y0, h_s_cla16_and287_y0, h_s_cla16_and289_y0);
  and_gate and_gate_h_s_cla16_and290_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and290_y0);
  and_gate and_gate_h_s_cla16_and291_y0(h_s_cla16_and290_y0, h_s_cla16_and289_y0, h_s_cla16_and291_y0);
  and_gate and_gate_h_s_cla16_and292_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and292_y0);
  and_gate and_gate_h_s_cla16_and293_y0(h_s_cla16_and292_y0, h_s_cla16_and291_y0, h_s_cla16_and293_y0);
  and_gate and_gate_h_s_cla16_and294_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and294_y0);
  and_gate and_gate_h_s_cla16_and295_y0(h_s_cla16_and294_y0, h_s_cla16_and293_y0, h_s_cla16_and295_y0);
  and_gate and_gate_h_s_cla16_and296_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and296_y0);
  and_gate and_gate_h_s_cla16_and297_y0(h_s_cla16_and296_y0, h_s_cla16_and295_y0, h_s_cla16_and297_y0);
  and_gate and_gate_h_s_cla16_and298_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and298_y0);
  and_gate and_gate_h_s_cla16_and299_y0(h_s_cla16_and298_y0, h_s_cla16_and297_y0, h_s_cla16_and299_y0);
  and_gate and_gate_h_s_cla16_and300_y0(h_s_cla16_pg_logic8_y0, constant_wire_0, h_s_cla16_and300_y0);
  and_gate and_gate_h_s_cla16_and301_y0(h_s_cla16_and300_y0, h_s_cla16_and299_y0, h_s_cla16_and301_y0);
  and_gate and_gate_h_s_cla16_and302_y0(h_s_cla16_pg_logic9_y0, constant_wire_0, h_s_cla16_and302_y0);
  and_gate and_gate_h_s_cla16_and303_y0(h_s_cla16_and302_y0, h_s_cla16_and301_y0, h_s_cla16_and303_y0);
  and_gate and_gate_h_s_cla16_and304_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and304_y0);
  and_gate and_gate_h_s_cla16_and305_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and305_y0);
  and_gate and_gate_h_s_cla16_and306_y0(h_s_cla16_and305_y0, h_s_cla16_and304_y0, h_s_cla16_and306_y0);
  and_gate and_gate_h_s_cla16_and307_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and307_y0);
  and_gate and_gate_h_s_cla16_and308_y0(h_s_cla16_and307_y0, h_s_cla16_and306_y0, h_s_cla16_and308_y0);
  and_gate and_gate_h_s_cla16_and309_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and309_y0);
  and_gate and_gate_h_s_cla16_and310_y0(h_s_cla16_and309_y0, h_s_cla16_and308_y0, h_s_cla16_and310_y0);
  and_gate and_gate_h_s_cla16_and311_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and311_y0);
  and_gate and_gate_h_s_cla16_and312_y0(h_s_cla16_and311_y0, h_s_cla16_and310_y0, h_s_cla16_and312_y0);
  and_gate and_gate_h_s_cla16_and313_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and313_y0);
  and_gate and_gate_h_s_cla16_and314_y0(h_s_cla16_and313_y0, h_s_cla16_and312_y0, h_s_cla16_and314_y0);
  and_gate and_gate_h_s_cla16_and315_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and315_y0);
  and_gate and_gate_h_s_cla16_and316_y0(h_s_cla16_and315_y0, h_s_cla16_and314_y0, h_s_cla16_and316_y0);
  and_gate and_gate_h_s_cla16_and317_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and317_y0);
  and_gate and_gate_h_s_cla16_and318_y0(h_s_cla16_and317_y0, h_s_cla16_and316_y0, h_s_cla16_and318_y0);
  and_gate and_gate_h_s_cla16_and319_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and319_y0);
  and_gate and_gate_h_s_cla16_and320_y0(h_s_cla16_and319_y0, h_s_cla16_and318_y0, h_s_cla16_and320_y0);
  and_gate and_gate_h_s_cla16_and321_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and321_y0);
  and_gate and_gate_h_s_cla16_and322_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and322_y0);
  and_gate and_gate_h_s_cla16_and323_y0(h_s_cla16_and322_y0, h_s_cla16_and321_y0, h_s_cla16_and323_y0);
  and_gate and_gate_h_s_cla16_and324_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and324_y0);
  and_gate and_gate_h_s_cla16_and325_y0(h_s_cla16_and324_y0, h_s_cla16_and323_y0, h_s_cla16_and325_y0);
  and_gate and_gate_h_s_cla16_and326_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and326_y0);
  and_gate and_gate_h_s_cla16_and327_y0(h_s_cla16_and326_y0, h_s_cla16_and325_y0, h_s_cla16_and327_y0);
  and_gate and_gate_h_s_cla16_and328_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and328_y0);
  and_gate and_gate_h_s_cla16_and329_y0(h_s_cla16_and328_y0, h_s_cla16_and327_y0, h_s_cla16_and329_y0);
  and_gate and_gate_h_s_cla16_and330_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and330_y0);
  and_gate and_gate_h_s_cla16_and331_y0(h_s_cla16_and330_y0, h_s_cla16_and329_y0, h_s_cla16_and331_y0);
  and_gate and_gate_h_s_cla16_and332_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and332_y0);
  and_gate and_gate_h_s_cla16_and333_y0(h_s_cla16_and332_y0, h_s_cla16_and331_y0, h_s_cla16_and333_y0);
  and_gate and_gate_h_s_cla16_and334_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and334_y0);
  and_gate and_gate_h_s_cla16_and335_y0(h_s_cla16_and334_y0, h_s_cla16_and333_y0, h_s_cla16_and335_y0);
  and_gate and_gate_h_s_cla16_and336_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and336_y0);
  and_gate and_gate_h_s_cla16_and337_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and337_y0);
  and_gate and_gate_h_s_cla16_and338_y0(h_s_cla16_and337_y0, h_s_cla16_and336_y0, h_s_cla16_and338_y0);
  and_gate and_gate_h_s_cla16_and339_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and339_y0);
  and_gate and_gate_h_s_cla16_and340_y0(h_s_cla16_and339_y0, h_s_cla16_and338_y0, h_s_cla16_and340_y0);
  and_gate and_gate_h_s_cla16_and341_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and341_y0);
  and_gate and_gate_h_s_cla16_and342_y0(h_s_cla16_and341_y0, h_s_cla16_and340_y0, h_s_cla16_and342_y0);
  and_gate and_gate_h_s_cla16_and343_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and343_y0);
  and_gate and_gate_h_s_cla16_and344_y0(h_s_cla16_and343_y0, h_s_cla16_and342_y0, h_s_cla16_and344_y0);
  and_gate and_gate_h_s_cla16_and345_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and345_y0);
  and_gate and_gate_h_s_cla16_and346_y0(h_s_cla16_and345_y0, h_s_cla16_and344_y0, h_s_cla16_and346_y0);
  and_gate and_gate_h_s_cla16_and347_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and347_y0);
  and_gate and_gate_h_s_cla16_and348_y0(h_s_cla16_and347_y0, h_s_cla16_and346_y0, h_s_cla16_and348_y0);
  and_gate and_gate_h_s_cla16_and349_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and349_y0);
  and_gate and_gate_h_s_cla16_and350_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and350_y0);
  and_gate and_gate_h_s_cla16_and351_y0(h_s_cla16_and350_y0, h_s_cla16_and349_y0, h_s_cla16_and351_y0);
  and_gate and_gate_h_s_cla16_and352_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and352_y0);
  and_gate and_gate_h_s_cla16_and353_y0(h_s_cla16_and352_y0, h_s_cla16_and351_y0, h_s_cla16_and353_y0);
  and_gate and_gate_h_s_cla16_and354_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and354_y0);
  and_gate and_gate_h_s_cla16_and355_y0(h_s_cla16_and354_y0, h_s_cla16_and353_y0, h_s_cla16_and355_y0);
  and_gate and_gate_h_s_cla16_and356_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and356_y0);
  and_gate and_gate_h_s_cla16_and357_y0(h_s_cla16_and356_y0, h_s_cla16_and355_y0, h_s_cla16_and357_y0);
  and_gate and_gate_h_s_cla16_and358_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and358_y0);
  and_gate and_gate_h_s_cla16_and359_y0(h_s_cla16_and358_y0, h_s_cla16_and357_y0, h_s_cla16_and359_y0);
  and_gate and_gate_h_s_cla16_and360_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and360_y0);
  and_gate and_gate_h_s_cla16_and361_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and361_y0);
  and_gate and_gate_h_s_cla16_and362_y0(h_s_cla16_and361_y0, h_s_cla16_and360_y0, h_s_cla16_and362_y0);
  and_gate and_gate_h_s_cla16_and363_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and363_y0);
  and_gate and_gate_h_s_cla16_and364_y0(h_s_cla16_and363_y0, h_s_cla16_and362_y0, h_s_cla16_and364_y0);
  and_gate and_gate_h_s_cla16_and365_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and365_y0);
  and_gate and_gate_h_s_cla16_and366_y0(h_s_cla16_and365_y0, h_s_cla16_and364_y0, h_s_cla16_and366_y0);
  and_gate and_gate_h_s_cla16_and367_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and367_y0);
  and_gate and_gate_h_s_cla16_and368_y0(h_s_cla16_and367_y0, h_s_cla16_and366_y0, h_s_cla16_and368_y0);
  and_gate and_gate_h_s_cla16_and369_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and369_y0);
  and_gate and_gate_h_s_cla16_and370_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and370_y0);
  and_gate and_gate_h_s_cla16_and371_y0(h_s_cla16_and370_y0, h_s_cla16_and369_y0, h_s_cla16_and371_y0);
  and_gate and_gate_h_s_cla16_and372_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and372_y0);
  and_gate and_gate_h_s_cla16_and373_y0(h_s_cla16_and372_y0, h_s_cla16_and371_y0, h_s_cla16_and373_y0);
  and_gate and_gate_h_s_cla16_and374_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and374_y0);
  and_gate and_gate_h_s_cla16_and375_y0(h_s_cla16_and374_y0, h_s_cla16_and373_y0, h_s_cla16_and375_y0);
  and_gate and_gate_h_s_cla16_and376_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and376_y0);
  and_gate and_gate_h_s_cla16_and377_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and377_y0);
  and_gate and_gate_h_s_cla16_and378_y0(h_s_cla16_and377_y0, h_s_cla16_and376_y0, h_s_cla16_and378_y0);
  and_gate and_gate_h_s_cla16_and379_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and379_y0);
  and_gate and_gate_h_s_cla16_and380_y0(h_s_cla16_and379_y0, h_s_cla16_and378_y0, h_s_cla16_and380_y0);
  and_gate and_gate_h_s_cla16_and381_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and381_y0);
  and_gate and_gate_h_s_cla16_and382_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and382_y0);
  and_gate and_gate_h_s_cla16_and383_y0(h_s_cla16_and382_y0, h_s_cla16_and381_y0, h_s_cla16_and383_y0);
  and_gate and_gate_h_s_cla16_and384_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and384_y0);
  or_gate or_gate_h_s_cla16_or45_y0(h_s_cla16_and384_y0, h_s_cla16_and303_y0, h_s_cla16_or45_y0);
  or_gate or_gate_h_s_cla16_or46_y0(h_s_cla16_or45_y0, h_s_cla16_and320_y0, h_s_cla16_or46_y0);
  or_gate or_gate_h_s_cla16_or47_y0(h_s_cla16_or46_y0, h_s_cla16_and335_y0, h_s_cla16_or47_y0);
  or_gate or_gate_h_s_cla16_or48_y0(h_s_cla16_or47_y0, h_s_cla16_and348_y0, h_s_cla16_or48_y0);
  or_gate or_gate_h_s_cla16_or49_y0(h_s_cla16_or48_y0, h_s_cla16_and359_y0, h_s_cla16_or49_y0);
  or_gate or_gate_h_s_cla16_or50_y0(h_s_cla16_or49_y0, h_s_cla16_and368_y0, h_s_cla16_or50_y0);
  or_gate or_gate_h_s_cla16_or51_y0(h_s_cla16_or50_y0, h_s_cla16_and375_y0, h_s_cla16_or51_y0);
  or_gate or_gate_h_s_cla16_or52_y0(h_s_cla16_or51_y0, h_s_cla16_and380_y0, h_s_cla16_or52_y0);
  or_gate or_gate_h_s_cla16_or53_y0(h_s_cla16_or52_y0, h_s_cla16_and383_y0, h_s_cla16_or53_y0);
  or_gate or_gate_h_s_cla16_or54_y0(h_s_cla16_pg_logic9_y1, h_s_cla16_or53_y0, h_s_cla16_or54_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic10_y0(a_10, b_10, h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_pg_logic10_y2);
  xor_gate xor_gate_h_s_cla16_xor10_y0(h_s_cla16_pg_logic10_y2, h_s_cla16_or54_y0, h_s_cla16_xor10_y0);
  and_gate and_gate_h_s_cla16_and385_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and385_y0);
  and_gate and_gate_h_s_cla16_and386_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and386_y0);
  and_gate and_gate_h_s_cla16_and387_y0(h_s_cla16_and386_y0, h_s_cla16_and385_y0, h_s_cla16_and387_y0);
  and_gate and_gate_h_s_cla16_and388_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and388_y0);
  and_gate and_gate_h_s_cla16_and389_y0(h_s_cla16_and388_y0, h_s_cla16_and387_y0, h_s_cla16_and389_y0);
  and_gate and_gate_h_s_cla16_and390_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and390_y0);
  and_gate and_gate_h_s_cla16_and391_y0(h_s_cla16_and390_y0, h_s_cla16_and389_y0, h_s_cla16_and391_y0);
  and_gate and_gate_h_s_cla16_and392_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and392_y0);
  and_gate and_gate_h_s_cla16_and393_y0(h_s_cla16_and392_y0, h_s_cla16_and391_y0, h_s_cla16_and393_y0);
  and_gate and_gate_h_s_cla16_and394_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and394_y0);
  and_gate and_gate_h_s_cla16_and395_y0(h_s_cla16_and394_y0, h_s_cla16_and393_y0, h_s_cla16_and395_y0);
  and_gate and_gate_h_s_cla16_and396_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and396_y0);
  and_gate and_gate_h_s_cla16_and397_y0(h_s_cla16_and396_y0, h_s_cla16_and395_y0, h_s_cla16_and397_y0);
  and_gate and_gate_h_s_cla16_and398_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and398_y0);
  and_gate and_gate_h_s_cla16_and399_y0(h_s_cla16_and398_y0, h_s_cla16_and397_y0, h_s_cla16_and399_y0);
  and_gate and_gate_h_s_cla16_and400_y0(h_s_cla16_pg_logic8_y0, constant_wire_0, h_s_cla16_and400_y0);
  and_gate and_gate_h_s_cla16_and401_y0(h_s_cla16_and400_y0, h_s_cla16_and399_y0, h_s_cla16_and401_y0);
  and_gate and_gate_h_s_cla16_and402_y0(h_s_cla16_pg_logic9_y0, constant_wire_0, h_s_cla16_and402_y0);
  and_gate and_gate_h_s_cla16_and403_y0(h_s_cla16_and402_y0, h_s_cla16_and401_y0, h_s_cla16_and403_y0);
  and_gate and_gate_h_s_cla16_and404_y0(h_s_cla16_pg_logic10_y0, constant_wire_0, h_s_cla16_and404_y0);
  and_gate and_gate_h_s_cla16_and405_y0(h_s_cla16_and404_y0, h_s_cla16_and403_y0, h_s_cla16_and405_y0);
  and_gate and_gate_h_s_cla16_and406_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and406_y0);
  and_gate and_gate_h_s_cla16_and407_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and407_y0);
  and_gate and_gate_h_s_cla16_and408_y0(h_s_cla16_and407_y0, h_s_cla16_and406_y0, h_s_cla16_and408_y0);
  and_gate and_gate_h_s_cla16_and409_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and409_y0);
  and_gate and_gate_h_s_cla16_and410_y0(h_s_cla16_and409_y0, h_s_cla16_and408_y0, h_s_cla16_and410_y0);
  and_gate and_gate_h_s_cla16_and411_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and411_y0);
  and_gate and_gate_h_s_cla16_and412_y0(h_s_cla16_and411_y0, h_s_cla16_and410_y0, h_s_cla16_and412_y0);
  and_gate and_gate_h_s_cla16_and413_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and413_y0);
  and_gate and_gate_h_s_cla16_and414_y0(h_s_cla16_and413_y0, h_s_cla16_and412_y0, h_s_cla16_and414_y0);
  and_gate and_gate_h_s_cla16_and415_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and415_y0);
  and_gate and_gate_h_s_cla16_and416_y0(h_s_cla16_and415_y0, h_s_cla16_and414_y0, h_s_cla16_and416_y0);
  and_gate and_gate_h_s_cla16_and417_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and417_y0);
  and_gate and_gate_h_s_cla16_and418_y0(h_s_cla16_and417_y0, h_s_cla16_and416_y0, h_s_cla16_and418_y0);
  and_gate and_gate_h_s_cla16_and419_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and419_y0);
  and_gate and_gate_h_s_cla16_and420_y0(h_s_cla16_and419_y0, h_s_cla16_and418_y0, h_s_cla16_and420_y0);
  and_gate and_gate_h_s_cla16_and421_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and421_y0);
  and_gate and_gate_h_s_cla16_and422_y0(h_s_cla16_and421_y0, h_s_cla16_and420_y0, h_s_cla16_and422_y0);
  and_gate and_gate_h_s_cla16_and423_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and423_y0);
  and_gate and_gate_h_s_cla16_and424_y0(h_s_cla16_and423_y0, h_s_cla16_and422_y0, h_s_cla16_and424_y0);
  and_gate and_gate_h_s_cla16_and425_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and425_y0);
  and_gate and_gate_h_s_cla16_and426_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and426_y0);
  and_gate and_gate_h_s_cla16_and427_y0(h_s_cla16_and426_y0, h_s_cla16_and425_y0, h_s_cla16_and427_y0);
  and_gate and_gate_h_s_cla16_and428_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and428_y0);
  and_gate and_gate_h_s_cla16_and429_y0(h_s_cla16_and428_y0, h_s_cla16_and427_y0, h_s_cla16_and429_y0);
  and_gate and_gate_h_s_cla16_and430_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and430_y0);
  and_gate and_gate_h_s_cla16_and431_y0(h_s_cla16_and430_y0, h_s_cla16_and429_y0, h_s_cla16_and431_y0);
  and_gate and_gate_h_s_cla16_and432_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and432_y0);
  and_gate and_gate_h_s_cla16_and433_y0(h_s_cla16_and432_y0, h_s_cla16_and431_y0, h_s_cla16_and433_y0);
  and_gate and_gate_h_s_cla16_and434_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and434_y0);
  and_gate and_gate_h_s_cla16_and435_y0(h_s_cla16_and434_y0, h_s_cla16_and433_y0, h_s_cla16_and435_y0);
  and_gate and_gate_h_s_cla16_and436_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and436_y0);
  and_gate and_gate_h_s_cla16_and437_y0(h_s_cla16_and436_y0, h_s_cla16_and435_y0, h_s_cla16_and437_y0);
  and_gate and_gate_h_s_cla16_and438_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and438_y0);
  and_gate and_gate_h_s_cla16_and439_y0(h_s_cla16_and438_y0, h_s_cla16_and437_y0, h_s_cla16_and439_y0);
  and_gate and_gate_h_s_cla16_and440_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and440_y0);
  and_gate and_gate_h_s_cla16_and441_y0(h_s_cla16_and440_y0, h_s_cla16_and439_y0, h_s_cla16_and441_y0);
  and_gate and_gate_h_s_cla16_and442_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and442_y0);
  and_gate and_gate_h_s_cla16_and443_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and443_y0);
  and_gate and_gate_h_s_cla16_and444_y0(h_s_cla16_and443_y0, h_s_cla16_and442_y0, h_s_cla16_and444_y0);
  and_gate and_gate_h_s_cla16_and445_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and445_y0);
  and_gate and_gate_h_s_cla16_and446_y0(h_s_cla16_and445_y0, h_s_cla16_and444_y0, h_s_cla16_and446_y0);
  and_gate and_gate_h_s_cla16_and447_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and447_y0);
  and_gate and_gate_h_s_cla16_and448_y0(h_s_cla16_and447_y0, h_s_cla16_and446_y0, h_s_cla16_and448_y0);
  and_gate and_gate_h_s_cla16_and449_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and449_y0);
  and_gate and_gate_h_s_cla16_and450_y0(h_s_cla16_and449_y0, h_s_cla16_and448_y0, h_s_cla16_and450_y0);
  and_gate and_gate_h_s_cla16_and451_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and451_y0);
  and_gate and_gate_h_s_cla16_and452_y0(h_s_cla16_and451_y0, h_s_cla16_and450_y0, h_s_cla16_and452_y0);
  and_gate and_gate_h_s_cla16_and453_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and453_y0);
  and_gate and_gate_h_s_cla16_and454_y0(h_s_cla16_and453_y0, h_s_cla16_and452_y0, h_s_cla16_and454_y0);
  and_gate and_gate_h_s_cla16_and455_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and455_y0);
  and_gate and_gate_h_s_cla16_and456_y0(h_s_cla16_and455_y0, h_s_cla16_and454_y0, h_s_cla16_and456_y0);
  and_gate and_gate_h_s_cla16_and457_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and457_y0);
  and_gate and_gate_h_s_cla16_and458_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and458_y0);
  and_gate and_gate_h_s_cla16_and459_y0(h_s_cla16_and458_y0, h_s_cla16_and457_y0, h_s_cla16_and459_y0);
  and_gate and_gate_h_s_cla16_and460_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and460_y0);
  and_gate and_gate_h_s_cla16_and461_y0(h_s_cla16_and460_y0, h_s_cla16_and459_y0, h_s_cla16_and461_y0);
  and_gate and_gate_h_s_cla16_and462_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and462_y0);
  and_gate and_gate_h_s_cla16_and463_y0(h_s_cla16_and462_y0, h_s_cla16_and461_y0, h_s_cla16_and463_y0);
  and_gate and_gate_h_s_cla16_and464_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and464_y0);
  and_gate and_gate_h_s_cla16_and465_y0(h_s_cla16_and464_y0, h_s_cla16_and463_y0, h_s_cla16_and465_y0);
  and_gate and_gate_h_s_cla16_and466_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and466_y0);
  and_gate and_gate_h_s_cla16_and467_y0(h_s_cla16_and466_y0, h_s_cla16_and465_y0, h_s_cla16_and467_y0);
  and_gate and_gate_h_s_cla16_and468_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and468_y0);
  and_gate and_gate_h_s_cla16_and469_y0(h_s_cla16_and468_y0, h_s_cla16_and467_y0, h_s_cla16_and469_y0);
  and_gate and_gate_h_s_cla16_and470_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and470_y0);
  and_gate and_gate_h_s_cla16_and471_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and471_y0);
  and_gate and_gate_h_s_cla16_and472_y0(h_s_cla16_and471_y0, h_s_cla16_and470_y0, h_s_cla16_and472_y0);
  and_gate and_gate_h_s_cla16_and473_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and473_y0);
  and_gate and_gate_h_s_cla16_and474_y0(h_s_cla16_and473_y0, h_s_cla16_and472_y0, h_s_cla16_and474_y0);
  and_gate and_gate_h_s_cla16_and475_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and475_y0);
  and_gate and_gate_h_s_cla16_and476_y0(h_s_cla16_and475_y0, h_s_cla16_and474_y0, h_s_cla16_and476_y0);
  and_gate and_gate_h_s_cla16_and477_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and477_y0);
  and_gate and_gate_h_s_cla16_and478_y0(h_s_cla16_and477_y0, h_s_cla16_and476_y0, h_s_cla16_and478_y0);
  and_gate and_gate_h_s_cla16_and479_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and479_y0);
  and_gate and_gate_h_s_cla16_and480_y0(h_s_cla16_and479_y0, h_s_cla16_and478_y0, h_s_cla16_and480_y0);
  and_gate and_gate_h_s_cla16_and481_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and481_y0);
  and_gate and_gate_h_s_cla16_and482_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and482_y0);
  and_gate and_gate_h_s_cla16_and483_y0(h_s_cla16_and482_y0, h_s_cla16_and481_y0, h_s_cla16_and483_y0);
  and_gate and_gate_h_s_cla16_and484_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and484_y0);
  and_gate and_gate_h_s_cla16_and485_y0(h_s_cla16_and484_y0, h_s_cla16_and483_y0, h_s_cla16_and485_y0);
  and_gate and_gate_h_s_cla16_and486_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and486_y0);
  and_gate and_gate_h_s_cla16_and487_y0(h_s_cla16_and486_y0, h_s_cla16_and485_y0, h_s_cla16_and487_y0);
  and_gate and_gate_h_s_cla16_and488_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and488_y0);
  and_gate and_gate_h_s_cla16_and489_y0(h_s_cla16_and488_y0, h_s_cla16_and487_y0, h_s_cla16_and489_y0);
  and_gate and_gate_h_s_cla16_and490_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and490_y0);
  and_gate and_gate_h_s_cla16_and491_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and491_y0);
  and_gate and_gate_h_s_cla16_and492_y0(h_s_cla16_and491_y0, h_s_cla16_and490_y0, h_s_cla16_and492_y0);
  and_gate and_gate_h_s_cla16_and493_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and493_y0);
  and_gate and_gate_h_s_cla16_and494_y0(h_s_cla16_and493_y0, h_s_cla16_and492_y0, h_s_cla16_and494_y0);
  and_gate and_gate_h_s_cla16_and495_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and495_y0);
  and_gate and_gate_h_s_cla16_and496_y0(h_s_cla16_and495_y0, h_s_cla16_and494_y0, h_s_cla16_and496_y0);
  and_gate and_gate_h_s_cla16_and497_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and497_y0);
  and_gate and_gate_h_s_cla16_and498_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and498_y0);
  and_gate and_gate_h_s_cla16_and499_y0(h_s_cla16_and498_y0, h_s_cla16_and497_y0, h_s_cla16_and499_y0);
  and_gate and_gate_h_s_cla16_and500_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and500_y0);
  and_gate and_gate_h_s_cla16_and501_y0(h_s_cla16_and500_y0, h_s_cla16_and499_y0, h_s_cla16_and501_y0);
  and_gate and_gate_h_s_cla16_and502_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and502_y0);
  and_gate and_gate_h_s_cla16_and503_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and503_y0);
  and_gate and_gate_h_s_cla16_and504_y0(h_s_cla16_and503_y0, h_s_cla16_and502_y0, h_s_cla16_and504_y0);
  and_gate and_gate_h_s_cla16_and505_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and505_y0);
  or_gate or_gate_h_s_cla16_or55_y0(h_s_cla16_and505_y0, h_s_cla16_and405_y0, h_s_cla16_or55_y0);
  or_gate or_gate_h_s_cla16_or56_y0(h_s_cla16_or55_y0, h_s_cla16_and424_y0, h_s_cla16_or56_y0);
  or_gate or_gate_h_s_cla16_or57_y0(h_s_cla16_or56_y0, h_s_cla16_and441_y0, h_s_cla16_or57_y0);
  or_gate or_gate_h_s_cla16_or58_y0(h_s_cla16_or57_y0, h_s_cla16_and456_y0, h_s_cla16_or58_y0);
  or_gate or_gate_h_s_cla16_or59_y0(h_s_cla16_or58_y0, h_s_cla16_and469_y0, h_s_cla16_or59_y0);
  or_gate or_gate_h_s_cla16_or60_y0(h_s_cla16_or59_y0, h_s_cla16_and480_y0, h_s_cla16_or60_y0);
  or_gate or_gate_h_s_cla16_or61_y0(h_s_cla16_or60_y0, h_s_cla16_and489_y0, h_s_cla16_or61_y0);
  or_gate or_gate_h_s_cla16_or62_y0(h_s_cla16_or61_y0, h_s_cla16_and496_y0, h_s_cla16_or62_y0);
  or_gate or_gate_h_s_cla16_or63_y0(h_s_cla16_or62_y0, h_s_cla16_and501_y0, h_s_cla16_or63_y0);
  or_gate or_gate_h_s_cla16_or64_y0(h_s_cla16_or63_y0, h_s_cla16_and504_y0, h_s_cla16_or64_y0);
  or_gate or_gate_h_s_cla16_or65_y0(h_s_cla16_pg_logic10_y1, h_s_cla16_or64_y0, h_s_cla16_or65_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic11_y0(a_11, b_11, h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_pg_logic11_y2);
  xor_gate xor_gate_h_s_cla16_xor11_y0(h_s_cla16_pg_logic11_y2, h_s_cla16_or65_y0, h_s_cla16_xor11_y0);
  and_gate and_gate_h_s_cla16_and506_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and506_y0);
  and_gate and_gate_h_s_cla16_and507_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and507_y0);
  and_gate and_gate_h_s_cla16_and508_y0(h_s_cla16_and507_y0, h_s_cla16_and506_y0, h_s_cla16_and508_y0);
  and_gate and_gate_h_s_cla16_and509_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and509_y0);
  and_gate and_gate_h_s_cla16_and510_y0(h_s_cla16_and509_y0, h_s_cla16_and508_y0, h_s_cla16_and510_y0);
  and_gate and_gate_h_s_cla16_and511_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and511_y0);
  and_gate and_gate_h_s_cla16_and512_y0(h_s_cla16_and511_y0, h_s_cla16_and510_y0, h_s_cla16_and512_y0);
  and_gate and_gate_h_s_cla16_and513_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and513_y0);
  and_gate and_gate_h_s_cla16_and514_y0(h_s_cla16_and513_y0, h_s_cla16_and512_y0, h_s_cla16_and514_y0);
  and_gate and_gate_h_s_cla16_and515_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and515_y0);
  and_gate and_gate_h_s_cla16_and516_y0(h_s_cla16_and515_y0, h_s_cla16_and514_y0, h_s_cla16_and516_y0);
  and_gate and_gate_h_s_cla16_and517_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and517_y0);
  and_gate and_gate_h_s_cla16_and518_y0(h_s_cla16_and517_y0, h_s_cla16_and516_y0, h_s_cla16_and518_y0);
  and_gate and_gate_h_s_cla16_and519_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and519_y0);
  and_gate and_gate_h_s_cla16_and520_y0(h_s_cla16_and519_y0, h_s_cla16_and518_y0, h_s_cla16_and520_y0);
  and_gate and_gate_h_s_cla16_and521_y0(h_s_cla16_pg_logic8_y0, constant_wire_0, h_s_cla16_and521_y0);
  and_gate and_gate_h_s_cla16_and522_y0(h_s_cla16_and521_y0, h_s_cla16_and520_y0, h_s_cla16_and522_y0);
  and_gate and_gate_h_s_cla16_and523_y0(h_s_cla16_pg_logic9_y0, constant_wire_0, h_s_cla16_and523_y0);
  and_gate and_gate_h_s_cla16_and524_y0(h_s_cla16_and523_y0, h_s_cla16_and522_y0, h_s_cla16_and524_y0);
  and_gate and_gate_h_s_cla16_and525_y0(h_s_cla16_pg_logic10_y0, constant_wire_0, h_s_cla16_and525_y0);
  and_gate and_gate_h_s_cla16_and526_y0(h_s_cla16_and525_y0, h_s_cla16_and524_y0, h_s_cla16_and526_y0);
  and_gate and_gate_h_s_cla16_and527_y0(h_s_cla16_pg_logic11_y0, constant_wire_0, h_s_cla16_and527_y0);
  and_gate and_gate_h_s_cla16_and528_y0(h_s_cla16_and527_y0, h_s_cla16_and526_y0, h_s_cla16_and528_y0);
  and_gate and_gate_h_s_cla16_and529_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and529_y0);
  and_gate and_gate_h_s_cla16_and530_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and530_y0);
  and_gate and_gate_h_s_cla16_and531_y0(h_s_cla16_and530_y0, h_s_cla16_and529_y0, h_s_cla16_and531_y0);
  and_gate and_gate_h_s_cla16_and532_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and532_y0);
  and_gate and_gate_h_s_cla16_and533_y0(h_s_cla16_and532_y0, h_s_cla16_and531_y0, h_s_cla16_and533_y0);
  and_gate and_gate_h_s_cla16_and534_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and534_y0);
  and_gate and_gate_h_s_cla16_and535_y0(h_s_cla16_and534_y0, h_s_cla16_and533_y0, h_s_cla16_and535_y0);
  and_gate and_gate_h_s_cla16_and536_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and536_y0);
  and_gate and_gate_h_s_cla16_and537_y0(h_s_cla16_and536_y0, h_s_cla16_and535_y0, h_s_cla16_and537_y0);
  and_gate and_gate_h_s_cla16_and538_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and538_y0);
  and_gate and_gate_h_s_cla16_and539_y0(h_s_cla16_and538_y0, h_s_cla16_and537_y0, h_s_cla16_and539_y0);
  and_gate and_gate_h_s_cla16_and540_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and540_y0);
  and_gate and_gate_h_s_cla16_and541_y0(h_s_cla16_and540_y0, h_s_cla16_and539_y0, h_s_cla16_and541_y0);
  and_gate and_gate_h_s_cla16_and542_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and542_y0);
  and_gate and_gate_h_s_cla16_and543_y0(h_s_cla16_and542_y0, h_s_cla16_and541_y0, h_s_cla16_and543_y0);
  and_gate and_gate_h_s_cla16_and544_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and544_y0);
  and_gate and_gate_h_s_cla16_and545_y0(h_s_cla16_and544_y0, h_s_cla16_and543_y0, h_s_cla16_and545_y0);
  and_gate and_gate_h_s_cla16_and546_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and546_y0);
  and_gate and_gate_h_s_cla16_and547_y0(h_s_cla16_and546_y0, h_s_cla16_and545_y0, h_s_cla16_and547_y0);
  and_gate and_gate_h_s_cla16_and548_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and548_y0);
  and_gate and_gate_h_s_cla16_and549_y0(h_s_cla16_and548_y0, h_s_cla16_and547_y0, h_s_cla16_and549_y0);
  and_gate and_gate_h_s_cla16_and550_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and550_y0);
  and_gate and_gate_h_s_cla16_and551_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and551_y0);
  and_gate and_gate_h_s_cla16_and552_y0(h_s_cla16_and551_y0, h_s_cla16_and550_y0, h_s_cla16_and552_y0);
  and_gate and_gate_h_s_cla16_and553_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and553_y0);
  and_gate and_gate_h_s_cla16_and554_y0(h_s_cla16_and553_y0, h_s_cla16_and552_y0, h_s_cla16_and554_y0);
  and_gate and_gate_h_s_cla16_and555_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and555_y0);
  and_gate and_gate_h_s_cla16_and556_y0(h_s_cla16_and555_y0, h_s_cla16_and554_y0, h_s_cla16_and556_y0);
  and_gate and_gate_h_s_cla16_and557_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and557_y0);
  and_gate and_gate_h_s_cla16_and558_y0(h_s_cla16_and557_y0, h_s_cla16_and556_y0, h_s_cla16_and558_y0);
  and_gate and_gate_h_s_cla16_and559_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and559_y0);
  and_gate and_gate_h_s_cla16_and560_y0(h_s_cla16_and559_y0, h_s_cla16_and558_y0, h_s_cla16_and560_y0);
  and_gate and_gate_h_s_cla16_and561_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and561_y0);
  and_gate and_gate_h_s_cla16_and562_y0(h_s_cla16_and561_y0, h_s_cla16_and560_y0, h_s_cla16_and562_y0);
  and_gate and_gate_h_s_cla16_and563_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and563_y0);
  and_gate and_gate_h_s_cla16_and564_y0(h_s_cla16_and563_y0, h_s_cla16_and562_y0, h_s_cla16_and564_y0);
  and_gate and_gate_h_s_cla16_and565_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and565_y0);
  and_gate and_gate_h_s_cla16_and566_y0(h_s_cla16_and565_y0, h_s_cla16_and564_y0, h_s_cla16_and566_y0);
  and_gate and_gate_h_s_cla16_and567_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and567_y0);
  and_gate and_gate_h_s_cla16_and568_y0(h_s_cla16_and567_y0, h_s_cla16_and566_y0, h_s_cla16_and568_y0);
  and_gate and_gate_h_s_cla16_and569_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and569_y0);
  and_gate and_gate_h_s_cla16_and570_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and570_y0);
  and_gate and_gate_h_s_cla16_and571_y0(h_s_cla16_and570_y0, h_s_cla16_and569_y0, h_s_cla16_and571_y0);
  and_gate and_gate_h_s_cla16_and572_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and572_y0);
  and_gate and_gate_h_s_cla16_and573_y0(h_s_cla16_and572_y0, h_s_cla16_and571_y0, h_s_cla16_and573_y0);
  and_gate and_gate_h_s_cla16_and574_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and574_y0);
  and_gate and_gate_h_s_cla16_and575_y0(h_s_cla16_and574_y0, h_s_cla16_and573_y0, h_s_cla16_and575_y0);
  and_gate and_gate_h_s_cla16_and576_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and576_y0);
  and_gate and_gate_h_s_cla16_and577_y0(h_s_cla16_and576_y0, h_s_cla16_and575_y0, h_s_cla16_and577_y0);
  and_gate and_gate_h_s_cla16_and578_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and578_y0);
  and_gate and_gate_h_s_cla16_and579_y0(h_s_cla16_and578_y0, h_s_cla16_and577_y0, h_s_cla16_and579_y0);
  and_gate and_gate_h_s_cla16_and580_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and580_y0);
  and_gate and_gate_h_s_cla16_and581_y0(h_s_cla16_and580_y0, h_s_cla16_and579_y0, h_s_cla16_and581_y0);
  and_gate and_gate_h_s_cla16_and582_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and582_y0);
  and_gate and_gate_h_s_cla16_and583_y0(h_s_cla16_and582_y0, h_s_cla16_and581_y0, h_s_cla16_and583_y0);
  and_gate and_gate_h_s_cla16_and584_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and584_y0);
  and_gate and_gate_h_s_cla16_and585_y0(h_s_cla16_and584_y0, h_s_cla16_and583_y0, h_s_cla16_and585_y0);
  and_gate and_gate_h_s_cla16_and586_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and586_y0);
  and_gate and_gate_h_s_cla16_and587_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and587_y0);
  and_gate and_gate_h_s_cla16_and588_y0(h_s_cla16_and587_y0, h_s_cla16_and586_y0, h_s_cla16_and588_y0);
  and_gate and_gate_h_s_cla16_and589_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and589_y0);
  and_gate and_gate_h_s_cla16_and590_y0(h_s_cla16_and589_y0, h_s_cla16_and588_y0, h_s_cla16_and590_y0);
  and_gate and_gate_h_s_cla16_and591_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and591_y0);
  and_gate and_gate_h_s_cla16_and592_y0(h_s_cla16_and591_y0, h_s_cla16_and590_y0, h_s_cla16_and592_y0);
  and_gate and_gate_h_s_cla16_and593_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and593_y0);
  and_gate and_gate_h_s_cla16_and594_y0(h_s_cla16_and593_y0, h_s_cla16_and592_y0, h_s_cla16_and594_y0);
  and_gate and_gate_h_s_cla16_and595_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and595_y0);
  and_gate and_gate_h_s_cla16_and596_y0(h_s_cla16_and595_y0, h_s_cla16_and594_y0, h_s_cla16_and596_y0);
  and_gate and_gate_h_s_cla16_and597_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and597_y0);
  and_gate and_gate_h_s_cla16_and598_y0(h_s_cla16_and597_y0, h_s_cla16_and596_y0, h_s_cla16_and598_y0);
  and_gate and_gate_h_s_cla16_and599_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and599_y0);
  and_gate and_gate_h_s_cla16_and600_y0(h_s_cla16_and599_y0, h_s_cla16_and598_y0, h_s_cla16_and600_y0);
  and_gate and_gate_h_s_cla16_and601_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and601_y0);
  and_gate and_gate_h_s_cla16_and602_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and602_y0);
  and_gate and_gate_h_s_cla16_and603_y0(h_s_cla16_and602_y0, h_s_cla16_and601_y0, h_s_cla16_and603_y0);
  and_gate and_gate_h_s_cla16_and604_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and604_y0);
  and_gate and_gate_h_s_cla16_and605_y0(h_s_cla16_and604_y0, h_s_cla16_and603_y0, h_s_cla16_and605_y0);
  and_gate and_gate_h_s_cla16_and606_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and606_y0);
  and_gate and_gate_h_s_cla16_and607_y0(h_s_cla16_and606_y0, h_s_cla16_and605_y0, h_s_cla16_and607_y0);
  and_gate and_gate_h_s_cla16_and608_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and608_y0);
  and_gate and_gate_h_s_cla16_and609_y0(h_s_cla16_and608_y0, h_s_cla16_and607_y0, h_s_cla16_and609_y0);
  and_gate and_gate_h_s_cla16_and610_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and610_y0);
  and_gate and_gate_h_s_cla16_and611_y0(h_s_cla16_and610_y0, h_s_cla16_and609_y0, h_s_cla16_and611_y0);
  and_gate and_gate_h_s_cla16_and612_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and612_y0);
  and_gate and_gate_h_s_cla16_and613_y0(h_s_cla16_and612_y0, h_s_cla16_and611_y0, h_s_cla16_and613_y0);
  and_gate and_gate_h_s_cla16_and614_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and614_y0);
  and_gate and_gate_h_s_cla16_and615_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and615_y0);
  and_gate and_gate_h_s_cla16_and616_y0(h_s_cla16_and615_y0, h_s_cla16_and614_y0, h_s_cla16_and616_y0);
  and_gate and_gate_h_s_cla16_and617_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and617_y0);
  and_gate and_gate_h_s_cla16_and618_y0(h_s_cla16_and617_y0, h_s_cla16_and616_y0, h_s_cla16_and618_y0);
  and_gate and_gate_h_s_cla16_and619_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and619_y0);
  and_gate and_gate_h_s_cla16_and620_y0(h_s_cla16_and619_y0, h_s_cla16_and618_y0, h_s_cla16_and620_y0);
  and_gate and_gate_h_s_cla16_and621_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and621_y0);
  and_gate and_gate_h_s_cla16_and622_y0(h_s_cla16_and621_y0, h_s_cla16_and620_y0, h_s_cla16_and622_y0);
  and_gate and_gate_h_s_cla16_and623_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and623_y0);
  and_gate and_gate_h_s_cla16_and624_y0(h_s_cla16_and623_y0, h_s_cla16_and622_y0, h_s_cla16_and624_y0);
  and_gate and_gate_h_s_cla16_and625_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and625_y0);
  and_gate and_gate_h_s_cla16_and626_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and626_y0);
  and_gate and_gate_h_s_cla16_and627_y0(h_s_cla16_and626_y0, h_s_cla16_and625_y0, h_s_cla16_and627_y0);
  and_gate and_gate_h_s_cla16_and628_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and628_y0);
  and_gate and_gate_h_s_cla16_and629_y0(h_s_cla16_and628_y0, h_s_cla16_and627_y0, h_s_cla16_and629_y0);
  and_gate and_gate_h_s_cla16_and630_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and630_y0);
  and_gate and_gate_h_s_cla16_and631_y0(h_s_cla16_and630_y0, h_s_cla16_and629_y0, h_s_cla16_and631_y0);
  and_gate and_gate_h_s_cla16_and632_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and632_y0);
  and_gate and_gate_h_s_cla16_and633_y0(h_s_cla16_and632_y0, h_s_cla16_and631_y0, h_s_cla16_and633_y0);
  and_gate and_gate_h_s_cla16_and634_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and634_y0);
  and_gate and_gate_h_s_cla16_and635_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and635_y0);
  and_gate and_gate_h_s_cla16_and636_y0(h_s_cla16_and635_y0, h_s_cla16_and634_y0, h_s_cla16_and636_y0);
  and_gate and_gate_h_s_cla16_and637_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and637_y0);
  and_gate and_gate_h_s_cla16_and638_y0(h_s_cla16_and637_y0, h_s_cla16_and636_y0, h_s_cla16_and638_y0);
  and_gate and_gate_h_s_cla16_and639_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and639_y0);
  and_gate and_gate_h_s_cla16_and640_y0(h_s_cla16_and639_y0, h_s_cla16_and638_y0, h_s_cla16_and640_y0);
  and_gate and_gate_h_s_cla16_and641_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and641_y0);
  and_gate and_gate_h_s_cla16_and642_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and642_y0);
  and_gate and_gate_h_s_cla16_and643_y0(h_s_cla16_and642_y0, h_s_cla16_and641_y0, h_s_cla16_and643_y0);
  and_gate and_gate_h_s_cla16_and644_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and644_y0);
  and_gate and_gate_h_s_cla16_and645_y0(h_s_cla16_and644_y0, h_s_cla16_and643_y0, h_s_cla16_and645_y0);
  and_gate and_gate_h_s_cla16_and646_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and646_y0);
  and_gate and_gate_h_s_cla16_and647_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and647_y0);
  and_gate and_gate_h_s_cla16_and648_y0(h_s_cla16_and647_y0, h_s_cla16_and646_y0, h_s_cla16_and648_y0);
  and_gate and_gate_h_s_cla16_and649_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and649_y0);
  or_gate or_gate_h_s_cla16_or66_y0(h_s_cla16_and649_y0, h_s_cla16_and528_y0, h_s_cla16_or66_y0);
  or_gate or_gate_h_s_cla16_or67_y0(h_s_cla16_or66_y0, h_s_cla16_and549_y0, h_s_cla16_or67_y0);
  or_gate or_gate_h_s_cla16_or68_y0(h_s_cla16_or67_y0, h_s_cla16_and568_y0, h_s_cla16_or68_y0);
  or_gate or_gate_h_s_cla16_or69_y0(h_s_cla16_or68_y0, h_s_cla16_and585_y0, h_s_cla16_or69_y0);
  or_gate or_gate_h_s_cla16_or70_y0(h_s_cla16_or69_y0, h_s_cla16_and600_y0, h_s_cla16_or70_y0);
  or_gate or_gate_h_s_cla16_or71_y0(h_s_cla16_or70_y0, h_s_cla16_and613_y0, h_s_cla16_or71_y0);
  or_gate or_gate_h_s_cla16_or72_y0(h_s_cla16_or71_y0, h_s_cla16_and624_y0, h_s_cla16_or72_y0);
  or_gate or_gate_h_s_cla16_or73_y0(h_s_cla16_or72_y0, h_s_cla16_and633_y0, h_s_cla16_or73_y0);
  or_gate or_gate_h_s_cla16_or74_y0(h_s_cla16_or73_y0, h_s_cla16_and640_y0, h_s_cla16_or74_y0);
  or_gate or_gate_h_s_cla16_or75_y0(h_s_cla16_or74_y0, h_s_cla16_and645_y0, h_s_cla16_or75_y0);
  or_gate or_gate_h_s_cla16_or76_y0(h_s_cla16_or75_y0, h_s_cla16_and648_y0, h_s_cla16_or76_y0);
  or_gate or_gate_h_s_cla16_or77_y0(h_s_cla16_pg_logic11_y1, h_s_cla16_or76_y0, h_s_cla16_or77_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic12_y0(a_12, b_12, h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic12_y1, h_s_cla16_pg_logic12_y2);
  xor_gate xor_gate_h_s_cla16_xor12_y0(h_s_cla16_pg_logic12_y2, h_s_cla16_or77_y0, h_s_cla16_xor12_y0);
  and_gate and_gate_h_s_cla16_and650_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and650_y0);
  and_gate and_gate_h_s_cla16_and651_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and651_y0);
  and_gate and_gate_h_s_cla16_and652_y0(h_s_cla16_and651_y0, h_s_cla16_and650_y0, h_s_cla16_and652_y0);
  and_gate and_gate_h_s_cla16_and653_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and653_y0);
  and_gate and_gate_h_s_cla16_and654_y0(h_s_cla16_and653_y0, h_s_cla16_and652_y0, h_s_cla16_and654_y0);
  and_gate and_gate_h_s_cla16_and655_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and655_y0);
  and_gate and_gate_h_s_cla16_and656_y0(h_s_cla16_and655_y0, h_s_cla16_and654_y0, h_s_cla16_and656_y0);
  and_gate and_gate_h_s_cla16_and657_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and657_y0);
  and_gate and_gate_h_s_cla16_and658_y0(h_s_cla16_and657_y0, h_s_cla16_and656_y0, h_s_cla16_and658_y0);
  and_gate and_gate_h_s_cla16_and659_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and659_y0);
  and_gate and_gate_h_s_cla16_and660_y0(h_s_cla16_and659_y0, h_s_cla16_and658_y0, h_s_cla16_and660_y0);
  and_gate and_gate_h_s_cla16_and661_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and661_y0);
  and_gate and_gate_h_s_cla16_and662_y0(h_s_cla16_and661_y0, h_s_cla16_and660_y0, h_s_cla16_and662_y0);
  and_gate and_gate_h_s_cla16_and663_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and663_y0);
  and_gate and_gate_h_s_cla16_and664_y0(h_s_cla16_and663_y0, h_s_cla16_and662_y0, h_s_cla16_and664_y0);
  and_gate and_gate_h_s_cla16_and665_y0(h_s_cla16_pg_logic8_y0, constant_wire_0, h_s_cla16_and665_y0);
  and_gate and_gate_h_s_cla16_and666_y0(h_s_cla16_and665_y0, h_s_cla16_and664_y0, h_s_cla16_and666_y0);
  and_gate and_gate_h_s_cla16_and667_y0(h_s_cla16_pg_logic9_y0, constant_wire_0, h_s_cla16_and667_y0);
  and_gate and_gate_h_s_cla16_and668_y0(h_s_cla16_and667_y0, h_s_cla16_and666_y0, h_s_cla16_and668_y0);
  and_gate and_gate_h_s_cla16_and669_y0(h_s_cla16_pg_logic10_y0, constant_wire_0, h_s_cla16_and669_y0);
  and_gate and_gate_h_s_cla16_and670_y0(h_s_cla16_and669_y0, h_s_cla16_and668_y0, h_s_cla16_and670_y0);
  and_gate and_gate_h_s_cla16_and671_y0(h_s_cla16_pg_logic11_y0, constant_wire_0, h_s_cla16_and671_y0);
  and_gate and_gate_h_s_cla16_and672_y0(h_s_cla16_and671_y0, h_s_cla16_and670_y0, h_s_cla16_and672_y0);
  and_gate and_gate_h_s_cla16_and673_y0(h_s_cla16_pg_logic12_y0, constant_wire_0, h_s_cla16_and673_y0);
  and_gate and_gate_h_s_cla16_and674_y0(h_s_cla16_and673_y0, h_s_cla16_and672_y0, h_s_cla16_and674_y0);
  and_gate and_gate_h_s_cla16_and675_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and675_y0);
  and_gate and_gate_h_s_cla16_and676_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and676_y0);
  and_gate and_gate_h_s_cla16_and677_y0(h_s_cla16_and676_y0, h_s_cla16_and675_y0, h_s_cla16_and677_y0);
  and_gate and_gate_h_s_cla16_and678_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and678_y0);
  and_gate and_gate_h_s_cla16_and679_y0(h_s_cla16_and678_y0, h_s_cla16_and677_y0, h_s_cla16_and679_y0);
  and_gate and_gate_h_s_cla16_and680_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and680_y0);
  and_gate and_gate_h_s_cla16_and681_y0(h_s_cla16_and680_y0, h_s_cla16_and679_y0, h_s_cla16_and681_y0);
  and_gate and_gate_h_s_cla16_and682_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and682_y0);
  and_gate and_gate_h_s_cla16_and683_y0(h_s_cla16_and682_y0, h_s_cla16_and681_y0, h_s_cla16_and683_y0);
  and_gate and_gate_h_s_cla16_and684_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and684_y0);
  and_gate and_gate_h_s_cla16_and685_y0(h_s_cla16_and684_y0, h_s_cla16_and683_y0, h_s_cla16_and685_y0);
  and_gate and_gate_h_s_cla16_and686_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and686_y0);
  and_gate and_gate_h_s_cla16_and687_y0(h_s_cla16_and686_y0, h_s_cla16_and685_y0, h_s_cla16_and687_y0);
  and_gate and_gate_h_s_cla16_and688_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and688_y0);
  and_gate and_gate_h_s_cla16_and689_y0(h_s_cla16_and688_y0, h_s_cla16_and687_y0, h_s_cla16_and689_y0);
  and_gate and_gate_h_s_cla16_and690_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and690_y0);
  and_gate and_gate_h_s_cla16_and691_y0(h_s_cla16_and690_y0, h_s_cla16_and689_y0, h_s_cla16_and691_y0);
  and_gate and_gate_h_s_cla16_and692_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and692_y0);
  and_gate and_gate_h_s_cla16_and693_y0(h_s_cla16_and692_y0, h_s_cla16_and691_y0, h_s_cla16_and693_y0);
  and_gate and_gate_h_s_cla16_and694_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and694_y0);
  and_gate and_gate_h_s_cla16_and695_y0(h_s_cla16_and694_y0, h_s_cla16_and693_y0, h_s_cla16_and695_y0);
  and_gate and_gate_h_s_cla16_and696_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and696_y0);
  and_gate and_gate_h_s_cla16_and697_y0(h_s_cla16_and696_y0, h_s_cla16_and695_y0, h_s_cla16_and697_y0);
  and_gate and_gate_h_s_cla16_and698_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and698_y0);
  and_gate and_gate_h_s_cla16_and699_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and699_y0);
  and_gate and_gate_h_s_cla16_and700_y0(h_s_cla16_and699_y0, h_s_cla16_and698_y0, h_s_cla16_and700_y0);
  and_gate and_gate_h_s_cla16_and701_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and701_y0);
  and_gate and_gate_h_s_cla16_and702_y0(h_s_cla16_and701_y0, h_s_cla16_and700_y0, h_s_cla16_and702_y0);
  and_gate and_gate_h_s_cla16_and703_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and703_y0);
  and_gate and_gate_h_s_cla16_and704_y0(h_s_cla16_and703_y0, h_s_cla16_and702_y0, h_s_cla16_and704_y0);
  and_gate and_gate_h_s_cla16_and705_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and705_y0);
  and_gate and_gate_h_s_cla16_and706_y0(h_s_cla16_and705_y0, h_s_cla16_and704_y0, h_s_cla16_and706_y0);
  and_gate and_gate_h_s_cla16_and707_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and707_y0);
  and_gate and_gate_h_s_cla16_and708_y0(h_s_cla16_and707_y0, h_s_cla16_and706_y0, h_s_cla16_and708_y0);
  and_gate and_gate_h_s_cla16_and709_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and709_y0);
  and_gate and_gate_h_s_cla16_and710_y0(h_s_cla16_and709_y0, h_s_cla16_and708_y0, h_s_cla16_and710_y0);
  and_gate and_gate_h_s_cla16_and711_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and711_y0);
  and_gate and_gate_h_s_cla16_and712_y0(h_s_cla16_and711_y0, h_s_cla16_and710_y0, h_s_cla16_and712_y0);
  and_gate and_gate_h_s_cla16_and713_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and713_y0);
  and_gate and_gate_h_s_cla16_and714_y0(h_s_cla16_and713_y0, h_s_cla16_and712_y0, h_s_cla16_and714_y0);
  and_gate and_gate_h_s_cla16_and715_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and715_y0);
  and_gate and_gate_h_s_cla16_and716_y0(h_s_cla16_and715_y0, h_s_cla16_and714_y0, h_s_cla16_and716_y0);
  and_gate and_gate_h_s_cla16_and717_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and717_y0);
  and_gate and_gate_h_s_cla16_and718_y0(h_s_cla16_and717_y0, h_s_cla16_and716_y0, h_s_cla16_and718_y0);
  and_gate and_gate_h_s_cla16_and719_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and719_y0);
  and_gate and_gate_h_s_cla16_and720_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and720_y0);
  and_gate and_gate_h_s_cla16_and721_y0(h_s_cla16_and720_y0, h_s_cla16_and719_y0, h_s_cla16_and721_y0);
  and_gate and_gate_h_s_cla16_and722_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and722_y0);
  and_gate and_gate_h_s_cla16_and723_y0(h_s_cla16_and722_y0, h_s_cla16_and721_y0, h_s_cla16_and723_y0);
  and_gate and_gate_h_s_cla16_and724_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and724_y0);
  and_gate and_gate_h_s_cla16_and725_y0(h_s_cla16_and724_y0, h_s_cla16_and723_y0, h_s_cla16_and725_y0);
  and_gate and_gate_h_s_cla16_and726_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and726_y0);
  and_gate and_gate_h_s_cla16_and727_y0(h_s_cla16_and726_y0, h_s_cla16_and725_y0, h_s_cla16_and727_y0);
  and_gate and_gate_h_s_cla16_and728_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and728_y0);
  and_gate and_gate_h_s_cla16_and729_y0(h_s_cla16_and728_y0, h_s_cla16_and727_y0, h_s_cla16_and729_y0);
  and_gate and_gate_h_s_cla16_and730_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and730_y0);
  and_gate and_gate_h_s_cla16_and731_y0(h_s_cla16_and730_y0, h_s_cla16_and729_y0, h_s_cla16_and731_y0);
  and_gate and_gate_h_s_cla16_and732_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and732_y0);
  and_gate and_gate_h_s_cla16_and733_y0(h_s_cla16_and732_y0, h_s_cla16_and731_y0, h_s_cla16_and733_y0);
  and_gate and_gate_h_s_cla16_and734_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and734_y0);
  and_gate and_gate_h_s_cla16_and735_y0(h_s_cla16_and734_y0, h_s_cla16_and733_y0, h_s_cla16_and735_y0);
  and_gate and_gate_h_s_cla16_and736_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and736_y0);
  and_gate and_gate_h_s_cla16_and737_y0(h_s_cla16_and736_y0, h_s_cla16_and735_y0, h_s_cla16_and737_y0);
  and_gate and_gate_h_s_cla16_and738_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and738_y0);
  and_gate and_gate_h_s_cla16_and739_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and739_y0);
  and_gate and_gate_h_s_cla16_and740_y0(h_s_cla16_and739_y0, h_s_cla16_and738_y0, h_s_cla16_and740_y0);
  and_gate and_gate_h_s_cla16_and741_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and741_y0);
  and_gate and_gate_h_s_cla16_and742_y0(h_s_cla16_and741_y0, h_s_cla16_and740_y0, h_s_cla16_and742_y0);
  and_gate and_gate_h_s_cla16_and743_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and743_y0);
  and_gate and_gate_h_s_cla16_and744_y0(h_s_cla16_and743_y0, h_s_cla16_and742_y0, h_s_cla16_and744_y0);
  and_gate and_gate_h_s_cla16_and745_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and745_y0);
  and_gate and_gate_h_s_cla16_and746_y0(h_s_cla16_and745_y0, h_s_cla16_and744_y0, h_s_cla16_and746_y0);
  and_gate and_gate_h_s_cla16_and747_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and747_y0);
  and_gate and_gate_h_s_cla16_and748_y0(h_s_cla16_and747_y0, h_s_cla16_and746_y0, h_s_cla16_and748_y0);
  and_gate and_gate_h_s_cla16_and749_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and749_y0);
  and_gate and_gate_h_s_cla16_and750_y0(h_s_cla16_and749_y0, h_s_cla16_and748_y0, h_s_cla16_and750_y0);
  and_gate and_gate_h_s_cla16_and751_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and751_y0);
  and_gate and_gate_h_s_cla16_and752_y0(h_s_cla16_and751_y0, h_s_cla16_and750_y0, h_s_cla16_and752_y0);
  and_gate and_gate_h_s_cla16_and753_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and753_y0);
  and_gate and_gate_h_s_cla16_and754_y0(h_s_cla16_and753_y0, h_s_cla16_and752_y0, h_s_cla16_and754_y0);
  and_gate and_gate_h_s_cla16_and755_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and755_y0);
  and_gate and_gate_h_s_cla16_and756_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and756_y0);
  and_gate and_gate_h_s_cla16_and757_y0(h_s_cla16_and756_y0, h_s_cla16_and755_y0, h_s_cla16_and757_y0);
  and_gate and_gate_h_s_cla16_and758_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and758_y0);
  and_gate and_gate_h_s_cla16_and759_y0(h_s_cla16_and758_y0, h_s_cla16_and757_y0, h_s_cla16_and759_y0);
  and_gate and_gate_h_s_cla16_and760_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and760_y0);
  and_gate and_gate_h_s_cla16_and761_y0(h_s_cla16_and760_y0, h_s_cla16_and759_y0, h_s_cla16_and761_y0);
  and_gate and_gate_h_s_cla16_and762_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and762_y0);
  and_gate and_gate_h_s_cla16_and763_y0(h_s_cla16_and762_y0, h_s_cla16_and761_y0, h_s_cla16_and763_y0);
  and_gate and_gate_h_s_cla16_and764_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and764_y0);
  and_gate and_gate_h_s_cla16_and765_y0(h_s_cla16_and764_y0, h_s_cla16_and763_y0, h_s_cla16_and765_y0);
  and_gate and_gate_h_s_cla16_and766_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and766_y0);
  and_gate and_gate_h_s_cla16_and767_y0(h_s_cla16_and766_y0, h_s_cla16_and765_y0, h_s_cla16_and767_y0);
  and_gate and_gate_h_s_cla16_and768_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and768_y0);
  and_gate and_gate_h_s_cla16_and769_y0(h_s_cla16_and768_y0, h_s_cla16_and767_y0, h_s_cla16_and769_y0);
  and_gate and_gate_h_s_cla16_and770_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and770_y0);
  and_gate and_gate_h_s_cla16_and771_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and771_y0);
  and_gate and_gate_h_s_cla16_and772_y0(h_s_cla16_and771_y0, h_s_cla16_and770_y0, h_s_cla16_and772_y0);
  and_gate and_gate_h_s_cla16_and773_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and773_y0);
  and_gate and_gate_h_s_cla16_and774_y0(h_s_cla16_and773_y0, h_s_cla16_and772_y0, h_s_cla16_and774_y0);
  and_gate and_gate_h_s_cla16_and775_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and775_y0);
  and_gate and_gate_h_s_cla16_and776_y0(h_s_cla16_and775_y0, h_s_cla16_and774_y0, h_s_cla16_and776_y0);
  and_gate and_gate_h_s_cla16_and777_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and777_y0);
  and_gate and_gate_h_s_cla16_and778_y0(h_s_cla16_and777_y0, h_s_cla16_and776_y0, h_s_cla16_and778_y0);
  and_gate and_gate_h_s_cla16_and779_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and779_y0);
  and_gate and_gate_h_s_cla16_and780_y0(h_s_cla16_and779_y0, h_s_cla16_and778_y0, h_s_cla16_and780_y0);
  and_gate and_gate_h_s_cla16_and781_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and781_y0);
  and_gate and_gate_h_s_cla16_and782_y0(h_s_cla16_and781_y0, h_s_cla16_and780_y0, h_s_cla16_and782_y0);
  and_gate and_gate_h_s_cla16_and783_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and783_y0);
  and_gate and_gate_h_s_cla16_and784_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and784_y0);
  and_gate and_gate_h_s_cla16_and785_y0(h_s_cla16_and784_y0, h_s_cla16_and783_y0, h_s_cla16_and785_y0);
  and_gate and_gate_h_s_cla16_and786_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and786_y0);
  and_gate and_gate_h_s_cla16_and787_y0(h_s_cla16_and786_y0, h_s_cla16_and785_y0, h_s_cla16_and787_y0);
  and_gate and_gate_h_s_cla16_and788_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and788_y0);
  and_gate and_gate_h_s_cla16_and789_y0(h_s_cla16_and788_y0, h_s_cla16_and787_y0, h_s_cla16_and789_y0);
  and_gate and_gate_h_s_cla16_and790_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and790_y0);
  and_gate and_gate_h_s_cla16_and791_y0(h_s_cla16_and790_y0, h_s_cla16_and789_y0, h_s_cla16_and791_y0);
  and_gate and_gate_h_s_cla16_and792_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and792_y0);
  and_gate and_gate_h_s_cla16_and793_y0(h_s_cla16_and792_y0, h_s_cla16_and791_y0, h_s_cla16_and793_y0);
  and_gate and_gate_h_s_cla16_and794_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and794_y0);
  and_gate and_gate_h_s_cla16_and795_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and795_y0);
  and_gate and_gate_h_s_cla16_and796_y0(h_s_cla16_and795_y0, h_s_cla16_and794_y0, h_s_cla16_and796_y0);
  and_gate and_gate_h_s_cla16_and797_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and797_y0);
  and_gate and_gate_h_s_cla16_and798_y0(h_s_cla16_and797_y0, h_s_cla16_and796_y0, h_s_cla16_and798_y0);
  and_gate and_gate_h_s_cla16_and799_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and799_y0);
  and_gate and_gate_h_s_cla16_and800_y0(h_s_cla16_and799_y0, h_s_cla16_and798_y0, h_s_cla16_and800_y0);
  and_gate and_gate_h_s_cla16_and801_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and801_y0);
  and_gate and_gate_h_s_cla16_and802_y0(h_s_cla16_and801_y0, h_s_cla16_and800_y0, h_s_cla16_and802_y0);
  and_gate and_gate_h_s_cla16_and803_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and803_y0);
  and_gate and_gate_h_s_cla16_and804_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and804_y0);
  and_gate and_gate_h_s_cla16_and805_y0(h_s_cla16_and804_y0, h_s_cla16_and803_y0, h_s_cla16_and805_y0);
  and_gate and_gate_h_s_cla16_and806_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and806_y0);
  and_gate and_gate_h_s_cla16_and807_y0(h_s_cla16_and806_y0, h_s_cla16_and805_y0, h_s_cla16_and807_y0);
  and_gate and_gate_h_s_cla16_and808_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and808_y0);
  and_gate and_gate_h_s_cla16_and809_y0(h_s_cla16_and808_y0, h_s_cla16_and807_y0, h_s_cla16_and809_y0);
  and_gate and_gate_h_s_cla16_and810_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and810_y0);
  and_gate and_gate_h_s_cla16_and811_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and811_y0);
  and_gate and_gate_h_s_cla16_and812_y0(h_s_cla16_and811_y0, h_s_cla16_and810_y0, h_s_cla16_and812_y0);
  and_gate and_gate_h_s_cla16_and813_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and813_y0);
  and_gate and_gate_h_s_cla16_and814_y0(h_s_cla16_and813_y0, h_s_cla16_and812_y0, h_s_cla16_and814_y0);
  and_gate and_gate_h_s_cla16_and815_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and815_y0);
  and_gate and_gate_h_s_cla16_and816_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and816_y0);
  and_gate and_gate_h_s_cla16_and817_y0(h_s_cla16_and816_y0, h_s_cla16_and815_y0, h_s_cla16_and817_y0);
  and_gate and_gate_h_s_cla16_and818_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and818_y0);
  or_gate or_gate_h_s_cla16_or78_y0(h_s_cla16_and818_y0, h_s_cla16_and674_y0, h_s_cla16_or78_y0);
  or_gate or_gate_h_s_cla16_or79_y0(h_s_cla16_or78_y0, h_s_cla16_and697_y0, h_s_cla16_or79_y0);
  or_gate or_gate_h_s_cla16_or80_y0(h_s_cla16_or79_y0, h_s_cla16_and718_y0, h_s_cla16_or80_y0);
  or_gate or_gate_h_s_cla16_or81_y0(h_s_cla16_or80_y0, h_s_cla16_and737_y0, h_s_cla16_or81_y0);
  or_gate or_gate_h_s_cla16_or82_y0(h_s_cla16_or81_y0, h_s_cla16_and754_y0, h_s_cla16_or82_y0);
  or_gate or_gate_h_s_cla16_or83_y0(h_s_cla16_or82_y0, h_s_cla16_and769_y0, h_s_cla16_or83_y0);
  or_gate or_gate_h_s_cla16_or84_y0(h_s_cla16_or83_y0, h_s_cla16_and782_y0, h_s_cla16_or84_y0);
  or_gate or_gate_h_s_cla16_or85_y0(h_s_cla16_or84_y0, h_s_cla16_and793_y0, h_s_cla16_or85_y0);
  or_gate or_gate_h_s_cla16_or86_y0(h_s_cla16_or85_y0, h_s_cla16_and802_y0, h_s_cla16_or86_y0);
  or_gate or_gate_h_s_cla16_or87_y0(h_s_cla16_or86_y0, h_s_cla16_and809_y0, h_s_cla16_or87_y0);
  or_gate or_gate_h_s_cla16_or88_y0(h_s_cla16_or87_y0, h_s_cla16_and814_y0, h_s_cla16_or88_y0);
  or_gate or_gate_h_s_cla16_or89_y0(h_s_cla16_or88_y0, h_s_cla16_and817_y0, h_s_cla16_or89_y0);
  or_gate or_gate_h_s_cla16_or90_y0(h_s_cla16_pg_logic12_y1, h_s_cla16_or89_y0, h_s_cla16_or90_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic13_y0(a_13, b_13, h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic13_y1, h_s_cla16_pg_logic13_y2);
  xor_gate xor_gate_h_s_cla16_xor13_y0(h_s_cla16_pg_logic13_y2, h_s_cla16_or90_y0, h_s_cla16_xor13_y0);
  and_gate and_gate_h_s_cla16_and819_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and819_y0);
  and_gate and_gate_h_s_cla16_and820_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and820_y0);
  and_gate and_gate_h_s_cla16_and821_y0(h_s_cla16_and820_y0, h_s_cla16_and819_y0, h_s_cla16_and821_y0);
  and_gate and_gate_h_s_cla16_and822_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and822_y0);
  and_gate and_gate_h_s_cla16_and823_y0(h_s_cla16_and822_y0, h_s_cla16_and821_y0, h_s_cla16_and823_y0);
  and_gate and_gate_h_s_cla16_and824_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and824_y0);
  and_gate and_gate_h_s_cla16_and825_y0(h_s_cla16_and824_y0, h_s_cla16_and823_y0, h_s_cla16_and825_y0);
  and_gate and_gate_h_s_cla16_and826_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and826_y0);
  and_gate and_gate_h_s_cla16_and827_y0(h_s_cla16_and826_y0, h_s_cla16_and825_y0, h_s_cla16_and827_y0);
  and_gate and_gate_h_s_cla16_and828_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and828_y0);
  and_gate and_gate_h_s_cla16_and829_y0(h_s_cla16_and828_y0, h_s_cla16_and827_y0, h_s_cla16_and829_y0);
  and_gate and_gate_h_s_cla16_and830_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and830_y0);
  and_gate and_gate_h_s_cla16_and831_y0(h_s_cla16_and830_y0, h_s_cla16_and829_y0, h_s_cla16_and831_y0);
  and_gate and_gate_h_s_cla16_and832_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and832_y0);
  and_gate and_gate_h_s_cla16_and833_y0(h_s_cla16_and832_y0, h_s_cla16_and831_y0, h_s_cla16_and833_y0);
  and_gate and_gate_h_s_cla16_and834_y0(h_s_cla16_pg_logic8_y0, constant_wire_0, h_s_cla16_and834_y0);
  and_gate and_gate_h_s_cla16_and835_y0(h_s_cla16_and834_y0, h_s_cla16_and833_y0, h_s_cla16_and835_y0);
  and_gate and_gate_h_s_cla16_and836_y0(h_s_cla16_pg_logic9_y0, constant_wire_0, h_s_cla16_and836_y0);
  and_gate and_gate_h_s_cla16_and837_y0(h_s_cla16_and836_y0, h_s_cla16_and835_y0, h_s_cla16_and837_y0);
  and_gate and_gate_h_s_cla16_and838_y0(h_s_cla16_pg_logic10_y0, constant_wire_0, h_s_cla16_and838_y0);
  and_gate and_gate_h_s_cla16_and839_y0(h_s_cla16_and838_y0, h_s_cla16_and837_y0, h_s_cla16_and839_y0);
  and_gate and_gate_h_s_cla16_and840_y0(h_s_cla16_pg_logic11_y0, constant_wire_0, h_s_cla16_and840_y0);
  and_gate and_gate_h_s_cla16_and841_y0(h_s_cla16_and840_y0, h_s_cla16_and839_y0, h_s_cla16_and841_y0);
  and_gate and_gate_h_s_cla16_and842_y0(h_s_cla16_pg_logic12_y0, constant_wire_0, h_s_cla16_and842_y0);
  and_gate and_gate_h_s_cla16_and843_y0(h_s_cla16_and842_y0, h_s_cla16_and841_y0, h_s_cla16_and843_y0);
  and_gate and_gate_h_s_cla16_and844_y0(h_s_cla16_pg_logic13_y0, constant_wire_0, h_s_cla16_and844_y0);
  and_gate and_gate_h_s_cla16_and845_y0(h_s_cla16_and844_y0, h_s_cla16_and843_y0, h_s_cla16_and845_y0);
  and_gate and_gate_h_s_cla16_and846_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and846_y0);
  and_gate and_gate_h_s_cla16_and847_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and847_y0);
  and_gate and_gate_h_s_cla16_and848_y0(h_s_cla16_and847_y0, h_s_cla16_and846_y0, h_s_cla16_and848_y0);
  and_gate and_gate_h_s_cla16_and849_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and849_y0);
  and_gate and_gate_h_s_cla16_and850_y0(h_s_cla16_and849_y0, h_s_cla16_and848_y0, h_s_cla16_and850_y0);
  and_gate and_gate_h_s_cla16_and851_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and851_y0);
  and_gate and_gate_h_s_cla16_and852_y0(h_s_cla16_and851_y0, h_s_cla16_and850_y0, h_s_cla16_and852_y0);
  and_gate and_gate_h_s_cla16_and853_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and853_y0);
  and_gate and_gate_h_s_cla16_and854_y0(h_s_cla16_and853_y0, h_s_cla16_and852_y0, h_s_cla16_and854_y0);
  and_gate and_gate_h_s_cla16_and855_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and855_y0);
  and_gate and_gate_h_s_cla16_and856_y0(h_s_cla16_and855_y0, h_s_cla16_and854_y0, h_s_cla16_and856_y0);
  and_gate and_gate_h_s_cla16_and857_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and857_y0);
  and_gate and_gate_h_s_cla16_and858_y0(h_s_cla16_and857_y0, h_s_cla16_and856_y0, h_s_cla16_and858_y0);
  and_gate and_gate_h_s_cla16_and859_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and859_y0);
  and_gate and_gate_h_s_cla16_and860_y0(h_s_cla16_and859_y0, h_s_cla16_and858_y0, h_s_cla16_and860_y0);
  and_gate and_gate_h_s_cla16_and861_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and861_y0);
  and_gate and_gate_h_s_cla16_and862_y0(h_s_cla16_and861_y0, h_s_cla16_and860_y0, h_s_cla16_and862_y0);
  and_gate and_gate_h_s_cla16_and863_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and863_y0);
  and_gate and_gate_h_s_cla16_and864_y0(h_s_cla16_and863_y0, h_s_cla16_and862_y0, h_s_cla16_and864_y0);
  and_gate and_gate_h_s_cla16_and865_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and865_y0);
  and_gate and_gate_h_s_cla16_and866_y0(h_s_cla16_and865_y0, h_s_cla16_and864_y0, h_s_cla16_and866_y0);
  and_gate and_gate_h_s_cla16_and867_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and867_y0);
  and_gate and_gate_h_s_cla16_and868_y0(h_s_cla16_and867_y0, h_s_cla16_and866_y0, h_s_cla16_and868_y0);
  and_gate and_gate_h_s_cla16_and869_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and869_y0);
  and_gate and_gate_h_s_cla16_and870_y0(h_s_cla16_and869_y0, h_s_cla16_and868_y0, h_s_cla16_and870_y0);
  and_gate and_gate_h_s_cla16_and871_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and871_y0);
  and_gate and_gate_h_s_cla16_and872_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and872_y0);
  and_gate and_gate_h_s_cla16_and873_y0(h_s_cla16_and872_y0, h_s_cla16_and871_y0, h_s_cla16_and873_y0);
  and_gate and_gate_h_s_cla16_and874_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and874_y0);
  and_gate and_gate_h_s_cla16_and875_y0(h_s_cla16_and874_y0, h_s_cla16_and873_y0, h_s_cla16_and875_y0);
  and_gate and_gate_h_s_cla16_and876_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and876_y0);
  and_gate and_gate_h_s_cla16_and877_y0(h_s_cla16_and876_y0, h_s_cla16_and875_y0, h_s_cla16_and877_y0);
  and_gate and_gate_h_s_cla16_and878_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and878_y0);
  and_gate and_gate_h_s_cla16_and879_y0(h_s_cla16_and878_y0, h_s_cla16_and877_y0, h_s_cla16_and879_y0);
  and_gate and_gate_h_s_cla16_and880_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and880_y0);
  and_gate and_gate_h_s_cla16_and881_y0(h_s_cla16_and880_y0, h_s_cla16_and879_y0, h_s_cla16_and881_y0);
  and_gate and_gate_h_s_cla16_and882_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and882_y0);
  and_gate and_gate_h_s_cla16_and883_y0(h_s_cla16_and882_y0, h_s_cla16_and881_y0, h_s_cla16_and883_y0);
  and_gate and_gate_h_s_cla16_and884_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and884_y0);
  and_gate and_gate_h_s_cla16_and885_y0(h_s_cla16_and884_y0, h_s_cla16_and883_y0, h_s_cla16_and885_y0);
  and_gate and_gate_h_s_cla16_and886_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and886_y0);
  and_gate and_gate_h_s_cla16_and887_y0(h_s_cla16_and886_y0, h_s_cla16_and885_y0, h_s_cla16_and887_y0);
  and_gate and_gate_h_s_cla16_and888_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and888_y0);
  and_gate and_gate_h_s_cla16_and889_y0(h_s_cla16_and888_y0, h_s_cla16_and887_y0, h_s_cla16_and889_y0);
  and_gate and_gate_h_s_cla16_and890_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and890_y0);
  and_gate and_gate_h_s_cla16_and891_y0(h_s_cla16_and890_y0, h_s_cla16_and889_y0, h_s_cla16_and891_y0);
  and_gate and_gate_h_s_cla16_and892_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and892_y0);
  and_gate and_gate_h_s_cla16_and893_y0(h_s_cla16_and892_y0, h_s_cla16_and891_y0, h_s_cla16_and893_y0);
  and_gate and_gate_h_s_cla16_and894_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and894_y0);
  and_gate and_gate_h_s_cla16_and895_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and895_y0);
  and_gate and_gate_h_s_cla16_and896_y0(h_s_cla16_and895_y0, h_s_cla16_and894_y0, h_s_cla16_and896_y0);
  and_gate and_gate_h_s_cla16_and897_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and897_y0);
  and_gate and_gate_h_s_cla16_and898_y0(h_s_cla16_and897_y0, h_s_cla16_and896_y0, h_s_cla16_and898_y0);
  and_gate and_gate_h_s_cla16_and899_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and899_y0);
  and_gate and_gate_h_s_cla16_and900_y0(h_s_cla16_and899_y0, h_s_cla16_and898_y0, h_s_cla16_and900_y0);
  and_gate and_gate_h_s_cla16_and901_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and901_y0);
  and_gate and_gate_h_s_cla16_and902_y0(h_s_cla16_and901_y0, h_s_cla16_and900_y0, h_s_cla16_and902_y0);
  and_gate and_gate_h_s_cla16_and903_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and903_y0);
  and_gate and_gate_h_s_cla16_and904_y0(h_s_cla16_and903_y0, h_s_cla16_and902_y0, h_s_cla16_and904_y0);
  and_gate and_gate_h_s_cla16_and905_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and905_y0);
  and_gate and_gate_h_s_cla16_and906_y0(h_s_cla16_and905_y0, h_s_cla16_and904_y0, h_s_cla16_and906_y0);
  and_gate and_gate_h_s_cla16_and907_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and907_y0);
  and_gate and_gate_h_s_cla16_and908_y0(h_s_cla16_and907_y0, h_s_cla16_and906_y0, h_s_cla16_and908_y0);
  and_gate and_gate_h_s_cla16_and909_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and909_y0);
  and_gate and_gate_h_s_cla16_and910_y0(h_s_cla16_and909_y0, h_s_cla16_and908_y0, h_s_cla16_and910_y0);
  and_gate and_gate_h_s_cla16_and911_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and911_y0);
  and_gate and_gate_h_s_cla16_and912_y0(h_s_cla16_and911_y0, h_s_cla16_and910_y0, h_s_cla16_and912_y0);
  and_gate and_gate_h_s_cla16_and913_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and913_y0);
  and_gate and_gate_h_s_cla16_and914_y0(h_s_cla16_and913_y0, h_s_cla16_and912_y0, h_s_cla16_and914_y0);
  and_gate and_gate_h_s_cla16_and915_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and915_y0);
  and_gate and_gate_h_s_cla16_and916_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and916_y0);
  and_gate and_gate_h_s_cla16_and917_y0(h_s_cla16_and916_y0, h_s_cla16_and915_y0, h_s_cla16_and917_y0);
  and_gate and_gate_h_s_cla16_and918_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and918_y0);
  and_gate and_gate_h_s_cla16_and919_y0(h_s_cla16_and918_y0, h_s_cla16_and917_y0, h_s_cla16_and919_y0);
  and_gate and_gate_h_s_cla16_and920_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and920_y0);
  and_gate and_gate_h_s_cla16_and921_y0(h_s_cla16_and920_y0, h_s_cla16_and919_y0, h_s_cla16_and921_y0);
  and_gate and_gate_h_s_cla16_and922_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and922_y0);
  and_gate and_gate_h_s_cla16_and923_y0(h_s_cla16_and922_y0, h_s_cla16_and921_y0, h_s_cla16_and923_y0);
  and_gate and_gate_h_s_cla16_and924_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and924_y0);
  and_gate and_gate_h_s_cla16_and925_y0(h_s_cla16_and924_y0, h_s_cla16_and923_y0, h_s_cla16_and925_y0);
  and_gate and_gate_h_s_cla16_and926_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and926_y0);
  and_gate and_gate_h_s_cla16_and927_y0(h_s_cla16_and926_y0, h_s_cla16_and925_y0, h_s_cla16_and927_y0);
  and_gate and_gate_h_s_cla16_and928_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and928_y0);
  and_gate and_gate_h_s_cla16_and929_y0(h_s_cla16_and928_y0, h_s_cla16_and927_y0, h_s_cla16_and929_y0);
  and_gate and_gate_h_s_cla16_and930_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and930_y0);
  and_gate and_gate_h_s_cla16_and931_y0(h_s_cla16_and930_y0, h_s_cla16_and929_y0, h_s_cla16_and931_y0);
  and_gate and_gate_h_s_cla16_and932_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and932_y0);
  and_gate and_gate_h_s_cla16_and933_y0(h_s_cla16_and932_y0, h_s_cla16_and931_y0, h_s_cla16_and933_y0);
  and_gate and_gate_h_s_cla16_and934_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and934_y0);
  and_gate and_gate_h_s_cla16_and935_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and935_y0);
  and_gate and_gate_h_s_cla16_and936_y0(h_s_cla16_and935_y0, h_s_cla16_and934_y0, h_s_cla16_and936_y0);
  and_gate and_gate_h_s_cla16_and937_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and937_y0);
  and_gate and_gate_h_s_cla16_and938_y0(h_s_cla16_and937_y0, h_s_cla16_and936_y0, h_s_cla16_and938_y0);
  and_gate and_gate_h_s_cla16_and939_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and939_y0);
  and_gate and_gate_h_s_cla16_and940_y0(h_s_cla16_and939_y0, h_s_cla16_and938_y0, h_s_cla16_and940_y0);
  and_gate and_gate_h_s_cla16_and941_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and941_y0);
  and_gate and_gate_h_s_cla16_and942_y0(h_s_cla16_and941_y0, h_s_cla16_and940_y0, h_s_cla16_and942_y0);
  and_gate and_gate_h_s_cla16_and943_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and943_y0);
  and_gate and_gate_h_s_cla16_and944_y0(h_s_cla16_and943_y0, h_s_cla16_and942_y0, h_s_cla16_and944_y0);
  and_gate and_gate_h_s_cla16_and945_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and945_y0);
  and_gate and_gate_h_s_cla16_and946_y0(h_s_cla16_and945_y0, h_s_cla16_and944_y0, h_s_cla16_and946_y0);
  and_gate and_gate_h_s_cla16_and947_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and947_y0);
  and_gate and_gate_h_s_cla16_and948_y0(h_s_cla16_and947_y0, h_s_cla16_and946_y0, h_s_cla16_and948_y0);
  and_gate and_gate_h_s_cla16_and949_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and949_y0);
  and_gate and_gate_h_s_cla16_and950_y0(h_s_cla16_and949_y0, h_s_cla16_and948_y0, h_s_cla16_and950_y0);
  and_gate and_gate_h_s_cla16_and951_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and951_y0);
  and_gate and_gate_h_s_cla16_and952_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and952_y0);
  and_gate and_gate_h_s_cla16_and953_y0(h_s_cla16_and952_y0, h_s_cla16_and951_y0, h_s_cla16_and953_y0);
  and_gate and_gate_h_s_cla16_and954_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and954_y0);
  and_gate and_gate_h_s_cla16_and955_y0(h_s_cla16_and954_y0, h_s_cla16_and953_y0, h_s_cla16_and955_y0);
  and_gate and_gate_h_s_cla16_and956_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and956_y0);
  and_gate and_gate_h_s_cla16_and957_y0(h_s_cla16_and956_y0, h_s_cla16_and955_y0, h_s_cla16_and957_y0);
  and_gate and_gate_h_s_cla16_and958_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and958_y0);
  and_gate and_gate_h_s_cla16_and959_y0(h_s_cla16_and958_y0, h_s_cla16_and957_y0, h_s_cla16_and959_y0);
  and_gate and_gate_h_s_cla16_and960_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and960_y0);
  and_gate and_gate_h_s_cla16_and961_y0(h_s_cla16_and960_y0, h_s_cla16_and959_y0, h_s_cla16_and961_y0);
  and_gate and_gate_h_s_cla16_and962_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and962_y0);
  and_gate and_gate_h_s_cla16_and963_y0(h_s_cla16_and962_y0, h_s_cla16_and961_y0, h_s_cla16_and963_y0);
  and_gate and_gate_h_s_cla16_and964_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and964_y0);
  and_gate and_gate_h_s_cla16_and965_y0(h_s_cla16_and964_y0, h_s_cla16_and963_y0, h_s_cla16_and965_y0);
  and_gate and_gate_h_s_cla16_and966_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and966_y0);
  and_gate and_gate_h_s_cla16_and967_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and967_y0);
  and_gate and_gate_h_s_cla16_and968_y0(h_s_cla16_and967_y0, h_s_cla16_and966_y0, h_s_cla16_and968_y0);
  and_gate and_gate_h_s_cla16_and969_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and969_y0);
  and_gate and_gate_h_s_cla16_and970_y0(h_s_cla16_and969_y0, h_s_cla16_and968_y0, h_s_cla16_and970_y0);
  and_gate and_gate_h_s_cla16_and971_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and971_y0);
  and_gate and_gate_h_s_cla16_and972_y0(h_s_cla16_and971_y0, h_s_cla16_and970_y0, h_s_cla16_and972_y0);
  and_gate and_gate_h_s_cla16_and973_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and973_y0);
  and_gate and_gate_h_s_cla16_and974_y0(h_s_cla16_and973_y0, h_s_cla16_and972_y0, h_s_cla16_and974_y0);
  and_gate and_gate_h_s_cla16_and975_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and975_y0);
  and_gate and_gate_h_s_cla16_and976_y0(h_s_cla16_and975_y0, h_s_cla16_and974_y0, h_s_cla16_and976_y0);
  and_gate and_gate_h_s_cla16_and977_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and977_y0);
  and_gate and_gate_h_s_cla16_and978_y0(h_s_cla16_and977_y0, h_s_cla16_and976_y0, h_s_cla16_and978_y0);
  and_gate and_gate_h_s_cla16_and979_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and979_y0);
  and_gate and_gate_h_s_cla16_and980_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and980_y0);
  and_gate and_gate_h_s_cla16_and981_y0(h_s_cla16_and980_y0, h_s_cla16_and979_y0, h_s_cla16_and981_y0);
  and_gate and_gate_h_s_cla16_and982_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and982_y0);
  and_gate and_gate_h_s_cla16_and983_y0(h_s_cla16_and982_y0, h_s_cla16_and981_y0, h_s_cla16_and983_y0);
  and_gate and_gate_h_s_cla16_and984_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and984_y0);
  and_gate and_gate_h_s_cla16_and985_y0(h_s_cla16_and984_y0, h_s_cla16_and983_y0, h_s_cla16_and985_y0);
  and_gate and_gate_h_s_cla16_and986_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and986_y0);
  and_gate and_gate_h_s_cla16_and987_y0(h_s_cla16_and986_y0, h_s_cla16_and985_y0, h_s_cla16_and987_y0);
  and_gate and_gate_h_s_cla16_and988_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and988_y0);
  and_gate and_gate_h_s_cla16_and989_y0(h_s_cla16_and988_y0, h_s_cla16_and987_y0, h_s_cla16_and989_y0);
  and_gate and_gate_h_s_cla16_and990_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and990_y0);
  and_gate and_gate_h_s_cla16_and991_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and991_y0);
  and_gate and_gate_h_s_cla16_and992_y0(h_s_cla16_and991_y0, h_s_cla16_and990_y0, h_s_cla16_and992_y0);
  and_gate and_gate_h_s_cla16_and993_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and993_y0);
  and_gate and_gate_h_s_cla16_and994_y0(h_s_cla16_and993_y0, h_s_cla16_and992_y0, h_s_cla16_and994_y0);
  and_gate and_gate_h_s_cla16_and995_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and995_y0);
  and_gate and_gate_h_s_cla16_and996_y0(h_s_cla16_and995_y0, h_s_cla16_and994_y0, h_s_cla16_and996_y0);
  and_gate and_gate_h_s_cla16_and997_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and997_y0);
  and_gate and_gate_h_s_cla16_and998_y0(h_s_cla16_and997_y0, h_s_cla16_and996_y0, h_s_cla16_and998_y0);
  and_gate and_gate_h_s_cla16_and999_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and999_y0);
  and_gate and_gate_h_s_cla16_and1000_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1000_y0);
  and_gate and_gate_h_s_cla16_and1001_y0(h_s_cla16_and1000_y0, h_s_cla16_and999_y0, h_s_cla16_and1001_y0);
  and_gate and_gate_h_s_cla16_and1002_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1002_y0);
  and_gate and_gate_h_s_cla16_and1003_y0(h_s_cla16_and1002_y0, h_s_cla16_and1001_y0, h_s_cla16_and1003_y0);
  and_gate and_gate_h_s_cla16_and1004_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1004_y0);
  and_gate and_gate_h_s_cla16_and1005_y0(h_s_cla16_and1004_y0, h_s_cla16_and1003_y0, h_s_cla16_and1005_y0);
  and_gate and_gate_h_s_cla16_and1006_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1006_y0);
  and_gate and_gate_h_s_cla16_and1007_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1007_y0);
  and_gate and_gate_h_s_cla16_and1008_y0(h_s_cla16_and1007_y0, h_s_cla16_and1006_y0, h_s_cla16_and1008_y0);
  and_gate and_gate_h_s_cla16_and1009_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1009_y0);
  and_gate and_gate_h_s_cla16_and1010_y0(h_s_cla16_and1009_y0, h_s_cla16_and1008_y0, h_s_cla16_and1010_y0);
  and_gate and_gate_h_s_cla16_and1011_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1011_y0);
  and_gate and_gate_h_s_cla16_and1012_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1012_y0);
  and_gate and_gate_h_s_cla16_and1013_y0(h_s_cla16_and1012_y0, h_s_cla16_and1011_y0, h_s_cla16_and1013_y0);
  and_gate and_gate_h_s_cla16_and1014_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic12_y1, h_s_cla16_and1014_y0);
  or_gate or_gate_h_s_cla16_or91_y0(h_s_cla16_and1014_y0, h_s_cla16_and845_y0, h_s_cla16_or91_y0);
  or_gate or_gate_h_s_cla16_or92_y0(h_s_cla16_or91_y0, h_s_cla16_and870_y0, h_s_cla16_or92_y0);
  or_gate or_gate_h_s_cla16_or93_y0(h_s_cla16_or92_y0, h_s_cla16_and893_y0, h_s_cla16_or93_y0);
  or_gate or_gate_h_s_cla16_or94_y0(h_s_cla16_or93_y0, h_s_cla16_and914_y0, h_s_cla16_or94_y0);
  or_gate or_gate_h_s_cla16_or95_y0(h_s_cla16_or94_y0, h_s_cla16_and933_y0, h_s_cla16_or95_y0);
  or_gate or_gate_h_s_cla16_or96_y0(h_s_cla16_or95_y0, h_s_cla16_and950_y0, h_s_cla16_or96_y0);
  or_gate or_gate_h_s_cla16_or97_y0(h_s_cla16_or96_y0, h_s_cla16_and965_y0, h_s_cla16_or97_y0);
  or_gate or_gate_h_s_cla16_or98_y0(h_s_cla16_or97_y0, h_s_cla16_and978_y0, h_s_cla16_or98_y0);
  or_gate or_gate_h_s_cla16_or99_y0(h_s_cla16_or98_y0, h_s_cla16_and989_y0, h_s_cla16_or99_y0);
  or_gate or_gate_h_s_cla16_or100_y0(h_s_cla16_or99_y0, h_s_cla16_and998_y0, h_s_cla16_or100_y0);
  or_gate or_gate_h_s_cla16_or101_y0(h_s_cla16_or100_y0, h_s_cla16_and1005_y0, h_s_cla16_or101_y0);
  or_gate or_gate_h_s_cla16_or102_y0(h_s_cla16_or101_y0, h_s_cla16_and1010_y0, h_s_cla16_or102_y0);
  or_gate or_gate_h_s_cla16_or103_y0(h_s_cla16_or102_y0, h_s_cla16_and1013_y0, h_s_cla16_or103_y0);
  or_gate or_gate_h_s_cla16_or104_y0(h_s_cla16_pg_logic13_y1, h_s_cla16_or103_y0, h_s_cla16_or104_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic14_y0(a_14, b_14, h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic14_y1, h_s_cla16_pg_logic14_y2);
  xor_gate xor_gate_h_s_cla16_xor14_y0(h_s_cla16_pg_logic14_y2, h_s_cla16_or104_y0, h_s_cla16_xor14_y0);
  and_gate and_gate_h_s_cla16_and1015_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and1015_y0);
  and_gate and_gate_h_s_cla16_and1016_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and1016_y0);
  and_gate and_gate_h_s_cla16_and1017_y0(h_s_cla16_and1016_y0, h_s_cla16_and1015_y0, h_s_cla16_and1017_y0);
  and_gate and_gate_h_s_cla16_and1018_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and1018_y0);
  and_gate and_gate_h_s_cla16_and1019_y0(h_s_cla16_and1018_y0, h_s_cla16_and1017_y0, h_s_cla16_and1019_y0);
  and_gate and_gate_h_s_cla16_and1020_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and1020_y0);
  and_gate and_gate_h_s_cla16_and1021_y0(h_s_cla16_and1020_y0, h_s_cla16_and1019_y0, h_s_cla16_and1021_y0);
  and_gate and_gate_h_s_cla16_and1022_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and1022_y0);
  and_gate and_gate_h_s_cla16_and1023_y0(h_s_cla16_and1022_y0, h_s_cla16_and1021_y0, h_s_cla16_and1023_y0);
  and_gate and_gate_h_s_cla16_and1024_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and1024_y0);
  and_gate and_gate_h_s_cla16_and1025_y0(h_s_cla16_and1024_y0, h_s_cla16_and1023_y0, h_s_cla16_and1025_y0);
  and_gate and_gate_h_s_cla16_and1026_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and1026_y0);
  and_gate and_gate_h_s_cla16_and1027_y0(h_s_cla16_and1026_y0, h_s_cla16_and1025_y0, h_s_cla16_and1027_y0);
  and_gate and_gate_h_s_cla16_and1028_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and1028_y0);
  and_gate and_gate_h_s_cla16_and1029_y0(h_s_cla16_and1028_y0, h_s_cla16_and1027_y0, h_s_cla16_and1029_y0);
  and_gate and_gate_h_s_cla16_and1030_y0(h_s_cla16_pg_logic8_y0, constant_wire_0, h_s_cla16_and1030_y0);
  and_gate and_gate_h_s_cla16_and1031_y0(h_s_cla16_and1030_y0, h_s_cla16_and1029_y0, h_s_cla16_and1031_y0);
  and_gate and_gate_h_s_cla16_and1032_y0(h_s_cla16_pg_logic9_y0, constant_wire_0, h_s_cla16_and1032_y0);
  and_gate and_gate_h_s_cla16_and1033_y0(h_s_cla16_and1032_y0, h_s_cla16_and1031_y0, h_s_cla16_and1033_y0);
  and_gate and_gate_h_s_cla16_and1034_y0(h_s_cla16_pg_logic10_y0, constant_wire_0, h_s_cla16_and1034_y0);
  and_gate and_gate_h_s_cla16_and1035_y0(h_s_cla16_and1034_y0, h_s_cla16_and1033_y0, h_s_cla16_and1035_y0);
  and_gate and_gate_h_s_cla16_and1036_y0(h_s_cla16_pg_logic11_y0, constant_wire_0, h_s_cla16_and1036_y0);
  and_gate and_gate_h_s_cla16_and1037_y0(h_s_cla16_and1036_y0, h_s_cla16_and1035_y0, h_s_cla16_and1037_y0);
  and_gate and_gate_h_s_cla16_and1038_y0(h_s_cla16_pg_logic12_y0, constant_wire_0, h_s_cla16_and1038_y0);
  and_gate and_gate_h_s_cla16_and1039_y0(h_s_cla16_and1038_y0, h_s_cla16_and1037_y0, h_s_cla16_and1039_y0);
  and_gate and_gate_h_s_cla16_and1040_y0(h_s_cla16_pg_logic13_y0, constant_wire_0, h_s_cla16_and1040_y0);
  and_gate and_gate_h_s_cla16_and1041_y0(h_s_cla16_and1040_y0, h_s_cla16_and1039_y0, h_s_cla16_and1041_y0);
  and_gate and_gate_h_s_cla16_and1042_y0(h_s_cla16_pg_logic14_y0, constant_wire_0, h_s_cla16_and1042_y0);
  and_gate and_gate_h_s_cla16_and1043_y0(h_s_cla16_and1042_y0, h_s_cla16_and1041_y0, h_s_cla16_and1043_y0);
  and_gate and_gate_h_s_cla16_and1044_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1044_y0);
  and_gate and_gate_h_s_cla16_and1045_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1045_y0);
  and_gate and_gate_h_s_cla16_and1046_y0(h_s_cla16_and1045_y0, h_s_cla16_and1044_y0, h_s_cla16_and1046_y0);
  and_gate and_gate_h_s_cla16_and1047_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1047_y0);
  and_gate and_gate_h_s_cla16_and1048_y0(h_s_cla16_and1047_y0, h_s_cla16_and1046_y0, h_s_cla16_and1048_y0);
  and_gate and_gate_h_s_cla16_and1049_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1049_y0);
  and_gate and_gate_h_s_cla16_and1050_y0(h_s_cla16_and1049_y0, h_s_cla16_and1048_y0, h_s_cla16_and1050_y0);
  and_gate and_gate_h_s_cla16_and1051_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1051_y0);
  and_gate and_gate_h_s_cla16_and1052_y0(h_s_cla16_and1051_y0, h_s_cla16_and1050_y0, h_s_cla16_and1052_y0);
  and_gate and_gate_h_s_cla16_and1053_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1053_y0);
  and_gate and_gate_h_s_cla16_and1054_y0(h_s_cla16_and1053_y0, h_s_cla16_and1052_y0, h_s_cla16_and1054_y0);
  and_gate and_gate_h_s_cla16_and1055_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1055_y0);
  and_gate and_gate_h_s_cla16_and1056_y0(h_s_cla16_and1055_y0, h_s_cla16_and1054_y0, h_s_cla16_and1056_y0);
  and_gate and_gate_h_s_cla16_and1057_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1057_y0);
  and_gate and_gate_h_s_cla16_and1058_y0(h_s_cla16_and1057_y0, h_s_cla16_and1056_y0, h_s_cla16_and1058_y0);
  and_gate and_gate_h_s_cla16_and1059_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1059_y0);
  and_gate and_gate_h_s_cla16_and1060_y0(h_s_cla16_and1059_y0, h_s_cla16_and1058_y0, h_s_cla16_and1060_y0);
  and_gate and_gate_h_s_cla16_and1061_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1061_y0);
  and_gate and_gate_h_s_cla16_and1062_y0(h_s_cla16_and1061_y0, h_s_cla16_and1060_y0, h_s_cla16_and1062_y0);
  and_gate and_gate_h_s_cla16_and1063_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1063_y0);
  and_gate and_gate_h_s_cla16_and1064_y0(h_s_cla16_and1063_y0, h_s_cla16_and1062_y0, h_s_cla16_and1064_y0);
  and_gate and_gate_h_s_cla16_and1065_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1065_y0);
  and_gate and_gate_h_s_cla16_and1066_y0(h_s_cla16_and1065_y0, h_s_cla16_and1064_y0, h_s_cla16_and1066_y0);
  and_gate and_gate_h_s_cla16_and1067_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1067_y0);
  and_gate and_gate_h_s_cla16_and1068_y0(h_s_cla16_and1067_y0, h_s_cla16_and1066_y0, h_s_cla16_and1068_y0);
  and_gate and_gate_h_s_cla16_and1069_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1069_y0);
  and_gate and_gate_h_s_cla16_and1070_y0(h_s_cla16_and1069_y0, h_s_cla16_and1068_y0, h_s_cla16_and1070_y0);
  and_gate and_gate_h_s_cla16_and1071_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1071_y0);
  and_gate and_gate_h_s_cla16_and1072_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1072_y0);
  and_gate and_gate_h_s_cla16_and1073_y0(h_s_cla16_and1072_y0, h_s_cla16_and1071_y0, h_s_cla16_and1073_y0);
  and_gate and_gate_h_s_cla16_and1074_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1074_y0);
  and_gate and_gate_h_s_cla16_and1075_y0(h_s_cla16_and1074_y0, h_s_cla16_and1073_y0, h_s_cla16_and1075_y0);
  and_gate and_gate_h_s_cla16_and1076_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1076_y0);
  and_gate and_gate_h_s_cla16_and1077_y0(h_s_cla16_and1076_y0, h_s_cla16_and1075_y0, h_s_cla16_and1077_y0);
  and_gate and_gate_h_s_cla16_and1078_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1078_y0);
  and_gate and_gate_h_s_cla16_and1079_y0(h_s_cla16_and1078_y0, h_s_cla16_and1077_y0, h_s_cla16_and1079_y0);
  and_gate and_gate_h_s_cla16_and1080_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1080_y0);
  and_gate and_gate_h_s_cla16_and1081_y0(h_s_cla16_and1080_y0, h_s_cla16_and1079_y0, h_s_cla16_and1081_y0);
  and_gate and_gate_h_s_cla16_and1082_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1082_y0);
  and_gate and_gate_h_s_cla16_and1083_y0(h_s_cla16_and1082_y0, h_s_cla16_and1081_y0, h_s_cla16_and1083_y0);
  and_gate and_gate_h_s_cla16_and1084_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1084_y0);
  and_gate and_gate_h_s_cla16_and1085_y0(h_s_cla16_and1084_y0, h_s_cla16_and1083_y0, h_s_cla16_and1085_y0);
  and_gate and_gate_h_s_cla16_and1086_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1086_y0);
  and_gate and_gate_h_s_cla16_and1087_y0(h_s_cla16_and1086_y0, h_s_cla16_and1085_y0, h_s_cla16_and1087_y0);
  and_gate and_gate_h_s_cla16_and1088_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1088_y0);
  and_gate and_gate_h_s_cla16_and1089_y0(h_s_cla16_and1088_y0, h_s_cla16_and1087_y0, h_s_cla16_and1089_y0);
  and_gate and_gate_h_s_cla16_and1090_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1090_y0);
  and_gate and_gate_h_s_cla16_and1091_y0(h_s_cla16_and1090_y0, h_s_cla16_and1089_y0, h_s_cla16_and1091_y0);
  and_gate and_gate_h_s_cla16_and1092_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1092_y0);
  and_gate and_gate_h_s_cla16_and1093_y0(h_s_cla16_and1092_y0, h_s_cla16_and1091_y0, h_s_cla16_and1093_y0);
  and_gate and_gate_h_s_cla16_and1094_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1094_y0);
  and_gate and_gate_h_s_cla16_and1095_y0(h_s_cla16_and1094_y0, h_s_cla16_and1093_y0, h_s_cla16_and1095_y0);
  and_gate and_gate_h_s_cla16_and1096_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1096_y0);
  and_gate and_gate_h_s_cla16_and1097_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1097_y0);
  and_gate and_gate_h_s_cla16_and1098_y0(h_s_cla16_and1097_y0, h_s_cla16_and1096_y0, h_s_cla16_and1098_y0);
  and_gate and_gate_h_s_cla16_and1099_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1099_y0);
  and_gate and_gate_h_s_cla16_and1100_y0(h_s_cla16_and1099_y0, h_s_cla16_and1098_y0, h_s_cla16_and1100_y0);
  and_gate and_gate_h_s_cla16_and1101_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1101_y0);
  and_gate and_gate_h_s_cla16_and1102_y0(h_s_cla16_and1101_y0, h_s_cla16_and1100_y0, h_s_cla16_and1102_y0);
  and_gate and_gate_h_s_cla16_and1103_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1103_y0);
  and_gate and_gate_h_s_cla16_and1104_y0(h_s_cla16_and1103_y0, h_s_cla16_and1102_y0, h_s_cla16_and1104_y0);
  and_gate and_gate_h_s_cla16_and1105_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1105_y0);
  and_gate and_gate_h_s_cla16_and1106_y0(h_s_cla16_and1105_y0, h_s_cla16_and1104_y0, h_s_cla16_and1106_y0);
  and_gate and_gate_h_s_cla16_and1107_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1107_y0);
  and_gate and_gate_h_s_cla16_and1108_y0(h_s_cla16_and1107_y0, h_s_cla16_and1106_y0, h_s_cla16_and1108_y0);
  and_gate and_gate_h_s_cla16_and1109_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1109_y0);
  and_gate and_gate_h_s_cla16_and1110_y0(h_s_cla16_and1109_y0, h_s_cla16_and1108_y0, h_s_cla16_and1110_y0);
  and_gate and_gate_h_s_cla16_and1111_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1111_y0);
  and_gate and_gate_h_s_cla16_and1112_y0(h_s_cla16_and1111_y0, h_s_cla16_and1110_y0, h_s_cla16_and1112_y0);
  and_gate and_gate_h_s_cla16_and1113_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1113_y0);
  and_gate and_gate_h_s_cla16_and1114_y0(h_s_cla16_and1113_y0, h_s_cla16_and1112_y0, h_s_cla16_and1114_y0);
  and_gate and_gate_h_s_cla16_and1115_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1115_y0);
  and_gate and_gate_h_s_cla16_and1116_y0(h_s_cla16_and1115_y0, h_s_cla16_and1114_y0, h_s_cla16_and1116_y0);
  and_gate and_gate_h_s_cla16_and1117_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1117_y0);
  and_gate and_gate_h_s_cla16_and1118_y0(h_s_cla16_and1117_y0, h_s_cla16_and1116_y0, h_s_cla16_and1118_y0);
  and_gate and_gate_h_s_cla16_and1119_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1119_y0);
  and_gate and_gate_h_s_cla16_and1120_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1120_y0);
  and_gate and_gate_h_s_cla16_and1121_y0(h_s_cla16_and1120_y0, h_s_cla16_and1119_y0, h_s_cla16_and1121_y0);
  and_gate and_gate_h_s_cla16_and1122_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1122_y0);
  and_gate and_gate_h_s_cla16_and1123_y0(h_s_cla16_and1122_y0, h_s_cla16_and1121_y0, h_s_cla16_and1123_y0);
  and_gate and_gate_h_s_cla16_and1124_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1124_y0);
  and_gate and_gate_h_s_cla16_and1125_y0(h_s_cla16_and1124_y0, h_s_cla16_and1123_y0, h_s_cla16_and1125_y0);
  and_gate and_gate_h_s_cla16_and1126_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1126_y0);
  and_gate and_gate_h_s_cla16_and1127_y0(h_s_cla16_and1126_y0, h_s_cla16_and1125_y0, h_s_cla16_and1127_y0);
  and_gate and_gate_h_s_cla16_and1128_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1128_y0);
  and_gate and_gate_h_s_cla16_and1129_y0(h_s_cla16_and1128_y0, h_s_cla16_and1127_y0, h_s_cla16_and1129_y0);
  and_gate and_gate_h_s_cla16_and1130_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1130_y0);
  and_gate and_gate_h_s_cla16_and1131_y0(h_s_cla16_and1130_y0, h_s_cla16_and1129_y0, h_s_cla16_and1131_y0);
  and_gate and_gate_h_s_cla16_and1132_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1132_y0);
  and_gate and_gate_h_s_cla16_and1133_y0(h_s_cla16_and1132_y0, h_s_cla16_and1131_y0, h_s_cla16_and1133_y0);
  and_gate and_gate_h_s_cla16_and1134_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1134_y0);
  and_gate and_gate_h_s_cla16_and1135_y0(h_s_cla16_and1134_y0, h_s_cla16_and1133_y0, h_s_cla16_and1135_y0);
  and_gate and_gate_h_s_cla16_and1136_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1136_y0);
  and_gate and_gate_h_s_cla16_and1137_y0(h_s_cla16_and1136_y0, h_s_cla16_and1135_y0, h_s_cla16_and1137_y0);
  and_gate and_gate_h_s_cla16_and1138_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1138_y0);
  and_gate and_gate_h_s_cla16_and1139_y0(h_s_cla16_and1138_y0, h_s_cla16_and1137_y0, h_s_cla16_and1139_y0);
  and_gate and_gate_h_s_cla16_and1140_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1140_y0);
  and_gate and_gate_h_s_cla16_and1141_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1141_y0);
  and_gate and_gate_h_s_cla16_and1142_y0(h_s_cla16_and1141_y0, h_s_cla16_and1140_y0, h_s_cla16_and1142_y0);
  and_gate and_gate_h_s_cla16_and1143_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1143_y0);
  and_gate and_gate_h_s_cla16_and1144_y0(h_s_cla16_and1143_y0, h_s_cla16_and1142_y0, h_s_cla16_and1144_y0);
  and_gate and_gate_h_s_cla16_and1145_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1145_y0);
  and_gate and_gate_h_s_cla16_and1146_y0(h_s_cla16_and1145_y0, h_s_cla16_and1144_y0, h_s_cla16_and1146_y0);
  and_gate and_gate_h_s_cla16_and1147_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1147_y0);
  and_gate and_gate_h_s_cla16_and1148_y0(h_s_cla16_and1147_y0, h_s_cla16_and1146_y0, h_s_cla16_and1148_y0);
  and_gate and_gate_h_s_cla16_and1149_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1149_y0);
  and_gate and_gate_h_s_cla16_and1150_y0(h_s_cla16_and1149_y0, h_s_cla16_and1148_y0, h_s_cla16_and1150_y0);
  and_gate and_gate_h_s_cla16_and1151_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1151_y0);
  and_gate and_gate_h_s_cla16_and1152_y0(h_s_cla16_and1151_y0, h_s_cla16_and1150_y0, h_s_cla16_and1152_y0);
  and_gate and_gate_h_s_cla16_and1153_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1153_y0);
  and_gate and_gate_h_s_cla16_and1154_y0(h_s_cla16_and1153_y0, h_s_cla16_and1152_y0, h_s_cla16_and1154_y0);
  and_gate and_gate_h_s_cla16_and1155_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1155_y0);
  and_gate and_gate_h_s_cla16_and1156_y0(h_s_cla16_and1155_y0, h_s_cla16_and1154_y0, h_s_cla16_and1156_y0);
  and_gate and_gate_h_s_cla16_and1157_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1157_y0);
  and_gate and_gate_h_s_cla16_and1158_y0(h_s_cla16_and1157_y0, h_s_cla16_and1156_y0, h_s_cla16_and1158_y0);
  and_gate and_gate_h_s_cla16_and1159_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1159_y0);
  and_gate and_gate_h_s_cla16_and1160_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1160_y0);
  and_gate and_gate_h_s_cla16_and1161_y0(h_s_cla16_and1160_y0, h_s_cla16_and1159_y0, h_s_cla16_and1161_y0);
  and_gate and_gate_h_s_cla16_and1162_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1162_y0);
  and_gate and_gate_h_s_cla16_and1163_y0(h_s_cla16_and1162_y0, h_s_cla16_and1161_y0, h_s_cla16_and1163_y0);
  and_gate and_gate_h_s_cla16_and1164_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1164_y0);
  and_gate and_gate_h_s_cla16_and1165_y0(h_s_cla16_and1164_y0, h_s_cla16_and1163_y0, h_s_cla16_and1165_y0);
  and_gate and_gate_h_s_cla16_and1166_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1166_y0);
  and_gate and_gate_h_s_cla16_and1167_y0(h_s_cla16_and1166_y0, h_s_cla16_and1165_y0, h_s_cla16_and1167_y0);
  and_gate and_gate_h_s_cla16_and1168_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1168_y0);
  and_gate and_gate_h_s_cla16_and1169_y0(h_s_cla16_and1168_y0, h_s_cla16_and1167_y0, h_s_cla16_and1169_y0);
  and_gate and_gate_h_s_cla16_and1170_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1170_y0);
  and_gate and_gate_h_s_cla16_and1171_y0(h_s_cla16_and1170_y0, h_s_cla16_and1169_y0, h_s_cla16_and1171_y0);
  and_gate and_gate_h_s_cla16_and1172_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1172_y0);
  and_gate and_gate_h_s_cla16_and1173_y0(h_s_cla16_and1172_y0, h_s_cla16_and1171_y0, h_s_cla16_and1173_y0);
  and_gate and_gate_h_s_cla16_and1174_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1174_y0);
  and_gate and_gate_h_s_cla16_and1175_y0(h_s_cla16_and1174_y0, h_s_cla16_and1173_y0, h_s_cla16_and1175_y0);
  and_gate and_gate_h_s_cla16_and1176_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1176_y0);
  and_gate and_gate_h_s_cla16_and1177_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1177_y0);
  and_gate and_gate_h_s_cla16_and1178_y0(h_s_cla16_and1177_y0, h_s_cla16_and1176_y0, h_s_cla16_and1178_y0);
  and_gate and_gate_h_s_cla16_and1179_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1179_y0);
  and_gate and_gate_h_s_cla16_and1180_y0(h_s_cla16_and1179_y0, h_s_cla16_and1178_y0, h_s_cla16_and1180_y0);
  and_gate and_gate_h_s_cla16_and1181_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1181_y0);
  and_gate and_gate_h_s_cla16_and1182_y0(h_s_cla16_and1181_y0, h_s_cla16_and1180_y0, h_s_cla16_and1182_y0);
  and_gate and_gate_h_s_cla16_and1183_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1183_y0);
  and_gate and_gate_h_s_cla16_and1184_y0(h_s_cla16_and1183_y0, h_s_cla16_and1182_y0, h_s_cla16_and1184_y0);
  and_gate and_gate_h_s_cla16_and1185_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1185_y0);
  and_gate and_gate_h_s_cla16_and1186_y0(h_s_cla16_and1185_y0, h_s_cla16_and1184_y0, h_s_cla16_and1186_y0);
  and_gate and_gate_h_s_cla16_and1187_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1187_y0);
  and_gate and_gate_h_s_cla16_and1188_y0(h_s_cla16_and1187_y0, h_s_cla16_and1186_y0, h_s_cla16_and1188_y0);
  and_gate and_gate_h_s_cla16_and1189_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1189_y0);
  and_gate and_gate_h_s_cla16_and1190_y0(h_s_cla16_and1189_y0, h_s_cla16_and1188_y0, h_s_cla16_and1190_y0);
  and_gate and_gate_h_s_cla16_and1191_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1191_y0);
  and_gate and_gate_h_s_cla16_and1192_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1192_y0);
  and_gate and_gate_h_s_cla16_and1193_y0(h_s_cla16_and1192_y0, h_s_cla16_and1191_y0, h_s_cla16_and1193_y0);
  and_gate and_gate_h_s_cla16_and1194_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1194_y0);
  and_gate and_gate_h_s_cla16_and1195_y0(h_s_cla16_and1194_y0, h_s_cla16_and1193_y0, h_s_cla16_and1195_y0);
  and_gate and_gate_h_s_cla16_and1196_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1196_y0);
  and_gate and_gate_h_s_cla16_and1197_y0(h_s_cla16_and1196_y0, h_s_cla16_and1195_y0, h_s_cla16_and1197_y0);
  and_gate and_gate_h_s_cla16_and1198_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1198_y0);
  and_gate and_gate_h_s_cla16_and1199_y0(h_s_cla16_and1198_y0, h_s_cla16_and1197_y0, h_s_cla16_and1199_y0);
  and_gate and_gate_h_s_cla16_and1200_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1200_y0);
  and_gate and_gate_h_s_cla16_and1201_y0(h_s_cla16_and1200_y0, h_s_cla16_and1199_y0, h_s_cla16_and1201_y0);
  and_gate and_gate_h_s_cla16_and1202_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1202_y0);
  and_gate and_gate_h_s_cla16_and1203_y0(h_s_cla16_and1202_y0, h_s_cla16_and1201_y0, h_s_cla16_and1203_y0);
  and_gate and_gate_h_s_cla16_and1204_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1204_y0);
  and_gate and_gate_h_s_cla16_and1205_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1205_y0);
  and_gate and_gate_h_s_cla16_and1206_y0(h_s_cla16_and1205_y0, h_s_cla16_and1204_y0, h_s_cla16_and1206_y0);
  and_gate and_gate_h_s_cla16_and1207_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1207_y0);
  and_gate and_gate_h_s_cla16_and1208_y0(h_s_cla16_and1207_y0, h_s_cla16_and1206_y0, h_s_cla16_and1208_y0);
  and_gate and_gate_h_s_cla16_and1209_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1209_y0);
  and_gate and_gate_h_s_cla16_and1210_y0(h_s_cla16_and1209_y0, h_s_cla16_and1208_y0, h_s_cla16_and1210_y0);
  and_gate and_gate_h_s_cla16_and1211_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1211_y0);
  and_gate and_gate_h_s_cla16_and1212_y0(h_s_cla16_and1211_y0, h_s_cla16_and1210_y0, h_s_cla16_and1212_y0);
  and_gate and_gate_h_s_cla16_and1213_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1213_y0);
  and_gate and_gate_h_s_cla16_and1214_y0(h_s_cla16_and1213_y0, h_s_cla16_and1212_y0, h_s_cla16_and1214_y0);
  and_gate and_gate_h_s_cla16_and1215_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1215_y0);
  and_gate and_gate_h_s_cla16_and1216_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1216_y0);
  and_gate and_gate_h_s_cla16_and1217_y0(h_s_cla16_and1216_y0, h_s_cla16_and1215_y0, h_s_cla16_and1217_y0);
  and_gate and_gate_h_s_cla16_and1218_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1218_y0);
  and_gate and_gate_h_s_cla16_and1219_y0(h_s_cla16_and1218_y0, h_s_cla16_and1217_y0, h_s_cla16_and1219_y0);
  and_gate and_gate_h_s_cla16_and1220_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1220_y0);
  and_gate and_gate_h_s_cla16_and1221_y0(h_s_cla16_and1220_y0, h_s_cla16_and1219_y0, h_s_cla16_and1221_y0);
  and_gate and_gate_h_s_cla16_and1222_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1222_y0);
  and_gate and_gate_h_s_cla16_and1223_y0(h_s_cla16_and1222_y0, h_s_cla16_and1221_y0, h_s_cla16_and1223_y0);
  and_gate and_gate_h_s_cla16_and1224_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1224_y0);
  and_gate and_gate_h_s_cla16_and1225_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1225_y0);
  and_gate and_gate_h_s_cla16_and1226_y0(h_s_cla16_and1225_y0, h_s_cla16_and1224_y0, h_s_cla16_and1226_y0);
  and_gate and_gate_h_s_cla16_and1227_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1227_y0);
  and_gate and_gate_h_s_cla16_and1228_y0(h_s_cla16_and1227_y0, h_s_cla16_and1226_y0, h_s_cla16_and1228_y0);
  and_gate and_gate_h_s_cla16_and1229_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1229_y0);
  and_gate and_gate_h_s_cla16_and1230_y0(h_s_cla16_and1229_y0, h_s_cla16_and1228_y0, h_s_cla16_and1230_y0);
  and_gate and_gate_h_s_cla16_and1231_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1231_y0);
  and_gate and_gate_h_s_cla16_and1232_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1232_y0);
  and_gate and_gate_h_s_cla16_and1233_y0(h_s_cla16_and1232_y0, h_s_cla16_and1231_y0, h_s_cla16_and1233_y0);
  and_gate and_gate_h_s_cla16_and1234_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1234_y0);
  and_gate and_gate_h_s_cla16_and1235_y0(h_s_cla16_and1234_y0, h_s_cla16_and1233_y0, h_s_cla16_and1235_y0);
  and_gate and_gate_h_s_cla16_and1236_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic12_y1, h_s_cla16_and1236_y0);
  and_gate and_gate_h_s_cla16_and1237_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic12_y1, h_s_cla16_and1237_y0);
  and_gate and_gate_h_s_cla16_and1238_y0(h_s_cla16_and1237_y0, h_s_cla16_and1236_y0, h_s_cla16_and1238_y0);
  and_gate and_gate_h_s_cla16_and1239_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic13_y1, h_s_cla16_and1239_y0);
  or_gate or_gate_h_s_cla16_or105_y0(h_s_cla16_and1239_y0, h_s_cla16_and1043_y0, h_s_cla16_or105_y0);
  or_gate or_gate_h_s_cla16_or106_y0(h_s_cla16_or105_y0, h_s_cla16_and1070_y0, h_s_cla16_or106_y0);
  or_gate or_gate_h_s_cla16_or107_y0(h_s_cla16_or106_y0, h_s_cla16_and1095_y0, h_s_cla16_or107_y0);
  or_gate or_gate_h_s_cla16_or108_y0(h_s_cla16_or107_y0, h_s_cla16_and1118_y0, h_s_cla16_or108_y0);
  or_gate or_gate_h_s_cla16_or109_y0(h_s_cla16_or108_y0, h_s_cla16_and1139_y0, h_s_cla16_or109_y0);
  or_gate or_gate_h_s_cla16_or110_y0(h_s_cla16_or109_y0, h_s_cla16_and1158_y0, h_s_cla16_or110_y0);
  or_gate or_gate_h_s_cla16_or111_y0(h_s_cla16_or110_y0, h_s_cla16_and1175_y0, h_s_cla16_or111_y0);
  or_gate or_gate_h_s_cla16_or112_y0(h_s_cla16_or111_y0, h_s_cla16_and1190_y0, h_s_cla16_or112_y0);
  or_gate or_gate_h_s_cla16_or113_y0(h_s_cla16_or112_y0, h_s_cla16_and1203_y0, h_s_cla16_or113_y0);
  or_gate or_gate_h_s_cla16_or114_y0(h_s_cla16_or113_y0, h_s_cla16_and1214_y0, h_s_cla16_or114_y0);
  or_gate or_gate_h_s_cla16_or115_y0(h_s_cla16_or114_y0, h_s_cla16_and1223_y0, h_s_cla16_or115_y0);
  or_gate or_gate_h_s_cla16_or116_y0(h_s_cla16_or115_y0, h_s_cla16_and1230_y0, h_s_cla16_or116_y0);
  or_gate or_gate_h_s_cla16_or117_y0(h_s_cla16_or116_y0, h_s_cla16_and1235_y0, h_s_cla16_or117_y0);
  or_gate or_gate_h_s_cla16_or118_y0(h_s_cla16_or117_y0, h_s_cla16_and1238_y0, h_s_cla16_or118_y0);
  or_gate or_gate_h_s_cla16_or119_y0(h_s_cla16_pg_logic14_y1, h_s_cla16_or118_y0, h_s_cla16_or119_y0);
  pg_logic pg_logic_h_s_cla16_pg_logic15_y0(a_15, b_15, h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic15_y1, h_s_cla16_pg_logic15_y2);
  xor_gate xor_gate_h_s_cla16_xor15_y0(h_s_cla16_pg_logic15_y2, h_s_cla16_or119_y0, h_s_cla16_xor15_y0);
  and_gate and_gate_h_s_cla16_and1240_y0(h_s_cla16_pg_logic0_y0, constant_wire_0, h_s_cla16_and1240_y0);
  and_gate and_gate_h_s_cla16_and1241_y0(h_s_cla16_pg_logic1_y0, constant_wire_0, h_s_cla16_and1241_y0);
  and_gate and_gate_h_s_cla16_and1242_y0(h_s_cla16_and1241_y0, h_s_cla16_and1240_y0, h_s_cla16_and1242_y0);
  and_gate and_gate_h_s_cla16_and1243_y0(h_s_cla16_pg_logic2_y0, constant_wire_0, h_s_cla16_and1243_y0);
  and_gate and_gate_h_s_cla16_and1244_y0(h_s_cla16_and1243_y0, h_s_cla16_and1242_y0, h_s_cla16_and1244_y0);
  and_gate and_gate_h_s_cla16_and1245_y0(h_s_cla16_pg_logic3_y0, constant_wire_0, h_s_cla16_and1245_y0);
  and_gate and_gate_h_s_cla16_and1246_y0(h_s_cla16_and1245_y0, h_s_cla16_and1244_y0, h_s_cla16_and1246_y0);
  and_gate and_gate_h_s_cla16_and1247_y0(h_s_cla16_pg_logic4_y0, constant_wire_0, h_s_cla16_and1247_y0);
  and_gate and_gate_h_s_cla16_and1248_y0(h_s_cla16_and1247_y0, h_s_cla16_and1246_y0, h_s_cla16_and1248_y0);
  and_gate and_gate_h_s_cla16_and1249_y0(h_s_cla16_pg_logic5_y0, constant_wire_0, h_s_cla16_and1249_y0);
  and_gate and_gate_h_s_cla16_and1250_y0(h_s_cla16_and1249_y0, h_s_cla16_and1248_y0, h_s_cla16_and1250_y0);
  and_gate and_gate_h_s_cla16_and1251_y0(h_s_cla16_pg_logic6_y0, constant_wire_0, h_s_cla16_and1251_y0);
  and_gate and_gate_h_s_cla16_and1252_y0(h_s_cla16_and1251_y0, h_s_cla16_and1250_y0, h_s_cla16_and1252_y0);
  and_gate and_gate_h_s_cla16_and1253_y0(h_s_cla16_pg_logic7_y0, constant_wire_0, h_s_cla16_and1253_y0);
  and_gate and_gate_h_s_cla16_and1254_y0(h_s_cla16_and1253_y0, h_s_cla16_and1252_y0, h_s_cla16_and1254_y0);
  and_gate and_gate_h_s_cla16_and1255_y0(h_s_cla16_pg_logic8_y0, constant_wire_0, h_s_cla16_and1255_y0);
  and_gate and_gate_h_s_cla16_and1256_y0(h_s_cla16_and1255_y0, h_s_cla16_and1254_y0, h_s_cla16_and1256_y0);
  and_gate and_gate_h_s_cla16_and1257_y0(h_s_cla16_pg_logic9_y0, constant_wire_0, h_s_cla16_and1257_y0);
  and_gate and_gate_h_s_cla16_and1258_y0(h_s_cla16_and1257_y0, h_s_cla16_and1256_y0, h_s_cla16_and1258_y0);
  and_gate and_gate_h_s_cla16_and1259_y0(h_s_cla16_pg_logic10_y0, constant_wire_0, h_s_cla16_and1259_y0);
  and_gate and_gate_h_s_cla16_and1260_y0(h_s_cla16_and1259_y0, h_s_cla16_and1258_y0, h_s_cla16_and1260_y0);
  and_gate and_gate_h_s_cla16_and1261_y0(h_s_cla16_pg_logic11_y0, constant_wire_0, h_s_cla16_and1261_y0);
  and_gate and_gate_h_s_cla16_and1262_y0(h_s_cla16_and1261_y0, h_s_cla16_and1260_y0, h_s_cla16_and1262_y0);
  and_gate and_gate_h_s_cla16_and1263_y0(h_s_cla16_pg_logic12_y0, constant_wire_0, h_s_cla16_and1263_y0);
  and_gate and_gate_h_s_cla16_and1264_y0(h_s_cla16_and1263_y0, h_s_cla16_and1262_y0, h_s_cla16_and1264_y0);
  and_gate and_gate_h_s_cla16_and1265_y0(h_s_cla16_pg_logic13_y0, constant_wire_0, h_s_cla16_and1265_y0);
  and_gate and_gate_h_s_cla16_and1266_y0(h_s_cla16_and1265_y0, h_s_cla16_and1264_y0, h_s_cla16_and1266_y0);
  and_gate and_gate_h_s_cla16_and1267_y0(h_s_cla16_pg_logic14_y0, constant_wire_0, h_s_cla16_and1267_y0);
  and_gate and_gate_h_s_cla16_and1268_y0(h_s_cla16_and1267_y0, h_s_cla16_and1266_y0, h_s_cla16_and1268_y0);
  and_gate and_gate_h_s_cla16_and1269_y0(h_s_cla16_pg_logic15_y0, constant_wire_0, h_s_cla16_and1269_y0);
  and_gate and_gate_h_s_cla16_and1270_y0(h_s_cla16_and1269_y0, h_s_cla16_and1268_y0, h_s_cla16_and1270_y0);
  and_gate and_gate_h_s_cla16_and1271_y0(h_s_cla16_pg_logic1_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1271_y0);
  and_gate and_gate_h_s_cla16_and1272_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1272_y0);
  and_gate and_gate_h_s_cla16_and1273_y0(h_s_cla16_and1272_y0, h_s_cla16_and1271_y0, h_s_cla16_and1273_y0);
  and_gate and_gate_h_s_cla16_and1274_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1274_y0);
  and_gate and_gate_h_s_cla16_and1275_y0(h_s_cla16_and1274_y0, h_s_cla16_and1273_y0, h_s_cla16_and1275_y0);
  and_gate and_gate_h_s_cla16_and1276_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1276_y0);
  and_gate and_gate_h_s_cla16_and1277_y0(h_s_cla16_and1276_y0, h_s_cla16_and1275_y0, h_s_cla16_and1277_y0);
  and_gate and_gate_h_s_cla16_and1278_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1278_y0);
  and_gate and_gate_h_s_cla16_and1279_y0(h_s_cla16_and1278_y0, h_s_cla16_and1277_y0, h_s_cla16_and1279_y0);
  and_gate and_gate_h_s_cla16_and1280_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1280_y0);
  and_gate and_gate_h_s_cla16_and1281_y0(h_s_cla16_and1280_y0, h_s_cla16_and1279_y0, h_s_cla16_and1281_y0);
  and_gate and_gate_h_s_cla16_and1282_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1282_y0);
  and_gate and_gate_h_s_cla16_and1283_y0(h_s_cla16_and1282_y0, h_s_cla16_and1281_y0, h_s_cla16_and1283_y0);
  and_gate and_gate_h_s_cla16_and1284_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1284_y0);
  and_gate and_gate_h_s_cla16_and1285_y0(h_s_cla16_and1284_y0, h_s_cla16_and1283_y0, h_s_cla16_and1285_y0);
  and_gate and_gate_h_s_cla16_and1286_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1286_y0);
  and_gate and_gate_h_s_cla16_and1287_y0(h_s_cla16_and1286_y0, h_s_cla16_and1285_y0, h_s_cla16_and1287_y0);
  and_gate and_gate_h_s_cla16_and1288_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1288_y0);
  and_gate and_gate_h_s_cla16_and1289_y0(h_s_cla16_and1288_y0, h_s_cla16_and1287_y0, h_s_cla16_and1289_y0);
  and_gate and_gate_h_s_cla16_and1290_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1290_y0);
  and_gate and_gate_h_s_cla16_and1291_y0(h_s_cla16_and1290_y0, h_s_cla16_and1289_y0, h_s_cla16_and1291_y0);
  and_gate and_gate_h_s_cla16_and1292_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1292_y0);
  and_gate and_gate_h_s_cla16_and1293_y0(h_s_cla16_and1292_y0, h_s_cla16_and1291_y0, h_s_cla16_and1293_y0);
  and_gate and_gate_h_s_cla16_and1294_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1294_y0);
  and_gate and_gate_h_s_cla16_and1295_y0(h_s_cla16_and1294_y0, h_s_cla16_and1293_y0, h_s_cla16_and1295_y0);
  and_gate and_gate_h_s_cla16_and1296_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1296_y0);
  and_gate and_gate_h_s_cla16_and1297_y0(h_s_cla16_and1296_y0, h_s_cla16_and1295_y0, h_s_cla16_and1297_y0);
  and_gate and_gate_h_s_cla16_and1298_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic0_y1, h_s_cla16_and1298_y0);
  and_gate and_gate_h_s_cla16_and1299_y0(h_s_cla16_and1298_y0, h_s_cla16_and1297_y0, h_s_cla16_and1299_y0);
  and_gate and_gate_h_s_cla16_and1300_y0(h_s_cla16_pg_logic2_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1300_y0);
  and_gate and_gate_h_s_cla16_and1301_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1301_y0);
  and_gate and_gate_h_s_cla16_and1302_y0(h_s_cla16_and1301_y0, h_s_cla16_and1300_y0, h_s_cla16_and1302_y0);
  and_gate and_gate_h_s_cla16_and1303_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1303_y0);
  and_gate and_gate_h_s_cla16_and1304_y0(h_s_cla16_and1303_y0, h_s_cla16_and1302_y0, h_s_cla16_and1304_y0);
  and_gate and_gate_h_s_cla16_and1305_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1305_y0);
  and_gate and_gate_h_s_cla16_and1306_y0(h_s_cla16_and1305_y0, h_s_cla16_and1304_y0, h_s_cla16_and1306_y0);
  and_gate and_gate_h_s_cla16_and1307_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1307_y0);
  and_gate and_gate_h_s_cla16_and1308_y0(h_s_cla16_and1307_y0, h_s_cla16_and1306_y0, h_s_cla16_and1308_y0);
  and_gate and_gate_h_s_cla16_and1309_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1309_y0);
  and_gate and_gate_h_s_cla16_and1310_y0(h_s_cla16_and1309_y0, h_s_cla16_and1308_y0, h_s_cla16_and1310_y0);
  and_gate and_gate_h_s_cla16_and1311_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1311_y0);
  and_gate and_gate_h_s_cla16_and1312_y0(h_s_cla16_and1311_y0, h_s_cla16_and1310_y0, h_s_cla16_and1312_y0);
  and_gate and_gate_h_s_cla16_and1313_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1313_y0);
  and_gate and_gate_h_s_cla16_and1314_y0(h_s_cla16_and1313_y0, h_s_cla16_and1312_y0, h_s_cla16_and1314_y0);
  and_gate and_gate_h_s_cla16_and1315_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1315_y0);
  and_gate and_gate_h_s_cla16_and1316_y0(h_s_cla16_and1315_y0, h_s_cla16_and1314_y0, h_s_cla16_and1316_y0);
  and_gate and_gate_h_s_cla16_and1317_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1317_y0);
  and_gate and_gate_h_s_cla16_and1318_y0(h_s_cla16_and1317_y0, h_s_cla16_and1316_y0, h_s_cla16_and1318_y0);
  and_gate and_gate_h_s_cla16_and1319_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1319_y0);
  and_gate and_gate_h_s_cla16_and1320_y0(h_s_cla16_and1319_y0, h_s_cla16_and1318_y0, h_s_cla16_and1320_y0);
  and_gate and_gate_h_s_cla16_and1321_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1321_y0);
  and_gate and_gate_h_s_cla16_and1322_y0(h_s_cla16_and1321_y0, h_s_cla16_and1320_y0, h_s_cla16_and1322_y0);
  and_gate and_gate_h_s_cla16_and1323_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1323_y0);
  and_gate and_gate_h_s_cla16_and1324_y0(h_s_cla16_and1323_y0, h_s_cla16_and1322_y0, h_s_cla16_and1324_y0);
  and_gate and_gate_h_s_cla16_and1325_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic1_y1, h_s_cla16_and1325_y0);
  and_gate and_gate_h_s_cla16_and1326_y0(h_s_cla16_and1325_y0, h_s_cla16_and1324_y0, h_s_cla16_and1326_y0);
  and_gate and_gate_h_s_cla16_and1327_y0(h_s_cla16_pg_logic3_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1327_y0);
  and_gate and_gate_h_s_cla16_and1328_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1328_y0);
  and_gate and_gate_h_s_cla16_and1329_y0(h_s_cla16_and1328_y0, h_s_cla16_and1327_y0, h_s_cla16_and1329_y0);
  and_gate and_gate_h_s_cla16_and1330_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1330_y0);
  and_gate and_gate_h_s_cla16_and1331_y0(h_s_cla16_and1330_y0, h_s_cla16_and1329_y0, h_s_cla16_and1331_y0);
  and_gate and_gate_h_s_cla16_and1332_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1332_y0);
  and_gate and_gate_h_s_cla16_and1333_y0(h_s_cla16_and1332_y0, h_s_cla16_and1331_y0, h_s_cla16_and1333_y0);
  and_gate and_gate_h_s_cla16_and1334_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1334_y0);
  and_gate and_gate_h_s_cla16_and1335_y0(h_s_cla16_and1334_y0, h_s_cla16_and1333_y0, h_s_cla16_and1335_y0);
  and_gate and_gate_h_s_cla16_and1336_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1336_y0);
  and_gate and_gate_h_s_cla16_and1337_y0(h_s_cla16_and1336_y0, h_s_cla16_and1335_y0, h_s_cla16_and1337_y0);
  and_gate and_gate_h_s_cla16_and1338_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1338_y0);
  and_gate and_gate_h_s_cla16_and1339_y0(h_s_cla16_and1338_y0, h_s_cla16_and1337_y0, h_s_cla16_and1339_y0);
  and_gate and_gate_h_s_cla16_and1340_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1340_y0);
  and_gate and_gate_h_s_cla16_and1341_y0(h_s_cla16_and1340_y0, h_s_cla16_and1339_y0, h_s_cla16_and1341_y0);
  and_gate and_gate_h_s_cla16_and1342_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1342_y0);
  and_gate and_gate_h_s_cla16_and1343_y0(h_s_cla16_and1342_y0, h_s_cla16_and1341_y0, h_s_cla16_and1343_y0);
  and_gate and_gate_h_s_cla16_and1344_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1344_y0);
  and_gate and_gate_h_s_cla16_and1345_y0(h_s_cla16_and1344_y0, h_s_cla16_and1343_y0, h_s_cla16_and1345_y0);
  and_gate and_gate_h_s_cla16_and1346_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1346_y0);
  and_gate and_gate_h_s_cla16_and1347_y0(h_s_cla16_and1346_y0, h_s_cla16_and1345_y0, h_s_cla16_and1347_y0);
  and_gate and_gate_h_s_cla16_and1348_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1348_y0);
  and_gate and_gate_h_s_cla16_and1349_y0(h_s_cla16_and1348_y0, h_s_cla16_and1347_y0, h_s_cla16_and1349_y0);
  and_gate and_gate_h_s_cla16_and1350_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic2_y1, h_s_cla16_and1350_y0);
  and_gate and_gate_h_s_cla16_and1351_y0(h_s_cla16_and1350_y0, h_s_cla16_and1349_y0, h_s_cla16_and1351_y0);
  and_gate and_gate_h_s_cla16_and1352_y0(h_s_cla16_pg_logic4_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1352_y0);
  and_gate and_gate_h_s_cla16_and1353_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1353_y0);
  and_gate and_gate_h_s_cla16_and1354_y0(h_s_cla16_and1353_y0, h_s_cla16_and1352_y0, h_s_cla16_and1354_y0);
  and_gate and_gate_h_s_cla16_and1355_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1355_y0);
  and_gate and_gate_h_s_cla16_and1356_y0(h_s_cla16_and1355_y0, h_s_cla16_and1354_y0, h_s_cla16_and1356_y0);
  and_gate and_gate_h_s_cla16_and1357_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1357_y0);
  and_gate and_gate_h_s_cla16_and1358_y0(h_s_cla16_and1357_y0, h_s_cla16_and1356_y0, h_s_cla16_and1358_y0);
  and_gate and_gate_h_s_cla16_and1359_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1359_y0);
  and_gate and_gate_h_s_cla16_and1360_y0(h_s_cla16_and1359_y0, h_s_cla16_and1358_y0, h_s_cla16_and1360_y0);
  and_gate and_gate_h_s_cla16_and1361_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1361_y0);
  and_gate and_gate_h_s_cla16_and1362_y0(h_s_cla16_and1361_y0, h_s_cla16_and1360_y0, h_s_cla16_and1362_y0);
  and_gate and_gate_h_s_cla16_and1363_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1363_y0);
  and_gate and_gate_h_s_cla16_and1364_y0(h_s_cla16_and1363_y0, h_s_cla16_and1362_y0, h_s_cla16_and1364_y0);
  and_gate and_gate_h_s_cla16_and1365_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1365_y0);
  and_gate and_gate_h_s_cla16_and1366_y0(h_s_cla16_and1365_y0, h_s_cla16_and1364_y0, h_s_cla16_and1366_y0);
  and_gate and_gate_h_s_cla16_and1367_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1367_y0);
  and_gate and_gate_h_s_cla16_and1368_y0(h_s_cla16_and1367_y0, h_s_cla16_and1366_y0, h_s_cla16_and1368_y0);
  and_gate and_gate_h_s_cla16_and1369_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1369_y0);
  and_gate and_gate_h_s_cla16_and1370_y0(h_s_cla16_and1369_y0, h_s_cla16_and1368_y0, h_s_cla16_and1370_y0);
  and_gate and_gate_h_s_cla16_and1371_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1371_y0);
  and_gate and_gate_h_s_cla16_and1372_y0(h_s_cla16_and1371_y0, h_s_cla16_and1370_y0, h_s_cla16_and1372_y0);
  and_gate and_gate_h_s_cla16_and1373_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic3_y1, h_s_cla16_and1373_y0);
  and_gate and_gate_h_s_cla16_and1374_y0(h_s_cla16_and1373_y0, h_s_cla16_and1372_y0, h_s_cla16_and1374_y0);
  and_gate and_gate_h_s_cla16_and1375_y0(h_s_cla16_pg_logic5_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1375_y0);
  and_gate and_gate_h_s_cla16_and1376_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1376_y0);
  and_gate and_gate_h_s_cla16_and1377_y0(h_s_cla16_and1376_y0, h_s_cla16_and1375_y0, h_s_cla16_and1377_y0);
  and_gate and_gate_h_s_cla16_and1378_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1378_y0);
  and_gate and_gate_h_s_cla16_and1379_y0(h_s_cla16_and1378_y0, h_s_cla16_and1377_y0, h_s_cla16_and1379_y0);
  and_gate and_gate_h_s_cla16_and1380_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1380_y0);
  and_gate and_gate_h_s_cla16_and1381_y0(h_s_cla16_and1380_y0, h_s_cla16_and1379_y0, h_s_cla16_and1381_y0);
  and_gate and_gate_h_s_cla16_and1382_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1382_y0);
  and_gate and_gate_h_s_cla16_and1383_y0(h_s_cla16_and1382_y0, h_s_cla16_and1381_y0, h_s_cla16_and1383_y0);
  and_gate and_gate_h_s_cla16_and1384_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1384_y0);
  and_gate and_gate_h_s_cla16_and1385_y0(h_s_cla16_and1384_y0, h_s_cla16_and1383_y0, h_s_cla16_and1385_y0);
  and_gate and_gate_h_s_cla16_and1386_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1386_y0);
  and_gate and_gate_h_s_cla16_and1387_y0(h_s_cla16_and1386_y0, h_s_cla16_and1385_y0, h_s_cla16_and1387_y0);
  and_gate and_gate_h_s_cla16_and1388_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1388_y0);
  and_gate and_gate_h_s_cla16_and1389_y0(h_s_cla16_and1388_y0, h_s_cla16_and1387_y0, h_s_cla16_and1389_y0);
  and_gate and_gate_h_s_cla16_and1390_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1390_y0);
  and_gate and_gate_h_s_cla16_and1391_y0(h_s_cla16_and1390_y0, h_s_cla16_and1389_y0, h_s_cla16_and1391_y0);
  and_gate and_gate_h_s_cla16_and1392_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1392_y0);
  and_gate and_gate_h_s_cla16_and1393_y0(h_s_cla16_and1392_y0, h_s_cla16_and1391_y0, h_s_cla16_and1393_y0);
  and_gate and_gate_h_s_cla16_and1394_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic4_y1, h_s_cla16_and1394_y0);
  and_gate and_gate_h_s_cla16_and1395_y0(h_s_cla16_and1394_y0, h_s_cla16_and1393_y0, h_s_cla16_and1395_y0);
  and_gate and_gate_h_s_cla16_and1396_y0(h_s_cla16_pg_logic6_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1396_y0);
  and_gate and_gate_h_s_cla16_and1397_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1397_y0);
  and_gate and_gate_h_s_cla16_and1398_y0(h_s_cla16_and1397_y0, h_s_cla16_and1396_y0, h_s_cla16_and1398_y0);
  and_gate and_gate_h_s_cla16_and1399_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1399_y0);
  and_gate and_gate_h_s_cla16_and1400_y0(h_s_cla16_and1399_y0, h_s_cla16_and1398_y0, h_s_cla16_and1400_y0);
  and_gate and_gate_h_s_cla16_and1401_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1401_y0);
  and_gate and_gate_h_s_cla16_and1402_y0(h_s_cla16_and1401_y0, h_s_cla16_and1400_y0, h_s_cla16_and1402_y0);
  and_gate and_gate_h_s_cla16_and1403_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1403_y0);
  and_gate and_gate_h_s_cla16_and1404_y0(h_s_cla16_and1403_y0, h_s_cla16_and1402_y0, h_s_cla16_and1404_y0);
  and_gate and_gate_h_s_cla16_and1405_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1405_y0);
  and_gate and_gate_h_s_cla16_and1406_y0(h_s_cla16_and1405_y0, h_s_cla16_and1404_y0, h_s_cla16_and1406_y0);
  and_gate and_gate_h_s_cla16_and1407_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1407_y0);
  and_gate and_gate_h_s_cla16_and1408_y0(h_s_cla16_and1407_y0, h_s_cla16_and1406_y0, h_s_cla16_and1408_y0);
  and_gate and_gate_h_s_cla16_and1409_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1409_y0);
  and_gate and_gate_h_s_cla16_and1410_y0(h_s_cla16_and1409_y0, h_s_cla16_and1408_y0, h_s_cla16_and1410_y0);
  and_gate and_gate_h_s_cla16_and1411_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1411_y0);
  and_gate and_gate_h_s_cla16_and1412_y0(h_s_cla16_and1411_y0, h_s_cla16_and1410_y0, h_s_cla16_and1412_y0);
  and_gate and_gate_h_s_cla16_and1413_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic5_y1, h_s_cla16_and1413_y0);
  and_gate and_gate_h_s_cla16_and1414_y0(h_s_cla16_and1413_y0, h_s_cla16_and1412_y0, h_s_cla16_and1414_y0);
  and_gate and_gate_h_s_cla16_and1415_y0(h_s_cla16_pg_logic7_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1415_y0);
  and_gate and_gate_h_s_cla16_and1416_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1416_y0);
  and_gate and_gate_h_s_cla16_and1417_y0(h_s_cla16_and1416_y0, h_s_cla16_and1415_y0, h_s_cla16_and1417_y0);
  and_gate and_gate_h_s_cla16_and1418_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1418_y0);
  and_gate and_gate_h_s_cla16_and1419_y0(h_s_cla16_and1418_y0, h_s_cla16_and1417_y0, h_s_cla16_and1419_y0);
  and_gate and_gate_h_s_cla16_and1420_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1420_y0);
  and_gate and_gate_h_s_cla16_and1421_y0(h_s_cla16_and1420_y0, h_s_cla16_and1419_y0, h_s_cla16_and1421_y0);
  and_gate and_gate_h_s_cla16_and1422_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1422_y0);
  and_gate and_gate_h_s_cla16_and1423_y0(h_s_cla16_and1422_y0, h_s_cla16_and1421_y0, h_s_cla16_and1423_y0);
  and_gate and_gate_h_s_cla16_and1424_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1424_y0);
  and_gate and_gate_h_s_cla16_and1425_y0(h_s_cla16_and1424_y0, h_s_cla16_and1423_y0, h_s_cla16_and1425_y0);
  and_gate and_gate_h_s_cla16_and1426_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1426_y0);
  and_gate and_gate_h_s_cla16_and1427_y0(h_s_cla16_and1426_y0, h_s_cla16_and1425_y0, h_s_cla16_and1427_y0);
  and_gate and_gate_h_s_cla16_and1428_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1428_y0);
  and_gate and_gate_h_s_cla16_and1429_y0(h_s_cla16_and1428_y0, h_s_cla16_and1427_y0, h_s_cla16_and1429_y0);
  and_gate and_gate_h_s_cla16_and1430_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic6_y1, h_s_cla16_and1430_y0);
  and_gate and_gate_h_s_cla16_and1431_y0(h_s_cla16_and1430_y0, h_s_cla16_and1429_y0, h_s_cla16_and1431_y0);
  and_gate and_gate_h_s_cla16_and1432_y0(h_s_cla16_pg_logic8_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1432_y0);
  and_gate and_gate_h_s_cla16_and1433_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1433_y0);
  and_gate and_gate_h_s_cla16_and1434_y0(h_s_cla16_and1433_y0, h_s_cla16_and1432_y0, h_s_cla16_and1434_y0);
  and_gate and_gate_h_s_cla16_and1435_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1435_y0);
  and_gate and_gate_h_s_cla16_and1436_y0(h_s_cla16_and1435_y0, h_s_cla16_and1434_y0, h_s_cla16_and1436_y0);
  and_gate and_gate_h_s_cla16_and1437_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1437_y0);
  and_gate and_gate_h_s_cla16_and1438_y0(h_s_cla16_and1437_y0, h_s_cla16_and1436_y0, h_s_cla16_and1438_y0);
  and_gate and_gate_h_s_cla16_and1439_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1439_y0);
  and_gate and_gate_h_s_cla16_and1440_y0(h_s_cla16_and1439_y0, h_s_cla16_and1438_y0, h_s_cla16_and1440_y0);
  and_gate and_gate_h_s_cla16_and1441_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1441_y0);
  and_gate and_gate_h_s_cla16_and1442_y0(h_s_cla16_and1441_y0, h_s_cla16_and1440_y0, h_s_cla16_and1442_y0);
  and_gate and_gate_h_s_cla16_and1443_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1443_y0);
  and_gate and_gate_h_s_cla16_and1444_y0(h_s_cla16_and1443_y0, h_s_cla16_and1442_y0, h_s_cla16_and1444_y0);
  and_gate and_gate_h_s_cla16_and1445_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic7_y1, h_s_cla16_and1445_y0);
  and_gate and_gate_h_s_cla16_and1446_y0(h_s_cla16_and1445_y0, h_s_cla16_and1444_y0, h_s_cla16_and1446_y0);
  and_gate and_gate_h_s_cla16_and1447_y0(h_s_cla16_pg_logic9_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1447_y0);
  and_gate and_gate_h_s_cla16_and1448_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1448_y0);
  and_gate and_gate_h_s_cla16_and1449_y0(h_s_cla16_and1448_y0, h_s_cla16_and1447_y0, h_s_cla16_and1449_y0);
  and_gate and_gate_h_s_cla16_and1450_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1450_y0);
  and_gate and_gate_h_s_cla16_and1451_y0(h_s_cla16_and1450_y0, h_s_cla16_and1449_y0, h_s_cla16_and1451_y0);
  and_gate and_gate_h_s_cla16_and1452_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1452_y0);
  and_gate and_gate_h_s_cla16_and1453_y0(h_s_cla16_and1452_y0, h_s_cla16_and1451_y0, h_s_cla16_and1453_y0);
  and_gate and_gate_h_s_cla16_and1454_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1454_y0);
  and_gate and_gate_h_s_cla16_and1455_y0(h_s_cla16_and1454_y0, h_s_cla16_and1453_y0, h_s_cla16_and1455_y0);
  and_gate and_gate_h_s_cla16_and1456_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1456_y0);
  and_gate and_gate_h_s_cla16_and1457_y0(h_s_cla16_and1456_y0, h_s_cla16_and1455_y0, h_s_cla16_and1457_y0);
  and_gate and_gate_h_s_cla16_and1458_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic8_y1, h_s_cla16_and1458_y0);
  and_gate and_gate_h_s_cla16_and1459_y0(h_s_cla16_and1458_y0, h_s_cla16_and1457_y0, h_s_cla16_and1459_y0);
  and_gate and_gate_h_s_cla16_and1460_y0(h_s_cla16_pg_logic10_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1460_y0);
  and_gate and_gate_h_s_cla16_and1461_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1461_y0);
  and_gate and_gate_h_s_cla16_and1462_y0(h_s_cla16_and1461_y0, h_s_cla16_and1460_y0, h_s_cla16_and1462_y0);
  and_gate and_gate_h_s_cla16_and1463_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1463_y0);
  and_gate and_gate_h_s_cla16_and1464_y0(h_s_cla16_and1463_y0, h_s_cla16_and1462_y0, h_s_cla16_and1464_y0);
  and_gate and_gate_h_s_cla16_and1465_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1465_y0);
  and_gate and_gate_h_s_cla16_and1466_y0(h_s_cla16_and1465_y0, h_s_cla16_and1464_y0, h_s_cla16_and1466_y0);
  and_gate and_gate_h_s_cla16_and1467_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1467_y0);
  and_gate and_gate_h_s_cla16_and1468_y0(h_s_cla16_and1467_y0, h_s_cla16_and1466_y0, h_s_cla16_and1468_y0);
  and_gate and_gate_h_s_cla16_and1469_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic9_y1, h_s_cla16_and1469_y0);
  and_gate and_gate_h_s_cla16_and1470_y0(h_s_cla16_and1469_y0, h_s_cla16_and1468_y0, h_s_cla16_and1470_y0);
  and_gate and_gate_h_s_cla16_and1471_y0(h_s_cla16_pg_logic11_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1471_y0);
  and_gate and_gate_h_s_cla16_and1472_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1472_y0);
  and_gate and_gate_h_s_cla16_and1473_y0(h_s_cla16_and1472_y0, h_s_cla16_and1471_y0, h_s_cla16_and1473_y0);
  and_gate and_gate_h_s_cla16_and1474_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1474_y0);
  and_gate and_gate_h_s_cla16_and1475_y0(h_s_cla16_and1474_y0, h_s_cla16_and1473_y0, h_s_cla16_and1475_y0);
  and_gate and_gate_h_s_cla16_and1476_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1476_y0);
  and_gate and_gate_h_s_cla16_and1477_y0(h_s_cla16_and1476_y0, h_s_cla16_and1475_y0, h_s_cla16_and1477_y0);
  and_gate and_gate_h_s_cla16_and1478_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic10_y1, h_s_cla16_and1478_y0);
  and_gate and_gate_h_s_cla16_and1479_y0(h_s_cla16_and1478_y0, h_s_cla16_and1477_y0, h_s_cla16_and1479_y0);
  and_gate and_gate_h_s_cla16_and1480_y0(h_s_cla16_pg_logic12_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1480_y0);
  and_gate and_gate_h_s_cla16_and1481_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1481_y0);
  and_gate and_gate_h_s_cla16_and1482_y0(h_s_cla16_and1481_y0, h_s_cla16_and1480_y0, h_s_cla16_and1482_y0);
  and_gate and_gate_h_s_cla16_and1483_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1483_y0);
  and_gate and_gate_h_s_cla16_and1484_y0(h_s_cla16_and1483_y0, h_s_cla16_and1482_y0, h_s_cla16_and1484_y0);
  and_gate and_gate_h_s_cla16_and1485_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic11_y1, h_s_cla16_and1485_y0);
  and_gate and_gate_h_s_cla16_and1486_y0(h_s_cla16_and1485_y0, h_s_cla16_and1484_y0, h_s_cla16_and1486_y0);
  and_gate and_gate_h_s_cla16_and1487_y0(h_s_cla16_pg_logic13_y0, h_s_cla16_pg_logic12_y1, h_s_cla16_and1487_y0);
  and_gate and_gate_h_s_cla16_and1488_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic12_y1, h_s_cla16_and1488_y0);
  and_gate and_gate_h_s_cla16_and1489_y0(h_s_cla16_and1488_y0, h_s_cla16_and1487_y0, h_s_cla16_and1489_y0);
  and_gate and_gate_h_s_cla16_and1490_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic12_y1, h_s_cla16_and1490_y0);
  and_gate and_gate_h_s_cla16_and1491_y0(h_s_cla16_and1490_y0, h_s_cla16_and1489_y0, h_s_cla16_and1491_y0);
  and_gate and_gate_h_s_cla16_and1492_y0(h_s_cla16_pg_logic14_y0, h_s_cla16_pg_logic13_y1, h_s_cla16_and1492_y0);
  and_gate and_gate_h_s_cla16_and1493_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic13_y1, h_s_cla16_and1493_y0);
  and_gate and_gate_h_s_cla16_and1494_y0(h_s_cla16_and1493_y0, h_s_cla16_and1492_y0, h_s_cla16_and1494_y0);
  and_gate and_gate_h_s_cla16_and1495_y0(h_s_cla16_pg_logic15_y0, h_s_cla16_pg_logic14_y1, h_s_cla16_and1495_y0);
  or_gate or_gate_h_s_cla16_or120_y0(h_s_cla16_and1495_y0, h_s_cla16_and1270_y0, h_s_cla16_or120_y0);
  or_gate or_gate_h_s_cla16_or121_y0(h_s_cla16_or120_y0, h_s_cla16_and1299_y0, h_s_cla16_or121_y0);
  or_gate or_gate_h_s_cla16_or122_y0(h_s_cla16_or121_y0, h_s_cla16_and1326_y0, h_s_cla16_or122_y0);
  or_gate or_gate_h_s_cla16_or123_y0(h_s_cla16_or122_y0, h_s_cla16_and1351_y0, h_s_cla16_or123_y0);
  or_gate or_gate_h_s_cla16_or124_y0(h_s_cla16_or123_y0, h_s_cla16_and1374_y0, h_s_cla16_or124_y0);
  or_gate or_gate_h_s_cla16_or125_y0(h_s_cla16_or124_y0, h_s_cla16_and1395_y0, h_s_cla16_or125_y0);
  or_gate or_gate_h_s_cla16_or126_y0(h_s_cla16_or125_y0, h_s_cla16_and1414_y0, h_s_cla16_or126_y0);
  or_gate or_gate_h_s_cla16_or127_y0(h_s_cla16_or126_y0, h_s_cla16_and1431_y0, h_s_cla16_or127_y0);
  or_gate or_gate_h_s_cla16_or128_y0(h_s_cla16_or127_y0, h_s_cla16_and1446_y0, h_s_cla16_or128_y0);
  or_gate or_gate_h_s_cla16_or129_y0(h_s_cla16_or128_y0, h_s_cla16_and1459_y0, h_s_cla16_or129_y0);
  or_gate or_gate_h_s_cla16_or130_y0(h_s_cla16_or129_y0, h_s_cla16_and1470_y0, h_s_cla16_or130_y0);
  or_gate or_gate_h_s_cla16_or131_y0(h_s_cla16_or130_y0, h_s_cla16_and1479_y0, h_s_cla16_or131_y0);
  or_gate or_gate_h_s_cla16_or132_y0(h_s_cla16_or131_y0, h_s_cla16_and1486_y0, h_s_cla16_or132_y0);
  or_gate or_gate_h_s_cla16_or133_y0(h_s_cla16_or132_y0, h_s_cla16_and1491_y0, h_s_cla16_or133_y0);
  or_gate or_gate_h_s_cla16_or134_y0(h_s_cla16_or133_y0, h_s_cla16_and1494_y0, h_s_cla16_or134_y0);
  or_gate or_gate_h_s_cla16_or135_y0(h_s_cla16_pg_logic15_y1, h_s_cla16_or134_y0, h_s_cla16_or135_y0);
  xor_gate xor_gate_h_s_cla16_xor16_y0(a_15, b_15, h_s_cla16_xor16_y0);
  xor_gate xor_gate_h_s_cla16_xor17_y0(h_s_cla16_xor16_y0, h_s_cla16_or135_y0, h_s_cla16_xor17_y0);

  assign out[0] = h_s_cla16_xor0_y0;
  assign out[1] = h_s_cla16_xor1_y0;
  assign out[2] = h_s_cla16_xor2_y0;
  assign out[3] = h_s_cla16_xor3_y0;
  assign out[4] = h_s_cla16_xor4_y0;
  assign out[5] = h_s_cla16_xor5_y0;
  assign out[6] = h_s_cla16_xor6_y0;
  assign out[7] = h_s_cla16_xor7_y0;
  assign out[8] = h_s_cla16_xor8_y0;
  assign out[9] = h_s_cla16_xor9_y0;
  assign out[10] = h_s_cla16_xor10_y0;
  assign out[11] = h_s_cla16_xor11_y0;
  assign out[12] = h_s_cla16_xor12_y0;
  assign out[13] = h_s_cla16_xor13_y0;
  assign out[14] = h_s_cla16_xor14_y0;
  assign out[15] = h_s_cla16_xor15_y0;
  assign out[16] = h_s_cla16_xor17_y0;
endmodule