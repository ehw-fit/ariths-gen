module s_CSAwallace_cla16(input [15:0] a, input [15:0] b, output [31:0] s_CSAwallace_cla16_out);
  wire s_CSAwallace_cla16_and_0_0;
  wire s_CSAwallace_cla16_and_1_0;
  wire s_CSAwallace_cla16_and_2_0;
  wire s_CSAwallace_cla16_and_3_0;
  wire s_CSAwallace_cla16_and_4_0;
  wire s_CSAwallace_cla16_and_5_0;
  wire s_CSAwallace_cla16_and_6_0;
  wire s_CSAwallace_cla16_and_7_0;
  wire s_CSAwallace_cla16_and_8_0;
  wire s_CSAwallace_cla16_and_9_0;
  wire s_CSAwallace_cla16_and_10_0;
  wire s_CSAwallace_cla16_and_11_0;
  wire s_CSAwallace_cla16_and_12_0;
  wire s_CSAwallace_cla16_and_13_0;
  wire s_CSAwallace_cla16_and_14_0;
  wire s_CSAwallace_cla16_nand_15_0;
  wire s_CSAwallace_cla16_and_0_1;
  wire s_CSAwallace_cla16_and_1_1;
  wire s_CSAwallace_cla16_and_2_1;
  wire s_CSAwallace_cla16_and_3_1;
  wire s_CSAwallace_cla16_and_4_1;
  wire s_CSAwallace_cla16_and_5_1;
  wire s_CSAwallace_cla16_and_6_1;
  wire s_CSAwallace_cla16_and_7_1;
  wire s_CSAwallace_cla16_and_8_1;
  wire s_CSAwallace_cla16_and_9_1;
  wire s_CSAwallace_cla16_and_10_1;
  wire s_CSAwallace_cla16_and_11_1;
  wire s_CSAwallace_cla16_and_12_1;
  wire s_CSAwallace_cla16_and_13_1;
  wire s_CSAwallace_cla16_and_14_1;
  wire s_CSAwallace_cla16_nand_15_1;
  wire s_CSAwallace_cla16_and_0_2;
  wire s_CSAwallace_cla16_and_1_2;
  wire s_CSAwallace_cla16_and_2_2;
  wire s_CSAwallace_cla16_and_3_2;
  wire s_CSAwallace_cla16_and_4_2;
  wire s_CSAwallace_cla16_and_5_2;
  wire s_CSAwallace_cla16_and_6_2;
  wire s_CSAwallace_cla16_and_7_2;
  wire s_CSAwallace_cla16_and_8_2;
  wire s_CSAwallace_cla16_and_9_2;
  wire s_CSAwallace_cla16_and_10_2;
  wire s_CSAwallace_cla16_and_11_2;
  wire s_CSAwallace_cla16_and_12_2;
  wire s_CSAwallace_cla16_and_13_2;
  wire s_CSAwallace_cla16_and_14_2;
  wire s_CSAwallace_cla16_nand_15_2;
  wire s_CSAwallace_cla16_and_0_3;
  wire s_CSAwallace_cla16_and_1_3;
  wire s_CSAwallace_cla16_and_2_3;
  wire s_CSAwallace_cla16_and_3_3;
  wire s_CSAwallace_cla16_and_4_3;
  wire s_CSAwallace_cla16_and_5_3;
  wire s_CSAwallace_cla16_and_6_3;
  wire s_CSAwallace_cla16_and_7_3;
  wire s_CSAwallace_cla16_and_8_3;
  wire s_CSAwallace_cla16_and_9_3;
  wire s_CSAwallace_cla16_and_10_3;
  wire s_CSAwallace_cla16_and_11_3;
  wire s_CSAwallace_cla16_and_12_3;
  wire s_CSAwallace_cla16_and_13_3;
  wire s_CSAwallace_cla16_and_14_3;
  wire s_CSAwallace_cla16_nand_15_3;
  wire s_CSAwallace_cla16_and_0_4;
  wire s_CSAwallace_cla16_and_1_4;
  wire s_CSAwallace_cla16_and_2_4;
  wire s_CSAwallace_cla16_and_3_4;
  wire s_CSAwallace_cla16_and_4_4;
  wire s_CSAwallace_cla16_and_5_4;
  wire s_CSAwallace_cla16_and_6_4;
  wire s_CSAwallace_cla16_and_7_4;
  wire s_CSAwallace_cla16_and_8_4;
  wire s_CSAwallace_cla16_and_9_4;
  wire s_CSAwallace_cla16_and_10_4;
  wire s_CSAwallace_cla16_and_11_4;
  wire s_CSAwallace_cla16_and_12_4;
  wire s_CSAwallace_cla16_and_13_4;
  wire s_CSAwallace_cla16_and_14_4;
  wire s_CSAwallace_cla16_nand_15_4;
  wire s_CSAwallace_cla16_and_0_5;
  wire s_CSAwallace_cla16_and_1_5;
  wire s_CSAwallace_cla16_and_2_5;
  wire s_CSAwallace_cla16_and_3_5;
  wire s_CSAwallace_cla16_and_4_5;
  wire s_CSAwallace_cla16_and_5_5;
  wire s_CSAwallace_cla16_and_6_5;
  wire s_CSAwallace_cla16_and_7_5;
  wire s_CSAwallace_cla16_and_8_5;
  wire s_CSAwallace_cla16_and_9_5;
  wire s_CSAwallace_cla16_and_10_5;
  wire s_CSAwallace_cla16_and_11_5;
  wire s_CSAwallace_cla16_and_12_5;
  wire s_CSAwallace_cla16_and_13_5;
  wire s_CSAwallace_cla16_and_14_5;
  wire s_CSAwallace_cla16_nand_15_5;
  wire s_CSAwallace_cla16_and_0_6;
  wire s_CSAwallace_cla16_and_1_6;
  wire s_CSAwallace_cla16_and_2_6;
  wire s_CSAwallace_cla16_and_3_6;
  wire s_CSAwallace_cla16_and_4_6;
  wire s_CSAwallace_cla16_and_5_6;
  wire s_CSAwallace_cla16_and_6_6;
  wire s_CSAwallace_cla16_and_7_6;
  wire s_CSAwallace_cla16_and_8_6;
  wire s_CSAwallace_cla16_and_9_6;
  wire s_CSAwallace_cla16_and_10_6;
  wire s_CSAwallace_cla16_and_11_6;
  wire s_CSAwallace_cla16_and_12_6;
  wire s_CSAwallace_cla16_and_13_6;
  wire s_CSAwallace_cla16_and_14_6;
  wire s_CSAwallace_cla16_nand_15_6;
  wire s_CSAwallace_cla16_and_0_7;
  wire s_CSAwallace_cla16_and_1_7;
  wire s_CSAwallace_cla16_and_2_7;
  wire s_CSAwallace_cla16_and_3_7;
  wire s_CSAwallace_cla16_and_4_7;
  wire s_CSAwallace_cla16_and_5_7;
  wire s_CSAwallace_cla16_and_6_7;
  wire s_CSAwallace_cla16_and_7_7;
  wire s_CSAwallace_cla16_and_8_7;
  wire s_CSAwallace_cla16_and_9_7;
  wire s_CSAwallace_cla16_and_10_7;
  wire s_CSAwallace_cla16_and_11_7;
  wire s_CSAwallace_cla16_and_12_7;
  wire s_CSAwallace_cla16_and_13_7;
  wire s_CSAwallace_cla16_and_14_7;
  wire s_CSAwallace_cla16_nand_15_7;
  wire s_CSAwallace_cla16_and_0_8;
  wire s_CSAwallace_cla16_and_1_8;
  wire s_CSAwallace_cla16_and_2_8;
  wire s_CSAwallace_cla16_and_3_8;
  wire s_CSAwallace_cla16_and_4_8;
  wire s_CSAwallace_cla16_and_5_8;
  wire s_CSAwallace_cla16_and_6_8;
  wire s_CSAwallace_cla16_and_7_8;
  wire s_CSAwallace_cla16_and_8_8;
  wire s_CSAwallace_cla16_and_9_8;
  wire s_CSAwallace_cla16_and_10_8;
  wire s_CSAwallace_cla16_and_11_8;
  wire s_CSAwallace_cla16_and_12_8;
  wire s_CSAwallace_cla16_and_13_8;
  wire s_CSAwallace_cla16_and_14_8;
  wire s_CSAwallace_cla16_nand_15_8;
  wire s_CSAwallace_cla16_and_0_9;
  wire s_CSAwallace_cla16_and_1_9;
  wire s_CSAwallace_cla16_and_2_9;
  wire s_CSAwallace_cla16_and_3_9;
  wire s_CSAwallace_cla16_and_4_9;
  wire s_CSAwallace_cla16_and_5_9;
  wire s_CSAwallace_cla16_and_6_9;
  wire s_CSAwallace_cla16_and_7_9;
  wire s_CSAwallace_cla16_and_8_9;
  wire s_CSAwallace_cla16_and_9_9;
  wire s_CSAwallace_cla16_and_10_9;
  wire s_CSAwallace_cla16_and_11_9;
  wire s_CSAwallace_cla16_and_12_9;
  wire s_CSAwallace_cla16_and_13_9;
  wire s_CSAwallace_cla16_and_14_9;
  wire s_CSAwallace_cla16_nand_15_9;
  wire s_CSAwallace_cla16_and_0_10;
  wire s_CSAwallace_cla16_and_1_10;
  wire s_CSAwallace_cla16_and_2_10;
  wire s_CSAwallace_cla16_and_3_10;
  wire s_CSAwallace_cla16_and_4_10;
  wire s_CSAwallace_cla16_and_5_10;
  wire s_CSAwallace_cla16_and_6_10;
  wire s_CSAwallace_cla16_and_7_10;
  wire s_CSAwallace_cla16_and_8_10;
  wire s_CSAwallace_cla16_and_9_10;
  wire s_CSAwallace_cla16_and_10_10;
  wire s_CSAwallace_cla16_and_11_10;
  wire s_CSAwallace_cla16_and_12_10;
  wire s_CSAwallace_cla16_and_13_10;
  wire s_CSAwallace_cla16_and_14_10;
  wire s_CSAwallace_cla16_nand_15_10;
  wire s_CSAwallace_cla16_and_0_11;
  wire s_CSAwallace_cla16_and_1_11;
  wire s_CSAwallace_cla16_and_2_11;
  wire s_CSAwallace_cla16_and_3_11;
  wire s_CSAwallace_cla16_and_4_11;
  wire s_CSAwallace_cla16_and_5_11;
  wire s_CSAwallace_cla16_and_6_11;
  wire s_CSAwallace_cla16_and_7_11;
  wire s_CSAwallace_cla16_and_8_11;
  wire s_CSAwallace_cla16_and_9_11;
  wire s_CSAwallace_cla16_and_10_11;
  wire s_CSAwallace_cla16_and_11_11;
  wire s_CSAwallace_cla16_and_12_11;
  wire s_CSAwallace_cla16_and_13_11;
  wire s_CSAwallace_cla16_and_14_11;
  wire s_CSAwallace_cla16_nand_15_11;
  wire s_CSAwallace_cla16_and_0_12;
  wire s_CSAwallace_cla16_and_1_12;
  wire s_CSAwallace_cla16_and_2_12;
  wire s_CSAwallace_cla16_and_3_12;
  wire s_CSAwallace_cla16_and_4_12;
  wire s_CSAwallace_cla16_and_5_12;
  wire s_CSAwallace_cla16_and_6_12;
  wire s_CSAwallace_cla16_and_7_12;
  wire s_CSAwallace_cla16_and_8_12;
  wire s_CSAwallace_cla16_and_9_12;
  wire s_CSAwallace_cla16_and_10_12;
  wire s_CSAwallace_cla16_and_11_12;
  wire s_CSAwallace_cla16_and_12_12;
  wire s_CSAwallace_cla16_and_13_12;
  wire s_CSAwallace_cla16_and_14_12;
  wire s_CSAwallace_cla16_nand_15_12;
  wire s_CSAwallace_cla16_and_0_13;
  wire s_CSAwallace_cla16_and_1_13;
  wire s_CSAwallace_cla16_and_2_13;
  wire s_CSAwallace_cla16_and_3_13;
  wire s_CSAwallace_cla16_and_4_13;
  wire s_CSAwallace_cla16_and_5_13;
  wire s_CSAwallace_cla16_and_6_13;
  wire s_CSAwallace_cla16_and_7_13;
  wire s_CSAwallace_cla16_and_8_13;
  wire s_CSAwallace_cla16_and_9_13;
  wire s_CSAwallace_cla16_and_10_13;
  wire s_CSAwallace_cla16_and_11_13;
  wire s_CSAwallace_cla16_and_12_13;
  wire s_CSAwallace_cla16_and_13_13;
  wire s_CSAwallace_cla16_and_14_13;
  wire s_CSAwallace_cla16_nand_15_13;
  wire s_CSAwallace_cla16_and_0_14;
  wire s_CSAwallace_cla16_and_1_14;
  wire s_CSAwallace_cla16_and_2_14;
  wire s_CSAwallace_cla16_and_3_14;
  wire s_CSAwallace_cla16_and_4_14;
  wire s_CSAwallace_cla16_and_5_14;
  wire s_CSAwallace_cla16_and_6_14;
  wire s_CSAwallace_cla16_and_7_14;
  wire s_CSAwallace_cla16_and_8_14;
  wire s_CSAwallace_cla16_and_9_14;
  wire s_CSAwallace_cla16_and_10_14;
  wire s_CSAwallace_cla16_and_11_14;
  wire s_CSAwallace_cla16_and_12_14;
  wire s_CSAwallace_cla16_and_13_14;
  wire s_CSAwallace_cla16_and_14_14;
  wire s_CSAwallace_cla16_nand_15_14;
  wire s_CSAwallace_cla16_nand_0_15;
  wire s_CSAwallace_cla16_nand_1_15;
  wire s_CSAwallace_cla16_nand_2_15;
  wire s_CSAwallace_cla16_nand_3_15;
  wire s_CSAwallace_cla16_nand_4_15;
  wire s_CSAwallace_cla16_nand_5_15;
  wire s_CSAwallace_cla16_nand_6_15;
  wire s_CSAwallace_cla16_nand_7_15;
  wire s_CSAwallace_cla16_nand_8_15;
  wire s_CSAwallace_cla16_nand_9_15;
  wire s_CSAwallace_cla16_nand_10_15;
  wire s_CSAwallace_cla16_nand_11_15;
  wire s_CSAwallace_cla16_nand_12_15;
  wire s_CSAwallace_cla16_nand_13_15;
  wire s_CSAwallace_cla16_nand_14_15;
  wire s_CSAwallace_cla16_and_15_15;
  wire s_CSAwallace_cla16_csa0_csa_component_fa1_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa1_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa2_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa2_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa2_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa2_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa2_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa3_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa3_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa3_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa3_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa3_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa4_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa4_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa4_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa4_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa4_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa5_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa5_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa5_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa5_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa5_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa6_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa6_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa6_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa6_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa6_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa7_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa7_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa7_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa8_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa8_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa8_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa9_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa9_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa9_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa10_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa10_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa10_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa0_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa0_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa4_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa4_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa5_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa5_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa5_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa5_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa5_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa6_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa6_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa6_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa6_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa6_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa7_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa7_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa7_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa8_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa8_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa8_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa9_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa9_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa9_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa10_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa10_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa10_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa1_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa1_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa8_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa8_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa8_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa9_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa9_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa9_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa10_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa10_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa10_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa2_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa2_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa22_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa23_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa24_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa24_and0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa24_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa24_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa24_or0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa25_xor0;
  wire s_CSAwallace_cla16_csa3_csa_component_fa25_xor1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa25_and1;
  wire s_CSAwallace_cla16_csa3_csa_component_fa25_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa22_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa23_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa24_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa24_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa24_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa24_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa24_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa25_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa25_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa25_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa25_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa25_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa26_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa26_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa26_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa26_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa26_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa27_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa27_and0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa27_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa27_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa27_or0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa28_xor0;
  wire s_CSAwallace_cla16_csa4_csa_component_fa28_xor1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa28_and1;
  wire s_CSAwallace_cla16_csa4_csa_component_fa28_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa2_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa2_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa3_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa3_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa3_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa3_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa3_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa4_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa4_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa4_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa4_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa4_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa5_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa5_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa5_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa5_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa5_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa6_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa6_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa6_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa6_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa6_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa7_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa7_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa7_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa8_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa8_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa8_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa9_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa9_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa9_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa10_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa10_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa10_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa5_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa5_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa6_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa6_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa8_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa8_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa8_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa9_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa9_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa9_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa10_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa10_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa10_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa6_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa6_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa22_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa23_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa24_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa24_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa24_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa24_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa24_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa25_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa25_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa25_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa25_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa25_or0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa26_xor0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa26_and0;
  wire s_CSAwallace_cla16_csa7_csa_component_fa26_xor1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa26_and1;
  wire s_CSAwallace_cla16_csa7_csa_component_fa26_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa3_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa3_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa4_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa4_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa5_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa5_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa5_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa5_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa5_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa6_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa6_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa6_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa6_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa6_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa7_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa7_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa7_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa8_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa8_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa8_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa9_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa9_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa9_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa10_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa10_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa10_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa8_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa8_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa22_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa23_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa24_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa24_and0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa24_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa24_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa24_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa25_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa25_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa25_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa25_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa26_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa26_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa26_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa26_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa27_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa27_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa27_and1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa27_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa28_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa28_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa28_or0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa29_xor0;
  wire s_CSAwallace_cla16_csa9_csa_component_fa29_xor1;
  wire s_CSAwallace_cla16_csa9_csa_component_fa29_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa4_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa4_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa5_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa5_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa6_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa6_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa7_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa7_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa7_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa8_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa8_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa8_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa9_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa9_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa9_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa10_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa10_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa10_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa10_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa10_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa22_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa23_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa24_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa24_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa24_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa24_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa24_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa25_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa25_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa25_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa25_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa25_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa26_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa26_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa26_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa26_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa26_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa27_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa27_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa27_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa27_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa27_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa28_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa28_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa28_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa28_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa28_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa29_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa29_and0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa29_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa29_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa29_or0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa30_xor0;
  wire s_CSAwallace_cla16_csa11_csa_component_fa30_xor1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa30_and1;
  wire s_CSAwallace_cla16_csa11_csa_component_fa30_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa5_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa5_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa6_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa6_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa10_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa10_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa10_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa11_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa11_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa11_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa12_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa12_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa12_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa13_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa13_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa13_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa14_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa14_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa14_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa22_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa23_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa24_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa24_and0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa24_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa24_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa24_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa25_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa25_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa25_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa25_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa26_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa26_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa26_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa26_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa27_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa27_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa27_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa27_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa28_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa28_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa28_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa28_or0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa29_xor0;
  wire s_CSAwallace_cla16_csa12_csa_component_fa29_xor1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa29_and1;
  wire s_CSAwallace_cla16_csa12_csa_component_fa29_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa6_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa6_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa7_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa7_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa8_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa8_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa9_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa9_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa10_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa10_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa11_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa11_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa12_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa12_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa13_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa13_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa14_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa14_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa15_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa15_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa15_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa15_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa15_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa16_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa16_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa16_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa16_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa16_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa17_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa17_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa17_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa17_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa17_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa18_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa18_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa18_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa18_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa18_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa19_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa19_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa19_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa19_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa19_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa20_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa20_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa20_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa20_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa20_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa21_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa21_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa21_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa21_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa21_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa22_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa22_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa22_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa22_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa22_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa23_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa23_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa23_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa23_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa23_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa24_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa24_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa24_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa24_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa24_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa25_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa25_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa25_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa25_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa25_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa26_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa26_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa26_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa26_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa26_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa27_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa27_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa27_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa27_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa27_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa28_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa28_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa28_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa28_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa28_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa29_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa29_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa29_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa29_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa29_or0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa30_xor0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa30_and0;
  wire s_CSAwallace_cla16_csa13_csa_component_fa30_xor1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa30_and1;
  wire s_CSAwallace_cla16_csa13_csa_component_fa30_or0;
  wire s_CSAwallace_cla16_u_cla32_and0;
  wire s_CSAwallace_cla16_u_cla32_and1;
  wire s_CSAwallace_cla16_u_cla32_and2;
  wire s_CSAwallace_cla16_u_cla32_and3;
  wire s_CSAwallace_cla16_u_cla32_pg_logic7_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic7_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic7_xor0;
  wire s_CSAwallace_cla16_u_cla32_and4;
  wire s_CSAwallace_cla16_u_cla32_and5;
  wire s_CSAwallace_cla16_u_cla32_pg_logic8_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic8_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic8_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor8;
  wire s_CSAwallace_cla16_u_cla32_and6;
  wire s_CSAwallace_cla16_u_cla32_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic9_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic9_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic9_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor9;
  wire s_CSAwallace_cla16_u_cla32_and7;
  wire s_CSAwallace_cla16_u_cla32_and8;
  wire s_CSAwallace_cla16_u_cla32_and9;
  wire s_CSAwallace_cla16_u_cla32_or1;
  wire s_CSAwallace_cla16_u_cla32_or2;
  wire s_CSAwallace_cla16_u_cla32_pg_logic10_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic10_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic10_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor10;
  wire s_CSAwallace_cla16_u_cla32_and10;
  wire s_CSAwallace_cla16_u_cla32_and11;
  wire s_CSAwallace_cla16_u_cla32_and12;
  wire s_CSAwallace_cla16_u_cla32_and13;
  wire s_CSAwallace_cla16_u_cla32_and14;
  wire s_CSAwallace_cla16_u_cla32_and15;
  wire s_CSAwallace_cla16_u_cla32_or3;
  wire s_CSAwallace_cla16_u_cla32_or4;
  wire s_CSAwallace_cla16_u_cla32_or5;
  wire s_CSAwallace_cla16_u_cla32_pg_logic11_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic11_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic11_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor11;
  wire s_CSAwallace_cla16_u_cla32_and16;
  wire s_CSAwallace_cla16_u_cla32_and17;
  wire s_CSAwallace_cla16_u_cla32_and18;
  wire s_CSAwallace_cla16_u_cla32_and19;
  wire s_CSAwallace_cla16_u_cla32_and20;
  wire s_CSAwallace_cla16_u_cla32_and21;
  wire s_CSAwallace_cla16_u_cla32_and22;
  wire s_CSAwallace_cla16_u_cla32_and23;
  wire s_CSAwallace_cla16_u_cla32_and24;
  wire s_CSAwallace_cla16_u_cla32_and25;
  wire s_CSAwallace_cla16_u_cla32_or6;
  wire s_CSAwallace_cla16_u_cla32_or7;
  wire s_CSAwallace_cla16_u_cla32_or8;
  wire s_CSAwallace_cla16_u_cla32_or9;
  wire s_CSAwallace_cla16_u_cla32_pg_logic12_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic12_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic12_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor12;
  wire s_CSAwallace_cla16_u_cla32_and26;
  wire s_CSAwallace_cla16_u_cla32_or10;
  wire s_CSAwallace_cla16_u_cla32_pg_logic13_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic13_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic13_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor13;
  wire s_CSAwallace_cla16_u_cla32_and27;
  wire s_CSAwallace_cla16_u_cla32_and28;
  wire s_CSAwallace_cla16_u_cla32_and29;
  wire s_CSAwallace_cla16_u_cla32_or11;
  wire s_CSAwallace_cla16_u_cla32_or12;
  wire s_CSAwallace_cla16_u_cla32_pg_logic14_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic14_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic14_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor14;
  wire s_CSAwallace_cla16_u_cla32_and30;
  wire s_CSAwallace_cla16_u_cla32_and31;
  wire s_CSAwallace_cla16_u_cla32_and32;
  wire s_CSAwallace_cla16_u_cla32_and33;
  wire s_CSAwallace_cla16_u_cla32_and34;
  wire s_CSAwallace_cla16_u_cla32_and35;
  wire s_CSAwallace_cla16_u_cla32_or13;
  wire s_CSAwallace_cla16_u_cla32_or14;
  wire s_CSAwallace_cla16_u_cla32_or15;
  wire s_CSAwallace_cla16_u_cla32_pg_logic15_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic15_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic15_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor15;
  wire s_CSAwallace_cla16_u_cla32_and36;
  wire s_CSAwallace_cla16_u_cla32_and37;
  wire s_CSAwallace_cla16_u_cla32_and38;
  wire s_CSAwallace_cla16_u_cla32_and39;
  wire s_CSAwallace_cla16_u_cla32_and40;
  wire s_CSAwallace_cla16_u_cla32_and41;
  wire s_CSAwallace_cla16_u_cla32_and42;
  wire s_CSAwallace_cla16_u_cla32_and43;
  wire s_CSAwallace_cla16_u_cla32_and44;
  wire s_CSAwallace_cla16_u_cla32_and45;
  wire s_CSAwallace_cla16_u_cla32_or16;
  wire s_CSAwallace_cla16_u_cla32_or17;
  wire s_CSAwallace_cla16_u_cla32_or18;
  wire s_CSAwallace_cla16_u_cla32_or19;
  wire s_CSAwallace_cla16_u_cla32_pg_logic16_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic16_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic16_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor16;
  wire s_CSAwallace_cla16_u_cla32_and46;
  wire s_CSAwallace_cla16_u_cla32_or20;
  wire s_CSAwallace_cla16_u_cla32_pg_logic17_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic17_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic17_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor17;
  wire s_CSAwallace_cla16_u_cla32_and47;
  wire s_CSAwallace_cla16_u_cla32_and48;
  wire s_CSAwallace_cla16_u_cla32_and49;
  wire s_CSAwallace_cla16_u_cla32_or21;
  wire s_CSAwallace_cla16_u_cla32_or22;
  wire s_CSAwallace_cla16_u_cla32_pg_logic18_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic18_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic18_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor18;
  wire s_CSAwallace_cla16_u_cla32_and50;
  wire s_CSAwallace_cla16_u_cla32_and51;
  wire s_CSAwallace_cla16_u_cla32_and52;
  wire s_CSAwallace_cla16_u_cla32_and53;
  wire s_CSAwallace_cla16_u_cla32_and54;
  wire s_CSAwallace_cla16_u_cla32_and55;
  wire s_CSAwallace_cla16_u_cla32_or23;
  wire s_CSAwallace_cla16_u_cla32_or24;
  wire s_CSAwallace_cla16_u_cla32_or25;
  wire s_CSAwallace_cla16_u_cla32_pg_logic19_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic19_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic19_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor19;
  wire s_CSAwallace_cla16_u_cla32_and56;
  wire s_CSAwallace_cla16_u_cla32_and57;
  wire s_CSAwallace_cla16_u_cla32_and58;
  wire s_CSAwallace_cla16_u_cla32_and59;
  wire s_CSAwallace_cla16_u_cla32_and60;
  wire s_CSAwallace_cla16_u_cla32_and61;
  wire s_CSAwallace_cla16_u_cla32_and62;
  wire s_CSAwallace_cla16_u_cla32_and63;
  wire s_CSAwallace_cla16_u_cla32_and64;
  wire s_CSAwallace_cla16_u_cla32_and65;
  wire s_CSAwallace_cla16_u_cla32_or26;
  wire s_CSAwallace_cla16_u_cla32_or27;
  wire s_CSAwallace_cla16_u_cla32_or28;
  wire s_CSAwallace_cla16_u_cla32_or29;
  wire s_CSAwallace_cla16_u_cla32_pg_logic20_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic20_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic20_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor20;
  wire s_CSAwallace_cla16_u_cla32_and66;
  wire s_CSAwallace_cla16_u_cla32_or30;
  wire s_CSAwallace_cla16_u_cla32_pg_logic21_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic21_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic21_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor21;
  wire s_CSAwallace_cla16_u_cla32_and67;
  wire s_CSAwallace_cla16_u_cla32_and68;
  wire s_CSAwallace_cla16_u_cla32_and69;
  wire s_CSAwallace_cla16_u_cla32_or31;
  wire s_CSAwallace_cla16_u_cla32_or32;
  wire s_CSAwallace_cla16_u_cla32_pg_logic22_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic22_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic22_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor22;
  wire s_CSAwallace_cla16_u_cla32_and70;
  wire s_CSAwallace_cla16_u_cla32_and71;
  wire s_CSAwallace_cla16_u_cla32_and72;
  wire s_CSAwallace_cla16_u_cla32_and73;
  wire s_CSAwallace_cla16_u_cla32_and74;
  wire s_CSAwallace_cla16_u_cla32_and75;
  wire s_CSAwallace_cla16_u_cla32_or33;
  wire s_CSAwallace_cla16_u_cla32_or34;
  wire s_CSAwallace_cla16_u_cla32_or35;
  wire s_CSAwallace_cla16_u_cla32_pg_logic23_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic23_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic23_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor23;
  wire s_CSAwallace_cla16_u_cla32_and76;
  wire s_CSAwallace_cla16_u_cla32_and77;
  wire s_CSAwallace_cla16_u_cla32_and78;
  wire s_CSAwallace_cla16_u_cla32_and79;
  wire s_CSAwallace_cla16_u_cla32_and80;
  wire s_CSAwallace_cla16_u_cla32_and81;
  wire s_CSAwallace_cla16_u_cla32_and82;
  wire s_CSAwallace_cla16_u_cla32_and83;
  wire s_CSAwallace_cla16_u_cla32_and84;
  wire s_CSAwallace_cla16_u_cla32_and85;
  wire s_CSAwallace_cla16_u_cla32_or36;
  wire s_CSAwallace_cla16_u_cla32_or37;
  wire s_CSAwallace_cla16_u_cla32_or38;
  wire s_CSAwallace_cla16_u_cla32_or39;
  wire s_CSAwallace_cla16_u_cla32_pg_logic24_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic24_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic24_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor24;
  wire s_CSAwallace_cla16_u_cla32_and86;
  wire s_CSAwallace_cla16_u_cla32_or40;
  wire s_CSAwallace_cla16_u_cla32_pg_logic25_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic25_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic25_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor25;
  wire s_CSAwallace_cla16_u_cla32_and87;
  wire s_CSAwallace_cla16_u_cla32_and88;
  wire s_CSAwallace_cla16_u_cla32_and89;
  wire s_CSAwallace_cla16_u_cla32_or41;
  wire s_CSAwallace_cla16_u_cla32_or42;
  wire s_CSAwallace_cla16_u_cla32_pg_logic26_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic26_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic26_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor26;
  wire s_CSAwallace_cla16_u_cla32_and90;
  wire s_CSAwallace_cla16_u_cla32_and91;
  wire s_CSAwallace_cla16_u_cla32_and92;
  wire s_CSAwallace_cla16_u_cla32_and93;
  wire s_CSAwallace_cla16_u_cla32_and94;
  wire s_CSAwallace_cla16_u_cla32_and95;
  wire s_CSAwallace_cla16_u_cla32_or43;
  wire s_CSAwallace_cla16_u_cla32_or44;
  wire s_CSAwallace_cla16_u_cla32_or45;
  wire s_CSAwallace_cla16_u_cla32_pg_logic27_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic27_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic27_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor27;
  wire s_CSAwallace_cla16_u_cla32_and96;
  wire s_CSAwallace_cla16_u_cla32_and97;
  wire s_CSAwallace_cla16_u_cla32_and98;
  wire s_CSAwallace_cla16_u_cla32_and99;
  wire s_CSAwallace_cla16_u_cla32_and100;
  wire s_CSAwallace_cla16_u_cla32_and101;
  wire s_CSAwallace_cla16_u_cla32_and102;
  wire s_CSAwallace_cla16_u_cla32_and103;
  wire s_CSAwallace_cla16_u_cla32_and104;
  wire s_CSAwallace_cla16_u_cla32_and105;
  wire s_CSAwallace_cla16_u_cla32_or46;
  wire s_CSAwallace_cla16_u_cla32_or47;
  wire s_CSAwallace_cla16_u_cla32_or48;
  wire s_CSAwallace_cla16_u_cla32_or49;
  wire s_CSAwallace_cla16_u_cla32_pg_logic28_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic28_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic28_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor28;
  wire s_CSAwallace_cla16_u_cla32_and106;
  wire s_CSAwallace_cla16_u_cla32_or50;
  wire s_CSAwallace_cla16_u_cla32_pg_logic29_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic29_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic29_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor29;
  wire s_CSAwallace_cla16_u_cla32_and107;
  wire s_CSAwallace_cla16_u_cla32_and108;
  wire s_CSAwallace_cla16_u_cla32_and109;
  wire s_CSAwallace_cla16_u_cla32_or51;
  wire s_CSAwallace_cla16_u_cla32_or52;
  wire s_CSAwallace_cla16_u_cla32_pg_logic30_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic30_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic30_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor30;
  wire s_CSAwallace_cla16_u_cla32_and110;
  wire s_CSAwallace_cla16_u_cla32_and111;
  wire s_CSAwallace_cla16_u_cla32_and112;
  wire s_CSAwallace_cla16_u_cla32_and113;
  wire s_CSAwallace_cla16_u_cla32_and114;
  wire s_CSAwallace_cla16_u_cla32_and115;
  wire s_CSAwallace_cla16_u_cla32_or53;
  wire s_CSAwallace_cla16_u_cla32_or54;
  wire s_CSAwallace_cla16_u_cla32_or55;
  wire s_CSAwallace_cla16_u_cla32_pg_logic31_or0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic31_and0;
  wire s_CSAwallace_cla16_u_cla32_pg_logic31_xor0;
  wire s_CSAwallace_cla16_u_cla32_xor31;
  wire s_CSAwallace_cla16_u_cla32_and116;
  wire s_CSAwallace_cla16_u_cla32_and117;
  wire s_CSAwallace_cla16_u_cla32_and118;
  wire s_CSAwallace_cla16_u_cla32_and119;
  wire s_CSAwallace_cla16_u_cla32_and120;
  wire s_CSAwallace_cla16_u_cla32_and121;
  wire s_CSAwallace_cla16_u_cla32_and122;
  wire s_CSAwallace_cla16_u_cla32_and123;
  wire s_CSAwallace_cla16_u_cla32_and124;
  wire s_CSAwallace_cla16_u_cla32_and125;
  wire s_CSAwallace_cla16_u_cla32_or56;
  wire s_CSAwallace_cla16_u_cla32_or57;
  wire s_CSAwallace_cla16_u_cla32_or58;
  wire s_CSAwallace_cla16_u_cla32_or59;
  wire s_CSAwallace_cla16_xor0;

  assign s_CSAwallace_cla16_and_0_0 = a[0] & b[0];
  assign s_CSAwallace_cla16_and_1_0 = a[1] & b[0];
  assign s_CSAwallace_cla16_and_2_0 = a[2] & b[0];
  assign s_CSAwallace_cla16_and_3_0 = a[3] & b[0];
  assign s_CSAwallace_cla16_and_4_0 = a[4] & b[0];
  assign s_CSAwallace_cla16_and_5_0 = a[5] & b[0];
  assign s_CSAwallace_cla16_and_6_0 = a[6] & b[0];
  assign s_CSAwallace_cla16_and_7_0 = a[7] & b[0];
  assign s_CSAwallace_cla16_and_8_0 = a[8] & b[0];
  assign s_CSAwallace_cla16_and_9_0 = a[9] & b[0];
  assign s_CSAwallace_cla16_and_10_0 = a[10] & b[0];
  assign s_CSAwallace_cla16_and_11_0 = a[11] & b[0];
  assign s_CSAwallace_cla16_and_12_0 = a[12] & b[0];
  assign s_CSAwallace_cla16_and_13_0 = a[13] & b[0];
  assign s_CSAwallace_cla16_and_14_0 = a[14] & b[0];
  assign s_CSAwallace_cla16_nand_15_0 = ~(a[15] & b[0]);
  assign s_CSAwallace_cla16_and_0_1 = a[0] & b[1];
  assign s_CSAwallace_cla16_and_1_1 = a[1] & b[1];
  assign s_CSAwallace_cla16_and_2_1 = a[2] & b[1];
  assign s_CSAwallace_cla16_and_3_1 = a[3] & b[1];
  assign s_CSAwallace_cla16_and_4_1 = a[4] & b[1];
  assign s_CSAwallace_cla16_and_5_1 = a[5] & b[1];
  assign s_CSAwallace_cla16_and_6_1 = a[6] & b[1];
  assign s_CSAwallace_cla16_and_7_1 = a[7] & b[1];
  assign s_CSAwallace_cla16_and_8_1 = a[8] & b[1];
  assign s_CSAwallace_cla16_and_9_1 = a[9] & b[1];
  assign s_CSAwallace_cla16_and_10_1 = a[10] & b[1];
  assign s_CSAwallace_cla16_and_11_1 = a[11] & b[1];
  assign s_CSAwallace_cla16_and_12_1 = a[12] & b[1];
  assign s_CSAwallace_cla16_and_13_1 = a[13] & b[1];
  assign s_CSAwallace_cla16_and_14_1 = a[14] & b[1];
  assign s_CSAwallace_cla16_nand_15_1 = ~(a[15] & b[1]);
  assign s_CSAwallace_cla16_and_0_2 = a[0] & b[2];
  assign s_CSAwallace_cla16_and_1_2 = a[1] & b[2];
  assign s_CSAwallace_cla16_and_2_2 = a[2] & b[2];
  assign s_CSAwallace_cla16_and_3_2 = a[3] & b[2];
  assign s_CSAwallace_cla16_and_4_2 = a[4] & b[2];
  assign s_CSAwallace_cla16_and_5_2 = a[5] & b[2];
  assign s_CSAwallace_cla16_and_6_2 = a[6] & b[2];
  assign s_CSAwallace_cla16_and_7_2 = a[7] & b[2];
  assign s_CSAwallace_cla16_and_8_2 = a[8] & b[2];
  assign s_CSAwallace_cla16_and_9_2 = a[9] & b[2];
  assign s_CSAwallace_cla16_and_10_2 = a[10] & b[2];
  assign s_CSAwallace_cla16_and_11_2 = a[11] & b[2];
  assign s_CSAwallace_cla16_and_12_2 = a[12] & b[2];
  assign s_CSAwallace_cla16_and_13_2 = a[13] & b[2];
  assign s_CSAwallace_cla16_and_14_2 = a[14] & b[2];
  assign s_CSAwallace_cla16_nand_15_2 = ~(a[15] & b[2]);
  assign s_CSAwallace_cla16_and_0_3 = a[0] & b[3];
  assign s_CSAwallace_cla16_and_1_3 = a[1] & b[3];
  assign s_CSAwallace_cla16_and_2_3 = a[2] & b[3];
  assign s_CSAwallace_cla16_and_3_3 = a[3] & b[3];
  assign s_CSAwallace_cla16_and_4_3 = a[4] & b[3];
  assign s_CSAwallace_cla16_and_5_3 = a[5] & b[3];
  assign s_CSAwallace_cla16_and_6_3 = a[6] & b[3];
  assign s_CSAwallace_cla16_and_7_3 = a[7] & b[3];
  assign s_CSAwallace_cla16_and_8_3 = a[8] & b[3];
  assign s_CSAwallace_cla16_and_9_3 = a[9] & b[3];
  assign s_CSAwallace_cla16_and_10_3 = a[10] & b[3];
  assign s_CSAwallace_cla16_and_11_3 = a[11] & b[3];
  assign s_CSAwallace_cla16_and_12_3 = a[12] & b[3];
  assign s_CSAwallace_cla16_and_13_3 = a[13] & b[3];
  assign s_CSAwallace_cla16_and_14_3 = a[14] & b[3];
  assign s_CSAwallace_cla16_nand_15_3 = ~(a[15] & b[3]);
  assign s_CSAwallace_cla16_and_0_4 = a[0] & b[4];
  assign s_CSAwallace_cla16_and_1_4 = a[1] & b[4];
  assign s_CSAwallace_cla16_and_2_4 = a[2] & b[4];
  assign s_CSAwallace_cla16_and_3_4 = a[3] & b[4];
  assign s_CSAwallace_cla16_and_4_4 = a[4] & b[4];
  assign s_CSAwallace_cla16_and_5_4 = a[5] & b[4];
  assign s_CSAwallace_cla16_and_6_4 = a[6] & b[4];
  assign s_CSAwallace_cla16_and_7_4 = a[7] & b[4];
  assign s_CSAwallace_cla16_and_8_4 = a[8] & b[4];
  assign s_CSAwallace_cla16_and_9_4 = a[9] & b[4];
  assign s_CSAwallace_cla16_and_10_4 = a[10] & b[4];
  assign s_CSAwallace_cla16_and_11_4 = a[11] & b[4];
  assign s_CSAwallace_cla16_and_12_4 = a[12] & b[4];
  assign s_CSAwallace_cla16_and_13_4 = a[13] & b[4];
  assign s_CSAwallace_cla16_and_14_4 = a[14] & b[4];
  assign s_CSAwallace_cla16_nand_15_4 = ~(a[15] & b[4]);
  assign s_CSAwallace_cla16_and_0_5 = a[0] & b[5];
  assign s_CSAwallace_cla16_and_1_5 = a[1] & b[5];
  assign s_CSAwallace_cla16_and_2_5 = a[2] & b[5];
  assign s_CSAwallace_cla16_and_3_5 = a[3] & b[5];
  assign s_CSAwallace_cla16_and_4_5 = a[4] & b[5];
  assign s_CSAwallace_cla16_and_5_5 = a[5] & b[5];
  assign s_CSAwallace_cla16_and_6_5 = a[6] & b[5];
  assign s_CSAwallace_cla16_and_7_5 = a[7] & b[5];
  assign s_CSAwallace_cla16_and_8_5 = a[8] & b[5];
  assign s_CSAwallace_cla16_and_9_5 = a[9] & b[5];
  assign s_CSAwallace_cla16_and_10_5 = a[10] & b[5];
  assign s_CSAwallace_cla16_and_11_5 = a[11] & b[5];
  assign s_CSAwallace_cla16_and_12_5 = a[12] & b[5];
  assign s_CSAwallace_cla16_and_13_5 = a[13] & b[5];
  assign s_CSAwallace_cla16_and_14_5 = a[14] & b[5];
  assign s_CSAwallace_cla16_nand_15_5 = ~(a[15] & b[5]);
  assign s_CSAwallace_cla16_and_0_6 = a[0] & b[6];
  assign s_CSAwallace_cla16_and_1_6 = a[1] & b[6];
  assign s_CSAwallace_cla16_and_2_6 = a[2] & b[6];
  assign s_CSAwallace_cla16_and_3_6 = a[3] & b[6];
  assign s_CSAwallace_cla16_and_4_6 = a[4] & b[6];
  assign s_CSAwallace_cla16_and_5_6 = a[5] & b[6];
  assign s_CSAwallace_cla16_and_6_6 = a[6] & b[6];
  assign s_CSAwallace_cla16_and_7_6 = a[7] & b[6];
  assign s_CSAwallace_cla16_and_8_6 = a[8] & b[6];
  assign s_CSAwallace_cla16_and_9_6 = a[9] & b[6];
  assign s_CSAwallace_cla16_and_10_6 = a[10] & b[6];
  assign s_CSAwallace_cla16_and_11_6 = a[11] & b[6];
  assign s_CSAwallace_cla16_and_12_6 = a[12] & b[6];
  assign s_CSAwallace_cla16_and_13_6 = a[13] & b[6];
  assign s_CSAwallace_cla16_and_14_6 = a[14] & b[6];
  assign s_CSAwallace_cla16_nand_15_6 = ~(a[15] & b[6]);
  assign s_CSAwallace_cla16_and_0_7 = a[0] & b[7];
  assign s_CSAwallace_cla16_and_1_7 = a[1] & b[7];
  assign s_CSAwallace_cla16_and_2_7 = a[2] & b[7];
  assign s_CSAwallace_cla16_and_3_7 = a[3] & b[7];
  assign s_CSAwallace_cla16_and_4_7 = a[4] & b[7];
  assign s_CSAwallace_cla16_and_5_7 = a[5] & b[7];
  assign s_CSAwallace_cla16_and_6_7 = a[6] & b[7];
  assign s_CSAwallace_cla16_and_7_7 = a[7] & b[7];
  assign s_CSAwallace_cla16_and_8_7 = a[8] & b[7];
  assign s_CSAwallace_cla16_and_9_7 = a[9] & b[7];
  assign s_CSAwallace_cla16_and_10_7 = a[10] & b[7];
  assign s_CSAwallace_cla16_and_11_7 = a[11] & b[7];
  assign s_CSAwallace_cla16_and_12_7 = a[12] & b[7];
  assign s_CSAwallace_cla16_and_13_7 = a[13] & b[7];
  assign s_CSAwallace_cla16_and_14_7 = a[14] & b[7];
  assign s_CSAwallace_cla16_nand_15_7 = ~(a[15] & b[7]);
  assign s_CSAwallace_cla16_and_0_8 = a[0] & b[8];
  assign s_CSAwallace_cla16_and_1_8 = a[1] & b[8];
  assign s_CSAwallace_cla16_and_2_8 = a[2] & b[8];
  assign s_CSAwallace_cla16_and_3_8 = a[3] & b[8];
  assign s_CSAwallace_cla16_and_4_8 = a[4] & b[8];
  assign s_CSAwallace_cla16_and_5_8 = a[5] & b[8];
  assign s_CSAwallace_cla16_and_6_8 = a[6] & b[8];
  assign s_CSAwallace_cla16_and_7_8 = a[7] & b[8];
  assign s_CSAwallace_cla16_and_8_8 = a[8] & b[8];
  assign s_CSAwallace_cla16_and_9_8 = a[9] & b[8];
  assign s_CSAwallace_cla16_and_10_8 = a[10] & b[8];
  assign s_CSAwallace_cla16_and_11_8 = a[11] & b[8];
  assign s_CSAwallace_cla16_and_12_8 = a[12] & b[8];
  assign s_CSAwallace_cla16_and_13_8 = a[13] & b[8];
  assign s_CSAwallace_cla16_and_14_8 = a[14] & b[8];
  assign s_CSAwallace_cla16_nand_15_8 = ~(a[15] & b[8]);
  assign s_CSAwallace_cla16_and_0_9 = a[0] & b[9];
  assign s_CSAwallace_cla16_and_1_9 = a[1] & b[9];
  assign s_CSAwallace_cla16_and_2_9 = a[2] & b[9];
  assign s_CSAwallace_cla16_and_3_9 = a[3] & b[9];
  assign s_CSAwallace_cla16_and_4_9 = a[4] & b[9];
  assign s_CSAwallace_cla16_and_5_9 = a[5] & b[9];
  assign s_CSAwallace_cla16_and_6_9 = a[6] & b[9];
  assign s_CSAwallace_cla16_and_7_9 = a[7] & b[9];
  assign s_CSAwallace_cla16_and_8_9 = a[8] & b[9];
  assign s_CSAwallace_cla16_and_9_9 = a[9] & b[9];
  assign s_CSAwallace_cla16_and_10_9 = a[10] & b[9];
  assign s_CSAwallace_cla16_and_11_9 = a[11] & b[9];
  assign s_CSAwallace_cla16_and_12_9 = a[12] & b[9];
  assign s_CSAwallace_cla16_and_13_9 = a[13] & b[9];
  assign s_CSAwallace_cla16_and_14_9 = a[14] & b[9];
  assign s_CSAwallace_cla16_nand_15_9 = ~(a[15] & b[9]);
  assign s_CSAwallace_cla16_and_0_10 = a[0] & b[10];
  assign s_CSAwallace_cla16_and_1_10 = a[1] & b[10];
  assign s_CSAwallace_cla16_and_2_10 = a[2] & b[10];
  assign s_CSAwallace_cla16_and_3_10 = a[3] & b[10];
  assign s_CSAwallace_cla16_and_4_10 = a[4] & b[10];
  assign s_CSAwallace_cla16_and_5_10 = a[5] & b[10];
  assign s_CSAwallace_cla16_and_6_10 = a[6] & b[10];
  assign s_CSAwallace_cla16_and_7_10 = a[7] & b[10];
  assign s_CSAwallace_cla16_and_8_10 = a[8] & b[10];
  assign s_CSAwallace_cla16_and_9_10 = a[9] & b[10];
  assign s_CSAwallace_cla16_and_10_10 = a[10] & b[10];
  assign s_CSAwallace_cla16_and_11_10 = a[11] & b[10];
  assign s_CSAwallace_cla16_and_12_10 = a[12] & b[10];
  assign s_CSAwallace_cla16_and_13_10 = a[13] & b[10];
  assign s_CSAwallace_cla16_and_14_10 = a[14] & b[10];
  assign s_CSAwallace_cla16_nand_15_10 = ~(a[15] & b[10]);
  assign s_CSAwallace_cla16_and_0_11 = a[0] & b[11];
  assign s_CSAwallace_cla16_and_1_11 = a[1] & b[11];
  assign s_CSAwallace_cla16_and_2_11 = a[2] & b[11];
  assign s_CSAwallace_cla16_and_3_11 = a[3] & b[11];
  assign s_CSAwallace_cla16_and_4_11 = a[4] & b[11];
  assign s_CSAwallace_cla16_and_5_11 = a[5] & b[11];
  assign s_CSAwallace_cla16_and_6_11 = a[6] & b[11];
  assign s_CSAwallace_cla16_and_7_11 = a[7] & b[11];
  assign s_CSAwallace_cla16_and_8_11 = a[8] & b[11];
  assign s_CSAwallace_cla16_and_9_11 = a[9] & b[11];
  assign s_CSAwallace_cla16_and_10_11 = a[10] & b[11];
  assign s_CSAwallace_cla16_and_11_11 = a[11] & b[11];
  assign s_CSAwallace_cla16_and_12_11 = a[12] & b[11];
  assign s_CSAwallace_cla16_and_13_11 = a[13] & b[11];
  assign s_CSAwallace_cla16_and_14_11 = a[14] & b[11];
  assign s_CSAwallace_cla16_nand_15_11 = ~(a[15] & b[11]);
  assign s_CSAwallace_cla16_and_0_12 = a[0] & b[12];
  assign s_CSAwallace_cla16_and_1_12 = a[1] & b[12];
  assign s_CSAwallace_cla16_and_2_12 = a[2] & b[12];
  assign s_CSAwallace_cla16_and_3_12 = a[3] & b[12];
  assign s_CSAwallace_cla16_and_4_12 = a[4] & b[12];
  assign s_CSAwallace_cla16_and_5_12 = a[5] & b[12];
  assign s_CSAwallace_cla16_and_6_12 = a[6] & b[12];
  assign s_CSAwallace_cla16_and_7_12 = a[7] & b[12];
  assign s_CSAwallace_cla16_and_8_12 = a[8] & b[12];
  assign s_CSAwallace_cla16_and_9_12 = a[9] & b[12];
  assign s_CSAwallace_cla16_and_10_12 = a[10] & b[12];
  assign s_CSAwallace_cla16_and_11_12 = a[11] & b[12];
  assign s_CSAwallace_cla16_and_12_12 = a[12] & b[12];
  assign s_CSAwallace_cla16_and_13_12 = a[13] & b[12];
  assign s_CSAwallace_cla16_and_14_12 = a[14] & b[12];
  assign s_CSAwallace_cla16_nand_15_12 = ~(a[15] & b[12]);
  assign s_CSAwallace_cla16_and_0_13 = a[0] & b[13];
  assign s_CSAwallace_cla16_and_1_13 = a[1] & b[13];
  assign s_CSAwallace_cla16_and_2_13 = a[2] & b[13];
  assign s_CSAwallace_cla16_and_3_13 = a[3] & b[13];
  assign s_CSAwallace_cla16_and_4_13 = a[4] & b[13];
  assign s_CSAwallace_cla16_and_5_13 = a[5] & b[13];
  assign s_CSAwallace_cla16_and_6_13 = a[6] & b[13];
  assign s_CSAwallace_cla16_and_7_13 = a[7] & b[13];
  assign s_CSAwallace_cla16_and_8_13 = a[8] & b[13];
  assign s_CSAwallace_cla16_and_9_13 = a[9] & b[13];
  assign s_CSAwallace_cla16_and_10_13 = a[10] & b[13];
  assign s_CSAwallace_cla16_and_11_13 = a[11] & b[13];
  assign s_CSAwallace_cla16_and_12_13 = a[12] & b[13];
  assign s_CSAwallace_cla16_and_13_13 = a[13] & b[13];
  assign s_CSAwallace_cla16_and_14_13 = a[14] & b[13];
  assign s_CSAwallace_cla16_nand_15_13 = ~(a[15] & b[13]);
  assign s_CSAwallace_cla16_and_0_14 = a[0] & b[14];
  assign s_CSAwallace_cla16_and_1_14 = a[1] & b[14];
  assign s_CSAwallace_cla16_and_2_14 = a[2] & b[14];
  assign s_CSAwallace_cla16_and_3_14 = a[3] & b[14];
  assign s_CSAwallace_cla16_and_4_14 = a[4] & b[14];
  assign s_CSAwallace_cla16_and_5_14 = a[5] & b[14];
  assign s_CSAwallace_cla16_and_6_14 = a[6] & b[14];
  assign s_CSAwallace_cla16_and_7_14 = a[7] & b[14];
  assign s_CSAwallace_cla16_and_8_14 = a[8] & b[14];
  assign s_CSAwallace_cla16_and_9_14 = a[9] & b[14];
  assign s_CSAwallace_cla16_and_10_14 = a[10] & b[14];
  assign s_CSAwallace_cla16_and_11_14 = a[11] & b[14];
  assign s_CSAwallace_cla16_and_12_14 = a[12] & b[14];
  assign s_CSAwallace_cla16_and_13_14 = a[13] & b[14];
  assign s_CSAwallace_cla16_and_14_14 = a[14] & b[14];
  assign s_CSAwallace_cla16_nand_15_14 = ~(a[15] & b[14]);
  assign s_CSAwallace_cla16_nand_0_15 = ~(a[0] & b[15]);
  assign s_CSAwallace_cla16_nand_1_15 = ~(a[1] & b[15]);
  assign s_CSAwallace_cla16_nand_2_15 = ~(a[2] & b[15]);
  assign s_CSAwallace_cla16_nand_3_15 = ~(a[3] & b[15]);
  assign s_CSAwallace_cla16_nand_4_15 = ~(a[4] & b[15]);
  assign s_CSAwallace_cla16_nand_5_15 = ~(a[5] & b[15]);
  assign s_CSAwallace_cla16_nand_6_15 = ~(a[6] & b[15]);
  assign s_CSAwallace_cla16_nand_7_15 = ~(a[7] & b[15]);
  assign s_CSAwallace_cla16_nand_8_15 = ~(a[8] & b[15]);
  assign s_CSAwallace_cla16_nand_9_15 = ~(a[9] & b[15]);
  assign s_CSAwallace_cla16_nand_10_15 = ~(a[10] & b[15]);
  assign s_CSAwallace_cla16_nand_11_15 = ~(a[11] & b[15]);
  assign s_CSAwallace_cla16_nand_12_15 = ~(a[12] & b[15]);
  assign s_CSAwallace_cla16_nand_13_15 = ~(a[13] & b[15]);
  assign s_CSAwallace_cla16_nand_14_15 = ~(a[14] & b[15]);
  assign s_CSAwallace_cla16_and_15_15 = a[15] & b[15];
  assign s_CSAwallace_cla16_csa0_csa_component_fa1_xor0 = s_CSAwallace_cla16_and_1_0 ^ s_CSAwallace_cla16_and_0_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa1_and0 = s_CSAwallace_cla16_and_1_0 & s_CSAwallace_cla16_and_0_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa2_xor0 = s_CSAwallace_cla16_and_2_0 ^ s_CSAwallace_cla16_and_1_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa2_and0 = s_CSAwallace_cla16_and_2_0 & s_CSAwallace_cla16_and_1_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa2_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa2_xor0 ^ s_CSAwallace_cla16_and_0_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa2_and1 = s_CSAwallace_cla16_csa0_csa_component_fa2_xor0 & s_CSAwallace_cla16_and_0_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa2_or0 = s_CSAwallace_cla16_csa0_csa_component_fa2_and0 | s_CSAwallace_cla16_csa0_csa_component_fa2_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa3_xor0 = s_CSAwallace_cla16_and_3_0 ^ s_CSAwallace_cla16_and_2_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa3_and0 = s_CSAwallace_cla16_and_3_0 & s_CSAwallace_cla16_and_2_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa3_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa3_xor0 ^ s_CSAwallace_cla16_and_1_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa3_and1 = s_CSAwallace_cla16_csa0_csa_component_fa3_xor0 & s_CSAwallace_cla16_and_1_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa3_or0 = s_CSAwallace_cla16_csa0_csa_component_fa3_and0 | s_CSAwallace_cla16_csa0_csa_component_fa3_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa4_xor0 = s_CSAwallace_cla16_and_4_0 ^ s_CSAwallace_cla16_and_3_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa4_and0 = s_CSAwallace_cla16_and_4_0 & s_CSAwallace_cla16_and_3_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa4_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa4_xor0 ^ s_CSAwallace_cla16_and_2_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa4_and1 = s_CSAwallace_cla16_csa0_csa_component_fa4_xor0 & s_CSAwallace_cla16_and_2_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa4_or0 = s_CSAwallace_cla16_csa0_csa_component_fa4_and0 | s_CSAwallace_cla16_csa0_csa_component_fa4_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa5_xor0 = s_CSAwallace_cla16_and_5_0 ^ s_CSAwallace_cla16_and_4_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa5_and0 = s_CSAwallace_cla16_and_5_0 & s_CSAwallace_cla16_and_4_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa5_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa5_xor0 ^ s_CSAwallace_cla16_and_3_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa5_and1 = s_CSAwallace_cla16_csa0_csa_component_fa5_xor0 & s_CSAwallace_cla16_and_3_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa5_or0 = s_CSAwallace_cla16_csa0_csa_component_fa5_and0 | s_CSAwallace_cla16_csa0_csa_component_fa5_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa6_xor0 = s_CSAwallace_cla16_and_6_0 ^ s_CSAwallace_cla16_and_5_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa6_and0 = s_CSAwallace_cla16_and_6_0 & s_CSAwallace_cla16_and_5_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa6_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa6_xor0 ^ s_CSAwallace_cla16_and_4_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa6_and1 = s_CSAwallace_cla16_csa0_csa_component_fa6_xor0 & s_CSAwallace_cla16_and_4_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa6_or0 = s_CSAwallace_cla16_csa0_csa_component_fa6_and0 | s_CSAwallace_cla16_csa0_csa_component_fa6_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa7_xor0 = s_CSAwallace_cla16_and_7_0 ^ s_CSAwallace_cla16_and_6_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa7_and0 = s_CSAwallace_cla16_and_7_0 & s_CSAwallace_cla16_and_6_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa7_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa7_xor0 ^ s_CSAwallace_cla16_and_5_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa7_and1 = s_CSAwallace_cla16_csa0_csa_component_fa7_xor0 & s_CSAwallace_cla16_and_5_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa7_or0 = s_CSAwallace_cla16_csa0_csa_component_fa7_and0 | s_CSAwallace_cla16_csa0_csa_component_fa7_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa8_xor0 = s_CSAwallace_cla16_and_8_0 ^ s_CSAwallace_cla16_and_7_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa8_and0 = s_CSAwallace_cla16_and_8_0 & s_CSAwallace_cla16_and_7_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa8_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_and_6_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa8_and1 = s_CSAwallace_cla16_csa0_csa_component_fa8_xor0 & s_CSAwallace_cla16_and_6_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa8_or0 = s_CSAwallace_cla16_csa0_csa_component_fa8_and0 | s_CSAwallace_cla16_csa0_csa_component_fa8_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa9_xor0 = s_CSAwallace_cla16_and_9_0 ^ s_CSAwallace_cla16_and_8_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa9_and0 = s_CSAwallace_cla16_and_9_0 & s_CSAwallace_cla16_and_8_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa9_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_and_7_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa9_and1 = s_CSAwallace_cla16_csa0_csa_component_fa9_xor0 & s_CSAwallace_cla16_and_7_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa9_or0 = s_CSAwallace_cla16_csa0_csa_component_fa9_and0 | s_CSAwallace_cla16_csa0_csa_component_fa9_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa10_xor0 = s_CSAwallace_cla16_and_10_0 ^ s_CSAwallace_cla16_and_9_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa10_and0 = s_CSAwallace_cla16_and_10_0 & s_CSAwallace_cla16_and_9_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa10_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_and_8_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa10_and1 = s_CSAwallace_cla16_csa0_csa_component_fa10_xor0 & s_CSAwallace_cla16_and_8_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa10_or0 = s_CSAwallace_cla16_csa0_csa_component_fa10_and0 | s_CSAwallace_cla16_csa0_csa_component_fa10_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa11_xor0 = s_CSAwallace_cla16_and_11_0 ^ s_CSAwallace_cla16_and_10_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa11_and0 = s_CSAwallace_cla16_and_11_0 & s_CSAwallace_cla16_and_10_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_and_9_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa11_and1 = s_CSAwallace_cla16_csa0_csa_component_fa11_xor0 & s_CSAwallace_cla16_and_9_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa11_or0 = s_CSAwallace_cla16_csa0_csa_component_fa11_and0 | s_CSAwallace_cla16_csa0_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa12_xor0 = s_CSAwallace_cla16_and_12_0 ^ s_CSAwallace_cla16_and_11_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa12_and0 = s_CSAwallace_cla16_and_12_0 & s_CSAwallace_cla16_and_11_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_and_10_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa12_and1 = s_CSAwallace_cla16_csa0_csa_component_fa12_xor0 & s_CSAwallace_cla16_and_10_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa12_or0 = s_CSAwallace_cla16_csa0_csa_component_fa12_and0 | s_CSAwallace_cla16_csa0_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa13_xor0 = s_CSAwallace_cla16_and_13_0 ^ s_CSAwallace_cla16_and_12_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa13_and0 = s_CSAwallace_cla16_and_13_0 & s_CSAwallace_cla16_and_12_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_and_11_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa13_and1 = s_CSAwallace_cla16_csa0_csa_component_fa13_xor0 & s_CSAwallace_cla16_and_11_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa13_or0 = s_CSAwallace_cla16_csa0_csa_component_fa13_and0 | s_CSAwallace_cla16_csa0_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa14_xor0 = s_CSAwallace_cla16_and_14_0 ^ s_CSAwallace_cla16_and_13_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa14_and0 = s_CSAwallace_cla16_and_14_0 & s_CSAwallace_cla16_and_13_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_and_12_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa14_and1 = s_CSAwallace_cla16_csa0_csa_component_fa14_xor0 & s_CSAwallace_cla16_and_12_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa14_or0 = s_CSAwallace_cla16_csa0_csa_component_fa14_and0 | s_CSAwallace_cla16_csa0_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa15_xor0 = s_CSAwallace_cla16_nand_15_0 ^ s_CSAwallace_cla16_and_14_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa15_and0 = s_CSAwallace_cla16_nand_15_0 & s_CSAwallace_cla16_and_14_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_and_13_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa15_and1 = s_CSAwallace_cla16_csa0_csa_component_fa15_xor0 & s_CSAwallace_cla16_and_13_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa15_or0 = s_CSAwallace_cla16_csa0_csa_component_fa15_and0 | s_CSAwallace_cla16_csa0_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa16_xor0 = ~s_CSAwallace_cla16_nand_15_1;
  assign s_CSAwallace_cla16_csa0_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa0_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_and_14_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa16_and1 = s_CSAwallace_cla16_csa0_csa_component_fa16_xor0 & s_CSAwallace_cla16_and_14_2;
  assign s_CSAwallace_cla16_csa0_csa_component_fa16_or0 = s_CSAwallace_cla16_nand_15_1 | s_CSAwallace_cla16_csa0_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa4_xor0 = s_CSAwallace_cla16_and_1_3 ^ s_CSAwallace_cla16_and_0_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa4_and0 = s_CSAwallace_cla16_and_1_3 & s_CSAwallace_cla16_and_0_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa5_xor0 = s_CSAwallace_cla16_and_2_3 ^ s_CSAwallace_cla16_and_1_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa5_and0 = s_CSAwallace_cla16_and_2_3 & s_CSAwallace_cla16_and_1_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa5_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa5_xor0 ^ s_CSAwallace_cla16_and_0_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa5_and1 = s_CSAwallace_cla16_csa1_csa_component_fa5_xor0 & s_CSAwallace_cla16_and_0_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa5_or0 = s_CSAwallace_cla16_csa1_csa_component_fa5_and0 | s_CSAwallace_cla16_csa1_csa_component_fa5_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa6_xor0 = s_CSAwallace_cla16_and_3_3 ^ s_CSAwallace_cla16_and_2_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa6_and0 = s_CSAwallace_cla16_and_3_3 & s_CSAwallace_cla16_and_2_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa6_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa6_xor0 ^ s_CSAwallace_cla16_and_1_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa6_and1 = s_CSAwallace_cla16_csa1_csa_component_fa6_xor0 & s_CSAwallace_cla16_and_1_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa6_or0 = s_CSAwallace_cla16_csa1_csa_component_fa6_and0 | s_CSAwallace_cla16_csa1_csa_component_fa6_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa7_xor0 = s_CSAwallace_cla16_and_4_3 ^ s_CSAwallace_cla16_and_3_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa7_and0 = s_CSAwallace_cla16_and_4_3 & s_CSAwallace_cla16_and_3_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa7_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa7_xor0 ^ s_CSAwallace_cla16_and_2_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa7_and1 = s_CSAwallace_cla16_csa1_csa_component_fa7_xor0 & s_CSAwallace_cla16_and_2_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa7_or0 = s_CSAwallace_cla16_csa1_csa_component_fa7_and0 | s_CSAwallace_cla16_csa1_csa_component_fa7_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa8_xor0 = s_CSAwallace_cla16_and_5_3 ^ s_CSAwallace_cla16_and_4_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa8_and0 = s_CSAwallace_cla16_and_5_3 & s_CSAwallace_cla16_and_4_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa8_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_and_3_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa8_and1 = s_CSAwallace_cla16_csa1_csa_component_fa8_xor0 & s_CSAwallace_cla16_and_3_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa8_or0 = s_CSAwallace_cla16_csa1_csa_component_fa8_and0 | s_CSAwallace_cla16_csa1_csa_component_fa8_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa9_xor0 = s_CSAwallace_cla16_and_6_3 ^ s_CSAwallace_cla16_and_5_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa9_and0 = s_CSAwallace_cla16_and_6_3 & s_CSAwallace_cla16_and_5_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa9_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_and_4_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa9_and1 = s_CSAwallace_cla16_csa1_csa_component_fa9_xor0 & s_CSAwallace_cla16_and_4_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa9_or0 = s_CSAwallace_cla16_csa1_csa_component_fa9_and0 | s_CSAwallace_cla16_csa1_csa_component_fa9_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa10_xor0 = s_CSAwallace_cla16_and_7_3 ^ s_CSAwallace_cla16_and_6_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa10_and0 = s_CSAwallace_cla16_and_7_3 & s_CSAwallace_cla16_and_6_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa10_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_and_5_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa10_and1 = s_CSAwallace_cla16_csa1_csa_component_fa10_xor0 & s_CSAwallace_cla16_and_5_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa10_or0 = s_CSAwallace_cla16_csa1_csa_component_fa10_and0 | s_CSAwallace_cla16_csa1_csa_component_fa10_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa11_xor0 = s_CSAwallace_cla16_and_8_3 ^ s_CSAwallace_cla16_and_7_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa11_and0 = s_CSAwallace_cla16_and_8_3 & s_CSAwallace_cla16_and_7_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_and_6_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa11_and1 = s_CSAwallace_cla16_csa1_csa_component_fa11_xor0 & s_CSAwallace_cla16_and_6_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa11_or0 = s_CSAwallace_cla16_csa1_csa_component_fa11_and0 | s_CSAwallace_cla16_csa1_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa12_xor0 = s_CSAwallace_cla16_and_9_3 ^ s_CSAwallace_cla16_and_8_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa12_and0 = s_CSAwallace_cla16_and_9_3 & s_CSAwallace_cla16_and_8_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_and_7_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa12_and1 = s_CSAwallace_cla16_csa1_csa_component_fa12_xor0 & s_CSAwallace_cla16_and_7_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa12_or0 = s_CSAwallace_cla16_csa1_csa_component_fa12_and0 | s_CSAwallace_cla16_csa1_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa13_xor0 = s_CSAwallace_cla16_and_10_3 ^ s_CSAwallace_cla16_and_9_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa13_and0 = s_CSAwallace_cla16_and_10_3 & s_CSAwallace_cla16_and_9_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_and_8_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa13_and1 = s_CSAwallace_cla16_csa1_csa_component_fa13_xor0 & s_CSAwallace_cla16_and_8_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa13_or0 = s_CSAwallace_cla16_csa1_csa_component_fa13_and0 | s_CSAwallace_cla16_csa1_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa14_xor0 = s_CSAwallace_cla16_and_11_3 ^ s_CSAwallace_cla16_and_10_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa14_and0 = s_CSAwallace_cla16_and_11_3 & s_CSAwallace_cla16_and_10_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_and_9_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa14_and1 = s_CSAwallace_cla16_csa1_csa_component_fa14_xor0 & s_CSAwallace_cla16_and_9_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa14_or0 = s_CSAwallace_cla16_csa1_csa_component_fa14_and0 | s_CSAwallace_cla16_csa1_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa15_xor0 = s_CSAwallace_cla16_and_12_3 ^ s_CSAwallace_cla16_and_11_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa15_and0 = s_CSAwallace_cla16_and_12_3 & s_CSAwallace_cla16_and_11_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_and_10_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa15_and1 = s_CSAwallace_cla16_csa1_csa_component_fa15_xor0 & s_CSAwallace_cla16_and_10_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa15_or0 = s_CSAwallace_cla16_csa1_csa_component_fa15_and0 | s_CSAwallace_cla16_csa1_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa16_xor0 = s_CSAwallace_cla16_and_13_3 ^ s_CSAwallace_cla16_and_12_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa16_and0 = s_CSAwallace_cla16_and_13_3 & s_CSAwallace_cla16_and_12_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_and_11_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa16_and1 = s_CSAwallace_cla16_csa1_csa_component_fa16_xor0 & s_CSAwallace_cla16_and_11_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa16_or0 = s_CSAwallace_cla16_csa1_csa_component_fa16_and0 | s_CSAwallace_cla16_csa1_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa17_xor0 = s_CSAwallace_cla16_and_14_3 ^ s_CSAwallace_cla16_and_13_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa17_and0 = s_CSAwallace_cla16_and_14_3 & s_CSAwallace_cla16_and_13_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_and_12_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa17_and1 = s_CSAwallace_cla16_csa1_csa_component_fa17_xor0 & s_CSAwallace_cla16_and_12_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa17_or0 = s_CSAwallace_cla16_csa1_csa_component_fa17_and0 | s_CSAwallace_cla16_csa1_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa18_xor0 = s_CSAwallace_cla16_nand_15_3 ^ s_CSAwallace_cla16_and_14_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa18_and0 = s_CSAwallace_cla16_nand_15_3 & s_CSAwallace_cla16_and_14_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_and_13_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa18_and1 = s_CSAwallace_cla16_csa1_csa_component_fa18_xor0 & s_CSAwallace_cla16_and_13_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa18_or0 = s_CSAwallace_cla16_csa1_csa_component_fa18_and0 | s_CSAwallace_cla16_csa1_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa1_csa_component_fa19_xor0 = ~s_CSAwallace_cla16_nand_15_4;
  assign s_CSAwallace_cla16_csa1_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa1_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_and_14_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa19_and1 = s_CSAwallace_cla16_csa1_csa_component_fa19_xor0 & s_CSAwallace_cla16_and_14_5;
  assign s_CSAwallace_cla16_csa1_csa_component_fa19_or0 = s_CSAwallace_cla16_nand_15_4 | s_CSAwallace_cla16_csa1_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa7_xor0 = s_CSAwallace_cla16_and_1_6 ^ s_CSAwallace_cla16_and_0_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa7_and0 = s_CSAwallace_cla16_and_1_6 & s_CSAwallace_cla16_and_0_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa8_xor0 = s_CSAwallace_cla16_and_2_6 ^ s_CSAwallace_cla16_and_1_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa8_and0 = s_CSAwallace_cla16_and_2_6 & s_CSAwallace_cla16_and_1_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa8_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_and_0_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa8_and1 = s_CSAwallace_cla16_csa2_csa_component_fa8_xor0 & s_CSAwallace_cla16_and_0_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa8_or0 = s_CSAwallace_cla16_csa2_csa_component_fa8_and0 | s_CSAwallace_cla16_csa2_csa_component_fa8_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa9_xor0 = s_CSAwallace_cla16_and_3_6 ^ s_CSAwallace_cla16_and_2_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa9_and0 = s_CSAwallace_cla16_and_3_6 & s_CSAwallace_cla16_and_2_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa9_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_and_1_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa9_and1 = s_CSAwallace_cla16_csa2_csa_component_fa9_xor0 & s_CSAwallace_cla16_and_1_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa9_or0 = s_CSAwallace_cla16_csa2_csa_component_fa9_and0 | s_CSAwallace_cla16_csa2_csa_component_fa9_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa10_xor0 = s_CSAwallace_cla16_and_4_6 ^ s_CSAwallace_cla16_and_3_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa10_and0 = s_CSAwallace_cla16_and_4_6 & s_CSAwallace_cla16_and_3_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa10_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_and_2_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa10_and1 = s_CSAwallace_cla16_csa2_csa_component_fa10_xor0 & s_CSAwallace_cla16_and_2_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa10_or0 = s_CSAwallace_cla16_csa2_csa_component_fa10_and0 | s_CSAwallace_cla16_csa2_csa_component_fa10_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa11_xor0 = s_CSAwallace_cla16_and_5_6 ^ s_CSAwallace_cla16_and_4_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa11_and0 = s_CSAwallace_cla16_and_5_6 & s_CSAwallace_cla16_and_4_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_and_3_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa11_and1 = s_CSAwallace_cla16_csa2_csa_component_fa11_xor0 & s_CSAwallace_cla16_and_3_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa11_or0 = s_CSAwallace_cla16_csa2_csa_component_fa11_and0 | s_CSAwallace_cla16_csa2_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa12_xor0 = s_CSAwallace_cla16_and_6_6 ^ s_CSAwallace_cla16_and_5_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa12_and0 = s_CSAwallace_cla16_and_6_6 & s_CSAwallace_cla16_and_5_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_and_4_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa12_and1 = s_CSAwallace_cla16_csa2_csa_component_fa12_xor0 & s_CSAwallace_cla16_and_4_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa12_or0 = s_CSAwallace_cla16_csa2_csa_component_fa12_and0 | s_CSAwallace_cla16_csa2_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa13_xor0 = s_CSAwallace_cla16_and_7_6 ^ s_CSAwallace_cla16_and_6_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa13_and0 = s_CSAwallace_cla16_and_7_6 & s_CSAwallace_cla16_and_6_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_and_5_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa13_and1 = s_CSAwallace_cla16_csa2_csa_component_fa13_xor0 & s_CSAwallace_cla16_and_5_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa13_or0 = s_CSAwallace_cla16_csa2_csa_component_fa13_and0 | s_CSAwallace_cla16_csa2_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa14_xor0 = s_CSAwallace_cla16_and_8_6 ^ s_CSAwallace_cla16_and_7_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa14_and0 = s_CSAwallace_cla16_and_8_6 & s_CSAwallace_cla16_and_7_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_and_6_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa14_and1 = s_CSAwallace_cla16_csa2_csa_component_fa14_xor0 & s_CSAwallace_cla16_and_6_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa14_or0 = s_CSAwallace_cla16_csa2_csa_component_fa14_and0 | s_CSAwallace_cla16_csa2_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa15_xor0 = s_CSAwallace_cla16_and_9_6 ^ s_CSAwallace_cla16_and_8_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa15_and0 = s_CSAwallace_cla16_and_9_6 & s_CSAwallace_cla16_and_8_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_and_7_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa15_and1 = s_CSAwallace_cla16_csa2_csa_component_fa15_xor0 & s_CSAwallace_cla16_and_7_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa15_or0 = s_CSAwallace_cla16_csa2_csa_component_fa15_and0 | s_CSAwallace_cla16_csa2_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa16_xor0 = s_CSAwallace_cla16_and_10_6 ^ s_CSAwallace_cla16_and_9_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa16_and0 = s_CSAwallace_cla16_and_10_6 & s_CSAwallace_cla16_and_9_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_and_8_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa16_and1 = s_CSAwallace_cla16_csa2_csa_component_fa16_xor0 & s_CSAwallace_cla16_and_8_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa16_or0 = s_CSAwallace_cla16_csa2_csa_component_fa16_and0 | s_CSAwallace_cla16_csa2_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa17_xor0 = s_CSAwallace_cla16_and_11_6 ^ s_CSAwallace_cla16_and_10_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa17_and0 = s_CSAwallace_cla16_and_11_6 & s_CSAwallace_cla16_and_10_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_and_9_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa17_and1 = s_CSAwallace_cla16_csa2_csa_component_fa17_xor0 & s_CSAwallace_cla16_and_9_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa17_or0 = s_CSAwallace_cla16_csa2_csa_component_fa17_and0 | s_CSAwallace_cla16_csa2_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa18_xor0 = s_CSAwallace_cla16_and_12_6 ^ s_CSAwallace_cla16_and_11_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa18_and0 = s_CSAwallace_cla16_and_12_6 & s_CSAwallace_cla16_and_11_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_and_10_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa18_and1 = s_CSAwallace_cla16_csa2_csa_component_fa18_xor0 & s_CSAwallace_cla16_and_10_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa18_or0 = s_CSAwallace_cla16_csa2_csa_component_fa18_and0 | s_CSAwallace_cla16_csa2_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa19_xor0 = s_CSAwallace_cla16_and_13_6 ^ s_CSAwallace_cla16_and_12_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa19_and0 = s_CSAwallace_cla16_and_13_6 & s_CSAwallace_cla16_and_12_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_and_11_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa19_and1 = s_CSAwallace_cla16_csa2_csa_component_fa19_xor0 & s_CSAwallace_cla16_and_11_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa19_or0 = s_CSAwallace_cla16_csa2_csa_component_fa19_and0 | s_CSAwallace_cla16_csa2_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa20_xor0 = s_CSAwallace_cla16_and_14_6 ^ s_CSAwallace_cla16_and_13_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa20_and0 = s_CSAwallace_cla16_and_14_6 & s_CSAwallace_cla16_and_13_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_and_12_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa20_and1 = s_CSAwallace_cla16_csa2_csa_component_fa20_xor0 & s_CSAwallace_cla16_and_12_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa20_or0 = s_CSAwallace_cla16_csa2_csa_component_fa20_and0 | s_CSAwallace_cla16_csa2_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa21_xor0 = s_CSAwallace_cla16_nand_15_6 ^ s_CSAwallace_cla16_and_14_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa21_and0 = s_CSAwallace_cla16_nand_15_6 & s_CSAwallace_cla16_and_14_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_and_13_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa21_and1 = s_CSAwallace_cla16_csa2_csa_component_fa21_xor0 & s_CSAwallace_cla16_and_13_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa21_or0 = s_CSAwallace_cla16_csa2_csa_component_fa21_and0 | s_CSAwallace_cla16_csa2_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa2_csa_component_fa22_xor0 = ~s_CSAwallace_cla16_nand_15_7;
  assign s_CSAwallace_cla16_csa2_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa2_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_and_14_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa22_and1 = s_CSAwallace_cla16_csa2_csa_component_fa22_xor0 & s_CSAwallace_cla16_and_14_8;
  assign s_CSAwallace_cla16_csa2_csa_component_fa22_or0 = s_CSAwallace_cla16_nand_15_7 | s_CSAwallace_cla16_csa2_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa10_xor0 = s_CSAwallace_cla16_and_1_9 ^ s_CSAwallace_cla16_and_0_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa10_and0 = s_CSAwallace_cla16_and_1_9 & s_CSAwallace_cla16_and_0_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa11_xor0 = s_CSAwallace_cla16_and_2_9 ^ s_CSAwallace_cla16_and_1_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa11_and0 = s_CSAwallace_cla16_and_2_9 & s_CSAwallace_cla16_and_1_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_and_0_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa11_and1 = s_CSAwallace_cla16_csa3_csa_component_fa11_xor0 & s_CSAwallace_cla16_and_0_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa11_or0 = s_CSAwallace_cla16_csa3_csa_component_fa11_and0 | s_CSAwallace_cla16_csa3_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa12_xor0 = s_CSAwallace_cla16_and_3_9 ^ s_CSAwallace_cla16_and_2_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa12_and0 = s_CSAwallace_cla16_and_3_9 & s_CSAwallace_cla16_and_2_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_and_1_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa12_and1 = s_CSAwallace_cla16_csa3_csa_component_fa12_xor0 & s_CSAwallace_cla16_and_1_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa12_or0 = s_CSAwallace_cla16_csa3_csa_component_fa12_and0 | s_CSAwallace_cla16_csa3_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa13_xor0 = s_CSAwallace_cla16_and_4_9 ^ s_CSAwallace_cla16_and_3_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa13_and0 = s_CSAwallace_cla16_and_4_9 & s_CSAwallace_cla16_and_3_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_and_2_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa13_and1 = s_CSAwallace_cla16_csa3_csa_component_fa13_xor0 & s_CSAwallace_cla16_and_2_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa13_or0 = s_CSAwallace_cla16_csa3_csa_component_fa13_and0 | s_CSAwallace_cla16_csa3_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa14_xor0 = s_CSAwallace_cla16_and_5_9 ^ s_CSAwallace_cla16_and_4_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa14_and0 = s_CSAwallace_cla16_and_5_9 & s_CSAwallace_cla16_and_4_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_and_3_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa14_and1 = s_CSAwallace_cla16_csa3_csa_component_fa14_xor0 & s_CSAwallace_cla16_and_3_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa14_or0 = s_CSAwallace_cla16_csa3_csa_component_fa14_and0 | s_CSAwallace_cla16_csa3_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa15_xor0 = s_CSAwallace_cla16_and_6_9 ^ s_CSAwallace_cla16_and_5_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa15_and0 = s_CSAwallace_cla16_and_6_9 & s_CSAwallace_cla16_and_5_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_and_4_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa15_and1 = s_CSAwallace_cla16_csa3_csa_component_fa15_xor0 & s_CSAwallace_cla16_and_4_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa15_or0 = s_CSAwallace_cla16_csa3_csa_component_fa15_and0 | s_CSAwallace_cla16_csa3_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa16_xor0 = s_CSAwallace_cla16_and_7_9 ^ s_CSAwallace_cla16_and_6_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa16_and0 = s_CSAwallace_cla16_and_7_9 & s_CSAwallace_cla16_and_6_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_and_5_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa16_and1 = s_CSAwallace_cla16_csa3_csa_component_fa16_xor0 & s_CSAwallace_cla16_and_5_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa16_or0 = s_CSAwallace_cla16_csa3_csa_component_fa16_and0 | s_CSAwallace_cla16_csa3_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa17_xor0 = s_CSAwallace_cla16_and_8_9 ^ s_CSAwallace_cla16_and_7_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa17_and0 = s_CSAwallace_cla16_and_8_9 & s_CSAwallace_cla16_and_7_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_and_6_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa17_and1 = s_CSAwallace_cla16_csa3_csa_component_fa17_xor0 & s_CSAwallace_cla16_and_6_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa17_or0 = s_CSAwallace_cla16_csa3_csa_component_fa17_and0 | s_CSAwallace_cla16_csa3_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa18_xor0 = s_CSAwallace_cla16_and_9_9 ^ s_CSAwallace_cla16_and_8_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa18_and0 = s_CSAwallace_cla16_and_9_9 & s_CSAwallace_cla16_and_8_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_and_7_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa18_and1 = s_CSAwallace_cla16_csa3_csa_component_fa18_xor0 & s_CSAwallace_cla16_and_7_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa18_or0 = s_CSAwallace_cla16_csa3_csa_component_fa18_and0 | s_CSAwallace_cla16_csa3_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa19_xor0 = s_CSAwallace_cla16_and_10_9 ^ s_CSAwallace_cla16_and_9_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa19_and0 = s_CSAwallace_cla16_and_10_9 & s_CSAwallace_cla16_and_9_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_and_8_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa19_and1 = s_CSAwallace_cla16_csa3_csa_component_fa19_xor0 & s_CSAwallace_cla16_and_8_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa19_or0 = s_CSAwallace_cla16_csa3_csa_component_fa19_and0 | s_CSAwallace_cla16_csa3_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa20_xor0 = s_CSAwallace_cla16_and_11_9 ^ s_CSAwallace_cla16_and_10_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa20_and0 = s_CSAwallace_cla16_and_11_9 & s_CSAwallace_cla16_and_10_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_and_9_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa20_and1 = s_CSAwallace_cla16_csa3_csa_component_fa20_xor0 & s_CSAwallace_cla16_and_9_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa20_or0 = s_CSAwallace_cla16_csa3_csa_component_fa20_and0 | s_CSAwallace_cla16_csa3_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa21_xor0 = s_CSAwallace_cla16_and_12_9 ^ s_CSAwallace_cla16_and_11_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa21_and0 = s_CSAwallace_cla16_and_12_9 & s_CSAwallace_cla16_and_11_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_and_10_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa21_and1 = s_CSAwallace_cla16_csa3_csa_component_fa21_xor0 & s_CSAwallace_cla16_and_10_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa21_or0 = s_CSAwallace_cla16_csa3_csa_component_fa21_and0 | s_CSAwallace_cla16_csa3_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa22_xor0 = s_CSAwallace_cla16_and_13_9 ^ s_CSAwallace_cla16_and_12_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa22_and0 = s_CSAwallace_cla16_and_13_9 & s_CSAwallace_cla16_and_12_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_and_11_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa22_and1 = s_CSAwallace_cla16_csa3_csa_component_fa22_xor0 & s_CSAwallace_cla16_and_11_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa22_or0 = s_CSAwallace_cla16_csa3_csa_component_fa22_and0 | s_CSAwallace_cla16_csa3_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa23_xor0 = s_CSAwallace_cla16_and_14_9 ^ s_CSAwallace_cla16_and_13_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa23_and0 = s_CSAwallace_cla16_and_14_9 & s_CSAwallace_cla16_and_13_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_and_12_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa23_and1 = s_CSAwallace_cla16_csa3_csa_component_fa23_xor0 & s_CSAwallace_cla16_and_12_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa23_or0 = s_CSAwallace_cla16_csa3_csa_component_fa23_and0 | s_CSAwallace_cla16_csa3_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa24_xor0 = s_CSAwallace_cla16_nand_15_9 ^ s_CSAwallace_cla16_and_14_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa24_and0 = s_CSAwallace_cla16_nand_15_9 & s_CSAwallace_cla16_and_14_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa24_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa24_xor0 ^ s_CSAwallace_cla16_and_13_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa24_and1 = s_CSAwallace_cla16_csa3_csa_component_fa24_xor0 & s_CSAwallace_cla16_and_13_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa24_or0 = s_CSAwallace_cla16_csa3_csa_component_fa24_and0 | s_CSAwallace_cla16_csa3_csa_component_fa24_and1;
  assign s_CSAwallace_cla16_csa3_csa_component_fa25_xor0 = ~s_CSAwallace_cla16_nand_15_10;
  assign s_CSAwallace_cla16_csa3_csa_component_fa25_xor1 = s_CSAwallace_cla16_csa3_csa_component_fa25_xor0 ^ s_CSAwallace_cla16_and_14_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa25_and1 = s_CSAwallace_cla16_csa3_csa_component_fa25_xor0 & s_CSAwallace_cla16_and_14_11;
  assign s_CSAwallace_cla16_csa3_csa_component_fa25_or0 = s_CSAwallace_cla16_nand_15_10 | s_CSAwallace_cla16_csa3_csa_component_fa25_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa13_xor0 = s_CSAwallace_cla16_and_1_12 ^ s_CSAwallace_cla16_and_0_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa13_and0 = s_CSAwallace_cla16_and_1_12 & s_CSAwallace_cla16_and_0_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa14_xor0 = s_CSAwallace_cla16_and_2_12 ^ s_CSAwallace_cla16_and_1_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa14_and0 = s_CSAwallace_cla16_and_2_12 & s_CSAwallace_cla16_and_1_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_and_0_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa14_and1 = s_CSAwallace_cla16_csa4_csa_component_fa14_xor0 & s_CSAwallace_cla16_and_0_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa14_or0 = s_CSAwallace_cla16_csa4_csa_component_fa14_and0 | s_CSAwallace_cla16_csa4_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa15_xor0 = s_CSAwallace_cla16_and_3_12 ^ s_CSAwallace_cla16_and_2_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa15_and0 = s_CSAwallace_cla16_and_3_12 & s_CSAwallace_cla16_and_2_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_and_1_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa15_and1 = s_CSAwallace_cla16_csa4_csa_component_fa15_xor0 & s_CSAwallace_cla16_and_1_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa15_or0 = s_CSAwallace_cla16_csa4_csa_component_fa15_and0 | s_CSAwallace_cla16_csa4_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa16_xor0 = s_CSAwallace_cla16_and_4_12 ^ s_CSAwallace_cla16_and_3_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa16_and0 = s_CSAwallace_cla16_and_4_12 & s_CSAwallace_cla16_and_3_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_and_2_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa16_and1 = s_CSAwallace_cla16_csa4_csa_component_fa16_xor0 & s_CSAwallace_cla16_and_2_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa16_or0 = s_CSAwallace_cla16_csa4_csa_component_fa16_and0 | s_CSAwallace_cla16_csa4_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa17_xor0 = s_CSAwallace_cla16_and_5_12 ^ s_CSAwallace_cla16_and_4_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa17_and0 = s_CSAwallace_cla16_and_5_12 & s_CSAwallace_cla16_and_4_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_and_3_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa17_and1 = s_CSAwallace_cla16_csa4_csa_component_fa17_xor0 & s_CSAwallace_cla16_and_3_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa17_or0 = s_CSAwallace_cla16_csa4_csa_component_fa17_and0 | s_CSAwallace_cla16_csa4_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa18_xor0 = s_CSAwallace_cla16_and_6_12 ^ s_CSAwallace_cla16_and_5_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa18_and0 = s_CSAwallace_cla16_and_6_12 & s_CSAwallace_cla16_and_5_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_and_4_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa18_and1 = s_CSAwallace_cla16_csa4_csa_component_fa18_xor0 & s_CSAwallace_cla16_and_4_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa18_or0 = s_CSAwallace_cla16_csa4_csa_component_fa18_and0 | s_CSAwallace_cla16_csa4_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa19_xor0 = s_CSAwallace_cla16_and_7_12 ^ s_CSAwallace_cla16_and_6_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa19_and0 = s_CSAwallace_cla16_and_7_12 & s_CSAwallace_cla16_and_6_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_and_5_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa19_and1 = s_CSAwallace_cla16_csa4_csa_component_fa19_xor0 & s_CSAwallace_cla16_and_5_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa19_or0 = s_CSAwallace_cla16_csa4_csa_component_fa19_and0 | s_CSAwallace_cla16_csa4_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa20_xor0 = s_CSAwallace_cla16_and_8_12 ^ s_CSAwallace_cla16_and_7_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa20_and0 = s_CSAwallace_cla16_and_8_12 & s_CSAwallace_cla16_and_7_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_and_6_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa20_and1 = s_CSAwallace_cla16_csa4_csa_component_fa20_xor0 & s_CSAwallace_cla16_and_6_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa20_or0 = s_CSAwallace_cla16_csa4_csa_component_fa20_and0 | s_CSAwallace_cla16_csa4_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa21_xor0 = s_CSAwallace_cla16_and_9_12 ^ s_CSAwallace_cla16_and_8_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa21_and0 = s_CSAwallace_cla16_and_9_12 & s_CSAwallace_cla16_and_8_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_and_7_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa21_and1 = s_CSAwallace_cla16_csa4_csa_component_fa21_xor0 & s_CSAwallace_cla16_and_7_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa21_or0 = s_CSAwallace_cla16_csa4_csa_component_fa21_and0 | s_CSAwallace_cla16_csa4_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa22_xor0 = s_CSAwallace_cla16_and_10_12 ^ s_CSAwallace_cla16_and_9_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa22_and0 = s_CSAwallace_cla16_and_10_12 & s_CSAwallace_cla16_and_9_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_and_8_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa22_and1 = s_CSAwallace_cla16_csa4_csa_component_fa22_xor0 & s_CSAwallace_cla16_and_8_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa22_or0 = s_CSAwallace_cla16_csa4_csa_component_fa22_and0 | s_CSAwallace_cla16_csa4_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa23_xor0 = s_CSAwallace_cla16_and_11_12 ^ s_CSAwallace_cla16_and_10_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa23_and0 = s_CSAwallace_cla16_and_11_12 & s_CSAwallace_cla16_and_10_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_and_9_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa23_and1 = s_CSAwallace_cla16_csa4_csa_component_fa23_xor0 & s_CSAwallace_cla16_and_9_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa23_or0 = s_CSAwallace_cla16_csa4_csa_component_fa23_and0 | s_CSAwallace_cla16_csa4_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa24_xor0 = s_CSAwallace_cla16_and_12_12 ^ s_CSAwallace_cla16_and_11_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa24_and0 = s_CSAwallace_cla16_and_12_12 & s_CSAwallace_cla16_and_11_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa24_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa24_xor0 ^ s_CSAwallace_cla16_and_10_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa24_and1 = s_CSAwallace_cla16_csa4_csa_component_fa24_xor0 & s_CSAwallace_cla16_and_10_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa24_or0 = s_CSAwallace_cla16_csa4_csa_component_fa24_and0 | s_CSAwallace_cla16_csa4_csa_component_fa24_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa25_xor0 = s_CSAwallace_cla16_and_13_12 ^ s_CSAwallace_cla16_and_12_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa25_and0 = s_CSAwallace_cla16_and_13_12 & s_CSAwallace_cla16_and_12_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa25_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa25_xor0 ^ s_CSAwallace_cla16_and_11_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa25_and1 = s_CSAwallace_cla16_csa4_csa_component_fa25_xor0 & s_CSAwallace_cla16_and_11_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa25_or0 = s_CSAwallace_cla16_csa4_csa_component_fa25_and0 | s_CSAwallace_cla16_csa4_csa_component_fa25_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa26_xor0 = s_CSAwallace_cla16_and_14_12 ^ s_CSAwallace_cla16_and_13_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa26_and0 = s_CSAwallace_cla16_and_14_12 & s_CSAwallace_cla16_and_13_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa26_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa26_xor0 ^ s_CSAwallace_cla16_and_12_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa26_and1 = s_CSAwallace_cla16_csa4_csa_component_fa26_xor0 & s_CSAwallace_cla16_and_12_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa26_or0 = s_CSAwallace_cla16_csa4_csa_component_fa26_and0 | s_CSAwallace_cla16_csa4_csa_component_fa26_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa27_xor0 = s_CSAwallace_cla16_nand_15_12 ^ s_CSAwallace_cla16_and_14_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa27_and0 = s_CSAwallace_cla16_nand_15_12 & s_CSAwallace_cla16_and_14_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa27_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa27_xor0 ^ s_CSAwallace_cla16_and_13_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa27_and1 = s_CSAwallace_cla16_csa4_csa_component_fa27_xor0 & s_CSAwallace_cla16_and_13_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa27_or0 = s_CSAwallace_cla16_csa4_csa_component_fa27_and0 | s_CSAwallace_cla16_csa4_csa_component_fa27_and1;
  assign s_CSAwallace_cla16_csa4_csa_component_fa28_xor0 = ~s_CSAwallace_cla16_nand_15_13;
  assign s_CSAwallace_cla16_csa4_csa_component_fa28_xor1 = s_CSAwallace_cla16_csa4_csa_component_fa28_xor0 ^ s_CSAwallace_cla16_and_14_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa28_and1 = s_CSAwallace_cla16_csa4_csa_component_fa28_xor0 & s_CSAwallace_cla16_and_14_14;
  assign s_CSAwallace_cla16_csa4_csa_component_fa28_or0 = s_CSAwallace_cla16_nand_15_13 | s_CSAwallace_cla16_csa4_csa_component_fa28_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa2_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa2_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa1_and0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa2_and0 = s_CSAwallace_cla16_csa0_csa_component_fa2_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa1_and0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa3_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa3_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa2_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa3_and0 = s_CSAwallace_cla16_csa0_csa_component_fa3_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa2_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa3_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa3_xor0 ^ s_CSAwallace_cla16_and_0_3;
  assign s_CSAwallace_cla16_csa5_csa_component_fa3_and1 = s_CSAwallace_cla16_csa5_csa_component_fa3_xor0 & s_CSAwallace_cla16_and_0_3;
  assign s_CSAwallace_cla16_csa5_csa_component_fa3_or0 = s_CSAwallace_cla16_csa5_csa_component_fa3_and0 | s_CSAwallace_cla16_csa5_csa_component_fa3_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa4_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa4_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa3_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa4_and0 = s_CSAwallace_cla16_csa0_csa_component_fa4_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa3_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa4_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa4_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa4_xor0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa4_and1 = s_CSAwallace_cla16_csa5_csa_component_fa4_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa4_xor0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa4_or0 = s_CSAwallace_cla16_csa5_csa_component_fa4_and0 | s_CSAwallace_cla16_csa5_csa_component_fa4_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa5_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa5_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa4_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa5_and0 = s_CSAwallace_cla16_csa0_csa_component_fa5_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa4_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa5_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa5_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa5_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa5_and1 = s_CSAwallace_cla16_csa5_csa_component_fa5_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa5_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa5_or0 = s_CSAwallace_cla16_csa5_csa_component_fa5_and0 | s_CSAwallace_cla16_csa5_csa_component_fa5_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa6_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa6_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa5_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa6_and0 = s_CSAwallace_cla16_csa0_csa_component_fa6_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa5_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa6_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa6_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa6_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa6_and1 = s_CSAwallace_cla16_csa5_csa_component_fa6_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa6_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa6_or0 = s_CSAwallace_cla16_csa5_csa_component_fa6_and0 | s_CSAwallace_cla16_csa5_csa_component_fa6_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa7_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa7_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa6_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa7_and0 = s_CSAwallace_cla16_csa0_csa_component_fa7_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa6_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa7_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa7_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa7_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa7_and1 = s_CSAwallace_cla16_csa5_csa_component_fa7_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa7_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa7_or0 = s_CSAwallace_cla16_csa5_csa_component_fa7_and0 | s_CSAwallace_cla16_csa5_csa_component_fa7_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa8_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa8_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa7_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa8_and0 = s_CSAwallace_cla16_csa0_csa_component_fa8_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa7_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa8_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa8_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa8_and1 = s_CSAwallace_cla16_csa5_csa_component_fa8_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa8_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa8_or0 = s_CSAwallace_cla16_csa5_csa_component_fa8_and0 | s_CSAwallace_cla16_csa5_csa_component_fa8_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa9_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa9_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa9_and0 = s_CSAwallace_cla16_csa0_csa_component_fa9_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa9_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa9_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa9_and1 = s_CSAwallace_cla16_csa5_csa_component_fa9_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa9_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa9_or0 = s_CSAwallace_cla16_csa5_csa_component_fa9_and0 | s_CSAwallace_cla16_csa5_csa_component_fa9_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa10_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa10_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa10_and0 = s_CSAwallace_cla16_csa0_csa_component_fa10_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa10_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa10_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa10_and1 = s_CSAwallace_cla16_csa5_csa_component_fa10_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa10_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa10_or0 = s_CSAwallace_cla16_csa5_csa_component_fa10_and0 | s_CSAwallace_cla16_csa5_csa_component_fa10_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa11_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa11_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa11_and0 = s_CSAwallace_cla16_csa0_csa_component_fa11_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa11_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa11_and1 = s_CSAwallace_cla16_csa5_csa_component_fa11_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa11_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa11_or0 = s_CSAwallace_cla16_csa5_csa_component_fa11_and0 | s_CSAwallace_cla16_csa5_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa12_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa12_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa12_and0 = s_CSAwallace_cla16_csa0_csa_component_fa12_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa12_and1 = s_CSAwallace_cla16_csa5_csa_component_fa12_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa12_or0 = s_CSAwallace_cla16_csa5_csa_component_fa12_and0 | s_CSAwallace_cla16_csa5_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa13_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa13_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa13_and0 = s_CSAwallace_cla16_csa0_csa_component_fa13_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa13_and1 = s_CSAwallace_cla16_csa5_csa_component_fa13_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa13_or0 = s_CSAwallace_cla16_csa5_csa_component_fa13_and0 | s_CSAwallace_cla16_csa5_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa14_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa14_and0 = s_CSAwallace_cla16_csa0_csa_component_fa14_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa14_and1 = s_CSAwallace_cla16_csa5_csa_component_fa14_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa14_or0 = s_CSAwallace_cla16_csa5_csa_component_fa14_and0 | s_CSAwallace_cla16_csa5_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa15_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa15_and0 = s_CSAwallace_cla16_csa0_csa_component_fa15_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa15_and1 = s_CSAwallace_cla16_csa5_csa_component_fa15_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa15_or0 = s_CSAwallace_cla16_csa5_csa_component_fa15_and0 | s_CSAwallace_cla16_csa5_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa0_csa_component_fa16_xor1 ^ s_CSAwallace_cla16_csa0_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa16_and0 = s_CSAwallace_cla16_csa0_csa_component_fa16_xor1 & s_CSAwallace_cla16_csa0_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa16_and1 = s_CSAwallace_cla16_csa5_csa_component_fa16_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa16_or0 = s_CSAwallace_cla16_csa5_csa_component_fa16_and0 | s_CSAwallace_cla16_csa5_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa17_xor0 = s_CSAwallace_cla16_nand_15_2 ^ s_CSAwallace_cla16_csa0_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa17_and0 = s_CSAwallace_cla16_nand_15_2 & s_CSAwallace_cla16_csa0_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa5_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa5_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa17_and1 = s_CSAwallace_cla16_csa5_csa_component_fa17_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa5_csa_component_fa17_or0 = s_CSAwallace_cla16_csa5_csa_component_fa17_and0 | s_CSAwallace_cla16_csa5_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa6_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa5_or0 ^ s_CSAwallace_cla16_and_0_6;
  assign s_CSAwallace_cla16_csa6_csa_component_fa6_and0 = s_CSAwallace_cla16_csa1_csa_component_fa5_or0 & s_CSAwallace_cla16_and_0_6;
  assign s_CSAwallace_cla16_csa6_csa_component_fa7_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa6_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa7_xor0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa7_and0 = s_CSAwallace_cla16_csa1_csa_component_fa6_or0 & s_CSAwallace_cla16_csa2_csa_component_fa7_xor0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa8_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa7_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa8_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa8_and0 = s_CSAwallace_cla16_csa1_csa_component_fa7_or0 & s_CSAwallace_cla16_csa2_csa_component_fa8_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa8_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa8_and1 = s_CSAwallace_cla16_csa6_csa_component_fa8_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa8_or0 = s_CSAwallace_cla16_csa6_csa_component_fa8_and0 | s_CSAwallace_cla16_csa6_csa_component_fa8_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa9_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa8_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa9_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa9_and0 = s_CSAwallace_cla16_csa1_csa_component_fa8_or0 & s_CSAwallace_cla16_csa2_csa_component_fa9_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa9_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa9_and1 = s_CSAwallace_cla16_csa6_csa_component_fa9_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa9_or0 = s_CSAwallace_cla16_csa6_csa_component_fa9_and0 | s_CSAwallace_cla16_csa6_csa_component_fa9_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa10_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa9_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa10_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa10_and0 = s_CSAwallace_cla16_csa1_csa_component_fa9_or0 & s_CSAwallace_cla16_csa2_csa_component_fa10_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa10_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa10_and1 = s_CSAwallace_cla16_csa6_csa_component_fa10_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa10_or0 = s_CSAwallace_cla16_csa6_csa_component_fa10_and0 | s_CSAwallace_cla16_csa6_csa_component_fa10_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa11_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa10_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa11_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa11_and0 = s_CSAwallace_cla16_csa1_csa_component_fa10_or0 & s_CSAwallace_cla16_csa2_csa_component_fa11_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa11_and1 = s_CSAwallace_cla16_csa6_csa_component_fa11_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa11_or0 = s_CSAwallace_cla16_csa6_csa_component_fa11_and0 | s_CSAwallace_cla16_csa6_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa12_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa11_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa12_and0 = s_CSAwallace_cla16_csa1_csa_component_fa11_or0 & s_CSAwallace_cla16_csa2_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa12_and1 = s_CSAwallace_cla16_csa6_csa_component_fa12_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa12_or0 = s_CSAwallace_cla16_csa6_csa_component_fa12_and0 | s_CSAwallace_cla16_csa6_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa13_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa12_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa13_and0 = s_CSAwallace_cla16_csa1_csa_component_fa12_or0 & s_CSAwallace_cla16_csa2_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa13_and1 = s_CSAwallace_cla16_csa6_csa_component_fa13_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa13_or0 = s_CSAwallace_cla16_csa6_csa_component_fa13_and0 | s_CSAwallace_cla16_csa6_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa13_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa14_and0 = s_CSAwallace_cla16_csa1_csa_component_fa13_or0 & s_CSAwallace_cla16_csa2_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa14_and1 = s_CSAwallace_cla16_csa6_csa_component_fa14_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa14_or0 = s_CSAwallace_cla16_csa6_csa_component_fa14_and0 | s_CSAwallace_cla16_csa6_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa14_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa15_and0 = s_CSAwallace_cla16_csa1_csa_component_fa14_or0 & s_CSAwallace_cla16_csa2_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa15_and1 = s_CSAwallace_cla16_csa6_csa_component_fa15_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa15_or0 = s_CSAwallace_cla16_csa6_csa_component_fa15_and0 | s_CSAwallace_cla16_csa6_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa15_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa16_and0 = s_CSAwallace_cla16_csa1_csa_component_fa15_or0 & s_CSAwallace_cla16_csa2_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa16_and1 = s_CSAwallace_cla16_csa6_csa_component_fa16_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa16_or0 = s_CSAwallace_cla16_csa6_csa_component_fa16_and0 | s_CSAwallace_cla16_csa6_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa17_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa16_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa17_and0 = s_CSAwallace_cla16_csa1_csa_component_fa16_or0 & s_CSAwallace_cla16_csa2_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa17_and1 = s_CSAwallace_cla16_csa6_csa_component_fa17_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa17_or0 = s_CSAwallace_cla16_csa6_csa_component_fa17_and0 | s_CSAwallace_cla16_csa6_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa18_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa17_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa18_and0 = s_CSAwallace_cla16_csa1_csa_component_fa17_or0 & s_CSAwallace_cla16_csa2_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa18_and1 = s_CSAwallace_cla16_csa6_csa_component_fa18_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa18_or0 = s_CSAwallace_cla16_csa6_csa_component_fa18_and0 | s_CSAwallace_cla16_csa6_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa19_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa18_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa19_and0 = s_CSAwallace_cla16_csa1_csa_component_fa18_or0 & s_CSAwallace_cla16_csa2_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa19_and1 = s_CSAwallace_cla16_csa6_csa_component_fa19_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa19_or0 = s_CSAwallace_cla16_csa6_csa_component_fa19_and0 | s_CSAwallace_cla16_csa6_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa20_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa19_or0 ^ s_CSAwallace_cla16_csa2_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa20_and0 = s_CSAwallace_cla16_csa1_csa_component_fa19_or0 & s_CSAwallace_cla16_csa2_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa20_and1 = s_CSAwallace_cla16_csa6_csa_component_fa20_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa20_or0 = s_CSAwallace_cla16_csa6_csa_component_fa20_and0 | s_CSAwallace_cla16_csa6_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa21_xor0 = ~s_CSAwallace_cla16_csa2_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa21_and1 = s_CSAwallace_cla16_csa6_csa_component_fa21_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa21_or0 = s_CSAwallace_cla16_csa2_csa_component_fa21_xor1 | s_CSAwallace_cla16_csa6_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa22_xor0 = ~s_CSAwallace_cla16_csa2_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa22_and1 = s_CSAwallace_cla16_csa6_csa_component_fa22_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa22_or0 = s_CSAwallace_cla16_csa2_csa_component_fa22_xor1 | s_CSAwallace_cla16_csa6_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa6_csa_component_fa23_xor0 = ~s_CSAwallace_cla16_nand_15_8;
  assign s_CSAwallace_cla16_csa6_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa6_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_csa2_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa23_and1 = s_CSAwallace_cla16_csa6_csa_component_fa23_xor0 & s_CSAwallace_cla16_csa2_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa6_csa_component_fa23_or0 = s_CSAwallace_cla16_nand_15_8 | s_CSAwallace_cla16_csa6_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa11_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa11_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa10_and0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa11_and0 = s_CSAwallace_cla16_csa3_csa_component_fa11_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa10_and0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa12_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa12_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa12_and0 = s_CSAwallace_cla16_csa3_csa_component_fa12_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_and_0_12;
  assign s_CSAwallace_cla16_csa7_csa_component_fa12_and1 = s_CSAwallace_cla16_csa7_csa_component_fa12_xor0 & s_CSAwallace_cla16_and_0_12;
  assign s_CSAwallace_cla16_csa7_csa_component_fa12_or0 = s_CSAwallace_cla16_csa7_csa_component_fa12_and0 | s_CSAwallace_cla16_csa7_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa13_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa13_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa13_and0 = s_CSAwallace_cla16_csa3_csa_component_fa13_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa13_xor0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa13_and1 = s_CSAwallace_cla16_csa7_csa_component_fa13_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa13_xor0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa13_or0 = s_CSAwallace_cla16_csa7_csa_component_fa13_and0 | s_CSAwallace_cla16_csa7_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa14_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa14_and0 = s_CSAwallace_cla16_csa3_csa_component_fa14_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa14_and1 = s_CSAwallace_cla16_csa7_csa_component_fa14_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa14_or0 = s_CSAwallace_cla16_csa7_csa_component_fa14_and0 | s_CSAwallace_cla16_csa7_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa15_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa15_and0 = s_CSAwallace_cla16_csa3_csa_component_fa15_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa15_and1 = s_CSAwallace_cla16_csa7_csa_component_fa15_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa15_or0 = s_CSAwallace_cla16_csa7_csa_component_fa15_and0 | s_CSAwallace_cla16_csa7_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa16_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa16_and0 = s_CSAwallace_cla16_csa3_csa_component_fa16_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa16_and1 = s_CSAwallace_cla16_csa7_csa_component_fa16_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa16_or0 = s_CSAwallace_cla16_csa7_csa_component_fa16_and0 | s_CSAwallace_cla16_csa7_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa17_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa17_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa17_and0 = s_CSAwallace_cla16_csa3_csa_component_fa17_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa17_and1 = s_CSAwallace_cla16_csa7_csa_component_fa17_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa17_or0 = s_CSAwallace_cla16_csa7_csa_component_fa17_and0 | s_CSAwallace_cla16_csa7_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa18_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa18_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa18_and0 = s_CSAwallace_cla16_csa3_csa_component_fa18_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa18_and1 = s_CSAwallace_cla16_csa7_csa_component_fa18_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa18_or0 = s_CSAwallace_cla16_csa7_csa_component_fa18_and0 | s_CSAwallace_cla16_csa7_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa19_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa19_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa19_and0 = s_CSAwallace_cla16_csa3_csa_component_fa19_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa19_and1 = s_CSAwallace_cla16_csa7_csa_component_fa19_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa19_or0 = s_CSAwallace_cla16_csa7_csa_component_fa19_and0 | s_CSAwallace_cla16_csa7_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa20_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa20_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa20_and0 = s_CSAwallace_cla16_csa3_csa_component_fa20_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa20_and1 = s_CSAwallace_cla16_csa7_csa_component_fa20_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa20_or0 = s_CSAwallace_cla16_csa7_csa_component_fa20_and0 | s_CSAwallace_cla16_csa7_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa21_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa21_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa21_and0 = s_CSAwallace_cla16_csa3_csa_component_fa21_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa21_and1 = s_CSAwallace_cla16_csa7_csa_component_fa21_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa21_or0 = s_CSAwallace_cla16_csa7_csa_component_fa21_and0 | s_CSAwallace_cla16_csa7_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa22_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa22_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa22_and0 = s_CSAwallace_cla16_csa3_csa_component_fa22_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa22_and1 = s_CSAwallace_cla16_csa7_csa_component_fa22_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa22_or0 = s_CSAwallace_cla16_csa7_csa_component_fa22_and0 | s_CSAwallace_cla16_csa7_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa23_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa23_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa23_and0 = s_CSAwallace_cla16_csa3_csa_component_fa23_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa23_and1 = s_CSAwallace_cla16_csa7_csa_component_fa23_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa23_or0 = s_CSAwallace_cla16_csa7_csa_component_fa23_and0 | s_CSAwallace_cla16_csa7_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa24_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa24_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa24_and0 = s_CSAwallace_cla16_csa3_csa_component_fa24_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa24_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa24_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa24_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa24_and1 = s_CSAwallace_cla16_csa7_csa_component_fa24_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa24_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa24_or0 = s_CSAwallace_cla16_csa7_csa_component_fa24_and0 | s_CSAwallace_cla16_csa7_csa_component_fa24_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa25_xor0 = s_CSAwallace_cla16_csa3_csa_component_fa25_xor1 ^ s_CSAwallace_cla16_csa3_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa25_and0 = s_CSAwallace_cla16_csa3_csa_component_fa25_xor1 & s_CSAwallace_cla16_csa3_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa25_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa25_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa25_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa25_and1 = s_CSAwallace_cla16_csa7_csa_component_fa25_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa25_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa25_or0 = s_CSAwallace_cla16_csa7_csa_component_fa25_and0 | s_CSAwallace_cla16_csa7_csa_component_fa25_and1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa26_xor0 = s_CSAwallace_cla16_nand_15_11 ^ s_CSAwallace_cla16_csa3_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa26_and0 = s_CSAwallace_cla16_nand_15_11 & s_CSAwallace_cla16_csa3_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa7_csa_component_fa26_xor1 = s_CSAwallace_cla16_csa7_csa_component_fa26_xor0 ^ s_CSAwallace_cla16_csa4_csa_component_fa26_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa26_and1 = s_CSAwallace_cla16_csa7_csa_component_fa26_xor0 & s_CSAwallace_cla16_csa4_csa_component_fa26_xor1;
  assign s_CSAwallace_cla16_csa7_csa_component_fa26_or0 = s_CSAwallace_cla16_csa7_csa_component_fa26_and0 | s_CSAwallace_cla16_csa7_csa_component_fa26_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa3_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa3_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa2_and0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa3_and0 = s_CSAwallace_cla16_csa5_csa_component_fa3_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa2_and0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa4_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa4_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa3_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa4_and0 = s_CSAwallace_cla16_csa5_csa_component_fa4_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa3_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa5_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa5_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa4_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa5_and0 = s_CSAwallace_cla16_csa5_csa_component_fa5_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa4_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa5_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa5_xor0 ^ s_CSAwallace_cla16_csa1_csa_component_fa4_and0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa5_and1 = s_CSAwallace_cla16_csa8_csa_component_fa5_xor0 & s_CSAwallace_cla16_csa1_csa_component_fa4_and0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa5_or0 = s_CSAwallace_cla16_csa8_csa_component_fa5_and0 | s_CSAwallace_cla16_csa8_csa_component_fa5_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa6_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa6_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa5_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa6_and0 = s_CSAwallace_cla16_csa5_csa_component_fa6_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa5_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa6_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa6_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa6_xor0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa6_and1 = s_CSAwallace_cla16_csa8_csa_component_fa6_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa6_xor0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa6_or0 = s_CSAwallace_cla16_csa8_csa_component_fa6_and0 | s_CSAwallace_cla16_csa8_csa_component_fa6_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa7_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa7_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa6_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa7_and0 = s_CSAwallace_cla16_csa5_csa_component_fa7_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa6_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa7_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa7_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa7_xor0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa7_and1 = s_CSAwallace_cla16_csa8_csa_component_fa7_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa7_xor0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa7_or0 = s_CSAwallace_cla16_csa8_csa_component_fa7_and0 | s_CSAwallace_cla16_csa8_csa_component_fa7_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa8_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa8_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa7_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa8_and0 = s_CSAwallace_cla16_csa5_csa_component_fa8_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa7_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa8_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa8_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa8_and1 = s_CSAwallace_cla16_csa8_csa_component_fa8_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa8_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa8_or0 = s_CSAwallace_cla16_csa8_csa_component_fa8_and0 | s_CSAwallace_cla16_csa8_csa_component_fa8_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa9_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa9_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa9_and0 = s_CSAwallace_cla16_csa5_csa_component_fa9_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa9_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa9_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa9_and1 = s_CSAwallace_cla16_csa8_csa_component_fa9_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa9_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa9_or0 = s_CSAwallace_cla16_csa8_csa_component_fa9_and0 | s_CSAwallace_cla16_csa8_csa_component_fa9_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa10_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa10_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa10_and0 = s_CSAwallace_cla16_csa5_csa_component_fa10_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa10_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa10_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa10_and1 = s_CSAwallace_cla16_csa8_csa_component_fa10_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa10_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa10_or0 = s_CSAwallace_cla16_csa8_csa_component_fa10_and0 | s_CSAwallace_cla16_csa8_csa_component_fa10_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa11_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa11_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa11_and0 = s_CSAwallace_cla16_csa5_csa_component_fa11_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa11_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa11_and1 = s_CSAwallace_cla16_csa8_csa_component_fa11_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa11_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa11_or0 = s_CSAwallace_cla16_csa8_csa_component_fa11_and0 | s_CSAwallace_cla16_csa8_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa12_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa12_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa12_and0 = s_CSAwallace_cla16_csa5_csa_component_fa12_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa12_and1 = s_CSAwallace_cla16_csa8_csa_component_fa12_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa12_or0 = s_CSAwallace_cla16_csa8_csa_component_fa12_and0 | s_CSAwallace_cla16_csa8_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa13_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa13_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa13_and0 = s_CSAwallace_cla16_csa5_csa_component_fa13_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa13_and1 = s_CSAwallace_cla16_csa8_csa_component_fa13_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa13_or0 = s_CSAwallace_cla16_csa8_csa_component_fa13_and0 | s_CSAwallace_cla16_csa8_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa14_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa14_and0 = s_CSAwallace_cla16_csa5_csa_component_fa14_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa14_and1 = s_CSAwallace_cla16_csa8_csa_component_fa14_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa14_or0 = s_CSAwallace_cla16_csa8_csa_component_fa14_and0 | s_CSAwallace_cla16_csa8_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa15_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa15_and0 = s_CSAwallace_cla16_csa5_csa_component_fa15_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa15_and1 = s_CSAwallace_cla16_csa8_csa_component_fa15_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa15_or0 = s_CSAwallace_cla16_csa8_csa_component_fa15_and0 | s_CSAwallace_cla16_csa8_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa16_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa16_and0 = s_CSAwallace_cla16_csa5_csa_component_fa16_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa16_and1 = s_CSAwallace_cla16_csa8_csa_component_fa16_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa16_or0 = s_CSAwallace_cla16_csa8_csa_component_fa16_and0 | s_CSAwallace_cla16_csa8_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa17_xor0 = s_CSAwallace_cla16_csa5_csa_component_fa17_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa17_and0 = s_CSAwallace_cla16_csa5_csa_component_fa17_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa17_and1 = s_CSAwallace_cla16_csa8_csa_component_fa17_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa17_or0 = s_CSAwallace_cla16_csa8_csa_component_fa17_and0 | s_CSAwallace_cla16_csa8_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa18_xor0 = s_CSAwallace_cla16_csa1_csa_component_fa18_xor1 ^ s_CSAwallace_cla16_csa5_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa18_and0 = s_CSAwallace_cla16_csa1_csa_component_fa18_xor1 & s_CSAwallace_cla16_csa5_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa8_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa18_and1 = s_CSAwallace_cla16_csa8_csa_component_fa18_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa18_or0 = s_CSAwallace_cla16_csa8_csa_component_fa18_and0 | s_CSAwallace_cla16_csa8_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa19_xor0 = ~s_CSAwallace_cla16_csa1_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa19_and1 = s_CSAwallace_cla16_csa8_csa_component_fa19_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa19_or0 = s_CSAwallace_cla16_csa1_csa_component_fa19_xor1 | s_CSAwallace_cla16_csa8_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa20_xor0 = ~s_CSAwallace_cla16_nand_15_5;
  assign s_CSAwallace_cla16_csa8_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa8_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa20_and1 = s_CSAwallace_cla16_csa8_csa_component_fa20_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa8_csa_component_fa20_or0 = s_CSAwallace_cla16_nand_15_5 | s_CSAwallace_cla16_csa8_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa9_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa8_or0 ^ s_CSAwallace_cla16_and_0_9;
  assign s_CSAwallace_cla16_csa9_csa_component_fa9_and0 = s_CSAwallace_cla16_csa6_csa_component_fa8_or0 & s_CSAwallace_cla16_and_0_9;
  assign s_CSAwallace_cla16_csa9_csa_component_fa10_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa9_or0 ^ s_CSAwallace_cla16_csa3_csa_component_fa10_xor0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa10_and0 = s_CSAwallace_cla16_csa6_csa_component_fa9_or0 & s_CSAwallace_cla16_csa3_csa_component_fa10_xor0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa11_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa10_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa11_xor0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa11_and0 = s_CSAwallace_cla16_csa6_csa_component_fa10_or0 & s_CSAwallace_cla16_csa7_csa_component_fa11_xor0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa12_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa11_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa12_and0 = s_CSAwallace_cla16_csa6_csa_component_fa11_or0 & s_CSAwallace_cla16_csa7_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa11_and0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa12_and1 = s_CSAwallace_cla16_csa9_csa_component_fa12_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa11_and0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa12_or0 = s_CSAwallace_cla16_csa9_csa_component_fa12_and0 | s_CSAwallace_cla16_csa9_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa13_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa12_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa13_and0 = s_CSAwallace_cla16_csa6_csa_component_fa12_or0 & s_CSAwallace_cla16_csa7_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa13_and1 = s_CSAwallace_cla16_csa9_csa_component_fa13_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa13_or0 = s_CSAwallace_cla16_csa9_csa_component_fa13_and0 | s_CSAwallace_cla16_csa9_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa13_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa14_and0 = s_CSAwallace_cla16_csa6_csa_component_fa13_or0 & s_CSAwallace_cla16_csa7_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa14_and1 = s_CSAwallace_cla16_csa9_csa_component_fa14_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa14_or0 = s_CSAwallace_cla16_csa9_csa_component_fa14_and0 | s_CSAwallace_cla16_csa9_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa14_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa15_and0 = s_CSAwallace_cla16_csa6_csa_component_fa14_or0 & s_CSAwallace_cla16_csa7_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa15_and1 = s_CSAwallace_cla16_csa9_csa_component_fa15_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa15_or0 = s_CSAwallace_cla16_csa9_csa_component_fa15_and0 | s_CSAwallace_cla16_csa9_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa15_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa16_and0 = s_CSAwallace_cla16_csa6_csa_component_fa15_or0 & s_CSAwallace_cla16_csa7_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa16_and1 = s_CSAwallace_cla16_csa9_csa_component_fa16_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa16_or0 = s_CSAwallace_cla16_csa9_csa_component_fa16_and0 | s_CSAwallace_cla16_csa9_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa17_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa16_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa17_and0 = s_CSAwallace_cla16_csa6_csa_component_fa16_or0 & s_CSAwallace_cla16_csa7_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa17_and1 = s_CSAwallace_cla16_csa9_csa_component_fa17_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa17_or0 = s_CSAwallace_cla16_csa9_csa_component_fa17_and0 | s_CSAwallace_cla16_csa9_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa18_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa17_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa18_and0 = s_CSAwallace_cla16_csa6_csa_component_fa17_or0 & s_CSAwallace_cla16_csa7_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa18_and1 = s_CSAwallace_cla16_csa9_csa_component_fa18_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa18_or0 = s_CSAwallace_cla16_csa9_csa_component_fa18_and0 | s_CSAwallace_cla16_csa9_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa19_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa18_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa19_and0 = s_CSAwallace_cla16_csa6_csa_component_fa18_or0 & s_CSAwallace_cla16_csa7_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa19_and1 = s_CSAwallace_cla16_csa9_csa_component_fa19_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa19_or0 = s_CSAwallace_cla16_csa9_csa_component_fa19_and0 | s_CSAwallace_cla16_csa9_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa20_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa19_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa20_and0 = s_CSAwallace_cla16_csa6_csa_component_fa19_or0 & s_CSAwallace_cla16_csa7_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa20_and1 = s_CSAwallace_cla16_csa9_csa_component_fa20_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa20_or0 = s_CSAwallace_cla16_csa9_csa_component_fa20_and0 | s_CSAwallace_cla16_csa9_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa21_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa20_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa21_and0 = s_CSAwallace_cla16_csa6_csa_component_fa20_or0 & s_CSAwallace_cla16_csa7_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa21_and1 = s_CSAwallace_cla16_csa9_csa_component_fa21_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa21_or0 = s_CSAwallace_cla16_csa9_csa_component_fa21_and0 | s_CSAwallace_cla16_csa9_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa22_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa21_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa22_and0 = s_CSAwallace_cla16_csa6_csa_component_fa21_or0 & s_CSAwallace_cla16_csa7_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa22_and1 = s_CSAwallace_cla16_csa9_csa_component_fa22_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa22_or0 = s_CSAwallace_cla16_csa9_csa_component_fa22_and0 | s_CSAwallace_cla16_csa9_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa23_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa22_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa23_and0 = s_CSAwallace_cla16_csa6_csa_component_fa22_or0 & s_CSAwallace_cla16_csa7_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa23_and1 = s_CSAwallace_cla16_csa9_csa_component_fa23_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa23_or0 = s_CSAwallace_cla16_csa9_csa_component_fa23_and0 | s_CSAwallace_cla16_csa9_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa24_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa23_or0 ^ s_CSAwallace_cla16_csa7_csa_component_fa24_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa24_and0 = s_CSAwallace_cla16_csa6_csa_component_fa23_or0 & s_CSAwallace_cla16_csa7_csa_component_fa24_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa24_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa24_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa24_and1 = s_CSAwallace_cla16_csa9_csa_component_fa24_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa24_or0 = s_CSAwallace_cla16_csa9_csa_component_fa24_and0 | s_CSAwallace_cla16_csa9_csa_component_fa24_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa25_xor0 = ~s_CSAwallace_cla16_csa7_csa_component_fa25_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa25_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa25_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa25_and1 = s_CSAwallace_cla16_csa9_csa_component_fa25_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa25_or0 = s_CSAwallace_cla16_csa7_csa_component_fa25_xor1 | s_CSAwallace_cla16_csa9_csa_component_fa25_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa26_xor0 = ~s_CSAwallace_cla16_csa7_csa_component_fa26_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa26_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa26_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa26_and1 = s_CSAwallace_cla16_csa9_csa_component_fa26_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa26_or0 = s_CSAwallace_cla16_csa7_csa_component_fa26_xor1 | s_CSAwallace_cla16_csa9_csa_component_fa26_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa27_xor0 = ~s_CSAwallace_cla16_csa4_csa_component_fa27_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa27_xor1 = s_CSAwallace_cla16_csa9_csa_component_fa27_xor0 ^ s_CSAwallace_cla16_csa7_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa27_and1 = s_CSAwallace_cla16_csa9_csa_component_fa27_xor0 & s_CSAwallace_cla16_csa7_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa27_or0 = s_CSAwallace_cla16_csa4_csa_component_fa27_xor1 | s_CSAwallace_cla16_csa9_csa_component_fa27_and1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa28_xor0 = ~s_CSAwallace_cla16_csa4_csa_component_fa28_xor1;
  assign s_CSAwallace_cla16_csa9_csa_component_fa28_xor1 = ~s_CSAwallace_cla16_csa9_csa_component_fa28_xor0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa28_or0 = s_CSAwallace_cla16_csa4_csa_component_fa28_xor1 | s_CSAwallace_cla16_csa9_csa_component_fa28_xor0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa29_xor0 = ~s_CSAwallace_cla16_nand_15_14;
  assign s_CSAwallace_cla16_csa9_csa_component_fa29_xor1 = ~s_CSAwallace_cla16_csa9_csa_component_fa29_xor0;
  assign s_CSAwallace_cla16_csa9_csa_component_fa29_or0 = s_CSAwallace_cla16_nand_15_14 | s_CSAwallace_cla16_csa9_csa_component_fa29_xor0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa4_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa4_xor0 ^ s_CSAwallace_cla16_csa8_csa_component_fa3_and0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa4_and0 = s_CSAwallace_cla16_csa8_csa_component_fa4_xor0 & s_CSAwallace_cla16_csa8_csa_component_fa3_and0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa5_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa5_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa4_and0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa5_and0 = s_CSAwallace_cla16_csa8_csa_component_fa5_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa4_and0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa6_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa6_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa5_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa6_and0 = s_CSAwallace_cla16_csa8_csa_component_fa6_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa5_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa7_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa7_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa6_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa7_and0 = s_CSAwallace_cla16_csa8_csa_component_fa7_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa6_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa7_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa7_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa7_and1 = s_CSAwallace_cla16_csa10_csa_component_fa7_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa7_or0 = s_CSAwallace_cla16_csa10_csa_component_fa7_and0 | s_CSAwallace_cla16_csa10_csa_component_fa7_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa8_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa8_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa7_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa8_and0 = s_CSAwallace_cla16_csa8_csa_component_fa8_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa7_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa8_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_csa6_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa8_and1 = s_CSAwallace_cla16_csa10_csa_component_fa8_xor0 & s_CSAwallace_cla16_csa6_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa8_or0 = s_CSAwallace_cla16_csa10_csa_component_fa8_and0 | s_CSAwallace_cla16_csa10_csa_component_fa8_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa9_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa9_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa9_and0 = s_CSAwallace_cla16_csa8_csa_component_fa9_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa9_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa9_xor0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa9_and1 = s_CSAwallace_cla16_csa10_csa_component_fa9_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa9_xor0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa9_or0 = s_CSAwallace_cla16_csa10_csa_component_fa9_and0 | s_CSAwallace_cla16_csa10_csa_component_fa9_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa10_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa10_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa10_and0 = s_CSAwallace_cla16_csa8_csa_component_fa10_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa10_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa10_xor0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa10_and1 = s_CSAwallace_cla16_csa10_csa_component_fa10_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa10_xor0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa10_or0 = s_CSAwallace_cla16_csa10_csa_component_fa10_and0 | s_CSAwallace_cla16_csa10_csa_component_fa10_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa11_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa11_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa11_and0 = s_CSAwallace_cla16_csa8_csa_component_fa11_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa11_xor0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa11_and1 = s_CSAwallace_cla16_csa10_csa_component_fa11_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa11_xor0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa11_or0 = s_CSAwallace_cla16_csa10_csa_component_fa11_and0 | s_CSAwallace_cla16_csa10_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa12_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa12_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa12_and0 = s_CSAwallace_cla16_csa8_csa_component_fa12_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa12_and1 = s_CSAwallace_cla16_csa10_csa_component_fa12_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa12_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa12_or0 = s_CSAwallace_cla16_csa10_csa_component_fa12_and0 | s_CSAwallace_cla16_csa10_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa13_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa13_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa13_and0 = s_CSAwallace_cla16_csa8_csa_component_fa13_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa13_and1 = s_CSAwallace_cla16_csa10_csa_component_fa13_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa13_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa13_or0 = s_CSAwallace_cla16_csa10_csa_component_fa13_and0 | s_CSAwallace_cla16_csa10_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa14_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa14_and0 = s_CSAwallace_cla16_csa8_csa_component_fa14_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa14_and1 = s_CSAwallace_cla16_csa10_csa_component_fa14_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa14_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa14_or0 = s_CSAwallace_cla16_csa10_csa_component_fa14_and0 | s_CSAwallace_cla16_csa10_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa15_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa15_and0 = s_CSAwallace_cla16_csa8_csa_component_fa15_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa15_and1 = s_CSAwallace_cla16_csa10_csa_component_fa15_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa15_or0 = s_CSAwallace_cla16_csa10_csa_component_fa15_and0 | s_CSAwallace_cla16_csa10_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa16_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa16_and0 = s_CSAwallace_cla16_csa8_csa_component_fa16_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa16_and1 = s_CSAwallace_cla16_csa10_csa_component_fa16_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa16_or0 = s_CSAwallace_cla16_csa10_csa_component_fa16_and0 | s_CSAwallace_cla16_csa10_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa17_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa17_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa17_and0 = s_CSAwallace_cla16_csa8_csa_component_fa17_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa17_and1 = s_CSAwallace_cla16_csa10_csa_component_fa17_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa17_or0 = s_CSAwallace_cla16_csa10_csa_component_fa17_and0 | s_CSAwallace_cla16_csa10_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa18_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa18_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa18_and0 = s_CSAwallace_cla16_csa8_csa_component_fa18_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa18_and1 = s_CSAwallace_cla16_csa10_csa_component_fa18_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa18_or0 = s_CSAwallace_cla16_csa10_csa_component_fa18_and0 | s_CSAwallace_cla16_csa10_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa19_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa19_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa19_and0 = s_CSAwallace_cla16_csa8_csa_component_fa19_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa19_and1 = s_CSAwallace_cla16_csa10_csa_component_fa19_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa19_or0 = s_CSAwallace_cla16_csa10_csa_component_fa19_and0 | s_CSAwallace_cla16_csa10_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa20_xor0 = s_CSAwallace_cla16_csa8_csa_component_fa20_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa20_and0 = s_CSAwallace_cla16_csa8_csa_component_fa20_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa20_and1 = s_CSAwallace_cla16_csa10_csa_component_fa20_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa20_or0 = s_CSAwallace_cla16_csa10_csa_component_fa20_and0 | s_CSAwallace_cla16_csa10_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa21_xor0 = s_CSAwallace_cla16_csa6_csa_component_fa21_xor1 ^ s_CSAwallace_cla16_csa8_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa21_and0 = s_CSAwallace_cla16_csa6_csa_component_fa21_xor1 & s_CSAwallace_cla16_csa8_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa10_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa21_and1 = s_CSAwallace_cla16_csa10_csa_component_fa21_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa21_or0 = s_CSAwallace_cla16_csa10_csa_component_fa21_and0 | s_CSAwallace_cla16_csa10_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa22_xor0 = ~s_CSAwallace_cla16_csa6_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa22_and1 = s_CSAwallace_cla16_csa10_csa_component_fa22_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa22_or0 = s_CSAwallace_cla16_csa6_csa_component_fa22_xor1 | s_CSAwallace_cla16_csa10_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa23_xor0 = ~s_CSAwallace_cla16_csa6_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa10_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa23_and1 = s_CSAwallace_cla16_csa10_csa_component_fa23_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa10_csa_component_fa23_or0 = s_CSAwallace_cla16_csa6_csa_component_fa23_xor1 | s_CSAwallace_cla16_csa10_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa13_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa13_and0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa14_and0 = s_CSAwallace_cla16_csa9_csa_component_fa13_or0 & s_CSAwallace_cla16_csa4_csa_component_fa13_and0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa14_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa15_and0 = s_CSAwallace_cla16_csa9_csa_component_fa14_or0 & s_CSAwallace_cla16_csa4_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_nand_0_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa15_and1 = s_CSAwallace_cla16_csa11_csa_component_fa15_xor0 & s_CSAwallace_cla16_nand_0_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa15_or0 = s_CSAwallace_cla16_csa11_csa_component_fa15_and0 | s_CSAwallace_cla16_csa11_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa15_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa16_and0 = s_CSAwallace_cla16_csa9_csa_component_fa15_or0 & s_CSAwallace_cla16_csa4_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_nand_1_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa16_and1 = s_CSAwallace_cla16_csa11_csa_component_fa16_xor0 & s_CSAwallace_cla16_nand_1_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa16_or0 = s_CSAwallace_cla16_csa11_csa_component_fa16_and0 | s_CSAwallace_cla16_csa11_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa17_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa16_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa17_and0 = s_CSAwallace_cla16_csa9_csa_component_fa16_or0 & s_CSAwallace_cla16_csa4_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_nand_2_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa17_and1 = s_CSAwallace_cla16_csa11_csa_component_fa17_xor0 & s_CSAwallace_cla16_nand_2_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa17_or0 = s_CSAwallace_cla16_csa11_csa_component_fa17_and0 | s_CSAwallace_cla16_csa11_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa18_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa17_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa18_and0 = s_CSAwallace_cla16_csa9_csa_component_fa17_or0 & s_CSAwallace_cla16_csa4_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_nand_3_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa18_and1 = s_CSAwallace_cla16_csa11_csa_component_fa18_xor0 & s_CSAwallace_cla16_nand_3_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa18_or0 = s_CSAwallace_cla16_csa11_csa_component_fa18_and0 | s_CSAwallace_cla16_csa11_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa19_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa18_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa19_and0 = s_CSAwallace_cla16_csa9_csa_component_fa18_or0 & s_CSAwallace_cla16_csa4_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_nand_4_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa19_and1 = s_CSAwallace_cla16_csa11_csa_component_fa19_xor0 & s_CSAwallace_cla16_nand_4_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa19_or0 = s_CSAwallace_cla16_csa11_csa_component_fa19_and0 | s_CSAwallace_cla16_csa11_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa20_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa19_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa20_and0 = s_CSAwallace_cla16_csa9_csa_component_fa19_or0 & s_CSAwallace_cla16_csa4_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_nand_5_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa20_and1 = s_CSAwallace_cla16_csa11_csa_component_fa20_xor0 & s_CSAwallace_cla16_nand_5_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa20_or0 = s_CSAwallace_cla16_csa11_csa_component_fa20_and0 | s_CSAwallace_cla16_csa11_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa21_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa20_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa21_and0 = s_CSAwallace_cla16_csa9_csa_component_fa20_or0 & s_CSAwallace_cla16_csa4_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_nand_6_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa21_and1 = s_CSAwallace_cla16_csa11_csa_component_fa21_xor0 & s_CSAwallace_cla16_nand_6_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa21_or0 = s_CSAwallace_cla16_csa11_csa_component_fa21_and0 | s_CSAwallace_cla16_csa11_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa22_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa21_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa22_and0 = s_CSAwallace_cla16_csa9_csa_component_fa21_or0 & s_CSAwallace_cla16_csa4_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_nand_7_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa22_and1 = s_CSAwallace_cla16_csa11_csa_component_fa22_xor0 & s_CSAwallace_cla16_nand_7_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa22_or0 = s_CSAwallace_cla16_csa11_csa_component_fa22_and0 | s_CSAwallace_cla16_csa11_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa23_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa22_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa23_and0 = s_CSAwallace_cla16_csa9_csa_component_fa22_or0 & s_CSAwallace_cla16_csa4_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_nand_8_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa23_and1 = s_CSAwallace_cla16_csa11_csa_component_fa23_xor0 & s_CSAwallace_cla16_nand_8_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa23_or0 = s_CSAwallace_cla16_csa11_csa_component_fa23_and0 | s_CSAwallace_cla16_csa11_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa24_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa23_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa24_and0 = s_CSAwallace_cla16_csa9_csa_component_fa23_or0 & s_CSAwallace_cla16_csa4_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa24_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa24_xor0 ^ s_CSAwallace_cla16_nand_9_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa24_and1 = s_CSAwallace_cla16_csa11_csa_component_fa24_xor0 & s_CSAwallace_cla16_nand_9_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa24_or0 = s_CSAwallace_cla16_csa11_csa_component_fa24_and0 | s_CSAwallace_cla16_csa11_csa_component_fa24_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa25_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa24_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa25_and0 = s_CSAwallace_cla16_csa9_csa_component_fa24_or0 & s_CSAwallace_cla16_csa4_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa25_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa25_xor0 ^ s_CSAwallace_cla16_nand_10_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa25_and1 = s_CSAwallace_cla16_csa11_csa_component_fa25_xor0 & s_CSAwallace_cla16_nand_10_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa25_or0 = s_CSAwallace_cla16_csa11_csa_component_fa25_and0 | s_CSAwallace_cla16_csa11_csa_component_fa25_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa26_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa25_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa26_and0 = s_CSAwallace_cla16_csa9_csa_component_fa25_or0 & s_CSAwallace_cla16_csa4_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa26_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa26_xor0 ^ s_CSAwallace_cla16_nand_11_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa26_and1 = s_CSAwallace_cla16_csa11_csa_component_fa26_xor0 & s_CSAwallace_cla16_nand_11_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa26_or0 = s_CSAwallace_cla16_csa11_csa_component_fa26_and0 | s_CSAwallace_cla16_csa11_csa_component_fa26_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa27_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa26_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa27_and0 = s_CSAwallace_cla16_csa9_csa_component_fa26_or0 & s_CSAwallace_cla16_csa4_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa27_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa27_xor0 ^ s_CSAwallace_cla16_nand_12_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa27_and1 = s_CSAwallace_cla16_csa11_csa_component_fa27_xor0 & s_CSAwallace_cla16_nand_12_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa27_or0 = s_CSAwallace_cla16_csa11_csa_component_fa27_and0 | s_CSAwallace_cla16_csa11_csa_component_fa27_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa28_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa27_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa28_and0 = s_CSAwallace_cla16_csa9_csa_component_fa27_or0 & s_CSAwallace_cla16_csa4_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa28_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa28_xor0 ^ s_CSAwallace_cla16_nand_13_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa28_and1 = s_CSAwallace_cla16_csa11_csa_component_fa28_xor0 & s_CSAwallace_cla16_nand_13_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa28_or0 = s_CSAwallace_cla16_csa11_csa_component_fa28_and0 | s_CSAwallace_cla16_csa11_csa_component_fa28_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa29_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa28_or0 ^ s_CSAwallace_cla16_csa4_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa29_and0 = s_CSAwallace_cla16_csa9_csa_component_fa28_or0 & s_CSAwallace_cla16_csa4_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa29_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa29_xor0 ^ s_CSAwallace_cla16_nand_14_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa29_and1 = s_CSAwallace_cla16_csa11_csa_component_fa29_xor0 & s_CSAwallace_cla16_nand_14_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa29_or0 = s_CSAwallace_cla16_csa11_csa_component_fa29_and0 | s_CSAwallace_cla16_csa11_csa_component_fa29_and1;
  assign s_CSAwallace_cla16_csa11_csa_component_fa30_xor0 = ~s_CSAwallace_cla16_csa9_csa_component_fa29_or0;
  assign s_CSAwallace_cla16_csa11_csa_component_fa30_xor1 = s_CSAwallace_cla16_csa11_csa_component_fa30_xor0 ^ s_CSAwallace_cla16_and_15_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa30_and1 = s_CSAwallace_cla16_csa11_csa_component_fa30_xor0 & s_CSAwallace_cla16_and_15_15;
  assign s_CSAwallace_cla16_csa11_csa_component_fa30_or0 = s_CSAwallace_cla16_csa9_csa_component_fa29_or0 | s_CSAwallace_cla16_csa11_csa_component_fa30_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa5_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa5_xor0 ^ s_CSAwallace_cla16_csa10_csa_component_fa4_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa5_and0 = s_CSAwallace_cla16_csa10_csa_component_fa5_xor0 & s_CSAwallace_cla16_csa10_csa_component_fa4_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa6_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa6_xor0 ^ s_CSAwallace_cla16_csa10_csa_component_fa5_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa6_and0 = s_CSAwallace_cla16_csa10_csa_component_fa6_xor0 & s_CSAwallace_cla16_csa10_csa_component_fa5_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa7_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa7_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa7_and0 = s_CSAwallace_cla16_csa10_csa_component_fa7_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa8_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa8_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa7_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa8_and0 = s_CSAwallace_cla16_csa10_csa_component_fa8_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa7_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa9_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa9_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa9_and0 = s_CSAwallace_cla16_csa10_csa_component_fa9_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa8_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa10_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa10_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa10_and0 = s_CSAwallace_cla16_csa10_csa_component_fa10_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa9_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa10_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa9_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa10_and1 = s_CSAwallace_cla16_csa12_csa_component_fa10_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa9_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa10_or0 = s_CSAwallace_cla16_csa12_csa_component_fa10_and0 | s_CSAwallace_cla16_csa12_csa_component_fa10_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa11_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa11_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa11_and0 = s_CSAwallace_cla16_csa10_csa_component_fa11_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa11_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa10_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa11_and1 = s_CSAwallace_cla16_csa12_csa_component_fa11_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa10_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa11_or0 = s_CSAwallace_cla16_csa12_csa_component_fa11_and0 | s_CSAwallace_cla16_csa12_csa_component_fa11_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa12_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa12_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa12_and0 = s_CSAwallace_cla16_csa10_csa_component_fa12_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa12_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa11_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa12_and1 = s_CSAwallace_cla16_csa12_csa_component_fa12_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa11_and0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa12_or0 = s_CSAwallace_cla16_csa12_csa_component_fa12_and0 | s_CSAwallace_cla16_csa12_csa_component_fa12_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa13_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa13_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa13_and0 = s_CSAwallace_cla16_csa10_csa_component_fa13_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa13_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_csa9_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa13_and1 = s_CSAwallace_cla16_csa12_csa_component_fa13_xor0 & s_CSAwallace_cla16_csa9_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa13_or0 = s_CSAwallace_cla16_csa12_csa_component_fa13_and0 | s_CSAwallace_cla16_csa12_csa_component_fa13_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa14_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa14_and0 = s_CSAwallace_cla16_csa10_csa_component_fa14_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa14_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa14_xor0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa14_and1 = s_CSAwallace_cla16_csa12_csa_component_fa14_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa14_xor0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa14_or0 = s_CSAwallace_cla16_csa12_csa_component_fa14_and0 | s_CSAwallace_cla16_csa12_csa_component_fa14_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa15_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa15_and0 = s_CSAwallace_cla16_csa10_csa_component_fa15_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa15_and1 = s_CSAwallace_cla16_csa12_csa_component_fa15_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa15_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa15_or0 = s_CSAwallace_cla16_csa12_csa_component_fa15_and0 | s_CSAwallace_cla16_csa12_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa16_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa16_and0 = s_CSAwallace_cla16_csa10_csa_component_fa16_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa16_and1 = s_CSAwallace_cla16_csa12_csa_component_fa16_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa16_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa16_or0 = s_CSAwallace_cla16_csa12_csa_component_fa16_and0 | s_CSAwallace_cla16_csa12_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa17_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa17_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa17_and0 = s_CSAwallace_cla16_csa10_csa_component_fa17_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa17_and1 = s_CSAwallace_cla16_csa12_csa_component_fa17_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa17_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa17_or0 = s_CSAwallace_cla16_csa12_csa_component_fa17_and0 | s_CSAwallace_cla16_csa12_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa18_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa18_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa18_and0 = s_CSAwallace_cla16_csa10_csa_component_fa18_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa18_and1 = s_CSAwallace_cla16_csa12_csa_component_fa18_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa18_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa18_or0 = s_CSAwallace_cla16_csa12_csa_component_fa18_and0 | s_CSAwallace_cla16_csa12_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa19_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa19_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa19_and0 = s_CSAwallace_cla16_csa10_csa_component_fa19_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa19_and1 = s_CSAwallace_cla16_csa12_csa_component_fa19_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa19_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa19_or0 = s_CSAwallace_cla16_csa12_csa_component_fa19_and0 | s_CSAwallace_cla16_csa12_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa20_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa20_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa20_and0 = s_CSAwallace_cla16_csa10_csa_component_fa20_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa20_and1 = s_CSAwallace_cla16_csa12_csa_component_fa20_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa20_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa20_or0 = s_CSAwallace_cla16_csa12_csa_component_fa20_and0 | s_CSAwallace_cla16_csa12_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa21_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa21_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa21_and0 = s_CSAwallace_cla16_csa10_csa_component_fa21_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa21_and1 = s_CSAwallace_cla16_csa12_csa_component_fa21_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa21_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa21_or0 = s_CSAwallace_cla16_csa12_csa_component_fa21_and0 | s_CSAwallace_cla16_csa12_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa22_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa22_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa22_and0 = s_CSAwallace_cla16_csa10_csa_component_fa22_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa22_and1 = s_CSAwallace_cla16_csa12_csa_component_fa22_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa22_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa22_or0 = s_CSAwallace_cla16_csa12_csa_component_fa22_and0 | s_CSAwallace_cla16_csa12_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa23_xor0 = s_CSAwallace_cla16_csa10_csa_component_fa23_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa23_and0 = s_CSAwallace_cla16_csa10_csa_component_fa23_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa23_and1 = s_CSAwallace_cla16_csa12_csa_component_fa23_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa23_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa23_or0 = s_CSAwallace_cla16_csa12_csa_component_fa23_and0 | s_CSAwallace_cla16_csa12_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa24_xor0 = s_CSAwallace_cla16_csa9_csa_component_fa24_xor1 ^ s_CSAwallace_cla16_csa10_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa24_and0 = s_CSAwallace_cla16_csa9_csa_component_fa24_xor1 & s_CSAwallace_cla16_csa10_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa12_csa_component_fa24_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa24_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa24_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa24_and1 = s_CSAwallace_cla16_csa12_csa_component_fa24_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa24_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa24_or0 = s_CSAwallace_cla16_csa12_csa_component_fa24_and0 | s_CSAwallace_cla16_csa12_csa_component_fa24_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa25_xor0 = ~s_CSAwallace_cla16_csa9_csa_component_fa25_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa25_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa25_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa25_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa25_and1 = s_CSAwallace_cla16_csa12_csa_component_fa25_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa25_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa25_or0 = s_CSAwallace_cla16_csa9_csa_component_fa25_xor1 | s_CSAwallace_cla16_csa12_csa_component_fa25_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa26_xor0 = ~s_CSAwallace_cla16_csa9_csa_component_fa26_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa26_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa26_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa26_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa26_and1 = s_CSAwallace_cla16_csa12_csa_component_fa26_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa26_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa26_or0 = s_CSAwallace_cla16_csa9_csa_component_fa26_xor1 | s_CSAwallace_cla16_csa12_csa_component_fa26_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa27_xor0 = ~s_CSAwallace_cla16_csa9_csa_component_fa27_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa27_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa27_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa27_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa27_and1 = s_CSAwallace_cla16_csa12_csa_component_fa27_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa27_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa27_or0 = s_CSAwallace_cla16_csa9_csa_component_fa27_xor1 | s_CSAwallace_cla16_csa12_csa_component_fa27_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa28_xor0 = ~s_CSAwallace_cla16_csa9_csa_component_fa28_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa28_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa28_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa28_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa28_and1 = s_CSAwallace_cla16_csa12_csa_component_fa28_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa28_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa28_or0 = s_CSAwallace_cla16_csa9_csa_component_fa28_xor1 | s_CSAwallace_cla16_csa12_csa_component_fa28_and1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa29_xor0 = ~s_CSAwallace_cla16_csa9_csa_component_fa29_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa29_xor1 = s_CSAwallace_cla16_csa12_csa_component_fa29_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa29_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa29_and1 = s_CSAwallace_cla16_csa12_csa_component_fa29_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa29_xor1;
  assign s_CSAwallace_cla16_csa12_csa_component_fa29_or0 = s_CSAwallace_cla16_csa9_csa_component_fa29_xor1 | s_CSAwallace_cla16_csa12_csa_component_fa29_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa6_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa6_xor0 ^ s_CSAwallace_cla16_csa12_csa_component_fa5_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa6_and0 = s_CSAwallace_cla16_csa12_csa_component_fa6_xor0 & s_CSAwallace_cla16_csa12_csa_component_fa5_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa7_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa7_xor0 ^ s_CSAwallace_cla16_csa12_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa7_and0 = s_CSAwallace_cla16_csa12_csa_component_fa7_xor0 & s_CSAwallace_cla16_csa12_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa8_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_csa12_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa8_and0 = s_CSAwallace_cla16_csa12_csa_component_fa8_xor0 & s_CSAwallace_cla16_csa12_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa9_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_csa12_csa_component_fa8_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa9_and0 = s_CSAwallace_cla16_csa12_csa_component_fa9_xor0 & s_CSAwallace_cla16_csa12_csa_component_fa8_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa10_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa10_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa9_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa10_and0 = s_CSAwallace_cla16_csa12_csa_component_fa10_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa9_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa11_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa11_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa11_and0 = s_CSAwallace_cla16_csa12_csa_component_fa11_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa10_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa12_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa12_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa12_and0 = s_CSAwallace_cla16_csa12_csa_component_fa12_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa11_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa13_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa13_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa13_and0 = s_CSAwallace_cla16_csa12_csa_component_fa13_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa12_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa14_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa14_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa14_and0 = s_CSAwallace_cla16_csa12_csa_component_fa14_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa13_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa15_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa15_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa15_and0 = s_CSAwallace_cla16_csa12_csa_component_fa15_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa14_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa15_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa15_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa14_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa15_and1 = s_CSAwallace_cla16_csa13_csa_component_fa15_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa14_and0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa15_or0 = s_CSAwallace_cla16_csa13_csa_component_fa15_and0 | s_CSAwallace_cla16_csa13_csa_component_fa15_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa16_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa16_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa16_and0 = s_CSAwallace_cla16_csa12_csa_component_fa16_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa16_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa16_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa16_and1 = s_CSAwallace_cla16_csa13_csa_component_fa16_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa16_or0 = s_CSAwallace_cla16_csa13_csa_component_fa16_and0 | s_CSAwallace_cla16_csa13_csa_component_fa16_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa17_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa17_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa17_and0 = s_CSAwallace_cla16_csa12_csa_component_fa17_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa17_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa17_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa17_and1 = s_CSAwallace_cla16_csa13_csa_component_fa17_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa17_or0 = s_CSAwallace_cla16_csa13_csa_component_fa17_and0 | s_CSAwallace_cla16_csa13_csa_component_fa17_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa18_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa18_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa18_and0 = s_CSAwallace_cla16_csa12_csa_component_fa18_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa18_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa18_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa18_and1 = s_CSAwallace_cla16_csa13_csa_component_fa18_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa18_or0 = s_CSAwallace_cla16_csa13_csa_component_fa18_and0 | s_CSAwallace_cla16_csa13_csa_component_fa18_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa19_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa19_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa19_and0 = s_CSAwallace_cla16_csa12_csa_component_fa19_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa19_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa19_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa19_and1 = s_CSAwallace_cla16_csa13_csa_component_fa19_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa19_or0 = s_CSAwallace_cla16_csa13_csa_component_fa19_and0 | s_CSAwallace_cla16_csa13_csa_component_fa19_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa20_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa20_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa20_and0 = s_CSAwallace_cla16_csa12_csa_component_fa20_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa20_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa20_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa20_and1 = s_CSAwallace_cla16_csa13_csa_component_fa20_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa20_or0 = s_CSAwallace_cla16_csa13_csa_component_fa20_and0 | s_CSAwallace_cla16_csa13_csa_component_fa20_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa21_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa21_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa21_and0 = s_CSAwallace_cla16_csa12_csa_component_fa21_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa21_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa21_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa21_and1 = s_CSAwallace_cla16_csa13_csa_component_fa21_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa21_or0 = s_CSAwallace_cla16_csa13_csa_component_fa21_and0 | s_CSAwallace_cla16_csa13_csa_component_fa21_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa22_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa22_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa22_and0 = s_CSAwallace_cla16_csa12_csa_component_fa22_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa22_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa22_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa22_and1 = s_CSAwallace_cla16_csa13_csa_component_fa22_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa22_or0 = s_CSAwallace_cla16_csa13_csa_component_fa22_and0 | s_CSAwallace_cla16_csa13_csa_component_fa22_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa23_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa23_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa23_and0 = s_CSAwallace_cla16_csa12_csa_component_fa23_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa23_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa23_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa23_and1 = s_CSAwallace_cla16_csa13_csa_component_fa23_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa23_or0 = s_CSAwallace_cla16_csa13_csa_component_fa23_and0 | s_CSAwallace_cla16_csa13_csa_component_fa23_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa24_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa24_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa24_and0 = s_CSAwallace_cla16_csa12_csa_component_fa24_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa24_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa24_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa24_and1 = s_CSAwallace_cla16_csa13_csa_component_fa24_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa24_or0 = s_CSAwallace_cla16_csa13_csa_component_fa24_and0 | s_CSAwallace_cla16_csa13_csa_component_fa24_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa25_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa25_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa25_and0 = s_CSAwallace_cla16_csa12_csa_component_fa25_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa25_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa25_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa25_and1 = s_CSAwallace_cla16_csa13_csa_component_fa25_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa25_or0 = s_CSAwallace_cla16_csa13_csa_component_fa25_and0 | s_CSAwallace_cla16_csa13_csa_component_fa25_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa26_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa26_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa26_and0 = s_CSAwallace_cla16_csa12_csa_component_fa26_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa26_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa26_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa26_and1 = s_CSAwallace_cla16_csa13_csa_component_fa26_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa26_or0 = s_CSAwallace_cla16_csa13_csa_component_fa26_and0 | s_CSAwallace_cla16_csa13_csa_component_fa26_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa27_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa27_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa27_and0 = s_CSAwallace_cla16_csa12_csa_component_fa27_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa27_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa27_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa27_and1 = s_CSAwallace_cla16_csa13_csa_component_fa27_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa27_or0 = s_CSAwallace_cla16_csa13_csa_component_fa27_and0 | s_CSAwallace_cla16_csa13_csa_component_fa27_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa28_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa28_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa28_and0 = s_CSAwallace_cla16_csa12_csa_component_fa28_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa28_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa28_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa28_and1 = s_CSAwallace_cla16_csa13_csa_component_fa28_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa28_or0 = s_CSAwallace_cla16_csa13_csa_component_fa28_and0 | s_CSAwallace_cla16_csa13_csa_component_fa28_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa29_xor0 = s_CSAwallace_cla16_csa12_csa_component_fa29_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa29_and0 = s_CSAwallace_cla16_csa12_csa_component_fa29_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa29_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa29_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa29_and1 = s_CSAwallace_cla16_csa13_csa_component_fa29_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa29_or0 = s_CSAwallace_cla16_csa13_csa_component_fa29_and0 | s_CSAwallace_cla16_csa13_csa_component_fa29_and1;
  assign s_CSAwallace_cla16_csa13_csa_component_fa30_xor0 = s_CSAwallace_cla16_csa11_csa_component_fa30_xor1 ^ s_CSAwallace_cla16_csa12_csa_component_fa29_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa30_and0 = s_CSAwallace_cla16_csa11_csa_component_fa30_xor1 & s_CSAwallace_cla16_csa12_csa_component_fa29_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa30_xor1 = s_CSAwallace_cla16_csa13_csa_component_fa30_xor0 ^ s_CSAwallace_cla16_csa11_csa_component_fa29_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa30_and1 = s_CSAwallace_cla16_csa13_csa_component_fa30_xor0 & s_CSAwallace_cla16_csa11_csa_component_fa29_or0;
  assign s_CSAwallace_cla16_csa13_csa_component_fa30_or0 = s_CSAwallace_cla16_csa13_csa_component_fa30_and0 | s_CSAwallace_cla16_csa13_csa_component_fa30_and1;
  assign s_CSAwallace_cla16_u_cla32_and0 = s_CSAwallace_cla16_csa5_csa_component_fa2_xor0 & s_CSAwallace_cla16_and_0_0;
  assign s_CSAwallace_cla16_u_cla32_and1 = s_CSAwallace_cla16_csa8_csa_component_fa3_xor0 & s_CSAwallace_cla16_csa0_csa_component_fa1_xor0;
  assign s_CSAwallace_cla16_u_cla32_and2 = s_CSAwallace_cla16_csa8_csa_component_fa3_xor0 & s_CSAwallace_cla16_csa0_csa_component_fa1_xor0;
  assign s_CSAwallace_cla16_u_cla32_and3 = s_CSAwallace_cla16_csa13_csa_component_fa6_xor0 & s_CSAwallace_cla16_csa10_csa_component_fa4_xor0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic7_or0 = s_CSAwallace_cla16_csa13_csa_component_fa7_xor0 | s_CSAwallace_cla16_csa13_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic7_and0 = s_CSAwallace_cla16_csa13_csa_component_fa7_xor0 & s_CSAwallace_cla16_csa13_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic7_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa7_xor0 ^ s_CSAwallace_cla16_csa13_csa_component_fa6_and0;
  assign s_CSAwallace_cla16_u_cla32_and4 = s_CSAwallace_cla16_u_cla32_pg_logic7_or0 & s_CSAwallace_cla16_csa12_csa_component_fa5_xor0;
  assign s_CSAwallace_cla16_u_cla32_and5 = s_CSAwallace_cla16_u_cla32_pg_logic7_or0 & s_CSAwallace_cla16_csa12_csa_component_fa5_xor0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic8_or0 = s_CSAwallace_cla16_csa13_csa_component_fa8_xor0 | s_CSAwallace_cla16_csa13_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic8_and0 = s_CSAwallace_cla16_csa13_csa_component_fa8_xor0 & s_CSAwallace_cla16_csa13_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic8_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa8_xor0 ^ s_CSAwallace_cla16_csa13_csa_component_fa7_and0;
  assign s_CSAwallace_cla16_u_cla32_xor8 = s_CSAwallace_cla16_u_cla32_pg_logic8_xor0 ^ s_CSAwallace_cla16_u_cla32_pg_logic7_and0;
  assign s_CSAwallace_cla16_u_cla32_and6 = s_CSAwallace_cla16_u_cla32_pg_logic7_and0 & s_CSAwallace_cla16_u_cla32_pg_logic8_or0;
  assign s_CSAwallace_cla16_u_cla32_or0 = s_CSAwallace_cla16_u_cla32_pg_logic8_and0 | s_CSAwallace_cla16_u_cla32_and6;
  assign s_CSAwallace_cla16_u_cla32_pg_logic9_or0 = s_CSAwallace_cla16_csa13_csa_component_fa9_xor0 | s_CSAwallace_cla16_csa13_csa_component_fa8_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic9_and0 = s_CSAwallace_cla16_csa13_csa_component_fa9_xor0 & s_CSAwallace_cla16_csa13_csa_component_fa8_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic9_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa9_xor0 ^ s_CSAwallace_cla16_csa13_csa_component_fa8_and0;
  assign s_CSAwallace_cla16_u_cla32_xor9 = s_CSAwallace_cla16_u_cla32_pg_logic9_xor0 ^ s_CSAwallace_cla16_u_cla32_or0;
  assign s_CSAwallace_cla16_u_cla32_and7 = s_CSAwallace_cla16_u_cla32_pg_logic7_and0 & s_CSAwallace_cla16_u_cla32_pg_logic9_or0;
  assign s_CSAwallace_cla16_u_cla32_and8 = s_CSAwallace_cla16_u_cla32_and7 & s_CSAwallace_cla16_u_cla32_pg_logic8_or0;
  assign s_CSAwallace_cla16_u_cla32_and9 = s_CSAwallace_cla16_u_cla32_pg_logic8_and0 & s_CSAwallace_cla16_u_cla32_pg_logic9_or0;
  assign s_CSAwallace_cla16_u_cla32_or1 = s_CSAwallace_cla16_u_cla32_and8 | s_CSAwallace_cla16_u_cla32_and9;
  assign s_CSAwallace_cla16_u_cla32_or2 = s_CSAwallace_cla16_u_cla32_pg_logic9_and0 | s_CSAwallace_cla16_u_cla32_or1;
  assign s_CSAwallace_cla16_u_cla32_pg_logic10_or0 = s_CSAwallace_cla16_csa13_csa_component_fa10_xor0 | s_CSAwallace_cla16_csa13_csa_component_fa9_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic10_and0 = s_CSAwallace_cla16_csa13_csa_component_fa10_xor0 & s_CSAwallace_cla16_csa13_csa_component_fa9_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic10_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa10_xor0 ^ s_CSAwallace_cla16_csa13_csa_component_fa9_and0;
  assign s_CSAwallace_cla16_u_cla32_xor10 = s_CSAwallace_cla16_u_cla32_pg_logic10_xor0 ^ s_CSAwallace_cla16_u_cla32_or2;
  assign s_CSAwallace_cla16_u_cla32_and10 = s_CSAwallace_cla16_u_cla32_pg_logic7_and0 & s_CSAwallace_cla16_u_cla32_pg_logic9_or0;
  assign s_CSAwallace_cla16_u_cla32_and11 = s_CSAwallace_cla16_u_cla32_pg_logic10_or0 & s_CSAwallace_cla16_u_cla32_pg_logic8_or0;
  assign s_CSAwallace_cla16_u_cla32_and12 = s_CSAwallace_cla16_u_cla32_and10 & s_CSAwallace_cla16_u_cla32_and11;
  assign s_CSAwallace_cla16_u_cla32_and13 = s_CSAwallace_cla16_u_cla32_pg_logic8_and0 & s_CSAwallace_cla16_u_cla32_pg_logic10_or0;
  assign s_CSAwallace_cla16_u_cla32_and14 = s_CSAwallace_cla16_u_cla32_and13 & s_CSAwallace_cla16_u_cla32_pg_logic9_or0;
  assign s_CSAwallace_cla16_u_cla32_and15 = s_CSAwallace_cla16_u_cla32_pg_logic9_and0 & s_CSAwallace_cla16_u_cla32_pg_logic10_or0;
  assign s_CSAwallace_cla16_u_cla32_or3 = s_CSAwallace_cla16_u_cla32_and12 | s_CSAwallace_cla16_u_cla32_and14;
  assign s_CSAwallace_cla16_u_cla32_or4 = s_CSAwallace_cla16_u_cla32_or3 | s_CSAwallace_cla16_u_cla32_and15;
  assign s_CSAwallace_cla16_u_cla32_or5 = s_CSAwallace_cla16_u_cla32_pg_logic10_and0 | s_CSAwallace_cla16_u_cla32_or4;
  assign s_CSAwallace_cla16_u_cla32_pg_logic11_or0 = s_CSAwallace_cla16_csa13_csa_component_fa11_xor0 | s_CSAwallace_cla16_csa13_csa_component_fa10_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic11_and0 = s_CSAwallace_cla16_csa13_csa_component_fa11_xor0 & s_CSAwallace_cla16_csa13_csa_component_fa10_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic11_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa11_xor0 ^ s_CSAwallace_cla16_csa13_csa_component_fa10_and0;
  assign s_CSAwallace_cla16_u_cla32_xor11 = s_CSAwallace_cla16_u_cla32_pg_logic11_xor0 ^ s_CSAwallace_cla16_u_cla32_or5;
  assign s_CSAwallace_cla16_u_cla32_and16 = s_CSAwallace_cla16_u_cla32_pg_logic7_and0 & s_CSAwallace_cla16_u_cla32_pg_logic10_or0;
  assign s_CSAwallace_cla16_u_cla32_and17 = s_CSAwallace_cla16_u_cla32_pg_logic11_or0 & s_CSAwallace_cla16_u_cla32_pg_logic9_or0;
  assign s_CSAwallace_cla16_u_cla32_and18 = s_CSAwallace_cla16_u_cla32_and16 & s_CSAwallace_cla16_u_cla32_and17;
  assign s_CSAwallace_cla16_u_cla32_and19 = s_CSAwallace_cla16_u_cla32_and18 & s_CSAwallace_cla16_u_cla32_pg_logic8_or0;
  assign s_CSAwallace_cla16_u_cla32_and20 = s_CSAwallace_cla16_u_cla32_pg_logic8_and0 & s_CSAwallace_cla16_u_cla32_pg_logic10_or0;
  assign s_CSAwallace_cla16_u_cla32_and21 = s_CSAwallace_cla16_u_cla32_pg_logic11_or0 & s_CSAwallace_cla16_u_cla32_pg_logic9_or0;
  assign s_CSAwallace_cla16_u_cla32_and22 = s_CSAwallace_cla16_u_cla32_and20 & s_CSAwallace_cla16_u_cla32_and21;
  assign s_CSAwallace_cla16_u_cla32_and23 = s_CSAwallace_cla16_u_cla32_pg_logic9_and0 & s_CSAwallace_cla16_u_cla32_pg_logic11_or0;
  assign s_CSAwallace_cla16_u_cla32_and24 = s_CSAwallace_cla16_u_cla32_and23 & s_CSAwallace_cla16_u_cla32_pg_logic10_or0;
  assign s_CSAwallace_cla16_u_cla32_and25 = s_CSAwallace_cla16_u_cla32_pg_logic10_and0 & s_CSAwallace_cla16_u_cla32_pg_logic11_or0;
  assign s_CSAwallace_cla16_u_cla32_or6 = s_CSAwallace_cla16_u_cla32_and19 | s_CSAwallace_cla16_u_cla32_and24;
  assign s_CSAwallace_cla16_u_cla32_or7 = s_CSAwallace_cla16_u_cla32_and22 | s_CSAwallace_cla16_u_cla32_and25;
  assign s_CSAwallace_cla16_u_cla32_or8 = s_CSAwallace_cla16_u_cla32_or6 | s_CSAwallace_cla16_u_cla32_or7;
  assign s_CSAwallace_cla16_u_cla32_or9 = s_CSAwallace_cla16_u_cla32_pg_logic11_and0 | s_CSAwallace_cla16_u_cla32_or8;
  assign s_CSAwallace_cla16_u_cla32_pg_logic12_or0 = s_CSAwallace_cla16_csa13_csa_component_fa12_xor0 | s_CSAwallace_cla16_csa13_csa_component_fa11_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic12_and0 = s_CSAwallace_cla16_csa13_csa_component_fa12_xor0 & s_CSAwallace_cla16_csa13_csa_component_fa11_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic12_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa12_xor0 ^ s_CSAwallace_cla16_csa13_csa_component_fa11_and0;
  assign s_CSAwallace_cla16_u_cla32_xor12 = s_CSAwallace_cla16_u_cla32_pg_logic12_xor0 ^ s_CSAwallace_cla16_u_cla32_or9;
  assign s_CSAwallace_cla16_u_cla32_and26 = s_CSAwallace_cla16_u_cla32_or9 & s_CSAwallace_cla16_u_cla32_pg_logic12_or0;
  assign s_CSAwallace_cla16_u_cla32_or10 = s_CSAwallace_cla16_u_cla32_pg_logic12_and0 | s_CSAwallace_cla16_u_cla32_and26;
  assign s_CSAwallace_cla16_u_cla32_pg_logic13_or0 = s_CSAwallace_cla16_csa13_csa_component_fa13_xor0 | s_CSAwallace_cla16_csa13_csa_component_fa12_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic13_and0 = s_CSAwallace_cla16_csa13_csa_component_fa13_xor0 & s_CSAwallace_cla16_csa13_csa_component_fa12_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic13_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa13_xor0 ^ s_CSAwallace_cla16_csa13_csa_component_fa12_and0;
  assign s_CSAwallace_cla16_u_cla32_xor13 = s_CSAwallace_cla16_u_cla32_pg_logic13_xor0 ^ s_CSAwallace_cla16_u_cla32_or10;
  assign s_CSAwallace_cla16_u_cla32_and27 = s_CSAwallace_cla16_u_cla32_or9 & s_CSAwallace_cla16_u_cla32_pg_logic13_or0;
  assign s_CSAwallace_cla16_u_cla32_and28 = s_CSAwallace_cla16_u_cla32_and27 & s_CSAwallace_cla16_u_cla32_pg_logic12_or0;
  assign s_CSAwallace_cla16_u_cla32_and29 = s_CSAwallace_cla16_u_cla32_pg_logic12_and0 & s_CSAwallace_cla16_u_cla32_pg_logic13_or0;
  assign s_CSAwallace_cla16_u_cla32_or11 = s_CSAwallace_cla16_u_cla32_and28 | s_CSAwallace_cla16_u_cla32_and29;
  assign s_CSAwallace_cla16_u_cla32_or12 = s_CSAwallace_cla16_u_cla32_pg_logic13_and0 | s_CSAwallace_cla16_u_cla32_or11;
  assign s_CSAwallace_cla16_u_cla32_pg_logic14_or0 = s_CSAwallace_cla16_csa13_csa_component_fa14_xor0 | s_CSAwallace_cla16_csa13_csa_component_fa13_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic14_and0 = s_CSAwallace_cla16_csa13_csa_component_fa14_xor0 & s_CSAwallace_cla16_csa13_csa_component_fa13_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic14_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa14_xor0 ^ s_CSAwallace_cla16_csa13_csa_component_fa13_and0;
  assign s_CSAwallace_cla16_u_cla32_xor14 = s_CSAwallace_cla16_u_cla32_pg_logic14_xor0 ^ s_CSAwallace_cla16_u_cla32_or12;
  assign s_CSAwallace_cla16_u_cla32_and30 = s_CSAwallace_cla16_u_cla32_or9 & s_CSAwallace_cla16_u_cla32_pg_logic13_or0;
  assign s_CSAwallace_cla16_u_cla32_and31 = s_CSAwallace_cla16_u_cla32_pg_logic14_or0 & s_CSAwallace_cla16_u_cla32_pg_logic12_or0;
  assign s_CSAwallace_cla16_u_cla32_and32 = s_CSAwallace_cla16_u_cla32_and30 & s_CSAwallace_cla16_u_cla32_and31;
  assign s_CSAwallace_cla16_u_cla32_and33 = s_CSAwallace_cla16_u_cla32_pg_logic12_and0 & s_CSAwallace_cla16_u_cla32_pg_logic14_or0;
  assign s_CSAwallace_cla16_u_cla32_and34 = s_CSAwallace_cla16_u_cla32_and33 & s_CSAwallace_cla16_u_cla32_pg_logic13_or0;
  assign s_CSAwallace_cla16_u_cla32_and35 = s_CSAwallace_cla16_u_cla32_pg_logic13_and0 & s_CSAwallace_cla16_u_cla32_pg_logic14_or0;
  assign s_CSAwallace_cla16_u_cla32_or13 = s_CSAwallace_cla16_u_cla32_and32 | s_CSAwallace_cla16_u_cla32_and34;
  assign s_CSAwallace_cla16_u_cla32_or14 = s_CSAwallace_cla16_u_cla32_or13 | s_CSAwallace_cla16_u_cla32_and35;
  assign s_CSAwallace_cla16_u_cla32_or15 = s_CSAwallace_cla16_u_cla32_pg_logic14_and0 | s_CSAwallace_cla16_u_cla32_or14;
  assign s_CSAwallace_cla16_u_cla32_pg_logic15_or0 = s_CSAwallace_cla16_csa13_csa_component_fa15_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa14_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic15_and0 = s_CSAwallace_cla16_csa13_csa_component_fa15_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa14_and0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic15_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa15_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa14_and0;
  assign s_CSAwallace_cla16_u_cla32_xor15 = s_CSAwallace_cla16_u_cla32_pg_logic15_xor0 ^ s_CSAwallace_cla16_u_cla32_or15;
  assign s_CSAwallace_cla16_u_cla32_and36 = s_CSAwallace_cla16_u_cla32_or9 & s_CSAwallace_cla16_u_cla32_pg_logic14_or0;
  assign s_CSAwallace_cla16_u_cla32_and37 = s_CSAwallace_cla16_u_cla32_pg_logic15_or0 & s_CSAwallace_cla16_u_cla32_pg_logic13_or0;
  assign s_CSAwallace_cla16_u_cla32_and38 = s_CSAwallace_cla16_u_cla32_and36 & s_CSAwallace_cla16_u_cla32_and37;
  assign s_CSAwallace_cla16_u_cla32_and39 = s_CSAwallace_cla16_u_cla32_and38 & s_CSAwallace_cla16_u_cla32_pg_logic12_or0;
  assign s_CSAwallace_cla16_u_cla32_and40 = s_CSAwallace_cla16_u_cla32_pg_logic12_and0 & s_CSAwallace_cla16_u_cla32_pg_logic14_or0;
  assign s_CSAwallace_cla16_u_cla32_and41 = s_CSAwallace_cla16_u_cla32_pg_logic15_or0 & s_CSAwallace_cla16_u_cla32_pg_logic13_or0;
  assign s_CSAwallace_cla16_u_cla32_and42 = s_CSAwallace_cla16_u_cla32_and40 & s_CSAwallace_cla16_u_cla32_and41;
  assign s_CSAwallace_cla16_u_cla32_and43 = s_CSAwallace_cla16_u_cla32_pg_logic13_and0 & s_CSAwallace_cla16_u_cla32_pg_logic15_or0;
  assign s_CSAwallace_cla16_u_cla32_and44 = s_CSAwallace_cla16_u_cla32_and43 & s_CSAwallace_cla16_u_cla32_pg_logic14_or0;
  assign s_CSAwallace_cla16_u_cla32_and45 = s_CSAwallace_cla16_u_cla32_pg_logic14_and0 & s_CSAwallace_cla16_u_cla32_pg_logic15_or0;
  assign s_CSAwallace_cla16_u_cla32_or16 = s_CSAwallace_cla16_u_cla32_and39 | s_CSAwallace_cla16_u_cla32_and44;
  assign s_CSAwallace_cla16_u_cla32_or17 = s_CSAwallace_cla16_u_cla32_and42 | s_CSAwallace_cla16_u_cla32_and45;
  assign s_CSAwallace_cla16_u_cla32_or18 = s_CSAwallace_cla16_u_cla32_or16 | s_CSAwallace_cla16_u_cla32_or17;
  assign s_CSAwallace_cla16_u_cla32_or19 = s_CSAwallace_cla16_u_cla32_pg_logic15_and0 | s_CSAwallace_cla16_u_cla32_or18;
  assign s_CSAwallace_cla16_u_cla32_pg_logic16_or0 = s_CSAwallace_cla16_csa13_csa_component_fa16_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic16_and0 = s_CSAwallace_cla16_csa13_csa_component_fa16_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic16_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa16_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa15_or0;
  assign s_CSAwallace_cla16_u_cla32_xor16 = s_CSAwallace_cla16_u_cla32_pg_logic16_xor0 ^ s_CSAwallace_cla16_u_cla32_or19;
  assign s_CSAwallace_cla16_u_cla32_and46 = s_CSAwallace_cla16_u_cla32_or19 & s_CSAwallace_cla16_u_cla32_pg_logic16_or0;
  assign s_CSAwallace_cla16_u_cla32_or20 = s_CSAwallace_cla16_u_cla32_pg_logic16_and0 | s_CSAwallace_cla16_u_cla32_and46;
  assign s_CSAwallace_cla16_u_cla32_pg_logic17_or0 = s_CSAwallace_cla16_csa13_csa_component_fa17_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic17_and0 = s_CSAwallace_cla16_csa13_csa_component_fa17_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic17_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa17_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa16_or0;
  assign s_CSAwallace_cla16_u_cla32_xor17 = s_CSAwallace_cla16_u_cla32_pg_logic17_xor0 ^ s_CSAwallace_cla16_u_cla32_or20;
  assign s_CSAwallace_cla16_u_cla32_and47 = s_CSAwallace_cla16_u_cla32_or19 & s_CSAwallace_cla16_u_cla32_pg_logic17_or0;
  assign s_CSAwallace_cla16_u_cla32_and48 = s_CSAwallace_cla16_u_cla32_and47 & s_CSAwallace_cla16_u_cla32_pg_logic16_or0;
  assign s_CSAwallace_cla16_u_cla32_and49 = s_CSAwallace_cla16_u_cla32_pg_logic16_and0 & s_CSAwallace_cla16_u_cla32_pg_logic17_or0;
  assign s_CSAwallace_cla16_u_cla32_or21 = s_CSAwallace_cla16_u_cla32_and48 | s_CSAwallace_cla16_u_cla32_and49;
  assign s_CSAwallace_cla16_u_cla32_or22 = s_CSAwallace_cla16_u_cla32_pg_logic17_and0 | s_CSAwallace_cla16_u_cla32_or21;
  assign s_CSAwallace_cla16_u_cla32_pg_logic18_or0 = s_CSAwallace_cla16_csa13_csa_component_fa18_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic18_and0 = s_CSAwallace_cla16_csa13_csa_component_fa18_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic18_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa18_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa17_or0;
  assign s_CSAwallace_cla16_u_cla32_xor18 = s_CSAwallace_cla16_u_cla32_pg_logic18_xor0 ^ s_CSAwallace_cla16_u_cla32_or22;
  assign s_CSAwallace_cla16_u_cla32_and50 = s_CSAwallace_cla16_u_cla32_or19 & s_CSAwallace_cla16_u_cla32_pg_logic17_or0;
  assign s_CSAwallace_cla16_u_cla32_and51 = s_CSAwallace_cla16_u_cla32_pg_logic18_or0 & s_CSAwallace_cla16_u_cla32_pg_logic16_or0;
  assign s_CSAwallace_cla16_u_cla32_and52 = s_CSAwallace_cla16_u_cla32_and50 & s_CSAwallace_cla16_u_cla32_and51;
  assign s_CSAwallace_cla16_u_cla32_and53 = s_CSAwallace_cla16_u_cla32_pg_logic16_and0 & s_CSAwallace_cla16_u_cla32_pg_logic18_or0;
  assign s_CSAwallace_cla16_u_cla32_and54 = s_CSAwallace_cla16_u_cla32_and53 & s_CSAwallace_cla16_u_cla32_pg_logic17_or0;
  assign s_CSAwallace_cla16_u_cla32_and55 = s_CSAwallace_cla16_u_cla32_pg_logic17_and0 & s_CSAwallace_cla16_u_cla32_pg_logic18_or0;
  assign s_CSAwallace_cla16_u_cla32_or23 = s_CSAwallace_cla16_u_cla32_and52 | s_CSAwallace_cla16_u_cla32_and54;
  assign s_CSAwallace_cla16_u_cla32_or24 = s_CSAwallace_cla16_u_cla32_or23 | s_CSAwallace_cla16_u_cla32_and55;
  assign s_CSAwallace_cla16_u_cla32_or25 = s_CSAwallace_cla16_u_cla32_pg_logic18_and0 | s_CSAwallace_cla16_u_cla32_or24;
  assign s_CSAwallace_cla16_u_cla32_pg_logic19_or0 = s_CSAwallace_cla16_csa13_csa_component_fa19_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic19_and0 = s_CSAwallace_cla16_csa13_csa_component_fa19_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic19_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa19_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa18_or0;
  assign s_CSAwallace_cla16_u_cla32_xor19 = s_CSAwallace_cla16_u_cla32_pg_logic19_xor0 ^ s_CSAwallace_cla16_u_cla32_or25;
  assign s_CSAwallace_cla16_u_cla32_and56 = s_CSAwallace_cla16_u_cla32_or19 & s_CSAwallace_cla16_u_cla32_pg_logic18_or0;
  assign s_CSAwallace_cla16_u_cla32_and57 = s_CSAwallace_cla16_u_cla32_pg_logic19_or0 & s_CSAwallace_cla16_u_cla32_pg_logic17_or0;
  assign s_CSAwallace_cla16_u_cla32_and58 = s_CSAwallace_cla16_u_cla32_and56 & s_CSAwallace_cla16_u_cla32_and57;
  assign s_CSAwallace_cla16_u_cla32_and59 = s_CSAwallace_cla16_u_cla32_and58 & s_CSAwallace_cla16_u_cla32_pg_logic16_or0;
  assign s_CSAwallace_cla16_u_cla32_and60 = s_CSAwallace_cla16_u_cla32_pg_logic16_and0 & s_CSAwallace_cla16_u_cla32_pg_logic18_or0;
  assign s_CSAwallace_cla16_u_cla32_and61 = s_CSAwallace_cla16_u_cla32_pg_logic19_or0 & s_CSAwallace_cla16_u_cla32_pg_logic17_or0;
  assign s_CSAwallace_cla16_u_cla32_and62 = s_CSAwallace_cla16_u_cla32_and60 & s_CSAwallace_cla16_u_cla32_and61;
  assign s_CSAwallace_cla16_u_cla32_and63 = s_CSAwallace_cla16_u_cla32_pg_logic17_and0 & s_CSAwallace_cla16_u_cla32_pg_logic19_or0;
  assign s_CSAwallace_cla16_u_cla32_and64 = s_CSAwallace_cla16_u_cla32_and63 & s_CSAwallace_cla16_u_cla32_pg_logic18_or0;
  assign s_CSAwallace_cla16_u_cla32_and65 = s_CSAwallace_cla16_u_cla32_pg_logic18_and0 & s_CSAwallace_cla16_u_cla32_pg_logic19_or0;
  assign s_CSAwallace_cla16_u_cla32_or26 = s_CSAwallace_cla16_u_cla32_and59 | s_CSAwallace_cla16_u_cla32_and64;
  assign s_CSAwallace_cla16_u_cla32_or27 = s_CSAwallace_cla16_u_cla32_and62 | s_CSAwallace_cla16_u_cla32_and65;
  assign s_CSAwallace_cla16_u_cla32_or28 = s_CSAwallace_cla16_u_cla32_or26 | s_CSAwallace_cla16_u_cla32_or27;
  assign s_CSAwallace_cla16_u_cla32_or29 = s_CSAwallace_cla16_u_cla32_pg_logic19_and0 | s_CSAwallace_cla16_u_cla32_or28;
  assign s_CSAwallace_cla16_u_cla32_pg_logic20_or0 = s_CSAwallace_cla16_csa13_csa_component_fa20_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic20_and0 = s_CSAwallace_cla16_csa13_csa_component_fa20_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic20_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa20_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa19_or0;
  assign s_CSAwallace_cla16_u_cla32_xor20 = s_CSAwallace_cla16_u_cla32_pg_logic20_xor0 ^ s_CSAwallace_cla16_u_cla32_or29;
  assign s_CSAwallace_cla16_u_cla32_and66 = s_CSAwallace_cla16_u_cla32_or29 & s_CSAwallace_cla16_u_cla32_pg_logic20_or0;
  assign s_CSAwallace_cla16_u_cla32_or30 = s_CSAwallace_cla16_u_cla32_pg_logic20_and0 | s_CSAwallace_cla16_u_cla32_and66;
  assign s_CSAwallace_cla16_u_cla32_pg_logic21_or0 = s_CSAwallace_cla16_csa13_csa_component_fa21_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic21_and0 = s_CSAwallace_cla16_csa13_csa_component_fa21_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic21_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa21_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa20_or0;
  assign s_CSAwallace_cla16_u_cla32_xor21 = s_CSAwallace_cla16_u_cla32_pg_logic21_xor0 ^ s_CSAwallace_cla16_u_cla32_or30;
  assign s_CSAwallace_cla16_u_cla32_and67 = s_CSAwallace_cla16_u_cla32_or29 & s_CSAwallace_cla16_u_cla32_pg_logic21_or0;
  assign s_CSAwallace_cla16_u_cla32_and68 = s_CSAwallace_cla16_u_cla32_and67 & s_CSAwallace_cla16_u_cla32_pg_logic20_or0;
  assign s_CSAwallace_cla16_u_cla32_and69 = s_CSAwallace_cla16_u_cla32_pg_logic20_and0 & s_CSAwallace_cla16_u_cla32_pg_logic21_or0;
  assign s_CSAwallace_cla16_u_cla32_or31 = s_CSAwallace_cla16_u_cla32_and68 | s_CSAwallace_cla16_u_cla32_and69;
  assign s_CSAwallace_cla16_u_cla32_or32 = s_CSAwallace_cla16_u_cla32_pg_logic21_and0 | s_CSAwallace_cla16_u_cla32_or31;
  assign s_CSAwallace_cla16_u_cla32_pg_logic22_or0 = s_CSAwallace_cla16_csa13_csa_component_fa22_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic22_and0 = s_CSAwallace_cla16_csa13_csa_component_fa22_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic22_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa22_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa21_or0;
  assign s_CSAwallace_cla16_u_cla32_xor22 = s_CSAwallace_cla16_u_cla32_pg_logic22_xor0 ^ s_CSAwallace_cla16_u_cla32_or32;
  assign s_CSAwallace_cla16_u_cla32_and70 = s_CSAwallace_cla16_u_cla32_or29 & s_CSAwallace_cla16_u_cla32_pg_logic21_or0;
  assign s_CSAwallace_cla16_u_cla32_and71 = s_CSAwallace_cla16_u_cla32_pg_logic22_or0 & s_CSAwallace_cla16_u_cla32_pg_logic20_or0;
  assign s_CSAwallace_cla16_u_cla32_and72 = s_CSAwallace_cla16_u_cla32_and70 & s_CSAwallace_cla16_u_cla32_and71;
  assign s_CSAwallace_cla16_u_cla32_and73 = s_CSAwallace_cla16_u_cla32_pg_logic20_and0 & s_CSAwallace_cla16_u_cla32_pg_logic22_or0;
  assign s_CSAwallace_cla16_u_cla32_and74 = s_CSAwallace_cla16_u_cla32_and73 & s_CSAwallace_cla16_u_cla32_pg_logic21_or0;
  assign s_CSAwallace_cla16_u_cla32_and75 = s_CSAwallace_cla16_u_cla32_pg_logic21_and0 & s_CSAwallace_cla16_u_cla32_pg_logic22_or0;
  assign s_CSAwallace_cla16_u_cla32_or33 = s_CSAwallace_cla16_u_cla32_and72 | s_CSAwallace_cla16_u_cla32_and74;
  assign s_CSAwallace_cla16_u_cla32_or34 = s_CSAwallace_cla16_u_cla32_or33 | s_CSAwallace_cla16_u_cla32_and75;
  assign s_CSAwallace_cla16_u_cla32_or35 = s_CSAwallace_cla16_u_cla32_pg_logic22_and0 | s_CSAwallace_cla16_u_cla32_or34;
  assign s_CSAwallace_cla16_u_cla32_pg_logic23_or0 = s_CSAwallace_cla16_csa13_csa_component_fa23_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic23_and0 = s_CSAwallace_cla16_csa13_csa_component_fa23_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic23_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa23_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa22_or0;
  assign s_CSAwallace_cla16_u_cla32_xor23 = s_CSAwallace_cla16_u_cla32_pg_logic23_xor0 ^ s_CSAwallace_cla16_u_cla32_or35;
  assign s_CSAwallace_cla16_u_cla32_and76 = s_CSAwallace_cla16_u_cla32_or29 & s_CSAwallace_cla16_u_cla32_pg_logic22_or0;
  assign s_CSAwallace_cla16_u_cla32_and77 = s_CSAwallace_cla16_u_cla32_pg_logic23_or0 & s_CSAwallace_cla16_u_cla32_pg_logic21_or0;
  assign s_CSAwallace_cla16_u_cla32_and78 = s_CSAwallace_cla16_u_cla32_and76 & s_CSAwallace_cla16_u_cla32_and77;
  assign s_CSAwallace_cla16_u_cla32_and79 = s_CSAwallace_cla16_u_cla32_and78 & s_CSAwallace_cla16_u_cla32_pg_logic20_or0;
  assign s_CSAwallace_cla16_u_cla32_and80 = s_CSAwallace_cla16_u_cla32_pg_logic20_and0 & s_CSAwallace_cla16_u_cla32_pg_logic22_or0;
  assign s_CSAwallace_cla16_u_cla32_and81 = s_CSAwallace_cla16_u_cla32_pg_logic23_or0 & s_CSAwallace_cla16_u_cla32_pg_logic21_or0;
  assign s_CSAwallace_cla16_u_cla32_and82 = s_CSAwallace_cla16_u_cla32_and80 & s_CSAwallace_cla16_u_cla32_and81;
  assign s_CSAwallace_cla16_u_cla32_and83 = s_CSAwallace_cla16_u_cla32_pg_logic21_and0 & s_CSAwallace_cla16_u_cla32_pg_logic23_or0;
  assign s_CSAwallace_cla16_u_cla32_and84 = s_CSAwallace_cla16_u_cla32_and83 & s_CSAwallace_cla16_u_cla32_pg_logic22_or0;
  assign s_CSAwallace_cla16_u_cla32_and85 = s_CSAwallace_cla16_u_cla32_pg_logic22_and0 & s_CSAwallace_cla16_u_cla32_pg_logic23_or0;
  assign s_CSAwallace_cla16_u_cla32_or36 = s_CSAwallace_cla16_u_cla32_and79 | s_CSAwallace_cla16_u_cla32_and84;
  assign s_CSAwallace_cla16_u_cla32_or37 = s_CSAwallace_cla16_u_cla32_and82 | s_CSAwallace_cla16_u_cla32_and85;
  assign s_CSAwallace_cla16_u_cla32_or38 = s_CSAwallace_cla16_u_cla32_or36 | s_CSAwallace_cla16_u_cla32_or37;
  assign s_CSAwallace_cla16_u_cla32_or39 = s_CSAwallace_cla16_u_cla32_pg_logic23_and0 | s_CSAwallace_cla16_u_cla32_or38;
  assign s_CSAwallace_cla16_u_cla32_pg_logic24_or0 = s_CSAwallace_cla16_csa13_csa_component_fa24_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic24_and0 = s_CSAwallace_cla16_csa13_csa_component_fa24_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic24_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa24_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa23_or0;
  assign s_CSAwallace_cla16_u_cla32_xor24 = s_CSAwallace_cla16_u_cla32_pg_logic24_xor0 ^ s_CSAwallace_cla16_u_cla32_or39;
  assign s_CSAwallace_cla16_u_cla32_and86 = s_CSAwallace_cla16_u_cla32_or39 & s_CSAwallace_cla16_u_cla32_pg_logic24_or0;
  assign s_CSAwallace_cla16_u_cla32_or40 = s_CSAwallace_cla16_u_cla32_pg_logic24_and0 | s_CSAwallace_cla16_u_cla32_and86;
  assign s_CSAwallace_cla16_u_cla32_pg_logic25_or0 = s_CSAwallace_cla16_csa13_csa_component_fa25_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic25_and0 = s_CSAwallace_cla16_csa13_csa_component_fa25_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic25_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa25_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa24_or0;
  assign s_CSAwallace_cla16_u_cla32_xor25 = s_CSAwallace_cla16_u_cla32_pg_logic25_xor0 ^ s_CSAwallace_cla16_u_cla32_or40;
  assign s_CSAwallace_cla16_u_cla32_and87 = s_CSAwallace_cla16_u_cla32_or39 & s_CSAwallace_cla16_u_cla32_pg_logic25_or0;
  assign s_CSAwallace_cla16_u_cla32_and88 = s_CSAwallace_cla16_u_cla32_and87 & s_CSAwallace_cla16_u_cla32_pg_logic24_or0;
  assign s_CSAwallace_cla16_u_cla32_and89 = s_CSAwallace_cla16_u_cla32_pg_logic24_and0 & s_CSAwallace_cla16_u_cla32_pg_logic25_or0;
  assign s_CSAwallace_cla16_u_cla32_or41 = s_CSAwallace_cla16_u_cla32_and88 | s_CSAwallace_cla16_u_cla32_and89;
  assign s_CSAwallace_cla16_u_cla32_or42 = s_CSAwallace_cla16_u_cla32_pg_logic25_and0 | s_CSAwallace_cla16_u_cla32_or41;
  assign s_CSAwallace_cla16_u_cla32_pg_logic26_or0 = s_CSAwallace_cla16_csa13_csa_component_fa26_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic26_and0 = s_CSAwallace_cla16_csa13_csa_component_fa26_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic26_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa26_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa25_or0;
  assign s_CSAwallace_cla16_u_cla32_xor26 = s_CSAwallace_cla16_u_cla32_pg_logic26_xor0 ^ s_CSAwallace_cla16_u_cla32_or42;
  assign s_CSAwallace_cla16_u_cla32_and90 = s_CSAwallace_cla16_u_cla32_or39 & s_CSAwallace_cla16_u_cla32_pg_logic25_or0;
  assign s_CSAwallace_cla16_u_cla32_and91 = s_CSAwallace_cla16_u_cla32_pg_logic26_or0 & s_CSAwallace_cla16_u_cla32_pg_logic24_or0;
  assign s_CSAwallace_cla16_u_cla32_and92 = s_CSAwallace_cla16_u_cla32_and90 & s_CSAwallace_cla16_u_cla32_and91;
  assign s_CSAwallace_cla16_u_cla32_and93 = s_CSAwallace_cla16_u_cla32_pg_logic24_and0 & s_CSAwallace_cla16_u_cla32_pg_logic26_or0;
  assign s_CSAwallace_cla16_u_cla32_and94 = s_CSAwallace_cla16_u_cla32_and93 & s_CSAwallace_cla16_u_cla32_pg_logic25_or0;
  assign s_CSAwallace_cla16_u_cla32_and95 = s_CSAwallace_cla16_u_cla32_pg_logic25_and0 & s_CSAwallace_cla16_u_cla32_pg_logic26_or0;
  assign s_CSAwallace_cla16_u_cla32_or43 = s_CSAwallace_cla16_u_cla32_and92 | s_CSAwallace_cla16_u_cla32_and94;
  assign s_CSAwallace_cla16_u_cla32_or44 = s_CSAwallace_cla16_u_cla32_or43 | s_CSAwallace_cla16_u_cla32_and95;
  assign s_CSAwallace_cla16_u_cla32_or45 = s_CSAwallace_cla16_u_cla32_pg_logic26_and0 | s_CSAwallace_cla16_u_cla32_or44;
  assign s_CSAwallace_cla16_u_cla32_pg_logic27_or0 = s_CSAwallace_cla16_csa13_csa_component_fa27_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic27_and0 = s_CSAwallace_cla16_csa13_csa_component_fa27_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic27_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa27_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa26_or0;
  assign s_CSAwallace_cla16_u_cla32_xor27 = s_CSAwallace_cla16_u_cla32_pg_logic27_xor0 ^ s_CSAwallace_cla16_u_cla32_or45;
  assign s_CSAwallace_cla16_u_cla32_and96 = s_CSAwallace_cla16_u_cla32_or39 & s_CSAwallace_cla16_u_cla32_pg_logic26_or0;
  assign s_CSAwallace_cla16_u_cla32_and97 = s_CSAwallace_cla16_u_cla32_pg_logic27_or0 & s_CSAwallace_cla16_u_cla32_pg_logic25_or0;
  assign s_CSAwallace_cla16_u_cla32_and98 = s_CSAwallace_cla16_u_cla32_and96 & s_CSAwallace_cla16_u_cla32_and97;
  assign s_CSAwallace_cla16_u_cla32_and99 = s_CSAwallace_cla16_u_cla32_and98 & s_CSAwallace_cla16_u_cla32_pg_logic24_or0;
  assign s_CSAwallace_cla16_u_cla32_and100 = s_CSAwallace_cla16_u_cla32_pg_logic24_and0 & s_CSAwallace_cla16_u_cla32_pg_logic26_or0;
  assign s_CSAwallace_cla16_u_cla32_and101 = s_CSAwallace_cla16_u_cla32_pg_logic27_or0 & s_CSAwallace_cla16_u_cla32_pg_logic25_or0;
  assign s_CSAwallace_cla16_u_cla32_and102 = s_CSAwallace_cla16_u_cla32_and100 & s_CSAwallace_cla16_u_cla32_and101;
  assign s_CSAwallace_cla16_u_cla32_and103 = s_CSAwallace_cla16_u_cla32_pg_logic25_and0 & s_CSAwallace_cla16_u_cla32_pg_logic27_or0;
  assign s_CSAwallace_cla16_u_cla32_and104 = s_CSAwallace_cla16_u_cla32_and103 & s_CSAwallace_cla16_u_cla32_pg_logic26_or0;
  assign s_CSAwallace_cla16_u_cla32_and105 = s_CSAwallace_cla16_u_cla32_pg_logic26_and0 & s_CSAwallace_cla16_u_cla32_pg_logic27_or0;
  assign s_CSAwallace_cla16_u_cla32_or46 = s_CSAwallace_cla16_u_cla32_and99 | s_CSAwallace_cla16_u_cla32_and104;
  assign s_CSAwallace_cla16_u_cla32_or47 = s_CSAwallace_cla16_u_cla32_and102 | s_CSAwallace_cla16_u_cla32_and105;
  assign s_CSAwallace_cla16_u_cla32_or48 = s_CSAwallace_cla16_u_cla32_or46 | s_CSAwallace_cla16_u_cla32_or47;
  assign s_CSAwallace_cla16_u_cla32_or49 = s_CSAwallace_cla16_u_cla32_pg_logic27_and0 | s_CSAwallace_cla16_u_cla32_or48;
  assign s_CSAwallace_cla16_u_cla32_pg_logic28_or0 = s_CSAwallace_cla16_csa13_csa_component_fa28_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic28_and0 = s_CSAwallace_cla16_csa13_csa_component_fa28_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic28_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa28_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa27_or0;
  assign s_CSAwallace_cla16_u_cla32_xor28 = s_CSAwallace_cla16_u_cla32_pg_logic28_xor0 ^ s_CSAwallace_cla16_u_cla32_or49;
  assign s_CSAwallace_cla16_u_cla32_and106 = s_CSAwallace_cla16_u_cla32_or49 & s_CSAwallace_cla16_u_cla32_pg_logic28_or0;
  assign s_CSAwallace_cla16_u_cla32_or50 = s_CSAwallace_cla16_u_cla32_pg_logic28_and0 | s_CSAwallace_cla16_u_cla32_and106;
  assign s_CSAwallace_cla16_u_cla32_pg_logic29_or0 = s_CSAwallace_cla16_csa13_csa_component_fa29_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic29_and0 = s_CSAwallace_cla16_csa13_csa_component_fa29_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic29_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa29_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa28_or0;
  assign s_CSAwallace_cla16_u_cla32_xor29 = s_CSAwallace_cla16_u_cla32_pg_logic29_xor0 ^ s_CSAwallace_cla16_u_cla32_or50;
  assign s_CSAwallace_cla16_u_cla32_and107 = s_CSAwallace_cla16_u_cla32_or49 & s_CSAwallace_cla16_u_cla32_pg_logic29_or0;
  assign s_CSAwallace_cla16_u_cla32_and108 = s_CSAwallace_cla16_u_cla32_and107 & s_CSAwallace_cla16_u_cla32_pg_logic28_or0;
  assign s_CSAwallace_cla16_u_cla32_and109 = s_CSAwallace_cla16_u_cla32_pg_logic28_and0 & s_CSAwallace_cla16_u_cla32_pg_logic29_or0;
  assign s_CSAwallace_cla16_u_cla32_or51 = s_CSAwallace_cla16_u_cla32_and108 | s_CSAwallace_cla16_u_cla32_and109;
  assign s_CSAwallace_cla16_u_cla32_or52 = s_CSAwallace_cla16_u_cla32_pg_logic29_and0 | s_CSAwallace_cla16_u_cla32_or51;
  assign s_CSAwallace_cla16_u_cla32_pg_logic30_or0 = s_CSAwallace_cla16_csa13_csa_component_fa30_xor1 | s_CSAwallace_cla16_csa13_csa_component_fa29_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic30_and0 = s_CSAwallace_cla16_csa13_csa_component_fa30_xor1 & s_CSAwallace_cla16_csa13_csa_component_fa29_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic30_xor0 = s_CSAwallace_cla16_csa13_csa_component_fa30_xor1 ^ s_CSAwallace_cla16_csa13_csa_component_fa29_or0;
  assign s_CSAwallace_cla16_u_cla32_xor30 = s_CSAwallace_cla16_u_cla32_pg_logic30_xor0 ^ s_CSAwallace_cla16_u_cla32_or52;
  assign s_CSAwallace_cla16_u_cla32_and110 = s_CSAwallace_cla16_u_cla32_or49 & s_CSAwallace_cla16_u_cla32_pg_logic29_or0;
  assign s_CSAwallace_cla16_u_cla32_and111 = s_CSAwallace_cla16_u_cla32_pg_logic30_or0 & s_CSAwallace_cla16_u_cla32_pg_logic28_or0;
  assign s_CSAwallace_cla16_u_cla32_and112 = s_CSAwallace_cla16_u_cla32_and110 & s_CSAwallace_cla16_u_cla32_and111;
  assign s_CSAwallace_cla16_u_cla32_and113 = s_CSAwallace_cla16_u_cla32_pg_logic28_and0 & s_CSAwallace_cla16_u_cla32_pg_logic30_or0;
  assign s_CSAwallace_cla16_u_cla32_and114 = s_CSAwallace_cla16_u_cla32_and113 & s_CSAwallace_cla16_u_cla32_pg_logic29_or0;
  assign s_CSAwallace_cla16_u_cla32_and115 = s_CSAwallace_cla16_u_cla32_pg_logic29_and0 & s_CSAwallace_cla16_u_cla32_pg_logic30_or0;
  assign s_CSAwallace_cla16_u_cla32_or53 = s_CSAwallace_cla16_u_cla32_and112 | s_CSAwallace_cla16_u_cla32_and114;
  assign s_CSAwallace_cla16_u_cla32_or54 = s_CSAwallace_cla16_u_cla32_or53 | s_CSAwallace_cla16_u_cla32_and115;
  assign s_CSAwallace_cla16_u_cla32_or55 = s_CSAwallace_cla16_u_cla32_pg_logic30_and0 | s_CSAwallace_cla16_u_cla32_or54;
  assign s_CSAwallace_cla16_u_cla32_pg_logic31_or0 = s_CSAwallace_cla16_csa11_csa_component_fa30_or0 | s_CSAwallace_cla16_csa13_csa_component_fa30_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic31_and0 = s_CSAwallace_cla16_csa11_csa_component_fa30_or0 & s_CSAwallace_cla16_csa13_csa_component_fa30_or0;
  assign s_CSAwallace_cla16_u_cla32_pg_logic31_xor0 = s_CSAwallace_cla16_csa11_csa_component_fa30_or0 ^ s_CSAwallace_cla16_csa13_csa_component_fa30_or0;
  assign s_CSAwallace_cla16_u_cla32_xor31 = s_CSAwallace_cla16_u_cla32_pg_logic31_xor0 ^ s_CSAwallace_cla16_u_cla32_or55;
  assign s_CSAwallace_cla16_u_cla32_and116 = s_CSAwallace_cla16_u_cla32_or49 & s_CSAwallace_cla16_u_cla32_pg_logic30_or0;
  assign s_CSAwallace_cla16_u_cla32_and117 = s_CSAwallace_cla16_u_cla32_pg_logic31_or0 & s_CSAwallace_cla16_u_cla32_pg_logic29_or0;
  assign s_CSAwallace_cla16_u_cla32_and118 = s_CSAwallace_cla16_u_cla32_and116 & s_CSAwallace_cla16_u_cla32_and117;
  assign s_CSAwallace_cla16_u_cla32_and119 = s_CSAwallace_cla16_u_cla32_and118 & s_CSAwallace_cla16_u_cla32_pg_logic28_or0;
  assign s_CSAwallace_cla16_u_cla32_and120 = s_CSAwallace_cla16_u_cla32_pg_logic28_and0 & s_CSAwallace_cla16_u_cla32_pg_logic30_or0;
  assign s_CSAwallace_cla16_u_cla32_and121 = s_CSAwallace_cla16_u_cla32_pg_logic31_or0 & s_CSAwallace_cla16_u_cla32_pg_logic29_or0;
  assign s_CSAwallace_cla16_u_cla32_and122 = s_CSAwallace_cla16_u_cla32_and120 & s_CSAwallace_cla16_u_cla32_and121;
  assign s_CSAwallace_cla16_u_cla32_and123 = s_CSAwallace_cla16_u_cla32_pg_logic29_and0 & s_CSAwallace_cla16_u_cla32_pg_logic31_or0;
  assign s_CSAwallace_cla16_u_cla32_and124 = s_CSAwallace_cla16_u_cla32_and123 & s_CSAwallace_cla16_u_cla32_pg_logic30_or0;
  assign s_CSAwallace_cla16_u_cla32_and125 = s_CSAwallace_cla16_u_cla32_pg_logic30_and0 & s_CSAwallace_cla16_u_cla32_pg_logic31_or0;
  assign s_CSAwallace_cla16_u_cla32_or56 = s_CSAwallace_cla16_u_cla32_and119 | s_CSAwallace_cla16_u_cla32_and124;
  assign s_CSAwallace_cla16_u_cla32_or57 = s_CSAwallace_cla16_u_cla32_and122 | s_CSAwallace_cla16_u_cla32_and125;
  assign s_CSAwallace_cla16_u_cla32_or58 = s_CSAwallace_cla16_u_cla32_or56 | s_CSAwallace_cla16_u_cla32_or57;
  assign s_CSAwallace_cla16_u_cla32_or59 = s_CSAwallace_cla16_u_cla32_pg_logic31_and0 | s_CSAwallace_cla16_u_cla32_or58;
  assign s_CSAwallace_cla16_xor0 = ~s_CSAwallace_cla16_u_cla32_xor31;

  assign s_CSAwallace_cla16_out[0] = s_CSAwallace_cla16_and_0_0;
  assign s_CSAwallace_cla16_out[1] = s_CSAwallace_cla16_csa0_csa_component_fa1_xor0;
  assign s_CSAwallace_cla16_out[2] = s_CSAwallace_cla16_csa5_csa_component_fa2_xor0;
  assign s_CSAwallace_cla16_out[3] = s_CSAwallace_cla16_csa8_csa_component_fa3_xor0;
  assign s_CSAwallace_cla16_out[4] = s_CSAwallace_cla16_csa10_csa_component_fa4_xor0;
  assign s_CSAwallace_cla16_out[5] = s_CSAwallace_cla16_csa12_csa_component_fa5_xor0;
  assign s_CSAwallace_cla16_out[6] = s_CSAwallace_cla16_csa13_csa_component_fa6_xor0;
  assign s_CSAwallace_cla16_out[7] = s_CSAwallace_cla16_u_cla32_pg_logic7_xor0;
  assign s_CSAwallace_cla16_out[8] = s_CSAwallace_cla16_u_cla32_xor8;
  assign s_CSAwallace_cla16_out[9] = s_CSAwallace_cla16_u_cla32_xor9;
  assign s_CSAwallace_cla16_out[10] = s_CSAwallace_cla16_u_cla32_xor10;
  assign s_CSAwallace_cla16_out[11] = s_CSAwallace_cla16_u_cla32_xor11;
  assign s_CSAwallace_cla16_out[12] = s_CSAwallace_cla16_u_cla32_xor12;
  assign s_CSAwallace_cla16_out[13] = s_CSAwallace_cla16_u_cla32_xor13;
  assign s_CSAwallace_cla16_out[14] = s_CSAwallace_cla16_u_cla32_xor14;
  assign s_CSAwallace_cla16_out[15] = s_CSAwallace_cla16_u_cla32_xor15;
  assign s_CSAwallace_cla16_out[16] = s_CSAwallace_cla16_u_cla32_xor16;
  assign s_CSAwallace_cla16_out[17] = s_CSAwallace_cla16_u_cla32_xor17;
  assign s_CSAwallace_cla16_out[18] = s_CSAwallace_cla16_u_cla32_xor18;
  assign s_CSAwallace_cla16_out[19] = s_CSAwallace_cla16_u_cla32_xor19;
  assign s_CSAwallace_cla16_out[20] = s_CSAwallace_cla16_u_cla32_xor20;
  assign s_CSAwallace_cla16_out[21] = s_CSAwallace_cla16_u_cla32_xor21;
  assign s_CSAwallace_cla16_out[22] = s_CSAwallace_cla16_u_cla32_xor22;
  assign s_CSAwallace_cla16_out[23] = s_CSAwallace_cla16_u_cla32_xor23;
  assign s_CSAwallace_cla16_out[24] = s_CSAwallace_cla16_u_cla32_xor24;
  assign s_CSAwallace_cla16_out[25] = s_CSAwallace_cla16_u_cla32_xor25;
  assign s_CSAwallace_cla16_out[26] = s_CSAwallace_cla16_u_cla32_xor26;
  assign s_CSAwallace_cla16_out[27] = s_CSAwallace_cla16_u_cla32_xor27;
  assign s_CSAwallace_cla16_out[28] = s_CSAwallace_cla16_u_cla32_xor28;
  assign s_CSAwallace_cla16_out[29] = s_CSAwallace_cla16_u_cla32_xor29;
  assign s_CSAwallace_cla16_out[30] = s_CSAwallace_cla16_u_cla32_xor30;
  assign s_CSAwallace_cla16_out[31] = s_CSAwallace_cla16_xor0;
endmodule