module u_pg_rca12(input [11:0] a, input [11:0] b, output [12:0] u_pg_rca12_out);
  wire u_pg_rca12_pg_fa0_xor0;
  wire u_pg_rca12_pg_fa0_and0;
  wire u_pg_rca12_pg_fa1_xor0;
  wire u_pg_rca12_pg_fa1_and0;
  wire u_pg_rca12_pg_fa1_xor1;
  wire u_pg_rca12_and1;
  wire u_pg_rca12_or1;
  wire u_pg_rca12_pg_fa2_xor0;
  wire u_pg_rca12_pg_fa2_and0;
  wire u_pg_rca12_pg_fa2_xor1;
  wire u_pg_rca12_and2;
  wire u_pg_rca12_or2;
  wire u_pg_rca12_pg_fa3_xor0;
  wire u_pg_rca12_pg_fa3_and0;
  wire u_pg_rca12_pg_fa3_xor1;
  wire u_pg_rca12_and3;
  wire u_pg_rca12_or3;
  wire u_pg_rca12_pg_fa4_xor0;
  wire u_pg_rca12_pg_fa4_and0;
  wire u_pg_rca12_pg_fa4_xor1;
  wire u_pg_rca12_and4;
  wire u_pg_rca12_or4;
  wire u_pg_rca12_pg_fa5_xor0;
  wire u_pg_rca12_pg_fa5_and0;
  wire u_pg_rca12_pg_fa5_xor1;
  wire u_pg_rca12_and5;
  wire u_pg_rca12_or5;
  wire u_pg_rca12_pg_fa6_xor0;
  wire u_pg_rca12_pg_fa6_and0;
  wire u_pg_rca12_pg_fa6_xor1;
  wire u_pg_rca12_and6;
  wire u_pg_rca12_or6;
  wire u_pg_rca12_pg_fa7_xor0;
  wire u_pg_rca12_pg_fa7_and0;
  wire u_pg_rca12_pg_fa7_xor1;
  wire u_pg_rca12_and7;
  wire u_pg_rca12_or7;
  wire u_pg_rca12_pg_fa8_xor0;
  wire u_pg_rca12_pg_fa8_and0;
  wire u_pg_rca12_pg_fa8_xor1;
  wire u_pg_rca12_and8;
  wire u_pg_rca12_or8;
  wire u_pg_rca12_pg_fa9_xor0;
  wire u_pg_rca12_pg_fa9_and0;
  wire u_pg_rca12_pg_fa9_xor1;
  wire u_pg_rca12_and9;
  wire u_pg_rca12_or9;
  wire u_pg_rca12_pg_fa10_xor0;
  wire u_pg_rca12_pg_fa10_and0;
  wire u_pg_rca12_pg_fa10_xor1;
  wire u_pg_rca12_and10;
  wire u_pg_rca12_or10;
  wire u_pg_rca12_pg_fa11_xor0;
  wire u_pg_rca12_pg_fa11_and0;
  wire u_pg_rca12_pg_fa11_xor1;
  wire u_pg_rca12_and11;
  wire u_pg_rca12_or11;

  assign u_pg_rca12_pg_fa0_xor0 = a[0] ^ b[0];
  assign u_pg_rca12_pg_fa0_and0 = a[0] & b[0];
  assign u_pg_rca12_pg_fa1_xor0 = a[1] ^ b[1];
  assign u_pg_rca12_pg_fa1_and0 = a[1] & b[1];
  assign u_pg_rca12_pg_fa1_xor1 = u_pg_rca12_pg_fa1_xor0 ^ u_pg_rca12_pg_fa0_and0;
  assign u_pg_rca12_and1 = u_pg_rca12_pg_fa0_and0 & u_pg_rca12_pg_fa1_xor0;
  assign u_pg_rca12_or1 = u_pg_rca12_and1 | u_pg_rca12_pg_fa1_and0;
  assign u_pg_rca12_pg_fa2_xor0 = a[2] ^ b[2];
  assign u_pg_rca12_pg_fa2_and0 = a[2] & b[2];
  assign u_pg_rca12_pg_fa2_xor1 = u_pg_rca12_pg_fa2_xor0 ^ u_pg_rca12_or1;
  assign u_pg_rca12_and2 = u_pg_rca12_or1 & u_pg_rca12_pg_fa2_xor0;
  assign u_pg_rca12_or2 = u_pg_rca12_and2 | u_pg_rca12_pg_fa2_and0;
  assign u_pg_rca12_pg_fa3_xor0 = a[3] ^ b[3];
  assign u_pg_rca12_pg_fa3_and0 = a[3] & b[3];
  assign u_pg_rca12_pg_fa3_xor1 = u_pg_rca12_pg_fa3_xor0 ^ u_pg_rca12_or2;
  assign u_pg_rca12_and3 = u_pg_rca12_or2 & u_pg_rca12_pg_fa3_xor0;
  assign u_pg_rca12_or3 = u_pg_rca12_and3 | u_pg_rca12_pg_fa3_and0;
  assign u_pg_rca12_pg_fa4_xor0 = a[4] ^ b[4];
  assign u_pg_rca12_pg_fa4_and0 = a[4] & b[4];
  assign u_pg_rca12_pg_fa4_xor1 = u_pg_rca12_pg_fa4_xor0 ^ u_pg_rca12_or3;
  assign u_pg_rca12_and4 = u_pg_rca12_or3 & u_pg_rca12_pg_fa4_xor0;
  assign u_pg_rca12_or4 = u_pg_rca12_and4 | u_pg_rca12_pg_fa4_and0;
  assign u_pg_rca12_pg_fa5_xor0 = a[5] ^ b[5];
  assign u_pg_rca12_pg_fa5_and0 = a[5] & b[5];
  assign u_pg_rca12_pg_fa5_xor1 = u_pg_rca12_pg_fa5_xor0 ^ u_pg_rca12_or4;
  assign u_pg_rca12_and5 = u_pg_rca12_or4 & u_pg_rca12_pg_fa5_xor0;
  assign u_pg_rca12_or5 = u_pg_rca12_and5 | u_pg_rca12_pg_fa5_and0;
  assign u_pg_rca12_pg_fa6_xor0 = a[6] ^ b[6];
  assign u_pg_rca12_pg_fa6_and0 = a[6] & b[6];
  assign u_pg_rca12_pg_fa6_xor1 = u_pg_rca12_pg_fa6_xor0 ^ u_pg_rca12_or5;
  assign u_pg_rca12_and6 = u_pg_rca12_or5 & u_pg_rca12_pg_fa6_xor0;
  assign u_pg_rca12_or6 = u_pg_rca12_and6 | u_pg_rca12_pg_fa6_and0;
  assign u_pg_rca12_pg_fa7_xor0 = a[7] ^ b[7];
  assign u_pg_rca12_pg_fa7_and0 = a[7] & b[7];
  assign u_pg_rca12_pg_fa7_xor1 = u_pg_rca12_pg_fa7_xor0 ^ u_pg_rca12_or6;
  assign u_pg_rca12_and7 = u_pg_rca12_or6 & u_pg_rca12_pg_fa7_xor0;
  assign u_pg_rca12_or7 = u_pg_rca12_and7 | u_pg_rca12_pg_fa7_and0;
  assign u_pg_rca12_pg_fa8_xor0 = a[8] ^ b[8];
  assign u_pg_rca12_pg_fa8_and0 = a[8] & b[8];
  assign u_pg_rca12_pg_fa8_xor1 = u_pg_rca12_pg_fa8_xor0 ^ u_pg_rca12_or7;
  assign u_pg_rca12_and8 = u_pg_rca12_or7 & u_pg_rca12_pg_fa8_xor0;
  assign u_pg_rca12_or8 = u_pg_rca12_and8 | u_pg_rca12_pg_fa8_and0;
  assign u_pg_rca12_pg_fa9_xor0 = a[9] ^ b[9];
  assign u_pg_rca12_pg_fa9_and0 = a[9] & b[9];
  assign u_pg_rca12_pg_fa9_xor1 = u_pg_rca12_pg_fa9_xor0 ^ u_pg_rca12_or8;
  assign u_pg_rca12_and9 = u_pg_rca12_or8 & u_pg_rca12_pg_fa9_xor0;
  assign u_pg_rca12_or9 = u_pg_rca12_and9 | u_pg_rca12_pg_fa9_and0;
  assign u_pg_rca12_pg_fa10_xor0 = a[10] ^ b[10];
  assign u_pg_rca12_pg_fa10_and0 = a[10] & b[10];
  assign u_pg_rca12_pg_fa10_xor1 = u_pg_rca12_pg_fa10_xor0 ^ u_pg_rca12_or9;
  assign u_pg_rca12_and10 = u_pg_rca12_or9 & u_pg_rca12_pg_fa10_xor0;
  assign u_pg_rca12_or10 = u_pg_rca12_and10 | u_pg_rca12_pg_fa10_and0;
  assign u_pg_rca12_pg_fa11_xor0 = a[11] ^ b[11];
  assign u_pg_rca12_pg_fa11_and0 = a[11] & b[11];
  assign u_pg_rca12_pg_fa11_xor1 = u_pg_rca12_pg_fa11_xor0 ^ u_pg_rca12_or10;
  assign u_pg_rca12_and11 = u_pg_rca12_or10 & u_pg_rca12_pg_fa11_xor0;
  assign u_pg_rca12_or11 = u_pg_rca12_and11 | u_pg_rca12_pg_fa11_and0;

  assign u_pg_rca12_out[0] = u_pg_rca12_pg_fa0_xor0;
  assign u_pg_rca12_out[1] = u_pg_rca12_pg_fa1_xor1;
  assign u_pg_rca12_out[2] = u_pg_rca12_pg_fa2_xor1;
  assign u_pg_rca12_out[3] = u_pg_rca12_pg_fa3_xor1;
  assign u_pg_rca12_out[4] = u_pg_rca12_pg_fa4_xor1;
  assign u_pg_rca12_out[5] = u_pg_rca12_pg_fa5_xor1;
  assign u_pg_rca12_out[6] = u_pg_rca12_pg_fa6_xor1;
  assign u_pg_rca12_out[7] = u_pg_rca12_pg_fa7_xor1;
  assign u_pg_rca12_out[8] = u_pg_rca12_pg_fa8_xor1;
  assign u_pg_rca12_out[9] = u_pg_rca12_pg_fa9_xor1;
  assign u_pg_rca12_out[10] = u_pg_rca12_pg_fa10_xor1;
  assign u_pg_rca12_out[11] = u_pg_rca12_pg_fa11_xor1;
  assign u_pg_rca12_out[12] = u_pg_rca12_or11;
endmodule