module or_gate(input a, input b, output out);
  assign out = a | b;
endmodule

module and_gate(input a, input b, output out);
  assign out = a & b;
endmodule

module xor_gate(input a, input b, output out);
  assign out = a ^ b;
endmodule

module pg_logic(input [0:0] a, input [0:0] b, output [0:0] pg_logic_or0, output [0:0] pg_logic_and0, output [0:0] pg_logic_xor0);
  or_gate or_gate_pg_logic_or0(.a(a[0]), .b(b[0]), .out(pg_logic_or0));
  and_gate and_gate_pg_logic_and0(.a(a[0]), .b(b[0]), .out(pg_logic_and0));
  xor_gate xor_gate_pg_logic_xor0(.a(a[0]), .b(b[0]), .out(pg_logic_xor0));
endmodule

module h_s_cla32(input [31:0] a, input [31:0] b, output [32:0] h_s_cla32_out);
  wire [0:0] h_s_cla32_pg_logic0_or0;
  wire [0:0] h_s_cla32_pg_logic0_and0;
  wire [0:0] h_s_cla32_pg_logic0_xor0;
  wire [0:0] h_s_cla32_pg_logic1_or0;
  wire [0:0] h_s_cla32_pg_logic1_and0;
  wire [0:0] h_s_cla32_pg_logic1_xor0;
  wire [0:0] h_s_cla32_xor1;
  wire [0:0] h_s_cla32_and0;
  wire [0:0] h_s_cla32_or0;
  wire [0:0] h_s_cla32_pg_logic2_or0;
  wire [0:0] h_s_cla32_pg_logic2_and0;
  wire [0:0] h_s_cla32_pg_logic2_xor0;
  wire [0:0] h_s_cla32_xor2;
  wire [0:0] h_s_cla32_and1;
  wire [0:0] h_s_cla32_and2;
  wire [0:0] h_s_cla32_and3;
  wire [0:0] h_s_cla32_and4;
  wire [0:0] h_s_cla32_or1;
  wire [0:0] h_s_cla32_or2;
  wire [0:0] h_s_cla32_pg_logic3_or0;
  wire [0:0] h_s_cla32_pg_logic3_and0;
  wire [0:0] h_s_cla32_pg_logic3_xor0;
  wire [0:0] h_s_cla32_xor3;
  wire [0:0] h_s_cla32_and5;
  wire [0:0] h_s_cla32_and6;
  wire [0:0] h_s_cla32_and7;
  wire [0:0] h_s_cla32_and8;
  wire [0:0] h_s_cla32_and9;
  wire [0:0] h_s_cla32_and10;
  wire [0:0] h_s_cla32_and11;
  wire [0:0] h_s_cla32_or3;
  wire [0:0] h_s_cla32_or4;
  wire [0:0] h_s_cla32_or5;
  wire [0:0] h_s_cla32_pg_logic4_or0;
  wire [0:0] h_s_cla32_pg_logic4_and0;
  wire [0:0] h_s_cla32_pg_logic4_xor0;
  wire [0:0] h_s_cla32_xor4;
  wire [0:0] h_s_cla32_and12;
  wire [0:0] h_s_cla32_or6;
  wire [0:0] h_s_cla32_pg_logic5_or0;
  wire [0:0] h_s_cla32_pg_logic5_and0;
  wire [0:0] h_s_cla32_pg_logic5_xor0;
  wire [0:0] h_s_cla32_xor5;
  wire [0:0] h_s_cla32_and13;
  wire [0:0] h_s_cla32_and14;
  wire [0:0] h_s_cla32_and15;
  wire [0:0] h_s_cla32_or7;
  wire [0:0] h_s_cla32_or8;
  wire [0:0] h_s_cla32_pg_logic6_or0;
  wire [0:0] h_s_cla32_pg_logic6_and0;
  wire [0:0] h_s_cla32_pg_logic6_xor0;
  wire [0:0] h_s_cla32_xor6;
  wire [0:0] h_s_cla32_and16;
  wire [0:0] h_s_cla32_and17;
  wire [0:0] h_s_cla32_and18;
  wire [0:0] h_s_cla32_and19;
  wire [0:0] h_s_cla32_and20;
  wire [0:0] h_s_cla32_and21;
  wire [0:0] h_s_cla32_or9;
  wire [0:0] h_s_cla32_or10;
  wire [0:0] h_s_cla32_or11;
  wire [0:0] h_s_cla32_pg_logic7_or0;
  wire [0:0] h_s_cla32_pg_logic7_and0;
  wire [0:0] h_s_cla32_pg_logic7_xor0;
  wire [0:0] h_s_cla32_xor7;
  wire [0:0] h_s_cla32_and22;
  wire [0:0] h_s_cla32_and23;
  wire [0:0] h_s_cla32_and24;
  wire [0:0] h_s_cla32_and25;
  wire [0:0] h_s_cla32_and26;
  wire [0:0] h_s_cla32_and27;
  wire [0:0] h_s_cla32_and28;
  wire [0:0] h_s_cla32_and29;
  wire [0:0] h_s_cla32_and30;
  wire [0:0] h_s_cla32_and31;
  wire [0:0] h_s_cla32_or12;
  wire [0:0] h_s_cla32_or13;
  wire [0:0] h_s_cla32_or14;
  wire [0:0] h_s_cla32_or15;
  wire [0:0] h_s_cla32_pg_logic8_or0;
  wire [0:0] h_s_cla32_pg_logic8_and0;
  wire [0:0] h_s_cla32_pg_logic8_xor0;
  wire [0:0] h_s_cla32_xor8;
  wire [0:0] h_s_cla32_and32;
  wire [0:0] h_s_cla32_or16;
  wire [0:0] h_s_cla32_pg_logic9_or0;
  wire [0:0] h_s_cla32_pg_logic9_and0;
  wire [0:0] h_s_cla32_pg_logic9_xor0;
  wire [0:0] h_s_cla32_xor9;
  wire [0:0] h_s_cla32_and33;
  wire [0:0] h_s_cla32_and34;
  wire [0:0] h_s_cla32_and35;
  wire [0:0] h_s_cla32_or17;
  wire [0:0] h_s_cla32_or18;
  wire [0:0] h_s_cla32_pg_logic10_or0;
  wire [0:0] h_s_cla32_pg_logic10_and0;
  wire [0:0] h_s_cla32_pg_logic10_xor0;
  wire [0:0] h_s_cla32_xor10;
  wire [0:0] h_s_cla32_and36;
  wire [0:0] h_s_cla32_and37;
  wire [0:0] h_s_cla32_and38;
  wire [0:0] h_s_cla32_and39;
  wire [0:0] h_s_cla32_and40;
  wire [0:0] h_s_cla32_and41;
  wire [0:0] h_s_cla32_or19;
  wire [0:0] h_s_cla32_or20;
  wire [0:0] h_s_cla32_or21;
  wire [0:0] h_s_cla32_pg_logic11_or0;
  wire [0:0] h_s_cla32_pg_logic11_and0;
  wire [0:0] h_s_cla32_pg_logic11_xor0;
  wire [0:0] h_s_cla32_xor11;
  wire [0:0] h_s_cla32_and42;
  wire [0:0] h_s_cla32_and43;
  wire [0:0] h_s_cla32_and44;
  wire [0:0] h_s_cla32_and45;
  wire [0:0] h_s_cla32_and46;
  wire [0:0] h_s_cla32_and47;
  wire [0:0] h_s_cla32_and48;
  wire [0:0] h_s_cla32_and49;
  wire [0:0] h_s_cla32_and50;
  wire [0:0] h_s_cla32_and51;
  wire [0:0] h_s_cla32_or22;
  wire [0:0] h_s_cla32_or23;
  wire [0:0] h_s_cla32_or24;
  wire [0:0] h_s_cla32_or25;
  wire [0:0] h_s_cla32_pg_logic12_or0;
  wire [0:0] h_s_cla32_pg_logic12_and0;
  wire [0:0] h_s_cla32_pg_logic12_xor0;
  wire [0:0] h_s_cla32_xor12;
  wire [0:0] h_s_cla32_and52;
  wire [0:0] h_s_cla32_or26;
  wire [0:0] h_s_cla32_pg_logic13_or0;
  wire [0:0] h_s_cla32_pg_logic13_and0;
  wire [0:0] h_s_cla32_pg_logic13_xor0;
  wire [0:0] h_s_cla32_xor13;
  wire [0:0] h_s_cla32_and53;
  wire [0:0] h_s_cla32_and54;
  wire [0:0] h_s_cla32_and55;
  wire [0:0] h_s_cla32_or27;
  wire [0:0] h_s_cla32_or28;
  wire [0:0] h_s_cla32_pg_logic14_or0;
  wire [0:0] h_s_cla32_pg_logic14_and0;
  wire [0:0] h_s_cla32_pg_logic14_xor0;
  wire [0:0] h_s_cla32_xor14;
  wire [0:0] h_s_cla32_and56;
  wire [0:0] h_s_cla32_and57;
  wire [0:0] h_s_cla32_and58;
  wire [0:0] h_s_cla32_and59;
  wire [0:0] h_s_cla32_and60;
  wire [0:0] h_s_cla32_and61;
  wire [0:0] h_s_cla32_or29;
  wire [0:0] h_s_cla32_or30;
  wire [0:0] h_s_cla32_or31;
  wire [0:0] h_s_cla32_pg_logic15_or0;
  wire [0:0] h_s_cla32_pg_logic15_and0;
  wire [0:0] h_s_cla32_pg_logic15_xor0;
  wire [0:0] h_s_cla32_xor15;
  wire [0:0] h_s_cla32_and62;
  wire [0:0] h_s_cla32_and63;
  wire [0:0] h_s_cla32_and64;
  wire [0:0] h_s_cla32_and65;
  wire [0:0] h_s_cla32_and66;
  wire [0:0] h_s_cla32_and67;
  wire [0:0] h_s_cla32_and68;
  wire [0:0] h_s_cla32_and69;
  wire [0:0] h_s_cla32_and70;
  wire [0:0] h_s_cla32_and71;
  wire [0:0] h_s_cla32_or32;
  wire [0:0] h_s_cla32_or33;
  wire [0:0] h_s_cla32_or34;
  wire [0:0] h_s_cla32_or35;
  wire [0:0] h_s_cla32_pg_logic16_or0;
  wire [0:0] h_s_cla32_pg_logic16_and0;
  wire [0:0] h_s_cla32_pg_logic16_xor0;
  wire [0:0] h_s_cla32_xor16;
  wire [0:0] h_s_cla32_and72;
  wire [0:0] h_s_cla32_or36;
  wire [0:0] h_s_cla32_pg_logic17_or0;
  wire [0:0] h_s_cla32_pg_logic17_and0;
  wire [0:0] h_s_cla32_pg_logic17_xor0;
  wire [0:0] h_s_cla32_xor17;
  wire [0:0] h_s_cla32_and73;
  wire [0:0] h_s_cla32_and74;
  wire [0:0] h_s_cla32_and75;
  wire [0:0] h_s_cla32_or37;
  wire [0:0] h_s_cla32_or38;
  wire [0:0] h_s_cla32_pg_logic18_or0;
  wire [0:0] h_s_cla32_pg_logic18_and0;
  wire [0:0] h_s_cla32_pg_logic18_xor0;
  wire [0:0] h_s_cla32_xor18;
  wire [0:0] h_s_cla32_and76;
  wire [0:0] h_s_cla32_and77;
  wire [0:0] h_s_cla32_and78;
  wire [0:0] h_s_cla32_and79;
  wire [0:0] h_s_cla32_and80;
  wire [0:0] h_s_cla32_and81;
  wire [0:0] h_s_cla32_or39;
  wire [0:0] h_s_cla32_or40;
  wire [0:0] h_s_cla32_or41;
  wire [0:0] h_s_cla32_pg_logic19_or0;
  wire [0:0] h_s_cla32_pg_logic19_and0;
  wire [0:0] h_s_cla32_pg_logic19_xor0;
  wire [0:0] h_s_cla32_xor19;
  wire [0:0] h_s_cla32_and82;
  wire [0:0] h_s_cla32_and83;
  wire [0:0] h_s_cla32_and84;
  wire [0:0] h_s_cla32_and85;
  wire [0:0] h_s_cla32_and86;
  wire [0:0] h_s_cla32_and87;
  wire [0:0] h_s_cla32_and88;
  wire [0:0] h_s_cla32_and89;
  wire [0:0] h_s_cla32_and90;
  wire [0:0] h_s_cla32_and91;
  wire [0:0] h_s_cla32_or42;
  wire [0:0] h_s_cla32_or43;
  wire [0:0] h_s_cla32_or44;
  wire [0:0] h_s_cla32_or45;
  wire [0:0] h_s_cla32_pg_logic20_or0;
  wire [0:0] h_s_cla32_pg_logic20_and0;
  wire [0:0] h_s_cla32_pg_logic20_xor0;
  wire [0:0] h_s_cla32_xor20;
  wire [0:0] h_s_cla32_and92;
  wire [0:0] h_s_cla32_or46;
  wire [0:0] h_s_cla32_pg_logic21_or0;
  wire [0:0] h_s_cla32_pg_logic21_and0;
  wire [0:0] h_s_cla32_pg_logic21_xor0;
  wire [0:0] h_s_cla32_xor21;
  wire [0:0] h_s_cla32_and93;
  wire [0:0] h_s_cla32_and94;
  wire [0:0] h_s_cla32_and95;
  wire [0:0] h_s_cla32_or47;
  wire [0:0] h_s_cla32_or48;
  wire [0:0] h_s_cla32_pg_logic22_or0;
  wire [0:0] h_s_cla32_pg_logic22_and0;
  wire [0:0] h_s_cla32_pg_logic22_xor0;
  wire [0:0] h_s_cla32_xor22;
  wire [0:0] h_s_cla32_and96;
  wire [0:0] h_s_cla32_and97;
  wire [0:0] h_s_cla32_and98;
  wire [0:0] h_s_cla32_and99;
  wire [0:0] h_s_cla32_and100;
  wire [0:0] h_s_cla32_and101;
  wire [0:0] h_s_cla32_or49;
  wire [0:0] h_s_cla32_or50;
  wire [0:0] h_s_cla32_or51;
  wire [0:0] h_s_cla32_pg_logic23_or0;
  wire [0:0] h_s_cla32_pg_logic23_and0;
  wire [0:0] h_s_cla32_pg_logic23_xor0;
  wire [0:0] h_s_cla32_xor23;
  wire [0:0] h_s_cla32_and102;
  wire [0:0] h_s_cla32_and103;
  wire [0:0] h_s_cla32_and104;
  wire [0:0] h_s_cla32_and105;
  wire [0:0] h_s_cla32_and106;
  wire [0:0] h_s_cla32_and107;
  wire [0:0] h_s_cla32_and108;
  wire [0:0] h_s_cla32_and109;
  wire [0:0] h_s_cla32_and110;
  wire [0:0] h_s_cla32_and111;
  wire [0:0] h_s_cla32_or52;
  wire [0:0] h_s_cla32_or53;
  wire [0:0] h_s_cla32_or54;
  wire [0:0] h_s_cla32_or55;
  wire [0:0] h_s_cla32_pg_logic24_or0;
  wire [0:0] h_s_cla32_pg_logic24_and0;
  wire [0:0] h_s_cla32_pg_logic24_xor0;
  wire [0:0] h_s_cla32_xor24;
  wire [0:0] h_s_cla32_and112;
  wire [0:0] h_s_cla32_or56;
  wire [0:0] h_s_cla32_pg_logic25_or0;
  wire [0:0] h_s_cla32_pg_logic25_and0;
  wire [0:0] h_s_cla32_pg_logic25_xor0;
  wire [0:0] h_s_cla32_xor25;
  wire [0:0] h_s_cla32_and113;
  wire [0:0] h_s_cla32_and114;
  wire [0:0] h_s_cla32_and115;
  wire [0:0] h_s_cla32_or57;
  wire [0:0] h_s_cla32_or58;
  wire [0:0] h_s_cla32_pg_logic26_or0;
  wire [0:0] h_s_cla32_pg_logic26_and0;
  wire [0:0] h_s_cla32_pg_logic26_xor0;
  wire [0:0] h_s_cla32_xor26;
  wire [0:0] h_s_cla32_and116;
  wire [0:0] h_s_cla32_and117;
  wire [0:0] h_s_cla32_and118;
  wire [0:0] h_s_cla32_and119;
  wire [0:0] h_s_cla32_and120;
  wire [0:0] h_s_cla32_and121;
  wire [0:0] h_s_cla32_or59;
  wire [0:0] h_s_cla32_or60;
  wire [0:0] h_s_cla32_or61;
  wire [0:0] h_s_cla32_pg_logic27_or0;
  wire [0:0] h_s_cla32_pg_logic27_and0;
  wire [0:0] h_s_cla32_pg_logic27_xor0;
  wire [0:0] h_s_cla32_xor27;
  wire [0:0] h_s_cla32_and122;
  wire [0:0] h_s_cla32_and123;
  wire [0:0] h_s_cla32_and124;
  wire [0:0] h_s_cla32_and125;
  wire [0:0] h_s_cla32_and126;
  wire [0:0] h_s_cla32_and127;
  wire [0:0] h_s_cla32_and128;
  wire [0:0] h_s_cla32_and129;
  wire [0:0] h_s_cla32_and130;
  wire [0:0] h_s_cla32_and131;
  wire [0:0] h_s_cla32_or62;
  wire [0:0] h_s_cla32_or63;
  wire [0:0] h_s_cla32_or64;
  wire [0:0] h_s_cla32_or65;
  wire [0:0] h_s_cla32_pg_logic28_or0;
  wire [0:0] h_s_cla32_pg_logic28_and0;
  wire [0:0] h_s_cla32_pg_logic28_xor0;
  wire [0:0] h_s_cla32_xor28;
  wire [0:0] h_s_cla32_and132;
  wire [0:0] h_s_cla32_or66;
  wire [0:0] h_s_cla32_pg_logic29_or0;
  wire [0:0] h_s_cla32_pg_logic29_and0;
  wire [0:0] h_s_cla32_pg_logic29_xor0;
  wire [0:0] h_s_cla32_xor29;
  wire [0:0] h_s_cla32_and133;
  wire [0:0] h_s_cla32_and134;
  wire [0:0] h_s_cla32_and135;
  wire [0:0] h_s_cla32_or67;
  wire [0:0] h_s_cla32_or68;
  wire [0:0] h_s_cla32_pg_logic30_or0;
  wire [0:0] h_s_cla32_pg_logic30_and0;
  wire [0:0] h_s_cla32_pg_logic30_xor0;
  wire [0:0] h_s_cla32_xor30;
  wire [0:0] h_s_cla32_and136;
  wire [0:0] h_s_cla32_and137;
  wire [0:0] h_s_cla32_and138;
  wire [0:0] h_s_cla32_and139;
  wire [0:0] h_s_cla32_and140;
  wire [0:0] h_s_cla32_and141;
  wire [0:0] h_s_cla32_or69;
  wire [0:0] h_s_cla32_or70;
  wire [0:0] h_s_cla32_or71;
  wire [0:0] h_s_cla32_pg_logic31_or0;
  wire [0:0] h_s_cla32_pg_logic31_and0;
  wire [0:0] h_s_cla32_pg_logic31_xor0;
  wire [0:0] h_s_cla32_xor31;
  wire [0:0] h_s_cla32_and142;
  wire [0:0] h_s_cla32_and143;
  wire [0:0] h_s_cla32_and144;
  wire [0:0] h_s_cla32_and145;
  wire [0:0] h_s_cla32_and146;
  wire [0:0] h_s_cla32_and147;
  wire [0:0] h_s_cla32_and148;
  wire [0:0] h_s_cla32_and149;
  wire [0:0] h_s_cla32_and150;
  wire [0:0] h_s_cla32_and151;
  wire [0:0] h_s_cla32_or72;
  wire [0:0] h_s_cla32_or73;
  wire [0:0] h_s_cla32_or74;
  wire [0:0] h_s_cla32_or75;
  wire [0:0] h_s_cla32_xor32;
  wire [0:0] h_s_cla32_xor33;

  pg_logic pg_logic_h_s_cla32_pg_logic0_out(.a(a[0]), .b(b[0]), .pg_logic_or0(h_s_cla32_pg_logic0_or0), .pg_logic_and0(h_s_cla32_pg_logic0_and0), .pg_logic_xor0(h_s_cla32_pg_logic0_xor0));
  pg_logic pg_logic_h_s_cla32_pg_logic1_out(.a(a[1]), .b(b[1]), .pg_logic_or0(h_s_cla32_pg_logic1_or0), .pg_logic_and0(h_s_cla32_pg_logic1_and0), .pg_logic_xor0(h_s_cla32_pg_logic1_xor0));
  xor_gate xor_gate_h_s_cla32_xor1(.a(h_s_cla32_pg_logic1_xor0[0]), .b(h_s_cla32_pg_logic0_and0[0]), .out(h_s_cla32_xor1));
  and_gate and_gate_h_s_cla32_and0(.a(h_s_cla32_pg_logic0_and0[0]), .b(h_s_cla32_pg_logic1_or0[0]), .out(h_s_cla32_and0));
  or_gate or_gate_h_s_cla32_or0(.a(h_s_cla32_pg_logic1_and0[0]), .b(h_s_cla32_and0[0]), .out(h_s_cla32_or0));
  pg_logic pg_logic_h_s_cla32_pg_logic2_out(.a(a[2]), .b(b[2]), .pg_logic_or0(h_s_cla32_pg_logic2_or0), .pg_logic_and0(h_s_cla32_pg_logic2_and0), .pg_logic_xor0(h_s_cla32_pg_logic2_xor0));
  xor_gate xor_gate_h_s_cla32_xor2(.a(h_s_cla32_pg_logic2_xor0[0]), .b(h_s_cla32_or0[0]), .out(h_s_cla32_xor2));
  and_gate and_gate_h_s_cla32_and1(.a(h_s_cla32_pg_logic2_or0[0]), .b(h_s_cla32_pg_logic0_or0[0]), .out(h_s_cla32_and1));
  and_gate and_gate_h_s_cla32_and2(.a(h_s_cla32_pg_logic0_and0[0]), .b(h_s_cla32_pg_logic2_or0[0]), .out(h_s_cla32_and2));
  and_gate and_gate_h_s_cla32_and3(.a(h_s_cla32_and2[0]), .b(h_s_cla32_pg_logic1_or0[0]), .out(h_s_cla32_and3));
  and_gate and_gate_h_s_cla32_and4(.a(h_s_cla32_pg_logic1_and0[0]), .b(h_s_cla32_pg_logic2_or0[0]), .out(h_s_cla32_and4));
  or_gate or_gate_h_s_cla32_or1(.a(h_s_cla32_and3[0]), .b(h_s_cla32_and4[0]), .out(h_s_cla32_or1));
  or_gate or_gate_h_s_cla32_or2(.a(h_s_cla32_pg_logic2_and0[0]), .b(h_s_cla32_or1[0]), .out(h_s_cla32_or2));
  pg_logic pg_logic_h_s_cla32_pg_logic3_out(.a(a[3]), .b(b[3]), .pg_logic_or0(h_s_cla32_pg_logic3_or0), .pg_logic_and0(h_s_cla32_pg_logic3_and0), .pg_logic_xor0(h_s_cla32_pg_logic3_xor0));
  xor_gate xor_gate_h_s_cla32_xor3(.a(h_s_cla32_pg_logic3_xor0[0]), .b(h_s_cla32_or2[0]), .out(h_s_cla32_xor3));
  and_gate and_gate_h_s_cla32_and5(.a(h_s_cla32_pg_logic3_or0[0]), .b(h_s_cla32_pg_logic1_or0[0]), .out(h_s_cla32_and5));
  and_gate and_gate_h_s_cla32_and6(.a(h_s_cla32_pg_logic0_and0[0]), .b(h_s_cla32_pg_logic2_or0[0]), .out(h_s_cla32_and6));
  and_gate and_gate_h_s_cla32_and7(.a(h_s_cla32_pg_logic3_or0[0]), .b(h_s_cla32_pg_logic1_or0[0]), .out(h_s_cla32_and7));
  and_gate and_gate_h_s_cla32_and8(.a(h_s_cla32_and6[0]), .b(h_s_cla32_and7[0]), .out(h_s_cla32_and8));
  and_gate and_gate_h_s_cla32_and9(.a(h_s_cla32_pg_logic1_and0[0]), .b(h_s_cla32_pg_logic3_or0[0]), .out(h_s_cla32_and9));
  and_gate and_gate_h_s_cla32_and10(.a(h_s_cla32_and9[0]), .b(h_s_cla32_pg_logic2_or0[0]), .out(h_s_cla32_and10));
  and_gate and_gate_h_s_cla32_and11(.a(h_s_cla32_pg_logic2_and0[0]), .b(h_s_cla32_pg_logic3_or0[0]), .out(h_s_cla32_and11));
  or_gate or_gate_h_s_cla32_or3(.a(h_s_cla32_and8[0]), .b(h_s_cla32_and11[0]), .out(h_s_cla32_or3));
  or_gate or_gate_h_s_cla32_or4(.a(h_s_cla32_and10[0]), .b(h_s_cla32_or3[0]), .out(h_s_cla32_or4));
  or_gate or_gate_h_s_cla32_or5(.a(h_s_cla32_pg_logic3_and0[0]), .b(h_s_cla32_or4[0]), .out(h_s_cla32_or5));
  pg_logic pg_logic_h_s_cla32_pg_logic4_out(.a(a[4]), .b(b[4]), .pg_logic_or0(h_s_cla32_pg_logic4_or0), .pg_logic_and0(h_s_cla32_pg_logic4_and0), .pg_logic_xor0(h_s_cla32_pg_logic4_xor0));
  xor_gate xor_gate_h_s_cla32_xor4(.a(h_s_cla32_pg_logic4_xor0[0]), .b(h_s_cla32_or5[0]), .out(h_s_cla32_xor4));
  and_gate and_gate_h_s_cla32_and12(.a(h_s_cla32_or5[0]), .b(h_s_cla32_pg_logic4_or0[0]), .out(h_s_cla32_and12));
  or_gate or_gate_h_s_cla32_or6(.a(h_s_cla32_pg_logic4_and0[0]), .b(h_s_cla32_and12[0]), .out(h_s_cla32_or6));
  pg_logic pg_logic_h_s_cla32_pg_logic5_out(.a(a[5]), .b(b[5]), .pg_logic_or0(h_s_cla32_pg_logic5_or0), .pg_logic_and0(h_s_cla32_pg_logic5_and0), .pg_logic_xor0(h_s_cla32_pg_logic5_xor0));
  xor_gate xor_gate_h_s_cla32_xor5(.a(h_s_cla32_pg_logic5_xor0[0]), .b(h_s_cla32_or6[0]), .out(h_s_cla32_xor5));
  and_gate and_gate_h_s_cla32_and13(.a(h_s_cla32_or5[0]), .b(h_s_cla32_pg_logic5_or0[0]), .out(h_s_cla32_and13));
  and_gate and_gate_h_s_cla32_and14(.a(h_s_cla32_and13[0]), .b(h_s_cla32_pg_logic4_or0[0]), .out(h_s_cla32_and14));
  and_gate and_gate_h_s_cla32_and15(.a(h_s_cla32_pg_logic4_and0[0]), .b(h_s_cla32_pg_logic5_or0[0]), .out(h_s_cla32_and15));
  or_gate or_gate_h_s_cla32_or7(.a(h_s_cla32_and14[0]), .b(h_s_cla32_and15[0]), .out(h_s_cla32_or7));
  or_gate or_gate_h_s_cla32_or8(.a(h_s_cla32_pg_logic5_and0[0]), .b(h_s_cla32_or7[0]), .out(h_s_cla32_or8));
  pg_logic pg_logic_h_s_cla32_pg_logic6_out(.a(a[6]), .b(b[6]), .pg_logic_or0(h_s_cla32_pg_logic6_or0), .pg_logic_and0(h_s_cla32_pg_logic6_and0), .pg_logic_xor0(h_s_cla32_pg_logic6_xor0));
  xor_gate xor_gate_h_s_cla32_xor6(.a(h_s_cla32_pg_logic6_xor0[0]), .b(h_s_cla32_or8[0]), .out(h_s_cla32_xor6));
  and_gate and_gate_h_s_cla32_and16(.a(h_s_cla32_or5[0]), .b(h_s_cla32_pg_logic5_or0[0]), .out(h_s_cla32_and16));
  and_gate and_gate_h_s_cla32_and17(.a(h_s_cla32_pg_logic6_or0[0]), .b(h_s_cla32_pg_logic4_or0[0]), .out(h_s_cla32_and17));
  and_gate and_gate_h_s_cla32_and18(.a(h_s_cla32_and16[0]), .b(h_s_cla32_and17[0]), .out(h_s_cla32_and18));
  and_gate and_gate_h_s_cla32_and19(.a(h_s_cla32_pg_logic4_and0[0]), .b(h_s_cla32_pg_logic6_or0[0]), .out(h_s_cla32_and19));
  and_gate and_gate_h_s_cla32_and20(.a(h_s_cla32_and19[0]), .b(h_s_cla32_pg_logic5_or0[0]), .out(h_s_cla32_and20));
  and_gate and_gate_h_s_cla32_and21(.a(h_s_cla32_pg_logic5_and0[0]), .b(h_s_cla32_pg_logic6_or0[0]), .out(h_s_cla32_and21));
  or_gate or_gate_h_s_cla32_or9(.a(h_s_cla32_and18[0]), .b(h_s_cla32_and20[0]), .out(h_s_cla32_or9));
  or_gate or_gate_h_s_cla32_or10(.a(h_s_cla32_or9[0]), .b(h_s_cla32_and21[0]), .out(h_s_cla32_or10));
  or_gate or_gate_h_s_cla32_or11(.a(h_s_cla32_pg_logic6_and0[0]), .b(h_s_cla32_or10[0]), .out(h_s_cla32_or11));
  pg_logic pg_logic_h_s_cla32_pg_logic7_out(.a(a[7]), .b(b[7]), .pg_logic_or0(h_s_cla32_pg_logic7_or0), .pg_logic_and0(h_s_cla32_pg_logic7_and0), .pg_logic_xor0(h_s_cla32_pg_logic7_xor0));
  xor_gate xor_gate_h_s_cla32_xor7(.a(h_s_cla32_pg_logic7_xor0[0]), .b(h_s_cla32_or11[0]), .out(h_s_cla32_xor7));
  and_gate and_gate_h_s_cla32_and22(.a(h_s_cla32_or5[0]), .b(h_s_cla32_pg_logic6_or0[0]), .out(h_s_cla32_and22));
  and_gate and_gate_h_s_cla32_and23(.a(h_s_cla32_pg_logic7_or0[0]), .b(h_s_cla32_pg_logic5_or0[0]), .out(h_s_cla32_and23));
  and_gate and_gate_h_s_cla32_and24(.a(h_s_cla32_and22[0]), .b(h_s_cla32_and23[0]), .out(h_s_cla32_and24));
  and_gate and_gate_h_s_cla32_and25(.a(h_s_cla32_and24[0]), .b(h_s_cla32_pg_logic4_or0[0]), .out(h_s_cla32_and25));
  and_gate and_gate_h_s_cla32_and26(.a(h_s_cla32_pg_logic4_and0[0]), .b(h_s_cla32_pg_logic6_or0[0]), .out(h_s_cla32_and26));
  and_gate and_gate_h_s_cla32_and27(.a(h_s_cla32_pg_logic7_or0[0]), .b(h_s_cla32_pg_logic5_or0[0]), .out(h_s_cla32_and27));
  and_gate and_gate_h_s_cla32_and28(.a(h_s_cla32_and26[0]), .b(h_s_cla32_and27[0]), .out(h_s_cla32_and28));
  and_gate and_gate_h_s_cla32_and29(.a(h_s_cla32_pg_logic5_and0[0]), .b(h_s_cla32_pg_logic7_or0[0]), .out(h_s_cla32_and29));
  and_gate and_gate_h_s_cla32_and30(.a(h_s_cla32_and29[0]), .b(h_s_cla32_pg_logic6_or0[0]), .out(h_s_cla32_and30));
  and_gate and_gate_h_s_cla32_and31(.a(h_s_cla32_pg_logic6_and0[0]), .b(h_s_cla32_pg_logic7_or0[0]), .out(h_s_cla32_and31));
  or_gate or_gate_h_s_cla32_or12(.a(h_s_cla32_and25[0]), .b(h_s_cla32_and30[0]), .out(h_s_cla32_or12));
  or_gate or_gate_h_s_cla32_or13(.a(h_s_cla32_and28[0]), .b(h_s_cla32_and31[0]), .out(h_s_cla32_or13));
  or_gate or_gate_h_s_cla32_or14(.a(h_s_cla32_or12[0]), .b(h_s_cla32_or13[0]), .out(h_s_cla32_or14));
  or_gate or_gate_h_s_cla32_or15(.a(h_s_cla32_pg_logic7_and0[0]), .b(h_s_cla32_or14[0]), .out(h_s_cla32_or15));
  pg_logic pg_logic_h_s_cla32_pg_logic8_out(.a(a[8]), .b(b[8]), .pg_logic_or0(h_s_cla32_pg_logic8_or0), .pg_logic_and0(h_s_cla32_pg_logic8_and0), .pg_logic_xor0(h_s_cla32_pg_logic8_xor0));
  xor_gate xor_gate_h_s_cla32_xor8(.a(h_s_cla32_pg_logic8_xor0[0]), .b(h_s_cla32_or15[0]), .out(h_s_cla32_xor8));
  and_gate and_gate_h_s_cla32_and32(.a(h_s_cla32_or15[0]), .b(h_s_cla32_pg_logic8_or0[0]), .out(h_s_cla32_and32));
  or_gate or_gate_h_s_cla32_or16(.a(h_s_cla32_pg_logic8_and0[0]), .b(h_s_cla32_and32[0]), .out(h_s_cla32_or16));
  pg_logic pg_logic_h_s_cla32_pg_logic9_out(.a(a[9]), .b(b[9]), .pg_logic_or0(h_s_cla32_pg_logic9_or0), .pg_logic_and0(h_s_cla32_pg_logic9_and0), .pg_logic_xor0(h_s_cla32_pg_logic9_xor0));
  xor_gate xor_gate_h_s_cla32_xor9(.a(h_s_cla32_pg_logic9_xor0[0]), .b(h_s_cla32_or16[0]), .out(h_s_cla32_xor9));
  and_gate and_gate_h_s_cla32_and33(.a(h_s_cla32_or15[0]), .b(h_s_cla32_pg_logic9_or0[0]), .out(h_s_cla32_and33));
  and_gate and_gate_h_s_cla32_and34(.a(h_s_cla32_and33[0]), .b(h_s_cla32_pg_logic8_or0[0]), .out(h_s_cla32_and34));
  and_gate and_gate_h_s_cla32_and35(.a(h_s_cla32_pg_logic8_and0[0]), .b(h_s_cla32_pg_logic9_or0[0]), .out(h_s_cla32_and35));
  or_gate or_gate_h_s_cla32_or17(.a(h_s_cla32_and34[0]), .b(h_s_cla32_and35[0]), .out(h_s_cla32_or17));
  or_gate or_gate_h_s_cla32_or18(.a(h_s_cla32_pg_logic9_and0[0]), .b(h_s_cla32_or17[0]), .out(h_s_cla32_or18));
  pg_logic pg_logic_h_s_cla32_pg_logic10_out(.a(a[10]), .b(b[10]), .pg_logic_or0(h_s_cla32_pg_logic10_or0), .pg_logic_and0(h_s_cla32_pg_logic10_and0), .pg_logic_xor0(h_s_cla32_pg_logic10_xor0));
  xor_gate xor_gate_h_s_cla32_xor10(.a(h_s_cla32_pg_logic10_xor0[0]), .b(h_s_cla32_or18[0]), .out(h_s_cla32_xor10));
  and_gate and_gate_h_s_cla32_and36(.a(h_s_cla32_or15[0]), .b(h_s_cla32_pg_logic9_or0[0]), .out(h_s_cla32_and36));
  and_gate and_gate_h_s_cla32_and37(.a(h_s_cla32_pg_logic10_or0[0]), .b(h_s_cla32_pg_logic8_or0[0]), .out(h_s_cla32_and37));
  and_gate and_gate_h_s_cla32_and38(.a(h_s_cla32_and36[0]), .b(h_s_cla32_and37[0]), .out(h_s_cla32_and38));
  and_gate and_gate_h_s_cla32_and39(.a(h_s_cla32_pg_logic8_and0[0]), .b(h_s_cla32_pg_logic10_or0[0]), .out(h_s_cla32_and39));
  and_gate and_gate_h_s_cla32_and40(.a(h_s_cla32_and39[0]), .b(h_s_cla32_pg_logic9_or0[0]), .out(h_s_cla32_and40));
  and_gate and_gate_h_s_cla32_and41(.a(h_s_cla32_pg_logic9_and0[0]), .b(h_s_cla32_pg_logic10_or0[0]), .out(h_s_cla32_and41));
  or_gate or_gate_h_s_cla32_or19(.a(h_s_cla32_and38[0]), .b(h_s_cla32_and40[0]), .out(h_s_cla32_or19));
  or_gate or_gate_h_s_cla32_or20(.a(h_s_cla32_or19[0]), .b(h_s_cla32_and41[0]), .out(h_s_cla32_or20));
  or_gate or_gate_h_s_cla32_or21(.a(h_s_cla32_pg_logic10_and0[0]), .b(h_s_cla32_or20[0]), .out(h_s_cla32_or21));
  pg_logic pg_logic_h_s_cla32_pg_logic11_out(.a(a[11]), .b(b[11]), .pg_logic_or0(h_s_cla32_pg_logic11_or0), .pg_logic_and0(h_s_cla32_pg_logic11_and0), .pg_logic_xor0(h_s_cla32_pg_logic11_xor0));
  xor_gate xor_gate_h_s_cla32_xor11(.a(h_s_cla32_pg_logic11_xor0[0]), .b(h_s_cla32_or21[0]), .out(h_s_cla32_xor11));
  and_gate and_gate_h_s_cla32_and42(.a(h_s_cla32_or15[0]), .b(h_s_cla32_pg_logic10_or0[0]), .out(h_s_cla32_and42));
  and_gate and_gate_h_s_cla32_and43(.a(h_s_cla32_pg_logic11_or0[0]), .b(h_s_cla32_pg_logic9_or0[0]), .out(h_s_cla32_and43));
  and_gate and_gate_h_s_cla32_and44(.a(h_s_cla32_and42[0]), .b(h_s_cla32_and43[0]), .out(h_s_cla32_and44));
  and_gate and_gate_h_s_cla32_and45(.a(h_s_cla32_and44[0]), .b(h_s_cla32_pg_logic8_or0[0]), .out(h_s_cla32_and45));
  and_gate and_gate_h_s_cla32_and46(.a(h_s_cla32_pg_logic8_and0[0]), .b(h_s_cla32_pg_logic10_or0[0]), .out(h_s_cla32_and46));
  and_gate and_gate_h_s_cla32_and47(.a(h_s_cla32_pg_logic11_or0[0]), .b(h_s_cla32_pg_logic9_or0[0]), .out(h_s_cla32_and47));
  and_gate and_gate_h_s_cla32_and48(.a(h_s_cla32_and46[0]), .b(h_s_cla32_and47[0]), .out(h_s_cla32_and48));
  and_gate and_gate_h_s_cla32_and49(.a(h_s_cla32_pg_logic9_and0[0]), .b(h_s_cla32_pg_logic11_or0[0]), .out(h_s_cla32_and49));
  and_gate and_gate_h_s_cla32_and50(.a(h_s_cla32_and49[0]), .b(h_s_cla32_pg_logic10_or0[0]), .out(h_s_cla32_and50));
  and_gate and_gate_h_s_cla32_and51(.a(h_s_cla32_pg_logic10_and0[0]), .b(h_s_cla32_pg_logic11_or0[0]), .out(h_s_cla32_and51));
  or_gate or_gate_h_s_cla32_or22(.a(h_s_cla32_and45[0]), .b(h_s_cla32_and50[0]), .out(h_s_cla32_or22));
  or_gate or_gate_h_s_cla32_or23(.a(h_s_cla32_and48[0]), .b(h_s_cla32_and51[0]), .out(h_s_cla32_or23));
  or_gate or_gate_h_s_cla32_or24(.a(h_s_cla32_or22[0]), .b(h_s_cla32_or23[0]), .out(h_s_cla32_or24));
  or_gate or_gate_h_s_cla32_or25(.a(h_s_cla32_pg_logic11_and0[0]), .b(h_s_cla32_or24[0]), .out(h_s_cla32_or25));
  pg_logic pg_logic_h_s_cla32_pg_logic12_out(.a(a[12]), .b(b[12]), .pg_logic_or0(h_s_cla32_pg_logic12_or0), .pg_logic_and0(h_s_cla32_pg_logic12_and0), .pg_logic_xor0(h_s_cla32_pg_logic12_xor0));
  xor_gate xor_gate_h_s_cla32_xor12(.a(h_s_cla32_pg_logic12_xor0[0]), .b(h_s_cla32_or25[0]), .out(h_s_cla32_xor12));
  and_gate and_gate_h_s_cla32_and52(.a(h_s_cla32_or25[0]), .b(h_s_cla32_pg_logic12_or0[0]), .out(h_s_cla32_and52));
  or_gate or_gate_h_s_cla32_or26(.a(h_s_cla32_pg_logic12_and0[0]), .b(h_s_cla32_and52[0]), .out(h_s_cla32_or26));
  pg_logic pg_logic_h_s_cla32_pg_logic13_out(.a(a[13]), .b(b[13]), .pg_logic_or0(h_s_cla32_pg_logic13_or0), .pg_logic_and0(h_s_cla32_pg_logic13_and0), .pg_logic_xor0(h_s_cla32_pg_logic13_xor0));
  xor_gate xor_gate_h_s_cla32_xor13(.a(h_s_cla32_pg_logic13_xor0[0]), .b(h_s_cla32_or26[0]), .out(h_s_cla32_xor13));
  and_gate and_gate_h_s_cla32_and53(.a(h_s_cla32_or25[0]), .b(h_s_cla32_pg_logic13_or0[0]), .out(h_s_cla32_and53));
  and_gate and_gate_h_s_cla32_and54(.a(h_s_cla32_and53[0]), .b(h_s_cla32_pg_logic12_or0[0]), .out(h_s_cla32_and54));
  and_gate and_gate_h_s_cla32_and55(.a(h_s_cla32_pg_logic12_and0[0]), .b(h_s_cla32_pg_logic13_or0[0]), .out(h_s_cla32_and55));
  or_gate or_gate_h_s_cla32_or27(.a(h_s_cla32_and54[0]), .b(h_s_cla32_and55[0]), .out(h_s_cla32_or27));
  or_gate or_gate_h_s_cla32_or28(.a(h_s_cla32_pg_logic13_and0[0]), .b(h_s_cla32_or27[0]), .out(h_s_cla32_or28));
  pg_logic pg_logic_h_s_cla32_pg_logic14_out(.a(a[14]), .b(b[14]), .pg_logic_or0(h_s_cla32_pg_logic14_or0), .pg_logic_and0(h_s_cla32_pg_logic14_and0), .pg_logic_xor0(h_s_cla32_pg_logic14_xor0));
  xor_gate xor_gate_h_s_cla32_xor14(.a(h_s_cla32_pg_logic14_xor0[0]), .b(h_s_cla32_or28[0]), .out(h_s_cla32_xor14));
  and_gate and_gate_h_s_cla32_and56(.a(h_s_cla32_or25[0]), .b(h_s_cla32_pg_logic13_or0[0]), .out(h_s_cla32_and56));
  and_gate and_gate_h_s_cla32_and57(.a(h_s_cla32_pg_logic14_or0[0]), .b(h_s_cla32_pg_logic12_or0[0]), .out(h_s_cla32_and57));
  and_gate and_gate_h_s_cla32_and58(.a(h_s_cla32_and56[0]), .b(h_s_cla32_and57[0]), .out(h_s_cla32_and58));
  and_gate and_gate_h_s_cla32_and59(.a(h_s_cla32_pg_logic12_and0[0]), .b(h_s_cla32_pg_logic14_or0[0]), .out(h_s_cla32_and59));
  and_gate and_gate_h_s_cla32_and60(.a(h_s_cla32_and59[0]), .b(h_s_cla32_pg_logic13_or0[0]), .out(h_s_cla32_and60));
  and_gate and_gate_h_s_cla32_and61(.a(h_s_cla32_pg_logic13_and0[0]), .b(h_s_cla32_pg_logic14_or0[0]), .out(h_s_cla32_and61));
  or_gate or_gate_h_s_cla32_or29(.a(h_s_cla32_and58[0]), .b(h_s_cla32_and60[0]), .out(h_s_cla32_or29));
  or_gate or_gate_h_s_cla32_or30(.a(h_s_cla32_or29[0]), .b(h_s_cla32_and61[0]), .out(h_s_cla32_or30));
  or_gate or_gate_h_s_cla32_or31(.a(h_s_cla32_pg_logic14_and0[0]), .b(h_s_cla32_or30[0]), .out(h_s_cla32_or31));
  pg_logic pg_logic_h_s_cla32_pg_logic15_out(.a(a[15]), .b(b[15]), .pg_logic_or0(h_s_cla32_pg_logic15_or0), .pg_logic_and0(h_s_cla32_pg_logic15_and0), .pg_logic_xor0(h_s_cla32_pg_logic15_xor0));
  xor_gate xor_gate_h_s_cla32_xor15(.a(h_s_cla32_pg_logic15_xor0[0]), .b(h_s_cla32_or31[0]), .out(h_s_cla32_xor15));
  and_gate and_gate_h_s_cla32_and62(.a(h_s_cla32_or25[0]), .b(h_s_cla32_pg_logic14_or0[0]), .out(h_s_cla32_and62));
  and_gate and_gate_h_s_cla32_and63(.a(h_s_cla32_pg_logic15_or0[0]), .b(h_s_cla32_pg_logic13_or0[0]), .out(h_s_cla32_and63));
  and_gate and_gate_h_s_cla32_and64(.a(h_s_cla32_and62[0]), .b(h_s_cla32_and63[0]), .out(h_s_cla32_and64));
  and_gate and_gate_h_s_cla32_and65(.a(h_s_cla32_and64[0]), .b(h_s_cla32_pg_logic12_or0[0]), .out(h_s_cla32_and65));
  and_gate and_gate_h_s_cla32_and66(.a(h_s_cla32_pg_logic12_and0[0]), .b(h_s_cla32_pg_logic14_or0[0]), .out(h_s_cla32_and66));
  and_gate and_gate_h_s_cla32_and67(.a(h_s_cla32_pg_logic15_or0[0]), .b(h_s_cla32_pg_logic13_or0[0]), .out(h_s_cla32_and67));
  and_gate and_gate_h_s_cla32_and68(.a(h_s_cla32_and66[0]), .b(h_s_cla32_and67[0]), .out(h_s_cla32_and68));
  and_gate and_gate_h_s_cla32_and69(.a(h_s_cla32_pg_logic13_and0[0]), .b(h_s_cla32_pg_logic15_or0[0]), .out(h_s_cla32_and69));
  and_gate and_gate_h_s_cla32_and70(.a(h_s_cla32_and69[0]), .b(h_s_cla32_pg_logic14_or0[0]), .out(h_s_cla32_and70));
  and_gate and_gate_h_s_cla32_and71(.a(h_s_cla32_pg_logic14_and0[0]), .b(h_s_cla32_pg_logic15_or0[0]), .out(h_s_cla32_and71));
  or_gate or_gate_h_s_cla32_or32(.a(h_s_cla32_and65[0]), .b(h_s_cla32_and70[0]), .out(h_s_cla32_or32));
  or_gate or_gate_h_s_cla32_or33(.a(h_s_cla32_and68[0]), .b(h_s_cla32_and71[0]), .out(h_s_cla32_or33));
  or_gate or_gate_h_s_cla32_or34(.a(h_s_cla32_or32[0]), .b(h_s_cla32_or33[0]), .out(h_s_cla32_or34));
  or_gate or_gate_h_s_cla32_or35(.a(h_s_cla32_pg_logic15_and0[0]), .b(h_s_cla32_or34[0]), .out(h_s_cla32_or35));
  pg_logic pg_logic_h_s_cla32_pg_logic16_out(.a(a[16]), .b(b[16]), .pg_logic_or0(h_s_cla32_pg_logic16_or0), .pg_logic_and0(h_s_cla32_pg_logic16_and0), .pg_logic_xor0(h_s_cla32_pg_logic16_xor0));
  xor_gate xor_gate_h_s_cla32_xor16(.a(h_s_cla32_pg_logic16_xor0[0]), .b(h_s_cla32_or35[0]), .out(h_s_cla32_xor16));
  and_gate and_gate_h_s_cla32_and72(.a(h_s_cla32_or35[0]), .b(h_s_cla32_pg_logic16_or0[0]), .out(h_s_cla32_and72));
  or_gate or_gate_h_s_cla32_or36(.a(h_s_cla32_pg_logic16_and0[0]), .b(h_s_cla32_and72[0]), .out(h_s_cla32_or36));
  pg_logic pg_logic_h_s_cla32_pg_logic17_out(.a(a[17]), .b(b[17]), .pg_logic_or0(h_s_cla32_pg_logic17_or0), .pg_logic_and0(h_s_cla32_pg_logic17_and0), .pg_logic_xor0(h_s_cla32_pg_logic17_xor0));
  xor_gate xor_gate_h_s_cla32_xor17(.a(h_s_cla32_pg_logic17_xor0[0]), .b(h_s_cla32_or36[0]), .out(h_s_cla32_xor17));
  and_gate and_gate_h_s_cla32_and73(.a(h_s_cla32_or35[0]), .b(h_s_cla32_pg_logic17_or0[0]), .out(h_s_cla32_and73));
  and_gate and_gate_h_s_cla32_and74(.a(h_s_cla32_and73[0]), .b(h_s_cla32_pg_logic16_or0[0]), .out(h_s_cla32_and74));
  and_gate and_gate_h_s_cla32_and75(.a(h_s_cla32_pg_logic16_and0[0]), .b(h_s_cla32_pg_logic17_or0[0]), .out(h_s_cla32_and75));
  or_gate or_gate_h_s_cla32_or37(.a(h_s_cla32_and74[0]), .b(h_s_cla32_and75[0]), .out(h_s_cla32_or37));
  or_gate or_gate_h_s_cla32_or38(.a(h_s_cla32_pg_logic17_and0[0]), .b(h_s_cla32_or37[0]), .out(h_s_cla32_or38));
  pg_logic pg_logic_h_s_cla32_pg_logic18_out(.a(a[18]), .b(b[18]), .pg_logic_or0(h_s_cla32_pg_logic18_or0), .pg_logic_and0(h_s_cla32_pg_logic18_and0), .pg_logic_xor0(h_s_cla32_pg_logic18_xor0));
  xor_gate xor_gate_h_s_cla32_xor18(.a(h_s_cla32_pg_logic18_xor0[0]), .b(h_s_cla32_or38[0]), .out(h_s_cla32_xor18));
  and_gate and_gate_h_s_cla32_and76(.a(h_s_cla32_or35[0]), .b(h_s_cla32_pg_logic17_or0[0]), .out(h_s_cla32_and76));
  and_gate and_gate_h_s_cla32_and77(.a(h_s_cla32_pg_logic18_or0[0]), .b(h_s_cla32_pg_logic16_or0[0]), .out(h_s_cla32_and77));
  and_gate and_gate_h_s_cla32_and78(.a(h_s_cla32_and76[0]), .b(h_s_cla32_and77[0]), .out(h_s_cla32_and78));
  and_gate and_gate_h_s_cla32_and79(.a(h_s_cla32_pg_logic16_and0[0]), .b(h_s_cla32_pg_logic18_or0[0]), .out(h_s_cla32_and79));
  and_gate and_gate_h_s_cla32_and80(.a(h_s_cla32_and79[0]), .b(h_s_cla32_pg_logic17_or0[0]), .out(h_s_cla32_and80));
  and_gate and_gate_h_s_cla32_and81(.a(h_s_cla32_pg_logic17_and0[0]), .b(h_s_cla32_pg_logic18_or0[0]), .out(h_s_cla32_and81));
  or_gate or_gate_h_s_cla32_or39(.a(h_s_cla32_and78[0]), .b(h_s_cla32_and80[0]), .out(h_s_cla32_or39));
  or_gate or_gate_h_s_cla32_or40(.a(h_s_cla32_or39[0]), .b(h_s_cla32_and81[0]), .out(h_s_cla32_or40));
  or_gate or_gate_h_s_cla32_or41(.a(h_s_cla32_pg_logic18_and0[0]), .b(h_s_cla32_or40[0]), .out(h_s_cla32_or41));
  pg_logic pg_logic_h_s_cla32_pg_logic19_out(.a(a[19]), .b(b[19]), .pg_logic_or0(h_s_cla32_pg_logic19_or0), .pg_logic_and0(h_s_cla32_pg_logic19_and0), .pg_logic_xor0(h_s_cla32_pg_logic19_xor0));
  xor_gate xor_gate_h_s_cla32_xor19(.a(h_s_cla32_pg_logic19_xor0[0]), .b(h_s_cla32_or41[0]), .out(h_s_cla32_xor19));
  and_gate and_gate_h_s_cla32_and82(.a(h_s_cla32_or35[0]), .b(h_s_cla32_pg_logic18_or0[0]), .out(h_s_cla32_and82));
  and_gate and_gate_h_s_cla32_and83(.a(h_s_cla32_pg_logic19_or0[0]), .b(h_s_cla32_pg_logic17_or0[0]), .out(h_s_cla32_and83));
  and_gate and_gate_h_s_cla32_and84(.a(h_s_cla32_and82[0]), .b(h_s_cla32_and83[0]), .out(h_s_cla32_and84));
  and_gate and_gate_h_s_cla32_and85(.a(h_s_cla32_and84[0]), .b(h_s_cla32_pg_logic16_or0[0]), .out(h_s_cla32_and85));
  and_gate and_gate_h_s_cla32_and86(.a(h_s_cla32_pg_logic16_and0[0]), .b(h_s_cla32_pg_logic18_or0[0]), .out(h_s_cla32_and86));
  and_gate and_gate_h_s_cla32_and87(.a(h_s_cla32_pg_logic19_or0[0]), .b(h_s_cla32_pg_logic17_or0[0]), .out(h_s_cla32_and87));
  and_gate and_gate_h_s_cla32_and88(.a(h_s_cla32_and86[0]), .b(h_s_cla32_and87[0]), .out(h_s_cla32_and88));
  and_gate and_gate_h_s_cla32_and89(.a(h_s_cla32_pg_logic17_and0[0]), .b(h_s_cla32_pg_logic19_or0[0]), .out(h_s_cla32_and89));
  and_gate and_gate_h_s_cla32_and90(.a(h_s_cla32_and89[0]), .b(h_s_cla32_pg_logic18_or0[0]), .out(h_s_cla32_and90));
  and_gate and_gate_h_s_cla32_and91(.a(h_s_cla32_pg_logic18_and0[0]), .b(h_s_cla32_pg_logic19_or0[0]), .out(h_s_cla32_and91));
  or_gate or_gate_h_s_cla32_or42(.a(h_s_cla32_and85[0]), .b(h_s_cla32_and90[0]), .out(h_s_cla32_or42));
  or_gate or_gate_h_s_cla32_or43(.a(h_s_cla32_and88[0]), .b(h_s_cla32_and91[0]), .out(h_s_cla32_or43));
  or_gate or_gate_h_s_cla32_or44(.a(h_s_cla32_or42[0]), .b(h_s_cla32_or43[0]), .out(h_s_cla32_or44));
  or_gate or_gate_h_s_cla32_or45(.a(h_s_cla32_pg_logic19_and0[0]), .b(h_s_cla32_or44[0]), .out(h_s_cla32_or45));
  pg_logic pg_logic_h_s_cla32_pg_logic20_out(.a(a[20]), .b(b[20]), .pg_logic_or0(h_s_cla32_pg_logic20_or0), .pg_logic_and0(h_s_cla32_pg_logic20_and0), .pg_logic_xor0(h_s_cla32_pg_logic20_xor0));
  xor_gate xor_gate_h_s_cla32_xor20(.a(h_s_cla32_pg_logic20_xor0[0]), .b(h_s_cla32_or45[0]), .out(h_s_cla32_xor20));
  and_gate and_gate_h_s_cla32_and92(.a(h_s_cla32_or45[0]), .b(h_s_cla32_pg_logic20_or0[0]), .out(h_s_cla32_and92));
  or_gate or_gate_h_s_cla32_or46(.a(h_s_cla32_pg_logic20_and0[0]), .b(h_s_cla32_and92[0]), .out(h_s_cla32_or46));
  pg_logic pg_logic_h_s_cla32_pg_logic21_out(.a(a[21]), .b(b[21]), .pg_logic_or0(h_s_cla32_pg_logic21_or0), .pg_logic_and0(h_s_cla32_pg_logic21_and0), .pg_logic_xor0(h_s_cla32_pg_logic21_xor0));
  xor_gate xor_gate_h_s_cla32_xor21(.a(h_s_cla32_pg_logic21_xor0[0]), .b(h_s_cla32_or46[0]), .out(h_s_cla32_xor21));
  and_gate and_gate_h_s_cla32_and93(.a(h_s_cla32_or45[0]), .b(h_s_cla32_pg_logic21_or0[0]), .out(h_s_cla32_and93));
  and_gate and_gate_h_s_cla32_and94(.a(h_s_cla32_and93[0]), .b(h_s_cla32_pg_logic20_or0[0]), .out(h_s_cla32_and94));
  and_gate and_gate_h_s_cla32_and95(.a(h_s_cla32_pg_logic20_and0[0]), .b(h_s_cla32_pg_logic21_or0[0]), .out(h_s_cla32_and95));
  or_gate or_gate_h_s_cla32_or47(.a(h_s_cla32_and94[0]), .b(h_s_cla32_and95[0]), .out(h_s_cla32_or47));
  or_gate or_gate_h_s_cla32_or48(.a(h_s_cla32_pg_logic21_and0[0]), .b(h_s_cla32_or47[0]), .out(h_s_cla32_or48));
  pg_logic pg_logic_h_s_cla32_pg_logic22_out(.a(a[22]), .b(b[22]), .pg_logic_or0(h_s_cla32_pg_logic22_or0), .pg_logic_and0(h_s_cla32_pg_logic22_and0), .pg_logic_xor0(h_s_cla32_pg_logic22_xor0));
  xor_gate xor_gate_h_s_cla32_xor22(.a(h_s_cla32_pg_logic22_xor0[0]), .b(h_s_cla32_or48[0]), .out(h_s_cla32_xor22));
  and_gate and_gate_h_s_cla32_and96(.a(h_s_cla32_or45[0]), .b(h_s_cla32_pg_logic21_or0[0]), .out(h_s_cla32_and96));
  and_gate and_gate_h_s_cla32_and97(.a(h_s_cla32_pg_logic22_or0[0]), .b(h_s_cla32_pg_logic20_or0[0]), .out(h_s_cla32_and97));
  and_gate and_gate_h_s_cla32_and98(.a(h_s_cla32_and96[0]), .b(h_s_cla32_and97[0]), .out(h_s_cla32_and98));
  and_gate and_gate_h_s_cla32_and99(.a(h_s_cla32_pg_logic20_and0[0]), .b(h_s_cla32_pg_logic22_or0[0]), .out(h_s_cla32_and99));
  and_gate and_gate_h_s_cla32_and100(.a(h_s_cla32_and99[0]), .b(h_s_cla32_pg_logic21_or0[0]), .out(h_s_cla32_and100));
  and_gate and_gate_h_s_cla32_and101(.a(h_s_cla32_pg_logic21_and0[0]), .b(h_s_cla32_pg_logic22_or0[0]), .out(h_s_cla32_and101));
  or_gate or_gate_h_s_cla32_or49(.a(h_s_cla32_and98[0]), .b(h_s_cla32_and100[0]), .out(h_s_cla32_or49));
  or_gate or_gate_h_s_cla32_or50(.a(h_s_cla32_or49[0]), .b(h_s_cla32_and101[0]), .out(h_s_cla32_or50));
  or_gate or_gate_h_s_cla32_or51(.a(h_s_cla32_pg_logic22_and0[0]), .b(h_s_cla32_or50[0]), .out(h_s_cla32_or51));
  pg_logic pg_logic_h_s_cla32_pg_logic23_out(.a(a[23]), .b(b[23]), .pg_logic_or0(h_s_cla32_pg_logic23_or0), .pg_logic_and0(h_s_cla32_pg_logic23_and0), .pg_logic_xor0(h_s_cla32_pg_logic23_xor0));
  xor_gate xor_gate_h_s_cla32_xor23(.a(h_s_cla32_pg_logic23_xor0[0]), .b(h_s_cla32_or51[0]), .out(h_s_cla32_xor23));
  and_gate and_gate_h_s_cla32_and102(.a(h_s_cla32_or45[0]), .b(h_s_cla32_pg_logic22_or0[0]), .out(h_s_cla32_and102));
  and_gate and_gate_h_s_cla32_and103(.a(h_s_cla32_pg_logic23_or0[0]), .b(h_s_cla32_pg_logic21_or0[0]), .out(h_s_cla32_and103));
  and_gate and_gate_h_s_cla32_and104(.a(h_s_cla32_and102[0]), .b(h_s_cla32_and103[0]), .out(h_s_cla32_and104));
  and_gate and_gate_h_s_cla32_and105(.a(h_s_cla32_and104[0]), .b(h_s_cla32_pg_logic20_or0[0]), .out(h_s_cla32_and105));
  and_gate and_gate_h_s_cla32_and106(.a(h_s_cla32_pg_logic20_and0[0]), .b(h_s_cla32_pg_logic22_or0[0]), .out(h_s_cla32_and106));
  and_gate and_gate_h_s_cla32_and107(.a(h_s_cla32_pg_logic23_or0[0]), .b(h_s_cla32_pg_logic21_or0[0]), .out(h_s_cla32_and107));
  and_gate and_gate_h_s_cla32_and108(.a(h_s_cla32_and106[0]), .b(h_s_cla32_and107[0]), .out(h_s_cla32_and108));
  and_gate and_gate_h_s_cla32_and109(.a(h_s_cla32_pg_logic21_and0[0]), .b(h_s_cla32_pg_logic23_or0[0]), .out(h_s_cla32_and109));
  and_gate and_gate_h_s_cla32_and110(.a(h_s_cla32_and109[0]), .b(h_s_cla32_pg_logic22_or0[0]), .out(h_s_cla32_and110));
  and_gate and_gate_h_s_cla32_and111(.a(h_s_cla32_pg_logic22_and0[0]), .b(h_s_cla32_pg_logic23_or0[0]), .out(h_s_cla32_and111));
  or_gate or_gate_h_s_cla32_or52(.a(h_s_cla32_and105[0]), .b(h_s_cla32_and110[0]), .out(h_s_cla32_or52));
  or_gate or_gate_h_s_cla32_or53(.a(h_s_cla32_and108[0]), .b(h_s_cla32_and111[0]), .out(h_s_cla32_or53));
  or_gate or_gate_h_s_cla32_or54(.a(h_s_cla32_or52[0]), .b(h_s_cla32_or53[0]), .out(h_s_cla32_or54));
  or_gate or_gate_h_s_cla32_or55(.a(h_s_cla32_pg_logic23_and0[0]), .b(h_s_cla32_or54[0]), .out(h_s_cla32_or55));
  pg_logic pg_logic_h_s_cla32_pg_logic24_out(.a(a[24]), .b(b[24]), .pg_logic_or0(h_s_cla32_pg_logic24_or0), .pg_logic_and0(h_s_cla32_pg_logic24_and0), .pg_logic_xor0(h_s_cla32_pg_logic24_xor0));
  xor_gate xor_gate_h_s_cla32_xor24(.a(h_s_cla32_pg_logic24_xor0[0]), .b(h_s_cla32_or55[0]), .out(h_s_cla32_xor24));
  and_gate and_gate_h_s_cla32_and112(.a(h_s_cla32_or55[0]), .b(h_s_cla32_pg_logic24_or0[0]), .out(h_s_cla32_and112));
  or_gate or_gate_h_s_cla32_or56(.a(h_s_cla32_pg_logic24_and0[0]), .b(h_s_cla32_and112[0]), .out(h_s_cla32_or56));
  pg_logic pg_logic_h_s_cla32_pg_logic25_out(.a(a[25]), .b(b[25]), .pg_logic_or0(h_s_cla32_pg_logic25_or0), .pg_logic_and0(h_s_cla32_pg_logic25_and0), .pg_logic_xor0(h_s_cla32_pg_logic25_xor0));
  xor_gate xor_gate_h_s_cla32_xor25(.a(h_s_cla32_pg_logic25_xor0[0]), .b(h_s_cla32_or56[0]), .out(h_s_cla32_xor25));
  and_gate and_gate_h_s_cla32_and113(.a(h_s_cla32_or55[0]), .b(h_s_cla32_pg_logic25_or0[0]), .out(h_s_cla32_and113));
  and_gate and_gate_h_s_cla32_and114(.a(h_s_cla32_and113[0]), .b(h_s_cla32_pg_logic24_or0[0]), .out(h_s_cla32_and114));
  and_gate and_gate_h_s_cla32_and115(.a(h_s_cla32_pg_logic24_and0[0]), .b(h_s_cla32_pg_logic25_or0[0]), .out(h_s_cla32_and115));
  or_gate or_gate_h_s_cla32_or57(.a(h_s_cla32_and114[0]), .b(h_s_cla32_and115[0]), .out(h_s_cla32_or57));
  or_gate or_gate_h_s_cla32_or58(.a(h_s_cla32_pg_logic25_and0[0]), .b(h_s_cla32_or57[0]), .out(h_s_cla32_or58));
  pg_logic pg_logic_h_s_cla32_pg_logic26_out(.a(a[26]), .b(b[26]), .pg_logic_or0(h_s_cla32_pg_logic26_or0), .pg_logic_and0(h_s_cla32_pg_logic26_and0), .pg_logic_xor0(h_s_cla32_pg_logic26_xor0));
  xor_gate xor_gate_h_s_cla32_xor26(.a(h_s_cla32_pg_logic26_xor0[0]), .b(h_s_cla32_or58[0]), .out(h_s_cla32_xor26));
  and_gate and_gate_h_s_cla32_and116(.a(h_s_cla32_or55[0]), .b(h_s_cla32_pg_logic25_or0[0]), .out(h_s_cla32_and116));
  and_gate and_gate_h_s_cla32_and117(.a(h_s_cla32_pg_logic26_or0[0]), .b(h_s_cla32_pg_logic24_or0[0]), .out(h_s_cla32_and117));
  and_gate and_gate_h_s_cla32_and118(.a(h_s_cla32_and116[0]), .b(h_s_cla32_and117[0]), .out(h_s_cla32_and118));
  and_gate and_gate_h_s_cla32_and119(.a(h_s_cla32_pg_logic24_and0[0]), .b(h_s_cla32_pg_logic26_or0[0]), .out(h_s_cla32_and119));
  and_gate and_gate_h_s_cla32_and120(.a(h_s_cla32_and119[0]), .b(h_s_cla32_pg_logic25_or0[0]), .out(h_s_cla32_and120));
  and_gate and_gate_h_s_cla32_and121(.a(h_s_cla32_pg_logic25_and0[0]), .b(h_s_cla32_pg_logic26_or0[0]), .out(h_s_cla32_and121));
  or_gate or_gate_h_s_cla32_or59(.a(h_s_cla32_and118[0]), .b(h_s_cla32_and120[0]), .out(h_s_cla32_or59));
  or_gate or_gate_h_s_cla32_or60(.a(h_s_cla32_or59[0]), .b(h_s_cla32_and121[0]), .out(h_s_cla32_or60));
  or_gate or_gate_h_s_cla32_or61(.a(h_s_cla32_pg_logic26_and0[0]), .b(h_s_cla32_or60[0]), .out(h_s_cla32_or61));
  pg_logic pg_logic_h_s_cla32_pg_logic27_out(.a(a[27]), .b(b[27]), .pg_logic_or0(h_s_cla32_pg_logic27_or0), .pg_logic_and0(h_s_cla32_pg_logic27_and0), .pg_logic_xor0(h_s_cla32_pg_logic27_xor0));
  xor_gate xor_gate_h_s_cla32_xor27(.a(h_s_cla32_pg_logic27_xor0[0]), .b(h_s_cla32_or61[0]), .out(h_s_cla32_xor27));
  and_gate and_gate_h_s_cla32_and122(.a(h_s_cla32_or55[0]), .b(h_s_cla32_pg_logic26_or0[0]), .out(h_s_cla32_and122));
  and_gate and_gate_h_s_cla32_and123(.a(h_s_cla32_pg_logic27_or0[0]), .b(h_s_cla32_pg_logic25_or0[0]), .out(h_s_cla32_and123));
  and_gate and_gate_h_s_cla32_and124(.a(h_s_cla32_and122[0]), .b(h_s_cla32_and123[0]), .out(h_s_cla32_and124));
  and_gate and_gate_h_s_cla32_and125(.a(h_s_cla32_and124[0]), .b(h_s_cla32_pg_logic24_or0[0]), .out(h_s_cla32_and125));
  and_gate and_gate_h_s_cla32_and126(.a(h_s_cla32_pg_logic24_and0[0]), .b(h_s_cla32_pg_logic26_or0[0]), .out(h_s_cla32_and126));
  and_gate and_gate_h_s_cla32_and127(.a(h_s_cla32_pg_logic27_or0[0]), .b(h_s_cla32_pg_logic25_or0[0]), .out(h_s_cla32_and127));
  and_gate and_gate_h_s_cla32_and128(.a(h_s_cla32_and126[0]), .b(h_s_cla32_and127[0]), .out(h_s_cla32_and128));
  and_gate and_gate_h_s_cla32_and129(.a(h_s_cla32_pg_logic25_and0[0]), .b(h_s_cla32_pg_logic27_or0[0]), .out(h_s_cla32_and129));
  and_gate and_gate_h_s_cla32_and130(.a(h_s_cla32_and129[0]), .b(h_s_cla32_pg_logic26_or0[0]), .out(h_s_cla32_and130));
  and_gate and_gate_h_s_cla32_and131(.a(h_s_cla32_pg_logic26_and0[0]), .b(h_s_cla32_pg_logic27_or0[0]), .out(h_s_cla32_and131));
  or_gate or_gate_h_s_cla32_or62(.a(h_s_cla32_and125[0]), .b(h_s_cla32_and130[0]), .out(h_s_cla32_or62));
  or_gate or_gate_h_s_cla32_or63(.a(h_s_cla32_and128[0]), .b(h_s_cla32_and131[0]), .out(h_s_cla32_or63));
  or_gate or_gate_h_s_cla32_or64(.a(h_s_cla32_or62[0]), .b(h_s_cla32_or63[0]), .out(h_s_cla32_or64));
  or_gate or_gate_h_s_cla32_or65(.a(h_s_cla32_pg_logic27_and0[0]), .b(h_s_cla32_or64[0]), .out(h_s_cla32_or65));
  pg_logic pg_logic_h_s_cla32_pg_logic28_out(.a(a[28]), .b(b[28]), .pg_logic_or0(h_s_cla32_pg_logic28_or0), .pg_logic_and0(h_s_cla32_pg_logic28_and0), .pg_logic_xor0(h_s_cla32_pg_logic28_xor0));
  xor_gate xor_gate_h_s_cla32_xor28(.a(h_s_cla32_pg_logic28_xor0[0]), .b(h_s_cla32_or65[0]), .out(h_s_cla32_xor28));
  and_gate and_gate_h_s_cla32_and132(.a(h_s_cla32_or65[0]), .b(h_s_cla32_pg_logic28_or0[0]), .out(h_s_cla32_and132));
  or_gate or_gate_h_s_cla32_or66(.a(h_s_cla32_pg_logic28_and0[0]), .b(h_s_cla32_and132[0]), .out(h_s_cla32_or66));
  pg_logic pg_logic_h_s_cla32_pg_logic29_out(.a(a[29]), .b(b[29]), .pg_logic_or0(h_s_cla32_pg_logic29_or0), .pg_logic_and0(h_s_cla32_pg_logic29_and0), .pg_logic_xor0(h_s_cla32_pg_logic29_xor0));
  xor_gate xor_gate_h_s_cla32_xor29(.a(h_s_cla32_pg_logic29_xor0[0]), .b(h_s_cla32_or66[0]), .out(h_s_cla32_xor29));
  and_gate and_gate_h_s_cla32_and133(.a(h_s_cla32_or65[0]), .b(h_s_cla32_pg_logic29_or0[0]), .out(h_s_cla32_and133));
  and_gate and_gate_h_s_cla32_and134(.a(h_s_cla32_and133[0]), .b(h_s_cla32_pg_logic28_or0[0]), .out(h_s_cla32_and134));
  and_gate and_gate_h_s_cla32_and135(.a(h_s_cla32_pg_logic28_and0[0]), .b(h_s_cla32_pg_logic29_or0[0]), .out(h_s_cla32_and135));
  or_gate or_gate_h_s_cla32_or67(.a(h_s_cla32_and134[0]), .b(h_s_cla32_and135[0]), .out(h_s_cla32_or67));
  or_gate or_gate_h_s_cla32_or68(.a(h_s_cla32_pg_logic29_and0[0]), .b(h_s_cla32_or67[0]), .out(h_s_cla32_or68));
  pg_logic pg_logic_h_s_cla32_pg_logic30_out(.a(a[30]), .b(b[30]), .pg_logic_or0(h_s_cla32_pg_logic30_or0), .pg_logic_and0(h_s_cla32_pg_logic30_and0), .pg_logic_xor0(h_s_cla32_pg_logic30_xor0));
  xor_gate xor_gate_h_s_cla32_xor30(.a(h_s_cla32_pg_logic30_xor0[0]), .b(h_s_cla32_or68[0]), .out(h_s_cla32_xor30));
  and_gate and_gate_h_s_cla32_and136(.a(h_s_cla32_or65[0]), .b(h_s_cla32_pg_logic29_or0[0]), .out(h_s_cla32_and136));
  and_gate and_gate_h_s_cla32_and137(.a(h_s_cla32_pg_logic30_or0[0]), .b(h_s_cla32_pg_logic28_or0[0]), .out(h_s_cla32_and137));
  and_gate and_gate_h_s_cla32_and138(.a(h_s_cla32_and136[0]), .b(h_s_cla32_and137[0]), .out(h_s_cla32_and138));
  and_gate and_gate_h_s_cla32_and139(.a(h_s_cla32_pg_logic28_and0[0]), .b(h_s_cla32_pg_logic30_or0[0]), .out(h_s_cla32_and139));
  and_gate and_gate_h_s_cla32_and140(.a(h_s_cla32_and139[0]), .b(h_s_cla32_pg_logic29_or0[0]), .out(h_s_cla32_and140));
  and_gate and_gate_h_s_cla32_and141(.a(h_s_cla32_pg_logic29_and0[0]), .b(h_s_cla32_pg_logic30_or0[0]), .out(h_s_cla32_and141));
  or_gate or_gate_h_s_cla32_or69(.a(h_s_cla32_and138[0]), .b(h_s_cla32_and140[0]), .out(h_s_cla32_or69));
  or_gate or_gate_h_s_cla32_or70(.a(h_s_cla32_or69[0]), .b(h_s_cla32_and141[0]), .out(h_s_cla32_or70));
  or_gate or_gate_h_s_cla32_or71(.a(h_s_cla32_pg_logic30_and0[0]), .b(h_s_cla32_or70[0]), .out(h_s_cla32_or71));
  pg_logic pg_logic_h_s_cla32_pg_logic31_out(.a(a[31]), .b(b[31]), .pg_logic_or0(h_s_cla32_pg_logic31_or0), .pg_logic_and0(h_s_cla32_pg_logic31_and0), .pg_logic_xor0(h_s_cla32_pg_logic31_xor0));
  xor_gate xor_gate_h_s_cla32_xor31(.a(h_s_cla32_pg_logic31_xor0[0]), .b(h_s_cla32_or71[0]), .out(h_s_cla32_xor31));
  and_gate and_gate_h_s_cla32_and142(.a(h_s_cla32_or65[0]), .b(h_s_cla32_pg_logic30_or0[0]), .out(h_s_cla32_and142));
  and_gate and_gate_h_s_cla32_and143(.a(h_s_cla32_pg_logic31_or0[0]), .b(h_s_cla32_pg_logic29_or0[0]), .out(h_s_cla32_and143));
  and_gate and_gate_h_s_cla32_and144(.a(h_s_cla32_and142[0]), .b(h_s_cla32_and143[0]), .out(h_s_cla32_and144));
  and_gate and_gate_h_s_cla32_and145(.a(h_s_cla32_and144[0]), .b(h_s_cla32_pg_logic28_or0[0]), .out(h_s_cla32_and145));
  and_gate and_gate_h_s_cla32_and146(.a(h_s_cla32_pg_logic28_and0[0]), .b(h_s_cla32_pg_logic30_or0[0]), .out(h_s_cla32_and146));
  and_gate and_gate_h_s_cla32_and147(.a(h_s_cla32_pg_logic31_or0[0]), .b(h_s_cla32_pg_logic29_or0[0]), .out(h_s_cla32_and147));
  and_gate and_gate_h_s_cla32_and148(.a(h_s_cla32_and146[0]), .b(h_s_cla32_and147[0]), .out(h_s_cla32_and148));
  and_gate and_gate_h_s_cla32_and149(.a(h_s_cla32_pg_logic29_and0[0]), .b(h_s_cla32_pg_logic31_or0[0]), .out(h_s_cla32_and149));
  and_gate and_gate_h_s_cla32_and150(.a(h_s_cla32_and149[0]), .b(h_s_cla32_pg_logic30_or0[0]), .out(h_s_cla32_and150));
  and_gate and_gate_h_s_cla32_and151(.a(h_s_cla32_pg_logic30_and0[0]), .b(h_s_cla32_pg_logic31_or0[0]), .out(h_s_cla32_and151));
  or_gate or_gate_h_s_cla32_or72(.a(h_s_cla32_and145[0]), .b(h_s_cla32_and150[0]), .out(h_s_cla32_or72));
  or_gate or_gate_h_s_cla32_or73(.a(h_s_cla32_and148[0]), .b(h_s_cla32_and151[0]), .out(h_s_cla32_or73));
  or_gate or_gate_h_s_cla32_or74(.a(h_s_cla32_or72[0]), .b(h_s_cla32_or73[0]), .out(h_s_cla32_or74));
  or_gate or_gate_h_s_cla32_or75(.a(h_s_cla32_pg_logic31_and0[0]), .b(h_s_cla32_or74[0]), .out(h_s_cla32_or75));
  xor_gate xor_gate_h_s_cla32_xor32(.a(a[31]), .b(b[31]), .out(h_s_cla32_xor32));
  xor_gate xor_gate_h_s_cla32_xor33(.a(h_s_cla32_xor32[0]), .b(h_s_cla32_or75[0]), .out(h_s_cla32_xor33));

  assign h_s_cla32_out[0] = h_s_cla32_pg_logic0_xor0[0];
  assign h_s_cla32_out[1] = h_s_cla32_xor1[0];
  assign h_s_cla32_out[2] = h_s_cla32_xor2[0];
  assign h_s_cla32_out[3] = h_s_cla32_xor3[0];
  assign h_s_cla32_out[4] = h_s_cla32_xor4[0];
  assign h_s_cla32_out[5] = h_s_cla32_xor5[0];
  assign h_s_cla32_out[6] = h_s_cla32_xor6[0];
  assign h_s_cla32_out[7] = h_s_cla32_xor7[0];
  assign h_s_cla32_out[8] = h_s_cla32_xor8[0];
  assign h_s_cla32_out[9] = h_s_cla32_xor9[0];
  assign h_s_cla32_out[10] = h_s_cla32_xor10[0];
  assign h_s_cla32_out[11] = h_s_cla32_xor11[0];
  assign h_s_cla32_out[12] = h_s_cla32_xor12[0];
  assign h_s_cla32_out[13] = h_s_cla32_xor13[0];
  assign h_s_cla32_out[14] = h_s_cla32_xor14[0];
  assign h_s_cla32_out[15] = h_s_cla32_xor15[0];
  assign h_s_cla32_out[16] = h_s_cla32_xor16[0];
  assign h_s_cla32_out[17] = h_s_cla32_xor17[0];
  assign h_s_cla32_out[18] = h_s_cla32_xor18[0];
  assign h_s_cla32_out[19] = h_s_cla32_xor19[0];
  assign h_s_cla32_out[20] = h_s_cla32_xor20[0];
  assign h_s_cla32_out[21] = h_s_cla32_xor21[0];
  assign h_s_cla32_out[22] = h_s_cla32_xor22[0];
  assign h_s_cla32_out[23] = h_s_cla32_xor23[0];
  assign h_s_cla32_out[24] = h_s_cla32_xor24[0];
  assign h_s_cla32_out[25] = h_s_cla32_xor25[0];
  assign h_s_cla32_out[26] = h_s_cla32_xor26[0];
  assign h_s_cla32_out[27] = h_s_cla32_xor27[0];
  assign h_s_cla32_out[28] = h_s_cla32_xor28[0];
  assign h_s_cla32_out[29] = h_s_cla32_xor29[0];
  assign h_s_cla32_out[30] = h_s_cla32_xor30[0];
  assign h_s_cla32_out[31] = h_s_cla32_xor31[0];
  assign h_s_cla32_out[32] = h_s_cla32_xor33[0];
endmodule