module s_csamul_cla32(input [31:0] a, input [31:0] b, output [63:0] s_csamul_cla32_out);
  wire s_csamul_cla32_and0_0;
  wire s_csamul_cla32_and1_0;
  wire s_csamul_cla32_and2_0;
  wire s_csamul_cla32_and3_0;
  wire s_csamul_cla32_and4_0;
  wire s_csamul_cla32_and5_0;
  wire s_csamul_cla32_and6_0;
  wire s_csamul_cla32_and7_0;
  wire s_csamul_cla32_and8_0;
  wire s_csamul_cla32_and9_0;
  wire s_csamul_cla32_and10_0;
  wire s_csamul_cla32_and11_0;
  wire s_csamul_cla32_and12_0;
  wire s_csamul_cla32_and13_0;
  wire s_csamul_cla32_and14_0;
  wire s_csamul_cla32_and15_0;
  wire s_csamul_cla32_and16_0;
  wire s_csamul_cla32_and17_0;
  wire s_csamul_cla32_and18_0;
  wire s_csamul_cla32_and19_0;
  wire s_csamul_cla32_and20_0;
  wire s_csamul_cla32_and21_0;
  wire s_csamul_cla32_and22_0;
  wire s_csamul_cla32_and23_0;
  wire s_csamul_cla32_and24_0;
  wire s_csamul_cla32_and25_0;
  wire s_csamul_cla32_and26_0;
  wire s_csamul_cla32_and27_0;
  wire s_csamul_cla32_and28_0;
  wire s_csamul_cla32_and29_0;
  wire s_csamul_cla32_and30_0;
  wire s_csamul_cla32_nand31_0;
  wire s_csamul_cla32_and0_1;
  wire s_csamul_cla32_ha0_1_xor0;
  wire s_csamul_cla32_ha0_1_and0;
  wire s_csamul_cla32_and1_1;
  wire s_csamul_cla32_ha1_1_xor0;
  wire s_csamul_cla32_ha1_1_and0;
  wire s_csamul_cla32_and2_1;
  wire s_csamul_cla32_ha2_1_xor0;
  wire s_csamul_cla32_ha2_1_and0;
  wire s_csamul_cla32_and3_1;
  wire s_csamul_cla32_ha3_1_xor0;
  wire s_csamul_cla32_ha3_1_and0;
  wire s_csamul_cla32_and4_1;
  wire s_csamul_cla32_ha4_1_xor0;
  wire s_csamul_cla32_ha4_1_and0;
  wire s_csamul_cla32_and5_1;
  wire s_csamul_cla32_ha5_1_xor0;
  wire s_csamul_cla32_ha5_1_and0;
  wire s_csamul_cla32_and6_1;
  wire s_csamul_cla32_ha6_1_xor0;
  wire s_csamul_cla32_ha6_1_and0;
  wire s_csamul_cla32_and7_1;
  wire s_csamul_cla32_ha7_1_xor0;
  wire s_csamul_cla32_ha7_1_and0;
  wire s_csamul_cla32_and8_1;
  wire s_csamul_cla32_ha8_1_xor0;
  wire s_csamul_cla32_ha8_1_and0;
  wire s_csamul_cla32_and9_1;
  wire s_csamul_cla32_ha9_1_xor0;
  wire s_csamul_cla32_ha9_1_and0;
  wire s_csamul_cla32_and10_1;
  wire s_csamul_cla32_ha10_1_xor0;
  wire s_csamul_cla32_ha10_1_and0;
  wire s_csamul_cla32_and11_1;
  wire s_csamul_cla32_ha11_1_xor0;
  wire s_csamul_cla32_ha11_1_and0;
  wire s_csamul_cla32_and12_1;
  wire s_csamul_cla32_ha12_1_xor0;
  wire s_csamul_cla32_ha12_1_and0;
  wire s_csamul_cla32_and13_1;
  wire s_csamul_cla32_ha13_1_xor0;
  wire s_csamul_cla32_ha13_1_and0;
  wire s_csamul_cla32_and14_1;
  wire s_csamul_cla32_ha14_1_xor0;
  wire s_csamul_cla32_ha14_1_and0;
  wire s_csamul_cla32_and15_1;
  wire s_csamul_cla32_ha15_1_xor0;
  wire s_csamul_cla32_ha15_1_and0;
  wire s_csamul_cla32_and16_1;
  wire s_csamul_cla32_ha16_1_xor0;
  wire s_csamul_cla32_ha16_1_and0;
  wire s_csamul_cla32_and17_1;
  wire s_csamul_cla32_ha17_1_xor0;
  wire s_csamul_cla32_ha17_1_and0;
  wire s_csamul_cla32_and18_1;
  wire s_csamul_cla32_ha18_1_xor0;
  wire s_csamul_cla32_ha18_1_and0;
  wire s_csamul_cla32_and19_1;
  wire s_csamul_cla32_ha19_1_xor0;
  wire s_csamul_cla32_ha19_1_and0;
  wire s_csamul_cla32_and20_1;
  wire s_csamul_cla32_ha20_1_xor0;
  wire s_csamul_cla32_ha20_1_and0;
  wire s_csamul_cla32_and21_1;
  wire s_csamul_cla32_ha21_1_xor0;
  wire s_csamul_cla32_ha21_1_and0;
  wire s_csamul_cla32_and22_1;
  wire s_csamul_cla32_ha22_1_xor0;
  wire s_csamul_cla32_ha22_1_and0;
  wire s_csamul_cla32_and23_1;
  wire s_csamul_cla32_ha23_1_xor0;
  wire s_csamul_cla32_ha23_1_and0;
  wire s_csamul_cla32_and24_1;
  wire s_csamul_cla32_ha24_1_xor0;
  wire s_csamul_cla32_ha24_1_and0;
  wire s_csamul_cla32_and25_1;
  wire s_csamul_cla32_ha25_1_xor0;
  wire s_csamul_cla32_ha25_1_and0;
  wire s_csamul_cla32_and26_1;
  wire s_csamul_cla32_ha26_1_xor0;
  wire s_csamul_cla32_ha26_1_and0;
  wire s_csamul_cla32_and27_1;
  wire s_csamul_cla32_ha27_1_xor0;
  wire s_csamul_cla32_ha27_1_and0;
  wire s_csamul_cla32_and28_1;
  wire s_csamul_cla32_ha28_1_xor0;
  wire s_csamul_cla32_ha28_1_and0;
  wire s_csamul_cla32_and29_1;
  wire s_csamul_cla32_ha29_1_xor0;
  wire s_csamul_cla32_ha29_1_and0;
  wire s_csamul_cla32_and30_1;
  wire s_csamul_cla32_ha30_1_xor0;
  wire s_csamul_cla32_ha30_1_and0;
  wire s_csamul_cla32_nand31_1;
  wire s_csamul_cla32_ha31_1_xor0;
  wire s_csamul_cla32_and0_2;
  wire s_csamul_cla32_fa0_2_xor0;
  wire s_csamul_cla32_fa0_2_and0;
  wire s_csamul_cla32_fa0_2_xor1;
  wire s_csamul_cla32_fa0_2_and1;
  wire s_csamul_cla32_fa0_2_or0;
  wire s_csamul_cla32_and1_2;
  wire s_csamul_cla32_fa1_2_xor0;
  wire s_csamul_cla32_fa1_2_and0;
  wire s_csamul_cla32_fa1_2_xor1;
  wire s_csamul_cla32_fa1_2_and1;
  wire s_csamul_cla32_fa1_2_or0;
  wire s_csamul_cla32_and2_2;
  wire s_csamul_cla32_fa2_2_xor0;
  wire s_csamul_cla32_fa2_2_and0;
  wire s_csamul_cla32_fa2_2_xor1;
  wire s_csamul_cla32_fa2_2_and1;
  wire s_csamul_cla32_fa2_2_or0;
  wire s_csamul_cla32_and3_2;
  wire s_csamul_cla32_fa3_2_xor0;
  wire s_csamul_cla32_fa3_2_and0;
  wire s_csamul_cla32_fa3_2_xor1;
  wire s_csamul_cla32_fa3_2_and1;
  wire s_csamul_cla32_fa3_2_or0;
  wire s_csamul_cla32_and4_2;
  wire s_csamul_cla32_fa4_2_xor0;
  wire s_csamul_cla32_fa4_2_and0;
  wire s_csamul_cla32_fa4_2_xor1;
  wire s_csamul_cla32_fa4_2_and1;
  wire s_csamul_cla32_fa4_2_or0;
  wire s_csamul_cla32_and5_2;
  wire s_csamul_cla32_fa5_2_xor0;
  wire s_csamul_cla32_fa5_2_and0;
  wire s_csamul_cla32_fa5_2_xor1;
  wire s_csamul_cla32_fa5_2_and1;
  wire s_csamul_cla32_fa5_2_or0;
  wire s_csamul_cla32_and6_2;
  wire s_csamul_cla32_fa6_2_xor0;
  wire s_csamul_cla32_fa6_2_and0;
  wire s_csamul_cla32_fa6_2_xor1;
  wire s_csamul_cla32_fa6_2_and1;
  wire s_csamul_cla32_fa6_2_or0;
  wire s_csamul_cla32_and7_2;
  wire s_csamul_cla32_fa7_2_xor0;
  wire s_csamul_cla32_fa7_2_and0;
  wire s_csamul_cla32_fa7_2_xor1;
  wire s_csamul_cla32_fa7_2_and1;
  wire s_csamul_cla32_fa7_2_or0;
  wire s_csamul_cla32_and8_2;
  wire s_csamul_cla32_fa8_2_xor0;
  wire s_csamul_cla32_fa8_2_and0;
  wire s_csamul_cla32_fa8_2_xor1;
  wire s_csamul_cla32_fa8_2_and1;
  wire s_csamul_cla32_fa8_2_or0;
  wire s_csamul_cla32_and9_2;
  wire s_csamul_cla32_fa9_2_xor0;
  wire s_csamul_cla32_fa9_2_and0;
  wire s_csamul_cla32_fa9_2_xor1;
  wire s_csamul_cla32_fa9_2_and1;
  wire s_csamul_cla32_fa9_2_or0;
  wire s_csamul_cla32_and10_2;
  wire s_csamul_cla32_fa10_2_xor0;
  wire s_csamul_cla32_fa10_2_and0;
  wire s_csamul_cla32_fa10_2_xor1;
  wire s_csamul_cla32_fa10_2_and1;
  wire s_csamul_cla32_fa10_2_or0;
  wire s_csamul_cla32_and11_2;
  wire s_csamul_cla32_fa11_2_xor0;
  wire s_csamul_cla32_fa11_2_and0;
  wire s_csamul_cla32_fa11_2_xor1;
  wire s_csamul_cla32_fa11_2_and1;
  wire s_csamul_cla32_fa11_2_or0;
  wire s_csamul_cla32_and12_2;
  wire s_csamul_cla32_fa12_2_xor0;
  wire s_csamul_cla32_fa12_2_and0;
  wire s_csamul_cla32_fa12_2_xor1;
  wire s_csamul_cla32_fa12_2_and1;
  wire s_csamul_cla32_fa12_2_or0;
  wire s_csamul_cla32_and13_2;
  wire s_csamul_cla32_fa13_2_xor0;
  wire s_csamul_cla32_fa13_2_and0;
  wire s_csamul_cla32_fa13_2_xor1;
  wire s_csamul_cla32_fa13_2_and1;
  wire s_csamul_cla32_fa13_2_or0;
  wire s_csamul_cla32_and14_2;
  wire s_csamul_cla32_fa14_2_xor0;
  wire s_csamul_cla32_fa14_2_and0;
  wire s_csamul_cla32_fa14_2_xor1;
  wire s_csamul_cla32_fa14_2_and1;
  wire s_csamul_cla32_fa14_2_or0;
  wire s_csamul_cla32_and15_2;
  wire s_csamul_cla32_fa15_2_xor0;
  wire s_csamul_cla32_fa15_2_and0;
  wire s_csamul_cla32_fa15_2_xor1;
  wire s_csamul_cla32_fa15_2_and1;
  wire s_csamul_cla32_fa15_2_or0;
  wire s_csamul_cla32_and16_2;
  wire s_csamul_cla32_fa16_2_xor0;
  wire s_csamul_cla32_fa16_2_and0;
  wire s_csamul_cla32_fa16_2_xor1;
  wire s_csamul_cla32_fa16_2_and1;
  wire s_csamul_cla32_fa16_2_or0;
  wire s_csamul_cla32_and17_2;
  wire s_csamul_cla32_fa17_2_xor0;
  wire s_csamul_cla32_fa17_2_and0;
  wire s_csamul_cla32_fa17_2_xor1;
  wire s_csamul_cla32_fa17_2_and1;
  wire s_csamul_cla32_fa17_2_or0;
  wire s_csamul_cla32_and18_2;
  wire s_csamul_cla32_fa18_2_xor0;
  wire s_csamul_cla32_fa18_2_and0;
  wire s_csamul_cla32_fa18_2_xor1;
  wire s_csamul_cla32_fa18_2_and1;
  wire s_csamul_cla32_fa18_2_or0;
  wire s_csamul_cla32_and19_2;
  wire s_csamul_cla32_fa19_2_xor0;
  wire s_csamul_cla32_fa19_2_and0;
  wire s_csamul_cla32_fa19_2_xor1;
  wire s_csamul_cla32_fa19_2_and1;
  wire s_csamul_cla32_fa19_2_or0;
  wire s_csamul_cla32_and20_2;
  wire s_csamul_cla32_fa20_2_xor0;
  wire s_csamul_cla32_fa20_2_and0;
  wire s_csamul_cla32_fa20_2_xor1;
  wire s_csamul_cla32_fa20_2_and1;
  wire s_csamul_cla32_fa20_2_or0;
  wire s_csamul_cla32_and21_2;
  wire s_csamul_cla32_fa21_2_xor0;
  wire s_csamul_cla32_fa21_2_and0;
  wire s_csamul_cla32_fa21_2_xor1;
  wire s_csamul_cla32_fa21_2_and1;
  wire s_csamul_cla32_fa21_2_or0;
  wire s_csamul_cla32_and22_2;
  wire s_csamul_cla32_fa22_2_xor0;
  wire s_csamul_cla32_fa22_2_and0;
  wire s_csamul_cla32_fa22_2_xor1;
  wire s_csamul_cla32_fa22_2_and1;
  wire s_csamul_cla32_fa22_2_or0;
  wire s_csamul_cla32_and23_2;
  wire s_csamul_cla32_fa23_2_xor0;
  wire s_csamul_cla32_fa23_2_and0;
  wire s_csamul_cla32_fa23_2_xor1;
  wire s_csamul_cla32_fa23_2_and1;
  wire s_csamul_cla32_fa23_2_or0;
  wire s_csamul_cla32_and24_2;
  wire s_csamul_cla32_fa24_2_xor0;
  wire s_csamul_cla32_fa24_2_and0;
  wire s_csamul_cla32_fa24_2_xor1;
  wire s_csamul_cla32_fa24_2_and1;
  wire s_csamul_cla32_fa24_2_or0;
  wire s_csamul_cla32_and25_2;
  wire s_csamul_cla32_fa25_2_xor0;
  wire s_csamul_cla32_fa25_2_and0;
  wire s_csamul_cla32_fa25_2_xor1;
  wire s_csamul_cla32_fa25_2_and1;
  wire s_csamul_cla32_fa25_2_or0;
  wire s_csamul_cla32_and26_2;
  wire s_csamul_cla32_fa26_2_xor0;
  wire s_csamul_cla32_fa26_2_and0;
  wire s_csamul_cla32_fa26_2_xor1;
  wire s_csamul_cla32_fa26_2_and1;
  wire s_csamul_cla32_fa26_2_or0;
  wire s_csamul_cla32_and27_2;
  wire s_csamul_cla32_fa27_2_xor0;
  wire s_csamul_cla32_fa27_2_and0;
  wire s_csamul_cla32_fa27_2_xor1;
  wire s_csamul_cla32_fa27_2_and1;
  wire s_csamul_cla32_fa27_2_or0;
  wire s_csamul_cla32_and28_2;
  wire s_csamul_cla32_fa28_2_xor0;
  wire s_csamul_cla32_fa28_2_and0;
  wire s_csamul_cla32_fa28_2_xor1;
  wire s_csamul_cla32_fa28_2_and1;
  wire s_csamul_cla32_fa28_2_or0;
  wire s_csamul_cla32_and29_2;
  wire s_csamul_cla32_fa29_2_xor0;
  wire s_csamul_cla32_fa29_2_and0;
  wire s_csamul_cla32_fa29_2_xor1;
  wire s_csamul_cla32_fa29_2_and1;
  wire s_csamul_cla32_fa29_2_or0;
  wire s_csamul_cla32_and30_2;
  wire s_csamul_cla32_fa30_2_xor0;
  wire s_csamul_cla32_fa30_2_and0;
  wire s_csamul_cla32_fa30_2_xor1;
  wire s_csamul_cla32_fa30_2_and1;
  wire s_csamul_cla32_fa30_2_or0;
  wire s_csamul_cla32_nand31_2;
  wire s_csamul_cla32_ha31_2_xor0;
  wire s_csamul_cla32_ha31_2_and0;
  wire s_csamul_cla32_and0_3;
  wire s_csamul_cla32_fa0_3_xor0;
  wire s_csamul_cla32_fa0_3_and0;
  wire s_csamul_cla32_fa0_3_xor1;
  wire s_csamul_cla32_fa0_3_and1;
  wire s_csamul_cla32_fa0_3_or0;
  wire s_csamul_cla32_and1_3;
  wire s_csamul_cla32_fa1_3_xor0;
  wire s_csamul_cla32_fa1_3_and0;
  wire s_csamul_cla32_fa1_3_xor1;
  wire s_csamul_cla32_fa1_3_and1;
  wire s_csamul_cla32_fa1_3_or0;
  wire s_csamul_cla32_and2_3;
  wire s_csamul_cla32_fa2_3_xor0;
  wire s_csamul_cla32_fa2_3_and0;
  wire s_csamul_cla32_fa2_3_xor1;
  wire s_csamul_cla32_fa2_3_and1;
  wire s_csamul_cla32_fa2_3_or0;
  wire s_csamul_cla32_and3_3;
  wire s_csamul_cla32_fa3_3_xor0;
  wire s_csamul_cla32_fa3_3_and0;
  wire s_csamul_cla32_fa3_3_xor1;
  wire s_csamul_cla32_fa3_3_and1;
  wire s_csamul_cla32_fa3_3_or0;
  wire s_csamul_cla32_and4_3;
  wire s_csamul_cla32_fa4_3_xor0;
  wire s_csamul_cla32_fa4_3_and0;
  wire s_csamul_cla32_fa4_3_xor1;
  wire s_csamul_cla32_fa4_3_and1;
  wire s_csamul_cla32_fa4_3_or0;
  wire s_csamul_cla32_and5_3;
  wire s_csamul_cla32_fa5_3_xor0;
  wire s_csamul_cla32_fa5_3_and0;
  wire s_csamul_cla32_fa5_3_xor1;
  wire s_csamul_cla32_fa5_3_and1;
  wire s_csamul_cla32_fa5_3_or0;
  wire s_csamul_cla32_and6_3;
  wire s_csamul_cla32_fa6_3_xor0;
  wire s_csamul_cla32_fa6_3_and0;
  wire s_csamul_cla32_fa6_3_xor1;
  wire s_csamul_cla32_fa6_3_and1;
  wire s_csamul_cla32_fa6_3_or0;
  wire s_csamul_cla32_and7_3;
  wire s_csamul_cla32_fa7_3_xor0;
  wire s_csamul_cla32_fa7_3_and0;
  wire s_csamul_cla32_fa7_3_xor1;
  wire s_csamul_cla32_fa7_3_and1;
  wire s_csamul_cla32_fa7_3_or0;
  wire s_csamul_cla32_and8_3;
  wire s_csamul_cla32_fa8_3_xor0;
  wire s_csamul_cla32_fa8_3_and0;
  wire s_csamul_cla32_fa8_3_xor1;
  wire s_csamul_cla32_fa8_3_and1;
  wire s_csamul_cla32_fa8_3_or0;
  wire s_csamul_cla32_and9_3;
  wire s_csamul_cla32_fa9_3_xor0;
  wire s_csamul_cla32_fa9_3_and0;
  wire s_csamul_cla32_fa9_3_xor1;
  wire s_csamul_cla32_fa9_3_and1;
  wire s_csamul_cla32_fa9_3_or0;
  wire s_csamul_cla32_and10_3;
  wire s_csamul_cla32_fa10_3_xor0;
  wire s_csamul_cla32_fa10_3_and0;
  wire s_csamul_cla32_fa10_3_xor1;
  wire s_csamul_cla32_fa10_3_and1;
  wire s_csamul_cla32_fa10_3_or0;
  wire s_csamul_cla32_and11_3;
  wire s_csamul_cla32_fa11_3_xor0;
  wire s_csamul_cla32_fa11_3_and0;
  wire s_csamul_cla32_fa11_3_xor1;
  wire s_csamul_cla32_fa11_3_and1;
  wire s_csamul_cla32_fa11_3_or0;
  wire s_csamul_cla32_and12_3;
  wire s_csamul_cla32_fa12_3_xor0;
  wire s_csamul_cla32_fa12_3_and0;
  wire s_csamul_cla32_fa12_3_xor1;
  wire s_csamul_cla32_fa12_3_and1;
  wire s_csamul_cla32_fa12_3_or0;
  wire s_csamul_cla32_and13_3;
  wire s_csamul_cla32_fa13_3_xor0;
  wire s_csamul_cla32_fa13_3_and0;
  wire s_csamul_cla32_fa13_3_xor1;
  wire s_csamul_cla32_fa13_3_and1;
  wire s_csamul_cla32_fa13_3_or0;
  wire s_csamul_cla32_and14_3;
  wire s_csamul_cla32_fa14_3_xor0;
  wire s_csamul_cla32_fa14_3_and0;
  wire s_csamul_cla32_fa14_3_xor1;
  wire s_csamul_cla32_fa14_3_and1;
  wire s_csamul_cla32_fa14_3_or0;
  wire s_csamul_cla32_and15_3;
  wire s_csamul_cla32_fa15_3_xor0;
  wire s_csamul_cla32_fa15_3_and0;
  wire s_csamul_cla32_fa15_3_xor1;
  wire s_csamul_cla32_fa15_3_and1;
  wire s_csamul_cla32_fa15_3_or0;
  wire s_csamul_cla32_and16_3;
  wire s_csamul_cla32_fa16_3_xor0;
  wire s_csamul_cla32_fa16_3_and0;
  wire s_csamul_cla32_fa16_3_xor1;
  wire s_csamul_cla32_fa16_3_and1;
  wire s_csamul_cla32_fa16_3_or0;
  wire s_csamul_cla32_and17_3;
  wire s_csamul_cla32_fa17_3_xor0;
  wire s_csamul_cla32_fa17_3_and0;
  wire s_csamul_cla32_fa17_3_xor1;
  wire s_csamul_cla32_fa17_3_and1;
  wire s_csamul_cla32_fa17_3_or0;
  wire s_csamul_cla32_and18_3;
  wire s_csamul_cla32_fa18_3_xor0;
  wire s_csamul_cla32_fa18_3_and0;
  wire s_csamul_cla32_fa18_3_xor1;
  wire s_csamul_cla32_fa18_3_and1;
  wire s_csamul_cla32_fa18_3_or0;
  wire s_csamul_cla32_and19_3;
  wire s_csamul_cla32_fa19_3_xor0;
  wire s_csamul_cla32_fa19_3_and0;
  wire s_csamul_cla32_fa19_3_xor1;
  wire s_csamul_cla32_fa19_3_and1;
  wire s_csamul_cla32_fa19_3_or0;
  wire s_csamul_cla32_and20_3;
  wire s_csamul_cla32_fa20_3_xor0;
  wire s_csamul_cla32_fa20_3_and0;
  wire s_csamul_cla32_fa20_3_xor1;
  wire s_csamul_cla32_fa20_3_and1;
  wire s_csamul_cla32_fa20_3_or0;
  wire s_csamul_cla32_and21_3;
  wire s_csamul_cla32_fa21_3_xor0;
  wire s_csamul_cla32_fa21_3_and0;
  wire s_csamul_cla32_fa21_3_xor1;
  wire s_csamul_cla32_fa21_3_and1;
  wire s_csamul_cla32_fa21_3_or0;
  wire s_csamul_cla32_and22_3;
  wire s_csamul_cla32_fa22_3_xor0;
  wire s_csamul_cla32_fa22_3_and0;
  wire s_csamul_cla32_fa22_3_xor1;
  wire s_csamul_cla32_fa22_3_and1;
  wire s_csamul_cla32_fa22_3_or0;
  wire s_csamul_cla32_and23_3;
  wire s_csamul_cla32_fa23_3_xor0;
  wire s_csamul_cla32_fa23_3_and0;
  wire s_csamul_cla32_fa23_3_xor1;
  wire s_csamul_cla32_fa23_3_and1;
  wire s_csamul_cla32_fa23_3_or0;
  wire s_csamul_cla32_and24_3;
  wire s_csamul_cla32_fa24_3_xor0;
  wire s_csamul_cla32_fa24_3_and0;
  wire s_csamul_cla32_fa24_3_xor1;
  wire s_csamul_cla32_fa24_3_and1;
  wire s_csamul_cla32_fa24_3_or0;
  wire s_csamul_cla32_and25_3;
  wire s_csamul_cla32_fa25_3_xor0;
  wire s_csamul_cla32_fa25_3_and0;
  wire s_csamul_cla32_fa25_3_xor1;
  wire s_csamul_cla32_fa25_3_and1;
  wire s_csamul_cla32_fa25_3_or0;
  wire s_csamul_cla32_and26_3;
  wire s_csamul_cla32_fa26_3_xor0;
  wire s_csamul_cla32_fa26_3_and0;
  wire s_csamul_cla32_fa26_3_xor1;
  wire s_csamul_cla32_fa26_3_and1;
  wire s_csamul_cla32_fa26_3_or0;
  wire s_csamul_cla32_and27_3;
  wire s_csamul_cla32_fa27_3_xor0;
  wire s_csamul_cla32_fa27_3_and0;
  wire s_csamul_cla32_fa27_3_xor1;
  wire s_csamul_cla32_fa27_3_and1;
  wire s_csamul_cla32_fa27_3_or0;
  wire s_csamul_cla32_and28_3;
  wire s_csamul_cla32_fa28_3_xor0;
  wire s_csamul_cla32_fa28_3_and0;
  wire s_csamul_cla32_fa28_3_xor1;
  wire s_csamul_cla32_fa28_3_and1;
  wire s_csamul_cla32_fa28_3_or0;
  wire s_csamul_cla32_and29_3;
  wire s_csamul_cla32_fa29_3_xor0;
  wire s_csamul_cla32_fa29_3_and0;
  wire s_csamul_cla32_fa29_3_xor1;
  wire s_csamul_cla32_fa29_3_and1;
  wire s_csamul_cla32_fa29_3_or0;
  wire s_csamul_cla32_and30_3;
  wire s_csamul_cla32_fa30_3_xor0;
  wire s_csamul_cla32_fa30_3_and0;
  wire s_csamul_cla32_fa30_3_xor1;
  wire s_csamul_cla32_fa30_3_and1;
  wire s_csamul_cla32_fa30_3_or0;
  wire s_csamul_cla32_nand31_3;
  wire s_csamul_cla32_ha31_3_xor0;
  wire s_csamul_cla32_ha31_3_and0;
  wire s_csamul_cla32_and0_4;
  wire s_csamul_cla32_fa0_4_xor0;
  wire s_csamul_cla32_fa0_4_and0;
  wire s_csamul_cla32_fa0_4_xor1;
  wire s_csamul_cla32_fa0_4_and1;
  wire s_csamul_cla32_fa0_4_or0;
  wire s_csamul_cla32_and1_4;
  wire s_csamul_cla32_fa1_4_xor0;
  wire s_csamul_cla32_fa1_4_and0;
  wire s_csamul_cla32_fa1_4_xor1;
  wire s_csamul_cla32_fa1_4_and1;
  wire s_csamul_cla32_fa1_4_or0;
  wire s_csamul_cla32_and2_4;
  wire s_csamul_cla32_fa2_4_xor0;
  wire s_csamul_cla32_fa2_4_and0;
  wire s_csamul_cla32_fa2_4_xor1;
  wire s_csamul_cla32_fa2_4_and1;
  wire s_csamul_cla32_fa2_4_or0;
  wire s_csamul_cla32_and3_4;
  wire s_csamul_cla32_fa3_4_xor0;
  wire s_csamul_cla32_fa3_4_and0;
  wire s_csamul_cla32_fa3_4_xor1;
  wire s_csamul_cla32_fa3_4_and1;
  wire s_csamul_cla32_fa3_4_or0;
  wire s_csamul_cla32_and4_4;
  wire s_csamul_cla32_fa4_4_xor0;
  wire s_csamul_cla32_fa4_4_and0;
  wire s_csamul_cla32_fa4_4_xor1;
  wire s_csamul_cla32_fa4_4_and1;
  wire s_csamul_cla32_fa4_4_or0;
  wire s_csamul_cla32_and5_4;
  wire s_csamul_cla32_fa5_4_xor0;
  wire s_csamul_cla32_fa5_4_and0;
  wire s_csamul_cla32_fa5_4_xor1;
  wire s_csamul_cla32_fa5_4_and1;
  wire s_csamul_cla32_fa5_4_or0;
  wire s_csamul_cla32_and6_4;
  wire s_csamul_cla32_fa6_4_xor0;
  wire s_csamul_cla32_fa6_4_and0;
  wire s_csamul_cla32_fa6_4_xor1;
  wire s_csamul_cla32_fa6_4_and1;
  wire s_csamul_cla32_fa6_4_or0;
  wire s_csamul_cla32_and7_4;
  wire s_csamul_cla32_fa7_4_xor0;
  wire s_csamul_cla32_fa7_4_and0;
  wire s_csamul_cla32_fa7_4_xor1;
  wire s_csamul_cla32_fa7_4_and1;
  wire s_csamul_cla32_fa7_4_or0;
  wire s_csamul_cla32_and8_4;
  wire s_csamul_cla32_fa8_4_xor0;
  wire s_csamul_cla32_fa8_4_and0;
  wire s_csamul_cla32_fa8_4_xor1;
  wire s_csamul_cla32_fa8_4_and1;
  wire s_csamul_cla32_fa8_4_or0;
  wire s_csamul_cla32_and9_4;
  wire s_csamul_cla32_fa9_4_xor0;
  wire s_csamul_cla32_fa9_4_and0;
  wire s_csamul_cla32_fa9_4_xor1;
  wire s_csamul_cla32_fa9_4_and1;
  wire s_csamul_cla32_fa9_4_or0;
  wire s_csamul_cla32_and10_4;
  wire s_csamul_cla32_fa10_4_xor0;
  wire s_csamul_cla32_fa10_4_and0;
  wire s_csamul_cla32_fa10_4_xor1;
  wire s_csamul_cla32_fa10_4_and1;
  wire s_csamul_cla32_fa10_4_or0;
  wire s_csamul_cla32_and11_4;
  wire s_csamul_cla32_fa11_4_xor0;
  wire s_csamul_cla32_fa11_4_and0;
  wire s_csamul_cla32_fa11_4_xor1;
  wire s_csamul_cla32_fa11_4_and1;
  wire s_csamul_cla32_fa11_4_or0;
  wire s_csamul_cla32_and12_4;
  wire s_csamul_cla32_fa12_4_xor0;
  wire s_csamul_cla32_fa12_4_and0;
  wire s_csamul_cla32_fa12_4_xor1;
  wire s_csamul_cla32_fa12_4_and1;
  wire s_csamul_cla32_fa12_4_or0;
  wire s_csamul_cla32_and13_4;
  wire s_csamul_cla32_fa13_4_xor0;
  wire s_csamul_cla32_fa13_4_and0;
  wire s_csamul_cla32_fa13_4_xor1;
  wire s_csamul_cla32_fa13_4_and1;
  wire s_csamul_cla32_fa13_4_or0;
  wire s_csamul_cla32_and14_4;
  wire s_csamul_cla32_fa14_4_xor0;
  wire s_csamul_cla32_fa14_4_and0;
  wire s_csamul_cla32_fa14_4_xor1;
  wire s_csamul_cla32_fa14_4_and1;
  wire s_csamul_cla32_fa14_4_or0;
  wire s_csamul_cla32_and15_4;
  wire s_csamul_cla32_fa15_4_xor0;
  wire s_csamul_cla32_fa15_4_and0;
  wire s_csamul_cla32_fa15_4_xor1;
  wire s_csamul_cla32_fa15_4_and1;
  wire s_csamul_cla32_fa15_4_or0;
  wire s_csamul_cla32_and16_4;
  wire s_csamul_cla32_fa16_4_xor0;
  wire s_csamul_cla32_fa16_4_and0;
  wire s_csamul_cla32_fa16_4_xor1;
  wire s_csamul_cla32_fa16_4_and1;
  wire s_csamul_cla32_fa16_4_or0;
  wire s_csamul_cla32_and17_4;
  wire s_csamul_cla32_fa17_4_xor0;
  wire s_csamul_cla32_fa17_4_and0;
  wire s_csamul_cla32_fa17_4_xor1;
  wire s_csamul_cla32_fa17_4_and1;
  wire s_csamul_cla32_fa17_4_or0;
  wire s_csamul_cla32_and18_4;
  wire s_csamul_cla32_fa18_4_xor0;
  wire s_csamul_cla32_fa18_4_and0;
  wire s_csamul_cla32_fa18_4_xor1;
  wire s_csamul_cla32_fa18_4_and1;
  wire s_csamul_cla32_fa18_4_or0;
  wire s_csamul_cla32_and19_4;
  wire s_csamul_cla32_fa19_4_xor0;
  wire s_csamul_cla32_fa19_4_and0;
  wire s_csamul_cla32_fa19_4_xor1;
  wire s_csamul_cla32_fa19_4_and1;
  wire s_csamul_cla32_fa19_4_or0;
  wire s_csamul_cla32_and20_4;
  wire s_csamul_cla32_fa20_4_xor0;
  wire s_csamul_cla32_fa20_4_and0;
  wire s_csamul_cla32_fa20_4_xor1;
  wire s_csamul_cla32_fa20_4_and1;
  wire s_csamul_cla32_fa20_4_or0;
  wire s_csamul_cla32_and21_4;
  wire s_csamul_cla32_fa21_4_xor0;
  wire s_csamul_cla32_fa21_4_and0;
  wire s_csamul_cla32_fa21_4_xor1;
  wire s_csamul_cla32_fa21_4_and1;
  wire s_csamul_cla32_fa21_4_or0;
  wire s_csamul_cla32_and22_4;
  wire s_csamul_cla32_fa22_4_xor0;
  wire s_csamul_cla32_fa22_4_and0;
  wire s_csamul_cla32_fa22_4_xor1;
  wire s_csamul_cla32_fa22_4_and1;
  wire s_csamul_cla32_fa22_4_or0;
  wire s_csamul_cla32_and23_4;
  wire s_csamul_cla32_fa23_4_xor0;
  wire s_csamul_cla32_fa23_4_and0;
  wire s_csamul_cla32_fa23_4_xor1;
  wire s_csamul_cla32_fa23_4_and1;
  wire s_csamul_cla32_fa23_4_or0;
  wire s_csamul_cla32_and24_4;
  wire s_csamul_cla32_fa24_4_xor0;
  wire s_csamul_cla32_fa24_4_and0;
  wire s_csamul_cla32_fa24_4_xor1;
  wire s_csamul_cla32_fa24_4_and1;
  wire s_csamul_cla32_fa24_4_or0;
  wire s_csamul_cla32_and25_4;
  wire s_csamul_cla32_fa25_4_xor0;
  wire s_csamul_cla32_fa25_4_and0;
  wire s_csamul_cla32_fa25_4_xor1;
  wire s_csamul_cla32_fa25_4_and1;
  wire s_csamul_cla32_fa25_4_or0;
  wire s_csamul_cla32_and26_4;
  wire s_csamul_cla32_fa26_4_xor0;
  wire s_csamul_cla32_fa26_4_and0;
  wire s_csamul_cla32_fa26_4_xor1;
  wire s_csamul_cla32_fa26_4_and1;
  wire s_csamul_cla32_fa26_4_or0;
  wire s_csamul_cla32_and27_4;
  wire s_csamul_cla32_fa27_4_xor0;
  wire s_csamul_cla32_fa27_4_and0;
  wire s_csamul_cla32_fa27_4_xor1;
  wire s_csamul_cla32_fa27_4_and1;
  wire s_csamul_cla32_fa27_4_or0;
  wire s_csamul_cla32_and28_4;
  wire s_csamul_cla32_fa28_4_xor0;
  wire s_csamul_cla32_fa28_4_and0;
  wire s_csamul_cla32_fa28_4_xor1;
  wire s_csamul_cla32_fa28_4_and1;
  wire s_csamul_cla32_fa28_4_or0;
  wire s_csamul_cla32_and29_4;
  wire s_csamul_cla32_fa29_4_xor0;
  wire s_csamul_cla32_fa29_4_and0;
  wire s_csamul_cla32_fa29_4_xor1;
  wire s_csamul_cla32_fa29_4_and1;
  wire s_csamul_cla32_fa29_4_or0;
  wire s_csamul_cla32_and30_4;
  wire s_csamul_cla32_fa30_4_xor0;
  wire s_csamul_cla32_fa30_4_and0;
  wire s_csamul_cla32_fa30_4_xor1;
  wire s_csamul_cla32_fa30_4_and1;
  wire s_csamul_cla32_fa30_4_or0;
  wire s_csamul_cla32_nand31_4;
  wire s_csamul_cla32_ha31_4_xor0;
  wire s_csamul_cla32_ha31_4_and0;
  wire s_csamul_cla32_and0_5;
  wire s_csamul_cla32_fa0_5_xor0;
  wire s_csamul_cla32_fa0_5_and0;
  wire s_csamul_cla32_fa0_5_xor1;
  wire s_csamul_cla32_fa0_5_and1;
  wire s_csamul_cla32_fa0_5_or0;
  wire s_csamul_cla32_and1_5;
  wire s_csamul_cla32_fa1_5_xor0;
  wire s_csamul_cla32_fa1_5_and0;
  wire s_csamul_cla32_fa1_5_xor1;
  wire s_csamul_cla32_fa1_5_and1;
  wire s_csamul_cla32_fa1_5_or0;
  wire s_csamul_cla32_and2_5;
  wire s_csamul_cla32_fa2_5_xor0;
  wire s_csamul_cla32_fa2_5_and0;
  wire s_csamul_cla32_fa2_5_xor1;
  wire s_csamul_cla32_fa2_5_and1;
  wire s_csamul_cla32_fa2_5_or0;
  wire s_csamul_cla32_and3_5;
  wire s_csamul_cla32_fa3_5_xor0;
  wire s_csamul_cla32_fa3_5_and0;
  wire s_csamul_cla32_fa3_5_xor1;
  wire s_csamul_cla32_fa3_5_and1;
  wire s_csamul_cla32_fa3_5_or0;
  wire s_csamul_cla32_and4_5;
  wire s_csamul_cla32_fa4_5_xor0;
  wire s_csamul_cla32_fa4_5_and0;
  wire s_csamul_cla32_fa4_5_xor1;
  wire s_csamul_cla32_fa4_5_and1;
  wire s_csamul_cla32_fa4_5_or0;
  wire s_csamul_cla32_and5_5;
  wire s_csamul_cla32_fa5_5_xor0;
  wire s_csamul_cla32_fa5_5_and0;
  wire s_csamul_cla32_fa5_5_xor1;
  wire s_csamul_cla32_fa5_5_and1;
  wire s_csamul_cla32_fa5_5_or0;
  wire s_csamul_cla32_and6_5;
  wire s_csamul_cla32_fa6_5_xor0;
  wire s_csamul_cla32_fa6_5_and0;
  wire s_csamul_cla32_fa6_5_xor1;
  wire s_csamul_cla32_fa6_5_and1;
  wire s_csamul_cla32_fa6_5_or0;
  wire s_csamul_cla32_and7_5;
  wire s_csamul_cla32_fa7_5_xor0;
  wire s_csamul_cla32_fa7_5_and0;
  wire s_csamul_cla32_fa7_5_xor1;
  wire s_csamul_cla32_fa7_5_and1;
  wire s_csamul_cla32_fa7_5_or0;
  wire s_csamul_cla32_and8_5;
  wire s_csamul_cla32_fa8_5_xor0;
  wire s_csamul_cla32_fa8_5_and0;
  wire s_csamul_cla32_fa8_5_xor1;
  wire s_csamul_cla32_fa8_5_and1;
  wire s_csamul_cla32_fa8_5_or0;
  wire s_csamul_cla32_and9_5;
  wire s_csamul_cla32_fa9_5_xor0;
  wire s_csamul_cla32_fa9_5_and0;
  wire s_csamul_cla32_fa9_5_xor1;
  wire s_csamul_cla32_fa9_5_and1;
  wire s_csamul_cla32_fa9_5_or0;
  wire s_csamul_cla32_and10_5;
  wire s_csamul_cla32_fa10_5_xor0;
  wire s_csamul_cla32_fa10_5_and0;
  wire s_csamul_cla32_fa10_5_xor1;
  wire s_csamul_cla32_fa10_5_and1;
  wire s_csamul_cla32_fa10_5_or0;
  wire s_csamul_cla32_and11_5;
  wire s_csamul_cla32_fa11_5_xor0;
  wire s_csamul_cla32_fa11_5_and0;
  wire s_csamul_cla32_fa11_5_xor1;
  wire s_csamul_cla32_fa11_5_and1;
  wire s_csamul_cla32_fa11_5_or0;
  wire s_csamul_cla32_and12_5;
  wire s_csamul_cla32_fa12_5_xor0;
  wire s_csamul_cla32_fa12_5_and0;
  wire s_csamul_cla32_fa12_5_xor1;
  wire s_csamul_cla32_fa12_5_and1;
  wire s_csamul_cla32_fa12_5_or0;
  wire s_csamul_cla32_and13_5;
  wire s_csamul_cla32_fa13_5_xor0;
  wire s_csamul_cla32_fa13_5_and0;
  wire s_csamul_cla32_fa13_5_xor1;
  wire s_csamul_cla32_fa13_5_and1;
  wire s_csamul_cla32_fa13_5_or0;
  wire s_csamul_cla32_and14_5;
  wire s_csamul_cla32_fa14_5_xor0;
  wire s_csamul_cla32_fa14_5_and0;
  wire s_csamul_cla32_fa14_5_xor1;
  wire s_csamul_cla32_fa14_5_and1;
  wire s_csamul_cla32_fa14_5_or0;
  wire s_csamul_cla32_and15_5;
  wire s_csamul_cla32_fa15_5_xor0;
  wire s_csamul_cla32_fa15_5_and0;
  wire s_csamul_cla32_fa15_5_xor1;
  wire s_csamul_cla32_fa15_5_and1;
  wire s_csamul_cla32_fa15_5_or0;
  wire s_csamul_cla32_and16_5;
  wire s_csamul_cla32_fa16_5_xor0;
  wire s_csamul_cla32_fa16_5_and0;
  wire s_csamul_cla32_fa16_5_xor1;
  wire s_csamul_cla32_fa16_5_and1;
  wire s_csamul_cla32_fa16_5_or0;
  wire s_csamul_cla32_and17_5;
  wire s_csamul_cla32_fa17_5_xor0;
  wire s_csamul_cla32_fa17_5_and0;
  wire s_csamul_cla32_fa17_5_xor1;
  wire s_csamul_cla32_fa17_5_and1;
  wire s_csamul_cla32_fa17_5_or0;
  wire s_csamul_cla32_and18_5;
  wire s_csamul_cla32_fa18_5_xor0;
  wire s_csamul_cla32_fa18_5_and0;
  wire s_csamul_cla32_fa18_5_xor1;
  wire s_csamul_cla32_fa18_5_and1;
  wire s_csamul_cla32_fa18_5_or0;
  wire s_csamul_cla32_and19_5;
  wire s_csamul_cla32_fa19_5_xor0;
  wire s_csamul_cla32_fa19_5_and0;
  wire s_csamul_cla32_fa19_5_xor1;
  wire s_csamul_cla32_fa19_5_and1;
  wire s_csamul_cla32_fa19_5_or0;
  wire s_csamul_cla32_and20_5;
  wire s_csamul_cla32_fa20_5_xor0;
  wire s_csamul_cla32_fa20_5_and0;
  wire s_csamul_cla32_fa20_5_xor1;
  wire s_csamul_cla32_fa20_5_and1;
  wire s_csamul_cla32_fa20_5_or0;
  wire s_csamul_cla32_and21_5;
  wire s_csamul_cla32_fa21_5_xor0;
  wire s_csamul_cla32_fa21_5_and0;
  wire s_csamul_cla32_fa21_5_xor1;
  wire s_csamul_cla32_fa21_5_and1;
  wire s_csamul_cla32_fa21_5_or0;
  wire s_csamul_cla32_and22_5;
  wire s_csamul_cla32_fa22_5_xor0;
  wire s_csamul_cla32_fa22_5_and0;
  wire s_csamul_cla32_fa22_5_xor1;
  wire s_csamul_cla32_fa22_5_and1;
  wire s_csamul_cla32_fa22_5_or0;
  wire s_csamul_cla32_and23_5;
  wire s_csamul_cla32_fa23_5_xor0;
  wire s_csamul_cla32_fa23_5_and0;
  wire s_csamul_cla32_fa23_5_xor1;
  wire s_csamul_cla32_fa23_5_and1;
  wire s_csamul_cla32_fa23_5_or0;
  wire s_csamul_cla32_and24_5;
  wire s_csamul_cla32_fa24_5_xor0;
  wire s_csamul_cla32_fa24_5_and0;
  wire s_csamul_cla32_fa24_5_xor1;
  wire s_csamul_cla32_fa24_5_and1;
  wire s_csamul_cla32_fa24_5_or0;
  wire s_csamul_cla32_and25_5;
  wire s_csamul_cla32_fa25_5_xor0;
  wire s_csamul_cla32_fa25_5_and0;
  wire s_csamul_cla32_fa25_5_xor1;
  wire s_csamul_cla32_fa25_5_and1;
  wire s_csamul_cla32_fa25_5_or0;
  wire s_csamul_cla32_and26_5;
  wire s_csamul_cla32_fa26_5_xor0;
  wire s_csamul_cla32_fa26_5_and0;
  wire s_csamul_cla32_fa26_5_xor1;
  wire s_csamul_cla32_fa26_5_and1;
  wire s_csamul_cla32_fa26_5_or0;
  wire s_csamul_cla32_and27_5;
  wire s_csamul_cla32_fa27_5_xor0;
  wire s_csamul_cla32_fa27_5_and0;
  wire s_csamul_cla32_fa27_5_xor1;
  wire s_csamul_cla32_fa27_5_and1;
  wire s_csamul_cla32_fa27_5_or0;
  wire s_csamul_cla32_and28_5;
  wire s_csamul_cla32_fa28_5_xor0;
  wire s_csamul_cla32_fa28_5_and0;
  wire s_csamul_cla32_fa28_5_xor1;
  wire s_csamul_cla32_fa28_5_and1;
  wire s_csamul_cla32_fa28_5_or0;
  wire s_csamul_cla32_and29_5;
  wire s_csamul_cla32_fa29_5_xor0;
  wire s_csamul_cla32_fa29_5_and0;
  wire s_csamul_cla32_fa29_5_xor1;
  wire s_csamul_cla32_fa29_5_and1;
  wire s_csamul_cla32_fa29_5_or0;
  wire s_csamul_cla32_and30_5;
  wire s_csamul_cla32_fa30_5_xor0;
  wire s_csamul_cla32_fa30_5_and0;
  wire s_csamul_cla32_fa30_5_xor1;
  wire s_csamul_cla32_fa30_5_and1;
  wire s_csamul_cla32_fa30_5_or0;
  wire s_csamul_cla32_nand31_5;
  wire s_csamul_cla32_ha31_5_xor0;
  wire s_csamul_cla32_ha31_5_and0;
  wire s_csamul_cla32_and0_6;
  wire s_csamul_cla32_fa0_6_xor0;
  wire s_csamul_cla32_fa0_6_and0;
  wire s_csamul_cla32_fa0_6_xor1;
  wire s_csamul_cla32_fa0_6_and1;
  wire s_csamul_cla32_fa0_6_or0;
  wire s_csamul_cla32_and1_6;
  wire s_csamul_cla32_fa1_6_xor0;
  wire s_csamul_cla32_fa1_6_and0;
  wire s_csamul_cla32_fa1_6_xor1;
  wire s_csamul_cla32_fa1_6_and1;
  wire s_csamul_cla32_fa1_6_or0;
  wire s_csamul_cla32_and2_6;
  wire s_csamul_cla32_fa2_6_xor0;
  wire s_csamul_cla32_fa2_6_and0;
  wire s_csamul_cla32_fa2_6_xor1;
  wire s_csamul_cla32_fa2_6_and1;
  wire s_csamul_cla32_fa2_6_or0;
  wire s_csamul_cla32_and3_6;
  wire s_csamul_cla32_fa3_6_xor0;
  wire s_csamul_cla32_fa3_6_and0;
  wire s_csamul_cla32_fa3_6_xor1;
  wire s_csamul_cla32_fa3_6_and1;
  wire s_csamul_cla32_fa3_6_or0;
  wire s_csamul_cla32_and4_6;
  wire s_csamul_cla32_fa4_6_xor0;
  wire s_csamul_cla32_fa4_6_and0;
  wire s_csamul_cla32_fa4_6_xor1;
  wire s_csamul_cla32_fa4_6_and1;
  wire s_csamul_cla32_fa4_6_or0;
  wire s_csamul_cla32_and5_6;
  wire s_csamul_cla32_fa5_6_xor0;
  wire s_csamul_cla32_fa5_6_and0;
  wire s_csamul_cla32_fa5_6_xor1;
  wire s_csamul_cla32_fa5_6_and1;
  wire s_csamul_cla32_fa5_6_or0;
  wire s_csamul_cla32_and6_6;
  wire s_csamul_cla32_fa6_6_xor0;
  wire s_csamul_cla32_fa6_6_and0;
  wire s_csamul_cla32_fa6_6_xor1;
  wire s_csamul_cla32_fa6_6_and1;
  wire s_csamul_cla32_fa6_6_or0;
  wire s_csamul_cla32_and7_6;
  wire s_csamul_cla32_fa7_6_xor0;
  wire s_csamul_cla32_fa7_6_and0;
  wire s_csamul_cla32_fa7_6_xor1;
  wire s_csamul_cla32_fa7_6_and1;
  wire s_csamul_cla32_fa7_6_or0;
  wire s_csamul_cla32_and8_6;
  wire s_csamul_cla32_fa8_6_xor0;
  wire s_csamul_cla32_fa8_6_and0;
  wire s_csamul_cla32_fa8_6_xor1;
  wire s_csamul_cla32_fa8_6_and1;
  wire s_csamul_cla32_fa8_6_or0;
  wire s_csamul_cla32_and9_6;
  wire s_csamul_cla32_fa9_6_xor0;
  wire s_csamul_cla32_fa9_6_and0;
  wire s_csamul_cla32_fa9_6_xor1;
  wire s_csamul_cla32_fa9_6_and1;
  wire s_csamul_cla32_fa9_6_or0;
  wire s_csamul_cla32_and10_6;
  wire s_csamul_cla32_fa10_6_xor0;
  wire s_csamul_cla32_fa10_6_and0;
  wire s_csamul_cla32_fa10_6_xor1;
  wire s_csamul_cla32_fa10_6_and1;
  wire s_csamul_cla32_fa10_6_or0;
  wire s_csamul_cla32_and11_6;
  wire s_csamul_cla32_fa11_6_xor0;
  wire s_csamul_cla32_fa11_6_and0;
  wire s_csamul_cla32_fa11_6_xor1;
  wire s_csamul_cla32_fa11_6_and1;
  wire s_csamul_cla32_fa11_6_or0;
  wire s_csamul_cla32_and12_6;
  wire s_csamul_cla32_fa12_6_xor0;
  wire s_csamul_cla32_fa12_6_and0;
  wire s_csamul_cla32_fa12_6_xor1;
  wire s_csamul_cla32_fa12_6_and1;
  wire s_csamul_cla32_fa12_6_or0;
  wire s_csamul_cla32_and13_6;
  wire s_csamul_cla32_fa13_6_xor0;
  wire s_csamul_cla32_fa13_6_and0;
  wire s_csamul_cla32_fa13_6_xor1;
  wire s_csamul_cla32_fa13_6_and1;
  wire s_csamul_cla32_fa13_6_or0;
  wire s_csamul_cla32_and14_6;
  wire s_csamul_cla32_fa14_6_xor0;
  wire s_csamul_cla32_fa14_6_and0;
  wire s_csamul_cla32_fa14_6_xor1;
  wire s_csamul_cla32_fa14_6_and1;
  wire s_csamul_cla32_fa14_6_or0;
  wire s_csamul_cla32_and15_6;
  wire s_csamul_cla32_fa15_6_xor0;
  wire s_csamul_cla32_fa15_6_and0;
  wire s_csamul_cla32_fa15_6_xor1;
  wire s_csamul_cla32_fa15_6_and1;
  wire s_csamul_cla32_fa15_6_or0;
  wire s_csamul_cla32_and16_6;
  wire s_csamul_cla32_fa16_6_xor0;
  wire s_csamul_cla32_fa16_6_and0;
  wire s_csamul_cla32_fa16_6_xor1;
  wire s_csamul_cla32_fa16_6_and1;
  wire s_csamul_cla32_fa16_6_or0;
  wire s_csamul_cla32_and17_6;
  wire s_csamul_cla32_fa17_6_xor0;
  wire s_csamul_cla32_fa17_6_and0;
  wire s_csamul_cla32_fa17_6_xor1;
  wire s_csamul_cla32_fa17_6_and1;
  wire s_csamul_cla32_fa17_6_or0;
  wire s_csamul_cla32_and18_6;
  wire s_csamul_cla32_fa18_6_xor0;
  wire s_csamul_cla32_fa18_6_and0;
  wire s_csamul_cla32_fa18_6_xor1;
  wire s_csamul_cla32_fa18_6_and1;
  wire s_csamul_cla32_fa18_6_or0;
  wire s_csamul_cla32_and19_6;
  wire s_csamul_cla32_fa19_6_xor0;
  wire s_csamul_cla32_fa19_6_and0;
  wire s_csamul_cla32_fa19_6_xor1;
  wire s_csamul_cla32_fa19_6_and1;
  wire s_csamul_cla32_fa19_6_or0;
  wire s_csamul_cla32_and20_6;
  wire s_csamul_cla32_fa20_6_xor0;
  wire s_csamul_cla32_fa20_6_and0;
  wire s_csamul_cla32_fa20_6_xor1;
  wire s_csamul_cla32_fa20_6_and1;
  wire s_csamul_cla32_fa20_6_or0;
  wire s_csamul_cla32_and21_6;
  wire s_csamul_cla32_fa21_6_xor0;
  wire s_csamul_cla32_fa21_6_and0;
  wire s_csamul_cla32_fa21_6_xor1;
  wire s_csamul_cla32_fa21_6_and1;
  wire s_csamul_cla32_fa21_6_or0;
  wire s_csamul_cla32_and22_6;
  wire s_csamul_cla32_fa22_6_xor0;
  wire s_csamul_cla32_fa22_6_and0;
  wire s_csamul_cla32_fa22_6_xor1;
  wire s_csamul_cla32_fa22_6_and1;
  wire s_csamul_cla32_fa22_6_or0;
  wire s_csamul_cla32_and23_6;
  wire s_csamul_cla32_fa23_6_xor0;
  wire s_csamul_cla32_fa23_6_and0;
  wire s_csamul_cla32_fa23_6_xor1;
  wire s_csamul_cla32_fa23_6_and1;
  wire s_csamul_cla32_fa23_6_or0;
  wire s_csamul_cla32_and24_6;
  wire s_csamul_cla32_fa24_6_xor0;
  wire s_csamul_cla32_fa24_6_and0;
  wire s_csamul_cla32_fa24_6_xor1;
  wire s_csamul_cla32_fa24_6_and1;
  wire s_csamul_cla32_fa24_6_or0;
  wire s_csamul_cla32_and25_6;
  wire s_csamul_cla32_fa25_6_xor0;
  wire s_csamul_cla32_fa25_6_and0;
  wire s_csamul_cla32_fa25_6_xor1;
  wire s_csamul_cla32_fa25_6_and1;
  wire s_csamul_cla32_fa25_6_or0;
  wire s_csamul_cla32_and26_6;
  wire s_csamul_cla32_fa26_6_xor0;
  wire s_csamul_cla32_fa26_6_and0;
  wire s_csamul_cla32_fa26_6_xor1;
  wire s_csamul_cla32_fa26_6_and1;
  wire s_csamul_cla32_fa26_6_or0;
  wire s_csamul_cla32_and27_6;
  wire s_csamul_cla32_fa27_6_xor0;
  wire s_csamul_cla32_fa27_6_and0;
  wire s_csamul_cla32_fa27_6_xor1;
  wire s_csamul_cla32_fa27_6_and1;
  wire s_csamul_cla32_fa27_6_or0;
  wire s_csamul_cla32_and28_6;
  wire s_csamul_cla32_fa28_6_xor0;
  wire s_csamul_cla32_fa28_6_and0;
  wire s_csamul_cla32_fa28_6_xor1;
  wire s_csamul_cla32_fa28_6_and1;
  wire s_csamul_cla32_fa28_6_or0;
  wire s_csamul_cla32_and29_6;
  wire s_csamul_cla32_fa29_6_xor0;
  wire s_csamul_cla32_fa29_6_and0;
  wire s_csamul_cla32_fa29_6_xor1;
  wire s_csamul_cla32_fa29_6_and1;
  wire s_csamul_cla32_fa29_6_or0;
  wire s_csamul_cla32_and30_6;
  wire s_csamul_cla32_fa30_6_xor0;
  wire s_csamul_cla32_fa30_6_and0;
  wire s_csamul_cla32_fa30_6_xor1;
  wire s_csamul_cla32_fa30_6_and1;
  wire s_csamul_cla32_fa30_6_or0;
  wire s_csamul_cla32_nand31_6;
  wire s_csamul_cla32_ha31_6_xor0;
  wire s_csamul_cla32_ha31_6_and0;
  wire s_csamul_cla32_and0_7;
  wire s_csamul_cla32_fa0_7_xor0;
  wire s_csamul_cla32_fa0_7_and0;
  wire s_csamul_cla32_fa0_7_xor1;
  wire s_csamul_cla32_fa0_7_and1;
  wire s_csamul_cla32_fa0_7_or0;
  wire s_csamul_cla32_and1_7;
  wire s_csamul_cla32_fa1_7_xor0;
  wire s_csamul_cla32_fa1_7_and0;
  wire s_csamul_cla32_fa1_7_xor1;
  wire s_csamul_cla32_fa1_7_and1;
  wire s_csamul_cla32_fa1_7_or0;
  wire s_csamul_cla32_and2_7;
  wire s_csamul_cla32_fa2_7_xor0;
  wire s_csamul_cla32_fa2_7_and0;
  wire s_csamul_cla32_fa2_7_xor1;
  wire s_csamul_cla32_fa2_7_and1;
  wire s_csamul_cla32_fa2_7_or0;
  wire s_csamul_cla32_and3_7;
  wire s_csamul_cla32_fa3_7_xor0;
  wire s_csamul_cla32_fa3_7_and0;
  wire s_csamul_cla32_fa3_7_xor1;
  wire s_csamul_cla32_fa3_7_and1;
  wire s_csamul_cla32_fa3_7_or0;
  wire s_csamul_cla32_and4_7;
  wire s_csamul_cla32_fa4_7_xor0;
  wire s_csamul_cla32_fa4_7_and0;
  wire s_csamul_cla32_fa4_7_xor1;
  wire s_csamul_cla32_fa4_7_and1;
  wire s_csamul_cla32_fa4_7_or0;
  wire s_csamul_cla32_and5_7;
  wire s_csamul_cla32_fa5_7_xor0;
  wire s_csamul_cla32_fa5_7_and0;
  wire s_csamul_cla32_fa5_7_xor1;
  wire s_csamul_cla32_fa5_7_and1;
  wire s_csamul_cla32_fa5_7_or0;
  wire s_csamul_cla32_and6_7;
  wire s_csamul_cla32_fa6_7_xor0;
  wire s_csamul_cla32_fa6_7_and0;
  wire s_csamul_cla32_fa6_7_xor1;
  wire s_csamul_cla32_fa6_7_and1;
  wire s_csamul_cla32_fa6_7_or0;
  wire s_csamul_cla32_and7_7;
  wire s_csamul_cla32_fa7_7_xor0;
  wire s_csamul_cla32_fa7_7_and0;
  wire s_csamul_cla32_fa7_7_xor1;
  wire s_csamul_cla32_fa7_7_and1;
  wire s_csamul_cla32_fa7_7_or0;
  wire s_csamul_cla32_and8_7;
  wire s_csamul_cla32_fa8_7_xor0;
  wire s_csamul_cla32_fa8_7_and0;
  wire s_csamul_cla32_fa8_7_xor1;
  wire s_csamul_cla32_fa8_7_and1;
  wire s_csamul_cla32_fa8_7_or0;
  wire s_csamul_cla32_and9_7;
  wire s_csamul_cla32_fa9_7_xor0;
  wire s_csamul_cla32_fa9_7_and0;
  wire s_csamul_cla32_fa9_7_xor1;
  wire s_csamul_cla32_fa9_7_and1;
  wire s_csamul_cla32_fa9_7_or0;
  wire s_csamul_cla32_and10_7;
  wire s_csamul_cla32_fa10_7_xor0;
  wire s_csamul_cla32_fa10_7_and0;
  wire s_csamul_cla32_fa10_7_xor1;
  wire s_csamul_cla32_fa10_7_and1;
  wire s_csamul_cla32_fa10_7_or0;
  wire s_csamul_cla32_and11_7;
  wire s_csamul_cla32_fa11_7_xor0;
  wire s_csamul_cla32_fa11_7_and0;
  wire s_csamul_cla32_fa11_7_xor1;
  wire s_csamul_cla32_fa11_7_and1;
  wire s_csamul_cla32_fa11_7_or0;
  wire s_csamul_cla32_and12_7;
  wire s_csamul_cla32_fa12_7_xor0;
  wire s_csamul_cla32_fa12_7_and0;
  wire s_csamul_cla32_fa12_7_xor1;
  wire s_csamul_cla32_fa12_7_and1;
  wire s_csamul_cla32_fa12_7_or0;
  wire s_csamul_cla32_and13_7;
  wire s_csamul_cla32_fa13_7_xor0;
  wire s_csamul_cla32_fa13_7_and0;
  wire s_csamul_cla32_fa13_7_xor1;
  wire s_csamul_cla32_fa13_7_and1;
  wire s_csamul_cla32_fa13_7_or0;
  wire s_csamul_cla32_and14_7;
  wire s_csamul_cla32_fa14_7_xor0;
  wire s_csamul_cla32_fa14_7_and0;
  wire s_csamul_cla32_fa14_7_xor1;
  wire s_csamul_cla32_fa14_7_and1;
  wire s_csamul_cla32_fa14_7_or0;
  wire s_csamul_cla32_and15_7;
  wire s_csamul_cla32_fa15_7_xor0;
  wire s_csamul_cla32_fa15_7_and0;
  wire s_csamul_cla32_fa15_7_xor1;
  wire s_csamul_cla32_fa15_7_and1;
  wire s_csamul_cla32_fa15_7_or0;
  wire s_csamul_cla32_and16_7;
  wire s_csamul_cla32_fa16_7_xor0;
  wire s_csamul_cla32_fa16_7_and0;
  wire s_csamul_cla32_fa16_7_xor1;
  wire s_csamul_cla32_fa16_7_and1;
  wire s_csamul_cla32_fa16_7_or0;
  wire s_csamul_cla32_and17_7;
  wire s_csamul_cla32_fa17_7_xor0;
  wire s_csamul_cla32_fa17_7_and0;
  wire s_csamul_cla32_fa17_7_xor1;
  wire s_csamul_cla32_fa17_7_and1;
  wire s_csamul_cla32_fa17_7_or0;
  wire s_csamul_cla32_and18_7;
  wire s_csamul_cla32_fa18_7_xor0;
  wire s_csamul_cla32_fa18_7_and0;
  wire s_csamul_cla32_fa18_7_xor1;
  wire s_csamul_cla32_fa18_7_and1;
  wire s_csamul_cla32_fa18_7_or0;
  wire s_csamul_cla32_and19_7;
  wire s_csamul_cla32_fa19_7_xor0;
  wire s_csamul_cla32_fa19_7_and0;
  wire s_csamul_cla32_fa19_7_xor1;
  wire s_csamul_cla32_fa19_7_and1;
  wire s_csamul_cla32_fa19_7_or0;
  wire s_csamul_cla32_and20_7;
  wire s_csamul_cla32_fa20_7_xor0;
  wire s_csamul_cla32_fa20_7_and0;
  wire s_csamul_cla32_fa20_7_xor1;
  wire s_csamul_cla32_fa20_7_and1;
  wire s_csamul_cla32_fa20_7_or0;
  wire s_csamul_cla32_and21_7;
  wire s_csamul_cla32_fa21_7_xor0;
  wire s_csamul_cla32_fa21_7_and0;
  wire s_csamul_cla32_fa21_7_xor1;
  wire s_csamul_cla32_fa21_7_and1;
  wire s_csamul_cla32_fa21_7_or0;
  wire s_csamul_cla32_and22_7;
  wire s_csamul_cla32_fa22_7_xor0;
  wire s_csamul_cla32_fa22_7_and0;
  wire s_csamul_cla32_fa22_7_xor1;
  wire s_csamul_cla32_fa22_7_and1;
  wire s_csamul_cla32_fa22_7_or0;
  wire s_csamul_cla32_and23_7;
  wire s_csamul_cla32_fa23_7_xor0;
  wire s_csamul_cla32_fa23_7_and0;
  wire s_csamul_cla32_fa23_7_xor1;
  wire s_csamul_cla32_fa23_7_and1;
  wire s_csamul_cla32_fa23_7_or0;
  wire s_csamul_cla32_and24_7;
  wire s_csamul_cla32_fa24_7_xor0;
  wire s_csamul_cla32_fa24_7_and0;
  wire s_csamul_cla32_fa24_7_xor1;
  wire s_csamul_cla32_fa24_7_and1;
  wire s_csamul_cla32_fa24_7_or0;
  wire s_csamul_cla32_and25_7;
  wire s_csamul_cla32_fa25_7_xor0;
  wire s_csamul_cla32_fa25_7_and0;
  wire s_csamul_cla32_fa25_7_xor1;
  wire s_csamul_cla32_fa25_7_and1;
  wire s_csamul_cla32_fa25_7_or0;
  wire s_csamul_cla32_and26_7;
  wire s_csamul_cla32_fa26_7_xor0;
  wire s_csamul_cla32_fa26_7_and0;
  wire s_csamul_cla32_fa26_7_xor1;
  wire s_csamul_cla32_fa26_7_and1;
  wire s_csamul_cla32_fa26_7_or0;
  wire s_csamul_cla32_and27_7;
  wire s_csamul_cla32_fa27_7_xor0;
  wire s_csamul_cla32_fa27_7_and0;
  wire s_csamul_cla32_fa27_7_xor1;
  wire s_csamul_cla32_fa27_7_and1;
  wire s_csamul_cla32_fa27_7_or0;
  wire s_csamul_cla32_and28_7;
  wire s_csamul_cla32_fa28_7_xor0;
  wire s_csamul_cla32_fa28_7_and0;
  wire s_csamul_cla32_fa28_7_xor1;
  wire s_csamul_cla32_fa28_7_and1;
  wire s_csamul_cla32_fa28_7_or0;
  wire s_csamul_cla32_and29_7;
  wire s_csamul_cla32_fa29_7_xor0;
  wire s_csamul_cla32_fa29_7_and0;
  wire s_csamul_cla32_fa29_7_xor1;
  wire s_csamul_cla32_fa29_7_and1;
  wire s_csamul_cla32_fa29_7_or0;
  wire s_csamul_cla32_and30_7;
  wire s_csamul_cla32_fa30_7_xor0;
  wire s_csamul_cla32_fa30_7_and0;
  wire s_csamul_cla32_fa30_7_xor1;
  wire s_csamul_cla32_fa30_7_and1;
  wire s_csamul_cla32_fa30_7_or0;
  wire s_csamul_cla32_nand31_7;
  wire s_csamul_cla32_ha31_7_xor0;
  wire s_csamul_cla32_ha31_7_and0;
  wire s_csamul_cla32_and0_8;
  wire s_csamul_cla32_fa0_8_xor0;
  wire s_csamul_cla32_fa0_8_and0;
  wire s_csamul_cla32_fa0_8_xor1;
  wire s_csamul_cla32_fa0_8_and1;
  wire s_csamul_cla32_fa0_8_or0;
  wire s_csamul_cla32_and1_8;
  wire s_csamul_cla32_fa1_8_xor0;
  wire s_csamul_cla32_fa1_8_and0;
  wire s_csamul_cla32_fa1_8_xor1;
  wire s_csamul_cla32_fa1_8_and1;
  wire s_csamul_cla32_fa1_8_or0;
  wire s_csamul_cla32_and2_8;
  wire s_csamul_cla32_fa2_8_xor0;
  wire s_csamul_cla32_fa2_8_and0;
  wire s_csamul_cla32_fa2_8_xor1;
  wire s_csamul_cla32_fa2_8_and1;
  wire s_csamul_cla32_fa2_8_or0;
  wire s_csamul_cla32_and3_8;
  wire s_csamul_cla32_fa3_8_xor0;
  wire s_csamul_cla32_fa3_8_and0;
  wire s_csamul_cla32_fa3_8_xor1;
  wire s_csamul_cla32_fa3_8_and1;
  wire s_csamul_cla32_fa3_8_or0;
  wire s_csamul_cla32_and4_8;
  wire s_csamul_cla32_fa4_8_xor0;
  wire s_csamul_cla32_fa4_8_and0;
  wire s_csamul_cla32_fa4_8_xor1;
  wire s_csamul_cla32_fa4_8_and1;
  wire s_csamul_cla32_fa4_8_or0;
  wire s_csamul_cla32_and5_8;
  wire s_csamul_cla32_fa5_8_xor0;
  wire s_csamul_cla32_fa5_8_and0;
  wire s_csamul_cla32_fa5_8_xor1;
  wire s_csamul_cla32_fa5_8_and1;
  wire s_csamul_cla32_fa5_8_or0;
  wire s_csamul_cla32_and6_8;
  wire s_csamul_cla32_fa6_8_xor0;
  wire s_csamul_cla32_fa6_8_and0;
  wire s_csamul_cla32_fa6_8_xor1;
  wire s_csamul_cla32_fa6_8_and1;
  wire s_csamul_cla32_fa6_8_or0;
  wire s_csamul_cla32_and7_8;
  wire s_csamul_cla32_fa7_8_xor0;
  wire s_csamul_cla32_fa7_8_and0;
  wire s_csamul_cla32_fa7_8_xor1;
  wire s_csamul_cla32_fa7_8_and1;
  wire s_csamul_cla32_fa7_8_or0;
  wire s_csamul_cla32_and8_8;
  wire s_csamul_cla32_fa8_8_xor0;
  wire s_csamul_cla32_fa8_8_and0;
  wire s_csamul_cla32_fa8_8_xor1;
  wire s_csamul_cla32_fa8_8_and1;
  wire s_csamul_cla32_fa8_8_or0;
  wire s_csamul_cla32_and9_8;
  wire s_csamul_cla32_fa9_8_xor0;
  wire s_csamul_cla32_fa9_8_and0;
  wire s_csamul_cla32_fa9_8_xor1;
  wire s_csamul_cla32_fa9_8_and1;
  wire s_csamul_cla32_fa9_8_or0;
  wire s_csamul_cla32_and10_8;
  wire s_csamul_cla32_fa10_8_xor0;
  wire s_csamul_cla32_fa10_8_and0;
  wire s_csamul_cla32_fa10_8_xor1;
  wire s_csamul_cla32_fa10_8_and1;
  wire s_csamul_cla32_fa10_8_or0;
  wire s_csamul_cla32_and11_8;
  wire s_csamul_cla32_fa11_8_xor0;
  wire s_csamul_cla32_fa11_8_and0;
  wire s_csamul_cla32_fa11_8_xor1;
  wire s_csamul_cla32_fa11_8_and1;
  wire s_csamul_cla32_fa11_8_or0;
  wire s_csamul_cla32_and12_8;
  wire s_csamul_cla32_fa12_8_xor0;
  wire s_csamul_cla32_fa12_8_and0;
  wire s_csamul_cla32_fa12_8_xor1;
  wire s_csamul_cla32_fa12_8_and1;
  wire s_csamul_cla32_fa12_8_or0;
  wire s_csamul_cla32_and13_8;
  wire s_csamul_cla32_fa13_8_xor0;
  wire s_csamul_cla32_fa13_8_and0;
  wire s_csamul_cla32_fa13_8_xor1;
  wire s_csamul_cla32_fa13_8_and1;
  wire s_csamul_cla32_fa13_8_or0;
  wire s_csamul_cla32_and14_8;
  wire s_csamul_cla32_fa14_8_xor0;
  wire s_csamul_cla32_fa14_8_and0;
  wire s_csamul_cla32_fa14_8_xor1;
  wire s_csamul_cla32_fa14_8_and1;
  wire s_csamul_cla32_fa14_8_or0;
  wire s_csamul_cla32_and15_8;
  wire s_csamul_cla32_fa15_8_xor0;
  wire s_csamul_cla32_fa15_8_and0;
  wire s_csamul_cla32_fa15_8_xor1;
  wire s_csamul_cla32_fa15_8_and1;
  wire s_csamul_cla32_fa15_8_or0;
  wire s_csamul_cla32_and16_8;
  wire s_csamul_cla32_fa16_8_xor0;
  wire s_csamul_cla32_fa16_8_and0;
  wire s_csamul_cla32_fa16_8_xor1;
  wire s_csamul_cla32_fa16_8_and1;
  wire s_csamul_cla32_fa16_8_or0;
  wire s_csamul_cla32_and17_8;
  wire s_csamul_cla32_fa17_8_xor0;
  wire s_csamul_cla32_fa17_8_and0;
  wire s_csamul_cla32_fa17_8_xor1;
  wire s_csamul_cla32_fa17_8_and1;
  wire s_csamul_cla32_fa17_8_or0;
  wire s_csamul_cla32_and18_8;
  wire s_csamul_cla32_fa18_8_xor0;
  wire s_csamul_cla32_fa18_8_and0;
  wire s_csamul_cla32_fa18_8_xor1;
  wire s_csamul_cla32_fa18_8_and1;
  wire s_csamul_cla32_fa18_8_or0;
  wire s_csamul_cla32_and19_8;
  wire s_csamul_cla32_fa19_8_xor0;
  wire s_csamul_cla32_fa19_8_and0;
  wire s_csamul_cla32_fa19_8_xor1;
  wire s_csamul_cla32_fa19_8_and1;
  wire s_csamul_cla32_fa19_8_or0;
  wire s_csamul_cla32_and20_8;
  wire s_csamul_cla32_fa20_8_xor0;
  wire s_csamul_cla32_fa20_8_and0;
  wire s_csamul_cla32_fa20_8_xor1;
  wire s_csamul_cla32_fa20_8_and1;
  wire s_csamul_cla32_fa20_8_or0;
  wire s_csamul_cla32_and21_8;
  wire s_csamul_cla32_fa21_8_xor0;
  wire s_csamul_cla32_fa21_8_and0;
  wire s_csamul_cla32_fa21_8_xor1;
  wire s_csamul_cla32_fa21_8_and1;
  wire s_csamul_cla32_fa21_8_or0;
  wire s_csamul_cla32_and22_8;
  wire s_csamul_cla32_fa22_8_xor0;
  wire s_csamul_cla32_fa22_8_and0;
  wire s_csamul_cla32_fa22_8_xor1;
  wire s_csamul_cla32_fa22_8_and1;
  wire s_csamul_cla32_fa22_8_or0;
  wire s_csamul_cla32_and23_8;
  wire s_csamul_cla32_fa23_8_xor0;
  wire s_csamul_cla32_fa23_8_and0;
  wire s_csamul_cla32_fa23_8_xor1;
  wire s_csamul_cla32_fa23_8_and1;
  wire s_csamul_cla32_fa23_8_or0;
  wire s_csamul_cla32_and24_8;
  wire s_csamul_cla32_fa24_8_xor0;
  wire s_csamul_cla32_fa24_8_and0;
  wire s_csamul_cla32_fa24_8_xor1;
  wire s_csamul_cla32_fa24_8_and1;
  wire s_csamul_cla32_fa24_8_or0;
  wire s_csamul_cla32_and25_8;
  wire s_csamul_cla32_fa25_8_xor0;
  wire s_csamul_cla32_fa25_8_and0;
  wire s_csamul_cla32_fa25_8_xor1;
  wire s_csamul_cla32_fa25_8_and1;
  wire s_csamul_cla32_fa25_8_or0;
  wire s_csamul_cla32_and26_8;
  wire s_csamul_cla32_fa26_8_xor0;
  wire s_csamul_cla32_fa26_8_and0;
  wire s_csamul_cla32_fa26_8_xor1;
  wire s_csamul_cla32_fa26_8_and1;
  wire s_csamul_cla32_fa26_8_or0;
  wire s_csamul_cla32_and27_8;
  wire s_csamul_cla32_fa27_8_xor0;
  wire s_csamul_cla32_fa27_8_and0;
  wire s_csamul_cla32_fa27_8_xor1;
  wire s_csamul_cla32_fa27_8_and1;
  wire s_csamul_cla32_fa27_8_or0;
  wire s_csamul_cla32_and28_8;
  wire s_csamul_cla32_fa28_8_xor0;
  wire s_csamul_cla32_fa28_8_and0;
  wire s_csamul_cla32_fa28_8_xor1;
  wire s_csamul_cla32_fa28_8_and1;
  wire s_csamul_cla32_fa28_8_or0;
  wire s_csamul_cla32_and29_8;
  wire s_csamul_cla32_fa29_8_xor0;
  wire s_csamul_cla32_fa29_8_and0;
  wire s_csamul_cla32_fa29_8_xor1;
  wire s_csamul_cla32_fa29_8_and1;
  wire s_csamul_cla32_fa29_8_or0;
  wire s_csamul_cla32_and30_8;
  wire s_csamul_cla32_fa30_8_xor0;
  wire s_csamul_cla32_fa30_8_and0;
  wire s_csamul_cla32_fa30_8_xor1;
  wire s_csamul_cla32_fa30_8_and1;
  wire s_csamul_cla32_fa30_8_or0;
  wire s_csamul_cla32_nand31_8;
  wire s_csamul_cla32_ha31_8_xor0;
  wire s_csamul_cla32_ha31_8_and0;
  wire s_csamul_cla32_and0_9;
  wire s_csamul_cla32_fa0_9_xor0;
  wire s_csamul_cla32_fa0_9_and0;
  wire s_csamul_cla32_fa0_9_xor1;
  wire s_csamul_cla32_fa0_9_and1;
  wire s_csamul_cla32_fa0_9_or0;
  wire s_csamul_cla32_and1_9;
  wire s_csamul_cla32_fa1_9_xor0;
  wire s_csamul_cla32_fa1_9_and0;
  wire s_csamul_cla32_fa1_9_xor1;
  wire s_csamul_cla32_fa1_9_and1;
  wire s_csamul_cla32_fa1_9_or0;
  wire s_csamul_cla32_and2_9;
  wire s_csamul_cla32_fa2_9_xor0;
  wire s_csamul_cla32_fa2_9_and0;
  wire s_csamul_cla32_fa2_9_xor1;
  wire s_csamul_cla32_fa2_9_and1;
  wire s_csamul_cla32_fa2_9_or0;
  wire s_csamul_cla32_and3_9;
  wire s_csamul_cla32_fa3_9_xor0;
  wire s_csamul_cla32_fa3_9_and0;
  wire s_csamul_cla32_fa3_9_xor1;
  wire s_csamul_cla32_fa3_9_and1;
  wire s_csamul_cla32_fa3_9_or0;
  wire s_csamul_cla32_and4_9;
  wire s_csamul_cla32_fa4_9_xor0;
  wire s_csamul_cla32_fa4_9_and0;
  wire s_csamul_cla32_fa4_9_xor1;
  wire s_csamul_cla32_fa4_9_and1;
  wire s_csamul_cla32_fa4_9_or0;
  wire s_csamul_cla32_and5_9;
  wire s_csamul_cla32_fa5_9_xor0;
  wire s_csamul_cla32_fa5_9_and0;
  wire s_csamul_cla32_fa5_9_xor1;
  wire s_csamul_cla32_fa5_9_and1;
  wire s_csamul_cla32_fa5_9_or0;
  wire s_csamul_cla32_and6_9;
  wire s_csamul_cla32_fa6_9_xor0;
  wire s_csamul_cla32_fa6_9_and0;
  wire s_csamul_cla32_fa6_9_xor1;
  wire s_csamul_cla32_fa6_9_and1;
  wire s_csamul_cla32_fa6_9_or0;
  wire s_csamul_cla32_and7_9;
  wire s_csamul_cla32_fa7_9_xor0;
  wire s_csamul_cla32_fa7_9_and0;
  wire s_csamul_cla32_fa7_9_xor1;
  wire s_csamul_cla32_fa7_9_and1;
  wire s_csamul_cla32_fa7_9_or0;
  wire s_csamul_cla32_and8_9;
  wire s_csamul_cla32_fa8_9_xor0;
  wire s_csamul_cla32_fa8_9_and0;
  wire s_csamul_cla32_fa8_9_xor1;
  wire s_csamul_cla32_fa8_9_and1;
  wire s_csamul_cla32_fa8_9_or0;
  wire s_csamul_cla32_and9_9;
  wire s_csamul_cla32_fa9_9_xor0;
  wire s_csamul_cla32_fa9_9_and0;
  wire s_csamul_cla32_fa9_9_xor1;
  wire s_csamul_cla32_fa9_9_and1;
  wire s_csamul_cla32_fa9_9_or0;
  wire s_csamul_cla32_and10_9;
  wire s_csamul_cla32_fa10_9_xor0;
  wire s_csamul_cla32_fa10_9_and0;
  wire s_csamul_cla32_fa10_9_xor1;
  wire s_csamul_cla32_fa10_9_and1;
  wire s_csamul_cla32_fa10_9_or0;
  wire s_csamul_cla32_and11_9;
  wire s_csamul_cla32_fa11_9_xor0;
  wire s_csamul_cla32_fa11_9_and0;
  wire s_csamul_cla32_fa11_9_xor1;
  wire s_csamul_cla32_fa11_9_and1;
  wire s_csamul_cla32_fa11_9_or0;
  wire s_csamul_cla32_and12_9;
  wire s_csamul_cla32_fa12_9_xor0;
  wire s_csamul_cla32_fa12_9_and0;
  wire s_csamul_cla32_fa12_9_xor1;
  wire s_csamul_cla32_fa12_9_and1;
  wire s_csamul_cla32_fa12_9_or0;
  wire s_csamul_cla32_and13_9;
  wire s_csamul_cla32_fa13_9_xor0;
  wire s_csamul_cla32_fa13_9_and0;
  wire s_csamul_cla32_fa13_9_xor1;
  wire s_csamul_cla32_fa13_9_and1;
  wire s_csamul_cla32_fa13_9_or0;
  wire s_csamul_cla32_and14_9;
  wire s_csamul_cla32_fa14_9_xor0;
  wire s_csamul_cla32_fa14_9_and0;
  wire s_csamul_cla32_fa14_9_xor1;
  wire s_csamul_cla32_fa14_9_and1;
  wire s_csamul_cla32_fa14_9_or0;
  wire s_csamul_cla32_and15_9;
  wire s_csamul_cla32_fa15_9_xor0;
  wire s_csamul_cla32_fa15_9_and0;
  wire s_csamul_cla32_fa15_9_xor1;
  wire s_csamul_cla32_fa15_9_and1;
  wire s_csamul_cla32_fa15_9_or0;
  wire s_csamul_cla32_and16_9;
  wire s_csamul_cla32_fa16_9_xor0;
  wire s_csamul_cla32_fa16_9_and0;
  wire s_csamul_cla32_fa16_9_xor1;
  wire s_csamul_cla32_fa16_9_and1;
  wire s_csamul_cla32_fa16_9_or0;
  wire s_csamul_cla32_and17_9;
  wire s_csamul_cla32_fa17_9_xor0;
  wire s_csamul_cla32_fa17_9_and0;
  wire s_csamul_cla32_fa17_9_xor1;
  wire s_csamul_cla32_fa17_9_and1;
  wire s_csamul_cla32_fa17_9_or0;
  wire s_csamul_cla32_and18_9;
  wire s_csamul_cla32_fa18_9_xor0;
  wire s_csamul_cla32_fa18_9_and0;
  wire s_csamul_cla32_fa18_9_xor1;
  wire s_csamul_cla32_fa18_9_and1;
  wire s_csamul_cla32_fa18_9_or0;
  wire s_csamul_cla32_and19_9;
  wire s_csamul_cla32_fa19_9_xor0;
  wire s_csamul_cla32_fa19_9_and0;
  wire s_csamul_cla32_fa19_9_xor1;
  wire s_csamul_cla32_fa19_9_and1;
  wire s_csamul_cla32_fa19_9_or0;
  wire s_csamul_cla32_and20_9;
  wire s_csamul_cla32_fa20_9_xor0;
  wire s_csamul_cla32_fa20_9_and0;
  wire s_csamul_cla32_fa20_9_xor1;
  wire s_csamul_cla32_fa20_9_and1;
  wire s_csamul_cla32_fa20_9_or0;
  wire s_csamul_cla32_and21_9;
  wire s_csamul_cla32_fa21_9_xor0;
  wire s_csamul_cla32_fa21_9_and0;
  wire s_csamul_cla32_fa21_9_xor1;
  wire s_csamul_cla32_fa21_9_and1;
  wire s_csamul_cla32_fa21_9_or0;
  wire s_csamul_cla32_and22_9;
  wire s_csamul_cla32_fa22_9_xor0;
  wire s_csamul_cla32_fa22_9_and0;
  wire s_csamul_cla32_fa22_9_xor1;
  wire s_csamul_cla32_fa22_9_and1;
  wire s_csamul_cla32_fa22_9_or0;
  wire s_csamul_cla32_and23_9;
  wire s_csamul_cla32_fa23_9_xor0;
  wire s_csamul_cla32_fa23_9_and0;
  wire s_csamul_cla32_fa23_9_xor1;
  wire s_csamul_cla32_fa23_9_and1;
  wire s_csamul_cla32_fa23_9_or0;
  wire s_csamul_cla32_and24_9;
  wire s_csamul_cla32_fa24_9_xor0;
  wire s_csamul_cla32_fa24_9_and0;
  wire s_csamul_cla32_fa24_9_xor1;
  wire s_csamul_cla32_fa24_9_and1;
  wire s_csamul_cla32_fa24_9_or0;
  wire s_csamul_cla32_and25_9;
  wire s_csamul_cla32_fa25_9_xor0;
  wire s_csamul_cla32_fa25_9_and0;
  wire s_csamul_cla32_fa25_9_xor1;
  wire s_csamul_cla32_fa25_9_and1;
  wire s_csamul_cla32_fa25_9_or0;
  wire s_csamul_cla32_and26_9;
  wire s_csamul_cla32_fa26_9_xor0;
  wire s_csamul_cla32_fa26_9_and0;
  wire s_csamul_cla32_fa26_9_xor1;
  wire s_csamul_cla32_fa26_9_and1;
  wire s_csamul_cla32_fa26_9_or0;
  wire s_csamul_cla32_and27_9;
  wire s_csamul_cla32_fa27_9_xor0;
  wire s_csamul_cla32_fa27_9_and0;
  wire s_csamul_cla32_fa27_9_xor1;
  wire s_csamul_cla32_fa27_9_and1;
  wire s_csamul_cla32_fa27_9_or0;
  wire s_csamul_cla32_and28_9;
  wire s_csamul_cla32_fa28_9_xor0;
  wire s_csamul_cla32_fa28_9_and0;
  wire s_csamul_cla32_fa28_9_xor1;
  wire s_csamul_cla32_fa28_9_and1;
  wire s_csamul_cla32_fa28_9_or0;
  wire s_csamul_cla32_and29_9;
  wire s_csamul_cla32_fa29_9_xor0;
  wire s_csamul_cla32_fa29_9_and0;
  wire s_csamul_cla32_fa29_9_xor1;
  wire s_csamul_cla32_fa29_9_and1;
  wire s_csamul_cla32_fa29_9_or0;
  wire s_csamul_cla32_and30_9;
  wire s_csamul_cla32_fa30_9_xor0;
  wire s_csamul_cla32_fa30_9_and0;
  wire s_csamul_cla32_fa30_9_xor1;
  wire s_csamul_cla32_fa30_9_and1;
  wire s_csamul_cla32_fa30_9_or0;
  wire s_csamul_cla32_nand31_9;
  wire s_csamul_cla32_ha31_9_xor0;
  wire s_csamul_cla32_ha31_9_and0;
  wire s_csamul_cla32_and0_10;
  wire s_csamul_cla32_fa0_10_xor0;
  wire s_csamul_cla32_fa0_10_and0;
  wire s_csamul_cla32_fa0_10_xor1;
  wire s_csamul_cla32_fa0_10_and1;
  wire s_csamul_cla32_fa0_10_or0;
  wire s_csamul_cla32_and1_10;
  wire s_csamul_cla32_fa1_10_xor0;
  wire s_csamul_cla32_fa1_10_and0;
  wire s_csamul_cla32_fa1_10_xor1;
  wire s_csamul_cla32_fa1_10_and1;
  wire s_csamul_cla32_fa1_10_or0;
  wire s_csamul_cla32_and2_10;
  wire s_csamul_cla32_fa2_10_xor0;
  wire s_csamul_cla32_fa2_10_and0;
  wire s_csamul_cla32_fa2_10_xor1;
  wire s_csamul_cla32_fa2_10_and1;
  wire s_csamul_cla32_fa2_10_or0;
  wire s_csamul_cla32_and3_10;
  wire s_csamul_cla32_fa3_10_xor0;
  wire s_csamul_cla32_fa3_10_and0;
  wire s_csamul_cla32_fa3_10_xor1;
  wire s_csamul_cla32_fa3_10_and1;
  wire s_csamul_cla32_fa3_10_or0;
  wire s_csamul_cla32_and4_10;
  wire s_csamul_cla32_fa4_10_xor0;
  wire s_csamul_cla32_fa4_10_and0;
  wire s_csamul_cla32_fa4_10_xor1;
  wire s_csamul_cla32_fa4_10_and1;
  wire s_csamul_cla32_fa4_10_or0;
  wire s_csamul_cla32_and5_10;
  wire s_csamul_cla32_fa5_10_xor0;
  wire s_csamul_cla32_fa5_10_and0;
  wire s_csamul_cla32_fa5_10_xor1;
  wire s_csamul_cla32_fa5_10_and1;
  wire s_csamul_cla32_fa5_10_or0;
  wire s_csamul_cla32_and6_10;
  wire s_csamul_cla32_fa6_10_xor0;
  wire s_csamul_cla32_fa6_10_and0;
  wire s_csamul_cla32_fa6_10_xor1;
  wire s_csamul_cla32_fa6_10_and1;
  wire s_csamul_cla32_fa6_10_or0;
  wire s_csamul_cla32_and7_10;
  wire s_csamul_cla32_fa7_10_xor0;
  wire s_csamul_cla32_fa7_10_and0;
  wire s_csamul_cla32_fa7_10_xor1;
  wire s_csamul_cla32_fa7_10_and1;
  wire s_csamul_cla32_fa7_10_or0;
  wire s_csamul_cla32_and8_10;
  wire s_csamul_cla32_fa8_10_xor0;
  wire s_csamul_cla32_fa8_10_and0;
  wire s_csamul_cla32_fa8_10_xor1;
  wire s_csamul_cla32_fa8_10_and1;
  wire s_csamul_cla32_fa8_10_or0;
  wire s_csamul_cla32_and9_10;
  wire s_csamul_cla32_fa9_10_xor0;
  wire s_csamul_cla32_fa9_10_and0;
  wire s_csamul_cla32_fa9_10_xor1;
  wire s_csamul_cla32_fa9_10_and1;
  wire s_csamul_cla32_fa9_10_or0;
  wire s_csamul_cla32_and10_10;
  wire s_csamul_cla32_fa10_10_xor0;
  wire s_csamul_cla32_fa10_10_and0;
  wire s_csamul_cla32_fa10_10_xor1;
  wire s_csamul_cla32_fa10_10_and1;
  wire s_csamul_cla32_fa10_10_or0;
  wire s_csamul_cla32_and11_10;
  wire s_csamul_cla32_fa11_10_xor0;
  wire s_csamul_cla32_fa11_10_and0;
  wire s_csamul_cla32_fa11_10_xor1;
  wire s_csamul_cla32_fa11_10_and1;
  wire s_csamul_cla32_fa11_10_or0;
  wire s_csamul_cla32_and12_10;
  wire s_csamul_cla32_fa12_10_xor0;
  wire s_csamul_cla32_fa12_10_and0;
  wire s_csamul_cla32_fa12_10_xor1;
  wire s_csamul_cla32_fa12_10_and1;
  wire s_csamul_cla32_fa12_10_or0;
  wire s_csamul_cla32_and13_10;
  wire s_csamul_cla32_fa13_10_xor0;
  wire s_csamul_cla32_fa13_10_and0;
  wire s_csamul_cla32_fa13_10_xor1;
  wire s_csamul_cla32_fa13_10_and1;
  wire s_csamul_cla32_fa13_10_or0;
  wire s_csamul_cla32_and14_10;
  wire s_csamul_cla32_fa14_10_xor0;
  wire s_csamul_cla32_fa14_10_and0;
  wire s_csamul_cla32_fa14_10_xor1;
  wire s_csamul_cla32_fa14_10_and1;
  wire s_csamul_cla32_fa14_10_or0;
  wire s_csamul_cla32_and15_10;
  wire s_csamul_cla32_fa15_10_xor0;
  wire s_csamul_cla32_fa15_10_and0;
  wire s_csamul_cla32_fa15_10_xor1;
  wire s_csamul_cla32_fa15_10_and1;
  wire s_csamul_cla32_fa15_10_or0;
  wire s_csamul_cla32_and16_10;
  wire s_csamul_cla32_fa16_10_xor0;
  wire s_csamul_cla32_fa16_10_and0;
  wire s_csamul_cla32_fa16_10_xor1;
  wire s_csamul_cla32_fa16_10_and1;
  wire s_csamul_cla32_fa16_10_or0;
  wire s_csamul_cla32_and17_10;
  wire s_csamul_cla32_fa17_10_xor0;
  wire s_csamul_cla32_fa17_10_and0;
  wire s_csamul_cla32_fa17_10_xor1;
  wire s_csamul_cla32_fa17_10_and1;
  wire s_csamul_cla32_fa17_10_or0;
  wire s_csamul_cla32_and18_10;
  wire s_csamul_cla32_fa18_10_xor0;
  wire s_csamul_cla32_fa18_10_and0;
  wire s_csamul_cla32_fa18_10_xor1;
  wire s_csamul_cla32_fa18_10_and1;
  wire s_csamul_cla32_fa18_10_or0;
  wire s_csamul_cla32_and19_10;
  wire s_csamul_cla32_fa19_10_xor0;
  wire s_csamul_cla32_fa19_10_and0;
  wire s_csamul_cla32_fa19_10_xor1;
  wire s_csamul_cla32_fa19_10_and1;
  wire s_csamul_cla32_fa19_10_or0;
  wire s_csamul_cla32_and20_10;
  wire s_csamul_cla32_fa20_10_xor0;
  wire s_csamul_cla32_fa20_10_and0;
  wire s_csamul_cla32_fa20_10_xor1;
  wire s_csamul_cla32_fa20_10_and1;
  wire s_csamul_cla32_fa20_10_or0;
  wire s_csamul_cla32_and21_10;
  wire s_csamul_cla32_fa21_10_xor0;
  wire s_csamul_cla32_fa21_10_and0;
  wire s_csamul_cla32_fa21_10_xor1;
  wire s_csamul_cla32_fa21_10_and1;
  wire s_csamul_cla32_fa21_10_or0;
  wire s_csamul_cla32_and22_10;
  wire s_csamul_cla32_fa22_10_xor0;
  wire s_csamul_cla32_fa22_10_and0;
  wire s_csamul_cla32_fa22_10_xor1;
  wire s_csamul_cla32_fa22_10_and1;
  wire s_csamul_cla32_fa22_10_or0;
  wire s_csamul_cla32_and23_10;
  wire s_csamul_cla32_fa23_10_xor0;
  wire s_csamul_cla32_fa23_10_and0;
  wire s_csamul_cla32_fa23_10_xor1;
  wire s_csamul_cla32_fa23_10_and1;
  wire s_csamul_cla32_fa23_10_or0;
  wire s_csamul_cla32_and24_10;
  wire s_csamul_cla32_fa24_10_xor0;
  wire s_csamul_cla32_fa24_10_and0;
  wire s_csamul_cla32_fa24_10_xor1;
  wire s_csamul_cla32_fa24_10_and1;
  wire s_csamul_cla32_fa24_10_or0;
  wire s_csamul_cla32_and25_10;
  wire s_csamul_cla32_fa25_10_xor0;
  wire s_csamul_cla32_fa25_10_and0;
  wire s_csamul_cla32_fa25_10_xor1;
  wire s_csamul_cla32_fa25_10_and1;
  wire s_csamul_cla32_fa25_10_or0;
  wire s_csamul_cla32_and26_10;
  wire s_csamul_cla32_fa26_10_xor0;
  wire s_csamul_cla32_fa26_10_and0;
  wire s_csamul_cla32_fa26_10_xor1;
  wire s_csamul_cla32_fa26_10_and1;
  wire s_csamul_cla32_fa26_10_or0;
  wire s_csamul_cla32_and27_10;
  wire s_csamul_cla32_fa27_10_xor0;
  wire s_csamul_cla32_fa27_10_and0;
  wire s_csamul_cla32_fa27_10_xor1;
  wire s_csamul_cla32_fa27_10_and1;
  wire s_csamul_cla32_fa27_10_or0;
  wire s_csamul_cla32_and28_10;
  wire s_csamul_cla32_fa28_10_xor0;
  wire s_csamul_cla32_fa28_10_and0;
  wire s_csamul_cla32_fa28_10_xor1;
  wire s_csamul_cla32_fa28_10_and1;
  wire s_csamul_cla32_fa28_10_or0;
  wire s_csamul_cla32_and29_10;
  wire s_csamul_cla32_fa29_10_xor0;
  wire s_csamul_cla32_fa29_10_and0;
  wire s_csamul_cla32_fa29_10_xor1;
  wire s_csamul_cla32_fa29_10_and1;
  wire s_csamul_cla32_fa29_10_or0;
  wire s_csamul_cla32_and30_10;
  wire s_csamul_cla32_fa30_10_xor0;
  wire s_csamul_cla32_fa30_10_and0;
  wire s_csamul_cla32_fa30_10_xor1;
  wire s_csamul_cla32_fa30_10_and1;
  wire s_csamul_cla32_fa30_10_or0;
  wire s_csamul_cla32_nand31_10;
  wire s_csamul_cla32_ha31_10_xor0;
  wire s_csamul_cla32_ha31_10_and0;
  wire s_csamul_cla32_and0_11;
  wire s_csamul_cla32_fa0_11_xor0;
  wire s_csamul_cla32_fa0_11_and0;
  wire s_csamul_cla32_fa0_11_xor1;
  wire s_csamul_cla32_fa0_11_and1;
  wire s_csamul_cla32_fa0_11_or0;
  wire s_csamul_cla32_and1_11;
  wire s_csamul_cla32_fa1_11_xor0;
  wire s_csamul_cla32_fa1_11_and0;
  wire s_csamul_cla32_fa1_11_xor1;
  wire s_csamul_cla32_fa1_11_and1;
  wire s_csamul_cla32_fa1_11_or0;
  wire s_csamul_cla32_and2_11;
  wire s_csamul_cla32_fa2_11_xor0;
  wire s_csamul_cla32_fa2_11_and0;
  wire s_csamul_cla32_fa2_11_xor1;
  wire s_csamul_cla32_fa2_11_and1;
  wire s_csamul_cla32_fa2_11_or0;
  wire s_csamul_cla32_and3_11;
  wire s_csamul_cla32_fa3_11_xor0;
  wire s_csamul_cla32_fa3_11_and0;
  wire s_csamul_cla32_fa3_11_xor1;
  wire s_csamul_cla32_fa3_11_and1;
  wire s_csamul_cla32_fa3_11_or0;
  wire s_csamul_cla32_and4_11;
  wire s_csamul_cla32_fa4_11_xor0;
  wire s_csamul_cla32_fa4_11_and0;
  wire s_csamul_cla32_fa4_11_xor1;
  wire s_csamul_cla32_fa4_11_and1;
  wire s_csamul_cla32_fa4_11_or0;
  wire s_csamul_cla32_and5_11;
  wire s_csamul_cla32_fa5_11_xor0;
  wire s_csamul_cla32_fa5_11_and0;
  wire s_csamul_cla32_fa5_11_xor1;
  wire s_csamul_cla32_fa5_11_and1;
  wire s_csamul_cla32_fa5_11_or0;
  wire s_csamul_cla32_and6_11;
  wire s_csamul_cla32_fa6_11_xor0;
  wire s_csamul_cla32_fa6_11_and0;
  wire s_csamul_cla32_fa6_11_xor1;
  wire s_csamul_cla32_fa6_11_and1;
  wire s_csamul_cla32_fa6_11_or0;
  wire s_csamul_cla32_and7_11;
  wire s_csamul_cla32_fa7_11_xor0;
  wire s_csamul_cla32_fa7_11_and0;
  wire s_csamul_cla32_fa7_11_xor1;
  wire s_csamul_cla32_fa7_11_and1;
  wire s_csamul_cla32_fa7_11_or0;
  wire s_csamul_cla32_and8_11;
  wire s_csamul_cla32_fa8_11_xor0;
  wire s_csamul_cla32_fa8_11_and0;
  wire s_csamul_cla32_fa8_11_xor1;
  wire s_csamul_cla32_fa8_11_and1;
  wire s_csamul_cla32_fa8_11_or0;
  wire s_csamul_cla32_and9_11;
  wire s_csamul_cla32_fa9_11_xor0;
  wire s_csamul_cla32_fa9_11_and0;
  wire s_csamul_cla32_fa9_11_xor1;
  wire s_csamul_cla32_fa9_11_and1;
  wire s_csamul_cla32_fa9_11_or0;
  wire s_csamul_cla32_and10_11;
  wire s_csamul_cla32_fa10_11_xor0;
  wire s_csamul_cla32_fa10_11_and0;
  wire s_csamul_cla32_fa10_11_xor1;
  wire s_csamul_cla32_fa10_11_and1;
  wire s_csamul_cla32_fa10_11_or0;
  wire s_csamul_cla32_and11_11;
  wire s_csamul_cla32_fa11_11_xor0;
  wire s_csamul_cla32_fa11_11_and0;
  wire s_csamul_cla32_fa11_11_xor1;
  wire s_csamul_cla32_fa11_11_and1;
  wire s_csamul_cla32_fa11_11_or0;
  wire s_csamul_cla32_and12_11;
  wire s_csamul_cla32_fa12_11_xor0;
  wire s_csamul_cla32_fa12_11_and0;
  wire s_csamul_cla32_fa12_11_xor1;
  wire s_csamul_cla32_fa12_11_and1;
  wire s_csamul_cla32_fa12_11_or0;
  wire s_csamul_cla32_and13_11;
  wire s_csamul_cla32_fa13_11_xor0;
  wire s_csamul_cla32_fa13_11_and0;
  wire s_csamul_cla32_fa13_11_xor1;
  wire s_csamul_cla32_fa13_11_and1;
  wire s_csamul_cla32_fa13_11_or0;
  wire s_csamul_cla32_and14_11;
  wire s_csamul_cla32_fa14_11_xor0;
  wire s_csamul_cla32_fa14_11_and0;
  wire s_csamul_cla32_fa14_11_xor1;
  wire s_csamul_cla32_fa14_11_and1;
  wire s_csamul_cla32_fa14_11_or0;
  wire s_csamul_cla32_and15_11;
  wire s_csamul_cla32_fa15_11_xor0;
  wire s_csamul_cla32_fa15_11_and0;
  wire s_csamul_cla32_fa15_11_xor1;
  wire s_csamul_cla32_fa15_11_and1;
  wire s_csamul_cla32_fa15_11_or0;
  wire s_csamul_cla32_and16_11;
  wire s_csamul_cla32_fa16_11_xor0;
  wire s_csamul_cla32_fa16_11_and0;
  wire s_csamul_cla32_fa16_11_xor1;
  wire s_csamul_cla32_fa16_11_and1;
  wire s_csamul_cla32_fa16_11_or0;
  wire s_csamul_cla32_and17_11;
  wire s_csamul_cla32_fa17_11_xor0;
  wire s_csamul_cla32_fa17_11_and0;
  wire s_csamul_cla32_fa17_11_xor1;
  wire s_csamul_cla32_fa17_11_and1;
  wire s_csamul_cla32_fa17_11_or0;
  wire s_csamul_cla32_and18_11;
  wire s_csamul_cla32_fa18_11_xor0;
  wire s_csamul_cla32_fa18_11_and0;
  wire s_csamul_cla32_fa18_11_xor1;
  wire s_csamul_cla32_fa18_11_and1;
  wire s_csamul_cla32_fa18_11_or0;
  wire s_csamul_cla32_and19_11;
  wire s_csamul_cla32_fa19_11_xor0;
  wire s_csamul_cla32_fa19_11_and0;
  wire s_csamul_cla32_fa19_11_xor1;
  wire s_csamul_cla32_fa19_11_and1;
  wire s_csamul_cla32_fa19_11_or0;
  wire s_csamul_cla32_and20_11;
  wire s_csamul_cla32_fa20_11_xor0;
  wire s_csamul_cla32_fa20_11_and0;
  wire s_csamul_cla32_fa20_11_xor1;
  wire s_csamul_cla32_fa20_11_and1;
  wire s_csamul_cla32_fa20_11_or0;
  wire s_csamul_cla32_and21_11;
  wire s_csamul_cla32_fa21_11_xor0;
  wire s_csamul_cla32_fa21_11_and0;
  wire s_csamul_cla32_fa21_11_xor1;
  wire s_csamul_cla32_fa21_11_and1;
  wire s_csamul_cla32_fa21_11_or0;
  wire s_csamul_cla32_and22_11;
  wire s_csamul_cla32_fa22_11_xor0;
  wire s_csamul_cla32_fa22_11_and0;
  wire s_csamul_cla32_fa22_11_xor1;
  wire s_csamul_cla32_fa22_11_and1;
  wire s_csamul_cla32_fa22_11_or0;
  wire s_csamul_cla32_and23_11;
  wire s_csamul_cla32_fa23_11_xor0;
  wire s_csamul_cla32_fa23_11_and0;
  wire s_csamul_cla32_fa23_11_xor1;
  wire s_csamul_cla32_fa23_11_and1;
  wire s_csamul_cla32_fa23_11_or0;
  wire s_csamul_cla32_and24_11;
  wire s_csamul_cla32_fa24_11_xor0;
  wire s_csamul_cla32_fa24_11_and0;
  wire s_csamul_cla32_fa24_11_xor1;
  wire s_csamul_cla32_fa24_11_and1;
  wire s_csamul_cla32_fa24_11_or0;
  wire s_csamul_cla32_and25_11;
  wire s_csamul_cla32_fa25_11_xor0;
  wire s_csamul_cla32_fa25_11_and0;
  wire s_csamul_cla32_fa25_11_xor1;
  wire s_csamul_cla32_fa25_11_and1;
  wire s_csamul_cla32_fa25_11_or0;
  wire s_csamul_cla32_and26_11;
  wire s_csamul_cla32_fa26_11_xor0;
  wire s_csamul_cla32_fa26_11_and0;
  wire s_csamul_cla32_fa26_11_xor1;
  wire s_csamul_cla32_fa26_11_and1;
  wire s_csamul_cla32_fa26_11_or0;
  wire s_csamul_cla32_and27_11;
  wire s_csamul_cla32_fa27_11_xor0;
  wire s_csamul_cla32_fa27_11_and0;
  wire s_csamul_cla32_fa27_11_xor1;
  wire s_csamul_cla32_fa27_11_and1;
  wire s_csamul_cla32_fa27_11_or0;
  wire s_csamul_cla32_and28_11;
  wire s_csamul_cla32_fa28_11_xor0;
  wire s_csamul_cla32_fa28_11_and0;
  wire s_csamul_cla32_fa28_11_xor1;
  wire s_csamul_cla32_fa28_11_and1;
  wire s_csamul_cla32_fa28_11_or0;
  wire s_csamul_cla32_and29_11;
  wire s_csamul_cla32_fa29_11_xor0;
  wire s_csamul_cla32_fa29_11_and0;
  wire s_csamul_cla32_fa29_11_xor1;
  wire s_csamul_cla32_fa29_11_and1;
  wire s_csamul_cla32_fa29_11_or0;
  wire s_csamul_cla32_and30_11;
  wire s_csamul_cla32_fa30_11_xor0;
  wire s_csamul_cla32_fa30_11_and0;
  wire s_csamul_cla32_fa30_11_xor1;
  wire s_csamul_cla32_fa30_11_and1;
  wire s_csamul_cla32_fa30_11_or0;
  wire s_csamul_cla32_nand31_11;
  wire s_csamul_cla32_ha31_11_xor0;
  wire s_csamul_cla32_ha31_11_and0;
  wire s_csamul_cla32_and0_12;
  wire s_csamul_cla32_fa0_12_xor0;
  wire s_csamul_cla32_fa0_12_and0;
  wire s_csamul_cla32_fa0_12_xor1;
  wire s_csamul_cla32_fa0_12_and1;
  wire s_csamul_cla32_fa0_12_or0;
  wire s_csamul_cla32_and1_12;
  wire s_csamul_cla32_fa1_12_xor0;
  wire s_csamul_cla32_fa1_12_and0;
  wire s_csamul_cla32_fa1_12_xor1;
  wire s_csamul_cla32_fa1_12_and1;
  wire s_csamul_cla32_fa1_12_or0;
  wire s_csamul_cla32_and2_12;
  wire s_csamul_cla32_fa2_12_xor0;
  wire s_csamul_cla32_fa2_12_and0;
  wire s_csamul_cla32_fa2_12_xor1;
  wire s_csamul_cla32_fa2_12_and1;
  wire s_csamul_cla32_fa2_12_or0;
  wire s_csamul_cla32_and3_12;
  wire s_csamul_cla32_fa3_12_xor0;
  wire s_csamul_cla32_fa3_12_and0;
  wire s_csamul_cla32_fa3_12_xor1;
  wire s_csamul_cla32_fa3_12_and1;
  wire s_csamul_cla32_fa3_12_or0;
  wire s_csamul_cla32_and4_12;
  wire s_csamul_cla32_fa4_12_xor0;
  wire s_csamul_cla32_fa4_12_and0;
  wire s_csamul_cla32_fa4_12_xor1;
  wire s_csamul_cla32_fa4_12_and1;
  wire s_csamul_cla32_fa4_12_or0;
  wire s_csamul_cla32_and5_12;
  wire s_csamul_cla32_fa5_12_xor0;
  wire s_csamul_cla32_fa5_12_and0;
  wire s_csamul_cla32_fa5_12_xor1;
  wire s_csamul_cla32_fa5_12_and1;
  wire s_csamul_cla32_fa5_12_or0;
  wire s_csamul_cla32_and6_12;
  wire s_csamul_cla32_fa6_12_xor0;
  wire s_csamul_cla32_fa6_12_and0;
  wire s_csamul_cla32_fa6_12_xor1;
  wire s_csamul_cla32_fa6_12_and1;
  wire s_csamul_cla32_fa6_12_or0;
  wire s_csamul_cla32_and7_12;
  wire s_csamul_cla32_fa7_12_xor0;
  wire s_csamul_cla32_fa7_12_and0;
  wire s_csamul_cla32_fa7_12_xor1;
  wire s_csamul_cla32_fa7_12_and1;
  wire s_csamul_cla32_fa7_12_or0;
  wire s_csamul_cla32_and8_12;
  wire s_csamul_cla32_fa8_12_xor0;
  wire s_csamul_cla32_fa8_12_and0;
  wire s_csamul_cla32_fa8_12_xor1;
  wire s_csamul_cla32_fa8_12_and1;
  wire s_csamul_cla32_fa8_12_or0;
  wire s_csamul_cla32_and9_12;
  wire s_csamul_cla32_fa9_12_xor0;
  wire s_csamul_cla32_fa9_12_and0;
  wire s_csamul_cla32_fa9_12_xor1;
  wire s_csamul_cla32_fa9_12_and1;
  wire s_csamul_cla32_fa9_12_or0;
  wire s_csamul_cla32_and10_12;
  wire s_csamul_cla32_fa10_12_xor0;
  wire s_csamul_cla32_fa10_12_and0;
  wire s_csamul_cla32_fa10_12_xor1;
  wire s_csamul_cla32_fa10_12_and1;
  wire s_csamul_cla32_fa10_12_or0;
  wire s_csamul_cla32_and11_12;
  wire s_csamul_cla32_fa11_12_xor0;
  wire s_csamul_cla32_fa11_12_and0;
  wire s_csamul_cla32_fa11_12_xor1;
  wire s_csamul_cla32_fa11_12_and1;
  wire s_csamul_cla32_fa11_12_or0;
  wire s_csamul_cla32_and12_12;
  wire s_csamul_cla32_fa12_12_xor0;
  wire s_csamul_cla32_fa12_12_and0;
  wire s_csamul_cla32_fa12_12_xor1;
  wire s_csamul_cla32_fa12_12_and1;
  wire s_csamul_cla32_fa12_12_or0;
  wire s_csamul_cla32_and13_12;
  wire s_csamul_cla32_fa13_12_xor0;
  wire s_csamul_cla32_fa13_12_and0;
  wire s_csamul_cla32_fa13_12_xor1;
  wire s_csamul_cla32_fa13_12_and1;
  wire s_csamul_cla32_fa13_12_or0;
  wire s_csamul_cla32_and14_12;
  wire s_csamul_cla32_fa14_12_xor0;
  wire s_csamul_cla32_fa14_12_and0;
  wire s_csamul_cla32_fa14_12_xor1;
  wire s_csamul_cla32_fa14_12_and1;
  wire s_csamul_cla32_fa14_12_or0;
  wire s_csamul_cla32_and15_12;
  wire s_csamul_cla32_fa15_12_xor0;
  wire s_csamul_cla32_fa15_12_and0;
  wire s_csamul_cla32_fa15_12_xor1;
  wire s_csamul_cla32_fa15_12_and1;
  wire s_csamul_cla32_fa15_12_or0;
  wire s_csamul_cla32_and16_12;
  wire s_csamul_cla32_fa16_12_xor0;
  wire s_csamul_cla32_fa16_12_and0;
  wire s_csamul_cla32_fa16_12_xor1;
  wire s_csamul_cla32_fa16_12_and1;
  wire s_csamul_cla32_fa16_12_or0;
  wire s_csamul_cla32_and17_12;
  wire s_csamul_cla32_fa17_12_xor0;
  wire s_csamul_cla32_fa17_12_and0;
  wire s_csamul_cla32_fa17_12_xor1;
  wire s_csamul_cla32_fa17_12_and1;
  wire s_csamul_cla32_fa17_12_or0;
  wire s_csamul_cla32_and18_12;
  wire s_csamul_cla32_fa18_12_xor0;
  wire s_csamul_cla32_fa18_12_and0;
  wire s_csamul_cla32_fa18_12_xor1;
  wire s_csamul_cla32_fa18_12_and1;
  wire s_csamul_cla32_fa18_12_or0;
  wire s_csamul_cla32_and19_12;
  wire s_csamul_cla32_fa19_12_xor0;
  wire s_csamul_cla32_fa19_12_and0;
  wire s_csamul_cla32_fa19_12_xor1;
  wire s_csamul_cla32_fa19_12_and1;
  wire s_csamul_cla32_fa19_12_or0;
  wire s_csamul_cla32_and20_12;
  wire s_csamul_cla32_fa20_12_xor0;
  wire s_csamul_cla32_fa20_12_and0;
  wire s_csamul_cla32_fa20_12_xor1;
  wire s_csamul_cla32_fa20_12_and1;
  wire s_csamul_cla32_fa20_12_or0;
  wire s_csamul_cla32_and21_12;
  wire s_csamul_cla32_fa21_12_xor0;
  wire s_csamul_cla32_fa21_12_and0;
  wire s_csamul_cla32_fa21_12_xor1;
  wire s_csamul_cla32_fa21_12_and1;
  wire s_csamul_cla32_fa21_12_or0;
  wire s_csamul_cla32_and22_12;
  wire s_csamul_cla32_fa22_12_xor0;
  wire s_csamul_cla32_fa22_12_and0;
  wire s_csamul_cla32_fa22_12_xor1;
  wire s_csamul_cla32_fa22_12_and1;
  wire s_csamul_cla32_fa22_12_or0;
  wire s_csamul_cla32_and23_12;
  wire s_csamul_cla32_fa23_12_xor0;
  wire s_csamul_cla32_fa23_12_and0;
  wire s_csamul_cla32_fa23_12_xor1;
  wire s_csamul_cla32_fa23_12_and1;
  wire s_csamul_cla32_fa23_12_or0;
  wire s_csamul_cla32_and24_12;
  wire s_csamul_cla32_fa24_12_xor0;
  wire s_csamul_cla32_fa24_12_and0;
  wire s_csamul_cla32_fa24_12_xor1;
  wire s_csamul_cla32_fa24_12_and1;
  wire s_csamul_cla32_fa24_12_or0;
  wire s_csamul_cla32_and25_12;
  wire s_csamul_cla32_fa25_12_xor0;
  wire s_csamul_cla32_fa25_12_and0;
  wire s_csamul_cla32_fa25_12_xor1;
  wire s_csamul_cla32_fa25_12_and1;
  wire s_csamul_cla32_fa25_12_or0;
  wire s_csamul_cla32_and26_12;
  wire s_csamul_cla32_fa26_12_xor0;
  wire s_csamul_cla32_fa26_12_and0;
  wire s_csamul_cla32_fa26_12_xor1;
  wire s_csamul_cla32_fa26_12_and1;
  wire s_csamul_cla32_fa26_12_or0;
  wire s_csamul_cla32_and27_12;
  wire s_csamul_cla32_fa27_12_xor0;
  wire s_csamul_cla32_fa27_12_and0;
  wire s_csamul_cla32_fa27_12_xor1;
  wire s_csamul_cla32_fa27_12_and1;
  wire s_csamul_cla32_fa27_12_or0;
  wire s_csamul_cla32_and28_12;
  wire s_csamul_cla32_fa28_12_xor0;
  wire s_csamul_cla32_fa28_12_and0;
  wire s_csamul_cla32_fa28_12_xor1;
  wire s_csamul_cla32_fa28_12_and1;
  wire s_csamul_cla32_fa28_12_or0;
  wire s_csamul_cla32_and29_12;
  wire s_csamul_cla32_fa29_12_xor0;
  wire s_csamul_cla32_fa29_12_and0;
  wire s_csamul_cla32_fa29_12_xor1;
  wire s_csamul_cla32_fa29_12_and1;
  wire s_csamul_cla32_fa29_12_or0;
  wire s_csamul_cla32_and30_12;
  wire s_csamul_cla32_fa30_12_xor0;
  wire s_csamul_cla32_fa30_12_and0;
  wire s_csamul_cla32_fa30_12_xor1;
  wire s_csamul_cla32_fa30_12_and1;
  wire s_csamul_cla32_fa30_12_or0;
  wire s_csamul_cla32_nand31_12;
  wire s_csamul_cla32_ha31_12_xor0;
  wire s_csamul_cla32_ha31_12_and0;
  wire s_csamul_cla32_and0_13;
  wire s_csamul_cla32_fa0_13_xor0;
  wire s_csamul_cla32_fa0_13_and0;
  wire s_csamul_cla32_fa0_13_xor1;
  wire s_csamul_cla32_fa0_13_and1;
  wire s_csamul_cla32_fa0_13_or0;
  wire s_csamul_cla32_and1_13;
  wire s_csamul_cla32_fa1_13_xor0;
  wire s_csamul_cla32_fa1_13_and0;
  wire s_csamul_cla32_fa1_13_xor1;
  wire s_csamul_cla32_fa1_13_and1;
  wire s_csamul_cla32_fa1_13_or0;
  wire s_csamul_cla32_and2_13;
  wire s_csamul_cla32_fa2_13_xor0;
  wire s_csamul_cla32_fa2_13_and0;
  wire s_csamul_cla32_fa2_13_xor1;
  wire s_csamul_cla32_fa2_13_and1;
  wire s_csamul_cla32_fa2_13_or0;
  wire s_csamul_cla32_and3_13;
  wire s_csamul_cla32_fa3_13_xor0;
  wire s_csamul_cla32_fa3_13_and0;
  wire s_csamul_cla32_fa3_13_xor1;
  wire s_csamul_cla32_fa3_13_and1;
  wire s_csamul_cla32_fa3_13_or0;
  wire s_csamul_cla32_and4_13;
  wire s_csamul_cla32_fa4_13_xor0;
  wire s_csamul_cla32_fa4_13_and0;
  wire s_csamul_cla32_fa4_13_xor1;
  wire s_csamul_cla32_fa4_13_and1;
  wire s_csamul_cla32_fa4_13_or0;
  wire s_csamul_cla32_and5_13;
  wire s_csamul_cla32_fa5_13_xor0;
  wire s_csamul_cla32_fa5_13_and0;
  wire s_csamul_cla32_fa5_13_xor1;
  wire s_csamul_cla32_fa5_13_and1;
  wire s_csamul_cla32_fa5_13_or0;
  wire s_csamul_cla32_and6_13;
  wire s_csamul_cla32_fa6_13_xor0;
  wire s_csamul_cla32_fa6_13_and0;
  wire s_csamul_cla32_fa6_13_xor1;
  wire s_csamul_cla32_fa6_13_and1;
  wire s_csamul_cla32_fa6_13_or0;
  wire s_csamul_cla32_and7_13;
  wire s_csamul_cla32_fa7_13_xor0;
  wire s_csamul_cla32_fa7_13_and0;
  wire s_csamul_cla32_fa7_13_xor1;
  wire s_csamul_cla32_fa7_13_and1;
  wire s_csamul_cla32_fa7_13_or0;
  wire s_csamul_cla32_and8_13;
  wire s_csamul_cla32_fa8_13_xor0;
  wire s_csamul_cla32_fa8_13_and0;
  wire s_csamul_cla32_fa8_13_xor1;
  wire s_csamul_cla32_fa8_13_and1;
  wire s_csamul_cla32_fa8_13_or0;
  wire s_csamul_cla32_and9_13;
  wire s_csamul_cla32_fa9_13_xor0;
  wire s_csamul_cla32_fa9_13_and0;
  wire s_csamul_cla32_fa9_13_xor1;
  wire s_csamul_cla32_fa9_13_and1;
  wire s_csamul_cla32_fa9_13_or0;
  wire s_csamul_cla32_and10_13;
  wire s_csamul_cla32_fa10_13_xor0;
  wire s_csamul_cla32_fa10_13_and0;
  wire s_csamul_cla32_fa10_13_xor1;
  wire s_csamul_cla32_fa10_13_and1;
  wire s_csamul_cla32_fa10_13_or0;
  wire s_csamul_cla32_and11_13;
  wire s_csamul_cla32_fa11_13_xor0;
  wire s_csamul_cla32_fa11_13_and0;
  wire s_csamul_cla32_fa11_13_xor1;
  wire s_csamul_cla32_fa11_13_and1;
  wire s_csamul_cla32_fa11_13_or0;
  wire s_csamul_cla32_and12_13;
  wire s_csamul_cla32_fa12_13_xor0;
  wire s_csamul_cla32_fa12_13_and0;
  wire s_csamul_cla32_fa12_13_xor1;
  wire s_csamul_cla32_fa12_13_and1;
  wire s_csamul_cla32_fa12_13_or0;
  wire s_csamul_cla32_and13_13;
  wire s_csamul_cla32_fa13_13_xor0;
  wire s_csamul_cla32_fa13_13_and0;
  wire s_csamul_cla32_fa13_13_xor1;
  wire s_csamul_cla32_fa13_13_and1;
  wire s_csamul_cla32_fa13_13_or0;
  wire s_csamul_cla32_and14_13;
  wire s_csamul_cla32_fa14_13_xor0;
  wire s_csamul_cla32_fa14_13_and0;
  wire s_csamul_cla32_fa14_13_xor1;
  wire s_csamul_cla32_fa14_13_and1;
  wire s_csamul_cla32_fa14_13_or0;
  wire s_csamul_cla32_and15_13;
  wire s_csamul_cla32_fa15_13_xor0;
  wire s_csamul_cla32_fa15_13_and0;
  wire s_csamul_cla32_fa15_13_xor1;
  wire s_csamul_cla32_fa15_13_and1;
  wire s_csamul_cla32_fa15_13_or0;
  wire s_csamul_cla32_and16_13;
  wire s_csamul_cla32_fa16_13_xor0;
  wire s_csamul_cla32_fa16_13_and0;
  wire s_csamul_cla32_fa16_13_xor1;
  wire s_csamul_cla32_fa16_13_and1;
  wire s_csamul_cla32_fa16_13_or0;
  wire s_csamul_cla32_and17_13;
  wire s_csamul_cla32_fa17_13_xor0;
  wire s_csamul_cla32_fa17_13_and0;
  wire s_csamul_cla32_fa17_13_xor1;
  wire s_csamul_cla32_fa17_13_and1;
  wire s_csamul_cla32_fa17_13_or0;
  wire s_csamul_cla32_and18_13;
  wire s_csamul_cla32_fa18_13_xor0;
  wire s_csamul_cla32_fa18_13_and0;
  wire s_csamul_cla32_fa18_13_xor1;
  wire s_csamul_cla32_fa18_13_and1;
  wire s_csamul_cla32_fa18_13_or0;
  wire s_csamul_cla32_and19_13;
  wire s_csamul_cla32_fa19_13_xor0;
  wire s_csamul_cla32_fa19_13_and0;
  wire s_csamul_cla32_fa19_13_xor1;
  wire s_csamul_cla32_fa19_13_and1;
  wire s_csamul_cla32_fa19_13_or0;
  wire s_csamul_cla32_and20_13;
  wire s_csamul_cla32_fa20_13_xor0;
  wire s_csamul_cla32_fa20_13_and0;
  wire s_csamul_cla32_fa20_13_xor1;
  wire s_csamul_cla32_fa20_13_and1;
  wire s_csamul_cla32_fa20_13_or0;
  wire s_csamul_cla32_and21_13;
  wire s_csamul_cla32_fa21_13_xor0;
  wire s_csamul_cla32_fa21_13_and0;
  wire s_csamul_cla32_fa21_13_xor1;
  wire s_csamul_cla32_fa21_13_and1;
  wire s_csamul_cla32_fa21_13_or0;
  wire s_csamul_cla32_and22_13;
  wire s_csamul_cla32_fa22_13_xor0;
  wire s_csamul_cla32_fa22_13_and0;
  wire s_csamul_cla32_fa22_13_xor1;
  wire s_csamul_cla32_fa22_13_and1;
  wire s_csamul_cla32_fa22_13_or0;
  wire s_csamul_cla32_and23_13;
  wire s_csamul_cla32_fa23_13_xor0;
  wire s_csamul_cla32_fa23_13_and0;
  wire s_csamul_cla32_fa23_13_xor1;
  wire s_csamul_cla32_fa23_13_and1;
  wire s_csamul_cla32_fa23_13_or0;
  wire s_csamul_cla32_and24_13;
  wire s_csamul_cla32_fa24_13_xor0;
  wire s_csamul_cla32_fa24_13_and0;
  wire s_csamul_cla32_fa24_13_xor1;
  wire s_csamul_cla32_fa24_13_and1;
  wire s_csamul_cla32_fa24_13_or0;
  wire s_csamul_cla32_and25_13;
  wire s_csamul_cla32_fa25_13_xor0;
  wire s_csamul_cla32_fa25_13_and0;
  wire s_csamul_cla32_fa25_13_xor1;
  wire s_csamul_cla32_fa25_13_and1;
  wire s_csamul_cla32_fa25_13_or0;
  wire s_csamul_cla32_and26_13;
  wire s_csamul_cla32_fa26_13_xor0;
  wire s_csamul_cla32_fa26_13_and0;
  wire s_csamul_cla32_fa26_13_xor1;
  wire s_csamul_cla32_fa26_13_and1;
  wire s_csamul_cla32_fa26_13_or0;
  wire s_csamul_cla32_and27_13;
  wire s_csamul_cla32_fa27_13_xor0;
  wire s_csamul_cla32_fa27_13_and0;
  wire s_csamul_cla32_fa27_13_xor1;
  wire s_csamul_cla32_fa27_13_and1;
  wire s_csamul_cla32_fa27_13_or0;
  wire s_csamul_cla32_and28_13;
  wire s_csamul_cla32_fa28_13_xor0;
  wire s_csamul_cla32_fa28_13_and0;
  wire s_csamul_cla32_fa28_13_xor1;
  wire s_csamul_cla32_fa28_13_and1;
  wire s_csamul_cla32_fa28_13_or0;
  wire s_csamul_cla32_and29_13;
  wire s_csamul_cla32_fa29_13_xor0;
  wire s_csamul_cla32_fa29_13_and0;
  wire s_csamul_cla32_fa29_13_xor1;
  wire s_csamul_cla32_fa29_13_and1;
  wire s_csamul_cla32_fa29_13_or0;
  wire s_csamul_cla32_and30_13;
  wire s_csamul_cla32_fa30_13_xor0;
  wire s_csamul_cla32_fa30_13_and0;
  wire s_csamul_cla32_fa30_13_xor1;
  wire s_csamul_cla32_fa30_13_and1;
  wire s_csamul_cla32_fa30_13_or0;
  wire s_csamul_cla32_nand31_13;
  wire s_csamul_cla32_ha31_13_xor0;
  wire s_csamul_cla32_ha31_13_and0;
  wire s_csamul_cla32_and0_14;
  wire s_csamul_cla32_fa0_14_xor0;
  wire s_csamul_cla32_fa0_14_and0;
  wire s_csamul_cla32_fa0_14_xor1;
  wire s_csamul_cla32_fa0_14_and1;
  wire s_csamul_cla32_fa0_14_or0;
  wire s_csamul_cla32_and1_14;
  wire s_csamul_cla32_fa1_14_xor0;
  wire s_csamul_cla32_fa1_14_and0;
  wire s_csamul_cla32_fa1_14_xor1;
  wire s_csamul_cla32_fa1_14_and1;
  wire s_csamul_cla32_fa1_14_or0;
  wire s_csamul_cla32_and2_14;
  wire s_csamul_cla32_fa2_14_xor0;
  wire s_csamul_cla32_fa2_14_and0;
  wire s_csamul_cla32_fa2_14_xor1;
  wire s_csamul_cla32_fa2_14_and1;
  wire s_csamul_cla32_fa2_14_or0;
  wire s_csamul_cla32_and3_14;
  wire s_csamul_cla32_fa3_14_xor0;
  wire s_csamul_cla32_fa3_14_and0;
  wire s_csamul_cla32_fa3_14_xor1;
  wire s_csamul_cla32_fa3_14_and1;
  wire s_csamul_cla32_fa3_14_or0;
  wire s_csamul_cla32_and4_14;
  wire s_csamul_cla32_fa4_14_xor0;
  wire s_csamul_cla32_fa4_14_and0;
  wire s_csamul_cla32_fa4_14_xor1;
  wire s_csamul_cla32_fa4_14_and1;
  wire s_csamul_cla32_fa4_14_or0;
  wire s_csamul_cla32_and5_14;
  wire s_csamul_cla32_fa5_14_xor0;
  wire s_csamul_cla32_fa5_14_and0;
  wire s_csamul_cla32_fa5_14_xor1;
  wire s_csamul_cla32_fa5_14_and1;
  wire s_csamul_cla32_fa5_14_or0;
  wire s_csamul_cla32_and6_14;
  wire s_csamul_cla32_fa6_14_xor0;
  wire s_csamul_cla32_fa6_14_and0;
  wire s_csamul_cla32_fa6_14_xor1;
  wire s_csamul_cla32_fa6_14_and1;
  wire s_csamul_cla32_fa6_14_or0;
  wire s_csamul_cla32_and7_14;
  wire s_csamul_cla32_fa7_14_xor0;
  wire s_csamul_cla32_fa7_14_and0;
  wire s_csamul_cla32_fa7_14_xor1;
  wire s_csamul_cla32_fa7_14_and1;
  wire s_csamul_cla32_fa7_14_or0;
  wire s_csamul_cla32_and8_14;
  wire s_csamul_cla32_fa8_14_xor0;
  wire s_csamul_cla32_fa8_14_and0;
  wire s_csamul_cla32_fa8_14_xor1;
  wire s_csamul_cla32_fa8_14_and1;
  wire s_csamul_cla32_fa8_14_or0;
  wire s_csamul_cla32_and9_14;
  wire s_csamul_cla32_fa9_14_xor0;
  wire s_csamul_cla32_fa9_14_and0;
  wire s_csamul_cla32_fa9_14_xor1;
  wire s_csamul_cla32_fa9_14_and1;
  wire s_csamul_cla32_fa9_14_or0;
  wire s_csamul_cla32_and10_14;
  wire s_csamul_cla32_fa10_14_xor0;
  wire s_csamul_cla32_fa10_14_and0;
  wire s_csamul_cla32_fa10_14_xor1;
  wire s_csamul_cla32_fa10_14_and1;
  wire s_csamul_cla32_fa10_14_or0;
  wire s_csamul_cla32_and11_14;
  wire s_csamul_cla32_fa11_14_xor0;
  wire s_csamul_cla32_fa11_14_and0;
  wire s_csamul_cla32_fa11_14_xor1;
  wire s_csamul_cla32_fa11_14_and1;
  wire s_csamul_cla32_fa11_14_or0;
  wire s_csamul_cla32_and12_14;
  wire s_csamul_cla32_fa12_14_xor0;
  wire s_csamul_cla32_fa12_14_and0;
  wire s_csamul_cla32_fa12_14_xor1;
  wire s_csamul_cla32_fa12_14_and1;
  wire s_csamul_cla32_fa12_14_or0;
  wire s_csamul_cla32_and13_14;
  wire s_csamul_cla32_fa13_14_xor0;
  wire s_csamul_cla32_fa13_14_and0;
  wire s_csamul_cla32_fa13_14_xor1;
  wire s_csamul_cla32_fa13_14_and1;
  wire s_csamul_cla32_fa13_14_or0;
  wire s_csamul_cla32_and14_14;
  wire s_csamul_cla32_fa14_14_xor0;
  wire s_csamul_cla32_fa14_14_and0;
  wire s_csamul_cla32_fa14_14_xor1;
  wire s_csamul_cla32_fa14_14_and1;
  wire s_csamul_cla32_fa14_14_or0;
  wire s_csamul_cla32_and15_14;
  wire s_csamul_cla32_fa15_14_xor0;
  wire s_csamul_cla32_fa15_14_and0;
  wire s_csamul_cla32_fa15_14_xor1;
  wire s_csamul_cla32_fa15_14_and1;
  wire s_csamul_cla32_fa15_14_or0;
  wire s_csamul_cla32_and16_14;
  wire s_csamul_cla32_fa16_14_xor0;
  wire s_csamul_cla32_fa16_14_and0;
  wire s_csamul_cla32_fa16_14_xor1;
  wire s_csamul_cla32_fa16_14_and1;
  wire s_csamul_cla32_fa16_14_or0;
  wire s_csamul_cla32_and17_14;
  wire s_csamul_cla32_fa17_14_xor0;
  wire s_csamul_cla32_fa17_14_and0;
  wire s_csamul_cla32_fa17_14_xor1;
  wire s_csamul_cla32_fa17_14_and1;
  wire s_csamul_cla32_fa17_14_or0;
  wire s_csamul_cla32_and18_14;
  wire s_csamul_cla32_fa18_14_xor0;
  wire s_csamul_cla32_fa18_14_and0;
  wire s_csamul_cla32_fa18_14_xor1;
  wire s_csamul_cla32_fa18_14_and1;
  wire s_csamul_cla32_fa18_14_or0;
  wire s_csamul_cla32_and19_14;
  wire s_csamul_cla32_fa19_14_xor0;
  wire s_csamul_cla32_fa19_14_and0;
  wire s_csamul_cla32_fa19_14_xor1;
  wire s_csamul_cla32_fa19_14_and1;
  wire s_csamul_cla32_fa19_14_or0;
  wire s_csamul_cla32_and20_14;
  wire s_csamul_cla32_fa20_14_xor0;
  wire s_csamul_cla32_fa20_14_and0;
  wire s_csamul_cla32_fa20_14_xor1;
  wire s_csamul_cla32_fa20_14_and1;
  wire s_csamul_cla32_fa20_14_or0;
  wire s_csamul_cla32_and21_14;
  wire s_csamul_cla32_fa21_14_xor0;
  wire s_csamul_cla32_fa21_14_and0;
  wire s_csamul_cla32_fa21_14_xor1;
  wire s_csamul_cla32_fa21_14_and1;
  wire s_csamul_cla32_fa21_14_or0;
  wire s_csamul_cla32_and22_14;
  wire s_csamul_cla32_fa22_14_xor0;
  wire s_csamul_cla32_fa22_14_and0;
  wire s_csamul_cla32_fa22_14_xor1;
  wire s_csamul_cla32_fa22_14_and1;
  wire s_csamul_cla32_fa22_14_or0;
  wire s_csamul_cla32_and23_14;
  wire s_csamul_cla32_fa23_14_xor0;
  wire s_csamul_cla32_fa23_14_and0;
  wire s_csamul_cla32_fa23_14_xor1;
  wire s_csamul_cla32_fa23_14_and1;
  wire s_csamul_cla32_fa23_14_or0;
  wire s_csamul_cla32_and24_14;
  wire s_csamul_cla32_fa24_14_xor0;
  wire s_csamul_cla32_fa24_14_and0;
  wire s_csamul_cla32_fa24_14_xor1;
  wire s_csamul_cla32_fa24_14_and1;
  wire s_csamul_cla32_fa24_14_or0;
  wire s_csamul_cla32_and25_14;
  wire s_csamul_cla32_fa25_14_xor0;
  wire s_csamul_cla32_fa25_14_and0;
  wire s_csamul_cla32_fa25_14_xor1;
  wire s_csamul_cla32_fa25_14_and1;
  wire s_csamul_cla32_fa25_14_or0;
  wire s_csamul_cla32_and26_14;
  wire s_csamul_cla32_fa26_14_xor0;
  wire s_csamul_cla32_fa26_14_and0;
  wire s_csamul_cla32_fa26_14_xor1;
  wire s_csamul_cla32_fa26_14_and1;
  wire s_csamul_cla32_fa26_14_or0;
  wire s_csamul_cla32_and27_14;
  wire s_csamul_cla32_fa27_14_xor0;
  wire s_csamul_cla32_fa27_14_and0;
  wire s_csamul_cla32_fa27_14_xor1;
  wire s_csamul_cla32_fa27_14_and1;
  wire s_csamul_cla32_fa27_14_or0;
  wire s_csamul_cla32_and28_14;
  wire s_csamul_cla32_fa28_14_xor0;
  wire s_csamul_cla32_fa28_14_and0;
  wire s_csamul_cla32_fa28_14_xor1;
  wire s_csamul_cla32_fa28_14_and1;
  wire s_csamul_cla32_fa28_14_or0;
  wire s_csamul_cla32_and29_14;
  wire s_csamul_cla32_fa29_14_xor0;
  wire s_csamul_cla32_fa29_14_and0;
  wire s_csamul_cla32_fa29_14_xor1;
  wire s_csamul_cla32_fa29_14_and1;
  wire s_csamul_cla32_fa29_14_or0;
  wire s_csamul_cla32_and30_14;
  wire s_csamul_cla32_fa30_14_xor0;
  wire s_csamul_cla32_fa30_14_and0;
  wire s_csamul_cla32_fa30_14_xor1;
  wire s_csamul_cla32_fa30_14_and1;
  wire s_csamul_cla32_fa30_14_or0;
  wire s_csamul_cla32_nand31_14;
  wire s_csamul_cla32_ha31_14_xor0;
  wire s_csamul_cla32_ha31_14_and0;
  wire s_csamul_cla32_and0_15;
  wire s_csamul_cla32_fa0_15_xor0;
  wire s_csamul_cla32_fa0_15_and0;
  wire s_csamul_cla32_fa0_15_xor1;
  wire s_csamul_cla32_fa0_15_and1;
  wire s_csamul_cla32_fa0_15_or0;
  wire s_csamul_cla32_and1_15;
  wire s_csamul_cla32_fa1_15_xor0;
  wire s_csamul_cla32_fa1_15_and0;
  wire s_csamul_cla32_fa1_15_xor1;
  wire s_csamul_cla32_fa1_15_and1;
  wire s_csamul_cla32_fa1_15_or0;
  wire s_csamul_cla32_and2_15;
  wire s_csamul_cla32_fa2_15_xor0;
  wire s_csamul_cla32_fa2_15_and0;
  wire s_csamul_cla32_fa2_15_xor1;
  wire s_csamul_cla32_fa2_15_and1;
  wire s_csamul_cla32_fa2_15_or0;
  wire s_csamul_cla32_and3_15;
  wire s_csamul_cla32_fa3_15_xor0;
  wire s_csamul_cla32_fa3_15_and0;
  wire s_csamul_cla32_fa3_15_xor1;
  wire s_csamul_cla32_fa3_15_and1;
  wire s_csamul_cla32_fa3_15_or0;
  wire s_csamul_cla32_and4_15;
  wire s_csamul_cla32_fa4_15_xor0;
  wire s_csamul_cla32_fa4_15_and0;
  wire s_csamul_cla32_fa4_15_xor1;
  wire s_csamul_cla32_fa4_15_and1;
  wire s_csamul_cla32_fa4_15_or0;
  wire s_csamul_cla32_and5_15;
  wire s_csamul_cla32_fa5_15_xor0;
  wire s_csamul_cla32_fa5_15_and0;
  wire s_csamul_cla32_fa5_15_xor1;
  wire s_csamul_cla32_fa5_15_and1;
  wire s_csamul_cla32_fa5_15_or0;
  wire s_csamul_cla32_and6_15;
  wire s_csamul_cla32_fa6_15_xor0;
  wire s_csamul_cla32_fa6_15_and0;
  wire s_csamul_cla32_fa6_15_xor1;
  wire s_csamul_cla32_fa6_15_and1;
  wire s_csamul_cla32_fa6_15_or0;
  wire s_csamul_cla32_and7_15;
  wire s_csamul_cla32_fa7_15_xor0;
  wire s_csamul_cla32_fa7_15_and0;
  wire s_csamul_cla32_fa7_15_xor1;
  wire s_csamul_cla32_fa7_15_and1;
  wire s_csamul_cla32_fa7_15_or0;
  wire s_csamul_cla32_and8_15;
  wire s_csamul_cla32_fa8_15_xor0;
  wire s_csamul_cla32_fa8_15_and0;
  wire s_csamul_cla32_fa8_15_xor1;
  wire s_csamul_cla32_fa8_15_and1;
  wire s_csamul_cla32_fa8_15_or0;
  wire s_csamul_cla32_and9_15;
  wire s_csamul_cla32_fa9_15_xor0;
  wire s_csamul_cla32_fa9_15_and0;
  wire s_csamul_cla32_fa9_15_xor1;
  wire s_csamul_cla32_fa9_15_and1;
  wire s_csamul_cla32_fa9_15_or0;
  wire s_csamul_cla32_and10_15;
  wire s_csamul_cla32_fa10_15_xor0;
  wire s_csamul_cla32_fa10_15_and0;
  wire s_csamul_cla32_fa10_15_xor1;
  wire s_csamul_cla32_fa10_15_and1;
  wire s_csamul_cla32_fa10_15_or0;
  wire s_csamul_cla32_and11_15;
  wire s_csamul_cla32_fa11_15_xor0;
  wire s_csamul_cla32_fa11_15_and0;
  wire s_csamul_cla32_fa11_15_xor1;
  wire s_csamul_cla32_fa11_15_and1;
  wire s_csamul_cla32_fa11_15_or0;
  wire s_csamul_cla32_and12_15;
  wire s_csamul_cla32_fa12_15_xor0;
  wire s_csamul_cla32_fa12_15_and0;
  wire s_csamul_cla32_fa12_15_xor1;
  wire s_csamul_cla32_fa12_15_and1;
  wire s_csamul_cla32_fa12_15_or0;
  wire s_csamul_cla32_and13_15;
  wire s_csamul_cla32_fa13_15_xor0;
  wire s_csamul_cla32_fa13_15_and0;
  wire s_csamul_cla32_fa13_15_xor1;
  wire s_csamul_cla32_fa13_15_and1;
  wire s_csamul_cla32_fa13_15_or0;
  wire s_csamul_cla32_and14_15;
  wire s_csamul_cla32_fa14_15_xor0;
  wire s_csamul_cla32_fa14_15_and0;
  wire s_csamul_cla32_fa14_15_xor1;
  wire s_csamul_cla32_fa14_15_and1;
  wire s_csamul_cla32_fa14_15_or0;
  wire s_csamul_cla32_and15_15;
  wire s_csamul_cla32_fa15_15_xor0;
  wire s_csamul_cla32_fa15_15_and0;
  wire s_csamul_cla32_fa15_15_xor1;
  wire s_csamul_cla32_fa15_15_and1;
  wire s_csamul_cla32_fa15_15_or0;
  wire s_csamul_cla32_and16_15;
  wire s_csamul_cla32_fa16_15_xor0;
  wire s_csamul_cla32_fa16_15_and0;
  wire s_csamul_cla32_fa16_15_xor1;
  wire s_csamul_cla32_fa16_15_and1;
  wire s_csamul_cla32_fa16_15_or0;
  wire s_csamul_cla32_and17_15;
  wire s_csamul_cla32_fa17_15_xor0;
  wire s_csamul_cla32_fa17_15_and0;
  wire s_csamul_cla32_fa17_15_xor1;
  wire s_csamul_cla32_fa17_15_and1;
  wire s_csamul_cla32_fa17_15_or0;
  wire s_csamul_cla32_and18_15;
  wire s_csamul_cla32_fa18_15_xor0;
  wire s_csamul_cla32_fa18_15_and0;
  wire s_csamul_cla32_fa18_15_xor1;
  wire s_csamul_cla32_fa18_15_and1;
  wire s_csamul_cla32_fa18_15_or0;
  wire s_csamul_cla32_and19_15;
  wire s_csamul_cla32_fa19_15_xor0;
  wire s_csamul_cla32_fa19_15_and0;
  wire s_csamul_cla32_fa19_15_xor1;
  wire s_csamul_cla32_fa19_15_and1;
  wire s_csamul_cla32_fa19_15_or0;
  wire s_csamul_cla32_and20_15;
  wire s_csamul_cla32_fa20_15_xor0;
  wire s_csamul_cla32_fa20_15_and0;
  wire s_csamul_cla32_fa20_15_xor1;
  wire s_csamul_cla32_fa20_15_and1;
  wire s_csamul_cla32_fa20_15_or0;
  wire s_csamul_cla32_and21_15;
  wire s_csamul_cla32_fa21_15_xor0;
  wire s_csamul_cla32_fa21_15_and0;
  wire s_csamul_cla32_fa21_15_xor1;
  wire s_csamul_cla32_fa21_15_and1;
  wire s_csamul_cla32_fa21_15_or0;
  wire s_csamul_cla32_and22_15;
  wire s_csamul_cla32_fa22_15_xor0;
  wire s_csamul_cla32_fa22_15_and0;
  wire s_csamul_cla32_fa22_15_xor1;
  wire s_csamul_cla32_fa22_15_and1;
  wire s_csamul_cla32_fa22_15_or0;
  wire s_csamul_cla32_and23_15;
  wire s_csamul_cla32_fa23_15_xor0;
  wire s_csamul_cla32_fa23_15_and0;
  wire s_csamul_cla32_fa23_15_xor1;
  wire s_csamul_cla32_fa23_15_and1;
  wire s_csamul_cla32_fa23_15_or0;
  wire s_csamul_cla32_and24_15;
  wire s_csamul_cla32_fa24_15_xor0;
  wire s_csamul_cla32_fa24_15_and0;
  wire s_csamul_cla32_fa24_15_xor1;
  wire s_csamul_cla32_fa24_15_and1;
  wire s_csamul_cla32_fa24_15_or0;
  wire s_csamul_cla32_and25_15;
  wire s_csamul_cla32_fa25_15_xor0;
  wire s_csamul_cla32_fa25_15_and0;
  wire s_csamul_cla32_fa25_15_xor1;
  wire s_csamul_cla32_fa25_15_and1;
  wire s_csamul_cla32_fa25_15_or0;
  wire s_csamul_cla32_and26_15;
  wire s_csamul_cla32_fa26_15_xor0;
  wire s_csamul_cla32_fa26_15_and0;
  wire s_csamul_cla32_fa26_15_xor1;
  wire s_csamul_cla32_fa26_15_and1;
  wire s_csamul_cla32_fa26_15_or0;
  wire s_csamul_cla32_and27_15;
  wire s_csamul_cla32_fa27_15_xor0;
  wire s_csamul_cla32_fa27_15_and0;
  wire s_csamul_cla32_fa27_15_xor1;
  wire s_csamul_cla32_fa27_15_and1;
  wire s_csamul_cla32_fa27_15_or0;
  wire s_csamul_cla32_and28_15;
  wire s_csamul_cla32_fa28_15_xor0;
  wire s_csamul_cla32_fa28_15_and0;
  wire s_csamul_cla32_fa28_15_xor1;
  wire s_csamul_cla32_fa28_15_and1;
  wire s_csamul_cla32_fa28_15_or0;
  wire s_csamul_cla32_and29_15;
  wire s_csamul_cla32_fa29_15_xor0;
  wire s_csamul_cla32_fa29_15_and0;
  wire s_csamul_cla32_fa29_15_xor1;
  wire s_csamul_cla32_fa29_15_and1;
  wire s_csamul_cla32_fa29_15_or0;
  wire s_csamul_cla32_and30_15;
  wire s_csamul_cla32_fa30_15_xor0;
  wire s_csamul_cla32_fa30_15_and0;
  wire s_csamul_cla32_fa30_15_xor1;
  wire s_csamul_cla32_fa30_15_and1;
  wire s_csamul_cla32_fa30_15_or0;
  wire s_csamul_cla32_nand31_15;
  wire s_csamul_cla32_ha31_15_xor0;
  wire s_csamul_cla32_ha31_15_and0;
  wire s_csamul_cla32_and0_16;
  wire s_csamul_cla32_fa0_16_xor0;
  wire s_csamul_cla32_fa0_16_and0;
  wire s_csamul_cla32_fa0_16_xor1;
  wire s_csamul_cla32_fa0_16_and1;
  wire s_csamul_cla32_fa0_16_or0;
  wire s_csamul_cla32_and1_16;
  wire s_csamul_cla32_fa1_16_xor0;
  wire s_csamul_cla32_fa1_16_and0;
  wire s_csamul_cla32_fa1_16_xor1;
  wire s_csamul_cla32_fa1_16_and1;
  wire s_csamul_cla32_fa1_16_or0;
  wire s_csamul_cla32_and2_16;
  wire s_csamul_cla32_fa2_16_xor0;
  wire s_csamul_cla32_fa2_16_and0;
  wire s_csamul_cla32_fa2_16_xor1;
  wire s_csamul_cla32_fa2_16_and1;
  wire s_csamul_cla32_fa2_16_or0;
  wire s_csamul_cla32_and3_16;
  wire s_csamul_cla32_fa3_16_xor0;
  wire s_csamul_cla32_fa3_16_and0;
  wire s_csamul_cla32_fa3_16_xor1;
  wire s_csamul_cla32_fa3_16_and1;
  wire s_csamul_cla32_fa3_16_or0;
  wire s_csamul_cla32_and4_16;
  wire s_csamul_cla32_fa4_16_xor0;
  wire s_csamul_cla32_fa4_16_and0;
  wire s_csamul_cla32_fa4_16_xor1;
  wire s_csamul_cla32_fa4_16_and1;
  wire s_csamul_cla32_fa4_16_or0;
  wire s_csamul_cla32_and5_16;
  wire s_csamul_cla32_fa5_16_xor0;
  wire s_csamul_cla32_fa5_16_and0;
  wire s_csamul_cla32_fa5_16_xor1;
  wire s_csamul_cla32_fa5_16_and1;
  wire s_csamul_cla32_fa5_16_or0;
  wire s_csamul_cla32_and6_16;
  wire s_csamul_cla32_fa6_16_xor0;
  wire s_csamul_cla32_fa6_16_and0;
  wire s_csamul_cla32_fa6_16_xor1;
  wire s_csamul_cla32_fa6_16_and1;
  wire s_csamul_cla32_fa6_16_or0;
  wire s_csamul_cla32_and7_16;
  wire s_csamul_cla32_fa7_16_xor0;
  wire s_csamul_cla32_fa7_16_and0;
  wire s_csamul_cla32_fa7_16_xor1;
  wire s_csamul_cla32_fa7_16_and1;
  wire s_csamul_cla32_fa7_16_or0;
  wire s_csamul_cla32_and8_16;
  wire s_csamul_cla32_fa8_16_xor0;
  wire s_csamul_cla32_fa8_16_and0;
  wire s_csamul_cla32_fa8_16_xor1;
  wire s_csamul_cla32_fa8_16_and1;
  wire s_csamul_cla32_fa8_16_or0;
  wire s_csamul_cla32_and9_16;
  wire s_csamul_cla32_fa9_16_xor0;
  wire s_csamul_cla32_fa9_16_and0;
  wire s_csamul_cla32_fa9_16_xor1;
  wire s_csamul_cla32_fa9_16_and1;
  wire s_csamul_cla32_fa9_16_or0;
  wire s_csamul_cla32_and10_16;
  wire s_csamul_cla32_fa10_16_xor0;
  wire s_csamul_cla32_fa10_16_and0;
  wire s_csamul_cla32_fa10_16_xor1;
  wire s_csamul_cla32_fa10_16_and1;
  wire s_csamul_cla32_fa10_16_or0;
  wire s_csamul_cla32_and11_16;
  wire s_csamul_cla32_fa11_16_xor0;
  wire s_csamul_cla32_fa11_16_and0;
  wire s_csamul_cla32_fa11_16_xor1;
  wire s_csamul_cla32_fa11_16_and1;
  wire s_csamul_cla32_fa11_16_or0;
  wire s_csamul_cla32_and12_16;
  wire s_csamul_cla32_fa12_16_xor0;
  wire s_csamul_cla32_fa12_16_and0;
  wire s_csamul_cla32_fa12_16_xor1;
  wire s_csamul_cla32_fa12_16_and1;
  wire s_csamul_cla32_fa12_16_or0;
  wire s_csamul_cla32_and13_16;
  wire s_csamul_cla32_fa13_16_xor0;
  wire s_csamul_cla32_fa13_16_and0;
  wire s_csamul_cla32_fa13_16_xor1;
  wire s_csamul_cla32_fa13_16_and1;
  wire s_csamul_cla32_fa13_16_or0;
  wire s_csamul_cla32_and14_16;
  wire s_csamul_cla32_fa14_16_xor0;
  wire s_csamul_cla32_fa14_16_and0;
  wire s_csamul_cla32_fa14_16_xor1;
  wire s_csamul_cla32_fa14_16_and1;
  wire s_csamul_cla32_fa14_16_or0;
  wire s_csamul_cla32_and15_16;
  wire s_csamul_cla32_fa15_16_xor0;
  wire s_csamul_cla32_fa15_16_and0;
  wire s_csamul_cla32_fa15_16_xor1;
  wire s_csamul_cla32_fa15_16_and1;
  wire s_csamul_cla32_fa15_16_or0;
  wire s_csamul_cla32_and16_16;
  wire s_csamul_cla32_fa16_16_xor0;
  wire s_csamul_cla32_fa16_16_and0;
  wire s_csamul_cla32_fa16_16_xor1;
  wire s_csamul_cla32_fa16_16_and1;
  wire s_csamul_cla32_fa16_16_or0;
  wire s_csamul_cla32_and17_16;
  wire s_csamul_cla32_fa17_16_xor0;
  wire s_csamul_cla32_fa17_16_and0;
  wire s_csamul_cla32_fa17_16_xor1;
  wire s_csamul_cla32_fa17_16_and1;
  wire s_csamul_cla32_fa17_16_or0;
  wire s_csamul_cla32_and18_16;
  wire s_csamul_cla32_fa18_16_xor0;
  wire s_csamul_cla32_fa18_16_and0;
  wire s_csamul_cla32_fa18_16_xor1;
  wire s_csamul_cla32_fa18_16_and1;
  wire s_csamul_cla32_fa18_16_or0;
  wire s_csamul_cla32_and19_16;
  wire s_csamul_cla32_fa19_16_xor0;
  wire s_csamul_cla32_fa19_16_and0;
  wire s_csamul_cla32_fa19_16_xor1;
  wire s_csamul_cla32_fa19_16_and1;
  wire s_csamul_cla32_fa19_16_or0;
  wire s_csamul_cla32_and20_16;
  wire s_csamul_cla32_fa20_16_xor0;
  wire s_csamul_cla32_fa20_16_and0;
  wire s_csamul_cla32_fa20_16_xor1;
  wire s_csamul_cla32_fa20_16_and1;
  wire s_csamul_cla32_fa20_16_or0;
  wire s_csamul_cla32_and21_16;
  wire s_csamul_cla32_fa21_16_xor0;
  wire s_csamul_cla32_fa21_16_and0;
  wire s_csamul_cla32_fa21_16_xor1;
  wire s_csamul_cla32_fa21_16_and1;
  wire s_csamul_cla32_fa21_16_or0;
  wire s_csamul_cla32_and22_16;
  wire s_csamul_cla32_fa22_16_xor0;
  wire s_csamul_cla32_fa22_16_and0;
  wire s_csamul_cla32_fa22_16_xor1;
  wire s_csamul_cla32_fa22_16_and1;
  wire s_csamul_cla32_fa22_16_or0;
  wire s_csamul_cla32_and23_16;
  wire s_csamul_cla32_fa23_16_xor0;
  wire s_csamul_cla32_fa23_16_and0;
  wire s_csamul_cla32_fa23_16_xor1;
  wire s_csamul_cla32_fa23_16_and1;
  wire s_csamul_cla32_fa23_16_or0;
  wire s_csamul_cla32_and24_16;
  wire s_csamul_cla32_fa24_16_xor0;
  wire s_csamul_cla32_fa24_16_and0;
  wire s_csamul_cla32_fa24_16_xor1;
  wire s_csamul_cla32_fa24_16_and1;
  wire s_csamul_cla32_fa24_16_or0;
  wire s_csamul_cla32_and25_16;
  wire s_csamul_cla32_fa25_16_xor0;
  wire s_csamul_cla32_fa25_16_and0;
  wire s_csamul_cla32_fa25_16_xor1;
  wire s_csamul_cla32_fa25_16_and1;
  wire s_csamul_cla32_fa25_16_or0;
  wire s_csamul_cla32_and26_16;
  wire s_csamul_cla32_fa26_16_xor0;
  wire s_csamul_cla32_fa26_16_and0;
  wire s_csamul_cla32_fa26_16_xor1;
  wire s_csamul_cla32_fa26_16_and1;
  wire s_csamul_cla32_fa26_16_or0;
  wire s_csamul_cla32_and27_16;
  wire s_csamul_cla32_fa27_16_xor0;
  wire s_csamul_cla32_fa27_16_and0;
  wire s_csamul_cla32_fa27_16_xor1;
  wire s_csamul_cla32_fa27_16_and1;
  wire s_csamul_cla32_fa27_16_or0;
  wire s_csamul_cla32_and28_16;
  wire s_csamul_cla32_fa28_16_xor0;
  wire s_csamul_cla32_fa28_16_and0;
  wire s_csamul_cla32_fa28_16_xor1;
  wire s_csamul_cla32_fa28_16_and1;
  wire s_csamul_cla32_fa28_16_or0;
  wire s_csamul_cla32_and29_16;
  wire s_csamul_cla32_fa29_16_xor0;
  wire s_csamul_cla32_fa29_16_and0;
  wire s_csamul_cla32_fa29_16_xor1;
  wire s_csamul_cla32_fa29_16_and1;
  wire s_csamul_cla32_fa29_16_or0;
  wire s_csamul_cla32_and30_16;
  wire s_csamul_cla32_fa30_16_xor0;
  wire s_csamul_cla32_fa30_16_and0;
  wire s_csamul_cla32_fa30_16_xor1;
  wire s_csamul_cla32_fa30_16_and1;
  wire s_csamul_cla32_fa30_16_or0;
  wire s_csamul_cla32_nand31_16;
  wire s_csamul_cla32_ha31_16_xor0;
  wire s_csamul_cla32_ha31_16_and0;
  wire s_csamul_cla32_and0_17;
  wire s_csamul_cla32_fa0_17_xor0;
  wire s_csamul_cla32_fa0_17_and0;
  wire s_csamul_cla32_fa0_17_xor1;
  wire s_csamul_cla32_fa0_17_and1;
  wire s_csamul_cla32_fa0_17_or0;
  wire s_csamul_cla32_and1_17;
  wire s_csamul_cla32_fa1_17_xor0;
  wire s_csamul_cla32_fa1_17_and0;
  wire s_csamul_cla32_fa1_17_xor1;
  wire s_csamul_cla32_fa1_17_and1;
  wire s_csamul_cla32_fa1_17_or0;
  wire s_csamul_cla32_and2_17;
  wire s_csamul_cla32_fa2_17_xor0;
  wire s_csamul_cla32_fa2_17_and0;
  wire s_csamul_cla32_fa2_17_xor1;
  wire s_csamul_cla32_fa2_17_and1;
  wire s_csamul_cla32_fa2_17_or0;
  wire s_csamul_cla32_and3_17;
  wire s_csamul_cla32_fa3_17_xor0;
  wire s_csamul_cla32_fa3_17_and0;
  wire s_csamul_cla32_fa3_17_xor1;
  wire s_csamul_cla32_fa3_17_and1;
  wire s_csamul_cla32_fa3_17_or0;
  wire s_csamul_cla32_and4_17;
  wire s_csamul_cla32_fa4_17_xor0;
  wire s_csamul_cla32_fa4_17_and0;
  wire s_csamul_cla32_fa4_17_xor1;
  wire s_csamul_cla32_fa4_17_and1;
  wire s_csamul_cla32_fa4_17_or0;
  wire s_csamul_cla32_and5_17;
  wire s_csamul_cla32_fa5_17_xor0;
  wire s_csamul_cla32_fa5_17_and0;
  wire s_csamul_cla32_fa5_17_xor1;
  wire s_csamul_cla32_fa5_17_and1;
  wire s_csamul_cla32_fa5_17_or0;
  wire s_csamul_cla32_and6_17;
  wire s_csamul_cla32_fa6_17_xor0;
  wire s_csamul_cla32_fa6_17_and0;
  wire s_csamul_cla32_fa6_17_xor1;
  wire s_csamul_cla32_fa6_17_and1;
  wire s_csamul_cla32_fa6_17_or0;
  wire s_csamul_cla32_and7_17;
  wire s_csamul_cla32_fa7_17_xor0;
  wire s_csamul_cla32_fa7_17_and0;
  wire s_csamul_cla32_fa7_17_xor1;
  wire s_csamul_cla32_fa7_17_and1;
  wire s_csamul_cla32_fa7_17_or0;
  wire s_csamul_cla32_and8_17;
  wire s_csamul_cla32_fa8_17_xor0;
  wire s_csamul_cla32_fa8_17_and0;
  wire s_csamul_cla32_fa8_17_xor1;
  wire s_csamul_cla32_fa8_17_and1;
  wire s_csamul_cla32_fa8_17_or0;
  wire s_csamul_cla32_and9_17;
  wire s_csamul_cla32_fa9_17_xor0;
  wire s_csamul_cla32_fa9_17_and0;
  wire s_csamul_cla32_fa9_17_xor1;
  wire s_csamul_cla32_fa9_17_and1;
  wire s_csamul_cla32_fa9_17_or0;
  wire s_csamul_cla32_and10_17;
  wire s_csamul_cla32_fa10_17_xor0;
  wire s_csamul_cla32_fa10_17_and0;
  wire s_csamul_cla32_fa10_17_xor1;
  wire s_csamul_cla32_fa10_17_and1;
  wire s_csamul_cla32_fa10_17_or0;
  wire s_csamul_cla32_and11_17;
  wire s_csamul_cla32_fa11_17_xor0;
  wire s_csamul_cla32_fa11_17_and0;
  wire s_csamul_cla32_fa11_17_xor1;
  wire s_csamul_cla32_fa11_17_and1;
  wire s_csamul_cla32_fa11_17_or0;
  wire s_csamul_cla32_and12_17;
  wire s_csamul_cla32_fa12_17_xor0;
  wire s_csamul_cla32_fa12_17_and0;
  wire s_csamul_cla32_fa12_17_xor1;
  wire s_csamul_cla32_fa12_17_and1;
  wire s_csamul_cla32_fa12_17_or0;
  wire s_csamul_cla32_and13_17;
  wire s_csamul_cla32_fa13_17_xor0;
  wire s_csamul_cla32_fa13_17_and0;
  wire s_csamul_cla32_fa13_17_xor1;
  wire s_csamul_cla32_fa13_17_and1;
  wire s_csamul_cla32_fa13_17_or0;
  wire s_csamul_cla32_and14_17;
  wire s_csamul_cla32_fa14_17_xor0;
  wire s_csamul_cla32_fa14_17_and0;
  wire s_csamul_cla32_fa14_17_xor1;
  wire s_csamul_cla32_fa14_17_and1;
  wire s_csamul_cla32_fa14_17_or0;
  wire s_csamul_cla32_and15_17;
  wire s_csamul_cla32_fa15_17_xor0;
  wire s_csamul_cla32_fa15_17_and0;
  wire s_csamul_cla32_fa15_17_xor1;
  wire s_csamul_cla32_fa15_17_and1;
  wire s_csamul_cla32_fa15_17_or0;
  wire s_csamul_cla32_and16_17;
  wire s_csamul_cla32_fa16_17_xor0;
  wire s_csamul_cla32_fa16_17_and0;
  wire s_csamul_cla32_fa16_17_xor1;
  wire s_csamul_cla32_fa16_17_and1;
  wire s_csamul_cla32_fa16_17_or0;
  wire s_csamul_cla32_and17_17;
  wire s_csamul_cla32_fa17_17_xor0;
  wire s_csamul_cla32_fa17_17_and0;
  wire s_csamul_cla32_fa17_17_xor1;
  wire s_csamul_cla32_fa17_17_and1;
  wire s_csamul_cla32_fa17_17_or0;
  wire s_csamul_cla32_and18_17;
  wire s_csamul_cla32_fa18_17_xor0;
  wire s_csamul_cla32_fa18_17_and0;
  wire s_csamul_cla32_fa18_17_xor1;
  wire s_csamul_cla32_fa18_17_and1;
  wire s_csamul_cla32_fa18_17_or0;
  wire s_csamul_cla32_and19_17;
  wire s_csamul_cla32_fa19_17_xor0;
  wire s_csamul_cla32_fa19_17_and0;
  wire s_csamul_cla32_fa19_17_xor1;
  wire s_csamul_cla32_fa19_17_and1;
  wire s_csamul_cla32_fa19_17_or0;
  wire s_csamul_cla32_and20_17;
  wire s_csamul_cla32_fa20_17_xor0;
  wire s_csamul_cla32_fa20_17_and0;
  wire s_csamul_cla32_fa20_17_xor1;
  wire s_csamul_cla32_fa20_17_and1;
  wire s_csamul_cla32_fa20_17_or0;
  wire s_csamul_cla32_and21_17;
  wire s_csamul_cla32_fa21_17_xor0;
  wire s_csamul_cla32_fa21_17_and0;
  wire s_csamul_cla32_fa21_17_xor1;
  wire s_csamul_cla32_fa21_17_and1;
  wire s_csamul_cla32_fa21_17_or0;
  wire s_csamul_cla32_and22_17;
  wire s_csamul_cla32_fa22_17_xor0;
  wire s_csamul_cla32_fa22_17_and0;
  wire s_csamul_cla32_fa22_17_xor1;
  wire s_csamul_cla32_fa22_17_and1;
  wire s_csamul_cla32_fa22_17_or0;
  wire s_csamul_cla32_and23_17;
  wire s_csamul_cla32_fa23_17_xor0;
  wire s_csamul_cla32_fa23_17_and0;
  wire s_csamul_cla32_fa23_17_xor1;
  wire s_csamul_cla32_fa23_17_and1;
  wire s_csamul_cla32_fa23_17_or0;
  wire s_csamul_cla32_and24_17;
  wire s_csamul_cla32_fa24_17_xor0;
  wire s_csamul_cla32_fa24_17_and0;
  wire s_csamul_cla32_fa24_17_xor1;
  wire s_csamul_cla32_fa24_17_and1;
  wire s_csamul_cla32_fa24_17_or0;
  wire s_csamul_cla32_and25_17;
  wire s_csamul_cla32_fa25_17_xor0;
  wire s_csamul_cla32_fa25_17_and0;
  wire s_csamul_cla32_fa25_17_xor1;
  wire s_csamul_cla32_fa25_17_and1;
  wire s_csamul_cla32_fa25_17_or0;
  wire s_csamul_cla32_and26_17;
  wire s_csamul_cla32_fa26_17_xor0;
  wire s_csamul_cla32_fa26_17_and0;
  wire s_csamul_cla32_fa26_17_xor1;
  wire s_csamul_cla32_fa26_17_and1;
  wire s_csamul_cla32_fa26_17_or0;
  wire s_csamul_cla32_and27_17;
  wire s_csamul_cla32_fa27_17_xor0;
  wire s_csamul_cla32_fa27_17_and0;
  wire s_csamul_cla32_fa27_17_xor1;
  wire s_csamul_cla32_fa27_17_and1;
  wire s_csamul_cla32_fa27_17_or0;
  wire s_csamul_cla32_and28_17;
  wire s_csamul_cla32_fa28_17_xor0;
  wire s_csamul_cla32_fa28_17_and0;
  wire s_csamul_cla32_fa28_17_xor1;
  wire s_csamul_cla32_fa28_17_and1;
  wire s_csamul_cla32_fa28_17_or0;
  wire s_csamul_cla32_and29_17;
  wire s_csamul_cla32_fa29_17_xor0;
  wire s_csamul_cla32_fa29_17_and0;
  wire s_csamul_cla32_fa29_17_xor1;
  wire s_csamul_cla32_fa29_17_and1;
  wire s_csamul_cla32_fa29_17_or0;
  wire s_csamul_cla32_and30_17;
  wire s_csamul_cla32_fa30_17_xor0;
  wire s_csamul_cla32_fa30_17_and0;
  wire s_csamul_cla32_fa30_17_xor1;
  wire s_csamul_cla32_fa30_17_and1;
  wire s_csamul_cla32_fa30_17_or0;
  wire s_csamul_cla32_nand31_17;
  wire s_csamul_cla32_ha31_17_xor0;
  wire s_csamul_cla32_ha31_17_and0;
  wire s_csamul_cla32_and0_18;
  wire s_csamul_cla32_fa0_18_xor0;
  wire s_csamul_cla32_fa0_18_and0;
  wire s_csamul_cla32_fa0_18_xor1;
  wire s_csamul_cla32_fa0_18_and1;
  wire s_csamul_cla32_fa0_18_or0;
  wire s_csamul_cla32_and1_18;
  wire s_csamul_cla32_fa1_18_xor0;
  wire s_csamul_cla32_fa1_18_and0;
  wire s_csamul_cla32_fa1_18_xor1;
  wire s_csamul_cla32_fa1_18_and1;
  wire s_csamul_cla32_fa1_18_or0;
  wire s_csamul_cla32_and2_18;
  wire s_csamul_cla32_fa2_18_xor0;
  wire s_csamul_cla32_fa2_18_and0;
  wire s_csamul_cla32_fa2_18_xor1;
  wire s_csamul_cla32_fa2_18_and1;
  wire s_csamul_cla32_fa2_18_or0;
  wire s_csamul_cla32_and3_18;
  wire s_csamul_cla32_fa3_18_xor0;
  wire s_csamul_cla32_fa3_18_and0;
  wire s_csamul_cla32_fa3_18_xor1;
  wire s_csamul_cla32_fa3_18_and1;
  wire s_csamul_cla32_fa3_18_or0;
  wire s_csamul_cla32_and4_18;
  wire s_csamul_cla32_fa4_18_xor0;
  wire s_csamul_cla32_fa4_18_and0;
  wire s_csamul_cla32_fa4_18_xor1;
  wire s_csamul_cla32_fa4_18_and1;
  wire s_csamul_cla32_fa4_18_or0;
  wire s_csamul_cla32_and5_18;
  wire s_csamul_cla32_fa5_18_xor0;
  wire s_csamul_cla32_fa5_18_and0;
  wire s_csamul_cla32_fa5_18_xor1;
  wire s_csamul_cla32_fa5_18_and1;
  wire s_csamul_cla32_fa5_18_or0;
  wire s_csamul_cla32_and6_18;
  wire s_csamul_cla32_fa6_18_xor0;
  wire s_csamul_cla32_fa6_18_and0;
  wire s_csamul_cla32_fa6_18_xor1;
  wire s_csamul_cla32_fa6_18_and1;
  wire s_csamul_cla32_fa6_18_or0;
  wire s_csamul_cla32_and7_18;
  wire s_csamul_cla32_fa7_18_xor0;
  wire s_csamul_cla32_fa7_18_and0;
  wire s_csamul_cla32_fa7_18_xor1;
  wire s_csamul_cla32_fa7_18_and1;
  wire s_csamul_cla32_fa7_18_or0;
  wire s_csamul_cla32_and8_18;
  wire s_csamul_cla32_fa8_18_xor0;
  wire s_csamul_cla32_fa8_18_and0;
  wire s_csamul_cla32_fa8_18_xor1;
  wire s_csamul_cla32_fa8_18_and1;
  wire s_csamul_cla32_fa8_18_or0;
  wire s_csamul_cla32_and9_18;
  wire s_csamul_cla32_fa9_18_xor0;
  wire s_csamul_cla32_fa9_18_and0;
  wire s_csamul_cla32_fa9_18_xor1;
  wire s_csamul_cla32_fa9_18_and1;
  wire s_csamul_cla32_fa9_18_or0;
  wire s_csamul_cla32_and10_18;
  wire s_csamul_cla32_fa10_18_xor0;
  wire s_csamul_cla32_fa10_18_and0;
  wire s_csamul_cla32_fa10_18_xor1;
  wire s_csamul_cla32_fa10_18_and1;
  wire s_csamul_cla32_fa10_18_or0;
  wire s_csamul_cla32_and11_18;
  wire s_csamul_cla32_fa11_18_xor0;
  wire s_csamul_cla32_fa11_18_and0;
  wire s_csamul_cla32_fa11_18_xor1;
  wire s_csamul_cla32_fa11_18_and1;
  wire s_csamul_cla32_fa11_18_or0;
  wire s_csamul_cla32_and12_18;
  wire s_csamul_cla32_fa12_18_xor0;
  wire s_csamul_cla32_fa12_18_and0;
  wire s_csamul_cla32_fa12_18_xor1;
  wire s_csamul_cla32_fa12_18_and1;
  wire s_csamul_cla32_fa12_18_or0;
  wire s_csamul_cla32_and13_18;
  wire s_csamul_cla32_fa13_18_xor0;
  wire s_csamul_cla32_fa13_18_and0;
  wire s_csamul_cla32_fa13_18_xor1;
  wire s_csamul_cla32_fa13_18_and1;
  wire s_csamul_cla32_fa13_18_or0;
  wire s_csamul_cla32_and14_18;
  wire s_csamul_cla32_fa14_18_xor0;
  wire s_csamul_cla32_fa14_18_and0;
  wire s_csamul_cla32_fa14_18_xor1;
  wire s_csamul_cla32_fa14_18_and1;
  wire s_csamul_cla32_fa14_18_or0;
  wire s_csamul_cla32_and15_18;
  wire s_csamul_cla32_fa15_18_xor0;
  wire s_csamul_cla32_fa15_18_and0;
  wire s_csamul_cla32_fa15_18_xor1;
  wire s_csamul_cla32_fa15_18_and1;
  wire s_csamul_cla32_fa15_18_or0;
  wire s_csamul_cla32_and16_18;
  wire s_csamul_cla32_fa16_18_xor0;
  wire s_csamul_cla32_fa16_18_and0;
  wire s_csamul_cla32_fa16_18_xor1;
  wire s_csamul_cla32_fa16_18_and1;
  wire s_csamul_cla32_fa16_18_or0;
  wire s_csamul_cla32_and17_18;
  wire s_csamul_cla32_fa17_18_xor0;
  wire s_csamul_cla32_fa17_18_and0;
  wire s_csamul_cla32_fa17_18_xor1;
  wire s_csamul_cla32_fa17_18_and1;
  wire s_csamul_cla32_fa17_18_or0;
  wire s_csamul_cla32_and18_18;
  wire s_csamul_cla32_fa18_18_xor0;
  wire s_csamul_cla32_fa18_18_and0;
  wire s_csamul_cla32_fa18_18_xor1;
  wire s_csamul_cla32_fa18_18_and1;
  wire s_csamul_cla32_fa18_18_or0;
  wire s_csamul_cla32_and19_18;
  wire s_csamul_cla32_fa19_18_xor0;
  wire s_csamul_cla32_fa19_18_and0;
  wire s_csamul_cla32_fa19_18_xor1;
  wire s_csamul_cla32_fa19_18_and1;
  wire s_csamul_cla32_fa19_18_or0;
  wire s_csamul_cla32_and20_18;
  wire s_csamul_cla32_fa20_18_xor0;
  wire s_csamul_cla32_fa20_18_and0;
  wire s_csamul_cla32_fa20_18_xor1;
  wire s_csamul_cla32_fa20_18_and1;
  wire s_csamul_cla32_fa20_18_or0;
  wire s_csamul_cla32_and21_18;
  wire s_csamul_cla32_fa21_18_xor0;
  wire s_csamul_cla32_fa21_18_and0;
  wire s_csamul_cla32_fa21_18_xor1;
  wire s_csamul_cla32_fa21_18_and1;
  wire s_csamul_cla32_fa21_18_or0;
  wire s_csamul_cla32_and22_18;
  wire s_csamul_cla32_fa22_18_xor0;
  wire s_csamul_cla32_fa22_18_and0;
  wire s_csamul_cla32_fa22_18_xor1;
  wire s_csamul_cla32_fa22_18_and1;
  wire s_csamul_cla32_fa22_18_or0;
  wire s_csamul_cla32_and23_18;
  wire s_csamul_cla32_fa23_18_xor0;
  wire s_csamul_cla32_fa23_18_and0;
  wire s_csamul_cla32_fa23_18_xor1;
  wire s_csamul_cla32_fa23_18_and1;
  wire s_csamul_cla32_fa23_18_or0;
  wire s_csamul_cla32_and24_18;
  wire s_csamul_cla32_fa24_18_xor0;
  wire s_csamul_cla32_fa24_18_and0;
  wire s_csamul_cla32_fa24_18_xor1;
  wire s_csamul_cla32_fa24_18_and1;
  wire s_csamul_cla32_fa24_18_or0;
  wire s_csamul_cla32_and25_18;
  wire s_csamul_cla32_fa25_18_xor0;
  wire s_csamul_cla32_fa25_18_and0;
  wire s_csamul_cla32_fa25_18_xor1;
  wire s_csamul_cla32_fa25_18_and1;
  wire s_csamul_cla32_fa25_18_or0;
  wire s_csamul_cla32_and26_18;
  wire s_csamul_cla32_fa26_18_xor0;
  wire s_csamul_cla32_fa26_18_and0;
  wire s_csamul_cla32_fa26_18_xor1;
  wire s_csamul_cla32_fa26_18_and1;
  wire s_csamul_cla32_fa26_18_or0;
  wire s_csamul_cla32_and27_18;
  wire s_csamul_cla32_fa27_18_xor0;
  wire s_csamul_cla32_fa27_18_and0;
  wire s_csamul_cla32_fa27_18_xor1;
  wire s_csamul_cla32_fa27_18_and1;
  wire s_csamul_cla32_fa27_18_or0;
  wire s_csamul_cla32_and28_18;
  wire s_csamul_cla32_fa28_18_xor0;
  wire s_csamul_cla32_fa28_18_and0;
  wire s_csamul_cla32_fa28_18_xor1;
  wire s_csamul_cla32_fa28_18_and1;
  wire s_csamul_cla32_fa28_18_or0;
  wire s_csamul_cla32_and29_18;
  wire s_csamul_cla32_fa29_18_xor0;
  wire s_csamul_cla32_fa29_18_and0;
  wire s_csamul_cla32_fa29_18_xor1;
  wire s_csamul_cla32_fa29_18_and1;
  wire s_csamul_cla32_fa29_18_or0;
  wire s_csamul_cla32_and30_18;
  wire s_csamul_cla32_fa30_18_xor0;
  wire s_csamul_cla32_fa30_18_and0;
  wire s_csamul_cla32_fa30_18_xor1;
  wire s_csamul_cla32_fa30_18_and1;
  wire s_csamul_cla32_fa30_18_or0;
  wire s_csamul_cla32_nand31_18;
  wire s_csamul_cla32_ha31_18_xor0;
  wire s_csamul_cla32_ha31_18_and0;
  wire s_csamul_cla32_and0_19;
  wire s_csamul_cla32_fa0_19_xor0;
  wire s_csamul_cla32_fa0_19_and0;
  wire s_csamul_cla32_fa0_19_xor1;
  wire s_csamul_cla32_fa0_19_and1;
  wire s_csamul_cla32_fa0_19_or0;
  wire s_csamul_cla32_and1_19;
  wire s_csamul_cla32_fa1_19_xor0;
  wire s_csamul_cla32_fa1_19_and0;
  wire s_csamul_cla32_fa1_19_xor1;
  wire s_csamul_cla32_fa1_19_and1;
  wire s_csamul_cla32_fa1_19_or0;
  wire s_csamul_cla32_and2_19;
  wire s_csamul_cla32_fa2_19_xor0;
  wire s_csamul_cla32_fa2_19_and0;
  wire s_csamul_cla32_fa2_19_xor1;
  wire s_csamul_cla32_fa2_19_and1;
  wire s_csamul_cla32_fa2_19_or0;
  wire s_csamul_cla32_and3_19;
  wire s_csamul_cla32_fa3_19_xor0;
  wire s_csamul_cla32_fa3_19_and0;
  wire s_csamul_cla32_fa3_19_xor1;
  wire s_csamul_cla32_fa3_19_and1;
  wire s_csamul_cla32_fa3_19_or0;
  wire s_csamul_cla32_and4_19;
  wire s_csamul_cla32_fa4_19_xor0;
  wire s_csamul_cla32_fa4_19_and0;
  wire s_csamul_cla32_fa4_19_xor1;
  wire s_csamul_cla32_fa4_19_and1;
  wire s_csamul_cla32_fa4_19_or0;
  wire s_csamul_cla32_and5_19;
  wire s_csamul_cla32_fa5_19_xor0;
  wire s_csamul_cla32_fa5_19_and0;
  wire s_csamul_cla32_fa5_19_xor1;
  wire s_csamul_cla32_fa5_19_and1;
  wire s_csamul_cla32_fa5_19_or0;
  wire s_csamul_cla32_and6_19;
  wire s_csamul_cla32_fa6_19_xor0;
  wire s_csamul_cla32_fa6_19_and0;
  wire s_csamul_cla32_fa6_19_xor1;
  wire s_csamul_cla32_fa6_19_and1;
  wire s_csamul_cla32_fa6_19_or0;
  wire s_csamul_cla32_and7_19;
  wire s_csamul_cla32_fa7_19_xor0;
  wire s_csamul_cla32_fa7_19_and0;
  wire s_csamul_cla32_fa7_19_xor1;
  wire s_csamul_cla32_fa7_19_and1;
  wire s_csamul_cla32_fa7_19_or0;
  wire s_csamul_cla32_and8_19;
  wire s_csamul_cla32_fa8_19_xor0;
  wire s_csamul_cla32_fa8_19_and0;
  wire s_csamul_cla32_fa8_19_xor1;
  wire s_csamul_cla32_fa8_19_and1;
  wire s_csamul_cla32_fa8_19_or0;
  wire s_csamul_cla32_and9_19;
  wire s_csamul_cla32_fa9_19_xor0;
  wire s_csamul_cla32_fa9_19_and0;
  wire s_csamul_cla32_fa9_19_xor1;
  wire s_csamul_cla32_fa9_19_and1;
  wire s_csamul_cla32_fa9_19_or0;
  wire s_csamul_cla32_and10_19;
  wire s_csamul_cla32_fa10_19_xor0;
  wire s_csamul_cla32_fa10_19_and0;
  wire s_csamul_cla32_fa10_19_xor1;
  wire s_csamul_cla32_fa10_19_and1;
  wire s_csamul_cla32_fa10_19_or0;
  wire s_csamul_cla32_and11_19;
  wire s_csamul_cla32_fa11_19_xor0;
  wire s_csamul_cla32_fa11_19_and0;
  wire s_csamul_cla32_fa11_19_xor1;
  wire s_csamul_cla32_fa11_19_and1;
  wire s_csamul_cla32_fa11_19_or0;
  wire s_csamul_cla32_and12_19;
  wire s_csamul_cla32_fa12_19_xor0;
  wire s_csamul_cla32_fa12_19_and0;
  wire s_csamul_cla32_fa12_19_xor1;
  wire s_csamul_cla32_fa12_19_and1;
  wire s_csamul_cla32_fa12_19_or0;
  wire s_csamul_cla32_and13_19;
  wire s_csamul_cla32_fa13_19_xor0;
  wire s_csamul_cla32_fa13_19_and0;
  wire s_csamul_cla32_fa13_19_xor1;
  wire s_csamul_cla32_fa13_19_and1;
  wire s_csamul_cla32_fa13_19_or0;
  wire s_csamul_cla32_and14_19;
  wire s_csamul_cla32_fa14_19_xor0;
  wire s_csamul_cla32_fa14_19_and0;
  wire s_csamul_cla32_fa14_19_xor1;
  wire s_csamul_cla32_fa14_19_and1;
  wire s_csamul_cla32_fa14_19_or0;
  wire s_csamul_cla32_and15_19;
  wire s_csamul_cla32_fa15_19_xor0;
  wire s_csamul_cla32_fa15_19_and0;
  wire s_csamul_cla32_fa15_19_xor1;
  wire s_csamul_cla32_fa15_19_and1;
  wire s_csamul_cla32_fa15_19_or0;
  wire s_csamul_cla32_and16_19;
  wire s_csamul_cla32_fa16_19_xor0;
  wire s_csamul_cla32_fa16_19_and0;
  wire s_csamul_cla32_fa16_19_xor1;
  wire s_csamul_cla32_fa16_19_and1;
  wire s_csamul_cla32_fa16_19_or0;
  wire s_csamul_cla32_and17_19;
  wire s_csamul_cla32_fa17_19_xor0;
  wire s_csamul_cla32_fa17_19_and0;
  wire s_csamul_cla32_fa17_19_xor1;
  wire s_csamul_cla32_fa17_19_and1;
  wire s_csamul_cla32_fa17_19_or0;
  wire s_csamul_cla32_and18_19;
  wire s_csamul_cla32_fa18_19_xor0;
  wire s_csamul_cla32_fa18_19_and0;
  wire s_csamul_cla32_fa18_19_xor1;
  wire s_csamul_cla32_fa18_19_and1;
  wire s_csamul_cla32_fa18_19_or0;
  wire s_csamul_cla32_and19_19;
  wire s_csamul_cla32_fa19_19_xor0;
  wire s_csamul_cla32_fa19_19_and0;
  wire s_csamul_cla32_fa19_19_xor1;
  wire s_csamul_cla32_fa19_19_and1;
  wire s_csamul_cla32_fa19_19_or0;
  wire s_csamul_cla32_and20_19;
  wire s_csamul_cla32_fa20_19_xor0;
  wire s_csamul_cla32_fa20_19_and0;
  wire s_csamul_cla32_fa20_19_xor1;
  wire s_csamul_cla32_fa20_19_and1;
  wire s_csamul_cla32_fa20_19_or0;
  wire s_csamul_cla32_and21_19;
  wire s_csamul_cla32_fa21_19_xor0;
  wire s_csamul_cla32_fa21_19_and0;
  wire s_csamul_cla32_fa21_19_xor1;
  wire s_csamul_cla32_fa21_19_and1;
  wire s_csamul_cla32_fa21_19_or0;
  wire s_csamul_cla32_and22_19;
  wire s_csamul_cla32_fa22_19_xor0;
  wire s_csamul_cla32_fa22_19_and0;
  wire s_csamul_cla32_fa22_19_xor1;
  wire s_csamul_cla32_fa22_19_and1;
  wire s_csamul_cla32_fa22_19_or0;
  wire s_csamul_cla32_and23_19;
  wire s_csamul_cla32_fa23_19_xor0;
  wire s_csamul_cla32_fa23_19_and0;
  wire s_csamul_cla32_fa23_19_xor1;
  wire s_csamul_cla32_fa23_19_and1;
  wire s_csamul_cla32_fa23_19_or0;
  wire s_csamul_cla32_and24_19;
  wire s_csamul_cla32_fa24_19_xor0;
  wire s_csamul_cla32_fa24_19_and0;
  wire s_csamul_cla32_fa24_19_xor1;
  wire s_csamul_cla32_fa24_19_and1;
  wire s_csamul_cla32_fa24_19_or0;
  wire s_csamul_cla32_and25_19;
  wire s_csamul_cla32_fa25_19_xor0;
  wire s_csamul_cla32_fa25_19_and0;
  wire s_csamul_cla32_fa25_19_xor1;
  wire s_csamul_cla32_fa25_19_and1;
  wire s_csamul_cla32_fa25_19_or0;
  wire s_csamul_cla32_and26_19;
  wire s_csamul_cla32_fa26_19_xor0;
  wire s_csamul_cla32_fa26_19_and0;
  wire s_csamul_cla32_fa26_19_xor1;
  wire s_csamul_cla32_fa26_19_and1;
  wire s_csamul_cla32_fa26_19_or0;
  wire s_csamul_cla32_and27_19;
  wire s_csamul_cla32_fa27_19_xor0;
  wire s_csamul_cla32_fa27_19_and0;
  wire s_csamul_cla32_fa27_19_xor1;
  wire s_csamul_cla32_fa27_19_and1;
  wire s_csamul_cla32_fa27_19_or0;
  wire s_csamul_cla32_and28_19;
  wire s_csamul_cla32_fa28_19_xor0;
  wire s_csamul_cla32_fa28_19_and0;
  wire s_csamul_cla32_fa28_19_xor1;
  wire s_csamul_cla32_fa28_19_and1;
  wire s_csamul_cla32_fa28_19_or0;
  wire s_csamul_cla32_and29_19;
  wire s_csamul_cla32_fa29_19_xor0;
  wire s_csamul_cla32_fa29_19_and0;
  wire s_csamul_cla32_fa29_19_xor1;
  wire s_csamul_cla32_fa29_19_and1;
  wire s_csamul_cla32_fa29_19_or0;
  wire s_csamul_cla32_and30_19;
  wire s_csamul_cla32_fa30_19_xor0;
  wire s_csamul_cla32_fa30_19_and0;
  wire s_csamul_cla32_fa30_19_xor1;
  wire s_csamul_cla32_fa30_19_and1;
  wire s_csamul_cla32_fa30_19_or0;
  wire s_csamul_cla32_nand31_19;
  wire s_csamul_cla32_ha31_19_xor0;
  wire s_csamul_cla32_ha31_19_and0;
  wire s_csamul_cla32_and0_20;
  wire s_csamul_cla32_fa0_20_xor0;
  wire s_csamul_cla32_fa0_20_and0;
  wire s_csamul_cla32_fa0_20_xor1;
  wire s_csamul_cla32_fa0_20_and1;
  wire s_csamul_cla32_fa0_20_or0;
  wire s_csamul_cla32_and1_20;
  wire s_csamul_cla32_fa1_20_xor0;
  wire s_csamul_cla32_fa1_20_and0;
  wire s_csamul_cla32_fa1_20_xor1;
  wire s_csamul_cla32_fa1_20_and1;
  wire s_csamul_cla32_fa1_20_or0;
  wire s_csamul_cla32_and2_20;
  wire s_csamul_cla32_fa2_20_xor0;
  wire s_csamul_cla32_fa2_20_and0;
  wire s_csamul_cla32_fa2_20_xor1;
  wire s_csamul_cla32_fa2_20_and1;
  wire s_csamul_cla32_fa2_20_or0;
  wire s_csamul_cla32_and3_20;
  wire s_csamul_cla32_fa3_20_xor0;
  wire s_csamul_cla32_fa3_20_and0;
  wire s_csamul_cla32_fa3_20_xor1;
  wire s_csamul_cla32_fa3_20_and1;
  wire s_csamul_cla32_fa3_20_or0;
  wire s_csamul_cla32_and4_20;
  wire s_csamul_cla32_fa4_20_xor0;
  wire s_csamul_cla32_fa4_20_and0;
  wire s_csamul_cla32_fa4_20_xor1;
  wire s_csamul_cla32_fa4_20_and1;
  wire s_csamul_cla32_fa4_20_or0;
  wire s_csamul_cla32_and5_20;
  wire s_csamul_cla32_fa5_20_xor0;
  wire s_csamul_cla32_fa5_20_and0;
  wire s_csamul_cla32_fa5_20_xor1;
  wire s_csamul_cla32_fa5_20_and1;
  wire s_csamul_cla32_fa5_20_or0;
  wire s_csamul_cla32_and6_20;
  wire s_csamul_cla32_fa6_20_xor0;
  wire s_csamul_cla32_fa6_20_and0;
  wire s_csamul_cla32_fa6_20_xor1;
  wire s_csamul_cla32_fa6_20_and1;
  wire s_csamul_cla32_fa6_20_or0;
  wire s_csamul_cla32_and7_20;
  wire s_csamul_cla32_fa7_20_xor0;
  wire s_csamul_cla32_fa7_20_and0;
  wire s_csamul_cla32_fa7_20_xor1;
  wire s_csamul_cla32_fa7_20_and1;
  wire s_csamul_cla32_fa7_20_or0;
  wire s_csamul_cla32_and8_20;
  wire s_csamul_cla32_fa8_20_xor0;
  wire s_csamul_cla32_fa8_20_and0;
  wire s_csamul_cla32_fa8_20_xor1;
  wire s_csamul_cla32_fa8_20_and1;
  wire s_csamul_cla32_fa8_20_or0;
  wire s_csamul_cla32_and9_20;
  wire s_csamul_cla32_fa9_20_xor0;
  wire s_csamul_cla32_fa9_20_and0;
  wire s_csamul_cla32_fa9_20_xor1;
  wire s_csamul_cla32_fa9_20_and1;
  wire s_csamul_cla32_fa9_20_or0;
  wire s_csamul_cla32_and10_20;
  wire s_csamul_cla32_fa10_20_xor0;
  wire s_csamul_cla32_fa10_20_and0;
  wire s_csamul_cla32_fa10_20_xor1;
  wire s_csamul_cla32_fa10_20_and1;
  wire s_csamul_cla32_fa10_20_or0;
  wire s_csamul_cla32_and11_20;
  wire s_csamul_cla32_fa11_20_xor0;
  wire s_csamul_cla32_fa11_20_and0;
  wire s_csamul_cla32_fa11_20_xor1;
  wire s_csamul_cla32_fa11_20_and1;
  wire s_csamul_cla32_fa11_20_or0;
  wire s_csamul_cla32_and12_20;
  wire s_csamul_cla32_fa12_20_xor0;
  wire s_csamul_cla32_fa12_20_and0;
  wire s_csamul_cla32_fa12_20_xor1;
  wire s_csamul_cla32_fa12_20_and1;
  wire s_csamul_cla32_fa12_20_or0;
  wire s_csamul_cla32_and13_20;
  wire s_csamul_cla32_fa13_20_xor0;
  wire s_csamul_cla32_fa13_20_and0;
  wire s_csamul_cla32_fa13_20_xor1;
  wire s_csamul_cla32_fa13_20_and1;
  wire s_csamul_cla32_fa13_20_or0;
  wire s_csamul_cla32_and14_20;
  wire s_csamul_cla32_fa14_20_xor0;
  wire s_csamul_cla32_fa14_20_and0;
  wire s_csamul_cla32_fa14_20_xor1;
  wire s_csamul_cla32_fa14_20_and1;
  wire s_csamul_cla32_fa14_20_or0;
  wire s_csamul_cla32_and15_20;
  wire s_csamul_cla32_fa15_20_xor0;
  wire s_csamul_cla32_fa15_20_and0;
  wire s_csamul_cla32_fa15_20_xor1;
  wire s_csamul_cla32_fa15_20_and1;
  wire s_csamul_cla32_fa15_20_or0;
  wire s_csamul_cla32_and16_20;
  wire s_csamul_cla32_fa16_20_xor0;
  wire s_csamul_cla32_fa16_20_and0;
  wire s_csamul_cla32_fa16_20_xor1;
  wire s_csamul_cla32_fa16_20_and1;
  wire s_csamul_cla32_fa16_20_or0;
  wire s_csamul_cla32_and17_20;
  wire s_csamul_cla32_fa17_20_xor0;
  wire s_csamul_cla32_fa17_20_and0;
  wire s_csamul_cla32_fa17_20_xor1;
  wire s_csamul_cla32_fa17_20_and1;
  wire s_csamul_cla32_fa17_20_or0;
  wire s_csamul_cla32_and18_20;
  wire s_csamul_cla32_fa18_20_xor0;
  wire s_csamul_cla32_fa18_20_and0;
  wire s_csamul_cla32_fa18_20_xor1;
  wire s_csamul_cla32_fa18_20_and1;
  wire s_csamul_cla32_fa18_20_or0;
  wire s_csamul_cla32_and19_20;
  wire s_csamul_cla32_fa19_20_xor0;
  wire s_csamul_cla32_fa19_20_and0;
  wire s_csamul_cla32_fa19_20_xor1;
  wire s_csamul_cla32_fa19_20_and1;
  wire s_csamul_cla32_fa19_20_or0;
  wire s_csamul_cla32_and20_20;
  wire s_csamul_cla32_fa20_20_xor0;
  wire s_csamul_cla32_fa20_20_and0;
  wire s_csamul_cla32_fa20_20_xor1;
  wire s_csamul_cla32_fa20_20_and1;
  wire s_csamul_cla32_fa20_20_or0;
  wire s_csamul_cla32_and21_20;
  wire s_csamul_cla32_fa21_20_xor0;
  wire s_csamul_cla32_fa21_20_and0;
  wire s_csamul_cla32_fa21_20_xor1;
  wire s_csamul_cla32_fa21_20_and1;
  wire s_csamul_cla32_fa21_20_or0;
  wire s_csamul_cla32_and22_20;
  wire s_csamul_cla32_fa22_20_xor0;
  wire s_csamul_cla32_fa22_20_and0;
  wire s_csamul_cla32_fa22_20_xor1;
  wire s_csamul_cla32_fa22_20_and1;
  wire s_csamul_cla32_fa22_20_or0;
  wire s_csamul_cla32_and23_20;
  wire s_csamul_cla32_fa23_20_xor0;
  wire s_csamul_cla32_fa23_20_and0;
  wire s_csamul_cla32_fa23_20_xor1;
  wire s_csamul_cla32_fa23_20_and1;
  wire s_csamul_cla32_fa23_20_or0;
  wire s_csamul_cla32_and24_20;
  wire s_csamul_cla32_fa24_20_xor0;
  wire s_csamul_cla32_fa24_20_and0;
  wire s_csamul_cla32_fa24_20_xor1;
  wire s_csamul_cla32_fa24_20_and1;
  wire s_csamul_cla32_fa24_20_or0;
  wire s_csamul_cla32_and25_20;
  wire s_csamul_cla32_fa25_20_xor0;
  wire s_csamul_cla32_fa25_20_and0;
  wire s_csamul_cla32_fa25_20_xor1;
  wire s_csamul_cla32_fa25_20_and1;
  wire s_csamul_cla32_fa25_20_or0;
  wire s_csamul_cla32_and26_20;
  wire s_csamul_cla32_fa26_20_xor0;
  wire s_csamul_cla32_fa26_20_and0;
  wire s_csamul_cla32_fa26_20_xor1;
  wire s_csamul_cla32_fa26_20_and1;
  wire s_csamul_cla32_fa26_20_or0;
  wire s_csamul_cla32_and27_20;
  wire s_csamul_cla32_fa27_20_xor0;
  wire s_csamul_cla32_fa27_20_and0;
  wire s_csamul_cla32_fa27_20_xor1;
  wire s_csamul_cla32_fa27_20_and1;
  wire s_csamul_cla32_fa27_20_or0;
  wire s_csamul_cla32_and28_20;
  wire s_csamul_cla32_fa28_20_xor0;
  wire s_csamul_cla32_fa28_20_and0;
  wire s_csamul_cla32_fa28_20_xor1;
  wire s_csamul_cla32_fa28_20_and1;
  wire s_csamul_cla32_fa28_20_or0;
  wire s_csamul_cla32_and29_20;
  wire s_csamul_cla32_fa29_20_xor0;
  wire s_csamul_cla32_fa29_20_and0;
  wire s_csamul_cla32_fa29_20_xor1;
  wire s_csamul_cla32_fa29_20_and1;
  wire s_csamul_cla32_fa29_20_or0;
  wire s_csamul_cla32_and30_20;
  wire s_csamul_cla32_fa30_20_xor0;
  wire s_csamul_cla32_fa30_20_and0;
  wire s_csamul_cla32_fa30_20_xor1;
  wire s_csamul_cla32_fa30_20_and1;
  wire s_csamul_cla32_fa30_20_or0;
  wire s_csamul_cla32_nand31_20;
  wire s_csamul_cla32_ha31_20_xor0;
  wire s_csamul_cla32_ha31_20_and0;
  wire s_csamul_cla32_and0_21;
  wire s_csamul_cla32_fa0_21_xor0;
  wire s_csamul_cla32_fa0_21_and0;
  wire s_csamul_cla32_fa0_21_xor1;
  wire s_csamul_cla32_fa0_21_and1;
  wire s_csamul_cla32_fa0_21_or0;
  wire s_csamul_cla32_and1_21;
  wire s_csamul_cla32_fa1_21_xor0;
  wire s_csamul_cla32_fa1_21_and0;
  wire s_csamul_cla32_fa1_21_xor1;
  wire s_csamul_cla32_fa1_21_and1;
  wire s_csamul_cla32_fa1_21_or0;
  wire s_csamul_cla32_and2_21;
  wire s_csamul_cla32_fa2_21_xor0;
  wire s_csamul_cla32_fa2_21_and0;
  wire s_csamul_cla32_fa2_21_xor1;
  wire s_csamul_cla32_fa2_21_and1;
  wire s_csamul_cla32_fa2_21_or0;
  wire s_csamul_cla32_and3_21;
  wire s_csamul_cla32_fa3_21_xor0;
  wire s_csamul_cla32_fa3_21_and0;
  wire s_csamul_cla32_fa3_21_xor1;
  wire s_csamul_cla32_fa3_21_and1;
  wire s_csamul_cla32_fa3_21_or0;
  wire s_csamul_cla32_and4_21;
  wire s_csamul_cla32_fa4_21_xor0;
  wire s_csamul_cla32_fa4_21_and0;
  wire s_csamul_cla32_fa4_21_xor1;
  wire s_csamul_cla32_fa4_21_and1;
  wire s_csamul_cla32_fa4_21_or0;
  wire s_csamul_cla32_and5_21;
  wire s_csamul_cla32_fa5_21_xor0;
  wire s_csamul_cla32_fa5_21_and0;
  wire s_csamul_cla32_fa5_21_xor1;
  wire s_csamul_cla32_fa5_21_and1;
  wire s_csamul_cla32_fa5_21_or0;
  wire s_csamul_cla32_and6_21;
  wire s_csamul_cla32_fa6_21_xor0;
  wire s_csamul_cla32_fa6_21_and0;
  wire s_csamul_cla32_fa6_21_xor1;
  wire s_csamul_cla32_fa6_21_and1;
  wire s_csamul_cla32_fa6_21_or0;
  wire s_csamul_cla32_and7_21;
  wire s_csamul_cla32_fa7_21_xor0;
  wire s_csamul_cla32_fa7_21_and0;
  wire s_csamul_cla32_fa7_21_xor1;
  wire s_csamul_cla32_fa7_21_and1;
  wire s_csamul_cla32_fa7_21_or0;
  wire s_csamul_cla32_and8_21;
  wire s_csamul_cla32_fa8_21_xor0;
  wire s_csamul_cla32_fa8_21_and0;
  wire s_csamul_cla32_fa8_21_xor1;
  wire s_csamul_cla32_fa8_21_and1;
  wire s_csamul_cla32_fa8_21_or0;
  wire s_csamul_cla32_and9_21;
  wire s_csamul_cla32_fa9_21_xor0;
  wire s_csamul_cla32_fa9_21_and0;
  wire s_csamul_cla32_fa9_21_xor1;
  wire s_csamul_cla32_fa9_21_and1;
  wire s_csamul_cla32_fa9_21_or0;
  wire s_csamul_cla32_and10_21;
  wire s_csamul_cla32_fa10_21_xor0;
  wire s_csamul_cla32_fa10_21_and0;
  wire s_csamul_cla32_fa10_21_xor1;
  wire s_csamul_cla32_fa10_21_and1;
  wire s_csamul_cla32_fa10_21_or0;
  wire s_csamul_cla32_and11_21;
  wire s_csamul_cla32_fa11_21_xor0;
  wire s_csamul_cla32_fa11_21_and0;
  wire s_csamul_cla32_fa11_21_xor1;
  wire s_csamul_cla32_fa11_21_and1;
  wire s_csamul_cla32_fa11_21_or0;
  wire s_csamul_cla32_and12_21;
  wire s_csamul_cla32_fa12_21_xor0;
  wire s_csamul_cla32_fa12_21_and0;
  wire s_csamul_cla32_fa12_21_xor1;
  wire s_csamul_cla32_fa12_21_and1;
  wire s_csamul_cla32_fa12_21_or0;
  wire s_csamul_cla32_and13_21;
  wire s_csamul_cla32_fa13_21_xor0;
  wire s_csamul_cla32_fa13_21_and0;
  wire s_csamul_cla32_fa13_21_xor1;
  wire s_csamul_cla32_fa13_21_and1;
  wire s_csamul_cla32_fa13_21_or0;
  wire s_csamul_cla32_and14_21;
  wire s_csamul_cla32_fa14_21_xor0;
  wire s_csamul_cla32_fa14_21_and0;
  wire s_csamul_cla32_fa14_21_xor1;
  wire s_csamul_cla32_fa14_21_and1;
  wire s_csamul_cla32_fa14_21_or0;
  wire s_csamul_cla32_and15_21;
  wire s_csamul_cla32_fa15_21_xor0;
  wire s_csamul_cla32_fa15_21_and0;
  wire s_csamul_cla32_fa15_21_xor1;
  wire s_csamul_cla32_fa15_21_and1;
  wire s_csamul_cla32_fa15_21_or0;
  wire s_csamul_cla32_and16_21;
  wire s_csamul_cla32_fa16_21_xor0;
  wire s_csamul_cla32_fa16_21_and0;
  wire s_csamul_cla32_fa16_21_xor1;
  wire s_csamul_cla32_fa16_21_and1;
  wire s_csamul_cla32_fa16_21_or0;
  wire s_csamul_cla32_and17_21;
  wire s_csamul_cla32_fa17_21_xor0;
  wire s_csamul_cla32_fa17_21_and0;
  wire s_csamul_cla32_fa17_21_xor1;
  wire s_csamul_cla32_fa17_21_and1;
  wire s_csamul_cla32_fa17_21_or0;
  wire s_csamul_cla32_and18_21;
  wire s_csamul_cla32_fa18_21_xor0;
  wire s_csamul_cla32_fa18_21_and0;
  wire s_csamul_cla32_fa18_21_xor1;
  wire s_csamul_cla32_fa18_21_and1;
  wire s_csamul_cla32_fa18_21_or0;
  wire s_csamul_cla32_and19_21;
  wire s_csamul_cla32_fa19_21_xor0;
  wire s_csamul_cla32_fa19_21_and0;
  wire s_csamul_cla32_fa19_21_xor1;
  wire s_csamul_cla32_fa19_21_and1;
  wire s_csamul_cla32_fa19_21_or0;
  wire s_csamul_cla32_and20_21;
  wire s_csamul_cla32_fa20_21_xor0;
  wire s_csamul_cla32_fa20_21_and0;
  wire s_csamul_cla32_fa20_21_xor1;
  wire s_csamul_cla32_fa20_21_and1;
  wire s_csamul_cla32_fa20_21_or0;
  wire s_csamul_cla32_and21_21;
  wire s_csamul_cla32_fa21_21_xor0;
  wire s_csamul_cla32_fa21_21_and0;
  wire s_csamul_cla32_fa21_21_xor1;
  wire s_csamul_cla32_fa21_21_and1;
  wire s_csamul_cla32_fa21_21_or0;
  wire s_csamul_cla32_and22_21;
  wire s_csamul_cla32_fa22_21_xor0;
  wire s_csamul_cla32_fa22_21_and0;
  wire s_csamul_cla32_fa22_21_xor1;
  wire s_csamul_cla32_fa22_21_and1;
  wire s_csamul_cla32_fa22_21_or0;
  wire s_csamul_cla32_and23_21;
  wire s_csamul_cla32_fa23_21_xor0;
  wire s_csamul_cla32_fa23_21_and0;
  wire s_csamul_cla32_fa23_21_xor1;
  wire s_csamul_cla32_fa23_21_and1;
  wire s_csamul_cla32_fa23_21_or0;
  wire s_csamul_cla32_and24_21;
  wire s_csamul_cla32_fa24_21_xor0;
  wire s_csamul_cla32_fa24_21_and0;
  wire s_csamul_cla32_fa24_21_xor1;
  wire s_csamul_cla32_fa24_21_and1;
  wire s_csamul_cla32_fa24_21_or0;
  wire s_csamul_cla32_and25_21;
  wire s_csamul_cla32_fa25_21_xor0;
  wire s_csamul_cla32_fa25_21_and0;
  wire s_csamul_cla32_fa25_21_xor1;
  wire s_csamul_cla32_fa25_21_and1;
  wire s_csamul_cla32_fa25_21_or0;
  wire s_csamul_cla32_and26_21;
  wire s_csamul_cla32_fa26_21_xor0;
  wire s_csamul_cla32_fa26_21_and0;
  wire s_csamul_cla32_fa26_21_xor1;
  wire s_csamul_cla32_fa26_21_and1;
  wire s_csamul_cla32_fa26_21_or0;
  wire s_csamul_cla32_and27_21;
  wire s_csamul_cla32_fa27_21_xor0;
  wire s_csamul_cla32_fa27_21_and0;
  wire s_csamul_cla32_fa27_21_xor1;
  wire s_csamul_cla32_fa27_21_and1;
  wire s_csamul_cla32_fa27_21_or0;
  wire s_csamul_cla32_and28_21;
  wire s_csamul_cla32_fa28_21_xor0;
  wire s_csamul_cla32_fa28_21_and0;
  wire s_csamul_cla32_fa28_21_xor1;
  wire s_csamul_cla32_fa28_21_and1;
  wire s_csamul_cla32_fa28_21_or0;
  wire s_csamul_cla32_and29_21;
  wire s_csamul_cla32_fa29_21_xor0;
  wire s_csamul_cla32_fa29_21_and0;
  wire s_csamul_cla32_fa29_21_xor1;
  wire s_csamul_cla32_fa29_21_and1;
  wire s_csamul_cla32_fa29_21_or0;
  wire s_csamul_cla32_and30_21;
  wire s_csamul_cla32_fa30_21_xor0;
  wire s_csamul_cla32_fa30_21_and0;
  wire s_csamul_cla32_fa30_21_xor1;
  wire s_csamul_cla32_fa30_21_and1;
  wire s_csamul_cla32_fa30_21_or0;
  wire s_csamul_cla32_nand31_21;
  wire s_csamul_cla32_ha31_21_xor0;
  wire s_csamul_cla32_ha31_21_and0;
  wire s_csamul_cla32_and0_22;
  wire s_csamul_cla32_fa0_22_xor0;
  wire s_csamul_cla32_fa0_22_and0;
  wire s_csamul_cla32_fa0_22_xor1;
  wire s_csamul_cla32_fa0_22_and1;
  wire s_csamul_cla32_fa0_22_or0;
  wire s_csamul_cla32_and1_22;
  wire s_csamul_cla32_fa1_22_xor0;
  wire s_csamul_cla32_fa1_22_and0;
  wire s_csamul_cla32_fa1_22_xor1;
  wire s_csamul_cla32_fa1_22_and1;
  wire s_csamul_cla32_fa1_22_or0;
  wire s_csamul_cla32_and2_22;
  wire s_csamul_cla32_fa2_22_xor0;
  wire s_csamul_cla32_fa2_22_and0;
  wire s_csamul_cla32_fa2_22_xor1;
  wire s_csamul_cla32_fa2_22_and1;
  wire s_csamul_cla32_fa2_22_or0;
  wire s_csamul_cla32_and3_22;
  wire s_csamul_cla32_fa3_22_xor0;
  wire s_csamul_cla32_fa3_22_and0;
  wire s_csamul_cla32_fa3_22_xor1;
  wire s_csamul_cla32_fa3_22_and1;
  wire s_csamul_cla32_fa3_22_or0;
  wire s_csamul_cla32_and4_22;
  wire s_csamul_cla32_fa4_22_xor0;
  wire s_csamul_cla32_fa4_22_and0;
  wire s_csamul_cla32_fa4_22_xor1;
  wire s_csamul_cla32_fa4_22_and1;
  wire s_csamul_cla32_fa4_22_or0;
  wire s_csamul_cla32_and5_22;
  wire s_csamul_cla32_fa5_22_xor0;
  wire s_csamul_cla32_fa5_22_and0;
  wire s_csamul_cla32_fa5_22_xor1;
  wire s_csamul_cla32_fa5_22_and1;
  wire s_csamul_cla32_fa5_22_or0;
  wire s_csamul_cla32_and6_22;
  wire s_csamul_cla32_fa6_22_xor0;
  wire s_csamul_cla32_fa6_22_and0;
  wire s_csamul_cla32_fa6_22_xor1;
  wire s_csamul_cla32_fa6_22_and1;
  wire s_csamul_cla32_fa6_22_or0;
  wire s_csamul_cla32_and7_22;
  wire s_csamul_cla32_fa7_22_xor0;
  wire s_csamul_cla32_fa7_22_and0;
  wire s_csamul_cla32_fa7_22_xor1;
  wire s_csamul_cla32_fa7_22_and1;
  wire s_csamul_cla32_fa7_22_or0;
  wire s_csamul_cla32_and8_22;
  wire s_csamul_cla32_fa8_22_xor0;
  wire s_csamul_cla32_fa8_22_and0;
  wire s_csamul_cla32_fa8_22_xor1;
  wire s_csamul_cla32_fa8_22_and1;
  wire s_csamul_cla32_fa8_22_or0;
  wire s_csamul_cla32_and9_22;
  wire s_csamul_cla32_fa9_22_xor0;
  wire s_csamul_cla32_fa9_22_and0;
  wire s_csamul_cla32_fa9_22_xor1;
  wire s_csamul_cla32_fa9_22_and1;
  wire s_csamul_cla32_fa9_22_or0;
  wire s_csamul_cla32_and10_22;
  wire s_csamul_cla32_fa10_22_xor0;
  wire s_csamul_cla32_fa10_22_and0;
  wire s_csamul_cla32_fa10_22_xor1;
  wire s_csamul_cla32_fa10_22_and1;
  wire s_csamul_cla32_fa10_22_or0;
  wire s_csamul_cla32_and11_22;
  wire s_csamul_cla32_fa11_22_xor0;
  wire s_csamul_cla32_fa11_22_and0;
  wire s_csamul_cla32_fa11_22_xor1;
  wire s_csamul_cla32_fa11_22_and1;
  wire s_csamul_cla32_fa11_22_or0;
  wire s_csamul_cla32_and12_22;
  wire s_csamul_cla32_fa12_22_xor0;
  wire s_csamul_cla32_fa12_22_and0;
  wire s_csamul_cla32_fa12_22_xor1;
  wire s_csamul_cla32_fa12_22_and1;
  wire s_csamul_cla32_fa12_22_or0;
  wire s_csamul_cla32_and13_22;
  wire s_csamul_cla32_fa13_22_xor0;
  wire s_csamul_cla32_fa13_22_and0;
  wire s_csamul_cla32_fa13_22_xor1;
  wire s_csamul_cla32_fa13_22_and1;
  wire s_csamul_cla32_fa13_22_or0;
  wire s_csamul_cla32_and14_22;
  wire s_csamul_cla32_fa14_22_xor0;
  wire s_csamul_cla32_fa14_22_and0;
  wire s_csamul_cla32_fa14_22_xor1;
  wire s_csamul_cla32_fa14_22_and1;
  wire s_csamul_cla32_fa14_22_or0;
  wire s_csamul_cla32_and15_22;
  wire s_csamul_cla32_fa15_22_xor0;
  wire s_csamul_cla32_fa15_22_and0;
  wire s_csamul_cla32_fa15_22_xor1;
  wire s_csamul_cla32_fa15_22_and1;
  wire s_csamul_cla32_fa15_22_or0;
  wire s_csamul_cla32_and16_22;
  wire s_csamul_cla32_fa16_22_xor0;
  wire s_csamul_cla32_fa16_22_and0;
  wire s_csamul_cla32_fa16_22_xor1;
  wire s_csamul_cla32_fa16_22_and1;
  wire s_csamul_cla32_fa16_22_or0;
  wire s_csamul_cla32_and17_22;
  wire s_csamul_cla32_fa17_22_xor0;
  wire s_csamul_cla32_fa17_22_and0;
  wire s_csamul_cla32_fa17_22_xor1;
  wire s_csamul_cla32_fa17_22_and1;
  wire s_csamul_cla32_fa17_22_or0;
  wire s_csamul_cla32_and18_22;
  wire s_csamul_cla32_fa18_22_xor0;
  wire s_csamul_cla32_fa18_22_and0;
  wire s_csamul_cla32_fa18_22_xor1;
  wire s_csamul_cla32_fa18_22_and1;
  wire s_csamul_cla32_fa18_22_or0;
  wire s_csamul_cla32_and19_22;
  wire s_csamul_cla32_fa19_22_xor0;
  wire s_csamul_cla32_fa19_22_and0;
  wire s_csamul_cla32_fa19_22_xor1;
  wire s_csamul_cla32_fa19_22_and1;
  wire s_csamul_cla32_fa19_22_or0;
  wire s_csamul_cla32_and20_22;
  wire s_csamul_cla32_fa20_22_xor0;
  wire s_csamul_cla32_fa20_22_and0;
  wire s_csamul_cla32_fa20_22_xor1;
  wire s_csamul_cla32_fa20_22_and1;
  wire s_csamul_cla32_fa20_22_or0;
  wire s_csamul_cla32_and21_22;
  wire s_csamul_cla32_fa21_22_xor0;
  wire s_csamul_cla32_fa21_22_and0;
  wire s_csamul_cla32_fa21_22_xor1;
  wire s_csamul_cla32_fa21_22_and1;
  wire s_csamul_cla32_fa21_22_or0;
  wire s_csamul_cla32_and22_22;
  wire s_csamul_cla32_fa22_22_xor0;
  wire s_csamul_cla32_fa22_22_and0;
  wire s_csamul_cla32_fa22_22_xor1;
  wire s_csamul_cla32_fa22_22_and1;
  wire s_csamul_cla32_fa22_22_or0;
  wire s_csamul_cla32_and23_22;
  wire s_csamul_cla32_fa23_22_xor0;
  wire s_csamul_cla32_fa23_22_and0;
  wire s_csamul_cla32_fa23_22_xor1;
  wire s_csamul_cla32_fa23_22_and1;
  wire s_csamul_cla32_fa23_22_or0;
  wire s_csamul_cla32_and24_22;
  wire s_csamul_cla32_fa24_22_xor0;
  wire s_csamul_cla32_fa24_22_and0;
  wire s_csamul_cla32_fa24_22_xor1;
  wire s_csamul_cla32_fa24_22_and1;
  wire s_csamul_cla32_fa24_22_or0;
  wire s_csamul_cla32_and25_22;
  wire s_csamul_cla32_fa25_22_xor0;
  wire s_csamul_cla32_fa25_22_and0;
  wire s_csamul_cla32_fa25_22_xor1;
  wire s_csamul_cla32_fa25_22_and1;
  wire s_csamul_cla32_fa25_22_or0;
  wire s_csamul_cla32_and26_22;
  wire s_csamul_cla32_fa26_22_xor0;
  wire s_csamul_cla32_fa26_22_and0;
  wire s_csamul_cla32_fa26_22_xor1;
  wire s_csamul_cla32_fa26_22_and1;
  wire s_csamul_cla32_fa26_22_or0;
  wire s_csamul_cla32_and27_22;
  wire s_csamul_cla32_fa27_22_xor0;
  wire s_csamul_cla32_fa27_22_and0;
  wire s_csamul_cla32_fa27_22_xor1;
  wire s_csamul_cla32_fa27_22_and1;
  wire s_csamul_cla32_fa27_22_or0;
  wire s_csamul_cla32_and28_22;
  wire s_csamul_cla32_fa28_22_xor0;
  wire s_csamul_cla32_fa28_22_and0;
  wire s_csamul_cla32_fa28_22_xor1;
  wire s_csamul_cla32_fa28_22_and1;
  wire s_csamul_cla32_fa28_22_or0;
  wire s_csamul_cla32_and29_22;
  wire s_csamul_cla32_fa29_22_xor0;
  wire s_csamul_cla32_fa29_22_and0;
  wire s_csamul_cla32_fa29_22_xor1;
  wire s_csamul_cla32_fa29_22_and1;
  wire s_csamul_cla32_fa29_22_or0;
  wire s_csamul_cla32_and30_22;
  wire s_csamul_cla32_fa30_22_xor0;
  wire s_csamul_cla32_fa30_22_and0;
  wire s_csamul_cla32_fa30_22_xor1;
  wire s_csamul_cla32_fa30_22_and1;
  wire s_csamul_cla32_fa30_22_or0;
  wire s_csamul_cla32_nand31_22;
  wire s_csamul_cla32_ha31_22_xor0;
  wire s_csamul_cla32_ha31_22_and0;
  wire s_csamul_cla32_and0_23;
  wire s_csamul_cla32_fa0_23_xor0;
  wire s_csamul_cla32_fa0_23_and0;
  wire s_csamul_cla32_fa0_23_xor1;
  wire s_csamul_cla32_fa0_23_and1;
  wire s_csamul_cla32_fa0_23_or0;
  wire s_csamul_cla32_and1_23;
  wire s_csamul_cla32_fa1_23_xor0;
  wire s_csamul_cla32_fa1_23_and0;
  wire s_csamul_cla32_fa1_23_xor1;
  wire s_csamul_cla32_fa1_23_and1;
  wire s_csamul_cla32_fa1_23_or0;
  wire s_csamul_cla32_and2_23;
  wire s_csamul_cla32_fa2_23_xor0;
  wire s_csamul_cla32_fa2_23_and0;
  wire s_csamul_cla32_fa2_23_xor1;
  wire s_csamul_cla32_fa2_23_and1;
  wire s_csamul_cla32_fa2_23_or0;
  wire s_csamul_cla32_and3_23;
  wire s_csamul_cla32_fa3_23_xor0;
  wire s_csamul_cla32_fa3_23_and0;
  wire s_csamul_cla32_fa3_23_xor1;
  wire s_csamul_cla32_fa3_23_and1;
  wire s_csamul_cla32_fa3_23_or0;
  wire s_csamul_cla32_and4_23;
  wire s_csamul_cla32_fa4_23_xor0;
  wire s_csamul_cla32_fa4_23_and0;
  wire s_csamul_cla32_fa4_23_xor1;
  wire s_csamul_cla32_fa4_23_and1;
  wire s_csamul_cla32_fa4_23_or0;
  wire s_csamul_cla32_and5_23;
  wire s_csamul_cla32_fa5_23_xor0;
  wire s_csamul_cla32_fa5_23_and0;
  wire s_csamul_cla32_fa5_23_xor1;
  wire s_csamul_cla32_fa5_23_and1;
  wire s_csamul_cla32_fa5_23_or0;
  wire s_csamul_cla32_and6_23;
  wire s_csamul_cla32_fa6_23_xor0;
  wire s_csamul_cla32_fa6_23_and0;
  wire s_csamul_cla32_fa6_23_xor1;
  wire s_csamul_cla32_fa6_23_and1;
  wire s_csamul_cla32_fa6_23_or0;
  wire s_csamul_cla32_and7_23;
  wire s_csamul_cla32_fa7_23_xor0;
  wire s_csamul_cla32_fa7_23_and0;
  wire s_csamul_cla32_fa7_23_xor1;
  wire s_csamul_cla32_fa7_23_and1;
  wire s_csamul_cla32_fa7_23_or0;
  wire s_csamul_cla32_and8_23;
  wire s_csamul_cla32_fa8_23_xor0;
  wire s_csamul_cla32_fa8_23_and0;
  wire s_csamul_cla32_fa8_23_xor1;
  wire s_csamul_cla32_fa8_23_and1;
  wire s_csamul_cla32_fa8_23_or0;
  wire s_csamul_cla32_and9_23;
  wire s_csamul_cla32_fa9_23_xor0;
  wire s_csamul_cla32_fa9_23_and0;
  wire s_csamul_cla32_fa9_23_xor1;
  wire s_csamul_cla32_fa9_23_and1;
  wire s_csamul_cla32_fa9_23_or0;
  wire s_csamul_cla32_and10_23;
  wire s_csamul_cla32_fa10_23_xor0;
  wire s_csamul_cla32_fa10_23_and0;
  wire s_csamul_cla32_fa10_23_xor1;
  wire s_csamul_cla32_fa10_23_and1;
  wire s_csamul_cla32_fa10_23_or0;
  wire s_csamul_cla32_and11_23;
  wire s_csamul_cla32_fa11_23_xor0;
  wire s_csamul_cla32_fa11_23_and0;
  wire s_csamul_cla32_fa11_23_xor1;
  wire s_csamul_cla32_fa11_23_and1;
  wire s_csamul_cla32_fa11_23_or0;
  wire s_csamul_cla32_and12_23;
  wire s_csamul_cla32_fa12_23_xor0;
  wire s_csamul_cla32_fa12_23_and0;
  wire s_csamul_cla32_fa12_23_xor1;
  wire s_csamul_cla32_fa12_23_and1;
  wire s_csamul_cla32_fa12_23_or0;
  wire s_csamul_cla32_and13_23;
  wire s_csamul_cla32_fa13_23_xor0;
  wire s_csamul_cla32_fa13_23_and0;
  wire s_csamul_cla32_fa13_23_xor1;
  wire s_csamul_cla32_fa13_23_and1;
  wire s_csamul_cla32_fa13_23_or0;
  wire s_csamul_cla32_and14_23;
  wire s_csamul_cla32_fa14_23_xor0;
  wire s_csamul_cla32_fa14_23_and0;
  wire s_csamul_cla32_fa14_23_xor1;
  wire s_csamul_cla32_fa14_23_and1;
  wire s_csamul_cla32_fa14_23_or0;
  wire s_csamul_cla32_and15_23;
  wire s_csamul_cla32_fa15_23_xor0;
  wire s_csamul_cla32_fa15_23_and0;
  wire s_csamul_cla32_fa15_23_xor1;
  wire s_csamul_cla32_fa15_23_and1;
  wire s_csamul_cla32_fa15_23_or0;
  wire s_csamul_cla32_and16_23;
  wire s_csamul_cla32_fa16_23_xor0;
  wire s_csamul_cla32_fa16_23_and0;
  wire s_csamul_cla32_fa16_23_xor1;
  wire s_csamul_cla32_fa16_23_and1;
  wire s_csamul_cla32_fa16_23_or0;
  wire s_csamul_cla32_and17_23;
  wire s_csamul_cla32_fa17_23_xor0;
  wire s_csamul_cla32_fa17_23_and0;
  wire s_csamul_cla32_fa17_23_xor1;
  wire s_csamul_cla32_fa17_23_and1;
  wire s_csamul_cla32_fa17_23_or0;
  wire s_csamul_cla32_and18_23;
  wire s_csamul_cla32_fa18_23_xor0;
  wire s_csamul_cla32_fa18_23_and0;
  wire s_csamul_cla32_fa18_23_xor1;
  wire s_csamul_cla32_fa18_23_and1;
  wire s_csamul_cla32_fa18_23_or0;
  wire s_csamul_cla32_and19_23;
  wire s_csamul_cla32_fa19_23_xor0;
  wire s_csamul_cla32_fa19_23_and0;
  wire s_csamul_cla32_fa19_23_xor1;
  wire s_csamul_cla32_fa19_23_and1;
  wire s_csamul_cla32_fa19_23_or0;
  wire s_csamul_cla32_and20_23;
  wire s_csamul_cla32_fa20_23_xor0;
  wire s_csamul_cla32_fa20_23_and0;
  wire s_csamul_cla32_fa20_23_xor1;
  wire s_csamul_cla32_fa20_23_and1;
  wire s_csamul_cla32_fa20_23_or0;
  wire s_csamul_cla32_and21_23;
  wire s_csamul_cla32_fa21_23_xor0;
  wire s_csamul_cla32_fa21_23_and0;
  wire s_csamul_cla32_fa21_23_xor1;
  wire s_csamul_cla32_fa21_23_and1;
  wire s_csamul_cla32_fa21_23_or0;
  wire s_csamul_cla32_and22_23;
  wire s_csamul_cla32_fa22_23_xor0;
  wire s_csamul_cla32_fa22_23_and0;
  wire s_csamul_cla32_fa22_23_xor1;
  wire s_csamul_cla32_fa22_23_and1;
  wire s_csamul_cla32_fa22_23_or0;
  wire s_csamul_cla32_and23_23;
  wire s_csamul_cla32_fa23_23_xor0;
  wire s_csamul_cla32_fa23_23_and0;
  wire s_csamul_cla32_fa23_23_xor1;
  wire s_csamul_cla32_fa23_23_and1;
  wire s_csamul_cla32_fa23_23_or0;
  wire s_csamul_cla32_and24_23;
  wire s_csamul_cla32_fa24_23_xor0;
  wire s_csamul_cla32_fa24_23_and0;
  wire s_csamul_cla32_fa24_23_xor1;
  wire s_csamul_cla32_fa24_23_and1;
  wire s_csamul_cla32_fa24_23_or0;
  wire s_csamul_cla32_and25_23;
  wire s_csamul_cla32_fa25_23_xor0;
  wire s_csamul_cla32_fa25_23_and0;
  wire s_csamul_cla32_fa25_23_xor1;
  wire s_csamul_cla32_fa25_23_and1;
  wire s_csamul_cla32_fa25_23_or0;
  wire s_csamul_cla32_and26_23;
  wire s_csamul_cla32_fa26_23_xor0;
  wire s_csamul_cla32_fa26_23_and0;
  wire s_csamul_cla32_fa26_23_xor1;
  wire s_csamul_cla32_fa26_23_and1;
  wire s_csamul_cla32_fa26_23_or0;
  wire s_csamul_cla32_and27_23;
  wire s_csamul_cla32_fa27_23_xor0;
  wire s_csamul_cla32_fa27_23_and0;
  wire s_csamul_cla32_fa27_23_xor1;
  wire s_csamul_cla32_fa27_23_and1;
  wire s_csamul_cla32_fa27_23_or0;
  wire s_csamul_cla32_and28_23;
  wire s_csamul_cla32_fa28_23_xor0;
  wire s_csamul_cla32_fa28_23_and0;
  wire s_csamul_cla32_fa28_23_xor1;
  wire s_csamul_cla32_fa28_23_and1;
  wire s_csamul_cla32_fa28_23_or0;
  wire s_csamul_cla32_and29_23;
  wire s_csamul_cla32_fa29_23_xor0;
  wire s_csamul_cla32_fa29_23_and0;
  wire s_csamul_cla32_fa29_23_xor1;
  wire s_csamul_cla32_fa29_23_and1;
  wire s_csamul_cla32_fa29_23_or0;
  wire s_csamul_cla32_and30_23;
  wire s_csamul_cla32_fa30_23_xor0;
  wire s_csamul_cla32_fa30_23_and0;
  wire s_csamul_cla32_fa30_23_xor1;
  wire s_csamul_cla32_fa30_23_and1;
  wire s_csamul_cla32_fa30_23_or0;
  wire s_csamul_cla32_nand31_23;
  wire s_csamul_cla32_ha31_23_xor0;
  wire s_csamul_cla32_ha31_23_and0;
  wire s_csamul_cla32_and0_24;
  wire s_csamul_cla32_fa0_24_xor0;
  wire s_csamul_cla32_fa0_24_and0;
  wire s_csamul_cla32_fa0_24_xor1;
  wire s_csamul_cla32_fa0_24_and1;
  wire s_csamul_cla32_fa0_24_or0;
  wire s_csamul_cla32_and1_24;
  wire s_csamul_cla32_fa1_24_xor0;
  wire s_csamul_cla32_fa1_24_and0;
  wire s_csamul_cla32_fa1_24_xor1;
  wire s_csamul_cla32_fa1_24_and1;
  wire s_csamul_cla32_fa1_24_or0;
  wire s_csamul_cla32_and2_24;
  wire s_csamul_cla32_fa2_24_xor0;
  wire s_csamul_cla32_fa2_24_and0;
  wire s_csamul_cla32_fa2_24_xor1;
  wire s_csamul_cla32_fa2_24_and1;
  wire s_csamul_cla32_fa2_24_or0;
  wire s_csamul_cla32_and3_24;
  wire s_csamul_cla32_fa3_24_xor0;
  wire s_csamul_cla32_fa3_24_and0;
  wire s_csamul_cla32_fa3_24_xor1;
  wire s_csamul_cla32_fa3_24_and1;
  wire s_csamul_cla32_fa3_24_or0;
  wire s_csamul_cla32_and4_24;
  wire s_csamul_cla32_fa4_24_xor0;
  wire s_csamul_cla32_fa4_24_and0;
  wire s_csamul_cla32_fa4_24_xor1;
  wire s_csamul_cla32_fa4_24_and1;
  wire s_csamul_cla32_fa4_24_or0;
  wire s_csamul_cla32_and5_24;
  wire s_csamul_cla32_fa5_24_xor0;
  wire s_csamul_cla32_fa5_24_and0;
  wire s_csamul_cla32_fa5_24_xor1;
  wire s_csamul_cla32_fa5_24_and1;
  wire s_csamul_cla32_fa5_24_or0;
  wire s_csamul_cla32_and6_24;
  wire s_csamul_cla32_fa6_24_xor0;
  wire s_csamul_cla32_fa6_24_and0;
  wire s_csamul_cla32_fa6_24_xor1;
  wire s_csamul_cla32_fa6_24_and1;
  wire s_csamul_cla32_fa6_24_or0;
  wire s_csamul_cla32_and7_24;
  wire s_csamul_cla32_fa7_24_xor0;
  wire s_csamul_cla32_fa7_24_and0;
  wire s_csamul_cla32_fa7_24_xor1;
  wire s_csamul_cla32_fa7_24_and1;
  wire s_csamul_cla32_fa7_24_or0;
  wire s_csamul_cla32_and8_24;
  wire s_csamul_cla32_fa8_24_xor0;
  wire s_csamul_cla32_fa8_24_and0;
  wire s_csamul_cla32_fa8_24_xor1;
  wire s_csamul_cla32_fa8_24_and1;
  wire s_csamul_cla32_fa8_24_or0;
  wire s_csamul_cla32_and9_24;
  wire s_csamul_cla32_fa9_24_xor0;
  wire s_csamul_cla32_fa9_24_and0;
  wire s_csamul_cla32_fa9_24_xor1;
  wire s_csamul_cla32_fa9_24_and1;
  wire s_csamul_cla32_fa9_24_or0;
  wire s_csamul_cla32_and10_24;
  wire s_csamul_cla32_fa10_24_xor0;
  wire s_csamul_cla32_fa10_24_and0;
  wire s_csamul_cla32_fa10_24_xor1;
  wire s_csamul_cla32_fa10_24_and1;
  wire s_csamul_cla32_fa10_24_or0;
  wire s_csamul_cla32_and11_24;
  wire s_csamul_cla32_fa11_24_xor0;
  wire s_csamul_cla32_fa11_24_and0;
  wire s_csamul_cla32_fa11_24_xor1;
  wire s_csamul_cla32_fa11_24_and1;
  wire s_csamul_cla32_fa11_24_or0;
  wire s_csamul_cla32_and12_24;
  wire s_csamul_cla32_fa12_24_xor0;
  wire s_csamul_cla32_fa12_24_and0;
  wire s_csamul_cla32_fa12_24_xor1;
  wire s_csamul_cla32_fa12_24_and1;
  wire s_csamul_cla32_fa12_24_or0;
  wire s_csamul_cla32_and13_24;
  wire s_csamul_cla32_fa13_24_xor0;
  wire s_csamul_cla32_fa13_24_and0;
  wire s_csamul_cla32_fa13_24_xor1;
  wire s_csamul_cla32_fa13_24_and1;
  wire s_csamul_cla32_fa13_24_or0;
  wire s_csamul_cla32_and14_24;
  wire s_csamul_cla32_fa14_24_xor0;
  wire s_csamul_cla32_fa14_24_and0;
  wire s_csamul_cla32_fa14_24_xor1;
  wire s_csamul_cla32_fa14_24_and1;
  wire s_csamul_cla32_fa14_24_or0;
  wire s_csamul_cla32_and15_24;
  wire s_csamul_cla32_fa15_24_xor0;
  wire s_csamul_cla32_fa15_24_and0;
  wire s_csamul_cla32_fa15_24_xor1;
  wire s_csamul_cla32_fa15_24_and1;
  wire s_csamul_cla32_fa15_24_or0;
  wire s_csamul_cla32_and16_24;
  wire s_csamul_cla32_fa16_24_xor0;
  wire s_csamul_cla32_fa16_24_and0;
  wire s_csamul_cla32_fa16_24_xor1;
  wire s_csamul_cla32_fa16_24_and1;
  wire s_csamul_cla32_fa16_24_or0;
  wire s_csamul_cla32_and17_24;
  wire s_csamul_cla32_fa17_24_xor0;
  wire s_csamul_cla32_fa17_24_and0;
  wire s_csamul_cla32_fa17_24_xor1;
  wire s_csamul_cla32_fa17_24_and1;
  wire s_csamul_cla32_fa17_24_or0;
  wire s_csamul_cla32_and18_24;
  wire s_csamul_cla32_fa18_24_xor0;
  wire s_csamul_cla32_fa18_24_and0;
  wire s_csamul_cla32_fa18_24_xor1;
  wire s_csamul_cla32_fa18_24_and1;
  wire s_csamul_cla32_fa18_24_or0;
  wire s_csamul_cla32_and19_24;
  wire s_csamul_cla32_fa19_24_xor0;
  wire s_csamul_cla32_fa19_24_and0;
  wire s_csamul_cla32_fa19_24_xor1;
  wire s_csamul_cla32_fa19_24_and1;
  wire s_csamul_cla32_fa19_24_or0;
  wire s_csamul_cla32_and20_24;
  wire s_csamul_cla32_fa20_24_xor0;
  wire s_csamul_cla32_fa20_24_and0;
  wire s_csamul_cla32_fa20_24_xor1;
  wire s_csamul_cla32_fa20_24_and1;
  wire s_csamul_cla32_fa20_24_or0;
  wire s_csamul_cla32_and21_24;
  wire s_csamul_cla32_fa21_24_xor0;
  wire s_csamul_cla32_fa21_24_and0;
  wire s_csamul_cla32_fa21_24_xor1;
  wire s_csamul_cla32_fa21_24_and1;
  wire s_csamul_cla32_fa21_24_or0;
  wire s_csamul_cla32_and22_24;
  wire s_csamul_cla32_fa22_24_xor0;
  wire s_csamul_cla32_fa22_24_and0;
  wire s_csamul_cla32_fa22_24_xor1;
  wire s_csamul_cla32_fa22_24_and1;
  wire s_csamul_cla32_fa22_24_or0;
  wire s_csamul_cla32_and23_24;
  wire s_csamul_cla32_fa23_24_xor0;
  wire s_csamul_cla32_fa23_24_and0;
  wire s_csamul_cla32_fa23_24_xor1;
  wire s_csamul_cla32_fa23_24_and1;
  wire s_csamul_cla32_fa23_24_or0;
  wire s_csamul_cla32_and24_24;
  wire s_csamul_cla32_fa24_24_xor0;
  wire s_csamul_cla32_fa24_24_and0;
  wire s_csamul_cla32_fa24_24_xor1;
  wire s_csamul_cla32_fa24_24_and1;
  wire s_csamul_cla32_fa24_24_or0;
  wire s_csamul_cla32_and25_24;
  wire s_csamul_cla32_fa25_24_xor0;
  wire s_csamul_cla32_fa25_24_and0;
  wire s_csamul_cla32_fa25_24_xor1;
  wire s_csamul_cla32_fa25_24_and1;
  wire s_csamul_cla32_fa25_24_or0;
  wire s_csamul_cla32_and26_24;
  wire s_csamul_cla32_fa26_24_xor0;
  wire s_csamul_cla32_fa26_24_and0;
  wire s_csamul_cla32_fa26_24_xor1;
  wire s_csamul_cla32_fa26_24_and1;
  wire s_csamul_cla32_fa26_24_or0;
  wire s_csamul_cla32_and27_24;
  wire s_csamul_cla32_fa27_24_xor0;
  wire s_csamul_cla32_fa27_24_and0;
  wire s_csamul_cla32_fa27_24_xor1;
  wire s_csamul_cla32_fa27_24_and1;
  wire s_csamul_cla32_fa27_24_or0;
  wire s_csamul_cla32_and28_24;
  wire s_csamul_cla32_fa28_24_xor0;
  wire s_csamul_cla32_fa28_24_and0;
  wire s_csamul_cla32_fa28_24_xor1;
  wire s_csamul_cla32_fa28_24_and1;
  wire s_csamul_cla32_fa28_24_or0;
  wire s_csamul_cla32_and29_24;
  wire s_csamul_cla32_fa29_24_xor0;
  wire s_csamul_cla32_fa29_24_and0;
  wire s_csamul_cla32_fa29_24_xor1;
  wire s_csamul_cla32_fa29_24_and1;
  wire s_csamul_cla32_fa29_24_or0;
  wire s_csamul_cla32_and30_24;
  wire s_csamul_cla32_fa30_24_xor0;
  wire s_csamul_cla32_fa30_24_and0;
  wire s_csamul_cla32_fa30_24_xor1;
  wire s_csamul_cla32_fa30_24_and1;
  wire s_csamul_cla32_fa30_24_or0;
  wire s_csamul_cla32_nand31_24;
  wire s_csamul_cla32_ha31_24_xor0;
  wire s_csamul_cla32_ha31_24_and0;
  wire s_csamul_cla32_and0_25;
  wire s_csamul_cla32_fa0_25_xor0;
  wire s_csamul_cla32_fa0_25_and0;
  wire s_csamul_cla32_fa0_25_xor1;
  wire s_csamul_cla32_fa0_25_and1;
  wire s_csamul_cla32_fa0_25_or0;
  wire s_csamul_cla32_and1_25;
  wire s_csamul_cla32_fa1_25_xor0;
  wire s_csamul_cla32_fa1_25_and0;
  wire s_csamul_cla32_fa1_25_xor1;
  wire s_csamul_cla32_fa1_25_and1;
  wire s_csamul_cla32_fa1_25_or0;
  wire s_csamul_cla32_and2_25;
  wire s_csamul_cla32_fa2_25_xor0;
  wire s_csamul_cla32_fa2_25_and0;
  wire s_csamul_cla32_fa2_25_xor1;
  wire s_csamul_cla32_fa2_25_and1;
  wire s_csamul_cla32_fa2_25_or0;
  wire s_csamul_cla32_and3_25;
  wire s_csamul_cla32_fa3_25_xor0;
  wire s_csamul_cla32_fa3_25_and0;
  wire s_csamul_cla32_fa3_25_xor1;
  wire s_csamul_cla32_fa3_25_and1;
  wire s_csamul_cla32_fa3_25_or0;
  wire s_csamul_cla32_and4_25;
  wire s_csamul_cla32_fa4_25_xor0;
  wire s_csamul_cla32_fa4_25_and0;
  wire s_csamul_cla32_fa4_25_xor1;
  wire s_csamul_cla32_fa4_25_and1;
  wire s_csamul_cla32_fa4_25_or0;
  wire s_csamul_cla32_and5_25;
  wire s_csamul_cla32_fa5_25_xor0;
  wire s_csamul_cla32_fa5_25_and0;
  wire s_csamul_cla32_fa5_25_xor1;
  wire s_csamul_cla32_fa5_25_and1;
  wire s_csamul_cla32_fa5_25_or0;
  wire s_csamul_cla32_and6_25;
  wire s_csamul_cla32_fa6_25_xor0;
  wire s_csamul_cla32_fa6_25_and0;
  wire s_csamul_cla32_fa6_25_xor1;
  wire s_csamul_cla32_fa6_25_and1;
  wire s_csamul_cla32_fa6_25_or0;
  wire s_csamul_cla32_and7_25;
  wire s_csamul_cla32_fa7_25_xor0;
  wire s_csamul_cla32_fa7_25_and0;
  wire s_csamul_cla32_fa7_25_xor1;
  wire s_csamul_cla32_fa7_25_and1;
  wire s_csamul_cla32_fa7_25_or0;
  wire s_csamul_cla32_and8_25;
  wire s_csamul_cla32_fa8_25_xor0;
  wire s_csamul_cla32_fa8_25_and0;
  wire s_csamul_cla32_fa8_25_xor1;
  wire s_csamul_cla32_fa8_25_and1;
  wire s_csamul_cla32_fa8_25_or0;
  wire s_csamul_cla32_and9_25;
  wire s_csamul_cla32_fa9_25_xor0;
  wire s_csamul_cla32_fa9_25_and0;
  wire s_csamul_cla32_fa9_25_xor1;
  wire s_csamul_cla32_fa9_25_and1;
  wire s_csamul_cla32_fa9_25_or0;
  wire s_csamul_cla32_and10_25;
  wire s_csamul_cla32_fa10_25_xor0;
  wire s_csamul_cla32_fa10_25_and0;
  wire s_csamul_cla32_fa10_25_xor1;
  wire s_csamul_cla32_fa10_25_and1;
  wire s_csamul_cla32_fa10_25_or0;
  wire s_csamul_cla32_and11_25;
  wire s_csamul_cla32_fa11_25_xor0;
  wire s_csamul_cla32_fa11_25_and0;
  wire s_csamul_cla32_fa11_25_xor1;
  wire s_csamul_cla32_fa11_25_and1;
  wire s_csamul_cla32_fa11_25_or0;
  wire s_csamul_cla32_and12_25;
  wire s_csamul_cla32_fa12_25_xor0;
  wire s_csamul_cla32_fa12_25_and0;
  wire s_csamul_cla32_fa12_25_xor1;
  wire s_csamul_cla32_fa12_25_and1;
  wire s_csamul_cla32_fa12_25_or0;
  wire s_csamul_cla32_and13_25;
  wire s_csamul_cla32_fa13_25_xor0;
  wire s_csamul_cla32_fa13_25_and0;
  wire s_csamul_cla32_fa13_25_xor1;
  wire s_csamul_cla32_fa13_25_and1;
  wire s_csamul_cla32_fa13_25_or0;
  wire s_csamul_cla32_and14_25;
  wire s_csamul_cla32_fa14_25_xor0;
  wire s_csamul_cla32_fa14_25_and0;
  wire s_csamul_cla32_fa14_25_xor1;
  wire s_csamul_cla32_fa14_25_and1;
  wire s_csamul_cla32_fa14_25_or0;
  wire s_csamul_cla32_and15_25;
  wire s_csamul_cla32_fa15_25_xor0;
  wire s_csamul_cla32_fa15_25_and0;
  wire s_csamul_cla32_fa15_25_xor1;
  wire s_csamul_cla32_fa15_25_and1;
  wire s_csamul_cla32_fa15_25_or0;
  wire s_csamul_cla32_and16_25;
  wire s_csamul_cla32_fa16_25_xor0;
  wire s_csamul_cla32_fa16_25_and0;
  wire s_csamul_cla32_fa16_25_xor1;
  wire s_csamul_cla32_fa16_25_and1;
  wire s_csamul_cla32_fa16_25_or0;
  wire s_csamul_cla32_and17_25;
  wire s_csamul_cla32_fa17_25_xor0;
  wire s_csamul_cla32_fa17_25_and0;
  wire s_csamul_cla32_fa17_25_xor1;
  wire s_csamul_cla32_fa17_25_and1;
  wire s_csamul_cla32_fa17_25_or0;
  wire s_csamul_cla32_and18_25;
  wire s_csamul_cla32_fa18_25_xor0;
  wire s_csamul_cla32_fa18_25_and0;
  wire s_csamul_cla32_fa18_25_xor1;
  wire s_csamul_cla32_fa18_25_and1;
  wire s_csamul_cla32_fa18_25_or0;
  wire s_csamul_cla32_and19_25;
  wire s_csamul_cla32_fa19_25_xor0;
  wire s_csamul_cla32_fa19_25_and0;
  wire s_csamul_cla32_fa19_25_xor1;
  wire s_csamul_cla32_fa19_25_and1;
  wire s_csamul_cla32_fa19_25_or0;
  wire s_csamul_cla32_and20_25;
  wire s_csamul_cla32_fa20_25_xor0;
  wire s_csamul_cla32_fa20_25_and0;
  wire s_csamul_cla32_fa20_25_xor1;
  wire s_csamul_cla32_fa20_25_and1;
  wire s_csamul_cla32_fa20_25_or0;
  wire s_csamul_cla32_and21_25;
  wire s_csamul_cla32_fa21_25_xor0;
  wire s_csamul_cla32_fa21_25_and0;
  wire s_csamul_cla32_fa21_25_xor1;
  wire s_csamul_cla32_fa21_25_and1;
  wire s_csamul_cla32_fa21_25_or0;
  wire s_csamul_cla32_and22_25;
  wire s_csamul_cla32_fa22_25_xor0;
  wire s_csamul_cla32_fa22_25_and0;
  wire s_csamul_cla32_fa22_25_xor1;
  wire s_csamul_cla32_fa22_25_and1;
  wire s_csamul_cla32_fa22_25_or0;
  wire s_csamul_cla32_and23_25;
  wire s_csamul_cla32_fa23_25_xor0;
  wire s_csamul_cla32_fa23_25_and0;
  wire s_csamul_cla32_fa23_25_xor1;
  wire s_csamul_cla32_fa23_25_and1;
  wire s_csamul_cla32_fa23_25_or0;
  wire s_csamul_cla32_and24_25;
  wire s_csamul_cla32_fa24_25_xor0;
  wire s_csamul_cla32_fa24_25_and0;
  wire s_csamul_cla32_fa24_25_xor1;
  wire s_csamul_cla32_fa24_25_and1;
  wire s_csamul_cla32_fa24_25_or0;
  wire s_csamul_cla32_and25_25;
  wire s_csamul_cla32_fa25_25_xor0;
  wire s_csamul_cla32_fa25_25_and0;
  wire s_csamul_cla32_fa25_25_xor1;
  wire s_csamul_cla32_fa25_25_and1;
  wire s_csamul_cla32_fa25_25_or0;
  wire s_csamul_cla32_and26_25;
  wire s_csamul_cla32_fa26_25_xor0;
  wire s_csamul_cla32_fa26_25_and0;
  wire s_csamul_cla32_fa26_25_xor1;
  wire s_csamul_cla32_fa26_25_and1;
  wire s_csamul_cla32_fa26_25_or0;
  wire s_csamul_cla32_and27_25;
  wire s_csamul_cla32_fa27_25_xor0;
  wire s_csamul_cla32_fa27_25_and0;
  wire s_csamul_cla32_fa27_25_xor1;
  wire s_csamul_cla32_fa27_25_and1;
  wire s_csamul_cla32_fa27_25_or0;
  wire s_csamul_cla32_and28_25;
  wire s_csamul_cla32_fa28_25_xor0;
  wire s_csamul_cla32_fa28_25_and0;
  wire s_csamul_cla32_fa28_25_xor1;
  wire s_csamul_cla32_fa28_25_and1;
  wire s_csamul_cla32_fa28_25_or0;
  wire s_csamul_cla32_and29_25;
  wire s_csamul_cla32_fa29_25_xor0;
  wire s_csamul_cla32_fa29_25_and0;
  wire s_csamul_cla32_fa29_25_xor1;
  wire s_csamul_cla32_fa29_25_and1;
  wire s_csamul_cla32_fa29_25_or0;
  wire s_csamul_cla32_and30_25;
  wire s_csamul_cla32_fa30_25_xor0;
  wire s_csamul_cla32_fa30_25_and0;
  wire s_csamul_cla32_fa30_25_xor1;
  wire s_csamul_cla32_fa30_25_and1;
  wire s_csamul_cla32_fa30_25_or0;
  wire s_csamul_cla32_nand31_25;
  wire s_csamul_cla32_ha31_25_xor0;
  wire s_csamul_cla32_ha31_25_and0;
  wire s_csamul_cla32_and0_26;
  wire s_csamul_cla32_fa0_26_xor0;
  wire s_csamul_cla32_fa0_26_and0;
  wire s_csamul_cla32_fa0_26_xor1;
  wire s_csamul_cla32_fa0_26_and1;
  wire s_csamul_cla32_fa0_26_or0;
  wire s_csamul_cla32_and1_26;
  wire s_csamul_cla32_fa1_26_xor0;
  wire s_csamul_cla32_fa1_26_and0;
  wire s_csamul_cla32_fa1_26_xor1;
  wire s_csamul_cla32_fa1_26_and1;
  wire s_csamul_cla32_fa1_26_or0;
  wire s_csamul_cla32_and2_26;
  wire s_csamul_cla32_fa2_26_xor0;
  wire s_csamul_cla32_fa2_26_and0;
  wire s_csamul_cla32_fa2_26_xor1;
  wire s_csamul_cla32_fa2_26_and1;
  wire s_csamul_cla32_fa2_26_or0;
  wire s_csamul_cla32_and3_26;
  wire s_csamul_cla32_fa3_26_xor0;
  wire s_csamul_cla32_fa3_26_and0;
  wire s_csamul_cla32_fa3_26_xor1;
  wire s_csamul_cla32_fa3_26_and1;
  wire s_csamul_cla32_fa3_26_or0;
  wire s_csamul_cla32_and4_26;
  wire s_csamul_cla32_fa4_26_xor0;
  wire s_csamul_cla32_fa4_26_and0;
  wire s_csamul_cla32_fa4_26_xor1;
  wire s_csamul_cla32_fa4_26_and1;
  wire s_csamul_cla32_fa4_26_or0;
  wire s_csamul_cla32_and5_26;
  wire s_csamul_cla32_fa5_26_xor0;
  wire s_csamul_cla32_fa5_26_and0;
  wire s_csamul_cla32_fa5_26_xor1;
  wire s_csamul_cla32_fa5_26_and1;
  wire s_csamul_cla32_fa5_26_or0;
  wire s_csamul_cla32_and6_26;
  wire s_csamul_cla32_fa6_26_xor0;
  wire s_csamul_cla32_fa6_26_and0;
  wire s_csamul_cla32_fa6_26_xor1;
  wire s_csamul_cla32_fa6_26_and1;
  wire s_csamul_cla32_fa6_26_or0;
  wire s_csamul_cla32_and7_26;
  wire s_csamul_cla32_fa7_26_xor0;
  wire s_csamul_cla32_fa7_26_and0;
  wire s_csamul_cla32_fa7_26_xor1;
  wire s_csamul_cla32_fa7_26_and1;
  wire s_csamul_cla32_fa7_26_or0;
  wire s_csamul_cla32_and8_26;
  wire s_csamul_cla32_fa8_26_xor0;
  wire s_csamul_cla32_fa8_26_and0;
  wire s_csamul_cla32_fa8_26_xor1;
  wire s_csamul_cla32_fa8_26_and1;
  wire s_csamul_cla32_fa8_26_or0;
  wire s_csamul_cla32_and9_26;
  wire s_csamul_cla32_fa9_26_xor0;
  wire s_csamul_cla32_fa9_26_and0;
  wire s_csamul_cla32_fa9_26_xor1;
  wire s_csamul_cla32_fa9_26_and1;
  wire s_csamul_cla32_fa9_26_or0;
  wire s_csamul_cla32_and10_26;
  wire s_csamul_cla32_fa10_26_xor0;
  wire s_csamul_cla32_fa10_26_and0;
  wire s_csamul_cla32_fa10_26_xor1;
  wire s_csamul_cla32_fa10_26_and1;
  wire s_csamul_cla32_fa10_26_or0;
  wire s_csamul_cla32_and11_26;
  wire s_csamul_cla32_fa11_26_xor0;
  wire s_csamul_cla32_fa11_26_and0;
  wire s_csamul_cla32_fa11_26_xor1;
  wire s_csamul_cla32_fa11_26_and1;
  wire s_csamul_cla32_fa11_26_or0;
  wire s_csamul_cla32_and12_26;
  wire s_csamul_cla32_fa12_26_xor0;
  wire s_csamul_cla32_fa12_26_and0;
  wire s_csamul_cla32_fa12_26_xor1;
  wire s_csamul_cla32_fa12_26_and1;
  wire s_csamul_cla32_fa12_26_or0;
  wire s_csamul_cla32_and13_26;
  wire s_csamul_cla32_fa13_26_xor0;
  wire s_csamul_cla32_fa13_26_and0;
  wire s_csamul_cla32_fa13_26_xor1;
  wire s_csamul_cla32_fa13_26_and1;
  wire s_csamul_cla32_fa13_26_or0;
  wire s_csamul_cla32_and14_26;
  wire s_csamul_cla32_fa14_26_xor0;
  wire s_csamul_cla32_fa14_26_and0;
  wire s_csamul_cla32_fa14_26_xor1;
  wire s_csamul_cla32_fa14_26_and1;
  wire s_csamul_cla32_fa14_26_or0;
  wire s_csamul_cla32_and15_26;
  wire s_csamul_cla32_fa15_26_xor0;
  wire s_csamul_cla32_fa15_26_and0;
  wire s_csamul_cla32_fa15_26_xor1;
  wire s_csamul_cla32_fa15_26_and1;
  wire s_csamul_cla32_fa15_26_or0;
  wire s_csamul_cla32_and16_26;
  wire s_csamul_cla32_fa16_26_xor0;
  wire s_csamul_cla32_fa16_26_and0;
  wire s_csamul_cla32_fa16_26_xor1;
  wire s_csamul_cla32_fa16_26_and1;
  wire s_csamul_cla32_fa16_26_or0;
  wire s_csamul_cla32_and17_26;
  wire s_csamul_cla32_fa17_26_xor0;
  wire s_csamul_cla32_fa17_26_and0;
  wire s_csamul_cla32_fa17_26_xor1;
  wire s_csamul_cla32_fa17_26_and1;
  wire s_csamul_cla32_fa17_26_or0;
  wire s_csamul_cla32_and18_26;
  wire s_csamul_cla32_fa18_26_xor0;
  wire s_csamul_cla32_fa18_26_and0;
  wire s_csamul_cla32_fa18_26_xor1;
  wire s_csamul_cla32_fa18_26_and1;
  wire s_csamul_cla32_fa18_26_or0;
  wire s_csamul_cla32_and19_26;
  wire s_csamul_cla32_fa19_26_xor0;
  wire s_csamul_cla32_fa19_26_and0;
  wire s_csamul_cla32_fa19_26_xor1;
  wire s_csamul_cla32_fa19_26_and1;
  wire s_csamul_cla32_fa19_26_or0;
  wire s_csamul_cla32_and20_26;
  wire s_csamul_cla32_fa20_26_xor0;
  wire s_csamul_cla32_fa20_26_and0;
  wire s_csamul_cla32_fa20_26_xor1;
  wire s_csamul_cla32_fa20_26_and1;
  wire s_csamul_cla32_fa20_26_or0;
  wire s_csamul_cla32_and21_26;
  wire s_csamul_cla32_fa21_26_xor0;
  wire s_csamul_cla32_fa21_26_and0;
  wire s_csamul_cla32_fa21_26_xor1;
  wire s_csamul_cla32_fa21_26_and1;
  wire s_csamul_cla32_fa21_26_or0;
  wire s_csamul_cla32_and22_26;
  wire s_csamul_cla32_fa22_26_xor0;
  wire s_csamul_cla32_fa22_26_and0;
  wire s_csamul_cla32_fa22_26_xor1;
  wire s_csamul_cla32_fa22_26_and1;
  wire s_csamul_cla32_fa22_26_or0;
  wire s_csamul_cla32_and23_26;
  wire s_csamul_cla32_fa23_26_xor0;
  wire s_csamul_cla32_fa23_26_and0;
  wire s_csamul_cla32_fa23_26_xor1;
  wire s_csamul_cla32_fa23_26_and1;
  wire s_csamul_cla32_fa23_26_or0;
  wire s_csamul_cla32_and24_26;
  wire s_csamul_cla32_fa24_26_xor0;
  wire s_csamul_cla32_fa24_26_and0;
  wire s_csamul_cla32_fa24_26_xor1;
  wire s_csamul_cla32_fa24_26_and1;
  wire s_csamul_cla32_fa24_26_or0;
  wire s_csamul_cla32_and25_26;
  wire s_csamul_cla32_fa25_26_xor0;
  wire s_csamul_cla32_fa25_26_and0;
  wire s_csamul_cla32_fa25_26_xor1;
  wire s_csamul_cla32_fa25_26_and1;
  wire s_csamul_cla32_fa25_26_or0;
  wire s_csamul_cla32_and26_26;
  wire s_csamul_cla32_fa26_26_xor0;
  wire s_csamul_cla32_fa26_26_and0;
  wire s_csamul_cla32_fa26_26_xor1;
  wire s_csamul_cla32_fa26_26_and1;
  wire s_csamul_cla32_fa26_26_or0;
  wire s_csamul_cla32_and27_26;
  wire s_csamul_cla32_fa27_26_xor0;
  wire s_csamul_cla32_fa27_26_and0;
  wire s_csamul_cla32_fa27_26_xor1;
  wire s_csamul_cla32_fa27_26_and1;
  wire s_csamul_cla32_fa27_26_or0;
  wire s_csamul_cla32_and28_26;
  wire s_csamul_cla32_fa28_26_xor0;
  wire s_csamul_cla32_fa28_26_and0;
  wire s_csamul_cla32_fa28_26_xor1;
  wire s_csamul_cla32_fa28_26_and1;
  wire s_csamul_cla32_fa28_26_or0;
  wire s_csamul_cla32_and29_26;
  wire s_csamul_cla32_fa29_26_xor0;
  wire s_csamul_cla32_fa29_26_and0;
  wire s_csamul_cla32_fa29_26_xor1;
  wire s_csamul_cla32_fa29_26_and1;
  wire s_csamul_cla32_fa29_26_or0;
  wire s_csamul_cla32_and30_26;
  wire s_csamul_cla32_fa30_26_xor0;
  wire s_csamul_cla32_fa30_26_and0;
  wire s_csamul_cla32_fa30_26_xor1;
  wire s_csamul_cla32_fa30_26_and1;
  wire s_csamul_cla32_fa30_26_or0;
  wire s_csamul_cla32_nand31_26;
  wire s_csamul_cla32_ha31_26_xor0;
  wire s_csamul_cla32_ha31_26_and0;
  wire s_csamul_cla32_and0_27;
  wire s_csamul_cla32_fa0_27_xor0;
  wire s_csamul_cla32_fa0_27_and0;
  wire s_csamul_cla32_fa0_27_xor1;
  wire s_csamul_cla32_fa0_27_and1;
  wire s_csamul_cla32_fa0_27_or0;
  wire s_csamul_cla32_and1_27;
  wire s_csamul_cla32_fa1_27_xor0;
  wire s_csamul_cla32_fa1_27_and0;
  wire s_csamul_cla32_fa1_27_xor1;
  wire s_csamul_cla32_fa1_27_and1;
  wire s_csamul_cla32_fa1_27_or0;
  wire s_csamul_cla32_and2_27;
  wire s_csamul_cla32_fa2_27_xor0;
  wire s_csamul_cla32_fa2_27_and0;
  wire s_csamul_cla32_fa2_27_xor1;
  wire s_csamul_cla32_fa2_27_and1;
  wire s_csamul_cla32_fa2_27_or0;
  wire s_csamul_cla32_and3_27;
  wire s_csamul_cla32_fa3_27_xor0;
  wire s_csamul_cla32_fa3_27_and0;
  wire s_csamul_cla32_fa3_27_xor1;
  wire s_csamul_cla32_fa3_27_and1;
  wire s_csamul_cla32_fa3_27_or0;
  wire s_csamul_cla32_and4_27;
  wire s_csamul_cla32_fa4_27_xor0;
  wire s_csamul_cla32_fa4_27_and0;
  wire s_csamul_cla32_fa4_27_xor1;
  wire s_csamul_cla32_fa4_27_and1;
  wire s_csamul_cla32_fa4_27_or0;
  wire s_csamul_cla32_and5_27;
  wire s_csamul_cla32_fa5_27_xor0;
  wire s_csamul_cla32_fa5_27_and0;
  wire s_csamul_cla32_fa5_27_xor1;
  wire s_csamul_cla32_fa5_27_and1;
  wire s_csamul_cla32_fa5_27_or0;
  wire s_csamul_cla32_and6_27;
  wire s_csamul_cla32_fa6_27_xor0;
  wire s_csamul_cla32_fa6_27_and0;
  wire s_csamul_cla32_fa6_27_xor1;
  wire s_csamul_cla32_fa6_27_and1;
  wire s_csamul_cla32_fa6_27_or0;
  wire s_csamul_cla32_and7_27;
  wire s_csamul_cla32_fa7_27_xor0;
  wire s_csamul_cla32_fa7_27_and0;
  wire s_csamul_cla32_fa7_27_xor1;
  wire s_csamul_cla32_fa7_27_and1;
  wire s_csamul_cla32_fa7_27_or0;
  wire s_csamul_cla32_and8_27;
  wire s_csamul_cla32_fa8_27_xor0;
  wire s_csamul_cla32_fa8_27_and0;
  wire s_csamul_cla32_fa8_27_xor1;
  wire s_csamul_cla32_fa8_27_and1;
  wire s_csamul_cla32_fa8_27_or0;
  wire s_csamul_cla32_and9_27;
  wire s_csamul_cla32_fa9_27_xor0;
  wire s_csamul_cla32_fa9_27_and0;
  wire s_csamul_cla32_fa9_27_xor1;
  wire s_csamul_cla32_fa9_27_and1;
  wire s_csamul_cla32_fa9_27_or0;
  wire s_csamul_cla32_and10_27;
  wire s_csamul_cla32_fa10_27_xor0;
  wire s_csamul_cla32_fa10_27_and0;
  wire s_csamul_cla32_fa10_27_xor1;
  wire s_csamul_cla32_fa10_27_and1;
  wire s_csamul_cla32_fa10_27_or0;
  wire s_csamul_cla32_and11_27;
  wire s_csamul_cla32_fa11_27_xor0;
  wire s_csamul_cla32_fa11_27_and0;
  wire s_csamul_cla32_fa11_27_xor1;
  wire s_csamul_cla32_fa11_27_and1;
  wire s_csamul_cla32_fa11_27_or0;
  wire s_csamul_cla32_and12_27;
  wire s_csamul_cla32_fa12_27_xor0;
  wire s_csamul_cla32_fa12_27_and0;
  wire s_csamul_cla32_fa12_27_xor1;
  wire s_csamul_cla32_fa12_27_and1;
  wire s_csamul_cla32_fa12_27_or0;
  wire s_csamul_cla32_and13_27;
  wire s_csamul_cla32_fa13_27_xor0;
  wire s_csamul_cla32_fa13_27_and0;
  wire s_csamul_cla32_fa13_27_xor1;
  wire s_csamul_cla32_fa13_27_and1;
  wire s_csamul_cla32_fa13_27_or0;
  wire s_csamul_cla32_and14_27;
  wire s_csamul_cla32_fa14_27_xor0;
  wire s_csamul_cla32_fa14_27_and0;
  wire s_csamul_cla32_fa14_27_xor1;
  wire s_csamul_cla32_fa14_27_and1;
  wire s_csamul_cla32_fa14_27_or0;
  wire s_csamul_cla32_and15_27;
  wire s_csamul_cla32_fa15_27_xor0;
  wire s_csamul_cla32_fa15_27_and0;
  wire s_csamul_cla32_fa15_27_xor1;
  wire s_csamul_cla32_fa15_27_and1;
  wire s_csamul_cla32_fa15_27_or0;
  wire s_csamul_cla32_and16_27;
  wire s_csamul_cla32_fa16_27_xor0;
  wire s_csamul_cla32_fa16_27_and0;
  wire s_csamul_cla32_fa16_27_xor1;
  wire s_csamul_cla32_fa16_27_and1;
  wire s_csamul_cla32_fa16_27_or0;
  wire s_csamul_cla32_and17_27;
  wire s_csamul_cla32_fa17_27_xor0;
  wire s_csamul_cla32_fa17_27_and0;
  wire s_csamul_cla32_fa17_27_xor1;
  wire s_csamul_cla32_fa17_27_and1;
  wire s_csamul_cla32_fa17_27_or0;
  wire s_csamul_cla32_and18_27;
  wire s_csamul_cla32_fa18_27_xor0;
  wire s_csamul_cla32_fa18_27_and0;
  wire s_csamul_cla32_fa18_27_xor1;
  wire s_csamul_cla32_fa18_27_and1;
  wire s_csamul_cla32_fa18_27_or0;
  wire s_csamul_cla32_and19_27;
  wire s_csamul_cla32_fa19_27_xor0;
  wire s_csamul_cla32_fa19_27_and0;
  wire s_csamul_cla32_fa19_27_xor1;
  wire s_csamul_cla32_fa19_27_and1;
  wire s_csamul_cla32_fa19_27_or0;
  wire s_csamul_cla32_and20_27;
  wire s_csamul_cla32_fa20_27_xor0;
  wire s_csamul_cla32_fa20_27_and0;
  wire s_csamul_cla32_fa20_27_xor1;
  wire s_csamul_cla32_fa20_27_and1;
  wire s_csamul_cla32_fa20_27_or0;
  wire s_csamul_cla32_and21_27;
  wire s_csamul_cla32_fa21_27_xor0;
  wire s_csamul_cla32_fa21_27_and0;
  wire s_csamul_cla32_fa21_27_xor1;
  wire s_csamul_cla32_fa21_27_and1;
  wire s_csamul_cla32_fa21_27_or0;
  wire s_csamul_cla32_and22_27;
  wire s_csamul_cla32_fa22_27_xor0;
  wire s_csamul_cla32_fa22_27_and0;
  wire s_csamul_cla32_fa22_27_xor1;
  wire s_csamul_cla32_fa22_27_and1;
  wire s_csamul_cla32_fa22_27_or0;
  wire s_csamul_cla32_and23_27;
  wire s_csamul_cla32_fa23_27_xor0;
  wire s_csamul_cla32_fa23_27_and0;
  wire s_csamul_cla32_fa23_27_xor1;
  wire s_csamul_cla32_fa23_27_and1;
  wire s_csamul_cla32_fa23_27_or0;
  wire s_csamul_cla32_and24_27;
  wire s_csamul_cla32_fa24_27_xor0;
  wire s_csamul_cla32_fa24_27_and0;
  wire s_csamul_cla32_fa24_27_xor1;
  wire s_csamul_cla32_fa24_27_and1;
  wire s_csamul_cla32_fa24_27_or0;
  wire s_csamul_cla32_and25_27;
  wire s_csamul_cla32_fa25_27_xor0;
  wire s_csamul_cla32_fa25_27_and0;
  wire s_csamul_cla32_fa25_27_xor1;
  wire s_csamul_cla32_fa25_27_and1;
  wire s_csamul_cla32_fa25_27_or0;
  wire s_csamul_cla32_and26_27;
  wire s_csamul_cla32_fa26_27_xor0;
  wire s_csamul_cla32_fa26_27_and0;
  wire s_csamul_cla32_fa26_27_xor1;
  wire s_csamul_cla32_fa26_27_and1;
  wire s_csamul_cla32_fa26_27_or0;
  wire s_csamul_cla32_and27_27;
  wire s_csamul_cla32_fa27_27_xor0;
  wire s_csamul_cla32_fa27_27_and0;
  wire s_csamul_cla32_fa27_27_xor1;
  wire s_csamul_cla32_fa27_27_and1;
  wire s_csamul_cla32_fa27_27_or0;
  wire s_csamul_cla32_and28_27;
  wire s_csamul_cla32_fa28_27_xor0;
  wire s_csamul_cla32_fa28_27_and0;
  wire s_csamul_cla32_fa28_27_xor1;
  wire s_csamul_cla32_fa28_27_and1;
  wire s_csamul_cla32_fa28_27_or0;
  wire s_csamul_cla32_and29_27;
  wire s_csamul_cla32_fa29_27_xor0;
  wire s_csamul_cla32_fa29_27_and0;
  wire s_csamul_cla32_fa29_27_xor1;
  wire s_csamul_cla32_fa29_27_and1;
  wire s_csamul_cla32_fa29_27_or0;
  wire s_csamul_cla32_and30_27;
  wire s_csamul_cla32_fa30_27_xor0;
  wire s_csamul_cla32_fa30_27_and0;
  wire s_csamul_cla32_fa30_27_xor1;
  wire s_csamul_cla32_fa30_27_and1;
  wire s_csamul_cla32_fa30_27_or0;
  wire s_csamul_cla32_nand31_27;
  wire s_csamul_cla32_ha31_27_xor0;
  wire s_csamul_cla32_ha31_27_and0;
  wire s_csamul_cla32_and0_28;
  wire s_csamul_cla32_fa0_28_xor0;
  wire s_csamul_cla32_fa0_28_and0;
  wire s_csamul_cla32_fa0_28_xor1;
  wire s_csamul_cla32_fa0_28_and1;
  wire s_csamul_cla32_fa0_28_or0;
  wire s_csamul_cla32_and1_28;
  wire s_csamul_cla32_fa1_28_xor0;
  wire s_csamul_cla32_fa1_28_and0;
  wire s_csamul_cla32_fa1_28_xor1;
  wire s_csamul_cla32_fa1_28_and1;
  wire s_csamul_cla32_fa1_28_or0;
  wire s_csamul_cla32_and2_28;
  wire s_csamul_cla32_fa2_28_xor0;
  wire s_csamul_cla32_fa2_28_and0;
  wire s_csamul_cla32_fa2_28_xor1;
  wire s_csamul_cla32_fa2_28_and1;
  wire s_csamul_cla32_fa2_28_or0;
  wire s_csamul_cla32_and3_28;
  wire s_csamul_cla32_fa3_28_xor0;
  wire s_csamul_cla32_fa3_28_and0;
  wire s_csamul_cla32_fa3_28_xor1;
  wire s_csamul_cla32_fa3_28_and1;
  wire s_csamul_cla32_fa3_28_or0;
  wire s_csamul_cla32_and4_28;
  wire s_csamul_cla32_fa4_28_xor0;
  wire s_csamul_cla32_fa4_28_and0;
  wire s_csamul_cla32_fa4_28_xor1;
  wire s_csamul_cla32_fa4_28_and1;
  wire s_csamul_cla32_fa4_28_or0;
  wire s_csamul_cla32_and5_28;
  wire s_csamul_cla32_fa5_28_xor0;
  wire s_csamul_cla32_fa5_28_and0;
  wire s_csamul_cla32_fa5_28_xor1;
  wire s_csamul_cla32_fa5_28_and1;
  wire s_csamul_cla32_fa5_28_or0;
  wire s_csamul_cla32_and6_28;
  wire s_csamul_cla32_fa6_28_xor0;
  wire s_csamul_cla32_fa6_28_and0;
  wire s_csamul_cla32_fa6_28_xor1;
  wire s_csamul_cla32_fa6_28_and1;
  wire s_csamul_cla32_fa6_28_or0;
  wire s_csamul_cla32_and7_28;
  wire s_csamul_cla32_fa7_28_xor0;
  wire s_csamul_cla32_fa7_28_and0;
  wire s_csamul_cla32_fa7_28_xor1;
  wire s_csamul_cla32_fa7_28_and1;
  wire s_csamul_cla32_fa7_28_or0;
  wire s_csamul_cla32_and8_28;
  wire s_csamul_cla32_fa8_28_xor0;
  wire s_csamul_cla32_fa8_28_and0;
  wire s_csamul_cla32_fa8_28_xor1;
  wire s_csamul_cla32_fa8_28_and1;
  wire s_csamul_cla32_fa8_28_or0;
  wire s_csamul_cla32_and9_28;
  wire s_csamul_cla32_fa9_28_xor0;
  wire s_csamul_cla32_fa9_28_and0;
  wire s_csamul_cla32_fa9_28_xor1;
  wire s_csamul_cla32_fa9_28_and1;
  wire s_csamul_cla32_fa9_28_or0;
  wire s_csamul_cla32_and10_28;
  wire s_csamul_cla32_fa10_28_xor0;
  wire s_csamul_cla32_fa10_28_and0;
  wire s_csamul_cla32_fa10_28_xor1;
  wire s_csamul_cla32_fa10_28_and1;
  wire s_csamul_cla32_fa10_28_or0;
  wire s_csamul_cla32_and11_28;
  wire s_csamul_cla32_fa11_28_xor0;
  wire s_csamul_cla32_fa11_28_and0;
  wire s_csamul_cla32_fa11_28_xor1;
  wire s_csamul_cla32_fa11_28_and1;
  wire s_csamul_cla32_fa11_28_or0;
  wire s_csamul_cla32_and12_28;
  wire s_csamul_cla32_fa12_28_xor0;
  wire s_csamul_cla32_fa12_28_and0;
  wire s_csamul_cla32_fa12_28_xor1;
  wire s_csamul_cla32_fa12_28_and1;
  wire s_csamul_cla32_fa12_28_or0;
  wire s_csamul_cla32_and13_28;
  wire s_csamul_cla32_fa13_28_xor0;
  wire s_csamul_cla32_fa13_28_and0;
  wire s_csamul_cla32_fa13_28_xor1;
  wire s_csamul_cla32_fa13_28_and1;
  wire s_csamul_cla32_fa13_28_or0;
  wire s_csamul_cla32_and14_28;
  wire s_csamul_cla32_fa14_28_xor0;
  wire s_csamul_cla32_fa14_28_and0;
  wire s_csamul_cla32_fa14_28_xor1;
  wire s_csamul_cla32_fa14_28_and1;
  wire s_csamul_cla32_fa14_28_or0;
  wire s_csamul_cla32_and15_28;
  wire s_csamul_cla32_fa15_28_xor0;
  wire s_csamul_cla32_fa15_28_and0;
  wire s_csamul_cla32_fa15_28_xor1;
  wire s_csamul_cla32_fa15_28_and1;
  wire s_csamul_cla32_fa15_28_or0;
  wire s_csamul_cla32_and16_28;
  wire s_csamul_cla32_fa16_28_xor0;
  wire s_csamul_cla32_fa16_28_and0;
  wire s_csamul_cla32_fa16_28_xor1;
  wire s_csamul_cla32_fa16_28_and1;
  wire s_csamul_cla32_fa16_28_or0;
  wire s_csamul_cla32_and17_28;
  wire s_csamul_cla32_fa17_28_xor0;
  wire s_csamul_cla32_fa17_28_and0;
  wire s_csamul_cla32_fa17_28_xor1;
  wire s_csamul_cla32_fa17_28_and1;
  wire s_csamul_cla32_fa17_28_or0;
  wire s_csamul_cla32_and18_28;
  wire s_csamul_cla32_fa18_28_xor0;
  wire s_csamul_cla32_fa18_28_and0;
  wire s_csamul_cla32_fa18_28_xor1;
  wire s_csamul_cla32_fa18_28_and1;
  wire s_csamul_cla32_fa18_28_or0;
  wire s_csamul_cla32_and19_28;
  wire s_csamul_cla32_fa19_28_xor0;
  wire s_csamul_cla32_fa19_28_and0;
  wire s_csamul_cla32_fa19_28_xor1;
  wire s_csamul_cla32_fa19_28_and1;
  wire s_csamul_cla32_fa19_28_or0;
  wire s_csamul_cla32_and20_28;
  wire s_csamul_cla32_fa20_28_xor0;
  wire s_csamul_cla32_fa20_28_and0;
  wire s_csamul_cla32_fa20_28_xor1;
  wire s_csamul_cla32_fa20_28_and1;
  wire s_csamul_cla32_fa20_28_or0;
  wire s_csamul_cla32_and21_28;
  wire s_csamul_cla32_fa21_28_xor0;
  wire s_csamul_cla32_fa21_28_and0;
  wire s_csamul_cla32_fa21_28_xor1;
  wire s_csamul_cla32_fa21_28_and1;
  wire s_csamul_cla32_fa21_28_or0;
  wire s_csamul_cla32_and22_28;
  wire s_csamul_cla32_fa22_28_xor0;
  wire s_csamul_cla32_fa22_28_and0;
  wire s_csamul_cla32_fa22_28_xor1;
  wire s_csamul_cla32_fa22_28_and1;
  wire s_csamul_cla32_fa22_28_or0;
  wire s_csamul_cla32_and23_28;
  wire s_csamul_cla32_fa23_28_xor0;
  wire s_csamul_cla32_fa23_28_and0;
  wire s_csamul_cla32_fa23_28_xor1;
  wire s_csamul_cla32_fa23_28_and1;
  wire s_csamul_cla32_fa23_28_or0;
  wire s_csamul_cla32_and24_28;
  wire s_csamul_cla32_fa24_28_xor0;
  wire s_csamul_cla32_fa24_28_and0;
  wire s_csamul_cla32_fa24_28_xor1;
  wire s_csamul_cla32_fa24_28_and1;
  wire s_csamul_cla32_fa24_28_or0;
  wire s_csamul_cla32_and25_28;
  wire s_csamul_cla32_fa25_28_xor0;
  wire s_csamul_cla32_fa25_28_and0;
  wire s_csamul_cla32_fa25_28_xor1;
  wire s_csamul_cla32_fa25_28_and1;
  wire s_csamul_cla32_fa25_28_or0;
  wire s_csamul_cla32_and26_28;
  wire s_csamul_cla32_fa26_28_xor0;
  wire s_csamul_cla32_fa26_28_and0;
  wire s_csamul_cla32_fa26_28_xor1;
  wire s_csamul_cla32_fa26_28_and1;
  wire s_csamul_cla32_fa26_28_or0;
  wire s_csamul_cla32_and27_28;
  wire s_csamul_cla32_fa27_28_xor0;
  wire s_csamul_cla32_fa27_28_and0;
  wire s_csamul_cla32_fa27_28_xor1;
  wire s_csamul_cla32_fa27_28_and1;
  wire s_csamul_cla32_fa27_28_or0;
  wire s_csamul_cla32_and28_28;
  wire s_csamul_cla32_fa28_28_xor0;
  wire s_csamul_cla32_fa28_28_and0;
  wire s_csamul_cla32_fa28_28_xor1;
  wire s_csamul_cla32_fa28_28_and1;
  wire s_csamul_cla32_fa28_28_or0;
  wire s_csamul_cla32_and29_28;
  wire s_csamul_cla32_fa29_28_xor0;
  wire s_csamul_cla32_fa29_28_and0;
  wire s_csamul_cla32_fa29_28_xor1;
  wire s_csamul_cla32_fa29_28_and1;
  wire s_csamul_cla32_fa29_28_or0;
  wire s_csamul_cla32_and30_28;
  wire s_csamul_cla32_fa30_28_xor0;
  wire s_csamul_cla32_fa30_28_and0;
  wire s_csamul_cla32_fa30_28_xor1;
  wire s_csamul_cla32_fa30_28_and1;
  wire s_csamul_cla32_fa30_28_or0;
  wire s_csamul_cla32_nand31_28;
  wire s_csamul_cla32_ha31_28_xor0;
  wire s_csamul_cla32_ha31_28_and0;
  wire s_csamul_cla32_and0_29;
  wire s_csamul_cla32_fa0_29_xor0;
  wire s_csamul_cla32_fa0_29_and0;
  wire s_csamul_cla32_fa0_29_xor1;
  wire s_csamul_cla32_fa0_29_and1;
  wire s_csamul_cla32_fa0_29_or0;
  wire s_csamul_cla32_and1_29;
  wire s_csamul_cla32_fa1_29_xor0;
  wire s_csamul_cla32_fa1_29_and0;
  wire s_csamul_cla32_fa1_29_xor1;
  wire s_csamul_cla32_fa1_29_and1;
  wire s_csamul_cla32_fa1_29_or0;
  wire s_csamul_cla32_and2_29;
  wire s_csamul_cla32_fa2_29_xor0;
  wire s_csamul_cla32_fa2_29_and0;
  wire s_csamul_cla32_fa2_29_xor1;
  wire s_csamul_cla32_fa2_29_and1;
  wire s_csamul_cla32_fa2_29_or0;
  wire s_csamul_cla32_and3_29;
  wire s_csamul_cla32_fa3_29_xor0;
  wire s_csamul_cla32_fa3_29_and0;
  wire s_csamul_cla32_fa3_29_xor1;
  wire s_csamul_cla32_fa3_29_and1;
  wire s_csamul_cla32_fa3_29_or0;
  wire s_csamul_cla32_and4_29;
  wire s_csamul_cla32_fa4_29_xor0;
  wire s_csamul_cla32_fa4_29_and0;
  wire s_csamul_cla32_fa4_29_xor1;
  wire s_csamul_cla32_fa4_29_and1;
  wire s_csamul_cla32_fa4_29_or0;
  wire s_csamul_cla32_and5_29;
  wire s_csamul_cla32_fa5_29_xor0;
  wire s_csamul_cla32_fa5_29_and0;
  wire s_csamul_cla32_fa5_29_xor1;
  wire s_csamul_cla32_fa5_29_and1;
  wire s_csamul_cla32_fa5_29_or0;
  wire s_csamul_cla32_and6_29;
  wire s_csamul_cla32_fa6_29_xor0;
  wire s_csamul_cla32_fa6_29_and0;
  wire s_csamul_cla32_fa6_29_xor1;
  wire s_csamul_cla32_fa6_29_and1;
  wire s_csamul_cla32_fa6_29_or0;
  wire s_csamul_cla32_and7_29;
  wire s_csamul_cla32_fa7_29_xor0;
  wire s_csamul_cla32_fa7_29_and0;
  wire s_csamul_cla32_fa7_29_xor1;
  wire s_csamul_cla32_fa7_29_and1;
  wire s_csamul_cla32_fa7_29_or0;
  wire s_csamul_cla32_and8_29;
  wire s_csamul_cla32_fa8_29_xor0;
  wire s_csamul_cla32_fa8_29_and0;
  wire s_csamul_cla32_fa8_29_xor1;
  wire s_csamul_cla32_fa8_29_and1;
  wire s_csamul_cla32_fa8_29_or0;
  wire s_csamul_cla32_and9_29;
  wire s_csamul_cla32_fa9_29_xor0;
  wire s_csamul_cla32_fa9_29_and0;
  wire s_csamul_cla32_fa9_29_xor1;
  wire s_csamul_cla32_fa9_29_and1;
  wire s_csamul_cla32_fa9_29_or0;
  wire s_csamul_cla32_and10_29;
  wire s_csamul_cla32_fa10_29_xor0;
  wire s_csamul_cla32_fa10_29_and0;
  wire s_csamul_cla32_fa10_29_xor1;
  wire s_csamul_cla32_fa10_29_and1;
  wire s_csamul_cla32_fa10_29_or0;
  wire s_csamul_cla32_and11_29;
  wire s_csamul_cla32_fa11_29_xor0;
  wire s_csamul_cla32_fa11_29_and0;
  wire s_csamul_cla32_fa11_29_xor1;
  wire s_csamul_cla32_fa11_29_and1;
  wire s_csamul_cla32_fa11_29_or0;
  wire s_csamul_cla32_and12_29;
  wire s_csamul_cla32_fa12_29_xor0;
  wire s_csamul_cla32_fa12_29_and0;
  wire s_csamul_cla32_fa12_29_xor1;
  wire s_csamul_cla32_fa12_29_and1;
  wire s_csamul_cla32_fa12_29_or0;
  wire s_csamul_cla32_and13_29;
  wire s_csamul_cla32_fa13_29_xor0;
  wire s_csamul_cla32_fa13_29_and0;
  wire s_csamul_cla32_fa13_29_xor1;
  wire s_csamul_cla32_fa13_29_and1;
  wire s_csamul_cla32_fa13_29_or0;
  wire s_csamul_cla32_and14_29;
  wire s_csamul_cla32_fa14_29_xor0;
  wire s_csamul_cla32_fa14_29_and0;
  wire s_csamul_cla32_fa14_29_xor1;
  wire s_csamul_cla32_fa14_29_and1;
  wire s_csamul_cla32_fa14_29_or0;
  wire s_csamul_cla32_and15_29;
  wire s_csamul_cla32_fa15_29_xor0;
  wire s_csamul_cla32_fa15_29_and0;
  wire s_csamul_cla32_fa15_29_xor1;
  wire s_csamul_cla32_fa15_29_and1;
  wire s_csamul_cla32_fa15_29_or0;
  wire s_csamul_cla32_and16_29;
  wire s_csamul_cla32_fa16_29_xor0;
  wire s_csamul_cla32_fa16_29_and0;
  wire s_csamul_cla32_fa16_29_xor1;
  wire s_csamul_cla32_fa16_29_and1;
  wire s_csamul_cla32_fa16_29_or0;
  wire s_csamul_cla32_and17_29;
  wire s_csamul_cla32_fa17_29_xor0;
  wire s_csamul_cla32_fa17_29_and0;
  wire s_csamul_cla32_fa17_29_xor1;
  wire s_csamul_cla32_fa17_29_and1;
  wire s_csamul_cla32_fa17_29_or0;
  wire s_csamul_cla32_and18_29;
  wire s_csamul_cla32_fa18_29_xor0;
  wire s_csamul_cla32_fa18_29_and0;
  wire s_csamul_cla32_fa18_29_xor1;
  wire s_csamul_cla32_fa18_29_and1;
  wire s_csamul_cla32_fa18_29_or0;
  wire s_csamul_cla32_and19_29;
  wire s_csamul_cla32_fa19_29_xor0;
  wire s_csamul_cla32_fa19_29_and0;
  wire s_csamul_cla32_fa19_29_xor1;
  wire s_csamul_cla32_fa19_29_and1;
  wire s_csamul_cla32_fa19_29_or0;
  wire s_csamul_cla32_and20_29;
  wire s_csamul_cla32_fa20_29_xor0;
  wire s_csamul_cla32_fa20_29_and0;
  wire s_csamul_cla32_fa20_29_xor1;
  wire s_csamul_cla32_fa20_29_and1;
  wire s_csamul_cla32_fa20_29_or0;
  wire s_csamul_cla32_and21_29;
  wire s_csamul_cla32_fa21_29_xor0;
  wire s_csamul_cla32_fa21_29_and0;
  wire s_csamul_cla32_fa21_29_xor1;
  wire s_csamul_cla32_fa21_29_and1;
  wire s_csamul_cla32_fa21_29_or0;
  wire s_csamul_cla32_and22_29;
  wire s_csamul_cla32_fa22_29_xor0;
  wire s_csamul_cla32_fa22_29_and0;
  wire s_csamul_cla32_fa22_29_xor1;
  wire s_csamul_cla32_fa22_29_and1;
  wire s_csamul_cla32_fa22_29_or0;
  wire s_csamul_cla32_and23_29;
  wire s_csamul_cla32_fa23_29_xor0;
  wire s_csamul_cla32_fa23_29_and0;
  wire s_csamul_cla32_fa23_29_xor1;
  wire s_csamul_cla32_fa23_29_and1;
  wire s_csamul_cla32_fa23_29_or0;
  wire s_csamul_cla32_and24_29;
  wire s_csamul_cla32_fa24_29_xor0;
  wire s_csamul_cla32_fa24_29_and0;
  wire s_csamul_cla32_fa24_29_xor1;
  wire s_csamul_cla32_fa24_29_and1;
  wire s_csamul_cla32_fa24_29_or0;
  wire s_csamul_cla32_and25_29;
  wire s_csamul_cla32_fa25_29_xor0;
  wire s_csamul_cla32_fa25_29_and0;
  wire s_csamul_cla32_fa25_29_xor1;
  wire s_csamul_cla32_fa25_29_and1;
  wire s_csamul_cla32_fa25_29_or0;
  wire s_csamul_cla32_and26_29;
  wire s_csamul_cla32_fa26_29_xor0;
  wire s_csamul_cla32_fa26_29_and0;
  wire s_csamul_cla32_fa26_29_xor1;
  wire s_csamul_cla32_fa26_29_and1;
  wire s_csamul_cla32_fa26_29_or0;
  wire s_csamul_cla32_and27_29;
  wire s_csamul_cla32_fa27_29_xor0;
  wire s_csamul_cla32_fa27_29_and0;
  wire s_csamul_cla32_fa27_29_xor1;
  wire s_csamul_cla32_fa27_29_and1;
  wire s_csamul_cla32_fa27_29_or0;
  wire s_csamul_cla32_and28_29;
  wire s_csamul_cla32_fa28_29_xor0;
  wire s_csamul_cla32_fa28_29_and0;
  wire s_csamul_cla32_fa28_29_xor1;
  wire s_csamul_cla32_fa28_29_and1;
  wire s_csamul_cla32_fa28_29_or0;
  wire s_csamul_cla32_and29_29;
  wire s_csamul_cla32_fa29_29_xor0;
  wire s_csamul_cla32_fa29_29_and0;
  wire s_csamul_cla32_fa29_29_xor1;
  wire s_csamul_cla32_fa29_29_and1;
  wire s_csamul_cla32_fa29_29_or0;
  wire s_csamul_cla32_and30_29;
  wire s_csamul_cla32_fa30_29_xor0;
  wire s_csamul_cla32_fa30_29_and0;
  wire s_csamul_cla32_fa30_29_xor1;
  wire s_csamul_cla32_fa30_29_and1;
  wire s_csamul_cla32_fa30_29_or0;
  wire s_csamul_cla32_nand31_29;
  wire s_csamul_cla32_ha31_29_xor0;
  wire s_csamul_cla32_ha31_29_and0;
  wire s_csamul_cla32_and0_30;
  wire s_csamul_cla32_fa0_30_xor0;
  wire s_csamul_cla32_fa0_30_and0;
  wire s_csamul_cla32_fa0_30_xor1;
  wire s_csamul_cla32_fa0_30_and1;
  wire s_csamul_cla32_fa0_30_or0;
  wire s_csamul_cla32_and1_30;
  wire s_csamul_cla32_fa1_30_xor0;
  wire s_csamul_cla32_fa1_30_and0;
  wire s_csamul_cla32_fa1_30_xor1;
  wire s_csamul_cla32_fa1_30_and1;
  wire s_csamul_cla32_fa1_30_or0;
  wire s_csamul_cla32_and2_30;
  wire s_csamul_cla32_fa2_30_xor0;
  wire s_csamul_cla32_fa2_30_and0;
  wire s_csamul_cla32_fa2_30_xor1;
  wire s_csamul_cla32_fa2_30_and1;
  wire s_csamul_cla32_fa2_30_or0;
  wire s_csamul_cla32_and3_30;
  wire s_csamul_cla32_fa3_30_xor0;
  wire s_csamul_cla32_fa3_30_and0;
  wire s_csamul_cla32_fa3_30_xor1;
  wire s_csamul_cla32_fa3_30_and1;
  wire s_csamul_cla32_fa3_30_or0;
  wire s_csamul_cla32_and4_30;
  wire s_csamul_cla32_fa4_30_xor0;
  wire s_csamul_cla32_fa4_30_and0;
  wire s_csamul_cla32_fa4_30_xor1;
  wire s_csamul_cla32_fa4_30_and1;
  wire s_csamul_cla32_fa4_30_or0;
  wire s_csamul_cla32_and5_30;
  wire s_csamul_cla32_fa5_30_xor0;
  wire s_csamul_cla32_fa5_30_and0;
  wire s_csamul_cla32_fa5_30_xor1;
  wire s_csamul_cla32_fa5_30_and1;
  wire s_csamul_cla32_fa5_30_or0;
  wire s_csamul_cla32_and6_30;
  wire s_csamul_cla32_fa6_30_xor0;
  wire s_csamul_cla32_fa6_30_and0;
  wire s_csamul_cla32_fa6_30_xor1;
  wire s_csamul_cla32_fa6_30_and1;
  wire s_csamul_cla32_fa6_30_or0;
  wire s_csamul_cla32_and7_30;
  wire s_csamul_cla32_fa7_30_xor0;
  wire s_csamul_cla32_fa7_30_and0;
  wire s_csamul_cla32_fa7_30_xor1;
  wire s_csamul_cla32_fa7_30_and1;
  wire s_csamul_cla32_fa7_30_or0;
  wire s_csamul_cla32_and8_30;
  wire s_csamul_cla32_fa8_30_xor0;
  wire s_csamul_cla32_fa8_30_and0;
  wire s_csamul_cla32_fa8_30_xor1;
  wire s_csamul_cla32_fa8_30_and1;
  wire s_csamul_cla32_fa8_30_or0;
  wire s_csamul_cla32_and9_30;
  wire s_csamul_cla32_fa9_30_xor0;
  wire s_csamul_cla32_fa9_30_and0;
  wire s_csamul_cla32_fa9_30_xor1;
  wire s_csamul_cla32_fa9_30_and1;
  wire s_csamul_cla32_fa9_30_or0;
  wire s_csamul_cla32_and10_30;
  wire s_csamul_cla32_fa10_30_xor0;
  wire s_csamul_cla32_fa10_30_and0;
  wire s_csamul_cla32_fa10_30_xor1;
  wire s_csamul_cla32_fa10_30_and1;
  wire s_csamul_cla32_fa10_30_or0;
  wire s_csamul_cla32_and11_30;
  wire s_csamul_cla32_fa11_30_xor0;
  wire s_csamul_cla32_fa11_30_and0;
  wire s_csamul_cla32_fa11_30_xor1;
  wire s_csamul_cla32_fa11_30_and1;
  wire s_csamul_cla32_fa11_30_or0;
  wire s_csamul_cla32_and12_30;
  wire s_csamul_cla32_fa12_30_xor0;
  wire s_csamul_cla32_fa12_30_and0;
  wire s_csamul_cla32_fa12_30_xor1;
  wire s_csamul_cla32_fa12_30_and1;
  wire s_csamul_cla32_fa12_30_or0;
  wire s_csamul_cla32_and13_30;
  wire s_csamul_cla32_fa13_30_xor0;
  wire s_csamul_cla32_fa13_30_and0;
  wire s_csamul_cla32_fa13_30_xor1;
  wire s_csamul_cla32_fa13_30_and1;
  wire s_csamul_cla32_fa13_30_or0;
  wire s_csamul_cla32_and14_30;
  wire s_csamul_cla32_fa14_30_xor0;
  wire s_csamul_cla32_fa14_30_and0;
  wire s_csamul_cla32_fa14_30_xor1;
  wire s_csamul_cla32_fa14_30_and1;
  wire s_csamul_cla32_fa14_30_or0;
  wire s_csamul_cla32_and15_30;
  wire s_csamul_cla32_fa15_30_xor0;
  wire s_csamul_cla32_fa15_30_and0;
  wire s_csamul_cla32_fa15_30_xor1;
  wire s_csamul_cla32_fa15_30_and1;
  wire s_csamul_cla32_fa15_30_or0;
  wire s_csamul_cla32_and16_30;
  wire s_csamul_cla32_fa16_30_xor0;
  wire s_csamul_cla32_fa16_30_and0;
  wire s_csamul_cla32_fa16_30_xor1;
  wire s_csamul_cla32_fa16_30_and1;
  wire s_csamul_cla32_fa16_30_or0;
  wire s_csamul_cla32_and17_30;
  wire s_csamul_cla32_fa17_30_xor0;
  wire s_csamul_cla32_fa17_30_and0;
  wire s_csamul_cla32_fa17_30_xor1;
  wire s_csamul_cla32_fa17_30_and1;
  wire s_csamul_cla32_fa17_30_or0;
  wire s_csamul_cla32_and18_30;
  wire s_csamul_cla32_fa18_30_xor0;
  wire s_csamul_cla32_fa18_30_and0;
  wire s_csamul_cla32_fa18_30_xor1;
  wire s_csamul_cla32_fa18_30_and1;
  wire s_csamul_cla32_fa18_30_or0;
  wire s_csamul_cla32_and19_30;
  wire s_csamul_cla32_fa19_30_xor0;
  wire s_csamul_cla32_fa19_30_and0;
  wire s_csamul_cla32_fa19_30_xor1;
  wire s_csamul_cla32_fa19_30_and1;
  wire s_csamul_cla32_fa19_30_or0;
  wire s_csamul_cla32_and20_30;
  wire s_csamul_cla32_fa20_30_xor0;
  wire s_csamul_cla32_fa20_30_and0;
  wire s_csamul_cla32_fa20_30_xor1;
  wire s_csamul_cla32_fa20_30_and1;
  wire s_csamul_cla32_fa20_30_or0;
  wire s_csamul_cla32_and21_30;
  wire s_csamul_cla32_fa21_30_xor0;
  wire s_csamul_cla32_fa21_30_and0;
  wire s_csamul_cla32_fa21_30_xor1;
  wire s_csamul_cla32_fa21_30_and1;
  wire s_csamul_cla32_fa21_30_or0;
  wire s_csamul_cla32_and22_30;
  wire s_csamul_cla32_fa22_30_xor0;
  wire s_csamul_cla32_fa22_30_and0;
  wire s_csamul_cla32_fa22_30_xor1;
  wire s_csamul_cla32_fa22_30_and1;
  wire s_csamul_cla32_fa22_30_or0;
  wire s_csamul_cla32_and23_30;
  wire s_csamul_cla32_fa23_30_xor0;
  wire s_csamul_cla32_fa23_30_and0;
  wire s_csamul_cla32_fa23_30_xor1;
  wire s_csamul_cla32_fa23_30_and1;
  wire s_csamul_cla32_fa23_30_or0;
  wire s_csamul_cla32_and24_30;
  wire s_csamul_cla32_fa24_30_xor0;
  wire s_csamul_cla32_fa24_30_and0;
  wire s_csamul_cla32_fa24_30_xor1;
  wire s_csamul_cla32_fa24_30_and1;
  wire s_csamul_cla32_fa24_30_or0;
  wire s_csamul_cla32_and25_30;
  wire s_csamul_cla32_fa25_30_xor0;
  wire s_csamul_cla32_fa25_30_and0;
  wire s_csamul_cla32_fa25_30_xor1;
  wire s_csamul_cla32_fa25_30_and1;
  wire s_csamul_cla32_fa25_30_or0;
  wire s_csamul_cla32_and26_30;
  wire s_csamul_cla32_fa26_30_xor0;
  wire s_csamul_cla32_fa26_30_and0;
  wire s_csamul_cla32_fa26_30_xor1;
  wire s_csamul_cla32_fa26_30_and1;
  wire s_csamul_cla32_fa26_30_or0;
  wire s_csamul_cla32_and27_30;
  wire s_csamul_cla32_fa27_30_xor0;
  wire s_csamul_cla32_fa27_30_and0;
  wire s_csamul_cla32_fa27_30_xor1;
  wire s_csamul_cla32_fa27_30_and1;
  wire s_csamul_cla32_fa27_30_or0;
  wire s_csamul_cla32_and28_30;
  wire s_csamul_cla32_fa28_30_xor0;
  wire s_csamul_cla32_fa28_30_and0;
  wire s_csamul_cla32_fa28_30_xor1;
  wire s_csamul_cla32_fa28_30_and1;
  wire s_csamul_cla32_fa28_30_or0;
  wire s_csamul_cla32_and29_30;
  wire s_csamul_cla32_fa29_30_xor0;
  wire s_csamul_cla32_fa29_30_and0;
  wire s_csamul_cla32_fa29_30_xor1;
  wire s_csamul_cla32_fa29_30_and1;
  wire s_csamul_cla32_fa29_30_or0;
  wire s_csamul_cla32_and30_30;
  wire s_csamul_cla32_fa30_30_xor0;
  wire s_csamul_cla32_fa30_30_and0;
  wire s_csamul_cla32_fa30_30_xor1;
  wire s_csamul_cla32_fa30_30_and1;
  wire s_csamul_cla32_fa30_30_or0;
  wire s_csamul_cla32_nand31_30;
  wire s_csamul_cla32_ha31_30_xor0;
  wire s_csamul_cla32_ha31_30_and0;
  wire s_csamul_cla32_nand0_31;
  wire s_csamul_cla32_fa0_31_xor0;
  wire s_csamul_cla32_fa0_31_and0;
  wire s_csamul_cla32_fa0_31_xor1;
  wire s_csamul_cla32_fa0_31_and1;
  wire s_csamul_cla32_fa0_31_or0;
  wire s_csamul_cla32_nand1_31;
  wire s_csamul_cla32_fa1_31_xor0;
  wire s_csamul_cla32_fa1_31_and0;
  wire s_csamul_cla32_fa1_31_xor1;
  wire s_csamul_cla32_fa1_31_and1;
  wire s_csamul_cla32_fa1_31_or0;
  wire s_csamul_cla32_nand2_31;
  wire s_csamul_cla32_fa2_31_xor0;
  wire s_csamul_cla32_fa2_31_and0;
  wire s_csamul_cla32_fa2_31_xor1;
  wire s_csamul_cla32_fa2_31_and1;
  wire s_csamul_cla32_fa2_31_or0;
  wire s_csamul_cla32_nand3_31;
  wire s_csamul_cla32_fa3_31_xor0;
  wire s_csamul_cla32_fa3_31_and0;
  wire s_csamul_cla32_fa3_31_xor1;
  wire s_csamul_cla32_fa3_31_and1;
  wire s_csamul_cla32_fa3_31_or0;
  wire s_csamul_cla32_nand4_31;
  wire s_csamul_cla32_fa4_31_xor0;
  wire s_csamul_cla32_fa4_31_and0;
  wire s_csamul_cla32_fa4_31_xor1;
  wire s_csamul_cla32_fa4_31_and1;
  wire s_csamul_cla32_fa4_31_or0;
  wire s_csamul_cla32_nand5_31;
  wire s_csamul_cla32_fa5_31_xor0;
  wire s_csamul_cla32_fa5_31_and0;
  wire s_csamul_cla32_fa5_31_xor1;
  wire s_csamul_cla32_fa5_31_and1;
  wire s_csamul_cla32_fa5_31_or0;
  wire s_csamul_cla32_nand6_31;
  wire s_csamul_cla32_fa6_31_xor0;
  wire s_csamul_cla32_fa6_31_and0;
  wire s_csamul_cla32_fa6_31_xor1;
  wire s_csamul_cla32_fa6_31_and1;
  wire s_csamul_cla32_fa6_31_or0;
  wire s_csamul_cla32_nand7_31;
  wire s_csamul_cla32_fa7_31_xor0;
  wire s_csamul_cla32_fa7_31_and0;
  wire s_csamul_cla32_fa7_31_xor1;
  wire s_csamul_cla32_fa7_31_and1;
  wire s_csamul_cla32_fa7_31_or0;
  wire s_csamul_cla32_nand8_31;
  wire s_csamul_cla32_fa8_31_xor0;
  wire s_csamul_cla32_fa8_31_and0;
  wire s_csamul_cla32_fa8_31_xor1;
  wire s_csamul_cla32_fa8_31_and1;
  wire s_csamul_cla32_fa8_31_or0;
  wire s_csamul_cla32_nand9_31;
  wire s_csamul_cla32_fa9_31_xor0;
  wire s_csamul_cla32_fa9_31_and0;
  wire s_csamul_cla32_fa9_31_xor1;
  wire s_csamul_cla32_fa9_31_and1;
  wire s_csamul_cla32_fa9_31_or0;
  wire s_csamul_cla32_nand10_31;
  wire s_csamul_cla32_fa10_31_xor0;
  wire s_csamul_cla32_fa10_31_and0;
  wire s_csamul_cla32_fa10_31_xor1;
  wire s_csamul_cla32_fa10_31_and1;
  wire s_csamul_cla32_fa10_31_or0;
  wire s_csamul_cla32_nand11_31;
  wire s_csamul_cla32_fa11_31_xor0;
  wire s_csamul_cla32_fa11_31_and0;
  wire s_csamul_cla32_fa11_31_xor1;
  wire s_csamul_cla32_fa11_31_and1;
  wire s_csamul_cla32_fa11_31_or0;
  wire s_csamul_cla32_nand12_31;
  wire s_csamul_cla32_fa12_31_xor0;
  wire s_csamul_cla32_fa12_31_and0;
  wire s_csamul_cla32_fa12_31_xor1;
  wire s_csamul_cla32_fa12_31_and1;
  wire s_csamul_cla32_fa12_31_or0;
  wire s_csamul_cla32_nand13_31;
  wire s_csamul_cla32_fa13_31_xor0;
  wire s_csamul_cla32_fa13_31_and0;
  wire s_csamul_cla32_fa13_31_xor1;
  wire s_csamul_cla32_fa13_31_and1;
  wire s_csamul_cla32_fa13_31_or0;
  wire s_csamul_cla32_nand14_31;
  wire s_csamul_cla32_fa14_31_xor0;
  wire s_csamul_cla32_fa14_31_and0;
  wire s_csamul_cla32_fa14_31_xor1;
  wire s_csamul_cla32_fa14_31_and1;
  wire s_csamul_cla32_fa14_31_or0;
  wire s_csamul_cla32_nand15_31;
  wire s_csamul_cla32_fa15_31_xor0;
  wire s_csamul_cla32_fa15_31_and0;
  wire s_csamul_cla32_fa15_31_xor1;
  wire s_csamul_cla32_fa15_31_and1;
  wire s_csamul_cla32_fa15_31_or0;
  wire s_csamul_cla32_nand16_31;
  wire s_csamul_cla32_fa16_31_xor0;
  wire s_csamul_cla32_fa16_31_and0;
  wire s_csamul_cla32_fa16_31_xor1;
  wire s_csamul_cla32_fa16_31_and1;
  wire s_csamul_cla32_fa16_31_or0;
  wire s_csamul_cla32_nand17_31;
  wire s_csamul_cla32_fa17_31_xor0;
  wire s_csamul_cla32_fa17_31_and0;
  wire s_csamul_cla32_fa17_31_xor1;
  wire s_csamul_cla32_fa17_31_and1;
  wire s_csamul_cla32_fa17_31_or0;
  wire s_csamul_cla32_nand18_31;
  wire s_csamul_cla32_fa18_31_xor0;
  wire s_csamul_cla32_fa18_31_and0;
  wire s_csamul_cla32_fa18_31_xor1;
  wire s_csamul_cla32_fa18_31_and1;
  wire s_csamul_cla32_fa18_31_or0;
  wire s_csamul_cla32_nand19_31;
  wire s_csamul_cla32_fa19_31_xor0;
  wire s_csamul_cla32_fa19_31_and0;
  wire s_csamul_cla32_fa19_31_xor1;
  wire s_csamul_cla32_fa19_31_and1;
  wire s_csamul_cla32_fa19_31_or0;
  wire s_csamul_cla32_nand20_31;
  wire s_csamul_cla32_fa20_31_xor0;
  wire s_csamul_cla32_fa20_31_and0;
  wire s_csamul_cla32_fa20_31_xor1;
  wire s_csamul_cla32_fa20_31_and1;
  wire s_csamul_cla32_fa20_31_or0;
  wire s_csamul_cla32_nand21_31;
  wire s_csamul_cla32_fa21_31_xor0;
  wire s_csamul_cla32_fa21_31_and0;
  wire s_csamul_cla32_fa21_31_xor1;
  wire s_csamul_cla32_fa21_31_and1;
  wire s_csamul_cla32_fa21_31_or0;
  wire s_csamul_cla32_nand22_31;
  wire s_csamul_cla32_fa22_31_xor0;
  wire s_csamul_cla32_fa22_31_and0;
  wire s_csamul_cla32_fa22_31_xor1;
  wire s_csamul_cla32_fa22_31_and1;
  wire s_csamul_cla32_fa22_31_or0;
  wire s_csamul_cla32_nand23_31;
  wire s_csamul_cla32_fa23_31_xor0;
  wire s_csamul_cla32_fa23_31_and0;
  wire s_csamul_cla32_fa23_31_xor1;
  wire s_csamul_cla32_fa23_31_and1;
  wire s_csamul_cla32_fa23_31_or0;
  wire s_csamul_cla32_nand24_31;
  wire s_csamul_cla32_fa24_31_xor0;
  wire s_csamul_cla32_fa24_31_and0;
  wire s_csamul_cla32_fa24_31_xor1;
  wire s_csamul_cla32_fa24_31_and1;
  wire s_csamul_cla32_fa24_31_or0;
  wire s_csamul_cla32_nand25_31;
  wire s_csamul_cla32_fa25_31_xor0;
  wire s_csamul_cla32_fa25_31_and0;
  wire s_csamul_cla32_fa25_31_xor1;
  wire s_csamul_cla32_fa25_31_and1;
  wire s_csamul_cla32_fa25_31_or0;
  wire s_csamul_cla32_nand26_31;
  wire s_csamul_cla32_fa26_31_xor0;
  wire s_csamul_cla32_fa26_31_and0;
  wire s_csamul_cla32_fa26_31_xor1;
  wire s_csamul_cla32_fa26_31_and1;
  wire s_csamul_cla32_fa26_31_or0;
  wire s_csamul_cla32_nand27_31;
  wire s_csamul_cla32_fa27_31_xor0;
  wire s_csamul_cla32_fa27_31_and0;
  wire s_csamul_cla32_fa27_31_xor1;
  wire s_csamul_cla32_fa27_31_and1;
  wire s_csamul_cla32_fa27_31_or0;
  wire s_csamul_cla32_nand28_31;
  wire s_csamul_cla32_fa28_31_xor0;
  wire s_csamul_cla32_fa28_31_and0;
  wire s_csamul_cla32_fa28_31_xor1;
  wire s_csamul_cla32_fa28_31_and1;
  wire s_csamul_cla32_fa28_31_or0;
  wire s_csamul_cla32_nand29_31;
  wire s_csamul_cla32_fa29_31_xor0;
  wire s_csamul_cla32_fa29_31_and0;
  wire s_csamul_cla32_fa29_31_xor1;
  wire s_csamul_cla32_fa29_31_and1;
  wire s_csamul_cla32_fa29_31_or0;
  wire s_csamul_cla32_nand30_31;
  wire s_csamul_cla32_fa30_31_xor0;
  wire s_csamul_cla32_fa30_31_and0;
  wire s_csamul_cla32_fa30_31_xor1;
  wire s_csamul_cla32_fa30_31_and1;
  wire s_csamul_cla32_fa30_31_or0;
  wire s_csamul_cla32_and31_31;
  wire s_csamul_cla32_ha31_31_xor0;
  wire s_csamul_cla32_ha31_31_and0;
  wire s_csamul_cla32_u_cla32_pg_logic0_or0;
  wire s_csamul_cla32_u_cla32_pg_logic0_and0;
  wire s_csamul_cla32_u_cla32_pg_logic0_xor0;
  wire s_csamul_cla32_u_cla32_pg_logic1_or0;
  wire s_csamul_cla32_u_cla32_pg_logic1_and0;
  wire s_csamul_cla32_u_cla32_pg_logic1_xor0;
  wire s_csamul_cla32_u_cla32_xor1;
  wire s_csamul_cla32_u_cla32_and0;
  wire s_csamul_cla32_u_cla32_or0;
  wire s_csamul_cla32_u_cla32_pg_logic2_or0;
  wire s_csamul_cla32_u_cla32_pg_logic2_and0;
  wire s_csamul_cla32_u_cla32_pg_logic2_xor0;
  wire s_csamul_cla32_u_cla32_xor2;
  wire s_csamul_cla32_u_cla32_and1;
  wire s_csamul_cla32_u_cla32_and2;
  wire s_csamul_cla32_u_cla32_and3;
  wire s_csamul_cla32_u_cla32_and4;
  wire s_csamul_cla32_u_cla32_or1;
  wire s_csamul_cla32_u_cla32_or2;
  wire s_csamul_cla32_u_cla32_pg_logic3_or0;
  wire s_csamul_cla32_u_cla32_pg_logic3_and0;
  wire s_csamul_cla32_u_cla32_pg_logic3_xor0;
  wire s_csamul_cla32_u_cla32_xor3;
  wire s_csamul_cla32_u_cla32_and5;
  wire s_csamul_cla32_u_cla32_and6;
  wire s_csamul_cla32_u_cla32_and7;
  wire s_csamul_cla32_u_cla32_and8;
  wire s_csamul_cla32_u_cla32_and9;
  wire s_csamul_cla32_u_cla32_and10;
  wire s_csamul_cla32_u_cla32_and11;
  wire s_csamul_cla32_u_cla32_or3;
  wire s_csamul_cla32_u_cla32_or4;
  wire s_csamul_cla32_u_cla32_or5;
  wire s_csamul_cla32_u_cla32_pg_logic4_or0;
  wire s_csamul_cla32_u_cla32_pg_logic4_and0;
  wire s_csamul_cla32_u_cla32_pg_logic4_xor0;
  wire s_csamul_cla32_u_cla32_xor4;
  wire s_csamul_cla32_u_cla32_and12;
  wire s_csamul_cla32_u_cla32_or6;
  wire s_csamul_cla32_u_cla32_pg_logic5_or0;
  wire s_csamul_cla32_u_cla32_pg_logic5_and0;
  wire s_csamul_cla32_u_cla32_pg_logic5_xor0;
  wire s_csamul_cla32_u_cla32_xor5;
  wire s_csamul_cla32_u_cla32_and13;
  wire s_csamul_cla32_u_cla32_and14;
  wire s_csamul_cla32_u_cla32_and15;
  wire s_csamul_cla32_u_cla32_or7;
  wire s_csamul_cla32_u_cla32_or8;
  wire s_csamul_cla32_u_cla32_pg_logic6_or0;
  wire s_csamul_cla32_u_cla32_pg_logic6_and0;
  wire s_csamul_cla32_u_cla32_pg_logic6_xor0;
  wire s_csamul_cla32_u_cla32_xor6;
  wire s_csamul_cla32_u_cla32_and16;
  wire s_csamul_cla32_u_cla32_and17;
  wire s_csamul_cla32_u_cla32_and18;
  wire s_csamul_cla32_u_cla32_and19;
  wire s_csamul_cla32_u_cla32_and20;
  wire s_csamul_cla32_u_cla32_and21;
  wire s_csamul_cla32_u_cla32_or9;
  wire s_csamul_cla32_u_cla32_or10;
  wire s_csamul_cla32_u_cla32_or11;
  wire s_csamul_cla32_u_cla32_pg_logic7_or0;
  wire s_csamul_cla32_u_cla32_pg_logic7_and0;
  wire s_csamul_cla32_u_cla32_pg_logic7_xor0;
  wire s_csamul_cla32_u_cla32_xor7;
  wire s_csamul_cla32_u_cla32_and22;
  wire s_csamul_cla32_u_cla32_and23;
  wire s_csamul_cla32_u_cla32_and24;
  wire s_csamul_cla32_u_cla32_and25;
  wire s_csamul_cla32_u_cla32_and26;
  wire s_csamul_cla32_u_cla32_and27;
  wire s_csamul_cla32_u_cla32_and28;
  wire s_csamul_cla32_u_cla32_and29;
  wire s_csamul_cla32_u_cla32_and30;
  wire s_csamul_cla32_u_cla32_and31;
  wire s_csamul_cla32_u_cla32_or12;
  wire s_csamul_cla32_u_cla32_or13;
  wire s_csamul_cla32_u_cla32_or14;
  wire s_csamul_cla32_u_cla32_or15;
  wire s_csamul_cla32_u_cla32_pg_logic8_or0;
  wire s_csamul_cla32_u_cla32_pg_logic8_and0;
  wire s_csamul_cla32_u_cla32_pg_logic8_xor0;
  wire s_csamul_cla32_u_cla32_xor8;
  wire s_csamul_cla32_u_cla32_and32;
  wire s_csamul_cla32_u_cla32_or16;
  wire s_csamul_cla32_u_cla32_pg_logic9_or0;
  wire s_csamul_cla32_u_cla32_pg_logic9_and0;
  wire s_csamul_cla32_u_cla32_pg_logic9_xor0;
  wire s_csamul_cla32_u_cla32_xor9;
  wire s_csamul_cla32_u_cla32_and33;
  wire s_csamul_cla32_u_cla32_and34;
  wire s_csamul_cla32_u_cla32_and35;
  wire s_csamul_cla32_u_cla32_or17;
  wire s_csamul_cla32_u_cla32_or18;
  wire s_csamul_cla32_u_cla32_pg_logic10_or0;
  wire s_csamul_cla32_u_cla32_pg_logic10_and0;
  wire s_csamul_cla32_u_cla32_pg_logic10_xor0;
  wire s_csamul_cla32_u_cla32_xor10;
  wire s_csamul_cla32_u_cla32_and36;
  wire s_csamul_cla32_u_cla32_and37;
  wire s_csamul_cla32_u_cla32_and38;
  wire s_csamul_cla32_u_cla32_and39;
  wire s_csamul_cla32_u_cla32_and40;
  wire s_csamul_cla32_u_cla32_and41;
  wire s_csamul_cla32_u_cla32_or19;
  wire s_csamul_cla32_u_cla32_or20;
  wire s_csamul_cla32_u_cla32_or21;
  wire s_csamul_cla32_u_cla32_pg_logic11_or0;
  wire s_csamul_cla32_u_cla32_pg_logic11_and0;
  wire s_csamul_cla32_u_cla32_pg_logic11_xor0;
  wire s_csamul_cla32_u_cla32_xor11;
  wire s_csamul_cla32_u_cla32_and42;
  wire s_csamul_cla32_u_cla32_and43;
  wire s_csamul_cla32_u_cla32_and44;
  wire s_csamul_cla32_u_cla32_and45;
  wire s_csamul_cla32_u_cla32_and46;
  wire s_csamul_cla32_u_cla32_and47;
  wire s_csamul_cla32_u_cla32_and48;
  wire s_csamul_cla32_u_cla32_and49;
  wire s_csamul_cla32_u_cla32_and50;
  wire s_csamul_cla32_u_cla32_and51;
  wire s_csamul_cla32_u_cla32_or22;
  wire s_csamul_cla32_u_cla32_or23;
  wire s_csamul_cla32_u_cla32_or24;
  wire s_csamul_cla32_u_cla32_or25;
  wire s_csamul_cla32_u_cla32_pg_logic12_or0;
  wire s_csamul_cla32_u_cla32_pg_logic12_and0;
  wire s_csamul_cla32_u_cla32_pg_logic12_xor0;
  wire s_csamul_cla32_u_cla32_xor12;
  wire s_csamul_cla32_u_cla32_and52;
  wire s_csamul_cla32_u_cla32_or26;
  wire s_csamul_cla32_u_cla32_pg_logic13_or0;
  wire s_csamul_cla32_u_cla32_pg_logic13_and0;
  wire s_csamul_cla32_u_cla32_pg_logic13_xor0;
  wire s_csamul_cla32_u_cla32_xor13;
  wire s_csamul_cla32_u_cla32_and53;
  wire s_csamul_cla32_u_cla32_and54;
  wire s_csamul_cla32_u_cla32_and55;
  wire s_csamul_cla32_u_cla32_or27;
  wire s_csamul_cla32_u_cla32_or28;
  wire s_csamul_cla32_u_cla32_pg_logic14_or0;
  wire s_csamul_cla32_u_cla32_pg_logic14_and0;
  wire s_csamul_cla32_u_cla32_pg_logic14_xor0;
  wire s_csamul_cla32_u_cla32_xor14;
  wire s_csamul_cla32_u_cla32_and56;
  wire s_csamul_cla32_u_cla32_and57;
  wire s_csamul_cla32_u_cla32_and58;
  wire s_csamul_cla32_u_cla32_and59;
  wire s_csamul_cla32_u_cla32_and60;
  wire s_csamul_cla32_u_cla32_and61;
  wire s_csamul_cla32_u_cla32_or29;
  wire s_csamul_cla32_u_cla32_or30;
  wire s_csamul_cla32_u_cla32_or31;
  wire s_csamul_cla32_u_cla32_pg_logic15_or0;
  wire s_csamul_cla32_u_cla32_pg_logic15_and0;
  wire s_csamul_cla32_u_cla32_pg_logic15_xor0;
  wire s_csamul_cla32_u_cla32_xor15;
  wire s_csamul_cla32_u_cla32_and62;
  wire s_csamul_cla32_u_cla32_and63;
  wire s_csamul_cla32_u_cla32_and64;
  wire s_csamul_cla32_u_cla32_and65;
  wire s_csamul_cla32_u_cla32_and66;
  wire s_csamul_cla32_u_cla32_and67;
  wire s_csamul_cla32_u_cla32_and68;
  wire s_csamul_cla32_u_cla32_and69;
  wire s_csamul_cla32_u_cla32_and70;
  wire s_csamul_cla32_u_cla32_and71;
  wire s_csamul_cla32_u_cla32_or32;
  wire s_csamul_cla32_u_cla32_or33;
  wire s_csamul_cla32_u_cla32_or34;
  wire s_csamul_cla32_u_cla32_or35;
  wire s_csamul_cla32_u_cla32_pg_logic16_or0;
  wire s_csamul_cla32_u_cla32_pg_logic16_and0;
  wire s_csamul_cla32_u_cla32_pg_logic16_xor0;
  wire s_csamul_cla32_u_cla32_xor16;
  wire s_csamul_cla32_u_cla32_and72;
  wire s_csamul_cla32_u_cla32_or36;
  wire s_csamul_cla32_u_cla32_pg_logic17_or0;
  wire s_csamul_cla32_u_cla32_pg_logic17_and0;
  wire s_csamul_cla32_u_cla32_pg_logic17_xor0;
  wire s_csamul_cla32_u_cla32_xor17;
  wire s_csamul_cla32_u_cla32_and73;
  wire s_csamul_cla32_u_cla32_and74;
  wire s_csamul_cla32_u_cla32_and75;
  wire s_csamul_cla32_u_cla32_or37;
  wire s_csamul_cla32_u_cla32_or38;
  wire s_csamul_cla32_u_cla32_pg_logic18_or0;
  wire s_csamul_cla32_u_cla32_pg_logic18_and0;
  wire s_csamul_cla32_u_cla32_pg_logic18_xor0;
  wire s_csamul_cla32_u_cla32_xor18;
  wire s_csamul_cla32_u_cla32_and76;
  wire s_csamul_cla32_u_cla32_and77;
  wire s_csamul_cla32_u_cla32_and78;
  wire s_csamul_cla32_u_cla32_and79;
  wire s_csamul_cla32_u_cla32_and80;
  wire s_csamul_cla32_u_cla32_and81;
  wire s_csamul_cla32_u_cla32_or39;
  wire s_csamul_cla32_u_cla32_or40;
  wire s_csamul_cla32_u_cla32_or41;
  wire s_csamul_cla32_u_cla32_pg_logic19_or0;
  wire s_csamul_cla32_u_cla32_pg_logic19_and0;
  wire s_csamul_cla32_u_cla32_pg_logic19_xor0;
  wire s_csamul_cla32_u_cla32_xor19;
  wire s_csamul_cla32_u_cla32_and82;
  wire s_csamul_cla32_u_cla32_and83;
  wire s_csamul_cla32_u_cla32_and84;
  wire s_csamul_cla32_u_cla32_and85;
  wire s_csamul_cla32_u_cla32_and86;
  wire s_csamul_cla32_u_cla32_and87;
  wire s_csamul_cla32_u_cla32_and88;
  wire s_csamul_cla32_u_cla32_and89;
  wire s_csamul_cla32_u_cla32_and90;
  wire s_csamul_cla32_u_cla32_and91;
  wire s_csamul_cla32_u_cla32_or42;
  wire s_csamul_cla32_u_cla32_or43;
  wire s_csamul_cla32_u_cla32_or44;
  wire s_csamul_cla32_u_cla32_or45;
  wire s_csamul_cla32_u_cla32_pg_logic20_or0;
  wire s_csamul_cla32_u_cla32_pg_logic20_and0;
  wire s_csamul_cla32_u_cla32_pg_logic20_xor0;
  wire s_csamul_cla32_u_cla32_xor20;
  wire s_csamul_cla32_u_cla32_and92;
  wire s_csamul_cla32_u_cla32_or46;
  wire s_csamul_cla32_u_cla32_pg_logic21_or0;
  wire s_csamul_cla32_u_cla32_pg_logic21_and0;
  wire s_csamul_cla32_u_cla32_pg_logic21_xor0;
  wire s_csamul_cla32_u_cla32_xor21;
  wire s_csamul_cla32_u_cla32_and93;
  wire s_csamul_cla32_u_cla32_and94;
  wire s_csamul_cla32_u_cla32_and95;
  wire s_csamul_cla32_u_cla32_or47;
  wire s_csamul_cla32_u_cla32_or48;
  wire s_csamul_cla32_u_cla32_pg_logic22_or0;
  wire s_csamul_cla32_u_cla32_pg_logic22_and0;
  wire s_csamul_cla32_u_cla32_pg_logic22_xor0;
  wire s_csamul_cla32_u_cla32_xor22;
  wire s_csamul_cla32_u_cla32_and96;
  wire s_csamul_cla32_u_cla32_and97;
  wire s_csamul_cla32_u_cla32_and98;
  wire s_csamul_cla32_u_cla32_and99;
  wire s_csamul_cla32_u_cla32_and100;
  wire s_csamul_cla32_u_cla32_and101;
  wire s_csamul_cla32_u_cla32_or49;
  wire s_csamul_cla32_u_cla32_or50;
  wire s_csamul_cla32_u_cla32_or51;
  wire s_csamul_cla32_u_cla32_pg_logic23_or0;
  wire s_csamul_cla32_u_cla32_pg_logic23_and0;
  wire s_csamul_cla32_u_cla32_pg_logic23_xor0;
  wire s_csamul_cla32_u_cla32_xor23;
  wire s_csamul_cla32_u_cla32_and102;
  wire s_csamul_cla32_u_cla32_and103;
  wire s_csamul_cla32_u_cla32_and104;
  wire s_csamul_cla32_u_cla32_and105;
  wire s_csamul_cla32_u_cla32_and106;
  wire s_csamul_cla32_u_cla32_and107;
  wire s_csamul_cla32_u_cla32_and108;
  wire s_csamul_cla32_u_cla32_and109;
  wire s_csamul_cla32_u_cla32_and110;
  wire s_csamul_cla32_u_cla32_and111;
  wire s_csamul_cla32_u_cla32_or52;
  wire s_csamul_cla32_u_cla32_or53;
  wire s_csamul_cla32_u_cla32_or54;
  wire s_csamul_cla32_u_cla32_or55;
  wire s_csamul_cla32_u_cla32_pg_logic24_or0;
  wire s_csamul_cla32_u_cla32_pg_logic24_and0;
  wire s_csamul_cla32_u_cla32_pg_logic24_xor0;
  wire s_csamul_cla32_u_cla32_xor24;
  wire s_csamul_cla32_u_cla32_and112;
  wire s_csamul_cla32_u_cla32_or56;
  wire s_csamul_cla32_u_cla32_pg_logic25_or0;
  wire s_csamul_cla32_u_cla32_pg_logic25_and0;
  wire s_csamul_cla32_u_cla32_pg_logic25_xor0;
  wire s_csamul_cla32_u_cla32_xor25;
  wire s_csamul_cla32_u_cla32_and113;
  wire s_csamul_cla32_u_cla32_and114;
  wire s_csamul_cla32_u_cla32_and115;
  wire s_csamul_cla32_u_cla32_or57;
  wire s_csamul_cla32_u_cla32_or58;
  wire s_csamul_cla32_u_cla32_pg_logic26_or0;
  wire s_csamul_cla32_u_cla32_pg_logic26_and0;
  wire s_csamul_cla32_u_cla32_pg_logic26_xor0;
  wire s_csamul_cla32_u_cla32_xor26;
  wire s_csamul_cla32_u_cla32_and116;
  wire s_csamul_cla32_u_cla32_and117;
  wire s_csamul_cla32_u_cla32_and118;
  wire s_csamul_cla32_u_cla32_and119;
  wire s_csamul_cla32_u_cla32_and120;
  wire s_csamul_cla32_u_cla32_and121;
  wire s_csamul_cla32_u_cla32_or59;
  wire s_csamul_cla32_u_cla32_or60;
  wire s_csamul_cla32_u_cla32_or61;
  wire s_csamul_cla32_u_cla32_pg_logic27_or0;
  wire s_csamul_cla32_u_cla32_pg_logic27_and0;
  wire s_csamul_cla32_u_cla32_pg_logic27_xor0;
  wire s_csamul_cla32_u_cla32_xor27;
  wire s_csamul_cla32_u_cla32_and122;
  wire s_csamul_cla32_u_cla32_and123;
  wire s_csamul_cla32_u_cla32_and124;
  wire s_csamul_cla32_u_cla32_and125;
  wire s_csamul_cla32_u_cla32_and126;
  wire s_csamul_cla32_u_cla32_and127;
  wire s_csamul_cla32_u_cla32_and128;
  wire s_csamul_cla32_u_cla32_and129;
  wire s_csamul_cla32_u_cla32_and130;
  wire s_csamul_cla32_u_cla32_and131;
  wire s_csamul_cla32_u_cla32_or62;
  wire s_csamul_cla32_u_cla32_or63;
  wire s_csamul_cla32_u_cla32_or64;
  wire s_csamul_cla32_u_cla32_or65;
  wire s_csamul_cla32_u_cla32_pg_logic28_or0;
  wire s_csamul_cla32_u_cla32_pg_logic28_and0;
  wire s_csamul_cla32_u_cla32_pg_logic28_xor0;
  wire s_csamul_cla32_u_cla32_xor28;
  wire s_csamul_cla32_u_cla32_and132;
  wire s_csamul_cla32_u_cla32_or66;
  wire s_csamul_cla32_u_cla32_pg_logic29_or0;
  wire s_csamul_cla32_u_cla32_pg_logic29_and0;
  wire s_csamul_cla32_u_cla32_pg_logic29_xor0;
  wire s_csamul_cla32_u_cla32_xor29;
  wire s_csamul_cla32_u_cla32_and133;
  wire s_csamul_cla32_u_cla32_and134;
  wire s_csamul_cla32_u_cla32_and135;
  wire s_csamul_cla32_u_cla32_or67;
  wire s_csamul_cla32_u_cla32_or68;
  wire s_csamul_cla32_u_cla32_pg_logic30_or0;
  wire s_csamul_cla32_u_cla32_pg_logic30_and0;
  wire s_csamul_cla32_u_cla32_pg_logic30_xor0;
  wire s_csamul_cla32_u_cla32_xor30;
  wire s_csamul_cla32_u_cla32_and136;
  wire s_csamul_cla32_u_cla32_and137;
  wire s_csamul_cla32_u_cla32_and138;
  wire s_csamul_cla32_u_cla32_and139;
  wire s_csamul_cla32_u_cla32_and140;
  wire s_csamul_cla32_u_cla32_and141;
  wire s_csamul_cla32_u_cla32_or69;
  wire s_csamul_cla32_u_cla32_or70;
  wire s_csamul_cla32_u_cla32_or71;
  wire s_csamul_cla32_u_cla32_pg_logic31_xor0;
  wire s_csamul_cla32_u_cla32_xor31;
  wire s_csamul_cla32_u_cla32_and142;
  wire s_csamul_cla32_u_cla32_and143;
  wire s_csamul_cla32_u_cla32_and144;
  wire s_csamul_cla32_u_cla32_and145;
  wire s_csamul_cla32_u_cla32_and146;
  wire s_csamul_cla32_u_cla32_and147;
  wire s_csamul_cla32_u_cla32_or72;
  wire s_csamul_cla32_u_cla32_or73;
  wire s_csamul_cla32_u_cla32_or74;
  wire s_csamul_cla32_u_cla32_or75;

  assign s_csamul_cla32_and0_0 = a[0] & b[0];
  assign s_csamul_cla32_and1_0 = a[1] & b[0];
  assign s_csamul_cla32_and2_0 = a[2] & b[0];
  assign s_csamul_cla32_and3_0 = a[3] & b[0];
  assign s_csamul_cla32_and4_0 = a[4] & b[0];
  assign s_csamul_cla32_and5_0 = a[5] & b[0];
  assign s_csamul_cla32_and6_0 = a[6] & b[0];
  assign s_csamul_cla32_and7_0 = a[7] & b[0];
  assign s_csamul_cla32_and8_0 = a[8] & b[0];
  assign s_csamul_cla32_and9_0 = a[9] & b[0];
  assign s_csamul_cla32_and10_0 = a[10] & b[0];
  assign s_csamul_cla32_and11_0 = a[11] & b[0];
  assign s_csamul_cla32_and12_0 = a[12] & b[0];
  assign s_csamul_cla32_and13_0 = a[13] & b[0];
  assign s_csamul_cla32_and14_0 = a[14] & b[0];
  assign s_csamul_cla32_and15_0 = a[15] & b[0];
  assign s_csamul_cla32_and16_0 = a[16] & b[0];
  assign s_csamul_cla32_and17_0 = a[17] & b[0];
  assign s_csamul_cla32_and18_0 = a[18] & b[0];
  assign s_csamul_cla32_and19_0 = a[19] & b[0];
  assign s_csamul_cla32_and20_0 = a[20] & b[0];
  assign s_csamul_cla32_and21_0 = a[21] & b[0];
  assign s_csamul_cla32_and22_0 = a[22] & b[0];
  assign s_csamul_cla32_and23_0 = a[23] & b[0];
  assign s_csamul_cla32_and24_0 = a[24] & b[0];
  assign s_csamul_cla32_and25_0 = a[25] & b[0];
  assign s_csamul_cla32_and26_0 = a[26] & b[0];
  assign s_csamul_cla32_and27_0 = a[27] & b[0];
  assign s_csamul_cla32_and28_0 = a[28] & b[0];
  assign s_csamul_cla32_and29_0 = a[29] & b[0];
  assign s_csamul_cla32_and30_0 = a[30] & b[0];
  assign s_csamul_cla32_nand31_0 = ~(a[31] & b[0]);
  assign s_csamul_cla32_and0_1 = a[0] & b[1];
  assign s_csamul_cla32_ha0_1_xor0 = s_csamul_cla32_and0_1 ^ s_csamul_cla32_and1_0;
  assign s_csamul_cla32_ha0_1_and0 = s_csamul_cla32_and0_1 & s_csamul_cla32_and1_0;
  assign s_csamul_cla32_and1_1 = a[1] & b[1];
  assign s_csamul_cla32_ha1_1_xor0 = s_csamul_cla32_and1_1 ^ s_csamul_cla32_and2_0;
  assign s_csamul_cla32_ha1_1_and0 = s_csamul_cla32_and1_1 & s_csamul_cla32_and2_0;
  assign s_csamul_cla32_and2_1 = a[2] & b[1];
  assign s_csamul_cla32_ha2_1_xor0 = s_csamul_cla32_and2_1 ^ s_csamul_cla32_and3_0;
  assign s_csamul_cla32_ha2_1_and0 = s_csamul_cla32_and2_1 & s_csamul_cla32_and3_0;
  assign s_csamul_cla32_and3_1 = a[3] & b[1];
  assign s_csamul_cla32_ha3_1_xor0 = s_csamul_cla32_and3_1 ^ s_csamul_cla32_and4_0;
  assign s_csamul_cla32_ha3_1_and0 = s_csamul_cla32_and3_1 & s_csamul_cla32_and4_0;
  assign s_csamul_cla32_and4_1 = a[4] & b[1];
  assign s_csamul_cla32_ha4_1_xor0 = s_csamul_cla32_and4_1 ^ s_csamul_cla32_and5_0;
  assign s_csamul_cla32_ha4_1_and0 = s_csamul_cla32_and4_1 & s_csamul_cla32_and5_0;
  assign s_csamul_cla32_and5_1 = a[5] & b[1];
  assign s_csamul_cla32_ha5_1_xor0 = s_csamul_cla32_and5_1 ^ s_csamul_cla32_and6_0;
  assign s_csamul_cla32_ha5_1_and0 = s_csamul_cla32_and5_1 & s_csamul_cla32_and6_0;
  assign s_csamul_cla32_and6_1 = a[6] & b[1];
  assign s_csamul_cla32_ha6_1_xor0 = s_csamul_cla32_and6_1 ^ s_csamul_cla32_and7_0;
  assign s_csamul_cla32_ha6_1_and0 = s_csamul_cla32_and6_1 & s_csamul_cla32_and7_0;
  assign s_csamul_cla32_and7_1 = a[7] & b[1];
  assign s_csamul_cla32_ha7_1_xor0 = s_csamul_cla32_and7_1 ^ s_csamul_cla32_and8_0;
  assign s_csamul_cla32_ha7_1_and0 = s_csamul_cla32_and7_1 & s_csamul_cla32_and8_0;
  assign s_csamul_cla32_and8_1 = a[8] & b[1];
  assign s_csamul_cla32_ha8_1_xor0 = s_csamul_cla32_and8_1 ^ s_csamul_cla32_and9_0;
  assign s_csamul_cla32_ha8_1_and0 = s_csamul_cla32_and8_1 & s_csamul_cla32_and9_0;
  assign s_csamul_cla32_and9_1 = a[9] & b[1];
  assign s_csamul_cla32_ha9_1_xor0 = s_csamul_cla32_and9_1 ^ s_csamul_cla32_and10_0;
  assign s_csamul_cla32_ha9_1_and0 = s_csamul_cla32_and9_1 & s_csamul_cla32_and10_0;
  assign s_csamul_cla32_and10_1 = a[10] & b[1];
  assign s_csamul_cla32_ha10_1_xor0 = s_csamul_cla32_and10_1 ^ s_csamul_cla32_and11_0;
  assign s_csamul_cla32_ha10_1_and0 = s_csamul_cla32_and10_1 & s_csamul_cla32_and11_0;
  assign s_csamul_cla32_and11_1 = a[11] & b[1];
  assign s_csamul_cla32_ha11_1_xor0 = s_csamul_cla32_and11_1 ^ s_csamul_cla32_and12_0;
  assign s_csamul_cla32_ha11_1_and0 = s_csamul_cla32_and11_1 & s_csamul_cla32_and12_0;
  assign s_csamul_cla32_and12_1 = a[12] & b[1];
  assign s_csamul_cla32_ha12_1_xor0 = s_csamul_cla32_and12_1 ^ s_csamul_cla32_and13_0;
  assign s_csamul_cla32_ha12_1_and0 = s_csamul_cla32_and12_1 & s_csamul_cla32_and13_0;
  assign s_csamul_cla32_and13_1 = a[13] & b[1];
  assign s_csamul_cla32_ha13_1_xor0 = s_csamul_cla32_and13_1 ^ s_csamul_cla32_and14_0;
  assign s_csamul_cla32_ha13_1_and0 = s_csamul_cla32_and13_1 & s_csamul_cla32_and14_0;
  assign s_csamul_cla32_and14_1 = a[14] & b[1];
  assign s_csamul_cla32_ha14_1_xor0 = s_csamul_cla32_and14_1 ^ s_csamul_cla32_and15_0;
  assign s_csamul_cla32_ha14_1_and0 = s_csamul_cla32_and14_1 & s_csamul_cla32_and15_0;
  assign s_csamul_cla32_and15_1 = a[15] & b[1];
  assign s_csamul_cla32_ha15_1_xor0 = s_csamul_cla32_and15_1 ^ s_csamul_cla32_and16_0;
  assign s_csamul_cla32_ha15_1_and0 = s_csamul_cla32_and15_1 & s_csamul_cla32_and16_0;
  assign s_csamul_cla32_and16_1 = a[16] & b[1];
  assign s_csamul_cla32_ha16_1_xor0 = s_csamul_cla32_and16_1 ^ s_csamul_cla32_and17_0;
  assign s_csamul_cla32_ha16_1_and0 = s_csamul_cla32_and16_1 & s_csamul_cla32_and17_0;
  assign s_csamul_cla32_and17_1 = a[17] & b[1];
  assign s_csamul_cla32_ha17_1_xor0 = s_csamul_cla32_and17_1 ^ s_csamul_cla32_and18_0;
  assign s_csamul_cla32_ha17_1_and0 = s_csamul_cla32_and17_1 & s_csamul_cla32_and18_0;
  assign s_csamul_cla32_and18_1 = a[18] & b[1];
  assign s_csamul_cla32_ha18_1_xor0 = s_csamul_cla32_and18_1 ^ s_csamul_cla32_and19_0;
  assign s_csamul_cla32_ha18_1_and0 = s_csamul_cla32_and18_1 & s_csamul_cla32_and19_0;
  assign s_csamul_cla32_and19_1 = a[19] & b[1];
  assign s_csamul_cla32_ha19_1_xor0 = s_csamul_cla32_and19_1 ^ s_csamul_cla32_and20_0;
  assign s_csamul_cla32_ha19_1_and0 = s_csamul_cla32_and19_1 & s_csamul_cla32_and20_0;
  assign s_csamul_cla32_and20_1 = a[20] & b[1];
  assign s_csamul_cla32_ha20_1_xor0 = s_csamul_cla32_and20_1 ^ s_csamul_cla32_and21_0;
  assign s_csamul_cla32_ha20_1_and0 = s_csamul_cla32_and20_1 & s_csamul_cla32_and21_0;
  assign s_csamul_cla32_and21_1 = a[21] & b[1];
  assign s_csamul_cla32_ha21_1_xor0 = s_csamul_cla32_and21_1 ^ s_csamul_cla32_and22_0;
  assign s_csamul_cla32_ha21_1_and0 = s_csamul_cla32_and21_1 & s_csamul_cla32_and22_0;
  assign s_csamul_cla32_and22_1 = a[22] & b[1];
  assign s_csamul_cla32_ha22_1_xor0 = s_csamul_cla32_and22_1 ^ s_csamul_cla32_and23_0;
  assign s_csamul_cla32_ha22_1_and0 = s_csamul_cla32_and22_1 & s_csamul_cla32_and23_0;
  assign s_csamul_cla32_and23_1 = a[23] & b[1];
  assign s_csamul_cla32_ha23_1_xor0 = s_csamul_cla32_and23_1 ^ s_csamul_cla32_and24_0;
  assign s_csamul_cla32_ha23_1_and0 = s_csamul_cla32_and23_1 & s_csamul_cla32_and24_0;
  assign s_csamul_cla32_and24_1 = a[24] & b[1];
  assign s_csamul_cla32_ha24_1_xor0 = s_csamul_cla32_and24_1 ^ s_csamul_cla32_and25_0;
  assign s_csamul_cla32_ha24_1_and0 = s_csamul_cla32_and24_1 & s_csamul_cla32_and25_0;
  assign s_csamul_cla32_and25_1 = a[25] & b[1];
  assign s_csamul_cla32_ha25_1_xor0 = s_csamul_cla32_and25_1 ^ s_csamul_cla32_and26_0;
  assign s_csamul_cla32_ha25_1_and0 = s_csamul_cla32_and25_1 & s_csamul_cla32_and26_0;
  assign s_csamul_cla32_and26_1 = a[26] & b[1];
  assign s_csamul_cla32_ha26_1_xor0 = s_csamul_cla32_and26_1 ^ s_csamul_cla32_and27_0;
  assign s_csamul_cla32_ha26_1_and0 = s_csamul_cla32_and26_1 & s_csamul_cla32_and27_0;
  assign s_csamul_cla32_and27_1 = a[27] & b[1];
  assign s_csamul_cla32_ha27_1_xor0 = s_csamul_cla32_and27_1 ^ s_csamul_cla32_and28_0;
  assign s_csamul_cla32_ha27_1_and0 = s_csamul_cla32_and27_1 & s_csamul_cla32_and28_0;
  assign s_csamul_cla32_and28_1 = a[28] & b[1];
  assign s_csamul_cla32_ha28_1_xor0 = s_csamul_cla32_and28_1 ^ s_csamul_cla32_and29_0;
  assign s_csamul_cla32_ha28_1_and0 = s_csamul_cla32_and28_1 & s_csamul_cla32_and29_0;
  assign s_csamul_cla32_and29_1 = a[29] & b[1];
  assign s_csamul_cla32_ha29_1_xor0 = s_csamul_cla32_and29_1 ^ s_csamul_cla32_and30_0;
  assign s_csamul_cla32_ha29_1_and0 = s_csamul_cla32_and29_1 & s_csamul_cla32_and30_0;
  assign s_csamul_cla32_and30_1 = a[30] & b[1];
  assign s_csamul_cla32_ha30_1_xor0 = s_csamul_cla32_and30_1 ^ s_csamul_cla32_nand31_0;
  assign s_csamul_cla32_ha30_1_and0 = s_csamul_cla32_and30_1 & s_csamul_cla32_nand31_0;
  assign s_csamul_cla32_nand31_1 = ~(a[31] & b[1]);
  assign s_csamul_cla32_ha31_1_xor0 = ~s_csamul_cla32_nand31_1;
  assign s_csamul_cla32_and0_2 = a[0] & b[2];
  assign s_csamul_cla32_fa0_2_xor0 = s_csamul_cla32_and0_2 ^ s_csamul_cla32_ha1_1_xor0;
  assign s_csamul_cla32_fa0_2_and0 = s_csamul_cla32_and0_2 & s_csamul_cla32_ha1_1_xor0;
  assign s_csamul_cla32_fa0_2_xor1 = s_csamul_cla32_fa0_2_xor0 ^ s_csamul_cla32_ha0_1_and0;
  assign s_csamul_cla32_fa0_2_and1 = s_csamul_cla32_fa0_2_xor0 & s_csamul_cla32_ha0_1_and0;
  assign s_csamul_cla32_fa0_2_or0 = s_csamul_cla32_fa0_2_and0 | s_csamul_cla32_fa0_2_and1;
  assign s_csamul_cla32_and1_2 = a[1] & b[2];
  assign s_csamul_cla32_fa1_2_xor0 = s_csamul_cla32_and1_2 ^ s_csamul_cla32_ha2_1_xor0;
  assign s_csamul_cla32_fa1_2_and0 = s_csamul_cla32_and1_2 & s_csamul_cla32_ha2_1_xor0;
  assign s_csamul_cla32_fa1_2_xor1 = s_csamul_cla32_fa1_2_xor0 ^ s_csamul_cla32_ha1_1_and0;
  assign s_csamul_cla32_fa1_2_and1 = s_csamul_cla32_fa1_2_xor0 & s_csamul_cla32_ha1_1_and0;
  assign s_csamul_cla32_fa1_2_or0 = s_csamul_cla32_fa1_2_and0 | s_csamul_cla32_fa1_2_and1;
  assign s_csamul_cla32_and2_2 = a[2] & b[2];
  assign s_csamul_cla32_fa2_2_xor0 = s_csamul_cla32_and2_2 ^ s_csamul_cla32_ha3_1_xor0;
  assign s_csamul_cla32_fa2_2_and0 = s_csamul_cla32_and2_2 & s_csamul_cla32_ha3_1_xor0;
  assign s_csamul_cla32_fa2_2_xor1 = s_csamul_cla32_fa2_2_xor0 ^ s_csamul_cla32_ha2_1_and0;
  assign s_csamul_cla32_fa2_2_and1 = s_csamul_cla32_fa2_2_xor0 & s_csamul_cla32_ha2_1_and0;
  assign s_csamul_cla32_fa2_2_or0 = s_csamul_cla32_fa2_2_and0 | s_csamul_cla32_fa2_2_and1;
  assign s_csamul_cla32_and3_2 = a[3] & b[2];
  assign s_csamul_cla32_fa3_2_xor0 = s_csamul_cla32_and3_2 ^ s_csamul_cla32_ha4_1_xor0;
  assign s_csamul_cla32_fa3_2_and0 = s_csamul_cla32_and3_2 & s_csamul_cla32_ha4_1_xor0;
  assign s_csamul_cla32_fa3_2_xor1 = s_csamul_cla32_fa3_2_xor0 ^ s_csamul_cla32_ha3_1_and0;
  assign s_csamul_cla32_fa3_2_and1 = s_csamul_cla32_fa3_2_xor0 & s_csamul_cla32_ha3_1_and0;
  assign s_csamul_cla32_fa3_2_or0 = s_csamul_cla32_fa3_2_and0 | s_csamul_cla32_fa3_2_and1;
  assign s_csamul_cla32_and4_2 = a[4] & b[2];
  assign s_csamul_cla32_fa4_2_xor0 = s_csamul_cla32_and4_2 ^ s_csamul_cla32_ha5_1_xor0;
  assign s_csamul_cla32_fa4_2_and0 = s_csamul_cla32_and4_2 & s_csamul_cla32_ha5_1_xor0;
  assign s_csamul_cla32_fa4_2_xor1 = s_csamul_cla32_fa4_2_xor0 ^ s_csamul_cla32_ha4_1_and0;
  assign s_csamul_cla32_fa4_2_and1 = s_csamul_cla32_fa4_2_xor0 & s_csamul_cla32_ha4_1_and0;
  assign s_csamul_cla32_fa4_2_or0 = s_csamul_cla32_fa4_2_and0 | s_csamul_cla32_fa4_2_and1;
  assign s_csamul_cla32_and5_2 = a[5] & b[2];
  assign s_csamul_cla32_fa5_2_xor0 = s_csamul_cla32_and5_2 ^ s_csamul_cla32_ha6_1_xor0;
  assign s_csamul_cla32_fa5_2_and0 = s_csamul_cla32_and5_2 & s_csamul_cla32_ha6_1_xor0;
  assign s_csamul_cla32_fa5_2_xor1 = s_csamul_cla32_fa5_2_xor0 ^ s_csamul_cla32_ha5_1_and0;
  assign s_csamul_cla32_fa5_2_and1 = s_csamul_cla32_fa5_2_xor0 & s_csamul_cla32_ha5_1_and0;
  assign s_csamul_cla32_fa5_2_or0 = s_csamul_cla32_fa5_2_and0 | s_csamul_cla32_fa5_2_and1;
  assign s_csamul_cla32_and6_2 = a[6] & b[2];
  assign s_csamul_cla32_fa6_2_xor0 = s_csamul_cla32_and6_2 ^ s_csamul_cla32_ha7_1_xor0;
  assign s_csamul_cla32_fa6_2_and0 = s_csamul_cla32_and6_2 & s_csamul_cla32_ha7_1_xor0;
  assign s_csamul_cla32_fa6_2_xor1 = s_csamul_cla32_fa6_2_xor0 ^ s_csamul_cla32_ha6_1_and0;
  assign s_csamul_cla32_fa6_2_and1 = s_csamul_cla32_fa6_2_xor0 & s_csamul_cla32_ha6_1_and0;
  assign s_csamul_cla32_fa6_2_or0 = s_csamul_cla32_fa6_2_and0 | s_csamul_cla32_fa6_2_and1;
  assign s_csamul_cla32_and7_2 = a[7] & b[2];
  assign s_csamul_cla32_fa7_2_xor0 = s_csamul_cla32_and7_2 ^ s_csamul_cla32_ha8_1_xor0;
  assign s_csamul_cla32_fa7_2_and0 = s_csamul_cla32_and7_2 & s_csamul_cla32_ha8_1_xor0;
  assign s_csamul_cla32_fa7_2_xor1 = s_csamul_cla32_fa7_2_xor0 ^ s_csamul_cla32_ha7_1_and0;
  assign s_csamul_cla32_fa7_2_and1 = s_csamul_cla32_fa7_2_xor0 & s_csamul_cla32_ha7_1_and0;
  assign s_csamul_cla32_fa7_2_or0 = s_csamul_cla32_fa7_2_and0 | s_csamul_cla32_fa7_2_and1;
  assign s_csamul_cla32_and8_2 = a[8] & b[2];
  assign s_csamul_cla32_fa8_2_xor0 = s_csamul_cla32_and8_2 ^ s_csamul_cla32_ha9_1_xor0;
  assign s_csamul_cla32_fa8_2_and0 = s_csamul_cla32_and8_2 & s_csamul_cla32_ha9_1_xor0;
  assign s_csamul_cla32_fa8_2_xor1 = s_csamul_cla32_fa8_2_xor0 ^ s_csamul_cla32_ha8_1_and0;
  assign s_csamul_cla32_fa8_2_and1 = s_csamul_cla32_fa8_2_xor0 & s_csamul_cla32_ha8_1_and0;
  assign s_csamul_cla32_fa8_2_or0 = s_csamul_cla32_fa8_2_and0 | s_csamul_cla32_fa8_2_and1;
  assign s_csamul_cla32_and9_2 = a[9] & b[2];
  assign s_csamul_cla32_fa9_2_xor0 = s_csamul_cla32_and9_2 ^ s_csamul_cla32_ha10_1_xor0;
  assign s_csamul_cla32_fa9_2_and0 = s_csamul_cla32_and9_2 & s_csamul_cla32_ha10_1_xor0;
  assign s_csamul_cla32_fa9_2_xor1 = s_csamul_cla32_fa9_2_xor0 ^ s_csamul_cla32_ha9_1_and0;
  assign s_csamul_cla32_fa9_2_and1 = s_csamul_cla32_fa9_2_xor0 & s_csamul_cla32_ha9_1_and0;
  assign s_csamul_cla32_fa9_2_or0 = s_csamul_cla32_fa9_2_and0 | s_csamul_cla32_fa9_2_and1;
  assign s_csamul_cla32_and10_2 = a[10] & b[2];
  assign s_csamul_cla32_fa10_2_xor0 = s_csamul_cla32_and10_2 ^ s_csamul_cla32_ha11_1_xor0;
  assign s_csamul_cla32_fa10_2_and0 = s_csamul_cla32_and10_2 & s_csamul_cla32_ha11_1_xor0;
  assign s_csamul_cla32_fa10_2_xor1 = s_csamul_cla32_fa10_2_xor0 ^ s_csamul_cla32_ha10_1_and0;
  assign s_csamul_cla32_fa10_2_and1 = s_csamul_cla32_fa10_2_xor0 & s_csamul_cla32_ha10_1_and0;
  assign s_csamul_cla32_fa10_2_or0 = s_csamul_cla32_fa10_2_and0 | s_csamul_cla32_fa10_2_and1;
  assign s_csamul_cla32_and11_2 = a[11] & b[2];
  assign s_csamul_cla32_fa11_2_xor0 = s_csamul_cla32_and11_2 ^ s_csamul_cla32_ha12_1_xor0;
  assign s_csamul_cla32_fa11_2_and0 = s_csamul_cla32_and11_2 & s_csamul_cla32_ha12_1_xor0;
  assign s_csamul_cla32_fa11_2_xor1 = s_csamul_cla32_fa11_2_xor0 ^ s_csamul_cla32_ha11_1_and0;
  assign s_csamul_cla32_fa11_2_and1 = s_csamul_cla32_fa11_2_xor0 & s_csamul_cla32_ha11_1_and0;
  assign s_csamul_cla32_fa11_2_or0 = s_csamul_cla32_fa11_2_and0 | s_csamul_cla32_fa11_2_and1;
  assign s_csamul_cla32_and12_2 = a[12] & b[2];
  assign s_csamul_cla32_fa12_2_xor0 = s_csamul_cla32_and12_2 ^ s_csamul_cla32_ha13_1_xor0;
  assign s_csamul_cla32_fa12_2_and0 = s_csamul_cla32_and12_2 & s_csamul_cla32_ha13_1_xor0;
  assign s_csamul_cla32_fa12_2_xor1 = s_csamul_cla32_fa12_2_xor0 ^ s_csamul_cla32_ha12_1_and0;
  assign s_csamul_cla32_fa12_2_and1 = s_csamul_cla32_fa12_2_xor0 & s_csamul_cla32_ha12_1_and0;
  assign s_csamul_cla32_fa12_2_or0 = s_csamul_cla32_fa12_2_and0 | s_csamul_cla32_fa12_2_and1;
  assign s_csamul_cla32_and13_2 = a[13] & b[2];
  assign s_csamul_cla32_fa13_2_xor0 = s_csamul_cla32_and13_2 ^ s_csamul_cla32_ha14_1_xor0;
  assign s_csamul_cla32_fa13_2_and0 = s_csamul_cla32_and13_2 & s_csamul_cla32_ha14_1_xor0;
  assign s_csamul_cla32_fa13_2_xor1 = s_csamul_cla32_fa13_2_xor0 ^ s_csamul_cla32_ha13_1_and0;
  assign s_csamul_cla32_fa13_2_and1 = s_csamul_cla32_fa13_2_xor0 & s_csamul_cla32_ha13_1_and0;
  assign s_csamul_cla32_fa13_2_or0 = s_csamul_cla32_fa13_2_and0 | s_csamul_cla32_fa13_2_and1;
  assign s_csamul_cla32_and14_2 = a[14] & b[2];
  assign s_csamul_cla32_fa14_2_xor0 = s_csamul_cla32_and14_2 ^ s_csamul_cla32_ha15_1_xor0;
  assign s_csamul_cla32_fa14_2_and0 = s_csamul_cla32_and14_2 & s_csamul_cla32_ha15_1_xor0;
  assign s_csamul_cla32_fa14_2_xor1 = s_csamul_cla32_fa14_2_xor0 ^ s_csamul_cla32_ha14_1_and0;
  assign s_csamul_cla32_fa14_2_and1 = s_csamul_cla32_fa14_2_xor0 & s_csamul_cla32_ha14_1_and0;
  assign s_csamul_cla32_fa14_2_or0 = s_csamul_cla32_fa14_2_and0 | s_csamul_cla32_fa14_2_and1;
  assign s_csamul_cla32_and15_2 = a[15] & b[2];
  assign s_csamul_cla32_fa15_2_xor0 = s_csamul_cla32_and15_2 ^ s_csamul_cla32_ha16_1_xor0;
  assign s_csamul_cla32_fa15_2_and0 = s_csamul_cla32_and15_2 & s_csamul_cla32_ha16_1_xor0;
  assign s_csamul_cla32_fa15_2_xor1 = s_csamul_cla32_fa15_2_xor0 ^ s_csamul_cla32_ha15_1_and0;
  assign s_csamul_cla32_fa15_2_and1 = s_csamul_cla32_fa15_2_xor0 & s_csamul_cla32_ha15_1_and0;
  assign s_csamul_cla32_fa15_2_or0 = s_csamul_cla32_fa15_2_and0 | s_csamul_cla32_fa15_2_and1;
  assign s_csamul_cla32_and16_2 = a[16] & b[2];
  assign s_csamul_cla32_fa16_2_xor0 = s_csamul_cla32_and16_2 ^ s_csamul_cla32_ha17_1_xor0;
  assign s_csamul_cla32_fa16_2_and0 = s_csamul_cla32_and16_2 & s_csamul_cla32_ha17_1_xor0;
  assign s_csamul_cla32_fa16_2_xor1 = s_csamul_cla32_fa16_2_xor0 ^ s_csamul_cla32_ha16_1_and0;
  assign s_csamul_cla32_fa16_2_and1 = s_csamul_cla32_fa16_2_xor0 & s_csamul_cla32_ha16_1_and0;
  assign s_csamul_cla32_fa16_2_or0 = s_csamul_cla32_fa16_2_and0 | s_csamul_cla32_fa16_2_and1;
  assign s_csamul_cla32_and17_2 = a[17] & b[2];
  assign s_csamul_cla32_fa17_2_xor0 = s_csamul_cla32_and17_2 ^ s_csamul_cla32_ha18_1_xor0;
  assign s_csamul_cla32_fa17_2_and0 = s_csamul_cla32_and17_2 & s_csamul_cla32_ha18_1_xor0;
  assign s_csamul_cla32_fa17_2_xor1 = s_csamul_cla32_fa17_2_xor0 ^ s_csamul_cla32_ha17_1_and0;
  assign s_csamul_cla32_fa17_2_and1 = s_csamul_cla32_fa17_2_xor0 & s_csamul_cla32_ha17_1_and0;
  assign s_csamul_cla32_fa17_2_or0 = s_csamul_cla32_fa17_2_and0 | s_csamul_cla32_fa17_2_and1;
  assign s_csamul_cla32_and18_2 = a[18] & b[2];
  assign s_csamul_cla32_fa18_2_xor0 = s_csamul_cla32_and18_2 ^ s_csamul_cla32_ha19_1_xor0;
  assign s_csamul_cla32_fa18_2_and0 = s_csamul_cla32_and18_2 & s_csamul_cla32_ha19_1_xor0;
  assign s_csamul_cla32_fa18_2_xor1 = s_csamul_cla32_fa18_2_xor0 ^ s_csamul_cla32_ha18_1_and0;
  assign s_csamul_cla32_fa18_2_and1 = s_csamul_cla32_fa18_2_xor0 & s_csamul_cla32_ha18_1_and0;
  assign s_csamul_cla32_fa18_2_or0 = s_csamul_cla32_fa18_2_and0 | s_csamul_cla32_fa18_2_and1;
  assign s_csamul_cla32_and19_2 = a[19] & b[2];
  assign s_csamul_cla32_fa19_2_xor0 = s_csamul_cla32_and19_2 ^ s_csamul_cla32_ha20_1_xor0;
  assign s_csamul_cla32_fa19_2_and0 = s_csamul_cla32_and19_2 & s_csamul_cla32_ha20_1_xor0;
  assign s_csamul_cla32_fa19_2_xor1 = s_csamul_cla32_fa19_2_xor0 ^ s_csamul_cla32_ha19_1_and0;
  assign s_csamul_cla32_fa19_2_and1 = s_csamul_cla32_fa19_2_xor0 & s_csamul_cla32_ha19_1_and0;
  assign s_csamul_cla32_fa19_2_or0 = s_csamul_cla32_fa19_2_and0 | s_csamul_cla32_fa19_2_and1;
  assign s_csamul_cla32_and20_2 = a[20] & b[2];
  assign s_csamul_cla32_fa20_2_xor0 = s_csamul_cla32_and20_2 ^ s_csamul_cla32_ha21_1_xor0;
  assign s_csamul_cla32_fa20_2_and0 = s_csamul_cla32_and20_2 & s_csamul_cla32_ha21_1_xor0;
  assign s_csamul_cla32_fa20_2_xor1 = s_csamul_cla32_fa20_2_xor0 ^ s_csamul_cla32_ha20_1_and0;
  assign s_csamul_cla32_fa20_2_and1 = s_csamul_cla32_fa20_2_xor0 & s_csamul_cla32_ha20_1_and0;
  assign s_csamul_cla32_fa20_2_or0 = s_csamul_cla32_fa20_2_and0 | s_csamul_cla32_fa20_2_and1;
  assign s_csamul_cla32_and21_2 = a[21] & b[2];
  assign s_csamul_cla32_fa21_2_xor0 = s_csamul_cla32_and21_2 ^ s_csamul_cla32_ha22_1_xor0;
  assign s_csamul_cla32_fa21_2_and0 = s_csamul_cla32_and21_2 & s_csamul_cla32_ha22_1_xor0;
  assign s_csamul_cla32_fa21_2_xor1 = s_csamul_cla32_fa21_2_xor0 ^ s_csamul_cla32_ha21_1_and0;
  assign s_csamul_cla32_fa21_2_and1 = s_csamul_cla32_fa21_2_xor0 & s_csamul_cla32_ha21_1_and0;
  assign s_csamul_cla32_fa21_2_or0 = s_csamul_cla32_fa21_2_and0 | s_csamul_cla32_fa21_2_and1;
  assign s_csamul_cla32_and22_2 = a[22] & b[2];
  assign s_csamul_cla32_fa22_2_xor0 = s_csamul_cla32_and22_2 ^ s_csamul_cla32_ha23_1_xor0;
  assign s_csamul_cla32_fa22_2_and0 = s_csamul_cla32_and22_2 & s_csamul_cla32_ha23_1_xor0;
  assign s_csamul_cla32_fa22_2_xor1 = s_csamul_cla32_fa22_2_xor0 ^ s_csamul_cla32_ha22_1_and0;
  assign s_csamul_cla32_fa22_2_and1 = s_csamul_cla32_fa22_2_xor0 & s_csamul_cla32_ha22_1_and0;
  assign s_csamul_cla32_fa22_2_or0 = s_csamul_cla32_fa22_2_and0 | s_csamul_cla32_fa22_2_and1;
  assign s_csamul_cla32_and23_2 = a[23] & b[2];
  assign s_csamul_cla32_fa23_2_xor0 = s_csamul_cla32_and23_2 ^ s_csamul_cla32_ha24_1_xor0;
  assign s_csamul_cla32_fa23_2_and0 = s_csamul_cla32_and23_2 & s_csamul_cla32_ha24_1_xor0;
  assign s_csamul_cla32_fa23_2_xor1 = s_csamul_cla32_fa23_2_xor0 ^ s_csamul_cla32_ha23_1_and0;
  assign s_csamul_cla32_fa23_2_and1 = s_csamul_cla32_fa23_2_xor0 & s_csamul_cla32_ha23_1_and0;
  assign s_csamul_cla32_fa23_2_or0 = s_csamul_cla32_fa23_2_and0 | s_csamul_cla32_fa23_2_and1;
  assign s_csamul_cla32_and24_2 = a[24] & b[2];
  assign s_csamul_cla32_fa24_2_xor0 = s_csamul_cla32_and24_2 ^ s_csamul_cla32_ha25_1_xor0;
  assign s_csamul_cla32_fa24_2_and0 = s_csamul_cla32_and24_2 & s_csamul_cla32_ha25_1_xor0;
  assign s_csamul_cla32_fa24_2_xor1 = s_csamul_cla32_fa24_2_xor0 ^ s_csamul_cla32_ha24_1_and0;
  assign s_csamul_cla32_fa24_2_and1 = s_csamul_cla32_fa24_2_xor0 & s_csamul_cla32_ha24_1_and0;
  assign s_csamul_cla32_fa24_2_or0 = s_csamul_cla32_fa24_2_and0 | s_csamul_cla32_fa24_2_and1;
  assign s_csamul_cla32_and25_2 = a[25] & b[2];
  assign s_csamul_cla32_fa25_2_xor0 = s_csamul_cla32_and25_2 ^ s_csamul_cla32_ha26_1_xor0;
  assign s_csamul_cla32_fa25_2_and0 = s_csamul_cla32_and25_2 & s_csamul_cla32_ha26_1_xor0;
  assign s_csamul_cla32_fa25_2_xor1 = s_csamul_cla32_fa25_2_xor0 ^ s_csamul_cla32_ha25_1_and0;
  assign s_csamul_cla32_fa25_2_and1 = s_csamul_cla32_fa25_2_xor0 & s_csamul_cla32_ha25_1_and0;
  assign s_csamul_cla32_fa25_2_or0 = s_csamul_cla32_fa25_2_and0 | s_csamul_cla32_fa25_2_and1;
  assign s_csamul_cla32_and26_2 = a[26] & b[2];
  assign s_csamul_cla32_fa26_2_xor0 = s_csamul_cla32_and26_2 ^ s_csamul_cla32_ha27_1_xor0;
  assign s_csamul_cla32_fa26_2_and0 = s_csamul_cla32_and26_2 & s_csamul_cla32_ha27_1_xor0;
  assign s_csamul_cla32_fa26_2_xor1 = s_csamul_cla32_fa26_2_xor0 ^ s_csamul_cla32_ha26_1_and0;
  assign s_csamul_cla32_fa26_2_and1 = s_csamul_cla32_fa26_2_xor0 & s_csamul_cla32_ha26_1_and0;
  assign s_csamul_cla32_fa26_2_or0 = s_csamul_cla32_fa26_2_and0 | s_csamul_cla32_fa26_2_and1;
  assign s_csamul_cla32_and27_2 = a[27] & b[2];
  assign s_csamul_cla32_fa27_2_xor0 = s_csamul_cla32_and27_2 ^ s_csamul_cla32_ha28_1_xor0;
  assign s_csamul_cla32_fa27_2_and0 = s_csamul_cla32_and27_2 & s_csamul_cla32_ha28_1_xor0;
  assign s_csamul_cla32_fa27_2_xor1 = s_csamul_cla32_fa27_2_xor0 ^ s_csamul_cla32_ha27_1_and0;
  assign s_csamul_cla32_fa27_2_and1 = s_csamul_cla32_fa27_2_xor0 & s_csamul_cla32_ha27_1_and0;
  assign s_csamul_cla32_fa27_2_or0 = s_csamul_cla32_fa27_2_and0 | s_csamul_cla32_fa27_2_and1;
  assign s_csamul_cla32_and28_2 = a[28] & b[2];
  assign s_csamul_cla32_fa28_2_xor0 = s_csamul_cla32_and28_2 ^ s_csamul_cla32_ha29_1_xor0;
  assign s_csamul_cla32_fa28_2_and0 = s_csamul_cla32_and28_2 & s_csamul_cla32_ha29_1_xor0;
  assign s_csamul_cla32_fa28_2_xor1 = s_csamul_cla32_fa28_2_xor0 ^ s_csamul_cla32_ha28_1_and0;
  assign s_csamul_cla32_fa28_2_and1 = s_csamul_cla32_fa28_2_xor0 & s_csamul_cla32_ha28_1_and0;
  assign s_csamul_cla32_fa28_2_or0 = s_csamul_cla32_fa28_2_and0 | s_csamul_cla32_fa28_2_and1;
  assign s_csamul_cla32_and29_2 = a[29] & b[2];
  assign s_csamul_cla32_fa29_2_xor0 = s_csamul_cla32_and29_2 ^ s_csamul_cla32_ha30_1_xor0;
  assign s_csamul_cla32_fa29_2_and0 = s_csamul_cla32_and29_2 & s_csamul_cla32_ha30_1_xor0;
  assign s_csamul_cla32_fa29_2_xor1 = s_csamul_cla32_fa29_2_xor0 ^ s_csamul_cla32_ha29_1_and0;
  assign s_csamul_cla32_fa29_2_and1 = s_csamul_cla32_fa29_2_xor0 & s_csamul_cla32_ha29_1_and0;
  assign s_csamul_cla32_fa29_2_or0 = s_csamul_cla32_fa29_2_and0 | s_csamul_cla32_fa29_2_and1;
  assign s_csamul_cla32_and30_2 = a[30] & b[2];
  assign s_csamul_cla32_fa30_2_xor0 = s_csamul_cla32_and30_2 ^ s_csamul_cla32_ha31_1_xor0;
  assign s_csamul_cla32_fa30_2_and0 = s_csamul_cla32_and30_2 & s_csamul_cla32_ha31_1_xor0;
  assign s_csamul_cla32_fa30_2_xor1 = s_csamul_cla32_fa30_2_xor0 ^ s_csamul_cla32_ha30_1_and0;
  assign s_csamul_cla32_fa30_2_and1 = s_csamul_cla32_fa30_2_xor0 & s_csamul_cla32_ha30_1_and0;
  assign s_csamul_cla32_fa30_2_or0 = s_csamul_cla32_fa30_2_and0 | s_csamul_cla32_fa30_2_and1;
  assign s_csamul_cla32_nand31_2 = ~(a[31] & b[2]);
  assign s_csamul_cla32_ha31_2_xor0 = s_csamul_cla32_nand31_2 ^ s_csamul_cla32_nand31_1;
  assign s_csamul_cla32_ha31_2_and0 = s_csamul_cla32_nand31_2 & s_csamul_cla32_nand31_1;
  assign s_csamul_cla32_and0_3 = a[0] & b[3];
  assign s_csamul_cla32_fa0_3_xor0 = s_csamul_cla32_and0_3 ^ s_csamul_cla32_fa1_2_xor1;
  assign s_csamul_cla32_fa0_3_and0 = s_csamul_cla32_and0_3 & s_csamul_cla32_fa1_2_xor1;
  assign s_csamul_cla32_fa0_3_xor1 = s_csamul_cla32_fa0_3_xor0 ^ s_csamul_cla32_fa0_2_or0;
  assign s_csamul_cla32_fa0_3_and1 = s_csamul_cla32_fa0_3_xor0 & s_csamul_cla32_fa0_2_or0;
  assign s_csamul_cla32_fa0_3_or0 = s_csamul_cla32_fa0_3_and0 | s_csamul_cla32_fa0_3_and1;
  assign s_csamul_cla32_and1_3 = a[1] & b[3];
  assign s_csamul_cla32_fa1_3_xor0 = s_csamul_cla32_and1_3 ^ s_csamul_cla32_fa2_2_xor1;
  assign s_csamul_cla32_fa1_3_and0 = s_csamul_cla32_and1_3 & s_csamul_cla32_fa2_2_xor1;
  assign s_csamul_cla32_fa1_3_xor1 = s_csamul_cla32_fa1_3_xor0 ^ s_csamul_cla32_fa1_2_or0;
  assign s_csamul_cla32_fa1_3_and1 = s_csamul_cla32_fa1_3_xor0 & s_csamul_cla32_fa1_2_or0;
  assign s_csamul_cla32_fa1_3_or0 = s_csamul_cla32_fa1_3_and0 | s_csamul_cla32_fa1_3_and1;
  assign s_csamul_cla32_and2_3 = a[2] & b[3];
  assign s_csamul_cla32_fa2_3_xor0 = s_csamul_cla32_and2_3 ^ s_csamul_cla32_fa3_2_xor1;
  assign s_csamul_cla32_fa2_3_and0 = s_csamul_cla32_and2_3 & s_csamul_cla32_fa3_2_xor1;
  assign s_csamul_cla32_fa2_3_xor1 = s_csamul_cla32_fa2_3_xor0 ^ s_csamul_cla32_fa2_2_or0;
  assign s_csamul_cla32_fa2_3_and1 = s_csamul_cla32_fa2_3_xor0 & s_csamul_cla32_fa2_2_or0;
  assign s_csamul_cla32_fa2_3_or0 = s_csamul_cla32_fa2_3_and0 | s_csamul_cla32_fa2_3_and1;
  assign s_csamul_cla32_and3_3 = a[3] & b[3];
  assign s_csamul_cla32_fa3_3_xor0 = s_csamul_cla32_and3_3 ^ s_csamul_cla32_fa4_2_xor1;
  assign s_csamul_cla32_fa3_3_and0 = s_csamul_cla32_and3_3 & s_csamul_cla32_fa4_2_xor1;
  assign s_csamul_cla32_fa3_3_xor1 = s_csamul_cla32_fa3_3_xor0 ^ s_csamul_cla32_fa3_2_or0;
  assign s_csamul_cla32_fa3_3_and1 = s_csamul_cla32_fa3_3_xor0 & s_csamul_cla32_fa3_2_or0;
  assign s_csamul_cla32_fa3_3_or0 = s_csamul_cla32_fa3_3_and0 | s_csamul_cla32_fa3_3_and1;
  assign s_csamul_cla32_and4_3 = a[4] & b[3];
  assign s_csamul_cla32_fa4_3_xor0 = s_csamul_cla32_and4_3 ^ s_csamul_cla32_fa5_2_xor1;
  assign s_csamul_cla32_fa4_3_and0 = s_csamul_cla32_and4_3 & s_csamul_cla32_fa5_2_xor1;
  assign s_csamul_cla32_fa4_3_xor1 = s_csamul_cla32_fa4_3_xor0 ^ s_csamul_cla32_fa4_2_or0;
  assign s_csamul_cla32_fa4_3_and1 = s_csamul_cla32_fa4_3_xor0 & s_csamul_cla32_fa4_2_or0;
  assign s_csamul_cla32_fa4_3_or0 = s_csamul_cla32_fa4_3_and0 | s_csamul_cla32_fa4_3_and1;
  assign s_csamul_cla32_and5_3 = a[5] & b[3];
  assign s_csamul_cla32_fa5_3_xor0 = s_csamul_cla32_and5_3 ^ s_csamul_cla32_fa6_2_xor1;
  assign s_csamul_cla32_fa5_3_and0 = s_csamul_cla32_and5_3 & s_csamul_cla32_fa6_2_xor1;
  assign s_csamul_cla32_fa5_3_xor1 = s_csamul_cla32_fa5_3_xor0 ^ s_csamul_cla32_fa5_2_or0;
  assign s_csamul_cla32_fa5_3_and1 = s_csamul_cla32_fa5_3_xor0 & s_csamul_cla32_fa5_2_or0;
  assign s_csamul_cla32_fa5_3_or0 = s_csamul_cla32_fa5_3_and0 | s_csamul_cla32_fa5_3_and1;
  assign s_csamul_cla32_and6_3 = a[6] & b[3];
  assign s_csamul_cla32_fa6_3_xor0 = s_csamul_cla32_and6_3 ^ s_csamul_cla32_fa7_2_xor1;
  assign s_csamul_cla32_fa6_3_and0 = s_csamul_cla32_and6_3 & s_csamul_cla32_fa7_2_xor1;
  assign s_csamul_cla32_fa6_3_xor1 = s_csamul_cla32_fa6_3_xor0 ^ s_csamul_cla32_fa6_2_or0;
  assign s_csamul_cla32_fa6_3_and1 = s_csamul_cla32_fa6_3_xor0 & s_csamul_cla32_fa6_2_or0;
  assign s_csamul_cla32_fa6_3_or0 = s_csamul_cla32_fa6_3_and0 | s_csamul_cla32_fa6_3_and1;
  assign s_csamul_cla32_and7_3 = a[7] & b[3];
  assign s_csamul_cla32_fa7_3_xor0 = s_csamul_cla32_and7_3 ^ s_csamul_cla32_fa8_2_xor1;
  assign s_csamul_cla32_fa7_3_and0 = s_csamul_cla32_and7_3 & s_csamul_cla32_fa8_2_xor1;
  assign s_csamul_cla32_fa7_3_xor1 = s_csamul_cla32_fa7_3_xor0 ^ s_csamul_cla32_fa7_2_or0;
  assign s_csamul_cla32_fa7_3_and1 = s_csamul_cla32_fa7_3_xor0 & s_csamul_cla32_fa7_2_or0;
  assign s_csamul_cla32_fa7_3_or0 = s_csamul_cla32_fa7_3_and0 | s_csamul_cla32_fa7_3_and1;
  assign s_csamul_cla32_and8_3 = a[8] & b[3];
  assign s_csamul_cla32_fa8_3_xor0 = s_csamul_cla32_and8_3 ^ s_csamul_cla32_fa9_2_xor1;
  assign s_csamul_cla32_fa8_3_and0 = s_csamul_cla32_and8_3 & s_csamul_cla32_fa9_2_xor1;
  assign s_csamul_cla32_fa8_3_xor1 = s_csamul_cla32_fa8_3_xor0 ^ s_csamul_cla32_fa8_2_or0;
  assign s_csamul_cla32_fa8_3_and1 = s_csamul_cla32_fa8_3_xor0 & s_csamul_cla32_fa8_2_or0;
  assign s_csamul_cla32_fa8_3_or0 = s_csamul_cla32_fa8_3_and0 | s_csamul_cla32_fa8_3_and1;
  assign s_csamul_cla32_and9_3 = a[9] & b[3];
  assign s_csamul_cla32_fa9_3_xor0 = s_csamul_cla32_and9_3 ^ s_csamul_cla32_fa10_2_xor1;
  assign s_csamul_cla32_fa9_3_and0 = s_csamul_cla32_and9_3 & s_csamul_cla32_fa10_2_xor1;
  assign s_csamul_cla32_fa9_3_xor1 = s_csamul_cla32_fa9_3_xor0 ^ s_csamul_cla32_fa9_2_or0;
  assign s_csamul_cla32_fa9_3_and1 = s_csamul_cla32_fa9_3_xor0 & s_csamul_cla32_fa9_2_or0;
  assign s_csamul_cla32_fa9_3_or0 = s_csamul_cla32_fa9_3_and0 | s_csamul_cla32_fa9_3_and1;
  assign s_csamul_cla32_and10_3 = a[10] & b[3];
  assign s_csamul_cla32_fa10_3_xor0 = s_csamul_cla32_and10_3 ^ s_csamul_cla32_fa11_2_xor1;
  assign s_csamul_cla32_fa10_3_and0 = s_csamul_cla32_and10_3 & s_csamul_cla32_fa11_2_xor1;
  assign s_csamul_cla32_fa10_3_xor1 = s_csamul_cla32_fa10_3_xor0 ^ s_csamul_cla32_fa10_2_or0;
  assign s_csamul_cla32_fa10_3_and1 = s_csamul_cla32_fa10_3_xor0 & s_csamul_cla32_fa10_2_or0;
  assign s_csamul_cla32_fa10_3_or0 = s_csamul_cla32_fa10_3_and0 | s_csamul_cla32_fa10_3_and1;
  assign s_csamul_cla32_and11_3 = a[11] & b[3];
  assign s_csamul_cla32_fa11_3_xor0 = s_csamul_cla32_and11_3 ^ s_csamul_cla32_fa12_2_xor1;
  assign s_csamul_cla32_fa11_3_and0 = s_csamul_cla32_and11_3 & s_csamul_cla32_fa12_2_xor1;
  assign s_csamul_cla32_fa11_3_xor1 = s_csamul_cla32_fa11_3_xor0 ^ s_csamul_cla32_fa11_2_or0;
  assign s_csamul_cla32_fa11_3_and1 = s_csamul_cla32_fa11_3_xor0 & s_csamul_cla32_fa11_2_or0;
  assign s_csamul_cla32_fa11_3_or0 = s_csamul_cla32_fa11_3_and0 | s_csamul_cla32_fa11_3_and1;
  assign s_csamul_cla32_and12_3 = a[12] & b[3];
  assign s_csamul_cla32_fa12_3_xor0 = s_csamul_cla32_and12_3 ^ s_csamul_cla32_fa13_2_xor1;
  assign s_csamul_cla32_fa12_3_and0 = s_csamul_cla32_and12_3 & s_csamul_cla32_fa13_2_xor1;
  assign s_csamul_cla32_fa12_3_xor1 = s_csamul_cla32_fa12_3_xor0 ^ s_csamul_cla32_fa12_2_or0;
  assign s_csamul_cla32_fa12_3_and1 = s_csamul_cla32_fa12_3_xor0 & s_csamul_cla32_fa12_2_or0;
  assign s_csamul_cla32_fa12_3_or0 = s_csamul_cla32_fa12_3_and0 | s_csamul_cla32_fa12_3_and1;
  assign s_csamul_cla32_and13_3 = a[13] & b[3];
  assign s_csamul_cla32_fa13_3_xor0 = s_csamul_cla32_and13_3 ^ s_csamul_cla32_fa14_2_xor1;
  assign s_csamul_cla32_fa13_3_and0 = s_csamul_cla32_and13_3 & s_csamul_cla32_fa14_2_xor1;
  assign s_csamul_cla32_fa13_3_xor1 = s_csamul_cla32_fa13_3_xor0 ^ s_csamul_cla32_fa13_2_or0;
  assign s_csamul_cla32_fa13_3_and1 = s_csamul_cla32_fa13_3_xor0 & s_csamul_cla32_fa13_2_or0;
  assign s_csamul_cla32_fa13_3_or0 = s_csamul_cla32_fa13_3_and0 | s_csamul_cla32_fa13_3_and1;
  assign s_csamul_cla32_and14_3 = a[14] & b[3];
  assign s_csamul_cla32_fa14_3_xor0 = s_csamul_cla32_and14_3 ^ s_csamul_cla32_fa15_2_xor1;
  assign s_csamul_cla32_fa14_3_and0 = s_csamul_cla32_and14_3 & s_csamul_cla32_fa15_2_xor1;
  assign s_csamul_cla32_fa14_3_xor1 = s_csamul_cla32_fa14_3_xor0 ^ s_csamul_cla32_fa14_2_or0;
  assign s_csamul_cla32_fa14_3_and1 = s_csamul_cla32_fa14_3_xor0 & s_csamul_cla32_fa14_2_or0;
  assign s_csamul_cla32_fa14_3_or0 = s_csamul_cla32_fa14_3_and0 | s_csamul_cla32_fa14_3_and1;
  assign s_csamul_cla32_and15_3 = a[15] & b[3];
  assign s_csamul_cla32_fa15_3_xor0 = s_csamul_cla32_and15_3 ^ s_csamul_cla32_fa16_2_xor1;
  assign s_csamul_cla32_fa15_3_and0 = s_csamul_cla32_and15_3 & s_csamul_cla32_fa16_2_xor1;
  assign s_csamul_cla32_fa15_3_xor1 = s_csamul_cla32_fa15_3_xor0 ^ s_csamul_cla32_fa15_2_or0;
  assign s_csamul_cla32_fa15_3_and1 = s_csamul_cla32_fa15_3_xor0 & s_csamul_cla32_fa15_2_or0;
  assign s_csamul_cla32_fa15_3_or0 = s_csamul_cla32_fa15_3_and0 | s_csamul_cla32_fa15_3_and1;
  assign s_csamul_cla32_and16_3 = a[16] & b[3];
  assign s_csamul_cla32_fa16_3_xor0 = s_csamul_cla32_and16_3 ^ s_csamul_cla32_fa17_2_xor1;
  assign s_csamul_cla32_fa16_3_and0 = s_csamul_cla32_and16_3 & s_csamul_cla32_fa17_2_xor1;
  assign s_csamul_cla32_fa16_3_xor1 = s_csamul_cla32_fa16_3_xor0 ^ s_csamul_cla32_fa16_2_or0;
  assign s_csamul_cla32_fa16_3_and1 = s_csamul_cla32_fa16_3_xor0 & s_csamul_cla32_fa16_2_or0;
  assign s_csamul_cla32_fa16_3_or0 = s_csamul_cla32_fa16_3_and0 | s_csamul_cla32_fa16_3_and1;
  assign s_csamul_cla32_and17_3 = a[17] & b[3];
  assign s_csamul_cla32_fa17_3_xor0 = s_csamul_cla32_and17_3 ^ s_csamul_cla32_fa18_2_xor1;
  assign s_csamul_cla32_fa17_3_and0 = s_csamul_cla32_and17_3 & s_csamul_cla32_fa18_2_xor1;
  assign s_csamul_cla32_fa17_3_xor1 = s_csamul_cla32_fa17_3_xor0 ^ s_csamul_cla32_fa17_2_or0;
  assign s_csamul_cla32_fa17_3_and1 = s_csamul_cla32_fa17_3_xor0 & s_csamul_cla32_fa17_2_or0;
  assign s_csamul_cla32_fa17_3_or0 = s_csamul_cla32_fa17_3_and0 | s_csamul_cla32_fa17_3_and1;
  assign s_csamul_cla32_and18_3 = a[18] & b[3];
  assign s_csamul_cla32_fa18_3_xor0 = s_csamul_cla32_and18_3 ^ s_csamul_cla32_fa19_2_xor1;
  assign s_csamul_cla32_fa18_3_and0 = s_csamul_cla32_and18_3 & s_csamul_cla32_fa19_2_xor1;
  assign s_csamul_cla32_fa18_3_xor1 = s_csamul_cla32_fa18_3_xor0 ^ s_csamul_cla32_fa18_2_or0;
  assign s_csamul_cla32_fa18_3_and1 = s_csamul_cla32_fa18_3_xor0 & s_csamul_cla32_fa18_2_or0;
  assign s_csamul_cla32_fa18_3_or0 = s_csamul_cla32_fa18_3_and0 | s_csamul_cla32_fa18_3_and1;
  assign s_csamul_cla32_and19_3 = a[19] & b[3];
  assign s_csamul_cla32_fa19_3_xor0 = s_csamul_cla32_and19_3 ^ s_csamul_cla32_fa20_2_xor1;
  assign s_csamul_cla32_fa19_3_and0 = s_csamul_cla32_and19_3 & s_csamul_cla32_fa20_2_xor1;
  assign s_csamul_cla32_fa19_3_xor1 = s_csamul_cla32_fa19_3_xor0 ^ s_csamul_cla32_fa19_2_or0;
  assign s_csamul_cla32_fa19_3_and1 = s_csamul_cla32_fa19_3_xor0 & s_csamul_cla32_fa19_2_or0;
  assign s_csamul_cla32_fa19_3_or0 = s_csamul_cla32_fa19_3_and0 | s_csamul_cla32_fa19_3_and1;
  assign s_csamul_cla32_and20_3 = a[20] & b[3];
  assign s_csamul_cla32_fa20_3_xor0 = s_csamul_cla32_and20_3 ^ s_csamul_cla32_fa21_2_xor1;
  assign s_csamul_cla32_fa20_3_and0 = s_csamul_cla32_and20_3 & s_csamul_cla32_fa21_2_xor1;
  assign s_csamul_cla32_fa20_3_xor1 = s_csamul_cla32_fa20_3_xor0 ^ s_csamul_cla32_fa20_2_or0;
  assign s_csamul_cla32_fa20_3_and1 = s_csamul_cla32_fa20_3_xor0 & s_csamul_cla32_fa20_2_or0;
  assign s_csamul_cla32_fa20_3_or0 = s_csamul_cla32_fa20_3_and0 | s_csamul_cla32_fa20_3_and1;
  assign s_csamul_cla32_and21_3 = a[21] & b[3];
  assign s_csamul_cla32_fa21_3_xor0 = s_csamul_cla32_and21_3 ^ s_csamul_cla32_fa22_2_xor1;
  assign s_csamul_cla32_fa21_3_and0 = s_csamul_cla32_and21_3 & s_csamul_cla32_fa22_2_xor1;
  assign s_csamul_cla32_fa21_3_xor1 = s_csamul_cla32_fa21_3_xor0 ^ s_csamul_cla32_fa21_2_or0;
  assign s_csamul_cla32_fa21_3_and1 = s_csamul_cla32_fa21_3_xor0 & s_csamul_cla32_fa21_2_or0;
  assign s_csamul_cla32_fa21_3_or0 = s_csamul_cla32_fa21_3_and0 | s_csamul_cla32_fa21_3_and1;
  assign s_csamul_cla32_and22_3 = a[22] & b[3];
  assign s_csamul_cla32_fa22_3_xor0 = s_csamul_cla32_and22_3 ^ s_csamul_cla32_fa23_2_xor1;
  assign s_csamul_cla32_fa22_3_and0 = s_csamul_cla32_and22_3 & s_csamul_cla32_fa23_2_xor1;
  assign s_csamul_cla32_fa22_3_xor1 = s_csamul_cla32_fa22_3_xor0 ^ s_csamul_cla32_fa22_2_or0;
  assign s_csamul_cla32_fa22_3_and1 = s_csamul_cla32_fa22_3_xor0 & s_csamul_cla32_fa22_2_or0;
  assign s_csamul_cla32_fa22_3_or0 = s_csamul_cla32_fa22_3_and0 | s_csamul_cla32_fa22_3_and1;
  assign s_csamul_cla32_and23_3 = a[23] & b[3];
  assign s_csamul_cla32_fa23_3_xor0 = s_csamul_cla32_and23_3 ^ s_csamul_cla32_fa24_2_xor1;
  assign s_csamul_cla32_fa23_3_and0 = s_csamul_cla32_and23_3 & s_csamul_cla32_fa24_2_xor1;
  assign s_csamul_cla32_fa23_3_xor1 = s_csamul_cla32_fa23_3_xor0 ^ s_csamul_cla32_fa23_2_or0;
  assign s_csamul_cla32_fa23_3_and1 = s_csamul_cla32_fa23_3_xor0 & s_csamul_cla32_fa23_2_or0;
  assign s_csamul_cla32_fa23_3_or0 = s_csamul_cla32_fa23_3_and0 | s_csamul_cla32_fa23_3_and1;
  assign s_csamul_cla32_and24_3 = a[24] & b[3];
  assign s_csamul_cla32_fa24_3_xor0 = s_csamul_cla32_and24_3 ^ s_csamul_cla32_fa25_2_xor1;
  assign s_csamul_cla32_fa24_3_and0 = s_csamul_cla32_and24_3 & s_csamul_cla32_fa25_2_xor1;
  assign s_csamul_cla32_fa24_3_xor1 = s_csamul_cla32_fa24_3_xor0 ^ s_csamul_cla32_fa24_2_or0;
  assign s_csamul_cla32_fa24_3_and1 = s_csamul_cla32_fa24_3_xor0 & s_csamul_cla32_fa24_2_or0;
  assign s_csamul_cla32_fa24_3_or0 = s_csamul_cla32_fa24_3_and0 | s_csamul_cla32_fa24_3_and1;
  assign s_csamul_cla32_and25_3 = a[25] & b[3];
  assign s_csamul_cla32_fa25_3_xor0 = s_csamul_cla32_and25_3 ^ s_csamul_cla32_fa26_2_xor1;
  assign s_csamul_cla32_fa25_3_and0 = s_csamul_cla32_and25_3 & s_csamul_cla32_fa26_2_xor1;
  assign s_csamul_cla32_fa25_3_xor1 = s_csamul_cla32_fa25_3_xor0 ^ s_csamul_cla32_fa25_2_or0;
  assign s_csamul_cla32_fa25_3_and1 = s_csamul_cla32_fa25_3_xor0 & s_csamul_cla32_fa25_2_or0;
  assign s_csamul_cla32_fa25_3_or0 = s_csamul_cla32_fa25_3_and0 | s_csamul_cla32_fa25_3_and1;
  assign s_csamul_cla32_and26_3 = a[26] & b[3];
  assign s_csamul_cla32_fa26_3_xor0 = s_csamul_cla32_and26_3 ^ s_csamul_cla32_fa27_2_xor1;
  assign s_csamul_cla32_fa26_3_and0 = s_csamul_cla32_and26_3 & s_csamul_cla32_fa27_2_xor1;
  assign s_csamul_cla32_fa26_3_xor1 = s_csamul_cla32_fa26_3_xor0 ^ s_csamul_cla32_fa26_2_or0;
  assign s_csamul_cla32_fa26_3_and1 = s_csamul_cla32_fa26_3_xor0 & s_csamul_cla32_fa26_2_or0;
  assign s_csamul_cla32_fa26_3_or0 = s_csamul_cla32_fa26_3_and0 | s_csamul_cla32_fa26_3_and1;
  assign s_csamul_cla32_and27_3 = a[27] & b[3];
  assign s_csamul_cla32_fa27_3_xor0 = s_csamul_cla32_and27_3 ^ s_csamul_cla32_fa28_2_xor1;
  assign s_csamul_cla32_fa27_3_and0 = s_csamul_cla32_and27_3 & s_csamul_cla32_fa28_2_xor1;
  assign s_csamul_cla32_fa27_3_xor1 = s_csamul_cla32_fa27_3_xor0 ^ s_csamul_cla32_fa27_2_or0;
  assign s_csamul_cla32_fa27_3_and1 = s_csamul_cla32_fa27_3_xor0 & s_csamul_cla32_fa27_2_or0;
  assign s_csamul_cla32_fa27_3_or0 = s_csamul_cla32_fa27_3_and0 | s_csamul_cla32_fa27_3_and1;
  assign s_csamul_cla32_and28_3 = a[28] & b[3];
  assign s_csamul_cla32_fa28_3_xor0 = s_csamul_cla32_and28_3 ^ s_csamul_cla32_fa29_2_xor1;
  assign s_csamul_cla32_fa28_3_and0 = s_csamul_cla32_and28_3 & s_csamul_cla32_fa29_2_xor1;
  assign s_csamul_cla32_fa28_3_xor1 = s_csamul_cla32_fa28_3_xor0 ^ s_csamul_cla32_fa28_2_or0;
  assign s_csamul_cla32_fa28_3_and1 = s_csamul_cla32_fa28_3_xor0 & s_csamul_cla32_fa28_2_or0;
  assign s_csamul_cla32_fa28_3_or0 = s_csamul_cla32_fa28_3_and0 | s_csamul_cla32_fa28_3_and1;
  assign s_csamul_cla32_and29_3 = a[29] & b[3];
  assign s_csamul_cla32_fa29_3_xor0 = s_csamul_cla32_and29_3 ^ s_csamul_cla32_fa30_2_xor1;
  assign s_csamul_cla32_fa29_3_and0 = s_csamul_cla32_and29_3 & s_csamul_cla32_fa30_2_xor1;
  assign s_csamul_cla32_fa29_3_xor1 = s_csamul_cla32_fa29_3_xor0 ^ s_csamul_cla32_fa29_2_or0;
  assign s_csamul_cla32_fa29_3_and1 = s_csamul_cla32_fa29_3_xor0 & s_csamul_cla32_fa29_2_or0;
  assign s_csamul_cla32_fa29_3_or0 = s_csamul_cla32_fa29_3_and0 | s_csamul_cla32_fa29_3_and1;
  assign s_csamul_cla32_and30_3 = a[30] & b[3];
  assign s_csamul_cla32_fa30_3_xor0 = s_csamul_cla32_and30_3 ^ s_csamul_cla32_ha31_2_xor0;
  assign s_csamul_cla32_fa30_3_and0 = s_csamul_cla32_and30_3 & s_csamul_cla32_ha31_2_xor0;
  assign s_csamul_cla32_fa30_3_xor1 = s_csamul_cla32_fa30_3_xor0 ^ s_csamul_cla32_fa30_2_or0;
  assign s_csamul_cla32_fa30_3_and1 = s_csamul_cla32_fa30_3_xor0 & s_csamul_cla32_fa30_2_or0;
  assign s_csamul_cla32_fa30_3_or0 = s_csamul_cla32_fa30_3_and0 | s_csamul_cla32_fa30_3_and1;
  assign s_csamul_cla32_nand31_3 = ~(a[31] & b[3]);
  assign s_csamul_cla32_ha31_3_xor0 = s_csamul_cla32_nand31_3 ^ s_csamul_cla32_ha31_2_and0;
  assign s_csamul_cla32_ha31_3_and0 = s_csamul_cla32_nand31_3 & s_csamul_cla32_ha31_2_and0;
  assign s_csamul_cla32_and0_4 = a[0] & b[4];
  assign s_csamul_cla32_fa0_4_xor0 = s_csamul_cla32_and0_4 ^ s_csamul_cla32_fa1_3_xor1;
  assign s_csamul_cla32_fa0_4_and0 = s_csamul_cla32_and0_4 & s_csamul_cla32_fa1_3_xor1;
  assign s_csamul_cla32_fa0_4_xor1 = s_csamul_cla32_fa0_4_xor0 ^ s_csamul_cla32_fa0_3_or0;
  assign s_csamul_cla32_fa0_4_and1 = s_csamul_cla32_fa0_4_xor0 & s_csamul_cla32_fa0_3_or0;
  assign s_csamul_cla32_fa0_4_or0 = s_csamul_cla32_fa0_4_and0 | s_csamul_cla32_fa0_4_and1;
  assign s_csamul_cla32_and1_4 = a[1] & b[4];
  assign s_csamul_cla32_fa1_4_xor0 = s_csamul_cla32_and1_4 ^ s_csamul_cla32_fa2_3_xor1;
  assign s_csamul_cla32_fa1_4_and0 = s_csamul_cla32_and1_4 & s_csamul_cla32_fa2_3_xor1;
  assign s_csamul_cla32_fa1_4_xor1 = s_csamul_cla32_fa1_4_xor0 ^ s_csamul_cla32_fa1_3_or0;
  assign s_csamul_cla32_fa1_4_and1 = s_csamul_cla32_fa1_4_xor0 & s_csamul_cla32_fa1_3_or0;
  assign s_csamul_cla32_fa1_4_or0 = s_csamul_cla32_fa1_4_and0 | s_csamul_cla32_fa1_4_and1;
  assign s_csamul_cla32_and2_4 = a[2] & b[4];
  assign s_csamul_cla32_fa2_4_xor0 = s_csamul_cla32_and2_4 ^ s_csamul_cla32_fa3_3_xor1;
  assign s_csamul_cla32_fa2_4_and0 = s_csamul_cla32_and2_4 & s_csamul_cla32_fa3_3_xor1;
  assign s_csamul_cla32_fa2_4_xor1 = s_csamul_cla32_fa2_4_xor0 ^ s_csamul_cla32_fa2_3_or0;
  assign s_csamul_cla32_fa2_4_and1 = s_csamul_cla32_fa2_4_xor0 & s_csamul_cla32_fa2_3_or0;
  assign s_csamul_cla32_fa2_4_or0 = s_csamul_cla32_fa2_4_and0 | s_csamul_cla32_fa2_4_and1;
  assign s_csamul_cla32_and3_4 = a[3] & b[4];
  assign s_csamul_cla32_fa3_4_xor0 = s_csamul_cla32_and3_4 ^ s_csamul_cla32_fa4_3_xor1;
  assign s_csamul_cla32_fa3_4_and0 = s_csamul_cla32_and3_4 & s_csamul_cla32_fa4_3_xor1;
  assign s_csamul_cla32_fa3_4_xor1 = s_csamul_cla32_fa3_4_xor0 ^ s_csamul_cla32_fa3_3_or0;
  assign s_csamul_cla32_fa3_4_and1 = s_csamul_cla32_fa3_4_xor0 & s_csamul_cla32_fa3_3_or0;
  assign s_csamul_cla32_fa3_4_or0 = s_csamul_cla32_fa3_4_and0 | s_csamul_cla32_fa3_4_and1;
  assign s_csamul_cla32_and4_4 = a[4] & b[4];
  assign s_csamul_cla32_fa4_4_xor0 = s_csamul_cla32_and4_4 ^ s_csamul_cla32_fa5_3_xor1;
  assign s_csamul_cla32_fa4_4_and0 = s_csamul_cla32_and4_4 & s_csamul_cla32_fa5_3_xor1;
  assign s_csamul_cla32_fa4_4_xor1 = s_csamul_cla32_fa4_4_xor0 ^ s_csamul_cla32_fa4_3_or0;
  assign s_csamul_cla32_fa4_4_and1 = s_csamul_cla32_fa4_4_xor0 & s_csamul_cla32_fa4_3_or0;
  assign s_csamul_cla32_fa4_4_or0 = s_csamul_cla32_fa4_4_and0 | s_csamul_cla32_fa4_4_and1;
  assign s_csamul_cla32_and5_4 = a[5] & b[4];
  assign s_csamul_cla32_fa5_4_xor0 = s_csamul_cla32_and5_4 ^ s_csamul_cla32_fa6_3_xor1;
  assign s_csamul_cla32_fa5_4_and0 = s_csamul_cla32_and5_4 & s_csamul_cla32_fa6_3_xor1;
  assign s_csamul_cla32_fa5_4_xor1 = s_csamul_cla32_fa5_4_xor0 ^ s_csamul_cla32_fa5_3_or0;
  assign s_csamul_cla32_fa5_4_and1 = s_csamul_cla32_fa5_4_xor0 & s_csamul_cla32_fa5_3_or0;
  assign s_csamul_cla32_fa5_4_or0 = s_csamul_cla32_fa5_4_and0 | s_csamul_cla32_fa5_4_and1;
  assign s_csamul_cla32_and6_4 = a[6] & b[4];
  assign s_csamul_cla32_fa6_4_xor0 = s_csamul_cla32_and6_4 ^ s_csamul_cla32_fa7_3_xor1;
  assign s_csamul_cla32_fa6_4_and0 = s_csamul_cla32_and6_4 & s_csamul_cla32_fa7_3_xor1;
  assign s_csamul_cla32_fa6_4_xor1 = s_csamul_cla32_fa6_4_xor0 ^ s_csamul_cla32_fa6_3_or0;
  assign s_csamul_cla32_fa6_4_and1 = s_csamul_cla32_fa6_4_xor0 & s_csamul_cla32_fa6_3_or0;
  assign s_csamul_cla32_fa6_4_or0 = s_csamul_cla32_fa6_4_and0 | s_csamul_cla32_fa6_4_and1;
  assign s_csamul_cla32_and7_4 = a[7] & b[4];
  assign s_csamul_cla32_fa7_4_xor0 = s_csamul_cla32_and7_4 ^ s_csamul_cla32_fa8_3_xor1;
  assign s_csamul_cla32_fa7_4_and0 = s_csamul_cla32_and7_4 & s_csamul_cla32_fa8_3_xor1;
  assign s_csamul_cla32_fa7_4_xor1 = s_csamul_cla32_fa7_4_xor0 ^ s_csamul_cla32_fa7_3_or0;
  assign s_csamul_cla32_fa7_4_and1 = s_csamul_cla32_fa7_4_xor0 & s_csamul_cla32_fa7_3_or0;
  assign s_csamul_cla32_fa7_4_or0 = s_csamul_cla32_fa7_4_and0 | s_csamul_cla32_fa7_4_and1;
  assign s_csamul_cla32_and8_4 = a[8] & b[4];
  assign s_csamul_cla32_fa8_4_xor0 = s_csamul_cla32_and8_4 ^ s_csamul_cla32_fa9_3_xor1;
  assign s_csamul_cla32_fa8_4_and0 = s_csamul_cla32_and8_4 & s_csamul_cla32_fa9_3_xor1;
  assign s_csamul_cla32_fa8_4_xor1 = s_csamul_cla32_fa8_4_xor0 ^ s_csamul_cla32_fa8_3_or0;
  assign s_csamul_cla32_fa8_4_and1 = s_csamul_cla32_fa8_4_xor0 & s_csamul_cla32_fa8_3_or0;
  assign s_csamul_cla32_fa8_4_or0 = s_csamul_cla32_fa8_4_and0 | s_csamul_cla32_fa8_4_and1;
  assign s_csamul_cla32_and9_4 = a[9] & b[4];
  assign s_csamul_cla32_fa9_4_xor0 = s_csamul_cla32_and9_4 ^ s_csamul_cla32_fa10_3_xor1;
  assign s_csamul_cla32_fa9_4_and0 = s_csamul_cla32_and9_4 & s_csamul_cla32_fa10_3_xor1;
  assign s_csamul_cla32_fa9_4_xor1 = s_csamul_cla32_fa9_4_xor0 ^ s_csamul_cla32_fa9_3_or0;
  assign s_csamul_cla32_fa9_4_and1 = s_csamul_cla32_fa9_4_xor0 & s_csamul_cla32_fa9_3_or0;
  assign s_csamul_cla32_fa9_4_or0 = s_csamul_cla32_fa9_4_and0 | s_csamul_cla32_fa9_4_and1;
  assign s_csamul_cla32_and10_4 = a[10] & b[4];
  assign s_csamul_cla32_fa10_4_xor0 = s_csamul_cla32_and10_4 ^ s_csamul_cla32_fa11_3_xor1;
  assign s_csamul_cla32_fa10_4_and0 = s_csamul_cla32_and10_4 & s_csamul_cla32_fa11_3_xor1;
  assign s_csamul_cla32_fa10_4_xor1 = s_csamul_cla32_fa10_4_xor0 ^ s_csamul_cla32_fa10_3_or0;
  assign s_csamul_cla32_fa10_4_and1 = s_csamul_cla32_fa10_4_xor0 & s_csamul_cla32_fa10_3_or0;
  assign s_csamul_cla32_fa10_4_or0 = s_csamul_cla32_fa10_4_and0 | s_csamul_cla32_fa10_4_and1;
  assign s_csamul_cla32_and11_4 = a[11] & b[4];
  assign s_csamul_cla32_fa11_4_xor0 = s_csamul_cla32_and11_4 ^ s_csamul_cla32_fa12_3_xor1;
  assign s_csamul_cla32_fa11_4_and0 = s_csamul_cla32_and11_4 & s_csamul_cla32_fa12_3_xor1;
  assign s_csamul_cla32_fa11_4_xor1 = s_csamul_cla32_fa11_4_xor0 ^ s_csamul_cla32_fa11_3_or0;
  assign s_csamul_cla32_fa11_4_and1 = s_csamul_cla32_fa11_4_xor0 & s_csamul_cla32_fa11_3_or0;
  assign s_csamul_cla32_fa11_4_or0 = s_csamul_cla32_fa11_4_and0 | s_csamul_cla32_fa11_4_and1;
  assign s_csamul_cla32_and12_4 = a[12] & b[4];
  assign s_csamul_cla32_fa12_4_xor0 = s_csamul_cla32_and12_4 ^ s_csamul_cla32_fa13_3_xor1;
  assign s_csamul_cla32_fa12_4_and0 = s_csamul_cla32_and12_4 & s_csamul_cla32_fa13_3_xor1;
  assign s_csamul_cla32_fa12_4_xor1 = s_csamul_cla32_fa12_4_xor0 ^ s_csamul_cla32_fa12_3_or0;
  assign s_csamul_cla32_fa12_4_and1 = s_csamul_cla32_fa12_4_xor0 & s_csamul_cla32_fa12_3_or0;
  assign s_csamul_cla32_fa12_4_or0 = s_csamul_cla32_fa12_4_and0 | s_csamul_cla32_fa12_4_and1;
  assign s_csamul_cla32_and13_4 = a[13] & b[4];
  assign s_csamul_cla32_fa13_4_xor0 = s_csamul_cla32_and13_4 ^ s_csamul_cla32_fa14_3_xor1;
  assign s_csamul_cla32_fa13_4_and0 = s_csamul_cla32_and13_4 & s_csamul_cla32_fa14_3_xor1;
  assign s_csamul_cla32_fa13_4_xor1 = s_csamul_cla32_fa13_4_xor0 ^ s_csamul_cla32_fa13_3_or0;
  assign s_csamul_cla32_fa13_4_and1 = s_csamul_cla32_fa13_4_xor0 & s_csamul_cla32_fa13_3_or0;
  assign s_csamul_cla32_fa13_4_or0 = s_csamul_cla32_fa13_4_and0 | s_csamul_cla32_fa13_4_and1;
  assign s_csamul_cla32_and14_4 = a[14] & b[4];
  assign s_csamul_cla32_fa14_4_xor0 = s_csamul_cla32_and14_4 ^ s_csamul_cla32_fa15_3_xor1;
  assign s_csamul_cla32_fa14_4_and0 = s_csamul_cla32_and14_4 & s_csamul_cla32_fa15_3_xor1;
  assign s_csamul_cla32_fa14_4_xor1 = s_csamul_cla32_fa14_4_xor0 ^ s_csamul_cla32_fa14_3_or0;
  assign s_csamul_cla32_fa14_4_and1 = s_csamul_cla32_fa14_4_xor0 & s_csamul_cla32_fa14_3_or0;
  assign s_csamul_cla32_fa14_4_or0 = s_csamul_cla32_fa14_4_and0 | s_csamul_cla32_fa14_4_and1;
  assign s_csamul_cla32_and15_4 = a[15] & b[4];
  assign s_csamul_cla32_fa15_4_xor0 = s_csamul_cla32_and15_4 ^ s_csamul_cla32_fa16_3_xor1;
  assign s_csamul_cla32_fa15_4_and0 = s_csamul_cla32_and15_4 & s_csamul_cla32_fa16_3_xor1;
  assign s_csamul_cla32_fa15_4_xor1 = s_csamul_cla32_fa15_4_xor0 ^ s_csamul_cla32_fa15_3_or0;
  assign s_csamul_cla32_fa15_4_and1 = s_csamul_cla32_fa15_4_xor0 & s_csamul_cla32_fa15_3_or0;
  assign s_csamul_cla32_fa15_4_or0 = s_csamul_cla32_fa15_4_and0 | s_csamul_cla32_fa15_4_and1;
  assign s_csamul_cla32_and16_4 = a[16] & b[4];
  assign s_csamul_cla32_fa16_4_xor0 = s_csamul_cla32_and16_4 ^ s_csamul_cla32_fa17_3_xor1;
  assign s_csamul_cla32_fa16_4_and0 = s_csamul_cla32_and16_4 & s_csamul_cla32_fa17_3_xor1;
  assign s_csamul_cla32_fa16_4_xor1 = s_csamul_cla32_fa16_4_xor0 ^ s_csamul_cla32_fa16_3_or0;
  assign s_csamul_cla32_fa16_4_and1 = s_csamul_cla32_fa16_4_xor0 & s_csamul_cla32_fa16_3_or0;
  assign s_csamul_cla32_fa16_4_or0 = s_csamul_cla32_fa16_4_and0 | s_csamul_cla32_fa16_4_and1;
  assign s_csamul_cla32_and17_4 = a[17] & b[4];
  assign s_csamul_cla32_fa17_4_xor0 = s_csamul_cla32_and17_4 ^ s_csamul_cla32_fa18_3_xor1;
  assign s_csamul_cla32_fa17_4_and0 = s_csamul_cla32_and17_4 & s_csamul_cla32_fa18_3_xor1;
  assign s_csamul_cla32_fa17_4_xor1 = s_csamul_cla32_fa17_4_xor0 ^ s_csamul_cla32_fa17_3_or0;
  assign s_csamul_cla32_fa17_4_and1 = s_csamul_cla32_fa17_4_xor0 & s_csamul_cla32_fa17_3_or0;
  assign s_csamul_cla32_fa17_4_or0 = s_csamul_cla32_fa17_4_and0 | s_csamul_cla32_fa17_4_and1;
  assign s_csamul_cla32_and18_4 = a[18] & b[4];
  assign s_csamul_cla32_fa18_4_xor0 = s_csamul_cla32_and18_4 ^ s_csamul_cla32_fa19_3_xor1;
  assign s_csamul_cla32_fa18_4_and0 = s_csamul_cla32_and18_4 & s_csamul_cla32_fa19_3_xor1;
  assign s_csamul_cla32_fa18_4_xor1 = s_csamul_cla32_fa18_4_xor0 ^ s_csamul_cla32_fa18_3_or0;
  assign s_csamul_cla32_fa18_4_and1 = s_csamul_cla32_fa18_4_xor0 & s_csamul_cla32_fa18_3_or0;
  assign s_csamul_cla32_fa18_4_or0 = s_csamul_cla32_fa18_4_and0 | s_csamul_cla32_fa18_4_and1;
  assign s_csamul_cla32_and19_4 = a[19] & b[4];
  assign s_csamul_cla32_fa19_4_xor0 = s_csamul_cla32_and19_4 ^ s_csamul_cla32_fa20_3_xor1;
  assign s_csamul_cla32_fa19_4_and0 = s_csamul_cla32_and19_4 & s_csamul_cla32_fa20_3_xor1;
  assign s_csamul_cla32_fa19_4_xor1 = s_csamul_cla32_fa19_4_xor0 ^ s_csamul_cla32_fa19_3_or0;
  assign s_csamul_cla32_fa19_4_and1 = s_csamul_cla32_fa19_4_xor0 & s_csamul_cla32_fa19_3_or0;
  assign s_csamul_cla32_fa19_4_or0 = s_csamul_cla32_fa19_4_and0 | s_csamul_cla32_fa19_4_and1;
  assign s_csamul_cla32_and20_4 = a[20] & b[4];
  assign s_csamul_cla32_fa20_4_xor0 = s_csamul_cla32_and20_4 ^ s_csamul_cla32_fa21_3_xor1;
  assign s_csamul_cla32_fa20_4_and0 = s_csamul_cla32_and20_4 & s_csamul_cla32_fa21_3_xor1;
  assign s_csamul_cla32_fa20_4_xor1 = s_csamul_cla32_fa20_4_xor0 ^ s_csamul_cla32_fa20_3_or0;
  assign s_csamul_cla32_fa20_4_and1 = s_csamul_cla32_fa20_4_xor0 & s_csamul_cla32_fa20_3_or0;
  assign s_csamul_cla32_fa20_4_or0 = s_csamul_cla32_fa20_4_and0 | s_csamul_cla32_fa20_4_and1;
  assign s_csamul_cla32_and21_4 = a[21] & b[4];
  assign s_csamul_cla32_fa21_4_xor0 = s_csamul_cla32_and21_4 ^ s_csamul_cla32_fa22_3_xor1;
  assign s_csamul_cla32_fa21_4_and0 = s_csamul_cla32_and21_4 & s_csamul_cla32_fa22_3_xor1;
  assign s_csamul_cla32_fa21_4_xor1 = s_csamul_cla32_fa21_4_xor0 ^ s_csamul_cla32_fa21_3_or0;
  assign s_csamul_cla32_fa21_4_and1 = s_csamul_cla32_fa21_4_xor0 & s_csamul_cla32_fa21_3_or0;
  assign s_csamul_cla32_fa21_4_or0 = s_csamul_cla32_fa21_4_and0 | s_csamul_cla32_fa21_4_and1;
  assign s_csamul_cla32_and22_4 = a[22] & b[4];
  assign s_csamul_cla32_fa22_4_xor0 = s_csamul_cla32_and22_4 ^ s_csamul_cla32_fa23_3_xor1;
  assign s_csamul_cla32_fa22_4_and0 = s_csamul_cla32_and22_4 & s_csamul_cla32_fa23_3_xor1;
  assign s_csamul_cla32_fa22_4_xor1 = s_csamul_cla32_fa22_4_xor0 ^ s_csamul_cla32_fa22_3_or0;
  assign s_csamul_cla32_fa22_4_and1 = s_csamul_cla32_fa22_4_xor0 & s_csamul_cla32_fa22_3_or0;
  assign s_csamul_cla32_fa22_4_or0 = s_csamul_cla32_fa22_4_and0 | s_csamul_cla32_fa22_4_and1;
  assign s_csamul_cla32_and23_4 = a[23] & b[4];
  assign s_csamul_cla32_fa23_4_xor0 = s_csamul_cla32_and23_4 ^ s_csamul_cla32_fa24_3_xor1;
  assign s_csamul_cla32_fa23_4_and0 = s_csamul_cla32_and23_4 & s_csamul_cla32_fa24_3_xor1;
  assign s_csamul_cla32_fa23_4_xor1 = s_csamul_cla32_fa23_4_xor0 ^ s_csamul_cla32_fa23_3_or0;
  assign s_csamul_cla32_fa23_4_and1 = s_csamul_cla32_fa23_4_xor0 & s_csamul_cla32_fa23_3_or0;
  assign s_csamul_cla32_fa23_4_or0 = s_csamul_cla32_fa23_4_and0 | s_csamul_cla32_fa23_4_and1;
  assign s_csamul_cla32_and24_4 = a[24] & b[4];
  assign s_csamul_cla32_fa24_4_xor0 = s_csamul_cla32_and24_4 ^ s_csamul_cla32_fa25_3_xor1;
  assign s_csamul_cla32_fa24_4_and0 = s_csamul_cla32_and24_4 & s_csamul_cla32_fa25_3_xor1;
  assign s_csamul_cla32_fa24_4_xor1 = s_csamul_cla32_fa24_4_xor0 ^ s_csamul_cla32_fa24_3_or0;
  assign s_csamul_cla32_fa24_4_and1 = s_csamul_cla32_fa24_4_xor0 & s_csamul_cla32_fa24_3_or0;
  assign s_csamul_cla32_fa24_4_or0 = s_csamul_cla32_fa24_4_and0 | s_csamul_cla32_fa24_4_and1;
  assign s_csamul_cla32_and25_4 = a[25] & b[4];
  assign s_csamul_cla32_fa25_4_xor0 = s_csamul_cla32_and25_4 ^ s_csamul_cla32_fa26_3_xor1;
  assign s_csamul_cla32_fa25_4_and0 = s_csamul_cla32_and25_4 & s_csamul_cla32_fa26_3_xor1;
  assign s_csamul_cla32_fa25_4_xor1 = s_csamul_cla32_fa25_4_xor0 ^ s_csamul_cla32_fa25_3_or0;
  assign s_csamul_cla32_fa25_4_and1 = s_csamul_cla32_fa25_4_xor0 & s_csamul_cla32_fa25_3_or0;
  assign s_csamul_cla32_fa25_4_or0 = s_csamul_cla32_fa25_4_and0 | s_csamul_cla32_fa25_4_and1;
  assign s_csamul_cla32_and26_4 = a[26] & b[4];
  assign s_csamul_cla32_fa26_4_xor0 = s_csamul_cla32_and26_4 ^ s_csamul_cla32_fa27_3_xor1;
  assign s_csamul_cla32_fa26_4_and0 = s_csamul_cla32_and26_4 & s_csamul_cla32_fa27_3_xor1;
  assign s_csamul_cla32_fa26_4_xor1 = s_csamul_cla32_fa26_4_xor0 ^ s_csamul_cla32_fa26_3_or0;
  assign s_csamul_cla32_fa26_4_and1 = s_csamul_cla32_fa26_4_xor0 & s_csamul_cla32_fa26_3_or0;
  assign s_csamul_cla32_fa26_4_or0 = s_csamul_cla32_fa26_4_and0 | s_csamul_cla32_fa26_4_and1;
  assign s_csamul_cla32_and27_4 = a[27] & b[4];
  assign s_csamul_cla32_fa27_4_xor0 = s_csamul_cla32_and27_4 ^ s_csamul_cla32_fa28_3_xor1;
  assign s_csamul_cla32_fa27_4_and0 = s_csamul_cla32_and27_4 & s_csamul_cla32_fa28_3_xor1;
  assign s_csamul_cla32_fa27_4_xor1 = s_csamul_cla32_fa27_4_xor0 ^ s_csamul_cla32_fa27_3_or0;
  assign s_csamul_cla32_fa27_4_and1 = s_csamul_cla32_fa27_4_xor0 & s_csamul_cla32_fa27_3_or0;
  assign s_csamul_cla32_fa27_4_or0 = s_csamul_cla32_fa27_4_and0 | s_csamul_cla32_fa27_4_and1;
  assign s_csamul_cla32_and28_4 = a[28] & b[4];
  assign s_csamul_cla32_fa28_4_xor0 = s_csamul_cla32_and28_4 ^ s_csamul_cla32_fa29_3_xor1;
  assign s_csamul_cla32_fa28_4_and0 = s_csamul_cla32_and28_4 & s_csamul_cla32_fa29_3_xor1;
  assign s_csamul_cla32_fa28_4_xor1 = s_csamul_cla32_fa28_4_xor0 ^ s_csamul_cla32_fa28_3_or0;
  assign s_csamul_cla32_fa28_4_and1 = s_csamul_cla32_fa28_4_xor0 & s_csamul_cla32_fa28_3_or0;
  assign s_csamul_cla32_fa28_4_or0 = s_csamul_cla32_fa28_4_and0 | s_csamul_cla32_fa28_4_and1;
  assign s_csamul_cla32_and29_4 = a[29] & b[4];
  assign s_csamul_cla32_fa29_4_xor0 = s_csamul_cla32_and29_4 ^ s_csamul_cla32_fa30_3_xor1;
  assign s_csamul_cla32_fa29_4_and0 = s_csamul_cla32_and29_4 & s_csamul_cla32_fa30_3_xor1;
  assign s_csamul_cla32_fa29_4_xor1 = s_csamul_cla32_fa29_4_xor0 ^ s_csamul_cla32_fa29_3_or0;
  assign s_csamul_cla32_fa29_4_and1 = s_csamul_cla32_fa29_4_xor0 & s_csamul_cla32_fa29_3_or0;
  assign s_csamul_cla32_fa29_4_or0 = s_csamul_cla32_fa29_4_and0 | s_csamul_cla32_fa29_4_and1;
  assign s_csamul_cla32_and30_4 = a[30] & b[4];
  assign s_csamul_cla32_fa30_4_xor0 = s_csamul_cla32_and30_4 ^ s_csamul_cla32_ha31_3_xor0;
  assign s_csamul_cla32_fa30_4_and0 = s_csamul_cla32_and30_4 & s_csamul_cla32_ha31_3_xor0;
  assign s_csamul_cla32_fa30_4_xor1 = s_csamul_cla32_fa30_4_xor0 ^ s_csamul_cla32_fa30_3_or0;
  assign s_csamul_cla32_fa30_4_and1 = s_csamul_cla32_fa30_4_xor0 & s_csamul_cla32_fa30_3_or0;
  assign s_csamul_cla32_fa30_4_or0 = s_csamul_cla32_fa30_4_and0 | s_csamul_cla32_fa30_4_and1;
  assign s_csamul_cla32_nand31_4 = ~(a[31] & b[4]);
  assign s_csamul_cla32_ha31_4_xor0 = s_csamul_cla32_nand31_4 ^ s_csamul_cla32_ha31_3_and0;
  assign s_csamul_cla32_ha31_4_and0 = s_csamul_cla32_nand31_4 & s_csamul_cla32_ha31_3_and0;
  assign s_csamul_cla32_and0_5 = a[0] & b[5];
  assign s_csamul_cla32_fa0_5_xor0 = s_csamul_cla32_and0_5 ^ s_csamul_cla32_fa1_4_xor1;
  assign s_csamul_cla32_fa0_5_and0 = s_csamul_cla32_and0_5 & s_csamul_cla32_fa1_4_xor1;
  assign s_csamul_cla32_fa0_5_xor1 = s_csamul_cla32_fa0_5_xor0 ^ s_csamul_cla32_fa0_4_or0;
  assign s_csamul_cla32_fa0_5_and1 = s_csamul_cla32_fa0_5_xor0 & s_csamul_cla32_fa0_4_or0;
  assign s_csamul_cla32_fa0_5_or0 = s_csamul_cla32_fa0_5_and0 | s_csamul_cla32_fa0_5_and1;
  assign s_csamul_cla32_and1_5 = a[1] & b[5];
  assign s_csamul_cla32_fa1_5_xor0 = s_csamul_cla32_and1_5 ^ s_csamul_cla32_fa2_4_xor1;
  assign s_csamul_cla32_fa1_5_and0 = s_csamul_cla32_and1_5 & s_csamul_cla32_fa2_4_xor1;
  assign s_csamul_cla32_fa1_5_xor1 = s_csamul_cla32_fa1_5_xor0 ^ s_csamul_cla32_fa1_4_or0;
  assign s_csamul_cla32_fa1_5_and1 = s_csamul_cla32_fa1_5_xor0 & s_csamul_cla32_fa1_4_or0;
  assign s_csamul_cla32_fa1_5_or0 = s_csamul_cla32_fa1_5_and0 | s_csamul_cla32_fa1_5_and1;
  assign s_csamul_cla32_and2_5 = a[2] & b[5];
  assign s_csamul_cla32_fa2_5_xor0 = s_csamul_cla32_and2_5 ^ s_csamul_cla32_fa3_4_xor1;
  assign s_csamul_cla32_fa2_5_and0 = s_csamul_cla32_and2_5 & s_csamul_cla32_fa3_4_xor1;
  assign s_csamul_cla32_fa2_5_xor1 = s_csamul_cla32_fa2_5_xor0 ^ s_csamul_cla32_fa2_4_or0;
  assign s_csamul_cla32_fa2_5_and1 = s_csamul_cla32_fa2_5_xor0 & s_csamul_cla32_fa2_4_or0;
  assign s_csamul_cla32_fa2_5_or0 = s_csamul_cla32_fa2_5_and0 | s_csamul_cla32_fa2_5_and1;
  assign s_csamul_cla32_and3_5 = a[3] & b[5];
  assign s_csamul_cla32_fa3_5_xor0 = s_csamul_cla32_and3_5 ^ s_csamul_cla32_fa4_4_xor1;
  assign s_csamul_cla32_fa3_5_and0 = s_csamul_cla32_and3_5 & s_csamul_cla32_fa4_4_xor1;
  assign s_csamul_cla32_fa3_5_xor1 = s_csamul_cla32_fa3_5_xor0 ^ s_csamul_cla32_fa3_4_or0;
  assign s_csamul_cla32_fa3_5_and1 = s_csamul_cla32_fa3_5_xor0 & s_csamul_cla32_fa3_4_or0;
  assign s_csamul_cla32_fa3_5_or0 = s_csamul_cla32_fa3_5_and0 | s_csamul_cla32_fa3_5_and1;
  assign s_csamul_cla32_and4_5 = a[4] & b[5];
  assign s_csamul_cla32_fa4_5_xor0 = s_csamul_cla32_and4_5 ^ s_csamul_cla32_fa5_4_xor1;
  assign s_csamul_cla32_fa4_5_and0 = s_csamul_cla32_and4_5 & s_csamul_cla32_fa5_4_xor1;
  assign s_csamul_cla32_fa4_5_xor1 = s_csamul_cla32_fa4_5_xor0 ^ s_csamul_cla32_fa4_4_or0;
  assign s_csamul_cla32_fa4_5_and1 = s_csamul_cla32_fa4_5_xor0 & s_csamul_cla32_fa4_4_or0;
  assign s_csamul_cla32_fa4_5_or0 = s_csamul_cla32_fa4_5_and0 | s_csamul_cla32_fa4_5_and1;
  assign s_csamul_cla32_and5_5 = a[5] & b[5];
  assign s_csamul_cla32_fa5_5_xor0 = s_csamul_cla32_and5_5 ^ s_csamul_cla32_fa6_4_xor1;
  assign s_csamul_cla32_fa5_5_and0 = s_csamul_cla32_and5_5 & s_csamul_cla32_fa6_4_xor1;
  assign s_csamul_cla32_fa5_5_xor1 = s_csamul_cla32_fa5_5_xor0 ^ s_csamul_cla32_fa5_4_or0;
  assign s_csamul_cla32_fa5_5_and1 = s_csamul_cla32_fa5_5_xor0 & s_csamul_cla32_fa5_4_or0;
  assign s_csamul_cla32_fa5_5_or0 = s_csamul_cla32_fa5_5_and0 | s_csamul_cla32_fa5_5_and1;
  assign s_csamul_cla32_and6_5 = a[6] & b[5];
  assign s_csamul_cla32_fa6_5_xor0 = s_csamul_cla32_and6_5 ^ s_csamul_cla32_fa7_4_xor1;
  assign s_csamul_cla32_fa6_5_and0 = s_csamul_cla32_and6_5 & s_csamul_cla32_fa7_4_xor1;
  assign s_csamul_cla32_fa6_5_xor1 = s_csamul_cla32_fa6_5_xor0 ^ s_csamul_cla32_fa6_4_or0;
  assign s_csamul_cla32_fa6_5_and1 = s_csamul_cla32_fa6_5_xor0 & s_csamul_cla32_fa6_4_or0;
  assign s_csamul_cla32_fa6_5_or0 = s_csamul_cla32_fa6_5_and0 | s_csamul_cla32_fa6_5_and1;
  assign s_csamul_cla32_and7_5 = a[7] & b[5];
  assign s_csamul_cla32_fa7_5_xor0 = s_csamul_cla32_and7_5 ^ s_csamul_cla32_fa8_4_xor1;
  assign s_csamul_cla32_fa7_5_and0 = s_csamul_cla32_and7_5 & s_csamul_cla32_fa8_4_xor1;
  assign s_csamul_cla32_fa7_5_xor1 = s_csamul_cla32_fa7_5_xor0 ^ s_csamul_cla32_fa7_4_or0;
  assign s_csamul_cla32_fa7_5_and1 = s_csamul_cla32_fa7_5_xor0 & s_csamul_cla32_fa7_4_or0;
  assign s_csamul_cla32_fa7_5_or0 = s_csamul_cla32_fa7_5_and0 | s_csamul_cla32_fa7_5_and1;
  assign s_csamul_cla32_and8_5 = a[8] & b[5];
  assign s_csamul_cla32_fa8_5_xor0 = s_csamul_cla32_and8_5 ^ s_csamul_cla32_fa9_4_xor1;
  assign s_csamul_cla32_fa8_5_and0 = s_csamul_cla32_and8_5 & s_csamul_cla32_fa9_4_xor1;
  assign s_csamul_cla32_fa8_5_xor1 = s_csamul_cla32_fa8_5_xor0 ^ s_csamul_cla32_fa8_4_or0;
  assign s_csamul_cla32_fa8_5_and1 = s_csamul_cla32_fa8_5_xor0 & s_csamul_cla32_fa8_4_or0;
  assign s_csamul_cla32_fa8_5_or0 = s_csamul_cla32_fa8_5_and0 | s_csamul_cla32_fa8_5_and1;
  assign s_csamul_cla32_and9_5 = a[9] & b[5];
  assign s_csamul_cla32_fa9_5_xor0 = s_csamul_cla32_and9_5 ^ s_csamul_cla32_fa10_4_xor1;
  assign s_csamul_cla32_fa9_5_and0 = s_csamul_cla32_and9_5 & s_csamul_cla32_fa10_4_xor1;
  assign s_csamul_cla32_fa9_5_xor1 = s_csamul_cla32_fa9_5_xor0 ^ s_csamul_cla32_fa9_4_or0;
  assign s_csamul_cla32_fa9_5_and1 = s_csamul_cla32_fa9_5_xor0 & s_csamul_cla32_fa9_4_or0;
  assign s_csamul_cla32_fa9_5_or0 = s_csamul_cla32_fa9_5_and0 | s_csamul_cla32_fa9_5_and1;
  assign s_csamul_cla32_and10_5 = a[10] & b[5];
  assign s_csamul_cla32_fa10_5_xor0 = s_csamul_cla32_and10_5 ^ s_csamul_cla32_fa11_4_xor1;
  assign s_csamul_cla32_fa10_5_and0 = s_csamul_cla32_and10_5 & s_csamul_cla32_fa11_4_xor1;
  assign s_csamul_cla32_fa10_5_xor1 = s_csamul_cla32_fa10_5_xor0 ^ s_csamul_cla32_fa10_4_or0;
  assign s_csamul_cla32_fa10_5_and1 = s_csamul_cla32_fa10_5_xor0 & s_csamul_cla32_fa10_4_or0;
  assign s_csamul_cla32_fa10_5_or0 = s_csamul_cla32_fa10_5_and0 | s_csamul_cla32_fa10_5_and1;
  assign s_csamul_cla32_and11_5 = a[11] & b[5];
  assign s_csamul_cla32_fa11_5_xor0 = s_csamul_cla32_and11_5 ^ s_csamul_cla32_fa12_4_xor1;
  assign s_csamul_cla32_fa11_5_and0 = s_csamul_cla32_and11_5 & s_csamul_cla32_fa12_4_xor1;
  assign s_csamul_cla32_fa11_5_xor1 = s_csamul_cla32_fa11_5_xor0 ^ s_csamul_cla32_fa11_4_or0;
  assign s_csamul_cla32_fa11_5_and1 = s_csamul_cla32_fa11_5_xor0 & s_csamul_cla32_fa11_4_or0;
  assign s_csamul_cla32_fa11_5_or0 = s_csamul_cla32_fa11_5_and0 | s_csamul_cla32_fa11_5_and1;
  assign s_csamul_cla32_and12_5 = a[12] & b[5];
  assign s_csamul_cla32_fa12_5_xor0 = s_csamul_cla32_and12_5 ^ s_csamul_cla32_fa13_4_xor1;
  assign s_csamul_cla32_fa12_5_and0 = s_csamul_cla32_and12_5 & s_csamul_cla32_fa13_4_xor1;
  assign s_csamul_cla32_fa12_5_xor1 = s_csamul_cla32_fa12_5_xor0 ^ s_csamul_cla32_fa12_4_or0;
  assign s_csamul_cla32_fa12_5_and1 = s_csamul_cla32_fa12_5_xor0 & s_csamul_cla32_fa12_4_or0;
  assign s_csamul_cla32_fa12_5_or0 = s_csamul_cla32_fa12_5_and0 | s_csamul_cla32_fa12_5_and1;
  assign s_csamul_cla32_and13_5 = a[13] & b[5];
  assign s_csamul_cla32_fa13_5_xor0 = s_csamul_cla32_and13_5 ^ s_csamul_cla32_fa14_4_xor1;
  assign s_csamul_cla32_fa13_5_and0 = s_csamul_cla32_and13_5 & s_csamul_cla32_fa14_4_xor1;
  assign s_csamul_cla32_fa13_5_xor1 = s_csamul_cla32_fa13_5_xor0 ^ s_csamul_cla32_fa13_4_or0;
  assign s_csamul_cla32_fa13_5_and1 = s_csamul_cla32_fa13_5_xor0 & s_csamul_cla32_fa13_4_or0;
  assign s_csamul_cla32_fa13_5_or0 = s_csamul_cla32_fa13_5_and0 | s_csamul_cla32_fa13_5_and1;
  assign s_csamul_cla32_and14_5 = a[14] & b[5];
  assign s_csamul_cla32_fa14_5_xor0 = s_csamul_cla32_and14_5 ^ s_csamul_cla32_fa15_4_xor1;
  assign s_csamul_cla32_fa14_5_and0 = s_csamul_cla32_and14_5 & s_csamul_cla32_fa15_4_xor1;
  assign s_csamul_cla32_fa14_5_xor1 = s_csamul_cla32_fa14_5_xor0 ^ s_csamul_cla32_fa14_4_or0;
  assign s_csamul_cla32_fa14_5_and1 = s_csamul_cla32_fa14_5_xor0 & s_csamul_cla32_fa14_4_or0;
  assign s_csamul_cla32_fa14_5_or0 = s_csamul_cla32_fa14_5_and0 | s_csamul_cla32_fa14_5_and1;
  assign s_csamul_cla32_and15_5 = a[15] & b[5];
  assign s_csamul_cla32_fa15_5_xor0 = s_csamul_cla32_and15_5 ^ s_csamul_cla32_fa16_4_xor1;
  assign s_csamul_cla32_fa15_5_and0 = s_csamul_cla32_and15_5 & s_csamul_cla32_fa16_4_xor1;
  assign s_csamul_cla32_fa15_5_xor1 = s_csamul_cla32_fa15_5_xor0 ^ s_csamul_cla32_fa15_4_or0;
  assign s_csamul_cla32_fa15_5_and1 = s_csamul_cla32_fa15_5_xor0 & s_csamul_cla32_fa15_4_or0;
  assign s_csamul_cla32_fa15_5_or0 = s_csamul_cla32_fa15_5_and0 | s_csamul_cla32_fa15_5_and1;
  assign s_csamul_cla32_and16_5 = a[16] & b[5];
  assign s_csamul_cla32_fa16_5_xor0 = s_csamul_cla32_and16_5 ^ s_csamul_cla32_fa17_4_xor1;
  assign s_csamul_cla32_fa16_5_and0 = s_csamul_cla32_and16_5 & s_csamul_cla32_fa17_4_xor1;
  assign s_csamul_cla32_fa16_5_xor1 = s_csamul_cla32_fa16_5_xor0 ^ s_csamul_cla32_fa16_4_or0;
  assign s_csamul_cla32_fa16_5_and1 = s_csamul_cla32_fa16_5_xor0 & s_csamul_cla32_fa16_4_or0;
  assign s_csamul_cla32_fa16_5_or0 = s_csamul_cla32_fa16_5_and0 | s_csamul_cla32_fa16_5_and1;
  assign s_csamul_cla32_and17_5 = a[17] & b[5];
  assign s_csamul_cla32_fa17_5_xor0 = s_csamul_cla32_and17_5 ^ s_csamul_cla32_fa18_4_xor1;
  assign s_csamul_cla32_fa17_5_and0 = s_csamul_cla32_and17_5 & s_csamul_cla32_fa18_4_xor1;
  assign s_csamul_cla32_fa17_5_xor1 = s_csamul_cla32_fa17_5_xor0 ^ s_csamul_cla32_fa17_4_or0;
  assign s_csamul_cla32_fa17_5_and1 = s_csamul_cla32_fa17_5_xor0 & s_csamul_cla32_fa17_4_or0;
  assign s_csamul_cla32_fa17_5_or0 = s_csamul_cla32_fa17_5_and0 | s_csamul_cla32_fa17_5_and1;
  assign s_csamul_cla32_and18_5 = a[18] & b[5];
  assign s_csamul_cla32_fa18_5_xor0 = s_csamul_cla32_and18_5 ^ s_csamul_cla32_fa19_4_xor1;
  assign s_csamul_cla32_fa18_5_and0 = s_csamul_cla32_and18_5 & s_csamul_cla32_fa19_4_xor1;
  assign s_csamul_cla32_fa18_5_xor1 = s_csamul_cla32_fa18_5_xor0 ^ s_csamul_cla32_fa18_4_or0;
  assign s_csamul_cla32_fa18_5_and1 = s_csamul_cla32_fa18_5_xor0 & s_csamul_cla32_fa18_4_or0;
  assign s_csamul_cla32_fa18_5_or0 = s_csamul_cla32_fa18_5_and0 | s_csamul_cla32_fa18_5_and1;
  assign s_csamul_cla32_and19_5 = a[19] & b[5];
  assign s_csamul_cla32_fa19_5_xor0 = s_csamul_cla32_and19_5 ^ s_csamul_cla32_fa20_4_xor1;
  assign s_csamul_cla32_fa19_5_and0 = s_csamul_cla32_and19_5 & s_csamul_cla32_fa20_4_xor1;
  assign s_csamul_cla32_fa19_5_xor1 = s_csamul_cla32_fa19_5_xor0 ^ s_csamul_cla32_fa19_4_or0;
  assign s_csamul_cla32_fa19_5_and1 = s_csamul_cla32_fa19_5_xor0 & s_csamul_cla32_fa19_4_or0;
  assign s_csamul_cla32_fa19_5_or0 = s_csamul_cla32_fa19_5_and0 | s_csamul_cla32_fa19_5_and1;
  assign s_csamul_cla32_and20_5 = a[20] & b[5];
  assign s_csamul_cla32_fa20_5_xor0 = s_csamul_cla32_and20_5 ^ s_csamul_cla32_fa21_4_xor1;
  assign s_csamul_cla32_fa20_5_and0 = s_csamul_cla32_and20_5 & s_csamul_cla32_fa21_4_xor1;
  assign s_csamul_cla32_fa20_5_xor1 = s_csamul_cla32_fa20_5_xor0 ^ s_csamul_cla32_fa20_4_or0;
  assign s_csamul_cla32_fa20_5_and1 = s_csamul_cla32_fa20_5_xor0 & s_csamul_cla32_fa20_4_or0;
  assign s_csamul_cla32_fa20_5_or0 = s_csamul_cla32_fa20_5_and0 | s_csamul_cla32_fa20_5_and1;
  assign s_csamul_cla32_and21_5 = a[21] & b[5];
  assign s_csamul_cla32_fa21_5_xor0 = s_csamul_cla32_and21_5 ^ s_csamul_cla32_fa22_4_xor1;
  assign s_csamul_cla32_fa21_5_and0 = s_csamul_cla32_and21_5 & s_csamul_cla32_fa22_4_xor1;
  assign s_csamul_cla32_fa21_5_xor1 = s_csamul_cla32_fa21_5_xor0 ^ s_csamul_cla32_fa21_4_or0;
  assign s_csamul_cla32_fa21_5_and1 = s_csamul_cla32_fa21_5_xor0 & s_csamul_cla32_fa21_4_or0;
  assign s_csamul_cla32_fa21_5_or0 = s_csamul_cla32_fa21_5_and0 | s_csamul_cla32_fa21_5_and1;
  assign s_csamul_cla32_and22_5 = a[22] & b[5];
  assign s_csamul_cla32_fa22_5_xor0 = s_csamul_cla32_and22_5 ^ s_csamul_cla32_fa23_4_xor1;
  assign s_csamul_cla32_fa22_5_and0 = s_csamul_cla32_and22_5 & s_csamul_cla32_fa23_4_xor1;
  assign s_csamul_cla32_fa22_5_xor1 = s_csamul_cla32_fa22_5_xor0 ^ s_csamul_cla32_fa22_4_or0;
  assign s_csamul_cla32_fa22_5_and1 = s_csamul_cla32_fa22_5_xor0 & s_csamul_cla32_fa22_4_or0;
  assign s_csamul_cla32_fa22_5_or0 = s_csamul_cla32_fa22_5_and0 | s_csamul_cla32_fa22_5_and1;
  assign s_csamul_cla32_and23_5 = a[23] & b[5];
  assign s_csamul_cla32_fa23_5_xor0 = s_csamul_cla32_and23_5 ^ s_csamul_cla32_fa24_4_xor1;
  assign s_csamul_cla32_fa23_5_and0 = s_csamul_cla32_and23_5 & s_csamul_cla32_fa24_4_xor1;
  assign s_csamul_cla32_fa23_5_xor1 = s_csamul_cla32_fa23_5_xor0 ^ s_csamul_cla32_fa23_4_or0;
  assign s_csamul_cla32_fa23_5_and1 = s_csamul_cla32_fa23_5_xor0 & s_csamul_cla32_fa23_4_or0;
  assign s_csamul_cla32_fa23_5_or0 = s_csamul_cla32_fa23_5_and0 | s_csamul_cla32_fa23_5_and1;
  assign s_csamul_cla32_and24_5 = a[24] & b[5];
  assign s_csamul_cla32_fa24_5_xor0 = s_csamul_cla32_and24_5 ^ s_csamul_cla32_fa25_4_xor1;
  assign s_csamul_cla32_fa24_5_and0 = s_csamul_cla32_and24_5 & s_csamul_cla32_fa25_4_xor1;
  assign s_csamul_cla32_fa24_5_xor1 = s_csamul_cla32_fa24_5_xor0 ^ s_csamul_cla32_fa24_4_or0;
  assign s_csamul_cla32_fa24_5_and1 = s_csamul_cla32_fa24_5_xor0 & s_csamul_cla32_fa24_4_or0;
  assign s_csamul_cla32_fa24_5_or0 = s_csamul_cla32_fa24_5_and0 | s_csamul_cla32_fa24_5_and1;
  assign s_csamul_cla32_and25_5 = a[25] & b[5];
  assign s_csamul_cla32_fa25_5_xor0 = s_csamul_cla32_and25_5 ^ s_csamul_cla32_fa26_4_xor1;
  assign s_csamul_cla32_fa25_5_and0 = s_csamul_cla32_and25_5 & s_csamul_cla32_fa26_4_xor1;
  assign s_csamul_cla32_fa25_5_xor1 = s_csamul_cla32_fa25_5_xor0 ^ s_csamul_cla32_fa25_4_or0;
  assign s_csamul_cla32_fa25_5_and1 = s_csamul_cla32_fa25_5_xor0 & s_csamul_cla32_fa25_4_or0;
  assign s_csamul_cla32_fa25_5_or0 = s_csamul_cla32_fa25_5_and0 | s_csamul_cla32_fa25_5_and1;
  assign s_csamul_cla32_and26_5 = a[26] & b[5];
  assign s_csamul_cla32_fa26_5_xor0 = s_csamul_cla32_and26_5 ^ s_csamul_cla32_fa27_4_xor1;
  assign s_csamul_cla32_fa26_5_and0 = s_csamul_cla32_and26_5 & s_csamul_cla32_fa27_4_xor1;
  assign s_csamul_cla32_fa26_5_xor1 = s_csamul_cla32_fa26_5_xor0 ^ s_csamul_cla32_fa26_4_or0;
  assign s_csamul_cla32_fa26_5_and1 = s_csamul_cla32_fa26_5_xor0 & s_csamul_cla32_fa26_4_or0;
  assign s_csamul_cla32_fa26_5_or0 = s_csamul_cla32_fa26_5_and0 | s_csamul_cla32_fa26_5_and1;
  assign s_csamul_cla32_and27_5 = a[27] & b[5];
  assign s_csamul_cla32_fa27_5_xor0 = s_csamul_cla32_and27_5 ^ s_csamul_cla32_fa28_4_xor1;
  assign s_csamul_cla32_fa27_5_and0 = s_csamul_cla32_and27_5 & s_csamul_cla32_fa28_4_xor1;
  assign s_csamul_cla32_fa27_5_xor1 = s_csamul_cla32_fa27_5_xor0 ^ s_csamul_cla32_fa27_4_or0;
  assign s_csamul_cla32_fa27_5_and1 = s_csamul_cla32_fa27_5_xor0 & s_csamul_cla32_fa27_4_or0;
  assign s_csamul_cla32_fa27_5_or0 = s_csamul_cla32_fa27_5_and0 | s_csamul_cla32_fa27_5_and1;
  assign s_csamul_cla32_and28_5 = a[28] & b[5];
  assign s_csamul_cla32_fa28_5_xor0 = s_csamul_cla32_and28_5 ^ s_csamul_cla32_fa29_4_xor1;
  assign s_csamul_cla32_fa28_5_and0 = s_csamul_cla32_and28_5 & s_csamul_cla32_fa29_4_xor1;
  assign s_csamul_cla32_fa28_5_xor1 = s_csamul_cla32_fa28_5_xor0 ^ s_csamul_cla32_fa28_4_or0;
  assign s_csamul_cla32_fa28_5_and1 = s_csamul_cla32_fa28_5_xor0 & s_csamul_cla32_fa28_4_or0;
  assign s_csamul_cla32_fa28_5_or0 = s_csamul_cla32_fa28_5_and0 | s_csamul_cla32_fa28_5_and1;
  assign s_csamul_cla32_and29_5 = a[29] & b[5];
  assign s_csamul_cla32_fa29_5_xor0 = s_csamul_cla32_and29_5 ^ s_csamul_cla32_fa30_4_xor1;
  assign s_csamul_cla32_fa29_5_and0 = s_csamul_cla32_and29_5 & s_csamul_cla32_fa30_4_xor1;
  assign s_csamul_cla32_fa29_5_xor1 = s_csamul_cla32_fa29_5_xor0 ^ s_csamul_cla32_fa29_4_or0;
  assign s_csamul_cla32_fa29_5_and1 = s_csamul_cla32_fa29_5_xor0 & s_csamul_cla32_fa29_4_or0;
  assign s_csamul_cla32_fa29_5_or0 = s_csamul_cla32_fa29_5_and0 | s_csamul_cla32_fa29_5_and1;
  assign s_csamul_cla32_and30_5 = a[30] & b[5];
  assign s_csamul_cla32_fa30_5_xor0 = s_csamul_cla32_and30_5 ^ s_csamul_cla32_ha31_4_xor0;
  assign s_csamul_cla32_fa30_5_and0 = s_csamul_cla32_and30_5 & s_csamul_cla32_ha31_4_xor0;
  assign s_csamul_cla32_fa30_5_xor1 = s_csamul_cla32_fa30_5_xor0 ^ s_csamul_cla32_fa30_4_or0;
  assign s_csamul_cla32_fa30_5_and1 = s_csamul_cla32_fa30_5_xor0 & s_csamul_cla32_fa30_4_or0;
  assign s_csamul_cla32_fa30_5_or0 = s_csamul_cla32_fa30_5_and0 | s_csamul_cla32_fa30_5_and1;
  assign s_csamul_cla32_nand31_5 = ~(a[31] & b[5]);
  assign s_csamul_cla32_ha31_5_xor0 = s_csamul_cla32_nand31_5 ^ s_csamul_cla32_ha31_4_and0;
  assign s_csamul_cla32_ha31_5_and0 = s_csamul_cla32_nand31_5 & s_csamul_cla32_ha31_4_and0;
  assign s_csamul_cla32_and0_6 = a[0] & b[6];
  assign s_csamul_cla32_fa0_6_xor0 = s_csamul_cla32_and0_6 ^ s_csamul_cla32_fa1_5_xor1;
  assign s_csamul_cla32_fa0_6_and0 = s_csamul_cla32_and0_6 & s_csamul_cla32_fa1_5_xor1;
  assign s_csamul_cla32_fa0_6_xor1 = s_csamul_cla32_fa0_6_xor0 ^ s_csamul_cla32_fa0_5_or0;
  assign s_csamul_cla32_fa0_6_and1 = s_csamul_cla32_fa0_6_xor0 & s_csamul_cla32_fa0_5_or0;
  assign s_csamul_cla32_fa0_6_or0 = s_csamul_cla32_fa0_6_and0 | s_csamul_cla32_fa0_6_and1;
  assign s_csamul_cla32_and1_6 = a[1] & b[6];
  assign s_csamul_cla32_fa1_6_xor0 = s_csamul_cla32_and1_6 ^ s_csamul_cla32_fa2_5_xor1;
  assign s_csamul_cla32_fa1_6_and0 = s_csamul_cla32_and1_6 & s_csamul_cla32_fa2_5_xor1;
  assign s_csamul_cla32_fa1_6_xor1 = s_csamul_cla32_fa1_6_xor0 ^ s_csamul_cla32_fa1_5_or0;
  assign s_csamul_cla32_fa1_6_and1 = s_csamul_cla32_fa1_6_xor0 & s_csamul_cla32_fa1_5_or0;
  assign s_csamul_cla32_fa1_6_or0 = s_csamul_cla32_fa1_6_and0 | s_csamul_cla32_fa1_6_and1;
  assign s_csamul_cla32_and2_6 = a[2] & b[6];
  assign s_csamul_cla32_fa2_6_xor0 = s_csamul_cla32_and2_6 ^ s_csamul_cla32_fa3_5_xor1;
  assign s_csamul_cla32_fa2_6_and0 = s_csamul_cla32_and2_6 & s_csamul_cla32_fa3_5_xor1;
  assign s_csamul_cla32_fa2_6_xor1 = s_csamul_cla32_fa2_6_xor0 ^ s_csamul_cla32_fa2_5_or0;
  assign s_csamul_cla32_fa2_6_and1 = s_csamul_cla32_fa2_6_xor0 & s_csamul_cla32_fa2_5_or0;
  assign s_csamul_cla32_fa2_6_or0 = s_csamul_cla32_fa2_6_and0 | s_csamul_cla32_fa2_6_and1;
  assign s_csamul_cla32_and3_6 = a[3] & b[6];
  assign s_csamul_cla32_fa3_6_xor0 = s_csamul_cla32_and3_6 ^ s_csamul_cla32_fa4_5_xor1;
  assign s_csamul_cla32_fa3_6_and0 = s_csamul_cla32_and3_6 & s_csamul_cla32_fa4_5_xor1;
  assign s_csamul_cla32_fa3_6_xor1 = s_csamul_cla32_fa3_6_xor0 ^ s_csamul_cla32_fa3_5_or0;
  assign s_csamul_cla32_fa3_6_and1 = s_csamul_cla32_fa3_6_xor0 & s_csamul_cla32_fa3_5_or0;
  assign s_csamul_cla32_fa3_6_or0 = s_csamul_cla32_fa3_6_and0 | s_csamul_cla32_fa3_6_and1;
  assign s_csamul_cla32_and4_6 = a[4] & b[6];
  assign s_csamul_cla32_fa4_6_xor0 = s_csamul_cla32_and4_6 ^ s_csamul_cla32_fa5_5_xor1;
  assign s_csamul_cla32_fa4_6_and0 = s_csamul_cla32_and4_6 & s_csamul_cla32_fa5_5_xor1;
  assign s_csamul_cla32_fa4_6_xor1 = s_csamul_cla32_fa4_6_xor0 ^ s_csamul_cla32_fa4_5_or0;
  assign s_csamul_cla32_fa4_6_and1 = s_csamul_cla32_fa4_6_xor0 & s_csamul_cla32_fa4_5_or0;
  assign s_csamul_cla32_fa4_6_or0 = s_csamul_cla32_fa4_6_and0 | s_csamul_cla32_fa4_6_and1;
  assign s_csamul_cla32_and5_6 = a[5] & b[6];
  assign s_csamul_cla32_fa5_6_xor0 = s_csamul_cla32_and5_6 ^ s_csamul_cla32_fa6_5_xor1;
  assign s_csamul_cla32_fa5_6_and0 = s_csamul_cla32_and5_6 & s_csamul_cla32_fa6_5_xor1;
  assign s_csamul_cla32_fa5_6_xor1 = s_csamul_cla32_fa5_6_xor0 ^ s_csamul_cla32_fa5_5_or0;
  assign s_csamul_cla32_fa5_6_and1 = s_csamul_cla32_fa5_6_xor0 & s_csamul_cla32_fa5_5_or0;
  assign s_csamul_cla32_fa5_6_or0 = s_csamul_cla32_fa5_6_and0 | s_csamul_cla32_fa5_6_and1;
  assign s_csamul_cla32_and6_6 = a[6] & b[6];
  assign s_csamul_cla32_fa6_6_xor0 = s_csamul_cla32_and6_6 ^ s_csamul_cla32_fa7_5_xor1;
  assign s_csamul_cla32_fa6_6_and0 = s_csamul_cla32_and6_6 & s_csamul_cla32_fa7_5_xor1;
  assign s_csamul_cla32_fa6_6_xor1 = s_csamul_cla32_fa6_6_xor0 ^ s_csamul_cla32_fa6_5_or0;
  assign s_csamul_cla32_fa6_6_and1 = s_csamul_cla32_fa6_6_xor0 & s_csamul_cla32_fa6_5_or0;
  assign s_csamul_cla32_fa6_6_or0 = s_csamul_cla32_fa6_6_and0 | s_csamul_cla32_fa6_6_and1;
  assign s_csamul_cla32_and7_6 = a[7] & b[6];
  assign s_csamul_cla32_fa7_6_xor0 = s_csamul_cla32_and7_6 ^ s_csamul_cla32_fa8_5_xor1;
  assign s_csamul_cla32_fa7_6_and0 = s_csamul_cla32_and7_6 & s_csamul_cla32_fa8_5_xor1;
  assign s_csamul_cla32_fa7_6_xor1 = s_csamul_cla32_fa7_6_xor0 ^ s_csamul_cla32_fa7_5_or0;
  assign s_csamul_cla32_fa7_6_and1 = s_csamul_cla32_fa7_6_xor0 & s_csamul_cla32_fa7_5_or0;
  assign s_csamul_cla32_fa7_6_or0 = s_csamul_cla32_fa7_6_and0 | s_csamul_cla32_fa7_6_and1;
  assign s_csamul_cla32_and8_6 = a[8] & b[6];
  assign s_csamul_cla32_fa8_6_xor0 = s_csamul_cla32_and8_6 ^ s_csamul_cla32_fa9_5_xor1;
  assign s_csamul_cla32_fa8_6_and0 = s_csamul_cla32_and8_6 & s_csamul_cla32_fa9_5_xor1;
  assign s_csamul_cla32_fa8_6_xor1 = s_csamul_cla32_fa8_6_xor0 ^ s_csamul_cla32_fa8_5_or0;
  assign s_csamul_cla32_fa8_6_and1 = s_csamul_cla32_fa8_6_xor0 & s_csamul_cla32_fa8_5_or0;
  assign s_csamul_cla32_fa8_6_or0 = s_csamul_cla32_fa8_6_and0 | s_csamul_cla32_fa8_6_and1;
  assign s_csamul_cla32_and9_6 = a[9] & b[6];
  assign s_csamul_cla32_fa9_6_xor0 = s_csamul_cla32_and9_6 ^ s_csamul_cla32_fa10_5_xor1;
  assign s_csamul_cla32_fa9_6_and0 = s_csamul_cla32_and9_6 & s_csamul_cla32_fa10_5_xor1;
  assign s_csamul_cla32_fa9_6_xor1 = s_csamul_cla32_fa9_6_xor0 ^ s_csamul_cla32_fa9_5_or0;
  assign s_csamul_cla32_fa9_6_and1 = s_csamul_cla32_fa9_6_xor0 & s_csamul_cla32_fa9_5_or0;
  assign s_csamul_cla32_fa9_6_or0 = s_csamul_cla32_fa9_6_and0 | s_csamul_cla32_fa9_6_and1;
  assign s_csamul_cla32_and10_6 = a[10] & b[6];
  assign s_csamul_cla32_fa10_6_xor0 = s_csamul_cla32_and10_6 ^ s_csamul_cla32_fa11_5_xor1;
  assign s_csamul_cla32_fa10_6_and0 = s_csamul_cla32_and10_6 & s_csamul_cla32_fa11_5_xor1;
  assign s_csamul_cla32_fa10_6_xor1 = s_csamul_cla32_fa10_6_xor0 ^ s_csamul_cla32_fa10_5_or0;
  assign s_csamul_cla32_fa10_6_and1 = s_csamul_cla32_fa10_6_xor0 & s_csamul_cla32_fa10_5_or0;
  assign s_csamul_cla32_fa10_6_or0 = s_csamul_cla32_fa10_6_and0 | s_csamul_cla32_fa10_6_and1;
  assign s_csamul_cla32_and11_6 = a[11] & b[6];
  assign s_csamul_cla32_fa11_6_xor0 = s_csamul_cla32_and11_6 ^ s_csamul_cla32_fa12_5_xor1;
  assign s_csamul_cla32_fa11_6_and0 = s_csamul_cla32_and11_6 & s_csamul_cla32_fa12_5_xor1;
  assign s_csamul_cla32_fa11_6_xor1 = s_csamul_cla32_fa11_6_xor0 ^ s_csamul_cla32_fa11_5_or0;
  assign s_csamul_cla32_fa11_6_and1 = s_csamul_cla32_fa11_6_xor0 & s_csamul_cla32_fa11_5_or0;
  assign s_csamul_cla32_fa11_6_or0 = s_csamul_cla32_fa11_6_and0 | s_csamul_cla32_fa11_6_and1;
  assign s_csamul_cla32_and12_6 = a[12] & b[6];
  assign s_csamul_cla32_fa12_6_xor0 = s_csamul_cla32_and12_6 ^ s_csamul_cla32_fa13_5_xor1;
  assign s_csamul_cla32_fa12_6_and0 = s_csamul_cla32_and12_6 & s_csamul_cla32_fa13_5_xor1;
  assign s_csamul_cla32_fa12_6_xor1 = s_csamul_cla32_fa12_6_xor0 ^ s_csamul_cla32_fa12_5_or0;
  assign s_csamul_cla32_fa12_6_and1 = s_csamul_cla32_fa12_6_xor0 & s_csamul_cla32_fa12_5_or0;
  assign s_csamul_cla32_fa12_6_or0 = s_csamul_cla32_fa12_6_and0 | s_csamul_cla32_fa12_6_and1;
  assign s_csamul_cla32_and13_6 = a[13] & b[6];
  assign s_csamul_cla32_fa13_6_xor0 = s_csamul_cla32_and13_6 ^ s_csamul_cla32_fa14_5_xor1;
  assign s_csamul_cla32_fa13_6_and0 = s_csamul_cla32_and13_6 & s_csamul_cla32_fa14_5_xor1;
  assign s_csamul_cla32_fa13_6_xor1 = s_csamul_cla32_fa13_6_xor0 ^ s_csamul_cla32_fa13_5_or0;
  assign s_csamul_cla32_fa13_6_and1 = s_csamul_cla32_fa13_6_xor0 & s_csamul_cla32_fa13_5_or0;
  assign s_csamul_cla32_fa13_6_or0 = s_csamul_cla32_fa13_6_and0 | s_csamul_cla32_fa13_6_and1;
  assign s_csamul_cla32_and14_6 = a[14] & b[6];
  assign s_csamul_cla32_fa14_6_xor0 = s_csamul_cla32_and14_6 ^ s_csamul_cla32_fa15_5_xor1;
  assign s_csamul_cla32_fa14_6_and0 = s_csamul_cla32_and14_6 & s_csamul_cla32_fa15_5_xor1;
  assign s_csamul_cla32_fa14_6_xor1 = s_csamul_cla32_fa14_6_xor0 ^ s_csamul_cla32_fa14_5_or0;
  assign s_csamul_cla32_fa14_6_and1 = s_csamul_cla32_fa14_6_xor0 & s_csamul_cla32_fa14_5_or0;
  assign s_csamul_cla32_fa14_6_or0 = s_csamul_cla32_fa14_6_and0 | s_csamul_cla32_fa14_6_and1;
  assign s_csamul_cla32_and15_6 = a[15] & b[6];
  assign s_csamul_cla32_fa15_6_xor0 = s_csamul_cla32_and15_6 ^ s_csamul_cla32_fa16_5_xor1;
  assign s_csamul_cla32_fa15_6_and0 = s_csamul_cla32_and15_6 & s_csamul_cla32_fa16_5_xor1;
  assign s_csamul_cla32_fa15_6_xor1 = s_csamul_cla32_fa15_6_xor0 ^ s_csamul_cla32_fa15_5_or0;
  assign s_csamul_cla32_fa15_6_and1 = s_csamul_cla32_fa15_6_xor0 & s_csamul_cla32_fa15_5_or0;
  assign s_csamul_cla32_fa15_6_or0 = s_csamul_cla32_fa15_6_and0 | s_csamul_cla32_fa15_6_and1;
  assign s_csamul_cla32_and16_6 = a[16] & b[6];
  assign s_csamul_cla32_fa16_6_xor0 = s_csamul_cla32_and16_6 ^ s_csamul_cla32_fa17_5_xor1;
  assign s_csamul_cla32_fa16_6_and0 = s_csamul_cla32_and16_6 & s_csamul_cla32_fa17_5_xor1;
  assign s_csamul_cla32_fa16_6_xor1 = s_csamul_cla32_fa16_6_xor0 ^ s_csamul_cla32_fa16_5_or0;
  assign s_csamul_cla32_fa16_6_and1 = s_csamul_cla32_fa16_6_xor0 & s_csamul_cla32_fa16_5_or0;
  assign s_csamul_cla32_fa16_6_or0 = s_csamul_cla32_fa16_6_and0 | s_csamul_cla32_fa16_6_and1;
  assign s_csamul_cla32_and17_6 = a[17] & b[6];
  assign s_csamul_cla32_fa17_6_xor0 = s_csamul_cla32_and17_6 ^ s_csamul_cla32_fa18_5_xor1;
  assign s_csamul_cla32_fa17_6_and0 = s_csamul_cla32_and17_6 & s_csamul_cla32_fa18_5_xor1;
  assign s_csamul_cla32_fa17_6_xor1 = s_csamul_cla32_fa17_6_xor0 ^ s_csamul_cla32_fa17_5_or0;
  assign s_csamul_cla32_fa17_6_and1 = s_csamul_cla32_fa17_6_xor0 & s_csamul_cla32_fa17_5_or0;
  assign s_csamul_cla32_fa17_6_or0 = s_csamul_cla32_fa17_6_and0 | s_csamul_cla32_fa17_6_and1;
  assign s_csamul_cla32_and18_6 = a[18] & b[6];
  assign s_csamul_cla32_fa18_6_xor0 = s_csamul_cla32_and18_6 ^ s_csamul_cla32_fa19_5_xor1;
  assign s_csamul_cla32_fa18_6_and0 = s_csamul_cla32_and18_6 & s_csamul_cla32_fa19_5_xor1;
  assign s_csamul_cla32_fa18_6_xor1 = s_csamul_cla32_fa18_6_xor0 ^ s_csamul_cla32_fa18_5_or0;
  assign s_csamul_cla32_fa18_6_and1 = s_csamul_cla32_fa18_6_xor0 & s_csamul_cla32_fa18_5_or0;
  assign s_csamul_cla32_fa18_6_or0 = s_csamul_cla32_fa18_6_and0 | s_csamul_cla32_fa18_6_and1;
  assign s_csamul_cla32_and19_6 = a[19] & b[6];
  assign s_csamul_cla32_fa19_6_xor0 = s_csamul_cla32_and19_6 ^ s_csamul_cla32_fa20_5_xor1;
  assign s_csamul_cla32_fa19_6_and0 = s_csamul_cla32_and19_6 & s_csamul_cla32_fa20_5_xor1;
  assign s_csamul_cla32_fa19_6_xor1 = s_csamul_cla32_fa19_6_xor0 ^ s_csamul_cla32_fa19_5_or0;
  assign s_csamul_cla32_fa19_6_and1 = s_csamul_cla32_fa19_6_xor0 & s_csamul_cla32_fa19_5_or0;
  assign s_csamul_cla32_fa19_6_or0 = s_csamul_cla32_fa19_6_and0 | s_csamul_cla32_fa19_6_and1;
  assign s_csamul_cla32_and20_6 = a[20] & b[6];
  assign s_csamul_cla32_fa20_6_xor0 = s_csamul_cla32_and20_6 ^ s_csamul_cla32_fa21_5_xor1;
  assign s_csamul_cla32_fa20_6_and0 = s_csamul_cla32_and20_6 & s_csamul_cla32_fa21_5_xor1;
  assign s_csamul_cla32_fa20_6_xor1 = s_csamul_cla32_fa20_6_xor0 ^ s_csamul_cla32_fa20_5_or0;
  assign s_csamul_cla32_fa20_6_and1 = s_csamul_cla32_fa20_6_xor0 & s_csamul_cla32_fa20_5_or0;
  assign s_csamul_cla32_fa20_6_or0 = s_csamul_cla32_fa20_6_and0 | s_csamul_cla32_fa20_6_and1;
  assign s_csamul_cla32_and21_6 = a[21] & b[6];
  assign s_csamul_cla32_fa21_6_xor0 = s_csamul_cla32_and21_6 ^ s_csamul_cla32_fa22_5_xor1;
  assign s_csamul_cla32_fa21_6_and0 = s_csamul_cla32_and21_6 & s_csamul_cla32_fa22_5_xor1;
  assign s_csamul_cla32_fa21_6_xor1 = s_csamul_cla32_fa21_6_xor0 ^ s_csamul_cla32_fa21_5_or0;
  assign s_csamul_cla32_fa21_6_and1 = s_csamul_cla32_fa21_6_xor0 & s_csamul_cla32_fa21_5_or0;
  assign s_csamul_cla32_fa21_6_or0 = s_csamul_cla32_fa21_6_and0 | s_csamul_cla32_fa21_6_and1;
  assign s_csamul_cla32_and22_6 = a[22] & b[6];
  assign s_csamul_cla32_fa22_6_xor0 = s_csamul_cla32_and22_6 ^ s_csamul_cla32_fa23_5_xor1;
  assign s_csamul_cla32_fa22_6_and0 = s_csamul_cla32_and22_6 & s_csamul_cla32_fa23_5_xor1;
  assign s_csamul_cla32_fa22_6_xor1 = s_csamul_cla32_fa22_6_xor0 ^ s_csamul_cla32_fa22_5_or0;
  assign s_csamul_cla32_fa22_6_and1 = s_csamul_cla32_fa22_6_xor0 & s_csamul_cla32_fa22_5_or0;
  assign s_csamul_cla32_fa22_6_or0 = s_csamul_cla32_fa22_6_and0 | s_csamul_cla32_fa22_6_and1;
  assign s_csamul_cla32_and23_6 = a[23] & b[6];
  assign s_csamul_cla32_fa23_6_xor0 = s_csamul_cla32_and23_6 ^ s_csamul_cla32_fa24_5_xor1;
  assign s_csamul_cla32_fa23_6_and0 = s_csamul_cla32_and23_6 & s_csamul_cla32_fa24_5_xor1;
  assign s_csamul_cla32_fa23_6_xor1 = s_csamul_cla32_fa23_6_xor0 ^ s_csamul_cla32_fa23_5_or0;
  assign s_csamul_cla32_fa23_6_and1 = s_csamul_cla32_fa23_6_xor0 & s_csamul_cla32_fa23_5_or0;
  assign s_csamul_cla32_fa23_6_or0 = s_csamul_cla32_fa23_6_and0 | s_csamul_cla32_fa23_6_and1;
  assign s_csamul_cla32_and24_6 = a[24] & b[6];
  assign s_csamul_cla32_fa24_6_xor0 = s_csamul_cla32_and24_6 ^ s_csamul_cla32_fa25_5_xor1;
  assign s_csamul_cla32_fa24_6_and0 = s_csamul_cla32_and24_6 & s_csamul_cla32_fa25_5_xor1;
  assign s_csamul_cla32_fa24_6_xor1 = s_csamul_cla32_fa24_6_xor0 ^ s_csamul_cla32_fa24_5_or0;
  assign s_csamul_cla32_fa24_6_and1 = s_csamul_cla32_fa24_6_xor0 & s_csamul_cla32_fa24_5_or0;
  assign s_csamul_cla32_fa24_6_or0 = s_csamul_cla32_fa24_6_and0 | s_csamul_cla32_fa24_6_and1;
  assign s_csamul_cla32_and25_6 = a[25] & b[6];
  assign s_csamul_cla32_fa25_6_xor0 = s_csamul_cla32_and25_6 ^ s_csamul_cla32_fa26_5_xor1;
  assign s_csamul_cla32_fa25_6_and0 = s_csamul_cla32_and25_6 & s_csamul_cla32_fa26_5_xor1;
  assign s_csamul_cla32_fa25_6_xor1 = s_csamul_cla32_fa25_6_xor0 ^ s_csamul_cla32_fa25_5_or0;
  assign s_csamul_cla32_fa25_6_and1 = s_csamul_cla32_fa25_6_xor0 & s_csamul_cla32_fa25_5_or0;
  assign s_csamul_cla32_fa25_6_or0 = s_csamul_cla32_fa25_6_and0 | s_csamul_cla32_fa25_6_and1;
  assign s_csamul_cla32_and26_6 = a[26] & b[6];
  assign s_csamul_cla32_fa26_6_xor0 = s_csamul_cla32_and26_6 ^ s_csamul_cla32_fa27_5_xor1;
  assign s_csamul_cla32_fa26_6_and0 = s_csamul_cla32_and26_6 & s_csamul_cla32_fa27_5_xor1;
  assign s_csamul_cla32_fa26_6_xor1 = s_csamul_cla32_fa26_6_xor0 ^ s_csamul_cla32_fa26_5_or0;
  assign s_csamul_cla32_fa26_6_and1 = s_csamul_cla32_fa26_6_xor0 & s_csamul_cla32_fa26_5_or0;
  assign s_csamul_cla32_fa26_6_or0 = s_csamul_cla32_fa26_6_and0 | s_csamul_cla32_fa26_6_and1;
  assign s_csamul_cla32_and27_6 = a[27] & b[6];
  assign s_csamul_cla32_fa27_6_xor0 = s_csamul_cla32_and27_6 ^ s_csamul_cla32_fa28_5_xor1;
  assign s_csamul_cla32_fa27_6_and0 = s_csamul_cla32_and27_6 & s_csamul_cla32_fa28_5_xor1;
  assign s_csamul_cla32_fa27_6_xor1 = s_csamul_cla32_fa27_6_xor0 ^ s_csamul_cla32_fa27_5_or0;
  assign s_csamul_cla32_fa27_6_and1 = s_csamul_cla32_fa27_6_xor0 & s_csamul_cla32_fa27_5_or0;
  assign s_csamul_cla32_fa27_6_or0 = s_csamul_cla32_fa27_6_and0 | s_csamul_cla32_fa27_6_and1;
  assign s_csamul_cla32_and28_6 = a[28] & b[6];
  assign s_csamul_cla32_fa28_6_xor0 = s_csamul_cla32_and28_6 ^ s_csamul_cla32_fa29_5_xor1;
  assign s_csamul_cla32_fa28_6_and0 = s_csamul_cla32_and28_6 & s_csamul_cla32_fa29_5_xor1;
  assign s_csamul_cla32_fa28_6_xor1 = s_csamul_cla32_fa28_6_xor0 ^ s_csamul_cla32_fa28_5_or0;
  assign s_csamul_cla32_fa28_6_and1 = s_csamul_cla32_fa28_6_xor0 & s_csamul_cla32_fa28_5_or0;
  assign s_csamul_cla32_fa28_6_or0 = s_csamul_cla32_fa28_6_and0 | s_csamul_cla32_fa28_6_and1;
  assign s_csamul_cla32_and29_6 = a[29] & b[6];
  assign s_csamul_cla32_fa29_6_xor0 = s_csamul_cla32_and29_6 ^ s_csamul_cla32_fa30_5_xor1;
  assign s_csamul_cla32_fa29_6_and0 = s_csamul_cla32_and29_6 & s_csamul_cla32_fa30_5_xor1;
  assign s_csamul_cla32_fa29_6_xor1 = s_csamul_cla32_fa29_6_xor0 ^ s_csamul_cla32_fa29_5_or0;
  assign s_csamul_cla32_fa29_6_and1 = s_csamul_cla32_fa29_6_xor0 & s_csamul_cla32_fa29_5_or0;
  assign s_csamul_cla32_fa29_6_or0 = s_csamul_cla32_fa29_6_and0 | s_csamul_cla32_fa29_6_and1;
  assign s_csamul_cla32_and30_6 = a[30] & b[6];
  assign s_csamul_cla32_fa30_6_xor0 = s_csamul_cla32_and30_6 ^ s_csamul_cla32_ha31_5_xor0;
  assign s_csamul_cla32_fa30_6_and0 = s_csamul_cla32_and30_6 & s_csamul_cla32_ha31_5_xor0;
  assign s_csamul_cla32_fa30_6_xor1 = s_csamul_cla32_fa30_6_xor0 ^ s_csamul_cla32_fa30_5_or0;
  assign s_csamul_cla32_fa30_6_and1 = s_csamul_cla32_fa30_6_xor0 & s_csamul_cla32_fa30_5_or0;
  assign s_csamul_cla32_fa30_6_or0 = s_csamul_cla32_fa30_6_and0 | s_csamul_cla32_fa30_6_and1;
  assign s_csamul_cla32_nand31_6 = ~(a[31] & b[6]);
  assign s_csamul_cla32_ha31_6_xor0 = s_csamul_cla32_nand31_6 ^ s_csamul_cla32_ha31_5_and0;
  assign s_csamul_cla32_ha31_6_and0 = s_csamul_cla32_nand31_6 & s_csamul_cla32_ha31_5_and0;
  assign s_csamul_cla32_and0_7 = a[0] & b[7];
  assign s_csamul_cla32_fa0_7_xor0 = s_csamul_cla32_and0_7 ^ s_csamul_cla32_fa1_6_xor1;
  assign s_csamul_cla32_fa0_7_and0 = s_csamul_cla32_and0_7 & s_csamul_cla32_fa1_6_xor1;
  assign s_csamul_cla32_fa0_7_xor1 = s_csamul_cla32_fa0_7_xor0 ^ s_csamul_cla32_fa0_6_or0;
  assign s_csamul_cla32_fa0_7_and1 = s_csamul_cla32_fa0_7_xor0 & s_csamul_cla32_fa0_6_or0;
  assign s_csamul_cla32_fa0_7_or0 = s_csamul_cla32_fa0_7_and0 | s_csamul_cla32_fa0_7_and1;
  assign s_csamul_cla32_and1_7 = a[1] & b[7];
  assign s_csamul_cla32_fa1_7_xor0 = s_csamul_cla32_and1_7 ^ s_csamul_cla32_fa2_6_xor1;
  assign s_csamul_cla32_fa1_7_and0 = s_csamul_cla32_and1_7 & s_csamul_cla32_fa2_6_xor1;
  assign s_csamul_cla32_fa1_7_xor1 = s_csamul_cla32_fa1_7_xor0 ^ s_csamul_cla32_fa1_6_or0;
  assign s_csamul_cla32_fa1_7_and1 = s_csamul_cla32_fa1_7_xor0 & s_csamul_cla32_fa1_6_or0;
  assign s_csamul_cla32_fa1_7_or0 = s_csamul_cla32_fa1_7_and0 | s_csamul_cla32_fa1_7_and1;
  assign s_csamul_cla32_and2_7 = a[2] & b[7];
  assign s_csamul_cla32_fa2_7_xor0 = s_csamul_cla32_and2_7 ^ s_csamul_cla32_fa3_6_xor1;
  assign s_csamul_cla32_fa2_7_and0 = s_csamul_cla32_and2_7 & s_csamul_cla32_fa3_6_xor1;
  assign s_csamul_cla32_fa2_7_xor1 = s_csamul_cla32_fa2_7_xor0 ^ s_csamul_cla32_fa2_6_or0;
  assign s_csamul_cla32_fa2_7_and1 = s_csamul_cla32_fa2_7_xor0 & s_csamul_cla32_fa2_6_or0;
  assign s_csamul_cla32_fa2_7_or0 = s_csamul_cla32_fa2_7_and0 | s_csamul_cla32_fa2_7_and1;
  assign s_csamul_cla32_and3_7 = a[3] & b[7];
  assign s_csamul_cla32_fa3_7_xor0 = s_csamul_cla32_and3_7 ^ s_csamul_cla32_fa4_6_xor1;
  assign s_csamul_cla32_fa3_7_and0 = s_csamul_cla32_and3_7 & s_csamul_cla32_fa4_6_xor1;
  assign s_csamul_cla32_fa3_7_xor1 = s_csamul_cla32_fa3_7_xor0 ^ s_csamul_cla32_fa3_6_or0;
  assign s_csamul_cla32_fa3_7_and1 = s_csamul_cla32_fa3_7_xor0 & s_csamul_cla32_fa3_6_or0;
  assign s_csamul_cla32_fa3_7_or0 = s_csamul_cla32_fa3_7_and0 | s_csamul_cla32_fa3_7_and1;
  assign s_csamul_cla32_and4_7 = a[4] & b[7];
  assign s_csamul_cla32_fa4_7_xor0 = s_csamul_cla32_and4_7 ^ s_csamul_cla32_fa5_6_xor1;
  assign s_csamul_cla32_fa4_7_and0 = s_csamul_cla32_and4_7 & s_csamul_cla32_fa5_6_xor1;
  assign s_csamul_cla32_fa4_7_xor1 = s_csamul_cla32_fa4_7_xor0 ^ s_csamul_cla32_fa4_6_or0;
  assign s_csamul_cla32_fa4_7_and1 = s_csamul_cla32_fa4_7_xor0 & s_csamul_cla32_fa4_6_or0;
  assign s_csamul_cla32_fa4_7_or0 = s_csamul_cla32_fa4_7_and0 | s_csamul_cla32_fa4_7_and1;
  assign s_csamul_cla32_and5_7 = a[5] & b[7];
  assign s_csamul_cla32_fa5_7_xor0 = s_csamul_cla32_and5_7 ^ s_csamul_cla32_fa6_6_xor1;
  assign s_csamul_cla32_fa5_7_and0 = s_csamul_cla32_and5_7 & s_csamul_cla32_fa6_6_xor1;
  assign s_csamul_cla32_fa5_7_xor1 = s_csamul_cla32_fa5_7_xor0 ^ s_csamul_cla32_fa5_6_or0;
  assign s_csamul_cla32_fa5_7_and1 = s_csamul_cla32_fa5_7_xor0 & s_csamul_cla32_fa5_6_or0;
  assign s_csamul_cla32_fa5_7_or0 = s_csamul_cla32_fa5_7_and0 | s_csamul_cla32_fa5_7_and1;
  assign s_csamul_cla32_and6_7 = a[6] & b[7];
  assign s_csamul_cla32_fa6_7_xor0 = s_csamul_cla32_and6_7 ^ s_csamul_cla32_fa7_6_xor1;
  assign s_csamul_cla32_fa6_7_and0 = s_csamul_cla32_and6_7 & s_csamul_cla32_fa7_6_xor1;
  assign s_csamul_cla32_fa6_7_xor1 = s_csamul_cla32_fa6_7_xor0 ^ s_csamul_cla32_fa6_6_or0;
  assign s_csamul_cla32_fa6_7_and1 = s_csamul_cla32_fa6_7_xor0 & s_csamul_cla32_fa6_6_or0;
  assign s_csamul_cla32_fa6_7_or0 = s_csamul_cla32_fa6_7_and0 | s_csamul_cla32_fa6_7_and1;
  assign s_csamul_cla32_and7_7 = a[7] & b[7];
  assign s_csamul_cla32_fa7_7_xor0 = s_csamul_cla32_and7_7 ^ s_csamul_cla32_fa8_6_xor1;
  assign s_csamul_cla32_fa7_7_and0 = s_csamul_cla32_and7_7 & s_csamul_cla32_fa8_6_xor1;
  assign s_csamul_cla32_fa7_7_xor1 = s_csamul_cla32_fa7_7_xor0 ^ s_csamul_cla32_fa7_6_or0;
  assign s_csamul_cla32_fa7_7_and1 = s_csamul_cla32_fa7_7_xor0 & s_csamul_cla32_fa7_6_or0;
  assign s_csamul_cla32_fa7_7_or0 = s_csamul_cla32_fa7_7_and0 | s_csamul_cla32_fa7_7_and1;
  assign s_csamul_cla32_and8_7 = a[8] & b[7];
  assign s_csamul_cla32_fa8_7_xor0 = s_csamul_cla32_and8_7 ^ s_csamul_cla32_fa9_6_xor1;
  assign s_csamul_cla32_fa8_7_and0 = s_csamul_cla32_and8_7 & s_csamul_cla32_fa9_6_xor1;
  assign s_csamul_cla32_fa8_7_xor1 = s_csamul_cla32_fa8_7_xor0 ^ s_csamul_cla32_fa8_6_or0;
  assign s_csamul_cla32_fa8_7_and1 = s_csamul_cla32_fa8_7_xor0 & s_csamul_cla32_fa8_6_or0;
  assign s_csamul_cla32_fa8_7_or0 = s_csamul_cla32_fa8_7_and0 | s_csamul_cla32_fa8_7_and1;
  assign s_csamul_cla32_and9_7 = a[9] & b[7];
  assign s_csamul_cla32_fa9_7_xor0 = s_csamul_cla32_and9_7 ^ s_csamul_cla32_fa10_6_xor1;
  assign s_csamul_cla32_fa9_7_and0 = s_csamul_cla32_and9_7 & s_csamul_cla32_fa10_6_xor1;
  assign s_csamul_cla32_fa9_7_xor1 = s_csamul_cla32_fa9_7_xor0 ^ s_csamul_cla32_fa9_6_or0;
  assign s_csamul_cla32_fa9_7_and1 = s_csamul_cla32_fa9_7_xor0 & s_csamul_cla32_fa9_6_or0;
  assign s_csamul_cla32_fa9_7_or0 = s_csamul_cla32_fa9_7_and0 | s_csamul_cla32_fa9_7_and1;
  assign s_csamul_cla32_and10_7 = a[10] & b[7];
  assign s_csamul_cla32_fa10_7_xor0 = s_csamul_cla32_and10_7 ^ s_csamul_cla32_fa11_6_xor1;
  assign s_csamul_cla32_fa10_7_and0 = s_csamul_cla32_and10_7 & s_csamul_cla32_fa11_6_xor1;
  assign s_csamul_cla32_fa10_7_xor1 = s_csamul_cla32_fa10_7_xor0 ^ s_csamul_cla32_fa10_6_or0;
  assign s_csamul_cla32_fa10_7_and1 = s_csamul_cla32_fa10_7_xor0 & s_csamul_cla32_fa10_6_or0;
  assign s_csamul_cla32_fa10_7_or0 = s_csamul_cla32_fa10_7_and0 | s_csamul_cla32_fa10_7_and1;
  assign s_csamul_cla32_and11_7 = a[11] & b[7];
  assign s_csamul_cla32_fa11_7_xor0 = s_csamul_cla32_and11_7 ^ s_csamul_cla32_fa12_6_xor1;
  assign s_csamul_cla32_fa11_7_and0 = s_csamul_cla32_and11_7 & s_csamul_cla32_fa12_6_xor1;
  assign s_csamul_cla32_fa11_7_xor1 = s_csamul_cla32_fa11_7_xor0 ^ s_csamul_cla32_fa11_6_or0;
  assign s_csamul_cla32_fa11_7_and1 = s_csamul_cla32_fa11_7_xor0 & s_csamul_cla32_fa11_6_or0;
  assign s_csamul_cla32_fa11_7_or0 = s_csamul_cla32_fa11_7_and0 | s_csamul_cla32_fa11_7_and1;
  assign s_csamul_cla32_and12_7 = a[12] & b[7];
  assign s_csamul_cla32_fa12_7_xor0 = s_csamul_cla32_and12_7 ^ s_csamul_cla32_fa13_6_xor1;
  assign s_csamul_cla32_fa12_7_and0 = s_csamul_cla32_and12_7 & s_csamul_cla32_fa13_6_xor1;
  assign s_csamul_cla32_fa12_7_xor1 = s_csamul_cla32_fa12_7_xor0 ^ s_csamul_cla32_fa12_6_or0;
  assign s_csamul_cla32_fa12_7_and1 = s_csamul_cla32_fa12_7_xor0 & s_csamul_cla32_fa12_6_or0;
  assign s_csamul_cla32_fa12_7_or0 = s_csamul_cla32_fa12_7_and0 | s_csamul_cla32_fa12_7_and1;
  assign s_csamul_cla32_and13_7 = a[13] & b[7];
  assign s_csamul_cla32_fa13_7_xor0 = s_csamul_cla32_and13_7 ^ s_csamul_cla32_fa14_6_xor1;
  assign s_csamul_cla32_fa13_7_and0 = s_csamul_cla32_and13_7 & s_csamul_cla32_fa14_6_xor1;
  assign s_csamul_cla32_fa13_7_xor1 = s_csamul_cla32_fa13_7_xor0 ^ s_csamul_cla32_fa13_6_or0;
  assign s_csamul_cla32_fa13_7_and1 = s_csamul_cla32_fa13_7_xor0 & s_csamul_cla32_fa13_6_or0;
  assign s_csamul_cla32_fa13_7_or0 = s_csamul_cla32_fa13_7_and0 | s_csamul_cla32_fa13_7_and1;
  assign s_csamul_cla32_and14_7 = a[14] & b[7];
  assign s_csamul_cla32_fa14_7_xor0 = s_csamul_cla32_and14_7 ^ s_csamul_cla32_fa15_6_xor1;
  assign s_csamul_cla32_fa14_7_and0 = s_csamul_cla32_and14_7 & s_csamul_cla32_fa15_6_xor1;
  assign s_csamul_cla32_fa14_7_xor1 = s_csamul_cla32_fa14_7_xor0 ^ s_csamul_cla32_fa14_6_or0;
  assign s_csamul_cla32_fa14_7_and1 = s_csamul_cla32_fa14_7_xor0 & s_csamul_cla32_fa14_6_or0;
  assign s_csamul_cla32_fa14_7_or0 = s_csamul_cla32_fa14_7_and0 | s_csamul_cla32_fa14_7_and1;
  assign s_csamul_cla32_and15_7 = a[15] & b[7];
  assign s_csamul_cla32_fa15_7_xor0 = s_csamul_cla32_and15_7 ^ s_csamul_cla32_fa16_6_xor1;
  assign s_csamul_cla32_fa15_7_and0 = s_csamul_cla32_and15_7 & s_csamul_cla32_fa16_6_xor1;
  assign s_csamul_cla32_fa15_7_xor1 = s_csamul_cla32_fa15_7_xor0 ^ s_csamul_cla32_fa15_6_or0;
  assign s_csamul_cla32_fa15_7_and1 = s_csamul_cla32_fa15_7_xor0 & s_csamul_cla32_fa15_6_or0;
  assign s_csamul_cla32_fa15_7_or0 = s_csamul_cla32_fa15_7_and0 | s_csamul_cla32_fa15_7_and1;
  assign s_csamul_cla32_and16_7 = a[16] & b[7];
  assign s_csamul_cla32_fa16_7_xor0 = s_csamul_cla32_and16_7 ^ s_csamul_cla32_fa17_6_xor1;
  assign s_csamul_cla32_fa16_7_and0 = s_csamul_cla32_and16_7 & s_csamul_cla32_fa17_6_xor1;
  assign s_csamul_cla32_fa16_7_xor1 = s_csamul_cla32_fa16_7_xor0 ^ s_csamul_cla32_fa16_6_or0;
  assign s_csamul_cla32_fa16_7_and1 = s_csamul_cla32_fa16_7_xor0 & s_csamul_cla32_fa16_6_or0;
  assign s_csamul_cla32_fa16_7_or0 = s_csamul_cla32_fa16_7_and0 | s_csamul_cla32_fa16_7_and1;
  assign s_csamul_cla32_and17_7 = a[17] & b[7];
  assign s_csamul_cla32_fa17_7_xor0 = s_csamul_cla32_and17_7 ^ s_csamul_cla32_fa18_6_xor1;
  assign s_csamul_cla32_fa17_7_and0 = s_csamul_cla32_and17_7 & s_csamul_cla32_fa18_6_xor1;
  assign s_csamul_cla32_fa17_7_xor1 = s_csamul_cla32_fa17_7_xor0 ^ s_csamul_cla32_fa17_6_or0;
  assign s_csamul_cla32_fa17_7_and1 = s_csamul_cla32_fa17_7_xor0 & s_csamul_cla32_fa17_6_or0;
  assign s_csamul_cla32_fa17_7_or0 = s_csamul_cla32_fa17_7_and0 | s_csamul_cla32_fa17_7_and1;
  assign s_csamul_cla32_and18_7 = a[18] & b[7];
  assign s_csamul_cla32_fa18_7_xor0 = s_csamul_cla32_and18_7 ^ s_csamul_cla32_fa19_6_xor1;
  assign s_csamul_cla32_fa18_7_and0 = s_csamul_cla32_and18_7 & s_csamul_cla32_fa19_6_xor1;
  assign s_csamul_cla32_fa18_7_xor1 = s_csamul_cla32_fa18_7_xor0 ^ s_csamul_cla32_fa18_6_or0;
  assign s_csamul_cla32_fa18_7_and1 = s_csamul_cla32_fa18_7_xor0 & s_csamul_cla32_fa18_6_or0;
  assign s_csamul_cla32_fa18_7_or0 = s_csamul_cla32_fa18_7_and0 | s_csamul_cla32_fa18_7_and1;
  assign s_csamul_cla32_and19_7 = a[19] & b[7];
  assign s_csamul_cla32_fa19_7_xor0 = s_csamul_cla32_and19_7 ^ s_csamul_cla32_fa20_6_xor1;
  assign s_csamul_cla32_fa19_7_and0 = s_csamul_cla32_and19_7 & s_csamul_cla32_fa20_6_xor1;
  assign s_csamul_cla32_fa19_7_xor1 = s_csamul_cla32_fa19_7_xor0 ^ s_csamul_cla32_fa19_6_or0;
  assign s_csamul_cla32_fa19_7_and1 = s_csamul_cla32_fa19_7_xor0 & s_csamul_cla32_fa19_6_or0;
  assign s_csamul_cla32_fa19_7_or0 = s_csamul_cla32_fa19_7_and0 | s_csamul_cla32_fa19_7_and1;
  assign s_csamul_cla32_and20_7 = a[20] & b[7];
  assign s_csamul_cla32_fa20_7_xor0 = s_csamul_cla32_and20_7 ^ s_csamul_cla32_fa21_6_xor1;
  assign s_csamul_cla32_fa20_7_and0 = s_csamul_cla32_and20_7 & s_csamul_cla32_fa21_6_xor1;
  assign s_csamul_cla32_fa20_7_xor1 = s_csamul_cla32_fa20_7_xor0 ^ s_csamul_cla32_fa20_6_or0;
  assign s_csamul_cla32_fa20_7_and1 = s_csamul_cla32_fa20_7_xor0 & s_csamul_cla32_fa20_6_or0;
  assign s_csamul_cla32_fa20_7_or0 = s_csamul_cla32_fa20_7_and0 | s_csamul_cla32_fa20_7_and1;
  assign s_csamul_cla32_and21_7 = a[21] & b[7];
  assign s_csamul_cla32_fa21_7_xor0 = s_csamul_cla32_and21_7 ^ s_csamul_cla32_fa22_6_xor1;
  assign s_csamul_cla32_fa21_7_and0 = s_csamul_cla32_and21_7 & s_csamul_cla32_fa22_6_xor1;
  assign s_csamul_cla32_fa21_7_xor1 = s_csamul_cla32_fa21_7_xor0 ^ s_csamul_cla32_fa21_6_or0;
  assign s_csamul_cla32_fa21_7_and1 = s_csamul_cla32_fa21_7_xor0 & s_csamul_cla32_fa21_6_or0;
  assign s_csamul_cla32_fa21_7_or0 = s_csamul_cla32_fa21_7_and0 | s_csamul_cla32_fa21_7_and1;
  assign s_csamul_cla32_and22_7 = a[22] & b[7];
  assign s_csamul_cla32_fa22_7_xor0 = s_csamul_cla32_and22_7 ^ s_csamul_cla32_fa23_6_xor1;
  assign s_csamul_cla32_fa22_7_and0 = s_csamul_cla32_and22_7 & s_csamul_cla32_fa23_6_xor1;
  assign s_csamul_cla32_fa22_7_xor1 = s_csamul_cla32_fa22_7_xor0 ^ s_csamul_cla32_fa22_6_or0;
  assign s_csamul_cla32_fa22_7_and1 = s_csamul_cla32_fa22_7_xor0 & s_csamul_cla32_fa22_6_or0;
  assign s_csamul_cla32_fa22_7_or0 = s_csamul_cla32_fa22_7_and0 | s_csamul_cla32_fa22_7_and1;
  assign s_csamul_cla32_and23_7 = a[23] & b[7];
  assign s_csamul_cla32_fa23_7_xor0 = s_csamul_cla32_and23_7 ^ s_csamul_cla32_fa24_6_xor1;
  assign s_csamul_cla32_fa23_7_and0 = s_csamul_cla32_and23_7 & s_csamul_cla32_fa24_6_xor1;
  assign s_csamul_cla32_fa23_7_xor1 = s_csamul_cla32_fa23_7_xor0 ^ s_csamul_cla32_fa23_6_or0;
  assign s_csamul_cla32_fa23_7_and1 = s_csamul_cla32_fa23_7_xor0 & s_csamul_cla32_fa23_6_or0;
  assign s_csamul_cla32_fa23_7_or0 = s_csamul_cla32_fa23_7_and0 | s_csamul_cla32_fa23_7_and1;
  assign s_csamul_cla32_and24_7 = a[24] & b[7];
  assign s_csamul_cla32_fa24_7_xor0 = s_csamul_cla32_and24_7 ^ s_csamul_cla32_fa25_6_xor1;
  assign s_csamul_cla32_fa24_7_and0 = s_csamul_cla32_and24_7 & s_csamul_cla32_fa25_6_xor1;
  assign s_csamul_cla32_fa24_7_xor1 = s_csamul_cla32_fa24_7_xor0 ^ s_csamul_cla32_fa24_6_or0;
  assign s_csamul_cla32_fa24_7_and1 = s_csamul_cla32_fa24_7_xor0 & s_csamul_cla32_fa24_6_or0;
  assign s_csamul_cla32_fa24_7_or0 = s_csamul_cla32_fa24_7_and0 | s_csamul_cla32_fa24_7_and1;
  assign s_csamul_cla32_and25_7 = a[25] & b[7];
  assign s_csamul_cla32_fa25_7_xor0 = s_csamul_cla32_and25_7 ^ s_csamul_cla32_fa26_6_xor1;
  assign s_csamul_cla32_fa25_7_and0 = s_csamul_cla32_and25_7 & s_csamul_cla32_fa26_6_xor1;
  assign s_csamul_cla32_fa25_7_xor1 = s_csamul_cla32_fa25_7_xor0 ^ s_csamul_cla32_fa25_6_or0;
  assign s_csamul_cla32_fa25_7_and1 = s_csamul_cla32_fa25_7_xor0 & s_csamul_cla32_fa25_6_or0;
  assign s_csamul_cla32_fa25_7_or0 = s_csamul_cla32_fa25_7_and0 | s_csamul_cla32_fa25_7_and1;
  assign s_csamul_cla32_and26_7 = a[26] & b[7];
  assign s_csamul_cla32_fa26_7_xor0 = s_csamul_cla32_and26_7 ^ s_csamul_cla32_fa27_6_xor1;
  assign s_csamul_cla32_fa26_7_and0 = s_csamul_cla32_and26_7 & s_csamul_cla32_fa27_6_xor1;
  assign s_csamul_cla32_fa26_7_xor1 = s_csamul_cla32_fa26_7_xor0 ^ s_csamul_cla32_fa26_6_or0;
  assign s_csamul_cla32_fa26_7_and1 = s_csamul_cla32_fa26_7_xor0 & s_csamul_cla32_fa26_6_or0;
  assign s_csamul_cla32_fa26_7_or0 = s_csamul_cla32_fa26_7_and0 | s_csamul_cla32_fa26_7_and1;
  assign s_csamul_cla32_and27_7 = a[27] & b[7];
  assign s_csamul_cla32_fa27_7_xor0 = s_csamul_cla32_and27_7 ^ s_csamul_cla32_fa28_6_xor1;
  assign s_csamul_cla32_fa27_7_and0 = s_csamul_cla32_and27_7 & s_csamul_cla32_fa28_6_xor1;
  assign s_csamul_cla32_fa27_7_xor1 = s_csamul_cla32_fa27_7_xor0 ^ s_csamul_cla32_fa27_6_or0;
  assign s_csamul_cla32_fa27_7_and1 = s_csamul_cla32_fa27_7_xor0 & s_csamul_cla32_fa27_6_or0;
  assign s_csamul_cla32_fa27_7_or0 = s_csamul_cla32_fa27_7_and0 | s_csamul_cla32_fa27_7_and1;
  assign s_csamul_cla32_and28_7 = a[28] & b[7];
  assign s_csamul_cla32_fa28_7_xor0 = s_csamul_cla32_and28_7 ^ s_csamul_cla32_fa29_6_xor1;
  assign s_csamul_cla32_fa28_7_and0 = s_csamul_cla32_and28_7 & s_csamul_cla32_fa29_6_xor1;
  assign s_csamul_cla32_fa28_7_xor1 = s_csamul_cla32_fa28_7_xor0 ^ s_csamul_cla32_fa28_6_or0;
  assign s_csamul_cla32_fa28_7_and1 = s_csamul_cla32_fa28_7_xor0 & s_csamul_cla32_fa28_6_or0;
  assign s_csamul_cla32_fa28_7_or0 = s_csamul_cla32_fa28_7_and0 | s_csamul_cla32_fa28_7_and1;
  assign s_csamul_cla32_and29_7 = a[29] & b[7];
  assign s_csamul_cla32_fa29_7_xor0 = s_csamul_cla32_and29_7 ^ s_csamul_cla32_fa30_6_xor1;
  assign s_csamul_cla32_fa29_7_and0 = s_csamul_cla32_and29_7 & s_csamul_cla32_fa30_6_xor1;
  assign s_csamul_cla32_fa29_7_xor1 = s_csamul_cla32_fa29_7_xor0 ^ s_csamul_cla32_fa29_6_or0;
  assign s_csamul_cla32_fa29_7_and1 = s_csamul_cla32_fa29_7_xor0 & s_csamul_cla32_fa29_6_or0;
  assign s_csamul_cla32_fa29_7_or0 = s_csamul_cla32_fa29_7_and0 | s_csamul_cla32_fa29_7_and1;
  assign s_csamul_cla32_and30_7 = a[30] & b[7];
  assign s_csamul_cla32_fa30_7_xor0 = s_csamul_cla32_and30_7 ^ s_csamul_cla32_ha31_6_xor0;
  assign s_csamul_cla32_fa30_7_and0 = s_csamul_cla32_and30_7 & s_csamul_cla32_ha31_6_xor0;
  assign s_csamul_cla32_fa30_7_xor1 = s_csamul_cla32_fa30_7_xor0 ^ s_csamul_cla32_fa30_6_or0;
  assign s_csamul_cla32_fa30_7_and1 = s_csamul_cla32_fa30_7_xor0 & s_csamul_cla32_fa30_6_or0;
  assign s_csamul_cla32_fa30_7_or0 = s_csamul_cla32_fa30_7_and0 | s_csamul_cla32_fa30_7_and1;
  assign s_csamul_cla32_nand31_7 = ~(a[31] & b[7]);
  assign s_csamul_cla32_ha31_7_xor0 = s_csamul_cla32_nand31_7 ^ s_csamul_cla32_ha31_6_and0;
  assign s_csamul_cla32_ha31_7_and0 = s_csamul_cla32_nand31_7 & s_csamul_cla32_ha31_6_and0;
  assign s_csamul_cla32_and0_8 = a[0] & b[8];
  assign s_csamul_cla32_fa0_8_xor0 = s_csamul_cla32_and0_8 ^ s_csamul_cla32_fa1_7_xor1;
  assign s_csamul_cla32_fa0_8_and0 = s_csamul_cla32_and0_8 & s_csamul_cla32_fa1_7_xor1;
  assign s_csamul_cla32_fa0_8_xor1 = s_csamul_cla32_fa0_8_xor0 ^ s_csamul_cla32_fa0_7_or0;
  assign s_csamul_cla32_fa0_8_and1 = s_csamul_cla32_fa0_8_xor0 & s_csamul_cla32_fa0_7_or0;
  assign s_csamul_cla32_fa0_8_or0 = s_csamul_cla32_fa0_8_and0 | s_csamul_cla32_fa0_8_and1;
  assign s_csamul_cla32_and1_8 = a[1] & b[8];
  assign s_csamul_cla32_fa1_8_xor0 = s_csamul_cla32_and1_8 ^ s_csamul_cla32_fa2_7_xor1;
  assign s_csamul_cla32_fa1_8_and0 = s_csamul_cla32_and1_8 & s_csamul_cla32_fa2_7_xor1;
  assign s_csamul_cla32_fa1_8_xor1 = s_csamul_cla32_fa1_8_xor0 ^ s_csamul_cla32_fa1_7_or0;
  assign s_csamul_cla32_fa1_8_and1 = s_csamul_cla32_fa1_8_xor0 & s_csamul_cla32_fa1_7_or0;
  assign s_csamul_cla32_fa1_8_or0 = s_csamul_cla32_fa1_8_and0 | s_csamul_cla32_fa1_8_and1;
  assign s_csamul_cla32_and2_8 = a[2] & b[8];
  assign s_csamul_cla32_fa2_8_xor0 = s_csamul_cla32_and2_8 ^ s_csamul_cla32_fa3_7_xor1;
  assign s_csamul_cla32_fa2_8_and0 = s_csamul_cla32_and2_8 & s_csamul_cla32_fa3_7_xor1;
  assign s_csamul_cla32_fa2_8_xor1 = s_csamul_cla32_fa2_8_xor0 ^ s_csamul_cla32_fa2_7_or0;
  assign s_csamul_cla32_fa2_8_and1 = s_csamul_cla32_fa2_8_xor0 & s_csamul_cla32_fa2_7_or0;
  assign s_csamul_cla32_fa2_8_or0 = s_csamul_cla32_fa2_8_and0 | s_csamul_cla32_fa2_8_and1;
  assign s_csamul_cla32_and3_8 = a[3] & b[8];
  assign s_csamul_cla32_fa3_8_xor0 = s_csamul_cla32_and3_8 ^ s_csamul_cla32_fa4_7_xor1;
  assign s_csamul_cla32_fa3_8_and0 = s_csamul_cla32_and3_8 & s_csamul_cla32_fa4_7_xor1;
  assign s_csamul_cla32_fa3_8_xor1 = s_csamul_cla32_fa3_8_xor0 ^ s_csamul_cla32_fa3_7_or0;
  assign s_csamul_cla32_fa3_8_and1 = s_csamul_cla32_fa3_8_xor0 & s_csamul_cla32_fa3_7_or0;
  assign s_csamul_cla32_fa3_8_or0 = s_csamul_cla32_fa3_8_and0 | s_csamul_cla32_fa3_8_and1;
  assign s_csamul_cla32_and4_8 = a[4] & b[8];
  assign s_csamul_cla32_fa4_8_xor0 = s_csamul_cla32_and4_8 ^ s_csamul_cla32_fa5_7_xor1;
  assign s_csamul_cla32_fa4_8_and0 = s_csamul_cla32_and4_8 & s_csamul_cla32_fa5_7_xor1;
  assign s_csamul_cla32_fa4_8_xor1 = s_csamul_cla32_fa4_8_xor0 ^ s_csamul_cla32_fa4_7_or0;
  assign s_csamul_cla32_fa4_8_and1 = s_csamul_cla32_fa4_8_xor0 & s_csamul_cla32_fa4_7_or0;
  assign s_csamul_cla32_fa4_8_or0 = s_csamul_cla32_fa4_8_and0 | s_csamul_cla32_fa4_8_and1;
  assign s_csamul_cla32_and5_8 = a[5] & b[8];
  assign s_csamul_cla32_fa5_8_xor0 = s_csamul_cla32_and5_8 ^ s_csamul_cla32_fa6_7_xor1;
  assign s_csamul_cla32_fa5_8_and0 = s_csamul_cla32_and5_8 & s_csamul_cla32_fa6_7_xor1;
  assign s_csamul_cla32_fa5_8_xor1 = s_csamul_cla32_fa5_8_xor0 ^ s_csamul_cla32_fa5_7_or0;
  assign s_csamul_cla32_fa5_8_and1 = s_csamul_cla32_fa5_8_xor0 & s_csamul_cla32_fa5_7_or0;
  assign s_csamul_cla32_fa5_8_or0 = s_csamul_cla32_fa5_8_and0 | s_csamul_cla32_fa5_8_and1;
  assign s_csamul_cla32_and6_8 = a[6] & b[8];
  assign s_csamul_cla32_fa6_8_xor0 = s_csamul_cla32_and6_8 ^ s_csamul_cla32_fa7_7_xor1;
  assign s_csamul_cla32_fa6_8_and0 = s_csamul_cla32_and6_8 & s_csamul_cla32_fa7_7_xor1;
  assign s_csamul_cla32_fa6_8_xor1 = s_csamul_cla32_fa6_8_xor0 ^ s_csamul_cla32_fa6_7_or0;
  assign s_csamul_cla32_fa6_8_and1 = s_csamul_cla32_fa6_8_xor0 & s_csamul_cla32_fa6_7_or0;
  assign s_csamul_cla32_fa6_8_or0 = s_csamul_cla32_fa6_8_and0 | s_csamul_cla32_fa6_8_and1;
  assign s_csamul_cla32_and7_8 = a[7] & b[8];
  assign s_csamul_cla32_fa7_8_xor0 = s_csamul_cla32_and7_8 ^ s_csamul_cla32_fa8_7_xor1;
  assign s_csamul_cla32_fa7_8_and0 = s_csamul_cla32_and7_8 & s_csamul_cla32_fa8_7_xor1;
  assign s_csamul_cla32_fa7_8_xor1 = s_csamul_cla32_fa7_8_xor0 ^ s_csamul_cla32_fa7_7_or0;
  assign s_csamul_cla32_fa7_8_and1 = s_csamul_cla32_fa7_8_xor0 & s_csamul_cla32_fa7_7_or0;
  assign s_csamul_cla32_fa7_8_or0 = s_csamul_cla32_fa7_8_and0 | s_csamul_cla32_fa7_8_and1;
  assign s_csamul_cla32_and8_8 = a[8] & b[8];
  assign s_csamul_cla32_fa8_8_xor0 = s_csamul_cla32_and8_8 ^ s_csamul_cla32_fa9_7_xor1;
  assign s_csamul_cla32_fa8_8_and0 = s_csamul_cla32_and8_8 & s_csamul_cla32_fa9_7_xor1;
  assign s_csamul_cla32_fa8_8_xor1 = s_csamul_cla32_fa8_8_xor0 ^ s_csamul_cla32_fa8_7_or0;
  assign s_csamul_cla32_fa8_8_and1 = s_csamul_cla32_fa8_8_xor0 & s_csamul_cla32_fa8_7_or0;
  assign s_csamul_cla32_fa8_8_or0 = s_csamul_cla32_fa8_8_and0 | s_csamul_cla32_fa8_8_and1;
  assign s_csamul_cla32_and9_8 = a[9] & b[8];
  assign s_csamul_cla32_fa9_8_xor0 = s_csamul_cla32_and9_8 ^ s_csamul_cla32_fa10_7_xor1;
  assign s_csamul_cla32_fa9_8_and0 = s_csamul_cla32_and9_8 & s_csamul_cla32_fa10_7_xor1;
  assign s_csamul_cla32_fa9_8_xor1 = s_csamul_cla32_fa9_8_xor0 ^ s_csamul_cla32_fa9_7_or0;
  assign s_csamul_cla32_fa9_8_and1 = s_csamul_cla32_fa9_8_xor0 & s_csamul_cla32_fa9_7_or0;
  assign s_csamul_cla32_fa9_8_or0 = s_csamul_cla32_fa9_8_and0 | s_csamul_cla32_fa9_8_and1;
  assign s_csamul_cla32_and10_8 = a[10] & b[8];
  assign s_csamul_cla32_fa10_8_xor0 = s_csamul_cla32_and10_8 ^ s_csamul_cla32_fa11_7_xor1;
  assign s_csamul_cla32_fa10_8_and0 = s_csamul_cla32_and10_8 & s_csamul_cla32_fa11_7_xor1;
  assign s_csamul_cla32_fa10_8_xor1 = s_csamul_cla32_fa10_8_xor0 ^ s_csamul_cla32_fa10_7_or0;
  assign s_csamul_cla32_fa10_8_and1 = s_csamul_cla32_fa10_8_xor0 & s_csamul_cla32_fa10_7_or0;
  assign s_csamul_cla32_fa10_8_or0 = s_csamul_cla32_fa10_8_and0 | s_csamul_cla32_fa10_8_and1;
  assign s_csamul_cla32_and11_8 = a[11] & b[8];
  assign s_csamul_cla32_fa11_8_xor0 = s_csamul_cla32_and11_8 ^ s_csamul_cla32_fa12_7_xor1;
  assign s_csamul_cla32_fa11_8_and0 = s_csamul_cla32_and11_8 & s_csamul_cla32_fa12_7_xor1;
  assign s_csamul_cla32_fa11_8_xor1 = s_csamul_cla32_fa11_8_xor0 ^ s_csamul_cla32_fa11_7_or0;
  assign s_csamul_cla32_fa11_8_and1 = s_csamul_cla32_fa11_8_xor0 & s_csamul_cla32_fa11_7_or0;
  assign s_csamul_cla32_fa11_8_or0 = s_csamul_cla32_fa11_8_and0 | s_csamul_cla32_fa11_8_and1;
  assign s_csamul_cla32_and12_8 = a[12] & b[8];
  assign s_csamul_cla32_fa12_8_xor0 = s_csamul_cla32_and12_8 ^ s_csamul_cla32_fa13_7_xor1;
  assign s_csamul_cla32_fa12_8_and0 = s_csamul_cla32_and12_8 & s_csamul_cla32_fa13_7_xor1;
  assign s_csamul_cla32_fa12_8_xor1 = s_csamul_cla32_fa12_8_xor0 ^ s_csamul_cla32_fa12_7_or0;
  assign s_csamul_cla32_fa12_8_and1 = s_csamul_cla32_fa12_8_xor0 & s_csamul_cla32_fa12_7_or0;
  assign s_csamul_cla32_fa12_8_or0 = s_csamul_cla32_fa12_8_and0 | s_csamul_cla32_fa12_8_and1;
  assign s_csamul_cla32_and13_8 = a[13] & b[8];
  assign s_csamul_cla32_fa13_8_xor0 = s_csamul_cla32_and13_8 ^ s_csamul_cla32_fa14_7_xor1;
  assign s_csamul_cla32_fa13_8_and0 = s_csamul_cla32_and13_8 & s_csamul_cla32_fa14_7_xor1;
  assign s_csamul_cla32_fa13_8_xor1 = s_csamul_cla32_fa13_8_xor0 ^ s_csamul_cla32_fa13_7_or0;
  assign s_csamul_cla32_fa13_8_and1 = s_csamul_cla32_fa13_8_xor0 & s_csamul_cla32_fa13_7_or0;
  assign s_csamul_cla32_fa13_8_or0 = s_csamul_cla32_fa13_8_and0 | s_csamul_cla32_fa13_8_and1;
  assign s_csamul_cla32_and14_8 = a[14] & b[8];
  assign s_csamul_cla32_fa14_8_xor0 = s_csamul_cla32_and14_8 ^ s_csamul_cla32_fa15_7_xor1;
  assign s_csamul_cla32_fa14_8_and0 = s_csamul_cla32_and14_8 & s_csamul_cla32_fa15_7_xor1;
  assign s_csamul_cla32_fa14_8_xor1 = s_csamul_cla32_fa14_8_xor0 ^ s_csamul_cla32_fa14_7_or0;
  assign s_csamul_cla32_fa14_8_and1 = s_csamul_cla32_fa14_8_xor0 & s_csamul_cla32_fa14_7_or0;
  assign s_csamul_cla32_fa14_8_or0 = s_csamul_cla32_fa14_8_and0 | s_csamul_cla32_fa14_8_and1;
  assign s_csamul_cla32_and15_8 = a[15] & b[8];
  assign s_csamul_cla32_fa15_8_xor0 = s_csamul_cla32_and15_8 ^ s_csamul_cla32_fa16_7_xor1;
  assign s_csamul_cla32_fa15_8_and0 = s_csamul_cla32_and15_8 & s_csamul_cla32_fa16_7_xor1;
  assign s_csamul_cla32_fa15_8_xor1 = s_csamul_cla32_fa15_8_xor0 ^ s_csamul_cla32_fa15_7_or0;
  assign s_csamul_cla32_fa15_8_and1 = s_csamul_cla32_fa15_8_xor0 & s_csamul_cla32_fa15_7_or0;
  assign s_csamul_cla32_fa15_8_or0 = s_csamul_cla32_fa15_8_and0 | s_csamul_cla32_fa15_8_and1;
  assign s_csamul_cla32_and16_8 = a[16] & b[8];
  assign s_csamul_cla32_fa16_8_xor0 = s_csamul_cla32_and16_8 ^ s_csamul_cla32_fa17_7_xor1;
  assign s_csamul_cla32_fa16_8_and0 = s_csamul_cla32_and16_8 & s_csamul_cla32_fa17_7_xor1;
  assign s_csamul_cla32_fa16_8_xor1 = s_csamul_cla32_fa16_8_xor0 ^ s_csamul_cla32_fa16_7_or0;
  assign s_csamul_cla32_fa16_8_and1 = s_csamul_cla32_fa16_8_xor0 & s_csamul_cla32_fa16_7_or0;
  assign s_csamul_cla32_fa16_8_or0 = s_csamul_cla32_fa16_8_and0 | s_csamul_cla32_fa16_8_and1;
  assign s_csamul_cla32_and17_8 = a[17] & b[8];
  assign s_csamul_cla32_fa17_8_xor0 = s_csamul_cla32_and17_8 ^ s_csamul_cla32_fa18_7_xor1;
  assign s_csamul_cla32_fa17_8_and0 = s_csamul_cla32_and17_8 & s_csamul_cla32_fa18_7_xor1;
  assign s_csamul_cla32_fa17_8_xor1 = s_csamul_cla32_fa17_8_xor0 ^ s_csamul_cla32_fa17_7_or0;
  assign s_csamul_cla32_fa17_8_and1 = s_csamul_cla32_fa17_8_xor0 & s_csamul_cla32_fa17_7_or0;
  assign s_csamul_cla32_fa17_8_or0 = s_csamul_cla32_fa17_8_and0 | s_csamul_cla32_fa17_8_and1;
  assign s_csamul_cla32_and18_8 = a[18] & b[8];
  assign s_csamul_cla32_fa18_8_xor0 = s_csamul_cla32_and18_8 ^ s_csamul_cla32_fa19_7_xor1;
  assign s_csamul_cla32_fa18_8_and0 = s_csamul_cla32_and18_8 & s_csamul_cla32_fa19_7_xor1;
  assign s_csamul_cla32_fa18_8_xor1 = s_csamul_cla32_fa18_8_xor0 ^ s_csamul_cla32_fa18_7_or0;
  assign s_csamul_cla32_fa18_8_and1 = s_csamul_cla32_fa18_8_xor0 & s_csamul_cla32_fa18_7_or0;
  assign s_csamul_cla32_fa18_8_or0 = s_csamul_cla32_fa18_8_and0 | s_csamul_cla32_fa18_8_and1;
  assign s_csamul_cla32_and19_8 = a[19] & b[8];
  assign s_csamul_cla32_fa19_8_xor0 = s_csamul_cla32_and19_8 ^ s_csamul_cla32_fa20_7_xor1;
  assign s_csamul_cla32_fa19_8_and0 = s_csamul_cla32_and19_8 & s_csamul_cla32_fa20_7_xor1;
  assign s_csamul_cla32_fa19_8_xor1 = s_csamul_cla32_fa19_8_xor0 ^ s_csamul_cla32_fa19_7_or0;
  assign s_csamul_cla32_fa19_8_and1 = s_csamul_cla32_fa19_8_xor0 & s_csamul_cla32_fa19_7_or0;
  assign s_csamul_cla32_fa19_8_or0 = s_csamul_cla32_fa19_8_and0 | s_csamul_cla32_fa19_8_and1;
  assign s_csamul_cla32_and20_8 = a[20] & b[8];
  assign s_csamul_cla32_fa20_8_xor0 = s_csamul_cla32_and20_8 ^ s_csamul_cla32_fa21_7_xor1;
  assign s_csamul_cla32_fa20_8_and0 = s_csamul_cla32_and20_8 & s_csamul_cla32_fa21_7_xor1;
  assign s_csamul_cla32_fa20_8_xor1 = s_csamul_cla32_fa20_8_xor0 ^ s_csamul_cla32_fa20_7_or0;
  assign s_csamul_cla32_fa20_8_and1 = s_csamul_cla32_fa20_8_xor0 & s_csamul_cla32_fa20_7_or0;
  assign s_csamul_cla32_fa20_8_or0 = s_csamul_cla32_fa20_8_and0 | s_csamul_cla32_fa20_8_and1;
  assign s_csamul_cla32_and21_8 = a[21] & b[8];
  assign s_csamul_cla32_fa21_8_xor0 = s_csamul_cla32_and21_8 ^ s_csamul_cla32_fa22_7_xor1;
  assign s_csamul_cla32_fa21_8_and0 = s_csamul_cla32_and21_8 & s_csamul_cla32_fa22_7_xor1;
  assign s_csamul_cla32_fa21_8_xor1 = s_csamul_cla32_fa21_8_xor0 ^ s_csamul_cla32_fa21_7_or0;
  assign s_csamul_cla32_fa21_8_and1 = s_csamul_cla32_fa21_8_xor0 & s_csamul_cla32_fa21_7_or0;
  assign s_csamul_cla32_fa21_8_or0 = s_csamul_cla32_fa21_8_and0 | s_csamul_cla32_fa21_8_and1;
  assign s_csamul_cla32_and22_8 = a[22] & b[8];
  assign s_csamul_cla32_fa22_8_xor0 = s_csamul_cla32_and22_8 ^ s_csamul_cla32_fa23_7_xor1;
  assign s_csamul_cla32_fa22_8_and0 = s_csamul_cla32_and22_8 & s_csamul_cla32_fa23_7_xor1;
  assign s_csamul_cla32_fa22_8_xor1 = s_csamul_cla32_fa22_8_xor0 ^ s_csamul_cla32_fa22_7_or0;
  assign s_csamul_cla32_fa22_8_and1 = s_csamul_cla32_fa22_8_xor0 & s_csamul_cla32_fa22_7_or0;
  assign s_csamul_cla32_fa22_8_or0 = s_csamul_cla32_fa22_8_and0 | s_csamul_cla32_fa22_8_and1;
  assign s_csamul_cla32_and23_8 = a[23] & b[8];
  assign s_csamul_cla32_fa23_8_xor0 = s_csamul_cla32_and23_8 ^ s_csamul_cla32_fa24_7_xor1;
  assign s_csamul_cla32_fa23_8_and0 = s_csamul_cla32_and23_8 & s_csamul_cla32_fa24_7_xor1;
  assign s_csamul_cla32_fa23_8_xor1 = s_csamul_cla32_fa23_8_xor0 ^ s_csamul_cla32_fa23_7_or0;
  assign s_csamul_cla32_fa23_8_and1 = s_csamul_cla32_fa23_8_xor0 & s_csamul_cla32_fa23_7_or0;
  assign s_csamul_cla32_fa23_8_or0 = s_csamul_cla32_fa23_8_and0 | s_csamul_cla32_fa23_8_and1;
  assign s_csamul_cla32_and24_8 = a[24] & b[8];
  assign s_csamul_cla32_fa24_8_xor0 = s_csamul_cla32_and24_8 ^ s_csamul_cla32_fa25_7_xor1;
  assign s_csamul_cla32_fa24_8_and0 = s_csamul_cla32_and24_8 & s_csamul_cla32_fa25_7_xor1;
  assign s_csamul_cla32_fa24_8_xor1 = s_csamul_cla32_fa24_8_xor0 ^ s_csamul_cla32_fa24_7_or0;
  assign s_csamul_cla32_fa24_8_and1 = s_csamul_cla32_fa24_8_xor0 & s_csamul_cla32_fa24_7_or0;
  assign s_csamul_cla32_fa24_8_or0 = s_csamul_cla32_fa24_8_and0 | s_csamul_cla32_fa24_8_and1;
  assign s_csamul_cla32_and25_8 = a[25] & b[8];
  assign s_csamul_cla32_fa25_8_xor0 = s_csamul_cla32_and25_8 ^ s_csamul_cla32_fa26_7_xor1;
  assign s_csamul_cla32_fa25_8_and0 = s_csamul_cla32_and25_8 & s_csamul_cla32_fa26_7_xor1;
  assign s_csamul_cla32_fa25_8_xor1 = s_csamul_cla32_fa25_8_xor0 ^ s_csamul_cla32_fa25_7_or0;
  assign s_csamul_cla32_fa25_8_and1 = s_csamul_cla32_fa25_8_xor0 & s_csamul_cla32_fa25_7_or0;
  assign s_csamul_cla32_fa25_8_or0 = s_csamul_cla32_fa25_8_and0 | s_csamul_cla32_fa25_8_and1;
  assign s_csamul_cla32_and26_8 = a[26] & b[8];
  assign s_csamul_cla32_fa26_8_xor0 = s_csamul_cla32_and26_8 ^ s_csamul_cla32_fa27_7_xor1;
  assign s_csamul_cla32_fa26_8_and0 = s_csamul_cla32_and26_8 & s_csamul_cla32_fa27_7_xor1;
  assign s_csamul_cla32_fa26_8_xor1 = s_csamul_cla32_fa26_8_xor0 ^ s_csamul_cla32_fa26_7_or0;
  assign s_csamul_cla32_fa26_8_and1 = s_csamul_cla32_fa26_8_xor0 & s_csamul_cla32_fa26_7_or0;
  assign s_csamul_cla32_fa26_8_or0 = s_csamul_cla32_fa26_8_and0 | s_csamul_cla32_fa26_8_and1;
  assign s_csamul_cla32_and27_8 = a[27] & b[8];
  assign s_csamul_cla32_fa27_8_xor0 = s_csamul_cla32_and27_8 ^ s_csamul_cla32_fa28_7_xor1;
  assign s_csamul_cla32_fa27_8_and0 = s_csamul_cla32_and27_8 & s_csamul_cla32_fa28_7_xor1;
  assign s_csamul_cla32_fa27_8_xor1 = s_csamul_cla32_fa27_8_xor0 ^ s_csamul_cla32_fa27_7_or0;
  assign s_csamul_cla32_fa27_8_and1 = s_csamul_cla32_fa27_8_xor0 & s_csamul_cla32_fa27_7_or0;
  assign s_csamul_cla32_fa27_8_or0 = s_csamul_cla32_fa27_8_and0 | s_csamul_cla32_fa27_8_and1;
  assign s_csamul_cla32_and28_8 = a[28] & b[8];
  assign s_csamul_cla32_fa28_8_xor0 = s_csamul_cla32_and28_8 ^ s_csamul_cla32_fa29_7_xor1;
  assign s_csamul_cla32_fa28_8_and0 = s_csamul_cla32_and28_8 & s_csamul_cla32_fa29_7_xor1;
  assign s_csamul_cla32_fa28_8_xor1 = s_csamul_cla32_fa28_8_xor0 ^ s_csamul_cla32_fa28_7_or0;
  assign s_csamul_cla32_fa28_8_and1 = s_csamul_cla32_fa28_8_xor0 & s_csamul_cla32_fa28_7_or0;
  assign s_csamul_cla32_fa28_8_or0 = s_csamul_cla32_fa28_8_and0 | s_csamul_cla32_fa28_8_and1;
  assign s_csamul_cla32_and29_8 = a[29] & b[8];
  assign s_csamul_cla32_fa29_8_xor0 = s_csamul_cla32_and29_8 ^ s_csamul_cla32_fa30_7_xor1;
  assign s_csamul_cla32_fa29_8_and0 = s_csamul_cla32_and29_8 & s_csamul_cla32_fa30_7_xor1;
  assign s_csamul_cla32_fa29_8_xor1 = s_csamul_cla32_fa29_8_xor0 ^ s_csamul_cla32_fa29_7_or0;
  assign s_csamul_cla32_fa29_8_and1 = s_csamul_cla32_fa29_8_xor0 & s_csamul_cla32_fa29_7_or0;
  assign s_csamul_cla32_fa29_8_or0 = s_csamul_cla32_fa29_8_and0 | s_csamul_cla32_fa29_8_and1;
  assign s_csamul_cla32_and30_8 = a[30] & b[8];
  assign s_csamul_cla32_fa30_8_xor0 = s_csamul_cla32_and30_8 ^ s_csamul_cla32_ha31_7_xor0;
  assign s_csamul_cla32_fa30_8_and0 = s_csamul_cla32_and30_8 & s_csamul_cla32_ha31_7_xor0;
  assign s_csamul_cla32_fa30_8_xor1 = s_csamul_cla32_fa30_8_xor0 ^ s_csamul_cla32_fa30_7_or0;
  assign s_csamul_cla32_fa30_8_and1 = s_csamul_cla32_fa30_8_xor0 & s_csamul_cla32_fa30_7_or0;
  assign s_csamul_cla32_fa30_8_or0 = s_csamul_cla32_fa30_8_and0 | s_csamul_cla32_fa30_8_and1;
  assign s_csamul_cla32_nand31_8 = ~(a[31] & b[8]);
  assign s_csamul_cla32_ha31_8_xor0 = s_csamul_cla32_nand31_8 ^ s_csamul_cla32_ha31_7_and0;
  assign s_csamul_cla32_ha31_8_and0 = s_csamul_cla32_nand31_8 & s_csamul_cla32_ha31_7_and0;
  assign s_csamul_cla32_and0_9 = a[0] & b[9];
  assign s_csamul_cla32_fa0_9_xor0 = s_csamul_cla32_and0_9 ^ s_csamul_cla32_fa1_8_xor1;
  assign s_csamul_cla32_fa0_9_and0 = s_csamul_cla32_and0_9 & s_csamul_cla32_fa1_8_xor1;
  assign s_csamul_cla32_fa0_9_xor1 = s_csamul_cla32_fa0_9_xor0 ^ s_csamul_cla32_fa0_8_or0;
  assign s_csamul_cla32_fa0_9_and1 = s_csamul_cla32_fa0_9_xor0 & s_csamul_cla32_fa0_8_or0;
  assign s_csamul_cla32_fa0_9_or0 = s_csamul_cla32_fa0_9_and0 | s_csamul_cla32_fa0_9_and1;
  assign s_csamul_cla32_and1_9 = a[1] & b[9];
  assign s_csamul_cla32_fa1_9_xor0 = s_csamul_cla32_and1_9 ^ s_csamul_cla32_fa2_8_xor1;
  assign s_csamul_cla32_fa1_9_and0 = s_csamul_cla32_and1_9 & s_csamul_cla32_fa2_8_xor1;
  assign s_csamul_cla32_fa1_9_xor1 = s_csamul_cla32_fa1_9_xor0 ^ s_csamul_cla32_fa1_8_or0;
  assign s_csamul_cla32_fa1_9_and1 = s_csamul_cla32_fa1_9_xor0 & s_csamul_cla32_fa1_8_or0;
  assign s_csamul_cla32_fa1_9_or0 = s_csamul_cla32_fa1_9_and0 | s_csamul_cla32_fa1_9_and1;
  assign s_csamul_cla32_and2_9 = a[2] & b[9];
  assign s_csamul_cla32_fa2_9_xor0 = s_csamul_cla32_and2_9 ^ s_csamul_cla32_fa3_8_xor1;
  assign s_csamul_cla32_fa2_9_and0 = s_csamul_cla32_and2_9 & s_csamul_cla32_fa3_8_xor1;
  assign s_csamul_cla32_fa2_9_xor1 = s_csamul_cla32_fa2_9_xor0 ^ s_csamul_cla32_fa2_8_or0;
  assign s_csamul_cla32_fa2_9_and1 = s_csamul_cla32_fa2_9_xor0 & s_csamul_cla32_fa2_8_or0;
  assign s_csamul_cla32_fa2_9_or0 = s_csamul_cla32_fa2_9_and0 | s_csamul_cla32_fa2_9_and1;
  assign s_csamul_cla32_and3_9 = a[3] & b[9];
  assign s_csamul_cla32_fa3_9_xor0 = s_csamul_cla32_and3_9 ^ s_csamul_cla32_fa4_8_xor1;
  assign s_csamul_cla32_fa3_9_and0 = s_csamul_cla32_and3_9 & s_csamul_cla32_fa4_8_xor1;
  assign s_csamul_cla32_fa3_9_xor1 = s_csamul_cla32_fa3_9_xor0 ^ s_csamul_cla32_fa3_8_or0;
  assign s_csamul_cla32_fa3_9_and1 = s_csamul_cla32_fa3_9_xor0 & s_csamul_cla32_fa3_8_or0;
  assign s_csamul_cla32_fa3_9_or0 = s_csamul_cla32_fa3_9_and0 | s_csamul_cla32_fa3_9_and1;
  assign s_csamul_cla32_and4_9 = a[4] & b[9];
  assign s_csamul_cla32_fa4_9_xor0 = s_csamul_cla32_and4_9 ^ s_csamul_cla32_fa5_8_xor1;
  assign s_csamul_cla32_fa4_9_and0 = s_csamul_cla32_and4_9 & s_csamul_cla32_fa5_8_xor1;
  assign s_csamul_cla32_fa4_9_xor1 = s_csamul_cla32_fa4_9_xor0 ^ s_csamul_cla32_fa4_8_or0;
  assign s_csamul_cla32_fa4_9_and1 = s_csamul_cla32_fa4_9_xor0 & s_csamul_cla32_fa4_8_or0;
  assign s_csamul_cla32_fa4_9_or0 = s_csamul_cla32_fa4_9_and0 | s_csamul_cla32_fa4_9_and1;
  assign s_csamul_cla32_and5_9 = a[5] & b[9];
  assign s_csamul_cla32_fa5_9_xor0 = s_csamul_cla32_and5_9 ^ s_csamul_cla32_fa6_8_xor1;
  assign s_csamul_cla32_fa5_9_and0 = s_csamul_cla32_and5_9 & s_csamul_cla32_fa6_8_xor1;
  assign s_csamul_cla32_fa5_9_xor1 = s_csamul_cla32_fa5_9_xor0 ^ s_csamul_cla32_fa5_8_or0;
  assign s_csamul_cla32_fa5_9_and1 = s_csamul_cla32_fa5_9_xor0 & s_csamul_cla32_fa5_8_or0;
  assign s_csamul_cla32_fa5_9_or0 = s_csamul_cla32_fa5_9_and0 | s_csamul_cla32_fa5_9_and1;
  assign s_csamul_cla32_and6_9 = a[6] & b[9];
  assign s_csamul_cla32_fa6_9_xor0 = s_csamul_cla32_and6_9 ^ s_csamul_cla32_fa7_8_xor1;
  assign s_csamul_cla32_fa6_9_and0 = s_csamul_cla32_and6_9 & s_csamul_cla32_fa7_8_xor1;
  assign s_csamul_cla32_fa6_9_xor1 = s_csamul_cla32_fa6_9_xor0 ^ s_csamul_cla32_fa6_8_or0;
  assign s_csamul_cla32_fa6_9_and1 = s_csamul_cla32_fa6_9_xor0 & s_csamul_cla32_fa6_8_or0;
  assign s_csamul_cla32_fa6_9_or0 = s_csamul_cla32_fa6_9_and0 | s_csamul_cla32_fa6_9_and1;
  assign s_csamul_cla32_and7_9 = a[7] & b[9];
  assign s_csamul_cla32_fa7_9_xor0 = s_csamul_cla32_and7_9 ^ s_csamul_cla32_fa8_8_xor1;
  assign s_csamul_cla32_fa7_9_and0 = s_csamul_cla32_and7_9 & s_csamul_cla32_fa8_8_xor1;
  assign s_csamul_cla32_fa7_9_xor1 = s_csamul_cla32_fa7_9_xor0 ^ s_csamul_cla32_fa7_8_or0;
  assign s_csamul_cla32_fa7_9_and1 = s_csamul_cla32_fa7_9_xor0 & s_csamul_cla32_fa7_8_or0;
  assign s_csamul_cla32_fa7_9_or0 = s_csamul_cla32_fa7_9_and0 | s_csamul_cla32_fa7_9_and1;
  assign s_csamul_cla32_and8_9 = a[8] & b[9];
  assign s_csamul_cla32_fa8_9_xor0 = s_csamul_cla32_and8_9 ^ s_csamul_cla32_fa9_8_xor1;
  assign s_csamul_cla32_fa8_9_and0 = s_csamul_cla32_and8_9 & s_csamul_cla32_fa9_8_xor1;
  assign s_csamul_cla32_fa8_9_xor1 = s_csamul_cla32_fa8_9_xor0 ^ s_csamul_cla32_fa8_8_or0;
  assign s_csamul_cla32_fa8_9_and1 = s_csamul_cla32_fa8_9_xor0 & s_csamul_cla32_fa8_8_or0;
  assign s_csamul_cla32_fa8_9_or0 = s_csamul_cla32_fa8_9_and0 | s_csamul_cla32_fa8_9_and1;
  assign s_csamul_cla32_and9_9 = a[9] & b[9];
  assign s_csamul_cla32_fa9_9_xor0 = s_csamul_cla32_and9_9 ^ s_csamul_cla32_fa10_8_xor1;
  assign s_csamul_cla32_fa9_9_and0 = s_csamul_cla32_and9_9 & s_csamul_cla32_fa10_8_xor1;
  assign s_csamul_cla32_fa9_9_xor1 = s_csamul_cla32_fa9_9_xor0 ^ s_csamul_cla32_fa9_8_or0;
  assign s_csamul_cla32_fa9_9_and1 = s_csamul_cla32_fa9_9_xor0 & s_csamul_cla32_fa9_8_or0;
  assign s_csamul_cla32_fa9_9_or0 = s_csamul_cla32_fa9_9_and0 | s_csamul_cla32_fa9_9_and1;
  assign s_csamul_cla32_and10_9 = a[10] & b[9];
  assign s_csamul_cla32_fa10_9_xor0 = s_csamul_cla32_and10_9 ^ s_csamul_cla32_fa11_8_xor1;
  assign s_csamul_cla32_fa10_9_and0 = s_csamul_cla32_and10_9 & s_csamul_cla32_fa11_8_xor1;
  assign s_csamul_cla32_fa10_9_xor1 = s_csamul_cla32_fa10_9_xor0 ^ s_csamul_cla32_fa10_8_or0;
  assign s_csamul_cla32_fa10_9_and1 = s_csamul_cla32_fa10_9_xor0 & s_csamul_cla32_fa10_8_or0;
  assign s_csamul_cla32_fa10_9_or0 = s_csamul_cla32_fa10_9_and0 | s_csamul_cla32_fa10_9_and1;
  assign s_csamul_cla32_and11_9 = a[11] & b[9];
  assign s_csamul_cla32_fa11_9_xor0 = s_csamul_cla32_and11_9 ^ s_csamul_cla32_fa12_8_xor1;
  assign s_csamul_cla32_fa11_9_and0 = s_csamul_cla32_and11_9 & s_csamul_cla32_fa12_8_xor1;
  assign s_csamul_cla32_fa11_9_xor1 = s_csamul_cla32_fa11_9_xor0 ^ s_csamul_cla32_fa11_8_or0;
  assign s_csamul_cla32_fa11_9_and1 = s_csamul_cla32_fa11_9_xor0 & s_csamul_cla32_fa11_8_or0;
  assign s_csamul_cla32_fa11_9_or0 = s_csamul_cla32_fa11_9_and0 | s_csamul_cla32_fa11_9_and1;
  assign s_csamul_cla32_and12_9 = a[12] & b[9];
  assign s_csamul_cla32_fa12_9_xor0 = s_csamul_cla32_and12_9 ^ s_csamul_cla32_fa13_8_xor1;
  assign s_csamul_cla32_fa12_9_and0 = s_csamul_cla32_and12_9 & s_csamul_cla32_fa13_8_xor1;
  assign s_csamul_cla32_fa12_9_xor1 = s_csamul_cla32_fa12_9_xor0 ^ s_csamul_cla32_fa12_8_or0;
  assign s_csamul_cla32_fa12_9_and1 = s_csamul_cla32_fa12_9_xor0 & s_csamul_cla32_fa12_8_or0;
  assign s_csamul_cla32_fa12_9_or0 = s_csamul_cla32_fa12_9_and0 | s_csamul_cla32_fa12_9_and1;
  assign s_csamul_cla32_and13_9 = a[13] & b[9];
  assign s_csamul_cla32_fa13_9_xor0 = s_csamul_cla32_and13_9 ^ s_csamul_cla32_fa14_8_xor1;
  assign s_csamul_cla32_fa13_9_and0 = s_csamul_cla32_and13_9 & s_csamul_cla32_fa14_8_xor1;
  assign s_csamul_cla32_fa13_9_xor1 = s_csamul_cla32_fa13_9_xor0 ^ s_csamul_cla32_fa13_8_or0;
  assign s_csamul_cla32_fa13_9_and1 = s_csamul_cla32_fa13_9_xor0 & s_csamul_cla32_fa13_8_or0;
  assign s_csamul_cla32_fa13_9_or0 = s_csamul_cla32_fa13_9_and0 | s_csamul_cla32_fa13_9_and1;
  assign s_csamul_cla32_and14_9 = a[14] & b[9];
  assign s_csamul_cla32_fa14_9_xor0 = s_csamul_cla32_and14_9 ^ s_csamul_cla32_fa15_8_xor1;
  assign s_csamul_cla32_fa14_9_and0 = s_csamul_cla32_and14_9 & s_csamul_cla32_fa15_8_xor1;
  assign s_csamul_cla32_fa14_9_xor1 = s_csamul_cla32_fa14_9_xor0 ^ s_csamul_cla32_fa14_8_or0;
  assign s_csamul_cla32_fa14_9_and1 = s_csamul_cla32_fa14_9_xor0 & s_csamul_cla32_fa14_8_or0;
  assign s_csamul_cla32_fa14_9_or0 = s_csamul_cla32_fa14_9_and0 | s_csamul_cla32_fa14_9_and1;
  assign s_csamul_cla32_and15_9 = a[15] & b[9];
  assign s_csamul_cla32_fa15_9_xor0 = s_csamul_cla32_and15_9 ^ s_csamul_cla32_fa16_8_xor1;
  assign s_csamul_cla32_fa15_9_and0 = s_csamul_cla32_and15_9 & s_csamul_cla32_fa16_8_xor1;
  assign s_csamul_cla32_fa15_9_xor1 = s_csamul_cla32_fa15_9_xor0 ^ s_csamul_cla32_fa15_8_or0;
  assign s_csamul_cla32_fa15_9_and1 = s_csamul_cla32_fa15_9_xor0 & s_csamul_cla32_fa15_8_or0;
  assign s_csamul_cla32_fa15_9_or0 = s_csamul_cla32_fa15_9_and0 | s_csamul_cla32_fa15_9_and1;
  assign s_csamul_cla32_and16_9 = a[16] & b[9];
  assign s_csamul_cla32_fa16_9_xor0 = s_csamul_cla32_and16_9 ^ s_csamul_cla32_fa17_8_xor1;
  assign s_csamul_cla32_fa16_9_and0 = s_csamul_cla32_and16_9 & s_csamul_cla32_fa17_8_xor1;
  assign s_csamul_cla32_fa16_9_xor1 = s_csamul_cla32_fa16_9_xor0 ^ s_csamul_cla32_fa16_8_or0;
  assign s_csamul_cla32_fa16_9_and1 = s_csamul_cla32_fa16_9_xor0 & s_csamul_cla32_fa16_8_or0;
  assign s_csamul_cla32_fa16_9_or0 = s_csamul_cla32_fa16_9_and0 | s_csamul_cla32_fa16_9_and1;
  assign s_csamul_cla32_and17_9 = a[17] & b[9];
  assign s_csamul_cla32_fa17_9_xor0 = s_csamul_cla32_and17_9 ^ s_csamul_cla32_fa18_8_xor1;
  assign s_csamul_cla32_fa17_9_and0 = s_csamul_cla32_and17_9 & s_csamul_cla32_fa18_8_xor1;
  assign s_csamul_cla32_fa17_9_xor1 = s_csamul_cla32_fa17_9_xor0 ^ s_csamul_cla32_fa17_8_or0;
  assign s_csamul_cla32_fa17_9_and1 = s_csamul_cla32_fa17_9_xor0 & s_csamul_cla32_fa17_8_or0;
  assign s_csamul_cla32_fa17_9_or0 = s_csamul_cla32_fa17_9_and0 | s_csamul_cla32_fa17_9_and1;
  assign s_csamul_cla32_and18_9 = a[18] & b[9];
  assign s_csamul_cla32_fa18_9_xor0 = s_csamul_cla32_and18_9 ^ s_csamul_cla32_fa19_8_xor1;
  assign s_csamul_cla32_fa18_9_and0 = s_csamul_cla32_and18_9 & s_csamul_cla32_fa19_8_xor1;
  assign s_csamul_cla32_fa18_9_xor1 = s_csamul_cla32_fa18_9_xor0 ^ s_csamul_cla32_fa18_8_or0;
  assign s_csamul_cla32_fa18_9_and1 = s_csamul_cla32_fa18_9_xor0 & s_csamul_cla32_fa18_8_or0;
  assign s_csamul_cla32_fa18_9_or0 = s_csamul_cla32_fa18_9_and0 | s_csamul_cla32_fa18_9_and1;
  assign s_csamul_cla32_and19_9 = a[19] & b[9];
  assign s_csamul_cla32_fa19_9_xor0 = s_csamul_cla32_and19_9 ^ s_csamul_cla32_fa20_8_xor1;
  assign s_csamul_cla32_fa19_9_and0 = s_csamul_cla32_and19_9 & s_csamul_cla32_fa20_8_xor1;
  assign s_csamul_cla32_fa19_9_xor1 = s_csamul_cla32_fa19_9_xor0 ^ s_csamul_cla32_fa19_8_or0;
  assign s_csamul_cla32_fa19_9_and1 = s_csamul_cla32_fa19_9_xor0 & s_csamul_cla32_fa19_8_or0;
  assign s_csamul_cla32_fa19_9_or0 = s_csamul_cla32_fa19_9_and0 | s_csamul_cla32_fa19_9_and1;
  assign s_csamul_cla32_and20_9 = a[20] & b[9];
  assign s_csamul_cla32_fa20_9_xor0 = s_csamul_cla32_and20_9 ^ s_csamul_cla32_fa21_8_xor1;
  assign s_csamul_cla32_fa20_9_and0 = s_csamul_cla32_and20_9 & s_csamul_cla32_fa21_8_xor1;
  assign s_csamul_cla32_fa20_9_xor1 = s_csamul_cla32_fa20_9_xor0 ^ s_csamul_cla32_fa20_8_or0;
  assign s_csamul_cla32_fa20_9_and1 = s_csamul_cla32_fa20_9_xor0 & s_csamul_cla32_fa20_8_or0;
  assign s_csamul_cla32_fa20_9_or0 = s_csamul_cla32_fa20_9_and0 | s_csamul_cla32_fa20_9_and1;
  assign s_csamul_cla32_and21_9 = a[21] & b[9];
  assign s_csamul_cla32_fa21_9_xor0 = s_csamul_cla32_and21_9 ^ s_csamul_cla32_fa22_8_xor1;
  assign s_csamul_cla32_fa21_9_and0 = s_csamul_cla32_and21_9 & s_csamul_cla32_fa22_8_xor1;
  assign s_csamul_cla32_fa21_9_xor1 = s_csamul_cla32_fa21_9_xor0 ^ s_csamul_cla32_fa21_8_or0;
  assign s_csamul_cla32_fa21_9_and1 = s_csamul_cla32_fa21_9_xor0 & s_csamul_cla32_fa21_8_or0;
  assign s_csamul_cla32_fa21_9_or0 = s_csamul_cla32_fa21_9_and0 | s_csamul_cla32_fa21_9_and1;
  assign s_csamul_cla32_and22_9 = a[22] & b[9];
  assign s_csamul_cla32_fa22_9_xor0 = s_csamul_cla32_and22_9 ^ s_csamul_cla32_fa23_8_xor1;
  assign s_csamul_cla32_fa22_9_and0 = s_csamul_cla32_and22_9 & s_csamul_cla32_fa23_8_xor1;
  assign s_csamul_cla32_fa22_9_xor1 = s_csamul_cla32_fa22_9_xor0 ^ s_csamul_cla32_fa22_8_or0;
  assign s_csamul_cla32_fa22_9_and1 = s_csamul_cla32_fa22_9_xor0 & s_csamul_cla32_fa22_8_or0;
  assign s_csamul_cla32_fa22_9_or0 = s_csamul_cla32_fa22_9_and0 | s_csamul_cla32_fa22_9_and1;
  assign s_csamul_cla32_and23_9 = a[23] & b[9];
  assign s_csamul_cla32_fa23_9_xor0 = s_csamul_cla32_and23_9 ^ s_csamul_cla32_fa24_8_xor1;
  assign s_csamul_cla32_fa23_9_and0 = s_csamul_cla32_and23_9 & s_csamul_cla32_fa24_8_xor1;
  assign s_csamul_cla32_fa23_9_xor1 = s_csamul_cla32_fa23_9_xor0 ^ s_csamul_cla32_fa23_8_or0;
  assign s_csamul_cla32_fa23_9_and1 = s_csamul_cla32_fa23_9_xor0 & s_csamul_cla32_fa23_8_or0;
  assign s_csamul_cla32_fa23_9_or0 = s_csamul_cla32_fa23_9_and0 | s_csamul_cla32_fa23_9_and1;
  assign s_csamul_cla32_and24_9 = a[24] & b[9];
  assign s_csamul_cla32_fa24_9_xor0 = s_csamul_cla32_and24_9 ^ s_csamul_cla32_fa25_8_xor1;
  assign s_csamul_cla32_fa24_9_and0 = s_csamul_cla32_and24_9 & s_csamul_cla32_fa25_8_xor1;
  assign s_csamul_cla32_fa24_9_xor1 = s_csamul_cla32_fa24_9_xor0 ^ s_csamul_cla32_fa24_8_or0;
  assign s_csamul_cla32_fa24_9_and1 = s_csamul_cla32_fa24_9_xor0 & s_csamul_cla32_fa24_8_or0;
  assign s_csamul_cla32_fa24_9_or0 = s_csamul_cla32_fa24_9_and0 | s_csamul_cla32_fa24_9_and1;
  assign s_csamul_cla32_and25_9 = a[25] & b[9];
  assign s_csamul_cla32_fa25_9_xor0 = s_csamul_cla32_and25_9 ^ s_csamul_cla32_fa26_8_xor1;
  assign s_csamul_cla32_fa25_9_and0 = s_csamul_cla32_and25_9 & s_csamul_cla32_fa26_8_xor1;
  assign s_csamul_cla32_fa25_9_xor1 = s_csamul_cla32_fa25_9_xor0 ^ s_csamul_cla32_fa25_8_or0;
  assign s_csamul_cla32_fa25_9_and1 = s_csamul_cla32_fa25_9_xor0 & s_csamul_cla32_fa25_8_or0;
  assign s_csamul_cla32_fa25_9_or0 = s_csamul_cla32_fa25_9_and0 | s_csamul_cla32_fa25_9_and1;
  assign s_csamul_cla32_and26_9 = a[26] & b[9];
  assign s_csamul_cla32_fa26_9_xor0 = s_csamul_cla32_and26_9 ^ s_csamul_cla32_fa27_8_xor1;
  assign s_csamul_cla32_fa26_9_and0 = s_csamul_cla32_and26_9 & s_csamul_cla32_fa27_8_xor1;
  assign s_csamul_cla32_fa26_9_xor1 = s_csamul_cla32_fa26_9_xor0 ^ s_csamul_cla32_fa26_8_or0;
  assign s_csamul_cla32_fa26_9_and1 = s_csamul_cla32_fa26_9_xor0 & s_csamul_cla32_fa26_8_or0;
  assign s_csamul_cla32_fa26_9_or0 = s_csamul_cla32_fa26_9_and0 | s_csamul_cla32_fa26_9_and1;
  assign s_csamul_cla32_and27_9 = a[27] & b[9];
  assign s_csamul_cla32_fa27_9_xor0 = s_csamul_cla32_and27_9 ^ s_csamul_cla32_fa28_8_xor1;
  assign s_csamul_cla32_fa27_9_and0 = s_csamul_cla32_and27_9 & s_csamul_cla32_fa28_8_xor1;
  assign s_csamul_cla32_fa27_9_xor1 = s_csamul_cla32_fa27_9_xor0 ^ s_csamul_cla32_fa27_8_or0;
  assign s_csamul_cla32_fa27_9_and1 = s_csamul_cla32_fa27_9_xor0 & s_csamul_cla32_fa27_8_or0;
  assign s_csamul_cla32_fa27_9_or0 = s_csamul_cla32_fa27_9_and0 | s_csamul_cla32_fa27_9_and1;
  assign s_csamul_cla32_and28_9 = a[28] & b[9];
  assign s_csamul_cla32_fa28_9_xor0 = s_csamul_cla32_and28_9 ^ s_csamul_cla32_fa29_8_xor1;
  assign s_csamul_cla32_fa28_9_and0 = s_csamul_cla32_and28_9 & s_csamul_cla32_fa29_8_xor1;
  assign s_csamul_cla32_fa28_9_xor1 = s_csamul_cla32_fa28_9_xor0 ^ s_csamul_cla32_fa28_8_or0;
  assign s_csamul_cla32_fa28_9_and1 = s_csamul_cla32_fa28_9_xor0 & s_csamul_cla32_fa28_8_or0;
  assign s_csamul_cla32_fa28_9_or0 = s_csamul_cla32_fa28_9_and0 | s_csamul_cla32_fa28_9_and1;
  assign s_csamul_cla32_and29_9 = a[29] & b[9];
  assign s_csamul_cla32_fa29_9_xor0 = s_csamul_cla32_and29_9 ^ s_csamul_cla32_fa30_8_xor1;
  assign s_csamul_cla32_fa29_9_and0 = s_csamul_cla32_and29_9 & s_csamul_cla32_fa30_8_xor1;
  assign s_csamul_cla32_fa29_9_xor1 = s_csamul_cla32_fa29_9_xor0 ^ s_csamul_cla32_fa29_8_or0;
  assign s_csamul_cla32_fa29_9_and1 = s_csamul_cla32_fa29_9_xor0 & s_csamul_cla32_fa29_8_or0;
  assign s_csamul_cla32_fa29_9_or0 = s_csamul_cla32_fa29_9_and0 | s_csamul_cla32_fa29_9_and1;
  assign s_csamul_cla32_and30_9 = a[30] & b[9];
  assign s_csamul_cla32_fa30_9_xor0 = s_csamul_cla32_and30_9 ^ s_csamul_cla32_ha31_8_xor0;
  assign s_csamul_cla32_fa30_9_and0 = s_csamul_cla32_and30_9 & s_csamul_cla32_ha31_8_xor0;
  assign s_csamul_cla32_fa30_9_xor1 = s_csamul_cla32_fa30_9_xor0 ^ s_csamul_cla32_fa30_8_or0;
  assign s_csamul_cla32_fa30_9_and1 = s_csamul_cla32_fa30_9_xor0 & s_csamul_cla32_fa30_8_or0;
  assign s_csamul_cla32_fa30_9_or0 = s_csamul_cla32_fa30_9_and0 | s_csamul_cla32_fa30_9_and1;
  assign s_csamul_cla32_nand31_9 = ~(a[31] & b[9]);
  assign s_csamul_cla32_ha31_9_xor0 = s_csamul_cla32_nand31_9 ^ s_csamul_cla32_ha31_8_and0;
  assign s_csamul_cla32_ha31_9_and0 = s_csamul_cla32_nand31_9 & s_csamul_cla32_ha31_8_and0;
  assign s_csamul_cla32_and0_10 = a[0] & b[10];
  assign s_csamul_cla32_fa0_10_xor0 = s_csamul_cla32_and0_10 ^ s_csamul_cla32_fa1_9_xor1;
  assign s_csamul_cla32_fa0_10_and0 = s_csamul_cla32_and0_10 & s_csamul_cla32_fa1_9_xor1;
  assign s_csamul_cla32_fa0_10_xor1 = s_csamul_cla32_fa0_10_xor0 ^ s_csamul_cla32_fa0_9_or0;
  assign s_csamul_cla32_fa0_10_and1 = s_csamul_cla32_fa0_10_xor0 & s_csamul_cla32_fa0_9_or0;
  assign s_csamul_cla32_fa0_10_or0 = s_csamul_cla32_fa0_10_and0 | s_csamul_cla32_fa0_10_and1;
  assign s_csamul_cla32_and1_10 = a[1] & b[10];
  assign s_csamul_cla32_fa1_10_xor0 = s_csamul_cla32_and1_10 ^ s_csamul_cla32_fa2_9_xor1;
  assign s_csamul_cla32_fa1_10_and0 = s_csamul_cla32_and1_10 & s_csamul_cla32_fa2_9_xor1;
  assign s_csamul_cla32_fa1_10_xor1 = s_csamul_cla32_fa1_10_xor0 ^ s_csamul_cla32_fa1_9_or0;
  assign s_csamul_cla32_fa1_10_and1 = s_csamul_cla32_fa1_10_xor0 & s_csamul_cla32_fa1_9_or0;
  assign s_csamul_cla32_fa1_10_or0 = s_csamul_cla32_fa1_10_and0 | s_csamul_cla32_fa1_10_and1;
  assign s_csamul_cla32_and2_10 = a[2] & b[10];
  assign s_csamul_cla32_fa2_10_xor0 = s_csamul_cla32_and2_10 ^ s_csamul_cla32_fa3_9_xor1;
  assign s_csamul_cla32_fa2_10_and0 = s_csamul_cla32_and2_10 & s_csamul_cla32_fa3_9_xor1;
  assign s_csamul_cla32_fa2_10_xor1 = s_csamul_cla32_fa2_10_xor0 ^ s_csamul_cla32_fa2_9_or0;
  assign s_csamul_cla32_fa2_10_and1 = s_csamul_cla32_fa2_10_xor0 & s_csamul_cla32_fa2_9_or0;
  assign s_csamul_cla32_fa2_10_or0 = s_csamul_cla32_fa2_10_and0 | s_csamul_cla32_fa2_10_and1;
  assign s_csamul_cla32_and3_10 = a[3] & b[10];
  assign s_csamul_cla32_fa3_10_xor0 = s_csamul_cla32_and3_10 ^ s_csamul_cla32_fa4_9_xor1;
  assign s_csamul_cla32_fa3_10_and0 = s_csamul_cla32_and3_10 & s_csamul_cla32_fa4_9_xor1;
  assign s_csamul_cla32_fa3_10_xor1 = s_csamul_cla32_fa3_10_xor0 ^ s_csamul_cla32_fa3_9_or0;
  assign s_csamul_cla32_fa3_10_and1 = s_csamul_cla32_fa3_10_xor0 & s_csamul_cla32_fa3_9_or0;
  assign s_csamul_cla32_fa3_10_or0 = s_csamul_cla32_fa3_10_and0 | s_csamul_cla32_fa3_10_and1;
  assign s_csamul_cla32_and4_10 = a[4] & b[10];
  assign s_csamul_cla32_fa4_10_xor0 = s_csamul_cla32_and4_10 ^ s_csamul_cla32_fa5_9_xor1;
  assign s_csamul_cla32_fa4_10_and0 = s_csamul_cla32_and4_10 & s_csamul_cla32_fa5_9_xor1;
  assign s_csamul_cla32_fa4_10_xor1 = s_csamul_cla32_fa4_10_xor0 ^ s_csamul_cla32_fa4_9_or0;
  assign s_csamul_cla32_fa4_10_and1 = s_csamul_cla32_fa4_10_xor0 & s_csamul_cla32_fa4_9_or0;
  assign s_csamul_cla32_fa4_10_or0 = s_csamul_cla32_fa4_10_and0 | s_csamul_cla32_fa4_10_and1;
  assign s_csamul_cla32_and5_10 = a[5] & b[10];
  assign s_csamul_cla32_fa5_10_xor0 = s_csamul_cla32_and5_10 ^ s_csamul_cla32_fa6_9_xor1;
  assign s_csamul_cla32_fa5_10_and0 = s_csamul_cla32_and5_10 & s_csamul_cla32_fa6_9_xor1;
  assign s_csamul_cla32_fa5_10_xor1 = s_csamul_cla32_fa5_10_xor0 ^ s_csamul_cla32_fa5_9_or0;
  assign s_csamul_cla32_fa5_10_and1 = s_csamul_cla32_fa5_10_xor0 & s_csamul_cla32_fa5_9_or0;
  assign s_csamul_cla32_fa5_10_or0 = s_csamul_cla32_fa5_10_and0 | s_csamul_cla32_fa5_10_and1;
  assign s_csamul_cla32_and6_10 = a[6] & b[10];
  assign s_csamul_cla32_fa6_10_xor0 = s_csamul_cla32_and6_10 ^ s_csamul_cla32_fa7_9_xor1;
  assign s_csamul_cla32_fa6_10_and0 = s_csamul_cla32_and6_10 & s_csamul_cla32_fa7_9_xor1;
  assign s_csamul_cla32_fa6_10_xor1 = s_csamul_cla32_fa6_10_xor0 ^ s_csamul_cla32_fa6_9_or0;
  assign s_csamul_cla32_fa6_10_and1 = s_csamul_cla32_fa6_10_xor0 & s_csamul_cla32_fa6_9_or0;
  assign s_csamul_cla32_fa6_10_or0 = s_csamul_cla32_fa6_10_and0 | s_csamul_cla32_fa6_10_and1;
  assign s_csamul_cla32_and7_10 = a[7] & b[10];
  assign s_csamul_cla32_fa7_10_xor0 = s_csamul_cla32_and7_10 ^ s_csamul_cla32_fa8_9_xor1;
  assign s_csamul_cla32_fa7_10_and0 = s_csamul_cla32_and7_10 & s_csamul_cla32_fa8_9_xor1;
  assign s_csamul_cla32_fa7_10_xor1 = s_csamul_cla32_fa7_10_xor0 ^ s_csamul_cla32_fa7_9_or0;
  assign s_csamul_cla32_fa7_10_and1 = s_csamul_cla32_fa7_10_xor0 & s_csamul_cla32_fa7_9_or0;
  assign s_csamul_cla32_fa7_10_or0 = s_csamul_cla32_fa7_10_and0 | s_csamul_cla32_fa7_10_and1;
  assign s_csamul_cla32_and8_10 = a[8] & b[10];
  assign s_csamul_cla32_fa8_10_xor0 = s_csamul_cla32_and8_10 ^ s_csamul_cla32_fa9_9_xor1;
  assign s_csamul_cla32_fa8_10_and0 = s_csamul_cla32_and8_10 & s_csamul_cla32_fa9_9_xor1;
  assign s_csamul_cla32_fa8_10_xor1 = s_csamul_cla32_fa8_10_xor0 ^ s_csamul_cla32_fa8_9_or0;
  assign s_csamul_cla32_fa8_10_and1 = s_csamul_cla32_fa8_10_xor0 & s_csamul_cla32_fa8_9_or0;
  assign s_csamul_cla32_fa8_10_or0 = s_csamul_cla32_fa8_10_and0 | s_csamul_cla32_fa8_10_and1;
  assign s_csamul_cla32_and9_10 = a[9] & b[10];
  assign s_csamul_cla32_fa9_10_xor0 = s_csamul_cla32_and9_10 ^ s_csamul_cla32_fa10_9_xor1;
  assign s_csamul_cla32_fa9_10_and0 = s_csamul_cla32_and9_10 & s_csamul_cla32_fa10_9_xor1;
  assign s_csamul_cla32_fa9_10_xor1 = s_csamul_cla32_fa9_10_xor0 ^ s_csamul_cla32_fa9_9_or0;
  assign s_csamul_cla32_fa9_10_and1 = s_csamul_cla32_fa9_10_xor0 & s_csamul_cla32_fa9_9_or0;
  assign s_csamul_cla32_fa9_10_or0 = s_csamul_cla32_fa9_10_and0 | s_csamul_cla32_fa9_10_and1;
  assign s_csamul_cla32_and10_10 = a[10] & b[10];
  assign s_csamul_cla32_fa10_10_xor0 = s_csamul_cla32_and10_10 ^ s_csamul_cla32_fa11_9_xor1;
  assign s_csamul_cla32_fa10_10_and0 = s_csamul_cla32_and10_10 & s_csamul_cla32_fa11_9_xor1;
  assign s_csamul_cla32_fa10_10_xor1 = s_csamul_cla32_fa10_10_xor0 ^ s_csamul_cla32_fa10_9_or0;
  assign s_csamul_cla32_fa10_10_and1 = s_csamul_cla32_fa10_10_xor0 & s_csamul_cla32_fa10_9_or0;
  assign s_csamul_cla32_fa10_10_or0 = s_csamul_cla32_fa10_10_and0 | s_csamul_cla32_fa10_10_and1;
  assign s_csamul_cla32_and11_10 = a[11] & b[10];
  assign s_csamul_cla32_fa11_10_xor0 = s_csamul_cla32_and11_10 ^ s_csamul_cla32_fa12_9_xor1;
  assign s_csamul_cla32_fa11_10_and0 = s_csamul_cla32_and11_10 & s_csamul_cla32_fa12_9_xor1;
  assign s_csamul_cla32_fa11_10_xor1 = s_csamul_cla32_fa11_10_xor0 ^ s_csamul_cla32_fa11_9_or0;
  assign s_csamul_cla32_fa11_10_and1 = s_csamul_cla32_fa11_10_xor0 & s_csamul_cla32_fa11_9_or0;
  assign s_csamul_cla32_fa11_10_or0 = s_csamul_cla32_fa11_10_and0 | s_csamul_cla32_fa11_10_and1;
  assign s_csamul_cla32_and12_10 = a[12] & b[10];
  assign s_csamul_cla32_fa12_10_xor0 = s_csamul_cla32_and12_10 ^ s_csamul_cla32_fa13_9_xor1;
  assign s_csamul_cla32_fa12_10_and0 = s_csamul_cla32_and12_10 & s_csamul_cla32_fa13_9_xor1;
  assign s_csamul_cla32_fa12_10_xor1 = s_csamul_cla32_fa12_10_xor0 ^ s_csamul_cla32_fa12_9_or0;
  assign s_csamul_cla32_fa12_10_and1 = s_csamul_cla32_fa12_10_xor0 & s_csamul_cla32_fa12_9_or0;
  assign s_csamul_cla32_fa12_10_or0 = s_csamul_cla32_fa12_10_and0 | s_csamul_cla32_fa12_10_and1;
  assign s_csamul_cla32_and13_10 = a[13] & b[10];
  assign s_csamul_cla32_fa13_10_xor0 = s_csamul_cla32_and13_10 ^ s_csamul_cla32_fa14_9_xor1;
  assign s_csamul_cla32_fa13_10_and0 = s_csamul_cla32_and13_10 & s_csamul_cla32_fa14_9_xor1;
  assign s_csamul_cla32_fa13_10_xor1 = s_csamul_cla32_fa13_10_xor0 ^ s_csamul_cla32_fa13_9_or0;
  assign s_csamul_cla32_fa13_10_and1 = s_csamul_cla32_fa13_10_xor0 & s_csamul_cla32_fa13_9_or0;
  assign s_csamul_cla32_fa13_10_or0 = s_csamul_cla32_fa13_10_and0 | s_csamul_cla32_fa13_10_and1;
  assign s_csamul_cla32_and14_10 = a[14] & b[10];
  assign s_csamul_cla32_fa14_10_xor0 = s_csamul_cla32_and14_10 ^ s_csamul_cla32_fa15_9_xor1;
  assign s_csamul_cla32_fa14_10_and0 = s_csamul_cla32_and14_10 & s_csamul_cla32_fa15_9_xor1;
  assign s_csamul_cla32_fa14_10_xor1 = s_csamul_cla32_fa14_10_xor0 ^ s_csamul_cla32_fa14_9_or0;
  assign s_csamul_cla32_fa14_10_and1 = s_csamul_cla32_fa14_10_xor0 & s_csamul_cla32_fa14_9_or0;
  assign s_csamul_cla32_fa14_10_or0 = s_csamul_cla32_fa14_10_and0 | s_csamul_cla32_fa14_10_and1;
  assign s_csamul_cla32_and15_10 = a[15] & b[10];
  assign s_csamul_cla32_fa15_10_xor0 = s_csamul_cla32_and15_10 ^ s_csamul_cla32_fa16_9_xor1;
  assign s_csamul_cla32_fa15_10_and0 = s_csamul_cla32_and15_10 & s_csamul_cla32_fa16_9_xor1;
  assign s_csamul_cla32_fa15_10_xor1 = s_csamul_cla32_fa15_10_xor0 ^ s_csamul_cla32_fa15_9_or0;
  assign s_csamul_cla32_fa15_10_and1 = s_csamul_cla32_fa15_10_xor0 & s_csamul_cla32_fa15_9_or0;
  assign s_csamul_cla32_fa15_10_or0 = s_csamul_cla32_fa15_10_and0 | s_csamul_cla32_fa15_10_and1;
  assign s_csamul_cla32_and16_10 = a[16] & b[10];
  assign s_csamul_cla32_fa16_10_xor0 = s_csamul_cla32_and16_10 ^ s_csamul_cla32_fa17_9_xor1;
  assign s_csamul_cla32_fa16_10_and0 = s_csamul_cla32_and16_10 & s_csamul_cla32_fa17_9_xor1;
  assign s_csamul_cla32_fa16_10_xor1 = s_csamul_cla32_fa16_10_xor0 ^ s_csamul_cla32_fa16_9_or0;
  assign s_csamul_cla32_fa16_10_and1 = s_csamul_cla32_fa16_10_xor0 & s_csamul_cla32_fa16_9_or0;
  assign s_csamul_cla32_fa16_10_or0 = s_csamul_cla32_fa16_10_and0 | s_csamul_cla32_fa16_10_and1;
  assign s_csamul_cla32_and17_10 = a[17] & b[10];
  assign s_csamul_cla32_fa17_10_xor0 = s_csamul_cla32_and17_10 ^ s_csamul_cla32_fa18_9_xor1;
  assign s_csamul_cla32_fa17_10_and0 = s_csamul_cla32_and17_10 & s_csamul_cla32_fa18_9_xor1;
  assign s_csamul_cla32_fa17_10_xor1 = s_csamul_cla32_fa17_10_xor0 ^ s_csamul_cla32_fa17_9_or0;
  assign s_csamul_cla32_fa17_10_and1 = s_csamul_cla32_fa17_10_xor0 & s_csamul_cla32_fa17_9_or0;
  assign s_csamul_cla32_fa17_10_or0 = s_csamul_cla32_fa17_10_and0 | s_csamul_cla32_fa17_10_and1;
  assign s_csamul_cla32_and18_10 = a[18] & b[10];
  assign s_csamul_cla32_fa18_10_xor0 = s_csamul_cla32_and18_10 ^ s_csamul_cla32_fa19_9_xor1;
  assign s_csamul_cla32_fa18_10_and0 = s_csamul_cla32_and18_10 & s_csamul_cla32_fa19_9_xor1;
  assign s_csamul_cla32_fa18_10_xor1 = s_csamul_cla32_fa18_10_xor0 ^ s_csamul_cla32_fa18_9_or0;
  assign s_csamul_cla32_fa18_10_and1 = s_csamul_cla32_fa18_10_xor0 & s_csamul_cla32_fa18_9_or0;
  assign s_csamul_cla32_fa18_10_or0 = s_csamul_cla32_fa18_10_and0 | s_csamul_cla32_fa18_10_and1;
  assign s_csamul_cla32_and19_10 = a[19] & b[10];
  assign s_csamul_cla32_fa19_10_xor0 = s_csamul_cla32_and19_10 ^ s_csamul_cla32_fa20_9_xor1;
  assign s_csamul_cla32_fa19_10_and0 = s_csamul_cla32_and19_10 & s_csamul_cla32_fa20_9_xor1;
  assign s_csamul_cla32_fa19_10_xor1 = s_csamul_cla32_fa19_10_xor0 ^ s_csamul_cla32_fa19_9_or0;
  assign s_csamul_cla32_fa19_10_and1 = s_csamul_cla32_fa19_10_xor0 & s_csamul_cla32_fa19_9_or0;
  assign s_csamul_cla32_fa19_10_or0 = s_csamul_cla32_fa19_10_and0 | s_csamul_cla32_fa19_10_and1;
  assign s_csamul_cla32_and20_10 = a[20] & b[10];
  assign s_csamul_cla32_fa20_10_xor0 = s_csamul_cla32_and20_10 ^ s_csamul_cla32_fa21_9_xor1;
  assign s_csamul_cla32_fa20_10_and0 = s_csamul_cla32_and20_10 & s_csamul_cla32_fa21_9_xor1;
  assign s_csamul_cla32_fa20_10_xor1 = s_csamul_cla32_fa20_10_xor0 ^ s_csamul_cla32_fa20_9_or0;
  assign s_csamul_cla32_fa20_10_and1 = s_csamul_cla32_fa20_10_xor0 & s_csamul_cla32_fa20_9_or0;
  assign s_csamul_cla32_fa20_10_or0 = s_csamul_cla32_fa20_10_and0 | s_csamul_cla32_fa20_10_and1;
  assign s_csamul_cla32_and21_10 = a[21] & b[10];
  assign s_csamul_cla32_fa21_10_xor0 = s_csamul_cla32_and21_10 ^ s_csamul_cla32_fa22_9_xor1;
  assign s_csamul_cla32_fa21_10_and0 = s_csamul_cla32_and21_10 & s_csamul_cla32_fa22_9_xor1;
  assign s_csamul_cla32_fa21_10_xor1 = s_csamul_cla32_fa21_10_xor0 ^ s_csamul_cla32_fa21_9_or0;
  assign s_csamul_cla32_fa21_10_and1 = s_csamul_cla32_fa21_10_xor0 & s_csamul_cla32_fa21_9_or0;
  assign s_csamul_cla32_fa21_10_or0 = s_csamul_cla32_fa21_10_and0 | s_csamul_cla32_fa21_10_and1;
  assign s_csamul_cla32_and22_10 = a[22] & b[10];
  assign s_csamul_cla32_fa22_10_xor0 = s_csamul_cla32_and22_10 ^ s_csamul_cla32_fa23_9_xor1;
  assign s_csamul_cla32_fa22_10_and0 = s_csamul_cla32_and22_10 & s_csamul_cla32_fa23_9_xor1;
  assign s_csamul_cla32_fa22_10_xor1 = s_csamul_cla32_fa22_10_xor0 ^ s_csamul_cla32_fa22_9_or0;
  assign s_csamul_cla32_fa22_10_and1 = s_csamul_cla32_fa22_10_xor0 & s_csamul_cla32_fa22_9_or0;
  assign s_csamul_cla32_fa22_10_or0 = s_csamul_cla32_fa22_10_and0 | s_csamul_cla32_fa22_10_and1;
  assign s_csamul_cla32_and23_10 = a[23] & b[10];
  assign s_csamul_cla32_fa23_10_xor0 = s_csamul_cla32_and23_10 ^ s_csamul_cla32_fa24_9_xor1;
  assign s_csamul_cla32_fa23_10_and0 = s_csamul_cla32_and23_10 & s_csamul_cla32_fa24_9_xor1;
  assign s_csamul_cla32_fa23_10_xor1 = s_csamul_cla32_fa23_10_xor0 ^ s_csamul_cla32_fa23_9_or0;
  assign s_csamul_cla32_fa23_10_and1 = s_csamul_cla32_fa23_10_xor0 & s_csamul_cla32_fa23_9_or0;
  assign s_csamul_cla32_fa23_10_or0 = s_csamul_cla32_fa23_10_and0 | s_csamul_cla32_fa23_10_and1;
  assign s_csamul_cla32_and24_10 = a[24] & b[10];
  assign s_csamul_cla32_fa24_10_xor0 = s_csamul_cla32_and24_10 ^ s_csamul_cla32_fa25_9_xor1;
  assign s_csamul_cla32_fa24_10_and0 = s_csamul_cla32_and24_10 & s_csamul_cla32_fa25_9_xor1;
  assign s_csamul_cla32_fa24_10_xor1 = s_csamul_cla32_fa24_10_xor0 ^ s_csamul_cla32_fa24_9_or0;
  assign s_csamul_cla32_fa24_10_and1 = s_csamul_cla32_fa24_10_xor0 & s_csamul_cla32_fa24_9_or0;
  assign s_csamul_cla32_fa24_10_or0 = s_csamul_cla32_fa24_10_and0 | s_csamul_cla32_fa24_10_and1;
  assign s_csamul_cla32_and25_10 = a[25] & b[10];
  assign s_csamul_cla32_fa25_10_xor0 = s_csamul_cla32_and25_10 ^ s_csamul_cla32_fa26_9_xor1;
  assign s_csamul_cla32_fa25_10_and0 = s_csamul_cla32_and25_10 & s_csamul_cla32_fa26_9_xor1;
  assign s_csamul_cla32_fa25_10_xor1 = s_csamul_cla32_fa25_10_xor0 ^ s_csamul_cla32_fa25_9_or0;
  assign s_csamul_cla32_fa25_10_and1 = s_csamul_cla32_fa25_10_xor0 & s_csamul_cla32_fa25_9_or0;
  assign s_csamul_cla32_fa25_10_or0 = s_csamul_cla32_fa25_10_and0 | s_csamul_cla32_fa25_10_and1;
  assign s_csamul_cla32_and26_10 = a[26] & b[10];
  assign s_csamul_cla32_fa26_10_xor0 = s_csamul_cla32_and26_10 ^ s_csamul_cla32_fa27_9_xor1;
  assign s_csamul_cla32_fa26_10_and0 = s_csamul_cla32_and26_10 & s_csamul_cla32_fa27_9_xor1;
  assign s_csamul_cla32_fa26_10_xor1 = s_csamul_cla32_fa26_10_xor0 ^ s_csamul_cla32_fa26_9_or0;
  assign s_csamul_cla32_fa26_10_and1 = s_csamul_cla32_fa26_10_xor0 & s_csamul_cla32_fa26_9_or0;
  assign s_csamul_cla32_fa26_10_or0 = s_csamul_cla32_fa26_10_and0 | s_csamul_cla32_fa26_10_and1;
  assign s_csamul_cla32_and27_10 = a[27] & b[10];
  assign s_csamul_cla32_fa27_10_xor0 = s_csamul_cla32_and27_10 ^ s_csamul_cla32_fa28_9_xor1;
  assign s_csamul_cla32_fa27_10_and0 = s_csamul_cla32_and27_10 & s_csamul_cla32_fa28_9_xor1;
  assign s_csamul_cla32_fa27_10_xor1 = s_csamul_cla32_fa27_10_xor0 ^ s_csamul_cla32_fa27_9_or0;
  assign s_csamul_cla32_fa27_10_and1 = s_csamul_cla32_fa27_10_xor0 & s_csamul_cla32_fa27_9_or0;
  assign s_csamul_cla32_fa27_10_or0 = s_csamul_cla32_fa27_10_and0 | s_csamul_cla32_fa27_10_and1;
  assign s_csamul_cla32_and28_10 = a[28] & b[10];
  assign s_csamul_cla32_fa28_10_xor0 = s_csamul_cla32_and28_10 ^ s_csamul_cla32_fa29_9_xor1;
  assign s_csamul_cla32_fa28_10_and0 = s_csamul_cla32_and28_10 & s_csamul_cla32_fa29_9_xor1;
  assign s_csamul_cla32_fa28_10_xor1 = s_csamul_cla32_fa28_10_xor0 ^ s_csamul_cla32_fa28_9_or0;
  assign s_csamul_cla32_fa28_10_and1 = s_csamul_cla32_fa28_10_xor0 & s_csamul_cla32_fa28_9_or0;
  assign s_csamul_cla32_fa28_10_or0 = s_csamul_cla32_fa28_10_and0 | s_csamul_cla32_fa28_10_and1;
  assign s_csamul_cla32_and29_10 = a[29] & b[10];
  assign s_csamul_cla32_fa29_10_xor0 = s_csamul_cla32_and29_10 ^ s_csamul_cla32_fa30_9_xor1;
  assign s_csamul_cla32_fa29_10_and0 = s_csamul_cla32_and29_10 & s_csamul_cla32_fa30_9_xor1;
  assign s_csamul_cla32_fa29_10_xor1 = s_csamul_cla32_fa29_10_xor0 ^ s_csamul_cla32_fa29_9_or0;
  assign s_csamul_cla32_fa29_10_and1 = s_csamul_cla32_fa29_10_xor0 & s_csamul_cla32_fa29_9_or0;
  assign s_csamul_cla32_fa29_10_or0 = s_csamul_cla32_fa29_10_and0 | s_csamul_cla32_fa29_10_and1;
  assign s_csamul_cla32_and30_10 = a[30] & b[10];
  assign s_csamul_cla32_fa30_10_xor0 = s_csamul_cla32_and30_10 ^ s_csamul_cla32_ha31_9_xor0;
  assign s_csamul_cla32_fa30_10_and0 = s_csamul_cla32_and30_10 & s_csamul_cla32_ha31_9_xor0;
  assign s_csamul_cla32_fa30_10_xor1 = s_csamul_cla32_fa30_10_xor0 ^ s_csamul_cla32_fa30_9_or0;
  assign s_csamul_cla32_fa30_10_and1 = s_csamul_cla32_fa30_10_xor0 & s_csamul_cla32_fa30_9_or0;
  assign s_csamul_cla32_fa30_10_or0 = s_csamul_cla32_fa30_10_and0 | s_csamul_cla32_fa30_10_and1;
  assign s_csamul_cla32_nand31_10 = ~(a[31] & b[10]);
  assign s_csamul_cla32_ha31_10_xor0 = s_csamul_cla32_nand31_10 ^ s_csamul_cla32_ha31_9_and0;
  assign s_csamul_cla32_ha31_10_and0 = s_csamul_cla32_nand31_10 & s_csamul_cla32_ha31_9_and0;
  assign s_csamul_cla32_and0_11 = a[0] & b[11];
  assign s_csamul_cla32_fa0_11_xor0 = s_csamul_cla32_and0_11 ^ s_csamul_cla32_fa1_10_xor1;
  assign s_csamul_cla32_fa0_11_and0 = s_csamul_cla32_and0_11 & s_csamul_cla32_fa1_10_xor1;
  assign s_csamul_cla32_fa0_11_xor1 = s_csamul_cla32_fa0_11_xor0 ^ s_csamul_cla32_fa0_10_or0;
  assign s_csamul_cla32_fa0_11_and1 = s_csamul_cla32_fa0_11_xor0 & s_csamul_cla32_fa0_10_or0;
  assign s_csamul_cla32_fa0_11_or0 = s_csamul_cla32_fa0_11_and0 | s_csamul_cla32_fa0_11_and1;
  assign s_csamul_cla32_and1_11 = a[1] & b[11];
  assign s_csamul_cla32_fa1_11_xor0 = s_csamul_cla32_and1_11 ^ s_csamul_cla32_fa2_10_xor1;
  assign s_csamul_cla32_fa1_11_and0 = s_csamul_cla32_and1_11 & s_csamul_cla32_fa2_10_xor1;
  assign s_csamul_cla32_fa1_11_xor1 = s_csamul_cla32_fa1_11_xor0 ^ s_csamul_cla32_fa1_10_or0;
  assign s_csamul_cla32_fa1_11_and1 = s_csamul_cla32_fa1_11_xor0 & s_csamul_cla32_fa1_10_or0;
  assign s_csamul_cla32_fa1_11_or0 = s_csamul_cla32_fa1_11_and0 | s_csamul_cla32_fa1_11_and1;
  assign s_csamul_cla32_and2_11 = a[2] & b[11];
  assign s_csamul_cla32_fa2_11_xor0 = s_csamul_cla32_and2_11 ^ s_csamul_cla32_fa3_10_xor1;
  assign s_csamul_cla32_fa2_11_and0 = s_csamul_cla32_and2_11 & s_csamul_cla32_fa3_10_xor1;
  assign s_csamul_cla32_fa2_11_xor1 = s_csamul_cla32_fa2_11_xor0 ^ s_csamul_cla32_fa2_10_or0;
  assign s_csamul_cla32_fa2_11_and1 = s_csamul_cla32_fa2_11_xor0 & s_csamul_cla32_fa2_10_or0;
  assign s_csamul_cla32_fa2_11_or0 = s_csamul_cla32_fa2_11_and0 | s_csamul_cla32_fa2_11_and1;
  assign s_csamul_cla32_and3_11 = a[3] & b[11];
  assign s_csamul_cla32_fa3_11_xor0 = s_csamul_cla32_and3_11 ^ s_csamul_cla32_fa4_10_xor1;
  assign s_csamul_cla32_fa3_11_and0 = s_csamul_cla32_and3_11 & s_csamul_cla32_fa4_10_xor1;
  assign s_csamul_cla32_fa3_11_xor1 = s_csamul_cla32_fa3_11_xor0 ^ s_csamul_cla32_fa3_10_or0;
  assign s_csamul_cla32_fa3_11_and1 = s_csamul_cla32_fa3_11_xor0 & s_csamul_cla32_fa3_10_or0;
  assign s_csamul_cla32_fa3_11_or0 = s_csamul_cla32_fa3_11_and0 | s_csamul_cla32_fa3_11_and1;
  assign s_csamul_cla32_and4_11 = a[4] & b[11];
  assign s_csamul_cla32_fa4_11_xor0 = s_csamul_cla32_and4_11 ^ s_csamul_cla32_fa5_10_xor1;
  assign s_csamul_cla32_fa4_11_and0 = s_csamul_cla32_and4_11 & s_csamul_cla32_fa5_10_xor1;
  assign s_csamul_cla32_fa4_11_xor1 = s_csamul_cla32_fa4_11_xor0 ^ s_csamul_cla32_fa4_10_or0;
  assign s_csamul_cla32_fa4_11_and1 = s_csamul_cla32_fa4_11_xor0 & s_csamul_cla32_fa4_10_or0;
  assign s_csamul_cla32_fa4_11_or0 = s_csamul_cla32_fa4_11_and0 | s_csamul_cla32_fa4_11_and1;
  assign s_csamul_cla32_and5_11 = a[5] & b[11];
  assign s_csamul_cla32_fa5_11_xor0 = s_csamul_cla32_and5_11 ^ s_csamul_cla32_fa6_10_xor1;
  assign s_csamul_cla32_fa5_11_and0 = s_csamul_cla32_and5_11 & s_csamul_cla32_fa6_10_xor1;
  assign s_csamul_cla32_fa5_11_xor1 = s_csamul_cla32_fa5_11_xor0 ^ s_csamul_cla32_fa5_10_or0;
  assign s_csamul_cla32_fa5_11_and1 = s_csamul_cla32_fa5_11_xor0 & s_csamul_cla32_fa5_10_or0;
  assign s_csamul_cla32_fa5_11_or0 = s_csamul_cla32_fa5_11_and0 | s_csamul_cla32_fa5_11_and1;
  assign s_csamul_cla32_and6_11 = a[6] & b[11];
  assign s_csamul_cla32_fa6_11_xor0 = s_csamul_cla32_and6_11 ^ s_csamul_cla32_fa7_10_xor1;
  assign s_csamul_cla32_fa6_11_and0 = s_csamul_cla32_and6_11 & s_csamul_cla32_fa7_10_xor1;
  assign s_csamul_cla32_fa6_11_xor1 = s_csamul_cla32_fa6_11_xor0 ^ s_csamul_cla32_fa6_10_or0;
  assign s_csamul_cla32_fa6_11_and1 = s_csamul_cla32_fa6_11_xor0 & s_csamul_cla32_fa6_10_or0;
  assign s_csamul_cla32_fa6_11_or0 = s_csamul_cla32_fa6_11_and0 | s_csamul_cla32_fa6_11_and1;
  assign s_csamul_cla32_and7_11 = a[7] & b[11];
  assign s_csamul_cla32_fa7_11_xor0 = s_csamul_cla32_and7_11 ^ s_csamul_cla32_fa8_10_xor1;
  assign s_csamul_cla32_fa7_11_and0 = s_csamul_cla32_and7_11 & s_csamul_cla32_fa8_10_xor1;
  assign s_csamul_cla32_fa7_11_xor1 = s_csamul_cla32_fa7_11_xor0 ^ s_csamul_cla32_fa7_10_or0;
  assign s_csamul_cla32_fa7_11_and1 = s_csamul_cla32_fa7_11_xor0 & s_csamul_cla32_fa7_10_or0;
  assign s_csamul_cla32_fa7_11_or0 = s_csamul_cla32_fa7_11_and0 | s_csamul_cla32_fa7_11_and1;
  assign s_csamul_cla32_and8_11 = a[8] & b[11];
  assign s_csamul_cla32_fa8_11_xor0 = s_csamul_cla32_and8_11 ^ s_csamul_cla32_fa9_10_xor1;
  assign s_csamul_cla32_fa8_11_and0 = s_csamul_cla32_and8_11 & s_csamul_cla32_fa9_10_xor1;
  assign s_csamul_cla32_fa8_11_xor1 = s_csamul_cla32_fa8_11_xor0 ^ s_csamul_cla32_fa8_10_or0;
  assign s_csamul_cla32_fa8_11_and1 = s_csamul_cla32_fa8_11_xor0 & s_csamul_cla32_fa8_10_or0;
  assign s_csamul_cla32_fa8_11_or0 = s_csamul_cla32_fa8_11_and0 | s_csamul_cla32_fa8_11_and1;
  assign s_csamul_cla32_and9_11 = a[9] & b[11];
  assign s_csamul_cla32_fa9_11_xor0 = s_csamul_cla32_and9_11 ^ s_csamul_cla32_fa10_10_xor1;
  assign s_csamul_cla32_fa9_11_and0 = s_csamul_cla32_and9_11 & s_csamul_cla32_fa10_10_xor1;
  assign s_csamul_cla32_fa9_11_xor1 = s_csamul_cla32_fa9_11_xor0 ^ s_csamul_cla32_fa9_10_or0;
  assign s_csamul_cla32_fa9_11_and1 = s_csamul_cla32_fa9_11_xor0 & s_csamul_cla32_fa9_10_or0;
  assign s_csamul_cla32_fa9_11_or0 = s_csamul_cla32_fa9_11_and0 | s_csamul_cla32_fa9_11_and1;
  assign s_csamul_cla32_and10_11 = a[10] & b[11];
  assign s_csamul_cla32_fa10_11_xor0 = s_csamul_cla32_and10_11 ^ s_csamul_cla32_fa11_10_xor1;
  assign s_csamul_cla32_fa10_11_and0 = s_csamul_cla32_and10_11 & s_csamul_cla32_fa11_10_xor1;
  assign s_csamul_cla32_fa10_11_xor1 = s_csamul_cla32_fa10_11_xor0 ^ s_csamul_cla32_fa10_10_or0;
  assign s_csamul_cla32_fa10_11_and1 = s_csamul_cla32_fa10_11_xor0 & s_csamul_cla32_fa10_10_or0;
  assign s_csamul_cla32_fa10_11_or0 = s_csamul_cla32_fa10_11_and0 | s_csamul_cla32_fa10_11_and1;
  assign s_csamul_cla32_and11_11 = a[11] & b[11];
  assign s_csamul_cla32_fa11_11_xor0 = s_csamul_cla32_and11_11 ^ s_csamul_cla32_fa12_10_xor1;
  assign s_csamul_cla32_fa11_11_and0 = s_csamul_cla32_and11_11 & s_csamul_cla32_fa12_10_xor1;
  assign s_csamul_cla32_fa11_11_xor1 = s_csamul_cla32_fa11_11_xor0 ^ s_csamul_cla32_fa11_10_or0;
  assign s_csamul_cla32_fa11_11_and1 = s_csamul_cla32_fa11_11_xor0 & s_csamul_cla32_fa11_10_or0;
  assign s_csamul_cla32_fa11_11_or0 = s_csamul_cla32_fa11_11_and0 | s_csamul_cla32_fa11_11_and1;
  assign s_csamul_cla32_and12_11 = a[12] & b[11];
  assign s_csamul_cla32_fa12_11_xor0 = s_csamul_cla32_and12_11 ^ s_csamul_cla32_fa13_10_xor1;
  assign s_csamul_cla32_fa12_11_and0 = s_csamul_cla32_and12_11 & s_csamul_cla32_fa13_10_xor1;
  assign s_csamul_cla32_fa12_11_xor1 = s_csamul_cla32_fa12_11_xor0 ^ s_csamul_cla32_fa12_10_or0;
  assign s_csamul_cla32_fa12_11_and1 = s_csamul_cla32_fa12_11_xor0 & s_csamul_cla32_fa12_10_or0;
  assign s_csamul_cla32_fa12_11_or0 = s_csamul_cla32_fa12_11_and0 | s_csamul_cla32_fa12_11_and1;
  assign s_csamul_cla32_and13_11 = a[13] & b[11];
  assign s_csamul_cla32_fa13_11_xor0 = s_csamul_cla32_and13_11 ^ s_csamul_cla32_fa14_10_xor1;
  assign s_csamul_cla32_fa13_11_and0 = s_csamul_cla32_and13_11 & s_csamul_cla32_fa14_10_xor1;
  assign s_csamul_cla32_fa13_11_xor1 = s_csamul_cla32_fa13_11_xor0 ^ s_csamul_cla32_fa13_10_or0;
  assign s_csamul_cla32_fa13_11_and1 = s_csamul_cla32_fa13_11_xor0 & s_csamul_cla32_fa13_10_or0;
  assign s_csamul_cla32_fa13_11_or0 = s_csamul_cla32_fa13_11_and0 | s_csamul_cla32_fa13_11_and1;
  assign s_csamul_cla32_and14_11 = a[14] & b[11];
  assign s_csamul_cla32_fa14_11_xor0 = s_csamul_cla32_and14_11 ^ s_csamul_cla32_fa15_10_xor1;
  assign s_csamul_cla32_fa14_11_and0 = s_csamul_cla32_and14_11 & s_csamul_cla32_fa15_10_xor1;
  assign s_csamul_cla32_fa14_11_xor1 = s_csamul_cla32_fa14_11_xor0 ^ s_csamul_cla32_fa14_10_or0;
  assign s_csamul_cla32_fa14_11_and1 = s_csamul_cla32_fa14_11_xor0 & s_csamul_cla32_fa14_10_or0;
  assign s_csamul_cla32_fa14_11_or0 = s_csamul_cla32_fa14_11_and0 | s_csamul_cla32_fa14_11_and1;
  assign s_csamul_cla32_and15_11 = a[15] & b[11];
  assign s_csamul_cla32_fa15_11_xor0 = s_csamul_cla32_and15_11 ^ s_csamul_cla32_fa16_10_xor1;
  assign s_csamul_cla32_fa15_11_and0 = s_csamul_cla32_and15_11 & s_csamul_cla32_fa16_10_xor1;
  assign s_csamul_cla32_fa15_11_xor1 = s_csamul_cla32_fa15_11_xor0 ^ s_csamul_cla32_fa15_10_or0;
  assign s_csamul_cla32_fa15_11_and1 = s_csamul_cla32_fa15_11_xor0 & s_csamul_cla32_fa15_10_or0;
  assign s_csamul_cla32_fa15_11_or0 = s_csamul_cla32_fa15_11_and0 | s_csamul_cla32_fa15_11_and1;
  assign s_csamul_cla32_and16_11 = a[16] & b[11];
  assign s_csamul_cla32_fa16_11_xor0 = s_csamul_cla32_and16_11 ^ s_csamul_cla32_fa17_10_xor1;
  assign s_csamul_cla32_fa16_11_and0 = s_csamul_cla32_and16_11 & s_csamul_cla32_fa17_10_xor1;
  assign s_csamul_cla32_fa16_11_xor1 = s_csamul_cla32_fa16_11_xor0 ^ s_csamul_cla32_fa16_10_or0;
  assign s_csamul_cla32_fa16_11_and1 = s_csamul_cla32_fa16_11_xor0 & s_csamul_cla32_fa16_10_or0;
  assign s_csamul_cla32_fa16_11_or0 = s_csamul_cla32_fa16_11_and0 | s_csamul_cla32_fa16_11_and1;
  assign s_csamul_cla32_and17_11 = a[17] & b[11];
  assign s_csamul_cla32_fa17_11_xor0 = s_csamul_cla32_and17_11 ^ s_csamul_cla32_fa18_10_xor1;
  assign s_csamul_cla32_fa17_11_and0 = s_csamul_cla32_and17_11 & s_csamul_cla32_fa18_10_xor1;
  assign s_csamul_cla32_fa17_11_xor1 = s_csamul_cla32_fa17_11_xor0 ^ s_csamul_cla32_fa17_10_or0;
  assign s_csamul_cla32_fa17_11_and1 = s_csamul_cla32_fa17_11_xor0 & s_csamul_cla32_fa17_10_or0;
  assign s_csamul_cla32_fa17_11_or0 = s_csamul_cla32_fa17_11_and0 | s_csamul_cla32_fa17_11_and1;
  assign s_csamul_cla32_and18_11 = a[18] & b[11];
  assign s_csamul_cla32_fa18_11_xor0 = s_csamul_cla32_and18_11 ^ s_csamul_cla32_fa19_10_xor1;
  assign s_csamul_cla32_fa18_11_and0 = s_csamul_cla32_and18_11 & s_csamul_cla32_fa19_10_xor1;
  assign s_csamul_cla32_fa18_11_xor1 = s_csamul_cla32_fa18_11_xor0 ^ s_csamul_cla32_fa18_10_or0;
  assign s_csamul_cla32_fa18_11_and1 = s_csamul_cla32_fa18_11_xor0 & s_csamul_cla32_fa18_10_or0;
  assign s_csamul_cla32_fa18_11_or0 = s_csamul_cla32_fa18_11_and0 | s_csamul_cla32_fa18_11_and1;
  assign s_csamul_cla32_and19_11 = a[19] & b[11];
  assign s_csamul_cla32_fa19_11_xor0 = s_csamul_cla32_and19_11 ^ s_csamul_cla32_fa20_10_xor1;
  assign s_csamul_cla32_fa19_11_and0 = s_csamul_cla32_and19_11 & s_csamul_cla32_fa20_10_xor1;
  assign s_csamul_cla32_fa19_11_xor1 = s_csamul_cla32_fa19_11_xor0 ^ s_csamul_cla32_fa19_10_or0;
  assign s_csamul_cla32_fa19_11_and1 = s_csamul_cla32_fa19_11_xor0 & s_csamul_cla32_fa19_10_or0;
  assign s_csamul_cla32_fa19_11_or0 = s_csamul_cla32_fa19_11_and0 | s_csamul_cla32_fa19_11_and1;
  assign s_csamul_cla32_and20_11 = a[20] & b[11];
  assign s_csamul_cla32_fa20_11_xor0 = s_csamul_cla32_and20_11 ^ s_csamul_cla32_fa21_10_xor1;
  assign s_csamul_cla32_fa20_11_and0 = s_csamul_cla32_and20_11 & s_csamul_cla32_fa21_10_xor1;
  assign s_csamul_cla32_fa20_11_xor1 = s_csamul_cla32_fa20_11_xor0 ^ s_csamul_cla32_fa20_10_or0;
  assign s_csamul_cla32_fa20_11_and1 = s_csamul_cla32_fa20_11_xor0 & s_csamul_cla32_fa20_10_or0;
  assign s_csamul_cla32_fa20_11_or0 = s_csamul_cla32_fa20_11_and0 | s_csamul_cla32_fa20_11_and1;
  assign s_csamul_cla32_and21_11 = a[21] & b[11];
  assign s_csamul_cla32_fa21_11_xor0 = s_csamul_cla32_and21_11 ^ s_csamul_cla32_fa22_10_xor1;
  assign s_csamul_cla32_fa21_11_and0 = s_csamul_cla32_and21_11 & s_csamul_cla32_fa22_10_xor1;
  assign s_csamul_cla32_fa21_11_xor1 = s_csamul_cla32_fa21_11_xor0 ^ s_csamul_cla32_fa21_10_or0;
  assign s_csamul_cla32_fa21_11_and1 = s_csamul_cla32_fa21_11_xor0 & s_csamul_cla32_fa21_10_or0;
  assign s_csamul_cla32_fa21_11_or0 = s_csamul_cla32_fa21_11_and0 | s_csamul_cla32_fa21_11_and1;
  assign s_csamul_cla32_and22_11 = a[22] & b[11];
  assign s_csamul_cla32_fa22_11_xor0 = s_csamul_cla32_and22_11 ^ s_csamul_cla32_fa23_10_xor1;
  assign s_csamul_cla32_fa22_11_and0 = s_csamul_cla32_and22_11 & s_csamul_cla32_fa23_10_xor1;
  assign s_csamul_cla32_fa22_11_xor1 = s_csamul_cla32_fa22_11_xor0 ^ s_csamul_cla32_fa22_10_or0;
  assign s_csamul_cla32_fa22_11_and1 = s_csamul_cla32_fa22_11_xor0 & s_csamul_cla32_fa22_10_or0;
  assign s_csamul_cla32_fa22_11_or0 = s_csamul_cla32_fa22_11_and0 | s_csamul_cla32_fa22_11_and1;
  assign s_csamul_cla32_and23_11 = a[23] & b[11];
  assign s_csamul_cla32_fa23_11_xor0 = s_csamul_cla32_and23_11 ^ s_csamul_cla32_fa24_10_xor1;
  assign s_csamul_cla32_fa23_11_and0 = s_csamul_cla32_and23_11 & s_csamul_cla32_fa24_10_xor1;
  assign s_csamul_cla32_fa23_11_xor1 = s_csamul_cla32_fa23_11_xor0 ^ s_csamul_cla32_fa23_10_or0;
  assign s_csamul_cla32_fa23_11_and1 = s_csamul_cla32_fa23_11_xor0 & s_csamul_cla32_fa23_10_or0;
  assign s_csamul_cla32_fa23_11_or0 = s_csamul_cla32_fa23_11_and0 | s_csamul_cla32_fa23_11_and1;
  assign s_csamul_cla32_and24_11 = a[24] & b[11];
  assign s_csamul_cla32_fa24_11_xor0 = s_csamul_cla32_and24_11 ^ s_csamul_cla32_fa25_10_xor1;
  assign s_csamul_cla32_fa24_11_and0 = s_csamul_cla32_and24_11 & s_csamul_cla32_fa25_10_xor1;
  assign s_csamul_cla32_fa24_11_xor1 = s_csamul_cla32_fa24_11_xor0 ^ s_csamul_cla32_fa24_10_or0;
  assign s_csamul_cla32_fa24_11_and1 = s_csamul_cla32_fa24_11_xor0 & s_csamul_cla32_fa24_10_or0;
  assign s_csamul_cla32_fa24_11_or0 = s_csamul_cla32_fa24_11_and0 | s_csamul_cla32_fa24_11_and1;
  assign s_csamul_cla32_and25_11 = a[25] & b[11];
  assign s_csamul_cla32_fa25_11_xor0 = s_csamul_cla32_and25_11 ^ s_csamul_cla32_fa26_10_xor1;
  assign s_csamul_cla32_fa25_11_and0 = s_csamul_cla32_and25_11 & s_csamul_cla32_fa26_10_xor1;
  assign s_csamul_cla32_fa25_11_xor1 = s_csamul_cla32_fa25_11_xor0 ^ s_csamul_cla32_fa25_10_or0;
  assign s_csamul_cla32_fa25_11_and1 = s_csamul_cla32_fa25_11_xor0 & s_csamul_cla32_fa25_10_or0;
  assign s_csamul_cla32_fa25_11_or0 = s_csamul_cla32_fa25_11_and0 | s_csamul_cla32_fa25_11_and1;
  assign s_csamul_cla32_and26_11 = a[26] & b[11];
  assign s_csamul_cla32_fa26_11_xor0 = s_csamul_cla32_and26_11 ^ s_csamul_cla32_fa27_10_xor1;
  assign s_csamul_cla32_fa26_11_and0 = s_csamul_cla32_and26_11 & s_csamul_cla32_fa27_10_xor1;
  assign s_csamul_cla32_fa26_11_xor1 = s_csamul_cla32_fa26_11_xor0 ^ s_csamul_cla32_fa26_10_or0;
  assign s_csamul_cla32_fa26_11_and1 = s_csamul_cla32_fa26_11_xor0 & s_csamul_cla32_fa26_10_or0;
  assign s_csamul_cla32_fa26_11_or0 = s_csamul_cla32_fa26_11_and0 | s_csamul_cla32_fa26_11_and1;
  assign s_csamul_cla32_and27_11 = a[27] & b[11];
  assign s_csamul_cla32_fa27_11_xor0 = s_csamul_cla32_and27_11 ^ s_csamul_cla32_fa28_10_xor1;
  assign s_csamul_cla32_fa27_11_and0 = s_csamul_cla32_and27_11 & s_csamul_cla32_fa28_10_xor1;
  assign s_csamul_cla32_fa27_11_xor1 = s_csamul_cla32_fa27_11_xor0 ^ s_csamul_cla32_fa27_10_or0;
  assign s_csamul_cla32_fa27_11_and1 = s_csamul_cla32_fa27_11_xor0 & s_csamul_cla32_fa27_10_or0;
  assign s_csamul_cla32_fa27_11_or0 = s_csamul_cla32_fa27_11_and0 | s_csamul_cla32_fa27_11_and1;
  assign s_csamul_cla32_and28_11 = a[28] & b[11];
  assign s_csamul_cla32_fa28_11_xor0 = s_csamul_cla32_and28_11 ^ s_csamul_cla32_fa29_10_xor1;
  assign s_csamul_cla32_fa28_11_and0 = s_csamul_cla32_and28_11 & s_csamul_cla32_fa29_10_xor1;
  assign s_csamul_cla32_fa28_11_xor1 = s_csamul_cla32_fa28_11_xor0 ^ s_csamul_cla32_fa28_10_or0;
  assign s_csamul_cla32_fa28_11_and1 = s_csamul_cla32_fa28_11_xor0 & s_csamul_cla32_fa28_10_or0;
  assign s_csamul_cla32_fa28_11_or0 = s_csamul_cla32_fa28_11_and0 | s_csamul_cla32_fa28_11_and1;
  assign s_csamul_cla32_and29_11 = a[29] & b[11];
  assign s_csamul_cla32_fa29_11_xor0 = s_csamul_cla32_and29_11 ^ s_csamul_cla32_fa30_10_xor1;
  assign s_csamul_cla32_fa29_11_and0 = s_csamul_cla32_and29_11 & s_csamul_cla32_fa30_10_xor1;
  assign s_csamul_cla32_fa29_11_xor1 = s_csamul_cla32_fa29_11_xor0 ^ s_csamul_cla32_fa29_10_or0;
  assign s_csamul_cla32_fa29_11_and1 = s_csamul_cla32_fa29_11_xor0 & s_csamul_cla32_fa29_10_or0;
  assign s_csamul_cla32_fa29_11_or0 = s_csamul_cla32_fa29_11_and0 | s_csamul_cla32_fa29_11_and1;
  assign s_csamul_cla32_and30_11 = a[30] & b[11];
  assign s_csamul_cla32_fa30_11_xor0 = s_csamul_cla32_and30_11 ^ s_csamul_cla32_ha31_10_xor0;
  assign s_csamul_cla32_fa30_11_and0 = s_csamul_cla32_and30_11 & s_csamul_cla32_ha31_10_xor0;
  assign s_csamul_cla32_fa30_11_xor1 = s_csamul_cla32_fa30_11_xor0 ^ s_csamul_cla32_fa30_10_or0;
  assign s_csamul_cla32_fa30_11_and1 = s_csamul_cla32_fa30_11_xor0 & s_csamul_cla32_fa30_10_or0;
  assign s_csamul_cla32_fa30_11_or0 = s_csamul_cla32_fa30_11_and0 | s_csamul_cla32_fa30_11_and1;
  assign s_csamul_cla32_nand31_11 = ~(a[31] & b[11]);
  assign s_csamul_cla32_ha31_11_xor0 = s_csamul_cla32_nand31_11 ^ s_csamul_cla32_ha31_10_and0;
  assign s_csamul_cla32_ha31_11_and0 = s_csamul_cla32_nand31_11 & s_csamul_cla32_ha31_10_and0;
  assign s_csamul_cla32_and0_12 = a[0] & b[12];
  assign s_csamul_cla32_fa0_12_xor0 = s_csamul_cla32_and0_12 ^ s_csamul_cla32_fa1_11_xor1;
  assign s_csamul_cla32_fa0_12_and0 = s_csamul_cla32_and0_12 & s_csamul_cla32_fa1_11_xor1;
  assign s_csamul_cla32_fa0_12_xor1 = s_csamul_cla32_fa0_12_xor0 ^ s_csamul_cla32_fa0_11_or0;
  assign s_csamul_cla32_fa0_12_and1 = s_csamul_cla32_fa0_12_xor0 & s_csamul_cla32_fa0_11_or0;
  assign s_csamul_cla32_fa0_12_or0 = s_csamul_cla32_fa0_12_and0 | s_csamul_cla32_fa0_12_and1;
  assign s_csamul_cla32_and1_12 = a[1] & b[12];
  assign s_csamul_cla32_fa1_12_xor0 = s_csamul_cla32_and1_12 ^ s_csamul_cla32_fa2_11_xor1;
  assign s_csamul_cla32_fa1_12_and0 = s_csamul_cla32_and1_12 & s_csamul_cla32_fa2_11_xor1;
  assign s_csamul_cla32_fa1_12_xor1 = s_csamul_cla32_fa1_12_xor0 ^ s_csamul_cla32_fa1_11_or0;
  assign s_csamul_cla32_fa1_12_and1 = s_csamul_cla32_fa1_12_xor0 & s_csamul_cla32_fa1_11_or0;
  assign s_csamul_cla32_fa1_12_or0 = s_csamul_cla32_fa1_12_and0 | s_csamul_cla32_fa1_12_and1;
  assign s_csamul_cla32_and2_12 = a[2] & b[12];
  assign s_csamul_cla32_fa2_12_xor0 = s_csamul_cla32_and2_12 ^ s_csamul_cla32_fa3_11_xor1;
  assign s_csamul_cla32_fa2_12_and0 = s_csamul_cla32_and2_12 & s_csamul_cla32_fa3_11_xor1;
  assign s_csamul_cla32_fa2_12_xor1 = s_csamul_cla32_fa2_12_xor0 ^ s_csamul_cla32_fa2_11_or0;
  assign s_csamul_cla32_fa2_12_and1 = s_csamul_cla32_fa2_12_xor0 & s_csamul_cla32_fa2_11_or0;
  assign s_csamul_cla32_fa2_12_or0 = s_csamul_cla32_fa2_12_and0 | s_csamul_cla32_fa2_12_and1;
  assign s_csamul_cla32_and3_12 = a[3] & b[12];
  assign s_csamul_cla32_fa3_12_xor0 = s_csamul_cla32_and3_12 ^ s_csamul_cla32_fa4_11_xor1;
  assign s_csamul_cla32_fa3_12_and0 = s_csamul_cla32_and3_12 & s_csamul_cla32_fa4_11_xor1;
  assign s_csamul_cla32_fa3_12_xor1 = s_csamul_cla32_fa3_12_xor0 ^ s_csamul_cla32_fa3_11_or0;
  assign s_csamul_cla32_fa3_12_and1 = s_csamul_cla32_fa3_12_xor0 & s_csamul_cla32_fa3_11_or0;
  assign s_csamul_cla32_fa3_12_or0 = s_csamul_cla32_fa3_12_and0 | s_csamul_cla32_fa3_12_and1;
  assign s_csamul_cla32_and4_12 = a[4] & b[12];
  assign s_csamul_cla32_fa4_12_xor0 = s_csamul_cla32_and4_12 ^ s_csamul_cla32_fa5_11_xor1;
  assign s_csamul_cla32_fa4_12_and0 = s_csamul_cla32_and4_12 & s_csamul_cla32_fa5_11_xor1;
  assign s_csamul_cla32_fa4_12_xor1 = s_csamul_cla32_fa4_12_xor0 ^ s_csamul_cla32_fa4_11_or0;
  assign s_csamul_cla32_fa4_12_and1 = s_csamul_cla32_fa4_12_xor0 & s_csamul_cla32_fa4_11_or0;
  assign s_csamul_cla32_fa4_12_or0 = s_csamul_cla32_fa4_12_and0 | s_csamul_cla32_fa4_12_and1;
  assign s_csamul_cla32_and5_12 = a[5] & b[12];
  assign s_csamul_cla32_fa5_12_xor0 = s_csamul_cla32_and5_12 ^ s_csamul_cla32_fa6_11_xor1;
  assign s_csamul_cla32_fa5_12_and0 = s_csamul_cla32_and5_12 & s_csamul_cla32_fa6_11_xor1;
  assign s_csamul_cla32_fa5_12_xor1 = s_csamul_cla32_fa5_12_xor0 ^ s_csamul_cla32_fa5_11_or0;
  assign s_csamul_cla32_fa5_12_and1 = s_csamul_cla32_fa5_12_xor0 & s_csamul_cla32_fa5_11_or0;
  assign s_csamul_cla32_fa5_12_or0 = s_csamul_cla32_fa5_12_and0 | s_csamul_cla32_fa5_12_and1;
  assign s_csamul_cla32_and6_12 = a[6] & b[12];
  assign s_csamul_cla32_fa6_12_xor0 = s_csamul_cla32_and6_12 ^ s_csamul_cla32_fa7_11_xor1;
  assign s_csamul_cla32_fa6_12_and0 = s_csamul_cla32_and6_12 & s_csamul_cla32_fa7_11_xor1;
  assign s_csamul_cla32_fa6_12_xor1 = s_csamul_cla32_fa6_12_xor0 ^ s_csamul_cla32_fa6_11_or0;
  assign s_csamul_cla32_fa6_12_and1 = s_csamul_cla32_fa6_12_xor0 & s_csamul_cla32_fa6_11_or0;
  assign s_csamul_cla32_fa6_12_or0 = s_csamul_cla32_fa6_12_and0 | s_csamul_cla32_fa6_12_and1;
  assign s_csamul_cla32_and7_12 = a[7] & b[12];
  assign s_csamul_cla32_fa7_12_xor0 = s_csamul_cla32_and7_12 ^ s_csamul_cla32_fa8_11_xor1;
  assign s_csamul_cla32_fa7_12_and0 = s_csamul_cla32_and7_12 & s_csamul_cla32_fa8_11_xor1;
  assign s_csamul_cla32_fa7_12_xor1 = s_csamul_cla32_fa7_12_xor0 ^ s_csamul_cla32_fa7_11_or0;
  assign s_csamul_cla32_fa7_12_and1 = s_csamul_cla32_fa7_12_xor0 & s_csamul_cla32_fa7_11_or0;
  assign s_csamul_cla32_fa7_12_or0 = s_csamul_cla32_fa7_12_and0 | s_csamul_cla32_fa7_12_and1;
  assign s_csamul_cla32_and8_12 = a[8] & b[12];
  assign s_csamul_cla32_fa8_12_xor0 = s_csamul_cla32_and8_12 ^ s_csamul_cla32_fa9_11_xor1;
  assign s_csamul_cla32_fa8_12_and0 = s_csamul_cla32_and8_12 & s_csamul_cla32_fa9_11_xor1;
  assign s_csamul_cla32_fa8_12_xor1 = s_csamul_cla32_fa8_12_xor0 ^ s_csamul_cla32_fa8_11_or0;
  assign s_csamul_cla32_fa8_12_and1 = s_csamul_cla32_fa8_12_xor0 & s_csamul_cla32_fa8_11_or0;
  assign s_csamul_cla32_fa8_12_or0 = s_csamul_cla32_fa8_12_and0 | s_csamul_cla32_fa8_12_and1;
  assign s_csamul_cla32_and9_12 = a[9] & b[12];
  assign s_csamul_cla32_fa9_12_xor0 = s_csamul_cla32_and9_12 ^ s_csamul_cla32_fa10_11_xor1;
  assign s_csamul_cla32_fa9_12_and0 = s_csamul_cla32_and9_12 & s_csamul_cla32_fa10_11_xor1;
  assign s_csamul_cla32_fa9_12_xor1 = s_csamul_cla32_fa9_12_xor0 ^ s_csamul_cla32_fa9_11_or0;
  assign s_csamul_cla32_fa9_12_and1 = s_csamul_cla32_fa9_12_xor0 & s_csamul_cla32_fa9_11_or0;
  assign s_csamul_cla32_fa9_12_or0 = s_csamul_cla32_fa9_12_and0 | s_csamul_cla32_fa9_12_and1;
  assign s_csamul_cla32_and10_12 = a[10] & b[12];
  assign s_csamul_cla32_fa10_12_xor0 = s_csamul_cla32_and10_12 ^ s_csamul_cla32_fa11_11_xor1;
  assign s_csamul_cla32_fa10_12_and0 = s_csamul_cla32_and10_12 & s_csamul_cla32_fa11_11_xor1;
  assign s_csamul_cla32_fa10_12_xor1 = s_csamul_cla32_fa10_12_xor0 ^ s_csamul_cla32_fa10_11_or0;
  assign s_csamul_cla32_fa10_12_and1 = s_csamul_cla32_fa10_12_xor0 & s_csamul_cla32_fa10_11_or0;
  assign s_csamul_cla32_fa10_12_or0 = s_csamul_cla32_fa10_12_and0 | s_csamul_cla32_fa10_12_and1;
  assign s_csamul_cla32_and11_12 = a[11] & b[12];
  assign s_csamul_cla32_fa11_12_xor0 = s_csamul_cla32_and11_12 ^ s_csamul_cla32_fa12_11_xor1;
  assign s_csamul_cla32_fa11_12_and0 = s_csamul_cla32_and11_12 & s_csamul_cla32_fa12_11_xor1;
  assign s_csamul_cla32_fa11_12_xor1 = s_csamul_cla32_fa11_12_xor0 ^ s_csamul_cla32_fa11_11_or0;
  assign s_csamul_cla32_fa11_12_and1 = s_csamul_cla32_fa11_12_xor0 & s_csamul_cla32_fa11_11_or0;
  assign s_csamul_cla32_fa11_12_or0 = s_csamul_cla32_fa11_12_and0 | s_csamul_cla32_fa11_12_and1;
  assign s_csamul_cla32_and12_12 = a[12] & b[12];
  assign s_csamul_cla32_fa12_12_xor0 = s_csamul_cla32_and12_12 ^ s_csamul_cla32_fa13_11_xor1;
  assign s_csamul_cla32_fa12_12_and0 = s_csamul_cla32_and12_12 & s_csamul_cla32_fa13_11_xor1;
  assign s_csamul_cla32_fa12_12_xor1 = s_csamul_cla32_fa12_12_xor0 ^ s_csamul_cla32_fa12_11_or0;
  assign s_csamul_cla32_fa12_12_and1 = s_csamul_cla32_fa12_12_xor0 & s_csamul_cla32_fa12_11_or0;
  assign s_csamul_cla32_fa12_12_or0 = s_csamul_cla32_fa12_12_and0 | s_csamul_cla32_fa12_12_and1;
  assign s_csamul_cla32_and13_12 = a[13] & b[12];
  assign s_csamul_cla32_fa13_12_xor0 = s_csamul_cla32_and13_12 ^ s_csamul_cla32_fa14_11_xor1;
  assign s_csamul_cla32_fa13_12_and0 = s_csamul_cla32_and13_12 & s_csamul_cla32_fa14_11_xor1;
  assign s_csamul_cla32_fa13_12_xor1 = s_csamul_cla32_fa13_12_xor0 ^ s_csamul_cla32_fa13_11_or0;
  assign s_csamul_cla32_fa13_12_and1 = s_csamul_cla32_fa13_12_xor0 & s_csamul_cla32_fa13_11_or0;
  assign s_csamul_cla32_fa13_12_or0 = s_csamul_cla32_fa13_12_and0 | s_csamul_cla32_fa13_12_and1;
  assign s_csamul_cla32_and14_12 = a[14] & b[12];
  assign s_csamul_cla32_fa14_12_xor0 = s_csamul_cla32_and14_12 ^ s_csamul_cla32_fa15_11_xor1;
  assign s_csamul_cla32_fa14_12_and0 = s_csamul_cla32_and14_12 & s_csamul_cla32_fa15_11_xor1;
  assign s_csamul_cla32_fa14_12_xor1 = s_csamul_cla32_fa14_12_xor0 ^ s_csamul_cla32_fa14_11_or0;
  assign s_csamul_cla32_fa14_12_and1 = s_csamul_cla32_fa14_12_xor0 & s_csamul_cla32_fa14_11_or0;
  assign s_csamul_cla32_fa14_12_or0 = s_csamul_cla32_fa14_12_and0 | s_csamul_cla32_fa14_12_and1;
  assign s_csamul_cla32_and15_12 = a[15] & b[12];
  assign s_csamul_cla32_fa15_12_xor0 = s_csamul_cla32_and15_12 ^ s_csamul_cla32_fa16_11_xor1;
  assign s_csamul_cla32_fa15_12_and0 = s_csamul_cla32_and15_12 & s_csamul_cla32_fa16_11_xor1;
  assign s_csamul_cla32_fa15_12_xor1 = s_csamul_cla32_fa15_12_xor0 ^ s_csamul_cla32_fa15_11_or0;
  assign s_csamul_cla32_fa15_12_and1 = s_csamul_cla32_fa15_12_xor0 & s_csamul_cla32_fa15_11_or0;
  assign s_csamul_cla32_fa15_12_or0 = s_csamul_cla32_fa15_12_and0 | s_csamul_cla32_fa15_12_and1;
  assign s_csamul_cla32_and16_12 = a[16] & b[12];
  assign s_csamul_cla32_fa16_12_xor0 = s_csamul_cla32_and16_12 ^ s_csamul_cla32_fa17_11_xor1;
  assign s_csamul_cla32_fa16_12_and0 = s_csamul_cla32_and16_12 & s_csamul_cla32_fa17_11_xor1;
  assign s_csamul_cla32_fa16_12_xor1 = s_csamul_cla32_fa16_12_xor0 ^ s_csamul_cla32_fa16_11_or0;
  assign s_csamul_cla32_fa16_12_and1 = s_csamul_cla32_fa16_12_xor0 & s_csamul_cla32_fa16_11_or0;
  assign s_csamul_cla32_fa16_12_or0 = s_csamul_cla32_fa16_12_and0 | s_csamul_cla32_fa16_12_and1;
  assign s_csamul_cla32_and17_12 = a[17] & b[12];
  assign s_csamul_cla32_fa17_12_xor0 = s_csamul_cla32_and17_12 ^ s_csamul_cla32_fa18_11_xor1;
  assign s_csamul_cla32_fa17_12_and0 = s_csamul_cla32_and17_12 & s_csamul_cla32_fa18_11_xor1;
  assign s_csamul_cla32_fa17_12_xor1 = s_csamul_cla32_fa17_12_xor0 ^ s_csamul_cla32_fa17_11_or0;
  assign s_csamul_cla32_fa17_12_and1 = s_csamul_cla32_fa17_12_xor0 & s_csamul_cla32_fa17_11_or0;
  assign s_csamul_cla32_fa17_12_or0 = s_csamul_cla32_fa17_12_and0 | s_csamul_cla32_fa17_12_and1;
  assign s_csamul_cla32_and18_12 = a[18] & b[12];
  assign s_csamul_cla32_fa18_12_xor0 = s_csamul_cla32_and18_12 ^ s_csamul_cla32_fa19_11_xor1;
  assign s_csamul_cla32_fa18_12_and0 = s_csamul_cla32_and18_12 & s_csamul_cla32_fa19_11_xor1;
  assign s_csamul_cla32_fa18_12_xor1 = s_csamul_cla32_fa18_12_xor0 ^ s_csamul_cla32_fa18_11_or0;
  assign s_csamul_cla32_fa18_12_and1 = s_csamul_cla32_fa18_12_xor0 & s_csamul_cla32_fa18_11_or0;
  assign s_csamul_cla32_fa18_12_or0 = s_csamul_cla32_fa18_12_and0 | s_csamul_cla32_fa18_12_and1;
  assign s_csamul_cla32_and19_12 = a[19] & b[12];
  assign s_csamul_cla32_fa19_12_xor0 = s_csamul_cla32_and19_12 ^ s_csamul_cla32_fa20_11_xor1;
  assign s_csamul_cla32_fa19_12_and0 = s_csamul_cla32_and19_12 & s_csamul_cla32_fa20_11_xor1;
  assign s_csamul_cla32_fa19_12_xor1 = s_csamul_cla32_fa19_12_xor0 ^ s_csamul_cla32_fa19_11_or0;
  assign s_csamul_cla32_fa19_12_and1 = s_csamul_cla32_fa19_12_xor0 & s_csamul_cla32_fa19_11_or0;
  assign s_csamul_cla32_fa19_12_or0 = s_csamul_cla32_fa19_12_and0 | s_csamul_cla32_fa19_12_and1;
  assign s_csamul_cla32_and20_12 = a[20] & b[12];
  assign s_csamul_cla32_fa20_12_xor0 = s_csamul_cla32_and20_12 ^ s_csamul_cla32_fa21_11_xor1;
  assign s_csamul_cla32_fa20_12_and0 = s_csamul_cla32_and20_12 & s_csamul_cla32_fa21_11_xor1;
  assign s_csamul_cla32_fa20_12_xor1 = s_csamul_cla32_fa20_12_xor0 ^ s_csamul_cla32_fa20_11_or0;
  assign s_csamul_cla32_fa20_12_and1 = s_csamul_cla32_fa20_12_xor0 & s_csamul_cla32_fa20_11_or0;
  assign s_csamul_cla32_fa20_12_or0 = s_csamul_cla32_fa20_12_and0 | s_csamul_cla32_fa20_12_and1;
  assign s_csamul_cla32_and21_12 = a[21] & b[12];
  assign s_csamul_cla32_fa21_12_xor0 = s_csamul_cla32_and21_12 ^ s_csamul_cla32_fa22_11_xor1;
  assign s_csamul_cla32_fa21_12_and0 = s_csamul_cla32_and21_12 & s_csamul_cla32_fa22_11_xor1;
  assign s_csamul_cla32_fa21_12_xor1 = s_csamul_cla32_fa21_12_xor0 ^ s_csamul_cla32_fa21_11_or0;
  assign s_csamul_cla32_fa21_12_and1 = s_csamul_cla32_fa21_12_xor0 & s_csamul_cla32_fa21_11_or0;
  assign s_csamul_cla32_fa21_12_or0 = s_csamul_cla32_fa21_12_and0 | s_csamul_cla32_fa21_12_and1;
  assign s_csamul_cla32_and22_12 = a[22] & b[12];
  assign s_csamul_cla32_fa22_12_xor0 = s_csamul_cla32_and22_12 ^ s_csamul_cla32_fa23_11_xor1;
  assign s_csamul_cla32_fa22_12_and0 = s_csamul_cla32_and22_12 & s_csamul_cla32_fa23_11_xor1;
  assign s_csamul_cla32_fa22_12_xor1 = s_csamul_cla32_fa22_12_xor0 ^ s_csamul_cla32_fa22_11_or0;
  assign s_csamul_cla32_fa22_12_and1 = s_csamul_cla32_fa22_12_xor0 & s_csamul_cla32_fa22_11_or0;
  assign s_csamul_cla32_fa22_12_or0 = s_csamul_cla32_fa22_12_and0 | s_csamul_cla32_fa22_12_and1;
  assign s_csamul_cla32_and23_12 = a[23] & b[12];
  assign s_csamul_cla32_fa23_12_xor0 = s_csamul_cla32_and23_12 ^ s_csamul_cla32_fa24_11_xor1;
  assign s_csamul_cla32_fa23_12_and0 = s_csamul_cla32_and23_12 & s_csamul_cla32_fa24_11_xor1;
  assign s_csamul_cla32_fa23_12_xor1 = s_csamul_cla32_fa23_12_xor0 ^ s_csamul_cla32_fa23_11_or0;
  assign s_csamul_cla32_fa23_12_and1 = s_csamul_cla32_fa23_12_xor0 & s_csamul_cla32_fa23_11_or0;
  assign s_csamul_cla32_fa23_12_or0 = s_csamul_cla32_fa23_12_and0 | s_csamul_cla32_fa23_12_and1;
  assign s_csamul_cla32_and24_12 = a[24] & b[12];
  assign s_csamul_cla32_fa24_12_xor0 = s_csamul_cla32_and24_12 ^ s_csamul_cla32_fa25_11_xor1;
  assign s_csamul_cla32_fa24_12_and0 = s_csamul_cla32_and24_12 & s_csamul_cla32_fa25_11_xor1;
  assign s_csamul_cla32_fa24_12_xor1 = s_csamul_cla32_fa24_12_xor0 ^ s_csamul_cla32_fa24_11_or0;
  assign s_csamul_cla32_fa24_12_and1 = s_csamul_cla32_fa24_12_xor0 & s_csamul_cla32_fa24_11_or0;
  assign s_csamul_cla32_fa24_12_or0 = s_csamul_cla32_fa24_12_and0 | s_csamul_cla32_fa24_12_and1;
  assign s_csamul_cla32_and25_12 = a[25] & b[12];
  assign s_csamul_cla32_fa25_12_xor0 = s_csamul_cla32_and25_12 ^ s_csamul_cla32_fa26_11_xor1;
  assign s_csamul_cla32_fa25_12_and0 = s_csamul_cla32_and25_12 & s_csamul_cla32_fa26_11_xor1;
  assign s_csamul_cla32_fa25_12_xor1 = s_csamul_cla32_fa25_12_xor0 ^ s_csamul_cla32_fa25_11_or0;
  assign s_csamul_cla32_fa25_12_and1 = s_csamul_cla32_fa25_12_xor0 & s_csamul_cla32_fa25_11_or0;
  assign s_csamul_cla32_fa25_12_or0 = s_csamul_cla32_fa25_12_and0 | s_csamul_cla32_fa25_12_and1;
  assign s_csamul_cla32_and26_12 = a[26] & b[12];
  assign s_csamul_cla32_fa26_12_xor0 = s_csamul_cla32_and26_12 ^ s_csamul_cla32_fa27_11_xor1;
  assign s_csamul_cla32_fa26_12_and0 = s_csamul_cla32_and26_12 & s_csamul_cla32_fa27_11_xor1;
  assign s_csamul_cla32_fa26_12_xor1 = s_csamul_cla32_fa26_12_xor0 ^ s_csamul_cla32_fa26_11_or0;
  assign s_csamul_cla32_fa26_12_and1 = s_csamul_cla32_fa26_12_xor0 & s_csamul_cla32_fa26_11_or0;
  assign s_csamul_cla32_fa26_12_or0 = s_csamul_cla32_fa26_12_and0 | s_csamul_cla32_fa26_12_and1;
  assign s_csamul_cla32_and27_12 = a[27] & b[12];
  assign s_csamul_cla32_fa27_12_xor0 = s_csamul_cla32_and27_12 ^ s_csamul_cla32_fa28_11_xor1;
  assign s_csamul_cla32_fa27_12_and0 = s_csamul_cla32_and27_12 & s_csamul_cla32_fa28_11_xor1;
  assign s_csamul_cla32_fa27_12_xor1 = s_csamul_cla32_fa27_12_xor0 ^ s_csamul_cla32_fa27_11_or0;
  assign s_csamul_cla32_fa27_12_and1 = s_csamul_cla32_fa27_12_xor0 & s_csamul_cla32_fa27_11_or0;
  assign s_csamul_cla32_fa27_12_or0 = s_csamul_cla32_fa27_12_and0 | s_csamul_cla32_fa27_12_and1;
  assign s_csamul_cla32_and28_12 = a[28] & b[12];
  assign s_csamul_cla32_fa28_12_xor0 = s_csamul_cla32_and28_12 ^ s_csamul_cla32_fa29_11_xor1;
  assign s_csamul_cla32_fa28_12_and0 = s_csamul_cla32_and28_12 & s_csamul_cla32_fa29_11_xor1;
  assign s_csamul_cla32_fa28_12_xor1 = s_csamul_cla32_fa28_12_xor0 ^ s_csamul_cla32_fa28_11_or0;
  assign s_csamul_cla32_fa28_12_and1 = s_csamul_cla32_fa28_12_xor0 & s_csamul_cla32_fa28_11_or0;
  assign s_csamul_cla32_fa28_12_or0 = s_csamul_cla32_fa28_12_and0 | s_csamul_cla32_fa28_12_and1;
  assign s_csamul_cla32_and29_12 = a[29] & b[12];
  assign s_csamul_cla32_fa29_12_xor0 = s_csamul_cla32_and29_12 ^ s_csamul_cla32_fa30_11_xor1;
  assign s_csamul_cla32_fa29_12_and0 = s_csamul_cla32_and29_12 & s_csamul_cla32_fa30_11_xor1;
  assign s_csamul_cla32_fa29_12_xor1 = s_csamul_cla32_fa29_12_xor0 ^ s_csamul_cla32_fa29_11_or0;
  assign s_csamul_cla32_fa29_12_and1 = s_csamul_cla32_fa29_12_xor0 & s_csamul_cla32_fa29_11_or0;
  assign s_csamul_cla32_fa29_12_or0 = s_csamul_cla32_fa29_12_and0 | s_csamul_cla32_fa29_12_and1;
  assign s_csamul_cla32_and30_12 = a[30] & b[12];
  assign s_csamul_cla32_fa30_12_xor0 = s_csamul_cla32_and30_12 ^ s_csamul_cla32_ha31_11_xor0;
  assign s_csamul_cla32_fa30_12_and0 = s_csamul_cla32_and30_12 & s_csamul_cla32_ha31_11_xor0;
  assign s_csamul_cla32_fa30_12_xor1 = s_csamul_cla32_fa30_12_xor0 ^ s_csamul_cla32_fa30_11_or0;
  assign s_csamul_cla32_fa30_12_and1 = s_csamul_cla32_fa30_12_xor0 & s_csamul_cla32_fa30_11_or0;
  assign s_csamul_cla32_fa30_12_or0 = s_csamul_cla32_fa30_12_and0 | s_csamul_cla32_fa30_12_and1;
  assign s_csamul_cla32_nand31_12 = ~(a[31] & b[12]);
  assign s_csamul_cla32_ha31_12_xor0 = s_csamul_cla32_nand31_12 ^ s_csamul_cla32_ha31_11_and0;
  assign s_csamul_cla32_ha31_12_and0 = s_csamul_cla32_nand31_12 & s_csamul_cla32_ha31_11_and0;
  assign s_csamul_cla32_and0_13 = a[0] & b[13];
  assign s_csamul_cla32_fa0_13_xor0 = s_csamul_cla32_and0_13 ^ s_csamul_cla32_fa1_12_xor1;
  assign s_csamul_cla32_fa0_13_and0 = s_csamul_cla32_and0_13 & s_csamul_cla32_fa1_12_xor1;
  assign s_csamul_cla32_fa0_13_xor1 = s_csamul_cla32_fa0_13_xor0 ^ s_csamul_cla32_fa0_12_or0;
  assign s_csamul_cla32_fa0_13_and1 = s_csamul_cla32_fa0_13_xor0 & s_csamul_cla32_fa0_12_or0;
  assign s_csamul_cla32_fa0_13_or0 = s_csamul_cla32_fa0_13_and0 | s_csamul_cla32_fa0_13_and1;
  assign s_csamul_cla32_and1_13 = a[1] & b[13];
  assign s_csamul_cla32_fa1_13_xor0 = s_csamul_cla32_and1_13 ^ s_csamul_cla32_fa2_12_xor1;
  assign s_csamul_cla32_fa1_13_and0 = s_csamul_cla32_and1_13 & s_csamul_cla32_fa2_12_xor1;
  assign s_csamul_cla32_fa1_13_xor1 = s_csamul_cla32_fa1_13_xor0 ^ s_csamul_cla32_fa1_12_or0;
  assign s_csamul_cla32_fa1_13_and1 = s_csamul_cla32_fa1_13_xor0 & s_csamul_cla32_fa1_12_or0;
  assign s_csamul_cla32_fa1_13_or0 = s_csamul_cla32_fa1_13_and0 | s_csamul_cla32_fa1_13_and1;
  assign s_csamul_cla32_and2_13 = a[2] & b[13];
  assign s_csamul_cla32_fa2_13_xor0 = s_csamul_cla32_and2_13 ^ s_csamul_cla32_fa3_12_xor1;
  assign s_csamul_cla32_fa2_13_and0 = s_csamul_cla32_and2_13 & s_csamul_cla32_fa3_12_xor1;
  assign s_csamul_cla32_fa2_13_xor1 = s_csamul_cla32_fa2_13_xor0 ^ s_csamul_cla32_fa2_12_or0;
  assign s_csamul_cla32_fa2_13_and1 = s_csamul_cla32_fa2_13_xor0 & s_csamul_cla32_fa2_12_or0;
  assign s_csamul_cla32_fa2_13_or0 = s_csamul_cla32_fa2_13_and0 | s_csamul_cla32_fa2_13_and1;
  assign s_csamul_cla32_and3_13 = a[3] & b[13];
  assign s_csamul_cla32_fa3_13_xor0 = s_csamul_cla32_and3_13 ^ s_csamul_cla32_fa4_12_xor1;
  assign s_csamul_cla32_fa3_13_and0 = s_csamul_cla32_and3_13 & s_csamul_cla32_fa4_12_xor1;
  assign s_csamul_cla32_fa3_13_xor1 = s_csamul_cla32_fa3_13_xor0 ^ s_csamul_cla32_fa3_12_or0;
  assign s_csamul_cla32_fa3_13_and1 = s_csamul_cla32_fa3_13_xor0 & s_csamul_cla32_fa3_12_or0;
  assign s_csamul_cla32_fa3_13_or0 = s_csamul_cla32_fa3_13_and0 | s_csamul_cla32_fa3_13_and1;
  assign s_csamul_cla32_and4_13 = a[4] & b[13];
  assign s_csamul_cla32_fa4_13_xor0 = s_csamul_cla32_and4_13 ^ s_csamul_cla32_fa5_12_xor1;
  assign s_csamul_cla32_fa4_13_and0 = s_csamul_cla32_and4_13 & s_csamul_cla32_fa5_12_xor1;
  assign s_csamul_cla32_fa4_13_xor1 = s_csamul_cla32_fa4_13_xor0 ^ s_csamul_cla32_fa4_12_or0;
  assign s_csamul_cla32_fa4_13_and1 = s_csamul_cla32_fa4_13_xor0 & s_csamul_cla32_fa4_12_or0;
  assign s_csamul_cla32_fa4_13_or0 = s_csamul_cla32_fa4_13_and0 | s_csamul_cla32_fa4_13_and1;
  assign s_csamul_cla32_and5_13 = a[5] & b[13];
  assign s_csamul_cla32_fa5_13_xor0 = s_csamul_cla32_and5_13 ^ s_csamul_cla32_fa6_12_xor1;
  assign s_csamul_cla32_fa5_13_and0 = s_csamul_cla32_and5_13 & s_csamul_cla32_fa6_12_xor1;
  assign s_csamul_cla32_fa5_13_xor1 = s_csamul_cla32_fa5_13_xor0 ^ s_csamul_cla32_fa5_12_or0;
  assign s_csamul_cla32_fa5_13_and1 = s_csamul_cla32_fa5_13_xor0 & s_csamul_cla32_fa5_12_or0;
  assign s_csamul_cla32_fa5_13_or0 = s_csamul_cla32_fa5_13_and0 | s_csamul_cla32_fa5_13_and1;
  assign s_csamul_cla32_and6_13 = a[6] & b[13];
  assign s_csamul_cla32_fa6_13_xor0 = s_csamul_cla32_and6_13 ^ s_csamul_cla32_fa7_12_xor1;
  assign s_csamul_cla32_fa6_13_and0 = s_csamul_cla32_and6_13 & s_csamul_cla32_fa7_12_xor1;
  assign s_csamul_cla32_fa6_13_xor1 = s_csamul_cla32_fa6_13_xor0 ^ s_csamul_cla32_fa6_12_or0;
  assign s_csamul_cla32_fa6_13_and1 = s_csamul_cla32_fa6_13_xor0 & s_csamul_cla32_fa6_12_or0;
  assign s_csamul_cla32_fa6_13_or0 = s_csamul_cla32_fa6_13_and0 | s_csamul_cla32_fa6_13_and1;
  assign s_csamul_cla32_and7_13 = a[7] & b[13];
  assign s_csamul_cla32_fa7_13_xor0 = s_csamul_cla32_and7_13 ^ s_csamul_cla32_fa8_12_xor1;
  assign s_csamul_cla32_fa7_13_and0 = s_csamul_cla32_and7_13 & s_csamul_cla32_fa8_12_xor1;
  assign s_csamul_cla32_fa7_13_xor1 = s_csamul_cla32_fa7_13_xor0 ^ s_csamul_cla32_fa7_12_or0;
  assign s_csamul_cla32_fa7_13_and1 = s_csamul_cla32_fa7_13_xor0 & s_csamul_cla32_fa7_12_or0;
  assign s_csamul_cla32_fa7_13_or0 = s_csamul_cla32_fa7_13_and0 | s_csamul_cla32_fa7_13_and1;
  assign s_csamul_cla32_and8_13 = a[8] & b[13];
  assign s_csamul_cla32_fa8_13_xor0 = s_csamul_cla32_and8_13 ^ s_csamul_cla32_fa9_12_xor1;
  assign s_csamul_cla32_fa8_13_and0 = s_csamul_cla32_and8_13 & s_csamul_cla32_fa9_12_xor1;
  assign s_csamul_cla32_fa8_13_xor1 = s_csamul_cla32_fa8_13_xor0 ^ s_csamul_cla32_fa8_12_or0;
  assign s_csamul_cla32_fa8_13_and1 = s_csamul_cla32_fa8_13_xor0 & s_csamul_cla32_fa8_12_or0;
  assign s_csamul_cla32_fa8_13_or0 = s_csamul_cla32_fa8_13_and0 | s_csamul_cla32_fa8_13_and1;
  assign s_csamul_cla32_and9_13 = a[9] & b[13];
  assign s_csamul_cla32_fa9_13_xor0 = s_csamul_cla32_and9_13 ^ s_csamul_cla32_fa10_12_xor1;
  assign s_csamul_cla32_fa9_13_and0 = s_csamul_cla32_and9_13 & s_csamul_cla32_fa10_12_xor1;
  assign s_csamul_cla32_fa9_13_xor1 = s_csamul_cla32_fa9_13_xor0 ^ s_csamul_cla32_fa9_12_or0;
  assign s_csamul_cla32_fa9_13_and1 = s_csamul_cla32_fa9_13_xor0 & s_csamul_cla32_fa9_12_or0;
  assign s_csamul_cla32_fa9_13_or0 = s_csamul_cla32_fa9_13_and0 | s_csamul_cla32_fa9_13_and1;
  assign s_csamul_cla32_and10_13 = a[10] & b[13];
  assign s_csamul_cla32_fa10_13_xor0 = s_csamul_cla32_and10_13 ^ s_csamul_cla32_fa11_12_xor1;
  assign s_csamul_cla32_fa10_13_and0 = s_csamul_cla32_and10_13 & s_csamul_cla32_fa11_12_xor1;
  assign s_csamul_cla32_fa10_13_xor1 = s_csamul_cla32_fa10_13_xor0 ^ s_csamul_cla32_fa10_12_or0;
  assign s_csamul_cla32_fa10_13_and1 = s_csamul_cla32_fa10_13_xor0 & s_csamul_cla32_fa10_12_or0;
  assign s_csamul_cla32_fa10_13_or0 = s_csamul_cla32_fa10_13_and0 | s_csamul_cla32_fa10_13_and1;
  assign s_csamul_cla32_and11_13 = a[11] & b[13];
  assign s_csamul_cla32_fa11_13_xor0 = s_csamul_cla32_and11_13 ^ s_csamul_cla32_fa12_12_xor1;
  assign s_csamul_cla32_fa11_13_and0 = s_csamul_cla32_and11_13 & s_csamul_cla32_fa12_12_xor1;
  assign s_csamul_cla32_fa11_13_xor1 = s_csamul_cla32_fa11_13_xor0 ^ s_csamul_cla32_fa11_12_or0;
  assign s_csamul_cla32_fa11_13_and1 = s_csamul_cla32_fa11_13_xor0 & s_csamul_cla32_fa11_12_or0;
  assign s_csamul_cla32_fa11_13_or0 = s_csamul_cla32_fa11_13_and0 | s_csamul_cla32_fa11_13_and1;
  assign s_csamul_cla32_and12_13 = a[12] & b[13];
  assign s_csamul_cla32_fa12_13_xor0 = s_csamul_cla32_and12_13 ^ s_csamul_cla32_fa13_12_xor1;
  assign s_csamul_cla32_fa12_13_and0 = s_csamul_cla32_and12_13 & s_csamul_cla32_fa13_12_xor1;
  assign s_csamul_cla32_fa12_13_xor1 = s_csamul_cla32_fa12_13_xor0 ^ s_csamul_cla32_fa12_12_or0;
  assign s_csamul_cla32_fa12_13_and1 = s_csamul_cla32_fa12_13_xor0 & s_csamul_cla32_fa12_12_or0;
  assign s_csamul_cla32_fa12_13_or0 = s_csamul_cla32_fa12_13_and0 | s_csamul_cla32_fa12_13_and1;
  assign s_csamul_cla32_and13_13 = a[13] & b[13];
  assign s_csamul_cla32_fa13_13_xor0 = s_csamul_cla32_and13_13 ^ s_csamul_cla32_fa14_12_xor1;
  assign s_csamul_cla32_fa13_13_and0 = s_csamul_cla32_and13_13 & s_csamul_cla32_fa14_12_xor1;
  assign s_csamul_cla32_fa13_13_xor1 = s_csamul_cla32_fa13_13_xor0 ^ s_csamul_cla32_fa13_12_or0;
  assign s_csamul_cla32_fa13_13_and1 = s_csamul_cla32_fa13_13_xor0 & s_csamul_cla32_fa13_12_or0;
  assign s_csamul_cla32_fa13_13_or0 = s_csamul_cla32_fa13_13_and0 | s_csamul_cla32_fa13_13_and1;
  assign s_csamul_cla32_and14_13 = a[14] & b[13];
  assign s_csamul_cla32_fa14_13_xor0 = s_csamul_cla32_and14_13 ^ s_csamul_cla32_fa15_12_xor1;
  assign s_csamul_cla32_fa14_13_and0 = s_csamul_cla32_and14_13 & s_csamul_cla32_fa15_12_xor1;
  assign s_csamul_cla32_fa14_13_xor1 = s_csamul_cla32_fa14_13_xor0 ^ s_csamul_cla32_fa14_12_or0;
  assign s_csamul_cla32_fa14_13_and1 = s_csamul_cla32_fa14_13_xor0 & s_csamul_cla32_fa14_12_or0;
  assign s_csamul_cla32_fa14_13_or0 = s_csamul_cla32_fa14_13_and0 | s_csamul_cla32_fa14_13_and1;
  assign s_csamul_cla32_and15_13 = a[15] & b[13];
  assign s_csamul_cla32_fa15_13_xor0 = s_csamul_cla32_and15_13 ^ s_csamul_cla32_fa16_12_xor1;
  assign s_csamul_cla32_fa15_13_and0 = s_csamul_cla32_and15_13 & s_csamul_cla32_fa16_12_xor1;
  assign s_csamul_cla32_fa15_13_xor1 = s_csamul_cla32_fa15_13_xor0 ^ s_csamul_cla32_fa15_12_or0;
  assign s_csamul_cla32_fa15_13_and1 = s_csamul_cla32_fa15_13_xor0 & s_csamul_cla32_fa15_12_or0;
  assign s_csamul_cla32_fa15_13_or0 = s_csamul_cla32_fa15_13_and0 | s_csamul_cla32_fa15_13_and1;
  assign s_csamul_cla32_and16_13 = a[16] & b[13];
  assign s_csamul_cla32_fa16_13_xor0 = s_csamul_cla32_and16_13 ^ s_csamul_cla32_fa17_12_xor1;
  assign s_csamul_cla32_fa16_13_and0 = s_csamul_cla32_and16_13 & s_csamul_cla32_fa17_12_xor1;
  assign s_csamul_cla32_fa16_13_xor1 = s_csamul_cla32_fa16_13_xor0 ^ s_csamul_cla32_fa16_12_or0;
  assign s_csamul_cla32_fa16_13_and1 = s_csamul_cla32_fa16_13_xor0 & s_csamul_cla32_fa16_12_or0;
  assign s_csamul_cla32_fa16_13_or0 = s_csamul_cla32_fa16_13_and0 | s_csamul_cla32_fa16_13_and1;
  assign s_csamul_cla32_and17_13 = a[17] & b[13];
  assign s_csamul_cla32_fa17_13_xor0 = s_csamul_cla32_and17_13 ^ s_csamul_cla32_fa18_12_xor1;
  assign s_csamul_cla32_fa17_13_and0 = s_csamul_cla32_and17_13 & s_csamul_cla32_fa18_12_xor1;
  assign s_csamul_cla32_fa17_13_xor1 = s_csamul_cla32_fa17_13_xor0 ^ s_csamul_cla32_fa17_12_or0;
  assign s_csamul_cla32_fa17_13_and1 = s_csamul_cla32_fa17_13_xor0 & s_csamul_cla32_fa17_12_or0;
  assign s_csamul_cla32_fa17_13_or0 = s_csamul_cla32_fa17_13_and0 | s_csamul_cla32_fa17_13_and1;
  assign s_csamul_cla32_and18_13 = a[18] & b[13];
  assign s_csamul_cla32_fa18_13_xor0 = s_csamul_cla32_and18_13 ^ s_csamul_cla32_fa19_12_xor1;
  assign s_csamul_cla32_fa18_13_and0 = s_csamul_cla32_and18_13 & s_csamul_cla32_fa19_12_xor1;
  assign s_csamul_cla32_fa18_13_xor1 = s_csamul_cla32_fa18_13_xor0 ^ s_csamul_cla32_fa18_12_or0;
  assign s_csamul_cla32_fa18_13_and1 = s_csamul_cla32_fa18_13_xor0 & s_csamul_cla32_fa18_12_or0;
  assign s_csamul_cla32_fa18_13_or0 = s_csamul_cla32_fa18_13_and0 | s_csamul_cla32_fa18_13_and1;
  assign s_csamul_cla32_and19_13 = a[19] & b[13];
  assign s_csamul_cla32_fa19_13_xor0 = s_csamul_cla32_and19_13 ^ s_csamul_cla32_fa20_12_xor1;
  assign s_csamul_cla32_fa19_13_and0 = s_csamul_cla32_and19_13 & s_csamul_cla32_fa20_12_xor1;
  assign s_csamul_cla32_fa19_13_xor1 = s_csamul_cla32_fa19_13_xor0 ^ s_csamul_cla32_fa19_12_or0;
  assign s_csamul_cla32_fa19_13_and1 = s_csamul_cla32_fa19_13_xor0 & s_csamul_cla32_fa19_12_or0;
  assign s_csamul_cla32_fa19_13_or0 = s_csamul_cla32_fa19_13_and0 | s_csamul_cla32_fa19_13_and1;
  assign s_csamul_cla32_and20_13 = a[20] & b[13];
  assign s_csamul_cla32_fa20_13_xor0 = s_csamul_cla32_and20_13 ^ s_csamul_cla32_fa21_12_xor1;
  assign s_csamul_cla32_fa20_13_and0 = s_csamul_cla32_and20_13 & s_csamul_cla32_fa21_12_xor1;
  assign s_csamul_cla32_fa20_13_xor1 = s_csamul_cla32_fa20_13_xor0 ^ s_csamul_cla32_fa20_12_or0;
  assign s_csamul_cla32_fa20_13_and1 = s_csamul_cla32_fa20_13_xor0 & s_csamul_cla32_fa20_12_or0;
  assign s_csamul_cla32_fa20_13_or0 = s_csamul_cla32_fa20_13_and0 | s_csamul_cla32_fa20_13_and1;
  assign s_csamul_cla32_and21_13 = a[21] & b[13];
  assign s_csamul_cla32_fa21_13_xor0 = s_csamul_cla32_and21_13 ^ s_csamul_cla32_fa22_12_xor1;
  assign s_csamul_cla32_fa21_13_and0 = s_csamul_cla32_and21_13 & s_csamul_cla32_fa22_12_xor1;
  assign s_csamul_cla32_fa21_13_xor1 = s_csamul_cla32_fa21_13_xor0 ^ s_csamul_cla32_fa21_12_or0;
  assign s_csamul_cla32_fa21_13_and1 = s_csamul_cla32_fa21_13_xor0 & s_csamul_cla32_fa21_12_or0;
  assign s_csamul_cla32_fa21_13_or0 = s_csamul_cla32_fa21_13_and0 | s_csamul_cla32_fa21_13_and1;
  assign s_csamul_cla32_and22_13 = a[22] & b[13];
  assign s_csamul_cla32_fa22_13_xor0 = s_csamul_cla32_and22_13 ^ s_csamul_cla32_fa23_12_xor1;
  assign s_csamul_cla32_fa22_13_and0 = s_csamul_cla32_and22_13 & s_csamul_cla32_fa23_12_xor1;
  assign s_csamul_cla32_fa22_13_xor1 = s_csamul_cla32_fa22_13_xor0 ^ s_csamul_cla32_fa22_12_or0;
  assign s_csamul_cla32_fa22_13_and1 = s_csamul_cla32_fa22_13_xor0 & s_csamul_cla32_fa22_12_or0;
  assign s_csamul_cla32_fa22_13_or0 = s_csamul_cla32_fa22_13_and0 | s_csamul_cla32_fa22_13_and1;
  assign s_csamul_cla32_and23_13 = a[23] & b[13];
  assign s_csamul_cla32_fa23_13_xor0 = s_csamul_cla32_and23_13 ^ s_csamul_cla32_fa24_12_xor1;
  assign s_csamul_cla32_fa23_13_and0 = s_csamul_cla32_and23_13 & s_csamul_cla32_fa24_12_xor1;
  assign s_csamul_cla32_fa23_13_xor1 = s_csamul_cla32_fa23_13_xor0 ^ s_csamul_cla32_fa23_12_or0;
  assign s_csamul_cla32_fa23_13_and1 = s_csamul_cla32_fa23_13_xor0 & s_csamul_cla32_fa23_12_or0;
  assign s_csamul_cla32_fa23_13_or0 = s_csamul_cla32_fa23_13_and0 | s_csamul_cla32_fa23_13_and1;
  assign s_csamul_cla32_and24_13 = a[24] & b[13];
  assign s_csamul_cla32_fa24_13_xor0 = s_csamul_cla32_and24_13 ^ s_csamul_cla32_fa25_12_xor1;
  assign s_csamul_cla32_fa24_13_and0 = s_csamul_cla32_and24_13 & s_csamul_cla32_fa25_12_xor1;
  assign s_csamul_cla32_fa24_13_xor1 = s_csamul_cla32_fa24_13_xor0 ^ s_csamul_cla32_fa24_12_or0;
  assign s_csamul_cla32_fa24_13_and1 = s_csamul_cla32_fa24_13_xor0 & s_csamul_cla32_fa24_12_or0;
  assign s_csamul_cla32_fa24_13_or0 = s_csamul_cla32_fa24_13_and0 | s_csamul_cla32_fa24_13_and1;
  assign s_csamul_cla32_and25_13 = a[25] & b[13];
  assign s_csamul_cla32_fa25_13_xor0 = s_csamul_cla32_and25_13 ^ s_csamul_cla32_fa26_12_xor1;
  assign s_csamul_cla32_fa25_13_and0 = s_csamul_cla32_and25_13 & s_csamul_cla32_fa26_12_xor1;
  assign s_csamul_cla32_fa25_13_xor1 = s_csamul_cla32_fa25_13_xor0 ^ s_csamul_cla32_fa25_12_or0;
  assign s_csamul_cla32_fa25_13_and1 = s_csamul_cla32_fa25_13_xor0 & s_csamul_cla32_fa25_12_or0;
  assign s_csamul_cla32_fa25_13_or0 = s_csamul_cla32_fa25_13_and0 | s_csamul_cla32_fa25_13_and1;
  assign s_csamul_cla32_and26_13 = a[26] & b[13];
  assign s_csamul_cla32_fa26_13_xor0 = s_csamul_cla32_and26_13 ^ s_csamul_cla32_fa27_12_xor1;
  assign s_csamul_cla32_fa26_13_and0 = s_csamul_cla32_and26_13 & s_csamul_cla32_fa27_12_xor1;
  assign s_csamul_cla32_fa26_13_xor1 = s_csamul_cla32_fa26_13_xor0 ^ s_csamul_cla32_fa26_12_or0;
  assign s_csamul_cla32_fa26_13_and1 = s_csamul_cla32_fa26_13_xor0 & s_csamul_cla32_fa26_12_or0;
  assign s_csamul_cla32_fa26_13_or0 = s_csamul_cla32_fa26_13_and0 | s_csamul_cla32_fa26_13_and1;
  assign s_csamul_cla32_and27_13 = a[27] & b[13];
  assign s_csamul_cla32_fa27_13_xor0 = s_csamul_cla32_and27_13 ^ s_csamul_cla32_fa28_12_xor1;
  assign s_csamul_cla32_fa27_13_and0 = s_csamul_cla32_and27_13 & s_csamul_cla32_fa28_12_xor1;
  assign s_csamul_cla32_fa27_13_xor1 = s_csamul_cla32_fa27_13_xor0 ^ s_csamul_cla32_fa27_12_or0;
  assign s_csamul_cla32_fa27_13_and1 = s_csamul_cla32_fa27_13_xor0 & s_csamul_cla32_fa27_12_or0;
  assign s_csamul_cla32_fa27_13_or0 = s_csamul_cla32_fa27_13_and0 | s_csamul_cla32_fa27_13_and1;
  assign s_csamul_cla32_and28_13 = a[28] & b[13];
  assign s_csamul_cla32_fa28_13_xor0 = s_csamul_cla32_and28_13 ^ s_csamul_cla32_fa29_12_xor1;
  assign s_csamul_cla32_fa28_13_and0 = s_csamul_cla32_and28_13 & s_csamul_cla32_fa29_12_xor1;
  assign s_csamul_cla32_fa28_13_xor1 = s_csamul_cla32_fa28_13_xor0 ^ s_csamul_cla32_fa28_12_or0;
  assign s_csamul_cla32_fa28_13_and1 = s_csamul_cla32_fa28_13_xor0 & s_csamul_cla32_fa28_12_or0;
  assign s_csamul_cla32_fa28_13_or0 = s_csamul_cla32_fa28_13_and0 | s_csamul_cla32_fa28_13_and1;
  assign s_csamul_cla32_and29_13 = a[29] & b[13];
  assign s_csamul_cla32_fa29_13_xor0 = s_csamul_cla32_and29_13 ^ s_csamul_cla32_fa30_12_xor1;
  assign s_csamul_cla32_fa29_13_and0 = s_csamul_cla32_and29_13 & s_csamul_cla32_fa30_12_xor1;
  assign s_csamul_cla32_fa29_13_xor1 = s_csamul_cla32_fa29_13_xor0 ^ s_csamul_cla32_fa29_12_or0;
  assign s_csamul_cla32_fa29_13_and1 = s_csamul_cla32_fa29_13_xor0 & s_csamul_cla32_fa29_12_or0;
  assign s_csamul_cla32_fa29_13_or0 = s_csamul_cla32_fa29_13_and0 | s_csamul_cla32_fa29_13_and1;
  assign s_csamul_cla32_and30_13 = a[30] & b[13];
  assign s_csamul_cla32_fa30_13_xor0 = s_csamul_cla32_and30_13 ^ s_csamul_cla32_ha31_12_xor0;
  assign s_csamul_cla32_fa30_13_and0 = s_csamul_cla32_and30_13 & s_csamul_cla32_ha31_12_xor0;
  assign s_csamul_cla32_fa30_13_xor1 = s_csamul_cla32_fa30_13_xor0 ^ s_csamul_cla32_fa30_12_or0;
  assign s_csamul_cla32_fa30_13_and1 = s_csamul_cla32_fa30_13_xor0 & s_csamul_cla32_fa30_12_or0;
  assign s_csamul_cla32_fa30_13_or0 = s_csamul_cla32_fa30_13_and0 | s_csamul_cla32_fa30_13_and1;
  assign s_csamul_cla32_nand31_13 = ~(a[31] & b[13]);
  assign s_csamul_cla32_ha31_13_xor0 = s_csamul_cla32_nand31_13 ^ s_csamul_cla32_ha31_12_and0;
  assign s_csamul_cla32_ha31_13_and0 = s_csamul_cla32_nand31_13 & s_csamul_cla32_ha31_12_and0;
  assign s_csamul_cla32_and0_14 = a[0] & b[14];
  assign s_csamul_cla32_fa0_14_xor0 = s_csamul_cla32_and0_14 ^ s_csamul_cla32_fa1_13_xor1;
  assign s_csamul_cla32_fa0_14_and0 = s_csamul_cla32_and0_14 & s_csamul_cla32_fa1_13_xor1;
  assign s_csamul_cla32_fa0_14_xor1 = s_csamul_cla32_fa0_14_xor0 ^ s_csamul_cla32_fa0_13_or0;
  assign s_csamul_cla32_fa0_14_and1 = s_csamul_cla32_fa0_14_xor0 & s_csamul_cla32_fa0_13_or0;
  assign s_csamul_cla32_fa0_14_or0 = s_csamul_cla32_fa0_14_and0 | s_csamul_cla32_fa0_14_and1;
  assign s_csamul_cla32_and1_14 = a[1] & b[14];
  assign s_csamul_cla32_fa1_14_xor0 = s_csamul_cla32_and1_14 ^ s_csamul_cla32_fa2_13_xor1;
  assign s_csamul_cla32_fa1_14_and0 = s_csamul_cla32_and1_14 & s_csamul_cla32_fa2_13_xor1;
  assign s_csamul_cla32_fa1_14_xor1 = s_csamul_cla32_fa1_14_xor0 ^ s_csamul_cla32_fa1_13_or0;
  assign s_csamul_cla32_fa1_14_and1 = s_csamul_cla32_fa1_14_xor0 & s_csamul_cla32_fa1_13_or0;
  assign s_csamul_cla32_fa1_14_or0 = s_csamul_cla32_fa1_14_and0 | s_csamul_cla32_fa1_14_and1;
  assign s_csamul_cla32_and2_14 = a[2] & b[14];
  assign s_csamul_cla32_fa2_14_xor0 = s_csamul_cla32_and2_14 ^ s_csamul_cla32_fa3_13_xor1;
  assign s_csamul_cla32_fa2_14_and0 = s_csamul_cla32_and2_14 & s_csamul_cla32_fa3_13_xor1;
  assign s_csamul_cla32_fa2_14_xor1 = s_csamul_cla32_fa2_14_xor0 ^ s_csamul_cla32_fa2_13_or0;
  assign s_csamul_cla32_fa2_14_and1 = s_csamul_cla32_fa2_14_xor0 & s_csamul_cla32_fa2_13_or0;
  assign s_csamul_cla32_fa2_14_or0 = s_csamul_cla32_fa2_14_and0 | s_csamul_cla32_fa2_14_and1;
  assign s_csamul_cla32_and3_14 = a[3] & b[14];
  assign s_csamul_cla32_fa3_14_xor0 = s_csamul_cla32_and3_14 ^ s_csamul_cla32_fa4_13_xor1;
  assign s_csamul_cla32_fa3_14_and0 = s_csamul_cla32_and3_14 & s_csamul_cla32_fa4_13_xor1;
  assign s_csamul_cla32_fa3_14_xor1 = s_csamul_cla32_fa3_14_xor0 ^ s_csamul_cla32_fa3_13_or0;
  assign s_csamul_cla32_fa3_14_and1 = s_csamul_cla32_fa3_14_xor0 & s_csamul_cla32_fa3_13_or0;
  assign s_csamul_cla32_fa3_14_or0 = s_csamul_cla32_fa3_14_and0 | s_csamul_cla32_fa3_14_and1;
  assign s_csamul_cla32_and4_14 = a[4] & b[14];
  assign s_csamul_cla32_fa4_14_xor0 = s_csamul_cla32_and4_14 ^ s_csamul_cla32_fa5_13_xor1;
  assign s_csamul_cla32_fa4_14_and0 = s_csamul_cla32_and4_14 & s_csamul_cla32_fa5_13_xor1;
  assign s_csamul_cla32_fa4_14_xor1 = s_csamul_cla32_fa4_14_xor0 ^ s_csamul_cla32_fa4_13_or0;
  assign s_csamul_cla32_fa4_14_and1 = s_csamul_cla32_fa4_14_xor0 & s_csamul_cla32_fa4_13_or0;
  assign s_csamul_cla32_fa4_14_or0 = s_csamul_cla32_fa4_14_and0 | s_csamul_cla32_fa4_14_and1;
  assign s_csamul_cla32_and5_14 = a[5] & b[14];
  assign s_csamul_cla32_fa5_14_xor0 = s_csamul_cla32_and5_14 ^ s_csamul_cla32_fa6_13_xor1;
  assign s_csamul_cla32_fa5_14_and0 = s_csamul_cla32_and5_14 & s_csamul_cla32_fa6_13_xor1;
  assign s_csamul_cla32_fa5_14_xor1 = s_csamul_cla32_fa5_14_xor0 ^ s_csamul_cla32_fa5_13_or0;
  assign s_csamul_cla32_fa5_14_and1 = s_csamul_cla32_fa5_14_xor0 & s_csamul_cla32_fa5_13_or0;
  assign s_csamul_cla32_fa5_14_or0 = s_csamul_cla32_fa5_14_and0 | s_csamul_cla32_fa5_14_and1;
  assign s_csamul_cla32_and6_14 = a[6] & b[14];
  assign s_csamul_cla32_fa6_14_xor0 = s_csamul_cla32_and6_14 ^ s_csamul_cla32_fa7_13_xor1;
  assign s_csamul_cla32_fa6_14_and0 = s_csamul_cla32_and6_14 & s_csamul_cla32_fa7_13_xor1;
  assign s_csamul_cla32_fa6_14_xor1 = s_csamul_cla32_fa6_14_xor0 ^ s_csamul_cla32_fa6_13_or0;
  assign s_csamul_cla32_fa6_14_and1 = s_csamul_cla32_fa6_14_xor0 & s_csamul_cla32_fa6_13_or0;
  assign s_csamul_cla32_fa6_14_or0 = s_csamul_cla32_fa6_14_and0 | s_csamul_cla32_fa6_14_and1;
  assign s_csamul_cla32_and7_14 = a[7] & b[14];
  assign s_csamul_cla32_fa7_14_xor0 = s_csamul_cla32_and7_14 ^ s_csamul_cla32_fa8_13_xor1;
  assign s_csamul_cla32_fa7_14_and0 = s_csamul_cla32_and7_14 & s_csamul_cla32_fa8_13_xor1;
  assign s_csamul_cla32_fa7_14_xor1 = s_csamul_cla32_fa7_14_xor0 ^ s_csamul_cla32_fa7_13_or0;
  assign s_csamul_cla32_fa7_14_and1 = s_csamul_cla32_fa7_14_xor0 & s_csamul_cla32_fa7_13_or0;
  assign s_csamul_cla32_fa7_14_or0 = s_csamul_cla32_fa7_14_and0 | s_csamul_cla32_fa7_14_and1;
  assign s_csamul_cla32_and8_14 = a[8] & b[14];
  assign s_csamul_cla32_fa8_14_xor0 = s_csamul_cla32_and8_14 ^ s_csamul_cla32_fa9_13_xor1;
  assign s_csamul_cla32_fa8_14_and0 = s_csamul_cla32_and8_14 & s_csamul_cla32_fa9_13_xor1;
  assign s_csamul_cla32_fa8_14_xor1 = s_csamul_cla32_fa8_14_xor0 ^ s_csamul_cla32_fa8_13_or0;
  assign s_csamul_cla32_fa8_14_and1 = s_csamul_cla32_fa8_14_xor0 & s_csamul_cla32_fa8_13_or0;
  assign s_csamul_cla32_fa8_14_or0 = s_csamul_cla32_fa8_14_and0 | s_csamul_cla32_fa8_14_and1;
  assign s_csamul_cla32_and9_14 = a[9] & b[14];
  assign s_csamul_cla32_fa9_14_xor0 = s_csamul_cla32_and9_14 ^ s_csamul_cla32_fa10_13_xor1;
  assign s_csamul_cla32_fa9_14_and0 = s_csamul_cla32_and9_14 & s_csamul_cla32_fa10_13_xor1;
  assign s_csamul_cla32_fa9_14_xor1 = s_csamul_cla32_fa9_14_xor0 ^ s_csamul_cla32_fa9_13_or0;
  assign s_csamul_cla32_fa9_14_and1 = s_csamul_cla32_fa9_14_xor0 & s_csamul_cla32_fa9_13_or0;
  assign s_csamul_cla32_fa9_14_or0 = s_csamul_cla32_fa9_14_and0 | s_csamul_cla32_fa9_14_and1;
  assign s_csamul_cla32_and10_14 = a[10] & b[14];
  assign s_csamul_cla32_fa10_14_xor0 = s_csamul_cla32_and10_14 ^ s_csamul_cla32_fa11_13_xor1;
  assign s_csamul_cla32_fa10_14_and0 = s_csamul_cla32_and10_14 & s_csamul_cla32_fa11_13_xor1;
  assign s_csamul_cla32_fa10_14_xor1 = s_csamul_cla32_fa10_14_xor0 ^ s_csamul_cla32_fa10_13_or0;
  assign s_csamul_cla32_fa10_14_and1 = s_csamul_cla32_fa10_14_xor0 & s_csamul_cla32_fa10_13_or0;
  assign s_csamul_cla32_fa10_14_or0 = s_csamul_cla32_fa10_14_and0 | s_csamul_cla32_fa10_14_and1;
  assign s_csamul_cla32_and11_14 = a[11] & b[14];
  assign s_csamul_cla32_fa11_14_xor0 = s_csamul_cla32_and11_14 ^ s_csamul_cla32_fa12_13_xor1;
  assign s_csamul_cla32_fa11_14_and0 = s_csamul_cla32_and11_14 & s_csamul_cla32_fa12_13_xor1;
  assign s_csamul_cla32_fa11_14_xor1 = s_csamul_cla32_fa11_14_xor0 ^ s_csamul_cla32_fa11_13_or0;
  assign s_csamul_cla32_fa11_14_and1 = s_csamul_cla32_fa11_14_xor0 & s_csamul_cla32_fa11_13_or0;
  assign s_csamul_cla32_fa11_14_or0 = s_csamul_cla32_fa11_14_and0 | s_csamul_cla32_fa11_14_and1;
  assign s_csamul_cla32_and12_14 = a[12] & b[14];
  assign s_csamul_cla32_fa12_14_xor0 = s_csamul_cla32_and12_14 ^ s_csamul_cla32_fa13_13_xor1;
  assign s_csamul_cla32_fa12_14_and0 = s_csamul_cla32_and12_14 & s_csamul_cla32_fa13_13_xor1;
  assign s_csamul_cla32_fa12_14_xor1 = s_csamul_cla32_fa12_14_xor0 ^ s_csamul_cla32_fa12_13_or0;
  assign s_csamul_cla32_fa12_14_and1 = s_csamul_cla32_fa12_14_xor0 & s_csamul_cla32_fa12_13_or0;
  assign s_csamul_cla32_fa12_14_or0 = s_csamul_cla32_fa12_14_and0 | s_csamul_cla32_fa12_14_and1;
  assign s_csamul_cla32_and13_14 = a[13] & b[14];
  assign s_csamul_cla32_fa13_14_xor0 = s_csamul_cla32_and13_14 ^ s_csamul_cla32_fa14_13_xor1;
  assign s_csamul_cla32_fa13_14_and0 = s_csamul_cla32_and13_14 & s_csamul_cla32_fa14_13_xor1;
  assign s_csamul_cla32_fa13_14_xor1 = s_csamul_cla32_fa13_14_xor0 ^ s_csamul_cla32_fa13_13_or0;
  assign s_csamul_cla32_fa13_14_and1 = s_csamul_cla32_fa13_14_xor0 & s_csamul_cla32_fa13_13_or0;
  assign s_csamul_cla32_fa13_14_or0 = s_csamul_cla32_fa13_14_and0 | s_csamul_cla32_fa13_14_and1;
  assign s_csamul_cla32_and14_14 = a[14] & b[14];
  assign s_csamul_cla32_fa14_14_xor0 = s_csamul_cla32_and14_14 ^ s_csamul_cla32_fa15_13_xor1;
  assign s_csamul_cla32_fa14_14_and0 = s_csamul_cla32_and14_14 & s_csamul_cla32_fa15_13_xor1;
  assign s_csamul_cla32_fa14_14_xor1 = s_csamul_cla32_fa14_14_xor0 ^ s_csamul_cla32_fa14_13_or0;
  assign s_csamul_cla32_fa14_14_and1 = s_csamul_cla32_fa14_14_xor0 & s_csamul_cla32_fa14_13_or0;
  assign s_csamul_cla32_fa14_14_or0 = s_csamul_cla32_fa14_14_and0 | s_csamul_cla32_fa14_14_and1;
  assign s_csamul_cla32_and15_14 = a[15] & b[14];
  assign s_csamul_cla32_fa15_14_xor0 = s_csamul_cla32_and15_14 ^ s_csamul_cla32_fa16_13_xor1;
  assign s_csamul_cla32_fa15_14_and0 = s_csamul_cla32_and15_14 & s_csamul_cla32_fa16_13_xor1;
  assign s_csamul_cla32_fa15_14_xor1 = s_csamul_cla32_fa15_14_xor0 ^ s_csamul_cla32_fa15_13_or0;
  assign s_csamul_cla32_fa15_14_and1 = s_csamul_cla32_fa15_14_xor0 & s_csamul_cla32_fa15_13_or0;
  assign s_csamul_cla32_fa15_14_or0 = s_csamul_cla32_fa15_14_and0 | s_csamul_cla32_fa15_14_and1;
  assign s_csamul_cla32_and16_14 = a[16] & b[14];
  assign s_csamul_cla32_fa16_14_xor0 = s_csamul_cla32_and16_14 ^ s_csamul_cla32_fa17_13_xor1;
  assign s_csamul_cla32_fa16_14_and0 = s_csamul_cla32_and16_14 & s_csamul_cla32_fa17_13_xor1;
  assign s_csamul_cla32_fa16_14_xor1 = s_csamul_cla32_fa16_14_xor0 ^ s_csamul_cla32_fa16_13_or0;
  assign s_csamul_cla32_fa16_14_and1 = s_csamul_cla32_fa16_14_xor0 & s_csamul_cla32_fa16_13_or0;
  assign s_csamul_cla32_fa16_14_or0 = s_csamul_cla32_fa16_14_and0 | s_csamul_cla32_fa16_14_and1;
  assign s_csamul_cla32_and17_14 = a[17] & b[14];
  assign s_csamul_cla32_fa17_14_xor0 = s_csamul_cla32_and17_14 ^ s_csamul_cla32_fa18_13_xor1;
  assign s_csamul_cla32_fa17_14_and0 = s_csamul_cla32_and17_14 & s_csamul_cla32_fa18_13_xor1;
  assign s_csamul_cla32_fa17_14_xor1 = s_csamul_cla32_fa17_14_xor0 ^ s_csamul_cla32_fa17_13_or0;
  assign s_csamul_cla32_fa17_14_and1 = s_csamul_cla32_fa17_14_xor0 & s_csamul_cla32_fa17_13_or0;
  assign s_csamul_cla32_fa17_14_or0 = s_csamul_cla32_fa17_14_and0 | s_csamul_cla32_fa17_14_and1;
  assign s_csamul_cla32_and18_14 = a[18] & b[14];
  assign s_csamul_cla32_fa18_14_xor0 = s_csamul_cla32_and18_14 ^ s_csamul_cla32_fa19_13_xor1;
  assign s_csamul_cla32_fa18_14_and0 = s_csamul_cla32_and18_14 & s_csamul_cla32_fa19_13_xor1;
  assign s_csamul_cla32_fa18_14_xor1 = s_csamul_cla32_fa18_14_xor0 ^ s_csamul_cla32_fa18_13_or0;
  assign s_csamul_cla32_fa18_14_and1 = s_csamul_cla32_fa18_14_xor0 & s_csamul_cla32_fa18_13_or0;
  assign s_csamul_cla32_fa18_14_or0 = s_csamul_cla32_fa18_14_and0 | s_csamul_cla32_fa18_14_and1;
  assign s_csamul_cla32_and19_14 = a[19] & b[14];
  assign s_csamul_cla32_fa19_14_xor0 = s_csamul_cla32_and19_14 ^ s_csamul_cla32_fa20_13_xor1;
  assign s_csamul_cla32_fa19_14_and0 = s_csamul_cla32_and19_14 & s_csamul_cla32_fa20_13_xor1;
  assign s_csamul_cla32_fa19_14_xor1 = s_csamul_cla32_fa19_14_xor0 ^ s_csamul_cla32_fa19_13_or0;
  assign s_csamul_cla32_fa19_14_and1 = s_csamul_cla32_fa19_14_xor0 & s_csamul_cla32_fa19_13_or0;
  assign s_csamul_cla32_fa19_14_or0 = s_csamul_cla32_fa19_14_and0 | s_csamul_cla32_fa19_14_and1;
  assign s_csamul_cla32_and20_14 = a[20] & b[14];
  assign s_csamul_cla32_fa20_14_xor0 = s_csamul_cla32_and20_14 ^ s_csamul_cla32_fa21_13_xor1;
  assign s_csamul_cla32_fa20_14_and0 = s_csamul_cla32_and20_14 & s_csamul_cla32_fa21_13_xor1;
  assign s_csamul_cla32_fa20_14_xor1 = s_csamul_cla32_fa20_14_xor0 ^ s_csamul_cla32_fa20_13_or0;
  assign s_csamul_cla32_fa20_14_and1 = s_csamul_cla32_fa20_14_xor0 & s_csamul_cla32_fa20_13_or0;
  assign s_csamul_cla32_fa20_14_or0 = s_csamul_cla32_fa20_14_and0 | s_csamul_cla32_fa20_14_and1;
  assign s_csamul_cla32_and21_14 = a[21] & b[14];
  assign s_csamul_cla32_fa21_14_xor0 = s_csamul_cla32_and21_14 ^ s_csamul_cla32_fa22_13_xor1;
  assign s_csamul_cla32_fa21_14_and0 = s_csamul_cla32_and21_14 & s_csamul_cla32_fa22_13_xor1;
  assign s_csamul_cla32_fa21_14_xor1 = s_csamul_cla32_fa21_14_xor0 ^ s_csamul_cla32_fa21_13_or0;
  assign s_csamul_cla32_fa21_14_and1 = s_csamul_cla32_fa21_14_xor0 & s_csamul_cla32_fa21_13_or0;
  assign s_csamul_cla32_fa21_14_or0 = s_csamul_cla32_fa21_14_and0 | s_csamul_cla32_fa21_14_and1;
  assign s_csamul_cla32_and22_14 = a[22] & b[14];
  assign s_csamul_cla32_fa22_14_xor0 = s_csamul_cla32_and22_14 ^ s_csamul_cla32_fa23_13_xor1;
  assign s_csamul_cla32_fa22_14_and0 = s_csamul_cla32_and22_14 & s_csamul_cla32_fa23_13_xor1;
  assign s_csamul_cla32_fa22_14_xor1 = s_csamul_cla32_fa22_14_xor0 ^ s_csamul_cla32_fa22_13_or0;
  assign s_csamul_cla32_fa22_14_and1 = s_csamul_cla32_fa22_14_xor0 & s_csamul_cla32_fa22_13_or0;
  assign s_csamul_cla32_fa22_14_or0 = s_csamul_cla32_fa22_14_and0 | s_csamul_cla32_fa22_14_and1;
  assign s_csamul_cla32_and23_14 = a[23] & b[14];
  assign s_csamul_cla32_fa23_14_xor0 = s_csamul_cla32_and23_14 ^ s_csamul_cla32_fa24_13_xor1;
  assign s_csamul_cla32_fa23_14_and0 = s_csamul_cla32_and23_14 & s_csamul_cla32_fa24_13_xor1;
  assign s_csamul_cla32_fa23_14_xor1 = s_csamul_cla32_fa23_14_xor0 ^ s_csamul_cla32_fa23_13_or0;
  assign s_csamul_cla32_fa23_14_and1 = s_csamul_cla32_fa23_14_xor0 & s_csamul_cla32_fa23_13_or0;
  assign s_csamul_cla32_fa23_14_or0 = s_csamul_cla32_fa23_14_and0 | s_csamul_cla32_fa23_14_and1;
  assign s_csamul_cla32_and24_14 = a[24] & b[14];
  assign s_csamul_cla32_fa24_14_xor0 = s_csamul_cla32_and24_14 ^ s_csamul_cla32_fa25_13_xor1;
  assign s_csamul_cla32_fa24_14_and0 = s_csamul_cla32_and24_14 & s_csamul_cla32_fa25_13_xor1;
  assign s_csamul_cla32_fa24_14_xor1 = s_csamul_cla32_fa24_14_xor0 ^ s_csamul_cla32_fa24_13_or0;
  assign s_csamul_cla32_fa24_14_and1 = s_csamul_cla32_fa24_14_xor0 & s_csamul_cla32_fa24_13_or0;
  assign s_csamul_cla32_fa24_14_or0 = s_csamul_cla32_fa24_14_and0 | s_csamul_cla32_fa24_14_and1;
  assign s_csamul_cla32_and25_14 = a[25] & b[14];
  assign s_csamul_cla32_fa25_14_xor0 = s_csamul_cla32_and25_14 ^ s_csamul_cla32_fa26_13_xor1;
  assign s_csamul_cla32_fa25_14_and0 = s_csamul_cla32_and25_14 & s_csamul_cla32_fa26_13_xor1;
  assign s_csamul_cla32_fa25_14_xor1 = s_csamul_cla32_fa25_14_xor0 ^ s_csamul_cla32_fa25_13_or0;
  assign s_csamul_cla32_fa25_14_and1 = s_csamul_cla32_fa25_14_xor0 & s_csamul_cla32_fa25_13_or0;
  assign s_csamul_cla32_fa25_14_or0 = s_csamul_cla32_fa25_14_and0 | s_csamul_cla32_fa25_14_and1;
  assign s_csamul_cla32_and26_14 = a[26] & b[14];
  assign s_csamul_cla32_fa26_14_xor0 = s_csamul_cla32_and26_14 ^ s_csamul_cla32_fa27_13_xor1;
  assign s_csamul_cla32_fa26_14_and0 = s_csamul_cla32_and26_14 & s_csamul_cla32_fa27_13_xor1;
  assign s_csamul_cla32_fa26_14_xor1 = s_csamul_cla32_fa26_14_xor0 ^ s_csamul_cla32_fa26_13_or0;
  assign s_csamul_cla32_fa26_14_and1 = s_csamul_cla32_fa26_14_xor0 & s_csamul_cla32_fa26_13_or0;
  assign s_csamul_cla32_fa26_14_or0 = s_csamul_cla32_fa26_14_and0 | s_csamul_cla32_fa26_14_and1;
  assign s_csamul_cla32_and27_14 = a[27] & b[14];
  assign s_csamul_cla32_fa27_14_xor0 = s_csamul_cla32_and27_14 ^ s_csamul_cla32_fa28_13_xor1;
  assign s_csamul_cla32_fa27_14_and0 = s_csamul_cla32_and27_14 & s_csamul_cla32_fa28_13_xor1;
  assign s_csamul_cla32_fa27_14_xor1 = s_csamul_cla32_fa27_14_xor0 ^ s_csamul_cla32_fa27_13_or0;
  assign s_csamul_cla32_fa27_14_and1 = s_csamul_cla32_fa27_14_xor0 & s_csamul_cla32_fa27_13_or0;
  assign s_csamul_cla32_fa27_14_or0 = s_csamul_cla32_fa27_14_and0 | s_csamul_cla32_fa27_14_and1;
  assign s_csamul_cla32_and28_14 = a[28] & b[14];
  assign s_csamul_cla32_fa28_14_xor0 = s_csamul_cla32_and28_14 ^ s_csamul_cla32_fa29_13_xor1;
  assign s_csamul_cla32_fa28_14_and0 = s_csamul_cla32_and28_14 & s_csamul_cla32_fa29_13_xor1;
  assign s_csamul_cla32_fa28_14_xor1 = s_csamul_cla32_fa28_14_xor0 ^ s_csamul_cla32_fa28_13_or0;
  assign s_csamul_cla32_fa28_14_and1 = s_csamul_cla32_fa28_14_xor0 & s_csamul_cla32_fa28_13_or0;
  assign s_csamul_cla32_fa28_14_or0 = s_csamul_cla32_fa28_14_and0 | s_csamul_cla32_fa28_14_and1;
  assign s_csamul_cla32_and29_14 = a[29] & b[14];
  assign s_csamul_cla32_fa29_14_xor0 = s_csamul_cla32_and29_14 ^ s_csamul_cla32_fa30_13_xor1;
  assign s_csamul_cla32_fa29_14_and0 = s_csamul_cla32_and29_14 & s_csamul_cla32_fa30_13_xor1;
  assign s_csamul_cla32_fa29_14_xor1 = s_csamul_cla32_fa29_14_xor0 ^ s_csamul_cla32_fa29_13_or0;
  assign s_csamul_cla32_fa29_14_and1 = s_csamul_cla32_fa29_14_xor0 & s_csamul_cla32_fa29_13_or0;
  assign s_csamul_cla32_fa29_14_or0 = s_csamul_cla32_fa29_14_and0 | s_csamul_cla32_fa29_14_and1;
  assign s_csamul_cla32_and30_14 = a[30] & b[14];
  assign s_csamul_cla32_fa30_14_xor0 = s_csamul_cla32_and30_14 ^ s_csamul_cla32_ha31_13_xor0;
  assign s_csamul_cla32_fa30_14_and0 = s_csamul_cla32_and30_14 & s_csamul_cla32_ha31_13_xor0;
  assign s_csamul_cla32_fa30_14_xor1 = s_csamul_cla32_fa30_14_xor0 ^ s_csamul_cla32_fa30_13_or0;
  assign s_csamul_cla32_fa30_14_and1 = s_csamul_cla32_fa30_14_xor0 & s_csamul_cla32_fa30_13_or0;
  assign s_csamul_cla32_fa30_14_or0 = s_csamul_cla32_fa30_14_and0 | s_csamul_cla32_fa30_14_and1;
  assign s_csamul_cla32_nand31_14 = ~(a[31] & b[14]);
  assign s_csamul_cla32_ha31_14_xor0 = s_csamul_cla32_nand31_14 ^ s_csamul_cla32_ha31_13_and0;
  assign s_csamul_cla32_ha31_14_and0 = s_csamul_cla32_nand31_14 & s_csamul_cla32_ha31_13_and0;
  assign s_csamul_cla32_and0_15 = a[0] & b[15];
  assign s_csamul_cla32_fa0_15_xor0 = s_csamul_cla32_and0_15 ^ s_csamul_cla32_fa1_14_xor1;
  assign s_csamul_cla32_fa0_15_and0 = s_csamul_cla32_and0_15 & s_csamul_cla32_fa1_14_xor1;
  assign s_csamul_cla32_fa0_15_xor1 = s_csamul_cla32_fa0_15_xor0 ^ s_csamul_cla32_fa0_14_or0;
  assign s_csamul_cla32_fa0_15_and1 = s_csamul_cla32_fa0_15_xor0 & s_csamul_cla32_fa0_14_or0;
  assign s_csamul_cla32_fa0_15_or0 = s_csamul_cla32_fa0_15_and0 | s_csamul_cla32_fa0_15_and1;
  assign s_csamul_cla32_and1_15 = a[1] & b[15];
  assign s_csamul_cla32_fa1_15_xor0 = s_csamul_cla32_and1_15 ^ s_csamul_cla32_fa2_14_xor1;
  assign s_csamul_cla32_fa1_15_and0 = s_csamul_cla32_and1_15 & s_csamul_cla32_fa2_14_xor1;
  assign s_csamul_cla32_fa1_15_xor1 = s_csamul_cla32_fa1_15_xor0 ^ s_csamul_cla32_fa1_14_or0;
  assign s_csamul_cla32_fa1_15_and1 = s_csamul_cla32_fa1_15_xor0 & s_csamul_cla32_fa1_14_or0;
  assign s_csamul_cla32_fa1_15_or0 = s_csamul_cla32_fa1_15_and0 | s_csamul_cla32_fa1_15_and1;
  assign s_csamul_cla32_and2_15 = a[2] & b[15];
  assign s_csamul_cla32_fa2_15_xor0 = s_csamul_cla32_and2_15 ^ s_csamul_cla32_fa3_14_xor1;
  assign s_csamul_cla32_fa2_15_and0 = s_csamul_cla32_and2_15 & s_csamul_cla32_fa3_14_xor1;
  assign s_csamul_cla32_fa2_15_xor1 = s_csamul_cla32_fa2_15_xor0 ^ s_csamul_cla32_fa2_14_or0;
  assign s_csamul_cla32_fa2_15_and1 = s_csamul_cla32_fa2_15_xor0 & s_csamul_cla32_fa2_14_or0;
  assign s_csamul_cla32_fa2_15_or0 = s_csamul_cla32_fa2_15_and0 | s_csamul_cla32_fa2_15_and1;
  assign s_csamul_cla32_and3_15 = a[3] & b[15];
  assign s_csamul_cla32_fa3_15_xor0 = s_csamul_cla32_and3_15 ^ s_csamul_cla32_fa4_14_xor1;
  assign s_csamul_cla32_fa3_15_and0 = s_csamul_cla32_and3_15 & s_csamul_cla32_fa4_14_xor1;
  assign s_csamul_cla32_fa3_15_xor1 = s_csamul_cla32_fa3_15_xor0 ^ s_csamul_cla32_fa3_14_or0;
  assign s_csamul_cla32_fa3_15_and1 = s_csamul_cla32_fa3_15_xor0 & s_csamul_cla32_fa3_14_or0;
  assign s_csamul_cla32_fa3_15_or0 = s_csamul_cla32_fa3_15_and0 | s_csamul_cla32_fa3_15_and1;
  assign s_csamul_cla32_and4_15 = a[4] & b[15];
  assign s_csamul_cla32_fa4_15_xor0 = s_csamul_cla32_and4_15 ^ s_csamul_cla32_fa5_14_xor1;
  assign s_csamul_cla32_fa4_15_and0 = s_csamul_cla32_and4_15 & s_csamul_cla32_fa5_14_xor1;
  assign s_csamul_cla32_fa4_15_xor1 = s_csamul_cla32_fa4_15_xor0 ^ s_csamul_cla32_fa4_14_or0;
  assign s_csamul_cla32_fa4_15_and1 = s_csamul_cla32_fa4_15_xor0 & s_csamul_cla32_fa4_14_or0;
  assign s_csamul_cla32_fa4_15_or0 = s_csamul_cla32_fa4_15_and0 | s_csamul_cla32_fa4_15_and1;
  assign s_csamul_cla32_and5_15 = a[5] & b[15];
  assign s_csamul_cla32_fa5_15_xor0 = s_csamul_cla32_and5_15 ^ s_csamul_cla32_fa6_14_xor1;
  assign s_csamul_cla32_fa5_15_and0 = s_csamul_cla32_and5_15 & s_csamul_cla32_fa6_14_xor1;
  assign s_csamul_cla32_fa5_15_xor1 = s_csamul_cla32_fa5_15_xor0 ^ s_csamul_cla32_fa5_14_or0;
  assign s_csamul_cla32_fa5_15_and1 = s_csamul_cla32_fa5_15_xor0 & s_csamul_cla32_fa5_14_or0;
  assign s_csamul_cla32_fa5_15_or0 = s_csamul_cla32_fa5_15_and0 | s_csamul_cla32_fa5_15_and1;
  assign s_csamul_cla32_and6_15 = a[6] & b[15];
  assign s_csamul_cla32_fa6_15_xor0 = s_csamul_cla32_and6_15 ^ s_csamul_cla32_fa7_14_xor1;
  assign s_csamul_cla32_fa6_15_and0 = s_csamul_cla32_and6_15 & s_csamul_cla32_fa7_14_xor1;
  assign s_csamul_cla32_fa6_15_xor1 = s_csamul_cla32_fa6_15_xor0 ^ s_csamul_cla32_fa6_14_or0;
  assign s_csamul_cla32_fa6_15_and1 = s_csamul_cla32_fa6_15_xor0 & s_csamul_cla32_fa6_14_or0;
  assign s_csamul_cla32_fa6_15_or0 = s_csamul_cla32_fa6_15_and0 | s_csamul_cla32_fa6_15_and1;
  assign s_csamul_cla32_and7_15 = a[7] & b[15];
  assign s_csamul_cla32_fa7_15_xor0 = s_csamul_cla32_and7_15 ^ s_csamul_cla32_fa8_14_xor1;
  assign s_csamul_cla32_fa7_15_and0 = s_csamul_cla32_and7_15 & s_csamul_cla32_fa8_14_xor1;
  assign s_csamul_cla32_fa7_15_xor1 = s_csamul_cla32_fa7_15_xor0 ^ s_csamul_cla32_fa7_14_or0;
  assign s_csamul_cla32_fa7_15_and1 = s_csamul_cla32_fa7_15_xor0 & s_csamul_cla32_fa7_14_or0;
  assign s_csamul_cla32_fa7_15_or0 = s_csamul_cla32_fa7_15_and0 | s_csamul_cla32_fa7_15_and1;
  assign s_csamul_cla32_and8_15 = a[8] & b[15];
  assign s_csamul_cla32_fa8_15_xor0 = s_csamul_cla32_and8_15 ^ s_csamul_cla32_fa9_14_xor1;
  assign s_csamul_cla32_fa8_15_and0 = s_csamul_cla32_and8_15 & s_csamul_cla32_fa9_14_xor1;
  assign s_csamul_cla32_fa8_15_xor1 = s_csamul_cla32_fa8_15_xor0 ^ s_csamul_cla32_fa8_14_or0;
  assign s_csamul_cla32_fa8_15_and1 = s_csamul_cla32_fa8_15_xor0 & s_csamul_cla32_fa8_14_or0;
  assign s_csamul_cla32_fa8_15_or0 = s_csamul_cla32_fa8_15_and0 | s_csamul_cla32_fa8_15_and1;
  assign s_csamul_cla32_and9_15 = a[9] & b[15];
  assign s_csamul_cla32_fa9_15_xor0 = s_csamul_cla32_and9_15 ^ s_csamul_cla32_fa10_14_xor1;
  assign s_csamul_cla32_fa9_15_and0 = s_csamul_cla32_and9_15 & s_csamul_cla32_fa10_14_xor1;
  assign s_csamul_cla32_fa9_15_xor1 = s_csamul_cla32_fa9_15_xor0 ^ s_csamul_cla32_fa9_14_or0;
  assign s_csamul_cla32_fa9_15_and1 = s_csamul_cla32_fa9_15_xor0 & s_csamul_cla32_fa9_14_or0;
  assign s_csamul_cla32_fa9_15_or0 = s_csamul_cla32_fa9_15_and0 | s_csamul_cla32_fa9_15_and1;
  assign s_csamul_cla32_and10_15 = a[10] & b[15];
  assign s_csamul_cla32_fa10_15_xor0 = s_csamul_cla32_and10_15 ^ s_csamul_cla32_fa11_14_xor1;
  assign s_csamul_cla32_fa10_15_and0 = s_csamul_cla32_and10_15 & s_csamul_cla32_fa11_14_xor1;
  assign s_csamul_cla32_fa10_15_xor1 = s_csamul_cla32_fa10_15_xor0 ^ s_csamul_cla32_fa10_14_or0;
  assign s_csamul_cla32_fa10_15_and1 = s_csamul_cla32_fa10_15_xor0 & s_csamul_cla32_fa10_14_or0;
  assign s_csamul_cla32_fa10_15_or0 = s_csamul_cla32_fa10_15_and0 | s_csamul_cla32_fa10_15_and1;
  assign s_csamul_cla32_and11_15 = a[11] & b[15];
  assign s_csamul_cla32_fa11_15_xor0 = s_csamul_cla32_and11_15 ^ s_csamul_cla32_fa12_14_xor1;
  assign s_csamul_cla32_fa11_15_and0 = s_csamul_cla32_and11_15 & s_csamul_cla32_fa12_14_xor1;
  assign s_csamul_cla32_fa11_15_xor1 = s_csamul_cla32_fa11_15_xor0 ^ s_csamul_cla32_fa11_14_or0;
  assign s_csamul_cla32_fa11_15_and1 = s_csamul_cla32_fa11_15_xor0 & s_csamul_cla32_fa11_14_or0;
  assign s_csamul_cla32_fa11_15_or0 = s_csamul_cla32_fa11_15_and0 | s_csamul_cla32_fa11_15_and1;
  assign s_csamul_cla32_and12_15 = a[12] & b[15];
  assign s_csamul_cla32_fa12_15_xor0 = s_csamul_cla32_and12_15 ^ s_csamul_cla32_fa13_14_xor1;
  assign s_csamul_cla32_fa12_15_and0 = s_csamul_cla32_and12_15 & s_csamul_cla32_fa13_14_xor1;
  assign s_csamul_cla32_fa12_15_xor1 = s_csamul_cla32_fa12_15_xor0 ^ s_csamul_cla32_fa12_14_or0;
  assign s_csamul_cla32_fa12_15_and1 = s_csamul_cla32_fa12_15_xor0 & s_csamul_cla32_fa12_14_or0;
  assign s_csamul_cla32_fa12_15_or0 = s_csamul_cla32_fa12_15_and0 | s_csamul_cla32_fa12_15_and1;
  assign s_csamul_cla32_and13_15 = a[13] & b[15];
  assign s_csamul_cla32_fa13_15_xor0 = s_csamul_cla32_and13_15 ^ s_csamul_cla32_fa14_14_xor1;
  assign s_csamul_cla32_fa13_15_and0 = s_csamul_cla32_and13_15 & s_csamul_cla32_fa14_14_xor1;
  assign s_csamul_cla32_fa13_15_xor1 = s_csamul_cla32_fa13_15_xor0 ^ s_csamul_cla32_fa13_14_or0;
  assign s_csamul_cla32_fa13_15_and1 = s_csamul_cla32_fa13_15_xor0 & s_csamul_cla32_fa13_14_or0;
  assign s_csamul_cla32_fa13_15_or0 = s_csamul_cla32_fa13_15_and0 | s_csamul_cla32_fa13_15_and1;
  assign s_csamul_cla32_and14_15 = a[14] & b[15];
  assign s_csamul_cla32_fa14_15_xor0 = s_csamul_cla32_and14_15 ^ s_csamul_cla32_fa15_14_xor1;
  assign s_csamul_cla32_fa14_15_and0 = s_csamul_cla32_and14_15 & s_csamul_cla32_fa15_14_xor1;
  assign s_csamul_cla32_fa14_15_xor1 = s_csamul_cla32_fa14_15_xor0 ^ s_csamul_cla32_fa14_14_or0;
  assign s_csamul_cla32_fa14_15_and1 = s_csamul_cla32_fa14_15_xor0 & s_csamul_cla32_fa14_14_or0;
  assign s_csamul_cla32_fa14_15_or0 = s_csamul_cla32_fa14_15_and0 | s_csamul_cla32_fa14_15_and1;
  assign s_csamul_cla32_and15_15 = a[15] & b[15];
  assign s_csamul_cla32_fa15_15_xor0 = s_csamul_cla32_and15_15 ^ s_csamul_cla32_fa16_14_xor1;
  assign s_csamul_cla32_fa15_15_and0 = s_csamul_cla32_and15_15 & s_csamul_cla32_fa16_14_xor1;
  assign s_csamul_cla32_fa15_15_xor1 = s_csamul_cla32_fa15_15_xor0 ^ s_csamul_cla32_fa15_14_or0;
  assign s_csamul_cla32_fa15_15_and1 = s_csamul_cla32_fa15_15_xor0 & s_csamul_cla32_fa15_14_or0;
  assign s_csamul_cla32_fa15_15_or0 = s_csamul_cla32_fa15_15_and0 | s_csamul_cla32_fa15_15_and1;
  assign s_csamul_cla32_and16_15 = a[16] & b[15];
  assign s_csamul_cla32_fa16_15_xor0 = s_csamul_cla32_and16_15 ^ s_csamul_cla32_fa17_14_xor1;
  assign s_csamul_cla32_fa16_15_and0 = s_csamul_cla32_and16_15 & s_csamul_cla32_fa17_14_xor1;
  assign s_csamul_cla32_fa16_15_xor1 = s_csamul_cla32_fa16_15_xor0 ^ s_csamul_cla32_fa16_14_or0;
  assign s_csamul_cla32_fa16_15_and1 = s_csamul_cla32_fa16_15_xor0 & s_csamul_cla32_fa16_14_or0;
  assign s_csamul_cla32_fa16_15_or0 = s_csamul_cla32_fa16_15_and0 | s_csamul_cla32_fa16_15_and1;
  assign s_csamul_cla32_and17_15 = a[17] & b[15];
  assign s_csamul_cla32_fa17_15_xor0 = s_csamul_cla32_and17_15 ^ s_csamul_cla32_fa18_14_xor1;
  assign s_csamul_cla32_fa17_15_and0 = s_csamul_cla32_and17_15 & s_csamul_cla32_fa18_14_xor1;
  assign s_csamul_cla32_fa17_15_xor1 = s_csamul_cla32_fa17_15_xor0 ^ s_csamul_cla32_fa17_14_or0;
  assign s_csamul_cla32_fa17_15_and1 = s_csamul_cla32_fa17_15_xor0 & s_csamul_cla32_fa17_14_or0;
  assign s_csamul_cla32_fa17_15_or0 = s_csamul_cla32_fa17_15_and0 | s_csamul_cla32_fa17_15_and1;
  assign s_csamul_cla32_and18_15 = a[18] & b[15];
  assign s_csamul_cla32_fa18_15_xor0 = s_csamul_cla32_and18_15 ^ s_csamul_cla32_fa19_14_xor1;
  assign s_csamul_cla32_fa18_15_and0 = s_csamul_cla32_and18_15 & s_csamul_cla32_fa19_14_xor1;
  assign s_csamul_cla32_fa18_15_xor1 = s_csamul_cla32_fa18_15_xor0 ^ s_csamul_cla32_fa18_14_or0;
  assign s_csamul_cla32_fa18_15_and1 = s_csamul_cla32_fa18_15_xor0 & s_csamul_cla32_fa18_14_or0;
  assign s_csamul_cla32_fa18_15_or0 = s_csamul_cla32_fa18_15_and0 | s_csamul_cla32_fa18_15_and1;
  assign s_csamul_cla32_and19_15 = a[19] & b[15];
  assign s_csamul_cla32_fa19_15_xor0 = s_csamul_cla32_and19_15 ^ s_csamul_cla32_fa20_14_xor1;
  assign s_csamul_cla32_fa19_15_and0 = s_csamul_cla32_and19_15 & s_csamul_cla32_fa20_14_xor1;
  assign s_csamul_cla32_fa19_15_xor1 = s_csamul_cla32_fa19_15_xor0 ^ s_csamul_cla32_fa19_14_or0;
  assign s_csamul_cla32_fa19_15_and1 = s_csamul_cla32_fa19_15_xor0 & s_csamul_cla32_fa19_14_or0;
  assign s_csamul_cla32_fa19_15_or0 = s_csamul_cla32_fa19_15_and0 | s_csamul_cla32_fa19_15_and1;
  assign s_csamul_cla32_and20_15 = a[20] & b[15];
  assign s_csamul_cla32_fa20_15_xor0 = s_csamul_cla32_and20_15 ^ s_csamul_cla32_fa21_14_xor1;
  assign s_csamul_cla32_fa20_15_and0 = s_csamul_cla32_and20_15 & s_csamul_cla32_fa21_14_xor1;
  assign s_csamul_cla32_fa20_15_xor1 = s_csamul_cla32_fa20_15_xor0 ^ s_csamul_cla32_fa20_14_or0;
  assign s_csamul_cla32_fa20_15_and1 = s_csamul_cla32_fa20_15_xor0 & s_csamul_cla32_fa20_14_or0;
  assign s_csamul_cla32_fa20_15_or0 = s_csamul_cla32_fa20_15_and0 | s_csamul_cla32_fa20_15_and1;
  assign s_csamul_cla32_and21_15 = a[21] & b[15];
  assign s_csamul_cla32_fa21_15_xor0 = s_csamul_cla32_and21_15 ^ s_csamul_cla32_fa22_14_xor1;
  assign s_csamul_cla32_fa21_15_and0 = s_csamul_cla32_and21_15 & s_csamul_cla32_fa22_14_xor1;
  assign s_csamul_cla32_fa21_15_xor1 = s_csamul_cla32_fa21_15_xor0 ^ s_csamul_cla32_fa21_14_or0;
  assign s_csamul_cla32_fa21_15_and1 = s_csamul_cla32_fa21_15_xor0 & s_csamul_cla32_fa21_14_or0;
  assign s_csamul_cla32_fa21_15_or0 = s_csamul_cla32_fa21_15_and0 | s_csamul_cla32_fa21_15_and1;
  assign s_csamul_cla32_and22_15 = a[22] & b[15];
  assign s_csamul_cla32_fa22_15_xor0 = s_csamul_cla32_and22_15 ^ s_csamul_cla32_fa23_14_xor1;
  assign s_csamul_cla32_fa22_15_and0 = s_csamul_cla32_and22_15 & s_csamul_cla32_fa23_14_xor1;
  assign s_csamul_cla32_fa22_15_xor1 = s_csamul_cla32_fa22_15_xor0 ^ s_csamul_cla32_fa22_14_or0;
  assign s_csamul_cla32_fa22_15_and1 = s_csamul_cla32_fa22_15_xor0 & s_csamul_cla32_fa22_14_or0;
  assign s_csamul_cla32_fa22_15_or0 = s_csamul_cla32_fa22_15_and0 | s_csamul_cla32_fa22_15_and1;
  assign s_csamul_cla32_and23_15 = a[23] & b[15];
  assign s_csamul_cla32_fa23_15_xor0 = s_csamul_cla32_and23_15 ^ s_csamul_cla32_fa24_14_xor1;
  assign s_csamul_cla32_fa23_15_and0 = s_csamul_cla32_and23_15 & s_csamul_cla32_fa24_14_xor1;
  assign s_csamul_cla32_fa23_15_xor1 = s_csamul_cla32_fa23_15_xor0 ^ s_csamul_cla32_fa23_14_or0;
  assign s_csamul_cla32_fa23_15_and1 = s_csamul_cla32_fa23_15_xor0 & s_csamul_cla32_fa23_14_or0;
  assign s_csamul_cla32_fa23_15_or0 = s_csamul_cla32_fa23_15_and0 | s_csamul_cla32_fa23_15_and1;
  assign s_csamul_cla32_and24_15 = a[24] & b[15];
  assign s_csamul_cla32_fa24_15_xor0 = s_csamul_cla32_and24_15 ^ s_csamul_cla32_fa25_14_xor1;
  assign s_csamul_cla32_fa24_15_and0 = s_csamul_cla32_and24_15 & s_csamul_cla32_fa25_14_xor1;
  assign s_csamul_cla32_fa24_15_xor1 = s_csamul_cla32_fa24_15_xor0 ^ s_csamul_cla32_fa24_14_or0;
  assign s_csamul_cla32_fa24_15_and1 = s_csamul_cla32_fa24_15_xor0 & s_csamul_cla32_fa24_14_or0;
  assign s_csamul_cla32_fa24_15_or0 = s_csamul_cla32_fa24_15_and0 | s_csamul_cla32_fa24_15_and1;
  assign s_csamul_cla32_and25_15 = a[25] & b[15];
  assign s_csamul_cla32_fa25_15_xor0 = s_csamul_cla32_and25_15 ^ s_csamul_cla32_fa26_14_xor1;
  assign s_csamul_cla32_fa25_15_and0 = s_csamul_cla32_and25_15 & s_csamul_cla32_fa26_14_xor1;
  assign s_csamul_cla32_fa25_15_xor1 = s_csamul_cla32_fa25_15_xor0 ^ s_csamul_cla32_fa25_14_or0;
  assign s_csamul_cla32_fa25_15_and1 = s_csamul_cla32_fa25_15_xor0 & s_csamul_cla32_fa25_14_or0;
  assign s_csamul_cla32_fa25_15_or0 = s_csamul_cla32_fa25_15_and0 | s_csamul_cla32_fa25_15_and1;
  assign s_csamul_cla32_and26_15 = a[26] & b[15];
  assign s_csamul_cla32_fa26_15_xor0 = s_csamul_cla32_and26_15 ^ s_csamul_cla32_fa27_14_xor1;
  assign s_csamul_cla32_fa26_15_and0 = s_csamul_cla32_and26_15 & s_csamul_cla32_fa27_14_xor1;
  assign s_csamul_cla32_fa26_15_xor1 = s_csamul_cla32_fa26_15_xor0 ^ s_csamul_cla32_fa26_14_or0;
  assign s_csamul_cla32_fa26_15_and1 = s_csamul_cla32_fa26_15_xor0 & s_csamul_cla32_fa26_14_or0;
  assign s_csamul_cla32_fa26_15_or0 = s_csamul_cla32_fa26_15_and0 | s_csamul_cla32_fa26_15_and1;
  assign s_csamul_cla32_and27_15 = a[27] & b[15];
  assign s_csamul_cla32_fa27_15_xor0 = s_csamul_cla32_and27_15 ^ s_csamul_cla32_fa28_14_xor1;
  assign s_csamul_cla32_fa27_15_and0 = s_csamul_cla32_and27_15 & s_csamul_cla32_fa28_14_xor1;
  assign s_csamul_cla32_fa27_15_xor1 = s_csamul_cla32_fa27_15_xor0 ^ s_csamul_cla32_fa27_14_or0;
  assign s_csamul_cla32_fa27_15_and1 = s_csamul_cla32_fa27_15_xor0 & s_csamul_cla32_fa27_14_or0;
  assign s_csamul_cla32_fa27_15_or0 = s_csamul_cla32_fa27_15_and0 | s_csamul_cla32_fa27_15_and1;
  assign s_csamul_cla32_and28_15 = a[28] & b[15];
  assign s_csamul_cla32_fa28_15_xor0 = s_csamul_cla32_and28_15 ^ s_csamul_cla32_fa29_14_xor1;
  assign s_csamul_cla32_fa28_15_and0 = s_csamul_cla32_and28_15 & s_csamul_cla32_fa29_14_xor1;
  assign s_csamul_cla32_fa28_15_xor1 = s_csamul_cla32_fa28_15_xor0 ^ s_csamul_cla32_fa28_14_or0;
  assign s_csamul_cla32_fa28_15_and1 = s_csamul_cla32_fa28_15_xor0 & s_csamul_cla32_fa28_14_or0;
  assign s_csamul_cla32_fa28_15_or0 = s_csamul_cla32_fa28_15_and0 | s_csamul_cla32_fa28_15_and1;
  assign s_csamul_cla32_and29_15 = a[29] & b[15];
  assign s_csamul_cla32_fa29_15_xor0 = s_csamul_cla32_and29_15 ^ s_csamul_cla32_fa30_14_xor1;
  assign s_csamul_cla32_fa29_15_and0 = s_csamul_cla32_and29_15 & s_csamul_cla32_fa30_14_xor1;
  assign s_csamul_cla32_fa29_15_xor1 = s_csamul_cla32_fa29_15_xor0 ^ s_csamul_cla32_fa29_14_or0;
  assign s_csamul_cla32_fa29_15_and1 = s_csamul_cla32_fa29_15_xor0 & s_csamul_cla32_fa29_14_or0;
  assign s_csamul_cla32_fa29_15_or0 = s_csamul_cla32_fa29_15_and0 | s_csamul_cla32_fa29_15_and1;
  assign s_csamul_cla32_and30_15 = a[30] & b[15];
  assign s_csamul_cla32_fa30_15_xor0 = s_csamul_cla32_and30_15 ^ s_csamul_cla32_ha31_14_xor0;
  assign s_csamul_cla32_fa30_15_and0 = s_csamul_cla32_and30_15 & s_csamul_cla32_ha31_14_xor0;
  assign s_csamul_cla32_fa30_15_xor1 = s_csamul_cla32_fa30_15_xor0 ^ s_csamul_cla32_fa30_14_or0;
  assign s_csamul_cla32_fa30_15_and1 = s_csamul_cla32_fa30_15_xor0 & s_csamul_cla32_fa30_14_or0;
  assign s_csamul_cla32_fa30_15_or0 = s_csamul_cla32_fa30_15_and0 | s_csamul_cla32_fa30_15_and1;
  assign s_csamul_cla32_nand31_15 = ~(a[31] & b[15]);
  assign s_csamul_cla32_ha31_15_xor0 = s_csamul_cla32_nand31_15 ^ s_csamul_cla32_ha31_14_and0;
  assign s_csamul_cla32_ha31_15_and0 = s_csamul_cla32_nand31_15 & s_csamul_cla32_ha31_14_and0;
  assign s_csamul_cla32_and0_16 = a[0] & b[16];
  assign s_csamul_cla32_fa0_16_xor0 = s_csamul_cla32_and0_16 ^ s_csamul_cla32_fa1_15_xor1;
  assign s_csamul_cla32_fa0_16_and0 = s_csamul_cla32_and0_16 & s_csamul_cla32_fa1_15_xor1;
  assign s_csamul_cla32_fa0_16_xor1 = s_csamul_cla32_fa0_16_xor0 ^ s_csamul_cla32_fa0_15_or0;
  assign s_csamul_cla32_fa0_16_and1 = s_csamul_cla32_fa0_16_xor0 & s_csamul_cla32_fa0_15_or0;
  assign s_csamul_cla32_fa0_16_or0 = s_csamul_cla32_fa0_16_and0 | s_csamul_cla32_fa0_16_and1;
  assign s_csamul_cla32_and1_16 = a[1] & b[16];
  assign s_csamul_cla32_fa1_16_xor0 = s_csamul_cla32_and1_16 ^ s_csamul_cla32_fa2_15_xor1;
  assign s_csamul_cla32_fa1_16_and0 = s_csamul_cla32_and1_16 & s_csamul_cla32_fa2_15_xor1;
  assign s_csamul_cla32_fa1_16_xor1 = s_csamul_cla32_fa1_16_xor0 ^ s_csamul_cla32_fa1_15_or0;
  assign s_csamul_cla32_fa1_16_and1 = s_csamul_cla32_fa1_16_xor0 & s_csamul_cla32_fa1_15_or0;
  assign s_csamul_cla32_fa1_16_or0 = s_csamul_cla32_fa1_16_and0 | s_csamul_cla32_fa1_16_and1;
  assign s_csamul_cla32_and2_16 = a[2] & b[16];
  assign s_csamul_cla32_fa2_16_xor0 = s_csamul_cla32_and2_16 ^ s_csamul_cla32_fa3_15_xor1;
  assign s_csamul_cla32_fa2_16_and0 = s_csamul_cla32_and2_16 & s_csamul_cla32_fa3_15_xor1;
  assign s_csamul_cla32_fa2_16_xor1 = s_csamul_cla32_fa2_16_xor0 ^ s_csamul_cla32_fa2_15_or0;
  assign s_csamul_cla32_fa2_16_and1 = s_csamul_cla32_fa2_16_xor0 & s_csamul_cla32_fa2_15_or0;
  assign s_csamul_cla32_fa2_16_or0 = s_csamul_cla32_fa2_16_and0 | s_csamul_cla32_fa2_16_and1;
  assign s_csamul_cla32_and3_16 = a[3] & b[16];
  assign s_csamul_cla32_fa3_16_xor0 = s_csamul_cla32_and3_16 ^ s_csamul_cla32_fa4_15_xor1;
  assign s_csamul_cla32_fa3_16_and0 = s_csamul_cla32_and3_16 & s_csamul_cla32_fa4_15_xor1;
  assign s_csamul_cla32_fa3_16_xor1 = s_csamul_cla32_fa3_16_xor0 ^ s_csamul_cla32_fa3_15_or0;
  assign s_csamul_cla32_fa3_16_and1 = s_csamul_cla32_fa3_16_xor0 & s_csamul_cla32_fa3_15_or0;
  assign s_csamul_cla32_fa3_16_or0 = s_csamul_cla32_fa3_16_and0 | s_csamul_cla32_fa3_16_and1;
  assign s_csamul_cla32_and4_16 = a[4] & b[16];
  assign s_csamul_cla32_fa4_16_xor0 = s_csamul_cla32_and4_16 ^ s_csamul_cla32_fa5_15_xor1;
  assign s_csamul_cla32_fa4_16_and0 = s_csamul_cla32_and4_16 & s_csamul_cla32_fa5_15_xor1;
  assign s_csamul_cla32_fa4_16_xor1 = s_csamul_cla32_fa4_16_xor0 ^ s_csamul_cla32_fa4_15_or0;
  assign s_csamul_cla32_fa4_16_and1 = s_csamul_cla32_fa4_16_xor0 & s_csamul_cla32_fa4_15_or0;
  assign s_csamul_cla32_fa4_16_or0 = s_csamul_cla32_fa4_16_and0 | s_csamul_cla32_fa4_16_and1;
  assign s_csamul_cla32_and5_16 = a[5] & b[16];
  assign s_csamul_cla32_fa5_16_xor0 = s_csamul_cla32_and5_16 ^ s_csamul_cla32_fa6_15_xor1;
  assign s_csamul_cla32_fa5_16_and0 = s_csamul_cla32_and5_16 & s_csamul_cla32_fa6_15_xor1;
  assign s_csamul_cla32_fa5_16_xor1 = s_csamul_cla32_fa5_16_xor0 ^ s_csamul_cla32_fa5_15_or0;
  assign s_csamul_cla32_fa5_16_and1 = s_csamul_cla32_fa5_16_xor0 & s_csamul_cla32_fa5_15_or0;
  assign s_csamul_cla32_fa5_16_or0 = s_csamul_cla32_fa5_16_and0 | s_csamul_cla32_fa5_16_and1;
  assign s_csamul_cla32_and6_16 = a[6] & b[16];
  assign s_csamul_cla32_fa6_16_xor0 = s_csamul_cla32_and6_16 ^ s_csamul_cla32_fa7_15_xor1;
  assign s_csamul_cla32_fa6_16_and0 = s_csamul_cla32_and6_16 & s_csamul_cla32_fa7_15_xor1;
  assign s_csamul_cla32_fa6_16_xor1 = s_csamul_cla32_fa6_16_xor0 ^ s_csamul_cla32_fa6_15_or0;
  assign s_csamul_cla32_fa6_16_and1 = s_csamul_cla32_fa6_16_xor0 & s_csamul_cla32_fa6_15_or0;
  assign s_csamul_cla32_fa6_16_or0 = s_csamul_cla32_fa6_16_and0 | s_csamul_cla32_fa6_16_and1;
  assign s_csamul_cla32_and7_16 = a[7] & b[16];
  assign s_csamul_cla32_fa7_16_xor0 = s_csamul_cla32_and7_16 ^ s_csamul_cla32_fa8_15_xor1;
  assign s_csamul_cla32_fa7_16_and0 = s_csamul_cla32_and7_16 & s_csamul_cla32_fa8_15_xor1;
  assign s_csamul_cla32_fa7_16_xor1 = s_csamul_cla32_fa7_16_xor0 ^ s_csamul_cla32_fa7_15_or0;
  assign s_csamul_cla32_fa7_16_and1 = s_csamul_cla32_fa7_16_xor0 & s_csamul_cla32_fa7_15_or0;
  assign s_csamul_cla32_fa7_16_or0 = s_csamul_cla32_fa7_16_and0 | s_csamul_cla32_fa7_16_and1;
  assign s_csamul_cla32_and8_16 = a[8] & b[16];
  assign s_csamul_cla32_fa8_16_xor0 = s_csamul_cla32_and8_16 ^ s_csamul_cla32_fa9_15_xor1;
  assign s_csamul_cla32_fa8_16_and0 = s_csamul_cla32_and8_16 & s_csamul_cla32_fa9_15_xor1;
  assign s_csamul_cla32_fa8_16_xor1 = s_csamul_cla32_fa8_16_xor0 ^ s_csamul_cla32_fa8_15_or0;
  assign s_csamul_cla32_fa8_16_and1 = s_csamul_cla32_fa8_16_xor0 & s_csamul_cla32_fa8_15_or0;
  assign s_csamul_cla32_fa8_16_or0 = s_csamul_cla32_fa8_16_and0 | s_csamul_cla32_fa8_16_and1;
  assign s_csamul_cla32_and9_16 = a[9] & b[16];
  assign s_csamul_cla32_fa9_16_xor0 = s_csamul_cla32_and9_16 ^ s_csamul_cla32_fa10_15_xor1;
  assign s_csamul_cla32_fa9_16_and0 = s_csamul_cla32_and9_16 & s_csamul_cla32_fa10_15_xor1;
  assign s_csamul_cla32_fa9_16_xor1 = s_csamul_cla32_fa9_16_xor0 ^ s_csamul_cla32_fa9_15_or0;
  assign s_csamul_cla32_fa9_16_and1 = s_csamul_cla32_fa9_16_xor0 & s_csamul_cla32_fa9_15_or0;
  assign s_csamul_cla32_fa9_16_or0 = s_csamul_cla32_fa9_16_and0 | s_csamul_cla32_fa9_16_and1;
  assign s_csamul_cla32_and10_16 = a[10] & b[16];
  assign s_csamul_cla32_fa10_16_xor0 = s_csamul_cla32_and10_16 ^ s_csamul_cla32_fa11_15_xor1;
  assign s_csamul_cla32_fa10_16_and0 = s_csamul_cla32_and10_16 & s_csamul_cla32_fa11_15_xor1;
  assign s_csamul_cla32_fa10_16_xor1 = s_csamul_cla32_fa10_16_xor0 ^ s_csamul_cla32_fa10_15_or0;
  assign s_csamul_cla32_fa10_16_and1 = s_csamul_cla32_fa10_16_xor0 & s_csamul_cla32_fa10_15_or0;
  assign s_csamul_cla32_fa10_16_or0 = s_csamul_cla32_fa10_16_and0 | s_csamul_cla32_fa10_16_and1;
  assign s_csamul_cla32_and11_16 = a[11] & b[16];
  assign s_csamul_cla32_fa11_16_xor0 = s_csamul_cla32_and11_16 ^ s_csamul_cla32_fa12_15_xor1;
  assign s_csamul_cla32_fa11_16_and0 = s_csamul_cla32_and11_16 & s_csamul_cla32_fa12_15_xor1;
  assign s_csamul_cla32_fa11_16_xor1 = s_csamul_cla32_fa11_16_xor0 ^ s_csamul_cla32_fa11_15_or0;
  assign s_csamul_cla32_fa11_16_and1 = s_csamul_cla32_fa11_16_xor0 & s_csamul_cla32_fa11_15_or0;
  assign s_csamul_cla32_fa11_16_or0 = s_csamul_cla32_fa11_16_and0 | s_csamul_cla32_fa11_16_and1;
  assign s_csamul_cla32_and12_16 = a[12] & b[16];
  assign s_csamul_cla32_fa12_16_xor0 = s_csamul_cla32_and12_16 ^ s_csamul_cla32_fa13_15_xor1;
  assign s_csamul_cla32_fa12_16_and0 = s_csamul_cla32_and12_16 & s_csamul_cla32_fa13_15_xor1;
  assign s_csamul_cla32_fa12_16_xor1 = s_csamul_cla32_fa12_16_xor0 ^ s_csamul_cla32_fa12_15_or0;
  assign s_csamul_cla32_fa12_16_and1 = s_csamul_cla32_fa12_16_xor0 & s_csamul_cla32_fa12_15_or0;
  assign s_csamul_cla32_fa12_16_or0 = s_csamul_cla32_fa12_16_and0 | s_csamul_cla32_fa12_16_and1;
  assign s_csamul_cla32_and13_16 = a[13] & b[16];
  assign s_csamul_cla32_fa13_16_xor0 = s_csamul_cla32_and13_16 ^ s_csamul_cla32_fa14_15_xor1;
  assign s_csamul_cla32_fa13_16_and0 = s_csamul_cla32_and13_16 & s_csamul_cla32_fa14_15_xor1;
  assign s_csamul_cla32_fa13_16_xor1 = s_csamul_cla32_fa13_16_xor0 ^ s_csamul_cla32_fa13_15_or0;
  assign s_csamul_cla32_fa13_16_and1 = s_csamul_cla32_fa13_16_xor0 & s_csamul_cla32_fa13_15_or0;
  assign s_csamul_cla32_fa13_16_or0 = s_csamul_cla32_fa13_16_and0 | s_csamul_cla32_fa13_16_and1;
  assign s_csamul_cla32_and14_16 = a[14] & b[16];
  assign s_csamul_cla32_fa14_16_xor0 = s_csamul_cla32_and14_16 ^ s_csamul_cla32_fa15_15_xor1;
  assign s_csamul_cla32_fa14_16_and0 = s_csamul_cla32_and14_16 & s_csamul_cla32_fa15_15_xor1;
  assign s_csamul_cla32_fa14_16_xor1 = s_csamul_cla32_fa14_16_xor0 ^ s_csamul_cla32_fa14_15_or0;
  assign s_csamul_cla32_fa14_16_and1 = s_csamul_cla32_fa14_16_xor0 & s_csamul_cla32_fa14_15_or0;
  assign s_csamul_cla32_fa14_16_or0 = s_csamul_cla32_fa14_16_and0 | s_csamul_cla32_fa14_16_and1;
  assign s_csamul_cla32_and15_16 = a[15] & b[16];
  assign s_csamul_cla32_fa15_16_xor0 = s_csamul_cla32_and15_16 ^ s_csamul_cla32_fa16_15_xor1;
  assign s_csamul_cla32_fa15_16_and0 = s_csamul_cla32_and15_16 & s_csamul_cla32_fa16_15_xor1;
  assign s_csamul_cla32_fa15_16_xor1 = s_csamul_cla32_fa15_16_xor0 ^ s_csamul_cla32_fa15_15_or0;
  assign s_csamul_cla32_fa15_16_and1 = s_csamul_cla32_fa15_16_xor0 & s_csamul_cla32_fa15_15_or0;
  assign s_csamul_cla32_fa15_16_or0 = s_csamul_cla32_fa15_16_and0 | s_csamul_cla32_fa15_16_and1;
  assign s_csamul_cla32_and16_16 = a[16] & b[16];
  assign s_csamul_cla32_fa16_16_xor0 = s_csamul_cla32_and16_16 ^ s_csamul_cla32_fa17_15_xor1;
  assign s_csamul_cla32_fa16_16_and0 = s_csamul_cla32_and16_16 & s_csamul_cla32_fa17_15_xor1;
  assign s_csamul_cla32_fa16_16_xor1 = s_csamul_cla32_fa16_16_xor0 ^ s_csamul_cla32_fa16_15_or0;
  assign s_csamul_cla32_fa16_16_and1 = s_csamul_cla32_fa16_16_xor0 & s_csamul_cla32_fa16_15_or0;
  assign s_csamul_cla32_fa16_16_or0 = s_csamul_cla32_fa16_16_and0 | s_csamul_cla32_fa16_16_and1;
  assign s_csamul_cla32_and17_16 = a[17] & b[16];
  assign s_csamul_cla32_fa17_16_xor0 = s_csamul_cla32_and17_16 ^ s_csamul_cla32_fa18_15_xor1;
  assign s_csamul_cla32_fa17_16_and0 = s_csamul_cla32_and17_16 & s_csamul_cla32_fa18_15_xor1;
  assign s_csamul_cla32_fa17_16_xor1 = s_csamul_cla32_fa17_16_xor0 ^ s_csamul_cla32_fa17_15_or0;
  assign s_csamul_cla32_fa17_16_and1 = s_csamul_cla32_fa17_16_xor0 & s_csamul_cla32_fa17_15_or0;
  assign s_csamul_cla32_fa17_16_or0 = s_csamul_cla32_fa17_16_and0 | s_csamul_cla32_fa17_16_and1;
  assign s_csamul_cla32_and18_16 = a[18] & b[16];
  assign s_csamul_cla32_fa18_16_xor0 = s_csamul_cla32_and18_16 ^ s_csamul_cla32_fa19_15_xor1;
  assign s_csamul_cla32_fa18_16_and0 = s_csamul_cla32_and18_16 & s_csamul_cla32_fa19_15_xor1;
  assign s_csamul_cla32_fa18_16_xor1 = s_csamul_cla32_fa18_16_xor0 ^ s_csamul_cla32_fa18_15_or0;
  assign s_csamul_cla32_fa18_16_and1 = s_csamul_cla32_fa18_16_xor0 & s_csamul_cla32_fa18_15_or0;
  assign s_csamul_cla32_fa18_16_or0 = s_csamul_cla32_fa18_16_and0 | s_csamul_cla32_fa18_16_and1;
  assign s_csamul_cla32_and19_16 = a[19] & b[16];
  assign s_csamul_cla32_fa19_16_xor0 = s_csamul_cla32_and19_16 ^ s_csamul_cla32_fa20_15_xor1;
  assign s_csamul_cla32_fa19_16_and0 = s_csamul_cla32_and19_16 & s_csamul_cla32_fa20_15_xor1;
  assign s_csamul_cla32_fa19_16_xor1 = s_csamul_cla32_fa19_16_xor0 ^ s_csamul_cla32_fa19_15_or0;
  assign s_csamul_cla32_fa19_16_and1 = s_csamul_cla32_fa19_16_xor0 & s_csamul_cla32_fa19_15_or0;
  assign s_csamul_cla32_fa19_16_or0 = s_csamul_cla32_fa19_16_and0 | s_csamul_cla32_fa19_16_and1;
  assign s_csamul_cla32_and20_16 = a[20] & b[16];
  assign s_csamul_cla32_fa20_16_xor0 = s_csamul_cla32_and20_16 ^ s_csamul_cla32_fa21_15_xor1;
  assign s_csamul_cla32_fa20_16_and0 = s_csamul_cla32_and20_16 & s_csamul_cla32_fa21_15_xor1;
  assign s_csamul_cla32_fa20_16_xor1 = s_csamul_cla32_fa20_16_xor0 ^ s_csamul_cla32_fa20_15_or0;
  assign s_csamul_cla32_fa20_16_and1 = s_csamul_cla32_fa20_16_xor0 & s_csamul_cla32_fa20_15_or0;
  assign s_csamul_cla32_fa20_16_or0 = s_csamul_cla32_fa20_16_and0 | s_csamul_cla32_fa20_16_and1;
  assign s_csamul_cla32_and21_16 = a[21] & b[16];
  assign s_csamul_cla32_fa21_16_xor0 = s_csamul_cla32_and21_16 ^ s_csamul_cla32_fa22_15_xor1;
  assign s_csamul_cla32_fa21_16_and0 = s_csamul_cla32_and21_16 & s_csamul_cla32_fa22_15_xor1;
  assign s_csamul_cla32_fa21_16_xor1 = s_csamul_cla32_fa21_16_xor0 ^ s_csamul_cla32_fa21_15_or0;
  assign s_csamul_cla32_fa21_16_and1 = s_csamul_cla32_fa21_16_xor0 & s_csamul_cla32_fa21_15_or0;
  assign s_csamul_cla32_fa21_16_or0 = s_csamul_cla32_fa21_16_and0 | s_csamul_cla32_fa21_16_and1;
  assign s_csamul_cla32_and22_16 = a[22] & b[16];
  assign s_csamul_cla32_fa22_16_xor0 = s_csamul_cla32_and22_16 ^ s_csamul_cla32_fa23_15_xor1;
  assign s_csamul_cla32_fa22_16_and0 = s_csamul_cla32_and22_16 & s_csamul_cla32_fa23_15_xor1;
  assign s_csamul_cla32_fa22_16_xor1 = s_csamul_cla32_fa22_16_xor0 ^ s_csamul_cla32_fa22_15_or0;
  assign s_csamul_cla32_fa22_16_and1 = s_csamul_cla32_fa22_16_xor0 & s_csamul_cla32_fa22_15_or0;
  assign s_csamul_cla32_fa22_16_or0 = s_csamul_cla32_fa22_16_and0 | s_csamul_cla32_fa22_16_and1;
  assign s_csamul_cla32_and23_16 = a[23] & b[16];
  assign s_csamul_cla32_fa23_16_xor0 = s_csamul_cla32_and23_16 ^ s_csamul_cla32_fa24_15_xor1;
  assign s_csamul_cla32_fa23_16_and0 = s_csamul_cla32_and23_16 & s_csamul_cla32_fa24_15_xor1;
  assign s_csamul_cla32_fa23_16_xor1 = s_csamul_cla32_fa23_16_xor0 ^ s_csamul_cla32_fa23_15_or0;
  assign s_csamul_cla32_fa23_16_and1 = s_csamul_cla32_fa23_16_xor0 & s_csamul_cla32_fa23_15_or0;
  assign s_csamul_cla32_fa23_16_or0 = s_csamul_cla32_fa23_16_and0 | s_csamul_cla32_fa23_16_and1;
  assign s_csamul_cla32_and24_16 = a[24] & b[16];
  assign s_csamul_cla32_fa24_16_xor0 = s_csamul_cla32_and24_16 ^ s_csamul_cla32_fa25_15_xor1;
  assign s_csamul_cla32_fa24_16_and0 = s_csamul_cla32_and24_16 & s_csamul_cla32_fa25_15_xor1;
  assign s_csamul_cla32_fa24_16_xor1 = s_csamul_cla32_fa24_16_xor0 ^ s_csamul_cla32_fa24_15_or0;
  assign s_csamul_cla32_fa24_16_and1 = s_csamul_cla32_fa24_16_xor0 & s_csamul_cla32_fa24_15_or0;
  assign s_csamul_cla32_fa24_16_or0 = s_csamul_cla32_fa24_16_and0 | s_csamul_cla32_fa24_16_and1;
  assign s_csamul_cla32_and25_16 = a[25] & b[16];
  assign s_csamul_cla32_fa25_16_xor0 = s_csamul_cla32_and25_16 ^ s_csamul_cla32_fa26_15_xor1;
  assign s_csamul_cla32_fa25_16_and0 = s_csamul_cla32_and25_16 & s_csamul_cla32_fa26_15_xor1;
  assign s_csamul_cla32_fa25_16_xor1 = s_csamul_cla32_fa25_16_xor0 ^ s_csamul_cla32_fa25_15_or0;
  assign s_csamul_cla32_fa25_16_and1 = s_csamul_cla32_fa25_16_xor0 & s_csamul_cla32_fa25_15_or0;
  assign s_csamul_cla32_fa25_16_or0 = s_csamul_cla32_fa25_16_and0 | s_csamul_cla32_fa25_16_and1;
  assign s_csamul_cla32_and26_16 = a[26] & b[16];
  assign s_csamul_cla32_fa26_16_xor0 = s_csamul_cla32_and26_16 ^ s_csamul_cla32_fa27_15_xor1;
  assign s_csamul_cla32_fa26_16_and0 = s_csamul_cla32_and26_16 & s_csamul_cla32_fa27_15_xor1;
  assign s_csamul_cla32_fa26_16_xor1 = s_csamul_cla32_fa26_16_xor0 ^ s_csamul_cla32_fa26_15_or0;
  assign s_csamul_cla32_fa26_16_and1 = s_csamul_cla32_fa26_16_xor0 & s_csamul_cla32_fa26_15_or0;
  assign s_csamul_cla32_fa26_16_or0 = s_csamul_cla32_fa26_16_and0 | s_csamul_cla32_fa26_16_and1;
  assign s_csamul_cla32_and27_16 = a[27] & b[16];
  assign s_csamul_cla32_fa27_16_xor0 = s_csamul_cla32_and27_16 ^ s_csamul_cla32_fa28_15_xor1;
  assign s_csamul_cla32_fa27_16_and0 = s_csamul_cla32_and27_16 & s_csamul_cla32_fa28_15_xor1;
  assign s_csamul_cla32_fa27_16_xor1 = s_csamul_cla32_fa27_16_xor0 ^ s_csamul_cla32_fa27_15_or0;
  assign s_csamul_cla32_fa27_16_and1 = s_csamul_cla32_fa27_16_xor0 & s_csamul_cla32_fa27_15_or0;
  assign s_csamul_cla32_fa27_16_or0 = s_csamul_cla32_fa27_16_and0 | s_csamul_cla32_fa27_16_and1;
  assign s_csamul_cla32_and28_16 = a[28] & b[16];
  assign s_csamul_cla32_fa28_16_xor0 = s_csamul_cla32_and28_16 ^ s_csamul_cla32_fa29_15_xor1;
  assign s_csamul_cla32_fa28_16_and0 = s_csamul_cla32_and28_16 & s_csamul_cla32_fa29_15_xor1;
  assign s_csamul_cla32_fa28_16_xor1 = s_csamul_cla32_fa28_16_xor0 ^ s_csamul_cla32_fa28_15_or0;
  assign s_csamul_cla32_fa28_16_and1 = s_csamul_cla32_fa28_16_xor0 & s_csamul_cla32_fa28_15_or0;
  assign s_csamul_cla32_fa28_16_or0 = s_csamul_cla32_fa28_16_and0 | s_csamul_cla32_fa28_16_and1;
  assign s_csamul_cla32_and29_16 = a[29] & b[16];
  assign s_csamul_cla32_fa29_16_xor0 = s_csamul_cla32_and29_16 ^ s_csamul_cla32_fa30_15_xor1;
  assign s_csamul_cla32_fa29_16_and0 = s_csamul_cla32_and29_16 & s_csamul_cla32_fa30_15_xor1;
  assign s_csamul_cla32_fa29_16_xor1 = s_csamul_cla32_fa29_16_xor0 ^ s_csamul_cla32_fa29_15_or0;
  assign s_csamul_cla32_fa29_16_and1 = s_csamul_cla32_fa29_16_xor0 & s_csamul_cla32_fa29_15_or0;
  assign s_csamul_cla32_fa29_16_or0 = s_csamul_cla32_fa29_16_and0 | s_csamul_cla32_fa29_16_and1;
  assign s_csamul_cla32_and30_16 = a[30] & b[16];
  assign s_csamul_cla32_fa30_16_xor0 = s_csamul_cla32_and30_16 ^ s_csamul_cla32_ha31_15_xor0;
  assign s_csamul_cla32_fa30_16_and0 = s_csamul_cla32_and30_16 & s_csamul_cla32_ha31_15_xor0;
  assign s_csamul_cla32_fa30_16_xor1 = s_csamul_cla32_fa30_16_xor0 ^ s_csamul_cla32_fa30_15_or0;
  assign s_csamul_cla32_fa30_16_and1 = s_csamul_cla32_fa30_16_xor0 & s_csamul_cla32_fa30_15_or0;
  assign s_csamul_cla32_fa30_16_or0 = s_csamul_cla32_fa30_16_and0 | s_csamul_cla32_fa30_16_and1;
  assign s_csamul_cla32_nand31_16 = ~(a[31] & b[16]);
  assign s_csamul_cla32_ha31_16_xor0 = s_csamul_cla32_nand31_16 ^ s_csamul_cla32_ha31_15_and0;
  assign s_csamul_cla32_ha31_16_and0 = s_csamul_cla32_nand31_16 & s_csamul_cla32_ha31_15_and0;
  assign s_csamul_cla32_and0_17 = a[0] & b[17];
  assign s_csamul_cla32_fa0_17_xor0 = s_csamul_cla32_and0_17 ^ s_csamul_cla32_fa1_16_xor1;
  assign s_csamul_cla32_fa0_17_and0 = s_csamul_cla32_and0_17 & s_csamul_cla32_fa1_16_xor1;
  assign s_csamul_cla32_fa0_17_xor1 = s_csamul_cla32_fa0_17_xor0 ^ s_csamul_cla32_fa0_16_or0;
  assign s_csamul_cla32_fa0_17_and1 = s_csamul_cla32_fa0_17_xor0 & s_csamul_cla32_fa0_16_or0;
  assign s_csamul_cla32_fa0_17_or0 = s_csamul_cla32_fa0_17_and0 | s_csamul_cla32_fa0_17_and1;
  assign s_csamul_cla32_and1_17 = a[1] & b[17];
  assign s_csamul_cla32_fa1_17_xor0 = s_csamul_cla32_and1_17 ^ s_csamul_cla32_fa2_16_xor1;
  assign s_csamul_cla32_fa1_17_and0 = s_csamul_cla32_and1_17 & s_csamul_cla32_fa2_16_xor1;
  assign s_csamul_cla32_fa1_17_xor1 = s_csamul_cla32_fa1_17_xor0 ^ s_csamul_cla32_fa1_16_or0;
  assign s_csamul_cla32_fa1_17_and1 = s_csamul_cla32_fa1_17_xor0 & s_csamul_cla32_fa1_16_or0;
  assign s_csamul_cla32_fa1_17_or0 = s_csamul_cla32_fa1_17_and0 | s_csamul_cla32_fa1_17_and1;
  assign s_csamul_cla32_and2_17 = a[2] & b[17];
  assign s_csamul_cla32_fa2_17_xor0 = s_csamul_cla32_and2_17 ^ s_csamul_cla32_fa3_16_xor1;
  assign s_csamul_cla32_fa2_17_and0 = s_csamul_cla32_and2_17 & s_csamul_cla32_fa3_16_xor1;
  assign s_csamul_cla32_fa2_17_xor1 = s_csamul_cla32_fa2_17_xor0 ^ s_csamul_cla32_fa2_16_or0;
  assign s_csamul_cla32_fa2_17_and1 = s_csamul_cla32_fa2_17_xor0 & s_csamul_cla32_fa2_16_or0;
  assign s_csamul_cla32_fa2_17_or0 = s_csamul_cla32_fa2_17_and0 | s_csamul_cla32_fa2_17_and1;
  assign s_csamul_cla32_and3_17 = a[3] & b[17];
  assign s_csamul_cla32_fa3_17_xor0 = s_csamul_cla32_and3_17 ^ s_csamul_cla32_fa4_16_xor1;
  assign s_csamul_cla32_fa3_17_and0 = s_csamul_cla32_and3_17 & s_csamul_cla32_fa4_16_xor1;
  assign s_csamul_cla32_fa3_17_xor1 = s_csamul_cla32_fa3_17_xor0 ^ s_csamul_cla32_fa3_16_or0;
  assign s_csamul_cla32_fa3_17_and1 = s_csamul_cla32_fa3_17_xor0 & s_csamul_cla32_fa3_16_or0;
  assign s_csamul_cla32_fa3_17_or0 = s_csamul_cla32_fa3_17_and0 | s_csamul_cla32_fa3_17_and1;
  assign s_csamul_cla32_and4_17 = a[4] & b[17];
  assign s_csamul_cla32_fa4_17_xor0 = s_csamul_cla32_and4_17 ^ s_csamul_cla32_fa5_16_xor1;
  assign s_csamul_cla32_fa4_17_and0 = s_csamul_cla32_and4_17 & s_csamul_cla32_fa5_16_xor1;
  assign s_csamul_cla32_fa4_17_xor1 = s_csamul_cla32_fa4_17_xor0 ^ s_csamul_cla32_fa4_16_or0;
  assign s_csamul_cla32_fa4_17_and1 = s_csamul_cla32_fa4_17_xor0 & s_csamul_cla32_fa4_16_or0;
  assign s_csamul_cla32_fa4_17_or0 = s_csamul_cla32_fa4_17_and0 | s_csamul_cla32_fa4_17_and1;
  assign s_csamul_cla32_and5_17 = a[5] & b[17];
  assign s_csamul_cla32_fa5_17_xor0 = s_csamul_cla32_and5_17 ^ s_csamul_cla32_fa6_16_xor1;
  assign s_csamul_cla32_fa5_17_and0 = s_csamul_cla32_and5_17 & s_csamul_cla32_fa6_16_xor1;
  assign s_csamul_cla32_fa5_17_xor1 = s_csamul_cla32_fa5_17_xor0 ^ s_csamul_cla32_fa5_16_or0;
  assign s_csamul_cla32_fa5_17_and1 = s_csamul_cla32_fa5_17_xor0 & s_csamul_cla32_fa5_16_or0;
  assign s_csamul_cla32_fa5_17_or0 = s_csamul_cla32_fa5_17_and0 | s_csamul_cla32_fa5_17_and1;
  assign s_csamul_cla32_and6_17 = a[6] & b[17];
  assign s_csamul_cla32_fa6_17_xor0 = s_csamul_cla32_and6_17 ^ s_csamul_cla32_fa7_16_xor1;
  assign s_csamul_cla32_fa6_17_and0 = s_csamul_cla32_and6_17 & s_csamul_cla32_fa7_16_xor1;
  assign s_csamul_cla32_fa6_17_xor1 = s_csamul_cla32_fa6_17_xor0 ^ s_csamul_cla32_fa6_16_or0;
  assign s_csamul_cla32_fa6_17_and1 = s_csamul_cla32_fa6_17_xor0 & s_csamul_cla32_fa6_16_or0;
  assign s_csamul_cla32_fa6_17_or0 = s_csamul_cla32_fa6_17_and0 | s_csamul_cla32_fa6_17_and1;
  assign s_csamul_cla32_and7_17 = a[7] & b[17];
  assign s_csamul_cla32_fa7_17_xor0 = s_csamul_cla32_and7_17 ^ s_csamul_cla32_fa8_16_xor1;
  assign s_csamul_cla32_fa7_17_and0 = s_csamul_cla32_and7_17 & s_csamul_cla32_fa8_16_xor1;
  assign s_csamul_cla32_fa7_17_xor1 = s_csamul_cla32_fa7_17_xor0 ^ s_csamul_cla32_fa7_16_or0;
  assign s_csamul_cla32_fa7_17_and1 = s_csamul_cla32_fa7_17_xor0 & s_csamul_cla32_fa7_16_or0;
  assign s_csamul_cla32_fa7_17_or0 = s_csamul_cla32_fa7_17_and0 | s_csamul_cla32_fa7_17_and1;
  assign s_csamul_cla32_and8_17 = a[8] & b[17];
  assign s_csamul_cla32_fa8_17_xor0 = s_csamul_cla32_and8_17 ^ s_csamul_cla32_fa9_16_xor1;
  assign s_csamul_cla32_fa8_17_and0 = s_csamul_cla32_and8_17 & s_csamul_cla32_fa9_16_xor1;
  assign s_csamul_cla32_fa8_17_xor1 = s_csamul_cla32_fa8_17_xor0 ^ s_csamul_cla32_fa8_16_or0;
  assign s_csamul_cla32_fa8_17_and1 = s_csamul_cla32_fa8_17_xor0 & s_csamul_cla32_fa8_16_or0;
  assign s_csamul_cla32_fa8_17_or0 = s_csamul_cla32_fa8_17_and0 | s_csamul_cla32_fa8_17_and1;
  assign s_csamul_cla32_and9_17 = a[9] & b[17];
  assign s_csamul_cla32_fa9_17_xor0 = s_csamul_cla32_and9_17 ^ s_csamul_cla32_fa10_16_xor1;
  assign s_csamul_cla32_fa9_17_and0 = s_csamul_cla32_and9_17 & s_csamul_cla32_fa10_16_xor1;
  assign s_csamul_cla32_fa9_17_xor1 = s_csamul_cla32_fa9_17_xor0 ^ s_csamul_cla32_fa9_16_or0;
  assign s_csamul_cla32_fa9_17_and1 = s_csamul_cla32_fa9_17_xor0 & s_csamul_cla32_fa9_16_or0;
  assign s_csamul_cla32_fa9_17_or0 = s_csamul_cla32_fa9_17_and0 | s_csamul_cla32_fa9_17_and1;
  assign s_csamul_cla32_and10_17 = a[10] & b[17];
  assign s_csamul_cla32_fa10_17_xor0 = s_csamul_cla32_and10_17 ^ s_csamul_cla32_fa11_16_xor1;
  assign s_csamul_cla32_fa10_17_and0 = s_csamul_cla32_and10_17 & s_csamul_cla32_fa11_16_xor1;
  assign s_csamul_cla32_fa10_17_xor1 = s_csamul_cla32_fa10_17_xor0 ^ s_csamul_cla32_fa10_16_or0;
  assign s_csamul_cla32_fa10_17_and1 = s_csamul_cla32_fa10_17_xor0 & s_csamul_cla32_fa10_16_or0;
  assign s_csamul_cla32_fa10_17_or0 = s_csamul_cla32_fa10_17_and0 | s_csamul_cla32_fa10_17_and1;
  assign s_csamul_cla32_and11_17 = a[11] & b[17];
  assign s_csamul_cla32_fa11_17_xor0 = s_csamul_cla32_and11_17 ^ s_csamul_cla32_fa12_16_xor1;
  assign s_csamul_cla32_fa11_17_and0 = s_csamul_cla32_and11_17 & s_csamul_cla32_fa12_16_xor1;
  assign s_csamul_cla32_fa11_17_xor1 = s_csamul_cla32_fa11_17_xor0 ^ s_csamul_cla32_fa11_16_or0;
  assign s_csamul_cla32_fa11_17_and1 = s_csamul_cla32_fa11_17_xor0 & s_csamul_cla32_fa11_16_or0;
  assign s_csamul_cla32_fa11_17_or0 = s_csamul_cla32_fa11_17_and0 | s_csamul_cla32_fa11_17_and1;
  assign s_csamul_cla32_and12_17 = a[12] & b[17];
  assign s_csamul_cla32_fa12_17_xor0 = s_csamul_cla32_and12_17 ^ s_csamul_cla32_fa13_16_xor1;
  assign s_csamul_cla32_fa12_17_and0 = s_csamul_cla32_and12_17 & s_csamul_cla32_fa13_16_xor1;
  assign s_csamul_cla32_fa12_17_xor1 = s_csamul_cla32_fa12_17_xor0 ^ s_csamul_cla32_fa12_16_or0;
  assign s_csamul_cla32_fa12_17_and1 = s_csamul_cla32_fa12_17_xor0 & s_csamul_cla32_fa12_16_or0;
  assign s_csamul_cla32_fa12_17_or0 = s_csamul_cla32_fa12_17_and0 | s_csamul_cla32_fa12_17_and1;
  assign s_csamul_cla32_and13_17 = a[13] & b[17];
  assign s_csamul_cla32_fa13_17_xor0 = s_csamul_cla32_and13_17 ^ s_csamul_cla32_fa14_16_xor1;
  assign s_csamul_cla32_fa13_17_and0 = s_csamul_cla32_and13_17 & s_csamul_cla32_fa14_16_xor1;
  assign s_csamul_cla32_fa13_17_xor1 = s_csamul_cla32_fa13_17_xor0 ^ s_csamul_cla32_fa13_16_or0;
  assign s_csamul_cla32_fa13_17_and1 = s_csamul_cla32_fa13_17_xor0 & s_csamul_cla32_fa13_16_or0;
  assign s_csamul_cla32_fa13_17_or0 = s_csamul_cla32_fa13_17_and0 | s_csamul_cla32_fa13_17_and1;
  assign s_csamul_cla32_and14_17 = a[14] & b[17];
  assign s_csamul_cla32_fa14_17_xor0 = s_csamul_cla32_and14_17 ^ s_csamul_cla32_fa15_16_xor1;
  assign s_csamul_cla32_fa14_17_and0 = s_csamul_cla32_and14_17 & s_csamul_cla32_fa15_16_xor1;
  assign s_csamul_cla32_fa14_17_xor1 = s_csamul_cla32_fa14_17_xor0 ^ s_csamul_cla32_fa14_16_or0;
  assign s_csamul_cla32_fa14_17_and1 = s_csamul_cla32_fa14_17_xor0 & s_csamul_cla32_fa14_16_or0;
  assign s_csamul_cla32_fa14_17_or0 = s_csamul_cla32_fa14_17_and0 | s_csamul_cla32_fa14_17_and1;
  assign s_csamul_cla32_and15_17 = a[15] & b[17];
  assign s_csamul_cla32_fa15_17_xor0 = s_csamul_cla32_and15_17 ^ s_csamul_cla32_fa16_16_xor1;
  assign s_csamul_cla32_fa15_17_and0 = s_csamul_cla32_and15_17 & s_csamul_cla32_fa16_16_xor1;
  assign s_csamul_cla32_fa15_17_xor1 = s_csamul_cla32_fa15_17_xor0 ^ s_csamul_cla32_fa15_16_or0;
  assign s_csamul_cla32_fa15_17_and1 = s_csamul_cla32_fa15_17_xor0 & s_csamul_cla32_fa15_16_or0;
  assign s_csamul_cla32_fa15_17_or0 = s_csamul_cla32_fa15_17_and0 | s_csamul_cla32_fa15_17_and1;
  assign s_csamul_cla32_and16_17 = a[16] & b[17];
  assign s_csamul_cla32_fa16_17_xor0 = s_csamul_cla32_and16_17 ^ s_csamul_cla32_fa17_16_xor1;
  assign s_csamul_cla32_fa16_17_and0 = s_csamul_cla32_and16_17 & s_csamul_cla32_fa17_16_xor1;
  assign s_csamul_cla32_fa16_17_xor1 = s_csamul_cla32_fa16_17_xor0 ^ s_csamul_cla32_fa16_16_or0;
  assign s_csamul_cla32_fa16_17_and1 = s_csamul_cla32_fa16_17_xor0 & s_csamul_cla32_fa16_16_or0;
  assign s_csamul_cla32_fa16_17_or0 = s_csamul_cla32_fa16_17_and0 | s_csamul_cla32_fa16_17_and1;
  assign s_csamul_cla32_and17_17 = a[17] & b[17];
  assign s_csamul_cla32_fa17_17_xor0 = s_csamul_cla32_and17_17 ^ s_csamul_cla32_fa18_16_xor1;
  assign s_csamul_cla32_fa17_17_and0 = s_csamul_cla32_and17_17 & s_csamul_cla32_fa18_16_xor1;
  assign s_csamul_cla32_fa17_17_xor1 = s_csamul_cla32_fa17_17_xor0 ^ s_csamul_cla32_fa17_16_or0;
  assign s_csamul_cla32_fa17_17_and1 = s_csamul_cla32_fa17_17_xor0 & s_csamul_cla32_fa17_16_or0;
  assign s_csamul_cla32_fa17_17_or0 = s_csamul_cla32_fa17_17_and0 | s_csamul_cla32_fa17_17_and1;
  assign s_csamul_cla32_and18_17 = a[18] & b[17];
  assign s_csamul_cla32_fa18_17_xor0 = s_csamul_cla32_and18_17 ^ s_csamul_cla32_fa19_16_xor1;
  assign s_csamul_cla32_fa18_17_and0 = s_csamul_cla32_and18_17 & s_csamul_cla32_fa19_16_xor1;
  assign s_csamul_cla32_fa18_17_xor1 = s_csamul_cla32_fa18_17_xor0 ^ s_csamul_cla32_fa18_16_or0;
  assign s_csamul_cla32_fa18_17_and1 = s_csamul_cla32_fa18_17_xor0 & s_csamul_cla32_fa18_16_or0;
  assign s_csamul_cla32_fa18_17_or0 = s_csamul_cla32_fa18_17_and0 | s_csamul_cla32_fa18_17_and1;
  assign s_csamul_cla32_and19_17 = a[19] & b[17];
  assign s_csamul_cla32_fa19_17_xor0 = s_csamul_cla32_and19_17 ^ s_csamul_cla32_fa20_16_xor1;
  assign s_csamul_cla32_fa19_17_and0 = s_csamul_cla32_and19_17 & s_csamul_cla32_fa20_16_xor1;
  assign s_csamul_cla32_fa19_17_xor1 = s_csamul_cla32_fa19_17_xor0 ^ s_csamul_cla32_fa19_16_or0;
  assign s_csamul_cla32_fa19_17_and1 = s_csamul_cla32_fa19_17_xor0 & s_csamul_cla32_fa19_16_or0;
  assign s_csamul_cla32_fa19_17_or0 = s_csamul_cla32_fa19_17_and0 | s_csamul_cla32_fa19_17_and1;
  assign s_csamul_cla32_and20_17 = a[20] & b[17];
  assign s_csamul_cla32_fa20_17_xor0 = s_csamul_cla32_and20_17 ^ s_csamul_cla32_fa21_16_xor1;
  assign s_csamul_cla32_fa20_17_and0 = s_csamul_cla32_and20_17 & s_csamul_cla32_fa21_16_xor1;
  assign s_csamul_cla32_fa20_17_xor1 = s_csamul_cla32_fa20_17_xor0 ^ s_csamul_cla32_fa20_16_or0;
  assign s_csamul_cla32_fa20_17_and1 = s_csamul_cla32_fa20_17_xor0 & s_csamul_cla32_fa20_16_or0;
  assign s_csamul_cla32_fa20_17_or0 = s_csamul_cla32_fa20_17_and0 | s_csamul_cla32_fa20_17_and1;
  assign s_csamul_cla32_and21_17 = a[21] & b[17];
  assign s_csamul_cla32_fa21_17_xor0 = s_csamul_cla32_and21_17 ^ s_csamul_cla32_fa22_16_xor1;
  assign s_csamul_cla32_fa21_17_and0 = s_csamul_cla32_and21_17 & s_csamul_cla32_fa22_16_xor1;
  assign s_csamul_cla32_fa21_17_xor1 = s_csamul_cla32_fa21_17_xor0 ^ s_csamul_cla32_fa21_16_or0;
  assign s_csamul_cla32_fa21_17_and1 = s_csamul_cla32_fa21_17_xor0 & s_csamul_cla32_fa21_16_or0;
  assign s_csamul_cla32_fa21_17_or0 = s_csamul_cla32_fa21_17_and0 | s_csamul_cla32_fa21_17_and1;
  assign s_csamul_cla32_and22_17 = a[22] & b[17];
  assign s_csamul_cla32_fa22_17_xor0 = s_csamul_cla32_and22_17 ^ s_csamul_cla32_fa23_16_xor1;
  assign s_csamul_cla32_fa22_17_and0 = s_csamul_cla32_and22_17 & s_csamul_cla32_fa23_16_xor1;
  assign s_csamul_cla32_fa22_17_xor1 = s_csamul_cla32_fa22_17_xor0 ^ s_csamul_cla32_fa22_16_or0;
  assign s_csamul_cla32_fa22_17_and1 = s_csamul_cla32_fa22_17_xor0 & s_csamul_cla32_fa22_16_or0;
  assign s_csamul_cla32_fa22_17_or0 = s_csamul_cla32_fa22_17_and0 | s_csamul_cla32_fa22_17_and1;
  assign s_csamul_cla32_and23_17 = a[23] & b[17];
  assign s_csamul_cla32_fa23_17_xor0 = s_csamul_cla32_and23_17 ^ s_csamul_cla32_fa24_16_xor1;
  assign s_csamul_cla32_fa23_17_and0 = s_csamul_cla32_and23_17 & s_csamul_cla32_fa24_16_xor1;
  assign s_csamul_cla32_fa23_17_xor1 = s_csamul_cla32_fa23_17_xor0 ^ s_csamul_cla32_fa23_16_or0;
  assign s_csamul_cla32_fa23_17_and1 = s_csamul_cla32_fa23_17_xor0 & s_csamul_cla32_fa23_16_or0;
  assign s_csamul_cla32_fa23_17_or0 = s_csamul_cla32_fa23_17_and0 | s_csamul_cla32_fa23_17_and1;
  assign s_csamul_cla32_and24_17 = a[24] & b[17];
  assign s_csamul_cla32_fa24_17_xor0 = s_csamul_cla32_and24_17 ^ s_csamul_cla32_fa25_16_xor1;
  assign s_csamul_cla32_fa24_17_and0 = s_csamul_cla32_and24_17 & s_csamul_cla32_fa25_16_xor1;
  assign s_csamul_cla32_fa24_17_xor1 = s_csamul_cla32_fa24_17_xor0 ^ s_csamul_cla32_fa24_16_or0;
  assign s_csamul_cla32_fa24_17_and1 = s_csamul_cla32_fa24_17_xor0 & s_csamul_cla32_fa24_16_or0;
  assign s_csamul_cla32_fa24_17_or0 = s_csamul_cla32_fa24_17_and0 | s_csamul_cla32_fa24_17_and1;
  assign s_csamul_cla32_and25_17 = a[25] & b[17];
  assign s_csamul_cla32_fa25_17_xor0 = s_csamul_cla32_and25_17 ^ s_csamul_cla32_fa26_16_xor1;
  assign s_csamul_cla32_fa25_17_and0 = s_csamul_cla32_and25_17 & s_csamul_cla32_fa26_16_xor1;
  assign s_csamul_cla32_fa25_17_xor1 = s_csamul_cla32_fa25_17_xor0 ^ s_csamul_cla32_fa25_16_or0;
  assign s_csamul_cla32_fa25_17_and1 = s_csamul_cla32_fa25_17_xor0 & s_csamul_cla32_fa25_16_or0;
  assign s_csamul_cla32_fa25_17_or0 = s_csamul_cla32_fa25_17_and0 | s_csamul_cla32_fa25_17_and1;
  assign s_csamul_cla32_and26_17 = a[26] & b[17];
  assign s_csamul_cla32_fa26_17_xor0 = s_csamul_cla32_and26_17 ^ s_csamul_cla32_fa27_16_xor1;
  assign s_csamul_cla32_fa26_17_and0 = s_csamul_cla32_and26_17 & s_csamul_cla32_fa27_16_xor1;
  assign s_csamul_cla32_fa26_17_xor1 = s_csamul_cla32_fa26_17_xor0 ^ s_csamul_cla32_fa26_16_or0;
  assign s_csamul_cla32_fa26_17_and1 = s_csamul_cla32_fa26_17_xor0 & s_csamul_cla32_fa26_16_or0;
  assign s_csamul_cla32_fa26_17_or0 = s_csamul_cla32_fa26_17_and0 | s_csamul_cla32_fa26_17_and1;
  assign s_csamul_cla32_and27_17 = a[27] & b[17];
  assign s_csamul_cla32_fa27_17_xor0 = s_csamul_cla32_and27_17 ^ s_csamul_cla32_fa28_16_xor1;
  assign s_csamul_cla32_fa27_17_and0 = s_csamul_cla32_and27_17 & s_csamul_cla32_fa28_16_xor1;
  assign s_csamul_cla32_fa27_17_xor1 = s_csamul_cla32_fa27_17_xor0 ^ s_csamul_cla32_fa27_16_or0;
  assign s_csamul_cla32_fa27_17_and1 = s_csamul_cla32_fa27_17_xor0 & s_csamul_cla32_fa27_16_or0;
  assign s_csamul_cla32_fa27_17_or0 = s_csamul_cla32_fa27_17_and0 | s_csamul_cla32_fa27_17_and1;
  assign s_csamul_cla32_and28_17 = a[28] & b[17];
  assign s_csamul_cla32_fa28_17_xor0 = s_csamul_cla32_and28_17 ^ s_csamul_cla32_fa29_16_xor1;
  assign s_csamul_cla32_fa28_17_and0 = s_csamul_cla32_and28_17 & s_csamul_cla32_fa29_16_xor1;
  assign s_csamul_cla32_fa28_17_xor1 = s_csamul_cla32_fa28_17_xor0 ^ s_csamul_cla32_fa28_16_or0;
  assign s_csamul_cla32_fa28_17_and1 = s_csamul_cla32_fa28_17_xor0 & s_csamul_cla32_fa28_16_or0;
  assign s_csamul_cla32_fa28_17_or0 = s_csamul_cla32_fa28_17_and0 | s_csamul_cla32_fa28_17_and1;
  assign s_csamul_cla32_and29_17 = a[29] & b[17];
  assign s_csamul_cla32_fa29_17_xor0 = s_csamul_cla32_and29_17 ^ s_csamul_cla32_fa30_16_xor1;
  assign s_csamul_cla32_fa29_17_and0 = s_csamul_cla32_and29_17 & s_csamul_cla32_fa30_16_xor1;
  assign s_csamul_cla32_fa29_17_xor1 = s_csamul_cla32_fa29_17_xor0 ^ s_csamul_cla32_fa29_16_or0;
  assign s_csamul_cla32_fa29_17_and1 = s_csamul_cla32_fa29_17_xor0 & s_csamul_cla32_fa29_16_or0;
  assign s_csamul_cla32_fa29_17_or0 = s_csamul_cla32_fa29_17_and0 | s_csamul_cla32_fa29_17_and1;
  assign s_csamul_cla32_and30_17 = a[30] & b[17];
  assign s_csamul_cla32_fa30_17_xor0 = s_csamul_cla32_and30_17 ^ s_csamul_cla32_ha31_16_xor0;
  assign s_csamul_cla32_fa30_17_and0 = s_csamul_cla32_and30_17 & s_csamul_cla32_ha31_16_xor0;
  assign s_csamul_cla32_fa30_17_xor1 = s_csamul_cla32_fa30_17_xor0 ^ s_csamul_cla32_fa30_16_or0;
  assign s_csamul_cla32_fa30_17_and1 = s_csamul_cla32_fa30_17_xor0 & s_csamul_cla32_fa30_16_or0;
  assign s_csamul_cla32_fa30_17_or0 = s_csamul_cla32_fa30_17_and0 | s_csamul_cla32_fa30_17_and1;
  assign s_csamul_cla32_nand31_17 = ~(a[31] & b[17]);
  assign s_csamul_cla32_ha31_17_xor0 = s_csamul_cla32_nand31_17 ^ s_csamul_cla32_ha31_16_and0;
  assign s_csamul_cla32_ha31_17_and0 = s_csamul_cla32_nand31_17 & s_csamul_cla32_ha31_16_and0;
  assign s_csamul_cla32_and0_18 = a[0] & b[18];
  assign s_csamul_cla32_fa0_18_xor0 = s_csamul_cla32_and0_18 ^ s_csamul_cla32_fa1_17_xor1;
  assign s_csamul_cla32_fa0_18_and0 = s_csamul_cla32_and0_18 & s_csamul_cla32_fa1_17_xor1;
  assign s_csamul_cla32_fa0_18_xor1 = s_csamul_cla32_fa0_18_xor0 ^ s_csamul_cla32_fa0_17_or0;
  assign s_csamul_cla32_fa0_18_and1 = s_csamul_cla32_fa0_18_xor0 & s_csamul_cla32_fa0_17_or0;
  assign s_csamul_cla32_fa0_18_or0 = s_csamul_cla32_fa0_18_and0 | s_csamul_cla32_fa0_18_and1;
  assign s_csamul_cla32_and1_18 = a[1] & b[18];
  assign s_csamul_cla32_fa1_18_xor0 = s_csamul_cla32_and1_18 ^ s_csamul_cla32_fa2_17_xor1;
  assign s_csamul_cla32_fa1_18_and0 = s_csamul_cla32_and1_18 & s_csamul_cla32_fa2_17_xor1;
  assign s_csamul_cla32_fa1_18_xor1 = s_csamul_cla32_fa1_18_xor0 ^ s_csamul_cla32_fa1_17_or0;
  assign s_csamul_cla32_fa1_18_and1 = s_csamul_cla32_fa1_18_xor0 & s_csamul_cla32_fa1_17_or0;
  assign s_csamul_cla32_fa1_18_or0 = s_csamul_cla32_fa1_18_and0 | s_csamul_cla32_fa1_18_and1;
  assign s_csamul_cla32_and2_18 = a[2] & b[18];
  assign s_csamul_cla32_fa2_18_xor0 = s_csamul_cla32_and2_18 ^ s_csamul_cla32_fa3_17_xor1;
  assign s_csamul_cla32_fa2_18_and0 = s_csamul_cla32_and2_18 & s_csamul_cla32_fa3_17_xor1;
  assign s_csamul_cla32_fa2_18_xor1 = s_csamul_cla32_fa2_18_xor0 ^ s_csamul_cla32_fa2_17_or0;
  assign s_csamul_cla32_fa2_18_and1 = s_csamul_cla32_fa2_18_xor0 & s_csamul_cla32_fa2_17_or0;
  assign s_csamul_cla32_fa2_18_or0 = s_csamul_cla32_fa2_18_and0 | s_csamul_cla32_fa2_18_and1;
  assign s_csamul_cla32_and3_18 = a[3] & b[18];
  assign s_csamul_cla32_fa3_18_xor0 = s_csamul_cla32_and3_18 ^ s_csamul_cla32_fa4_17_xor1;
  assign s_csamul_cla32_fa3_18_and0 = s_csamul_cla32_and3_18 & s_csamul_cla32_fa4_17_xor1;
  assign s_csamul_cla32_fa3_18_xor1 = s_csamul_cla32_fa3_18_xor0 ^ s_csamul_cla32_fa3_17_or0;
  assign s_csamul_cla32_fa3_18_and1 = s_csamul_cla32_fa3_18_xor0 & s_csamul_cla32_fa3_17_or0;
  assign s_csamul_cla32_fa3_18_or0 = s_csamul_cla32_fa3_18_and0 | s_csamul_cla32_fa3_18_and1;
  assign s_csamul_cla32_and4_18 = a[4] & b[18];
  assign s_csamul_cla32_fa4_18_xor0 = s_csamul_cla32_and4_18 ^ s_csamul_cla32_fa5_17_xor1;
  assign s_csamul_cla32_fa4_18_and0 = s_csamul_cla32_and4_18 & s_csamul_cla32_fa5_17_xor1;
  assign s_csamul_cla32_fa4_18_xor1 = s_csamul_cla32_fa4_18_xor0 ^ s_csamul_cla32_fa4_17_or0;
  assign s_csamul_cla32_fa4_18_and1 = s_csamul_cla32_fa4_18_xor0 & s_csamul_cla32_fa4_17_or0;
  assign s_csamul_cla32_fa4_18_or0 = s_csamul_cla32_fa4_18_and0 | s_csamul_cla32_fa4_18_and1;
  assign s_csamul_cla32_and5_18 = a[5] & b[18];
  assign s_csamul_cla32_fa5_18_xor0 = s_csamul_cla32_and5_18 ^ s_csamul_cla32_fa6_17_xor1;
  assign s_csamul_cla32_fa5_18_and0 = s_csamul_cla32_and5_18 & s_csamul_cla32_fa6_17_xor1;
  assign s_csamul_cla32_fa5_18_xor1 = s_csamul_cla32_fa5_18_xor0 ^ s_csamul_cla32_fa5_17_or0;
  assign s_csamul_cla32_fa5_18_and1 = s_csamul_cla32_fa5_18_xor0 & s_csamul_cla32_fa5_17_or0;
  assign s_csamul_cla32_fa5_18_or0 = s_csamul_cla32_fa5_18_and0 | s_csamul_cla32_fa5_18_and1;
  assign s_csamul_cla32_and6_18 = a[6] & b[18];
  assign s_csamul_cla32_fa6_18_xor0 = s_csamul_cla32_and6_18 ^ s_csamul_cla32_fa7_17_xor1;
  assign s_csamul_cla32_fa6_18_and0 = s_csamul_cla32_and6_18 & s_csamul_cla32_fa7_17_xor1;
  assign s_csamul_cla32_fa6_18_xor1 = s_csamul_cla32_fa6_18_xor0 ^ s_csamul_cla32_fa6_17_or0;
  assign s_csamul_cla32_fa6_18_and1 = s_csamul_cla32_fa6_18_xor0 & s_csamul_cla32_fa6_17_or0;
  assign s_csamul_cla32_fa6_18_or0 = s_csamul_cla32_fa6_18_and0 | s_csamul_cla32_fa6_18_and1;
  assign s_csamul_cla32_and7_18 = a[7] & b[18];
  assign s_csamul_cla32_fa7_18_xor0 = s_csamul_cla32_and7_18 ^ s_csamul_cla32_fa8_17_xor1;
  assign s_csamul_cla32_fa7_18_and0 = s_csamul_cla32_and7_18 & s_csamul_cla32_fa8_17_xor1;
  assign s_csamul_cla32_fa7_18_xor1 = s_csamul_cla32_fa7_18_xor0 ^ s_csamul_cla32_fa7_17_or0;
  assign s_csamul_cla32_fa7_18_and1 = s_csamul_cla32_fa7_18_xor0 & s_csamul_cla32_fa7_17_or0;
  assign s_csamul_cla32_fa7_18_or0 = s_csamul_cla32_fa7_18_and0 | s_csamul_cla32_fa7_18_and1;
  assign s_csamul_cla32_and8_18 = a[8] & b[18];
  assign s_csamul_cla32_fa8_18_xor0 = s_csamul_cla32_and8_18 ^ s_csamul_cla32_fa9_17_xor1;
  assign s_csamul_cla32_fa8_18_and0 = s_csamul_cla32_and8_18 & s_csamul_cla32_fa9_17_xor1;
  assign s_csamul_cla32_fa8_18_xor1 = s_csamul_cla32_fa8_18_xor0 ^ s_csamul_cla32_fa8_17_or0;
  assign s_csamul_cla32_fa8_18_and1 = s_csamul_cla32_fa8_18_xor0 & s_csamul_cla32_fa8_17_or0;
  assign s_csamul_cla32_fa8_18_or0 = s_csamul_cla32_fa8_18_and0 | s_csamul_cla32_fa8_18_and1;
  assign s_csamul_cla32_and9_18 = a[9] & b[18];
  assign s_csamul_cla32_fa9_18_xor0 = s_csamul_cla32_and9_18 ^ s_csamul_cla32_fa10_17_xor1;
  assign s_csamul_cla32_fa9_18_and0 = s_csamul_cla32_and9_18 & s_csamul_cla32_fa10_17_xor1;
  assign s_csamul_cla32_fa9_18_xor1 = s_csamul_cla32_fa9_18_xor0 ^ s_csamul_cla32_fa9_17_or0;
  assign s_csamul_cla32_fa9_18_and1 = s_csamul_cla32_fa9_18_xor0 & s_csamul_cla32_fa9_17_or0;
  assign s_csamul_cla32_fa9_18_or0 = s_csamul_cla32_fa9_18_and0 | s_csamul_cla32_fa9_18_and1;
  assign s_csamul_cla32_and10_18 = a[10] & b[18];
  assign s_csamul_cla32_fa10_18_xor0 = s_csamul_cla32_and10_18 ^ s_csamul_cla32_fa11_17_xor1;
  assign s_csamul_cla32_fa10_18_and0 = s_csamul_cla32_and10_18 & s_csamul_cla32_fa11_17_xor1;
  assign s_csamul_cla32_fa10_18_xor1 = s_csamul_cla32_fa10_18_xor0 ^ s_csamul_cla32_fa10_17_or0;
  assign s_csamul_cla32_fa10_18_and1 = s_csamul_cla32_fa10_18_xor0 & s_csamul_cla32_fa10_17_or0;
  assign s_csamul_cla32_fa10_18_or0 = s_csamul_cla32_fa10_18_and0 | s_csamul_cla32_fa10_18_and1;
  assign s_csamul_cla32_and11_18 = a[11] & b[18];
  assign s_csamul_cla32_fa11_18_xor0 = s_csamul_cla32_and11_18 ^ s_csamul_cla32_fa12_17_xor1;
  assign s_csamul_cla32_fa11_18_and0 = s_csamul_cla32_and11_18 & s_csamul_cla32_fa12_17_xor1;
  assign s_csamul_cla32_fa11_18_xor1 = s_csamul_cla32_fa11_18_xor0 ^ s_csamul_cla32_fa11_17_or0;
  assign s_csamul_cla32_fa11_18_and1 = s_csamul_cla32_fa11_18_xor0 & s_csamul_cla32_fa11_17_or0;
  assign s_csamul_cla32_fa11_18_or0 = s_csamul_cla32_fa11_18_and0 | s_csamul_cla32_fa11_18_and1;
  assign s_csamul_cla32_and12_18 = a[12] & b[18];
  assign s_csamul_cla32_fa12_18_xor0 = s_csamul_cla32_and12_18 ^ s_csamul_cla32_fa13_17_xor1;
  assign s_csamul_cla32_fa12_18_and0 = s_csamul_cla32_and12_18 & s_csamul_cla32_fa13_17_xor1;
  assign s_csamul_cla32_fa12_18_xor1 = s_csamul_cla32_fa12_18_xor0 ^ s_csamul_cla32_fa12_17_or0;
  assign s_csamul_cla32_fa12_18_and1 = s_csamul_cla32_fa12_18_xor0 & s_csamul_cla32_fa12_17_or0;
  assign s_csamul_cla32_fa12_18_or0 = s_csamul_cla32_fa12_18_and0 | s_csamul_cla32_fa12_18_and1;
  assign s_csamul_cla32_and13_18 = a[13] & b[18];
  assign s_csamul_cla32_fa13_18_xor0 = s_csamul_cla32_and13_18 ^ s_csamul_cla32_fa14_17_xor1;
  assign s_csamul_cla32_fa13_18_and0 = s_csamul_cla32_and13_18 & s_csamul_cla32_fa14_17_xor1;
  assign s_csamul_cla32_fa13_18_xor1 = s_csamul_cla32_fa13_18_xor0 ^ s_csamul_cla32_fa13_17_or0;
  assign s_csamul_cla32_fa13_18_and1 = s_csamul_cla32_fa13_18_xor0 & s_csamul_cla32_fa13_17_or0;
  assign s_csamul_cla32_fa13_18_or0 = s_csamul_cla32_fa13_18_and0 | s_csamul_cla32_fa13_18_and1;
  assign s_csamul_cla32_and14_18 = a[14] & b[18];
  assign s_csamul_cla32_fa14_18_xor0 = s_csamul_cla32_and14_18 ^ s_csamul_cla32_fa15_17_xor1;
  assign s_csamul_cla32_fa14_18_and0 = s_csamul_cla32_and14_18 & s_csamul_cla32_fa15_17_xor1;
  assign s_csamul_cla32_fa14_18_xor1 = s_csamul_cla32_fa14_18_xor0 ^ s_csamul_cla32_fa14_17_or0;
  assign s_csamul_cla32_fa14_18_and1 = s_csamul_cla32_fa14_18_xor0 & s_csamul_cla32_fa14_17_or0;
  assign s_csamul_cla32_fa14_18_or0 = s_csamul_cla32_fa14_18_and0 | s_csamul_cla32_fa14_18_and1;
  assign s_csamul_cla32_and15_18 = a[15] & b[18];
  assign s_csamul_cla32_fa15_18_xor0 = s_csamul_cla32_and15_18 ^ s_csamul_cla32_fa16_17_xor1;
  assign s_csamul_cla32_fa15_18_and0 = s_csamul_cla32_and15_18 & s_csamul_cla32_fa16_17_xor1;
  assign s_csamul_cla32_fa15_18_xor1 = s_csamul_cla32_fa15_18_xor0 ^ s_csamul_cla32_fa15_17_or0;
  assign s_csamul_cla32_fa15_18_and1 = s_csamul_cla32_fa15_18_xor0 & s_csamul_cla32_fa15_17_or0;
  assign s_csamul_cla32_fa15_18_or0 = s_csamul_cla32_fa15_18_and0 | s_csamul_cla32_fa15_18_and1;
  assign s_csamul_cla32_and16_18 = a[16] & b[18];
  assign s_csamul_cla32_fa16_18_xor0 = s_csamul_cla32_and16_18 ^ s_csamul_cla32_fa17_17_xor1;
  assign s_csamul_cla32_fa16_18_and0 = s_csamul_cla32_and16_18 & s_csamul_cla32_fa17_17_xor1;
  assign s_csamul_cla32_fa16_18_xor1 = s_csamul_cla32_fa16_18_xor0 ^ s_csamul_cla32_fa16_17_or0;
  assign s_csamul_cla32_fa16_18_and1 = s_csamul_cla32_fa16_18_xor0 & s_csamul_cla32_fa16_17_or0;
  assign s_csamul_cla32_fa16_18_or0 = s_csamul_cla32_fa16_18_and0 | s_csamul_cla32_fa16_18_and1;
  assign s_csamul_cla32_and17_18 = a[17] & b[18];
  assign s_csamul_cla32_fa17_18_xor0 = s_csamul_cla32_and17_18 ^ s_csamul_cla32_fa18_17_xor1;
  assign s_csamul_cla32_fa17_18_and0 = s_csamul_cla32_and17_18 & s_csamul_cla32_fa18_17_xor1;
  assign s_csamul_cla32_fa17_18_xor1 = s_csamul_cla32_fa17_18_xor0 ^ s_csamul_cla32_fa17_17_or0;
  assign s_csamul_cla32_fa17_18_and1 = s_csamul_cla32_fa17_18_xor0 & s_csamul_cla32_fa17_17_or0;
  assign s_csamul_cla32_fa17_18_or0 = s_csamul_cla32_fa17_18_and0 | s_csamul_cla32_fa17_18_and1;
  assign s_csamul_cla32_and18_18 = a[18] & b[18];
  assign s_csamul_cla32_fa18_18_xor0 = s_csamul_cla32_and18_18 ^ s_csamul_cla32_fa19_17_xor1;
  assign s_csamul_cla32_fa18_18_and0 = s_csamul_cla32_and18_18 & s_csamul_cla32_fa19_17_xor1;
  assign s_csamul_cla32_fa18_18_xor1 = s_csamul_cla32_fa18_18_xor0 ^ s_csamul_cla32_fa18_17_or0;
  assign s_csamul_cla32_fa18_18_and1 = s_csamul_cla32_fa18_18_xor0 & s_csamul_cla32_fa18_17_or0;
  assign s_csamul_cla32_fa18_18_or0 = s_csamul_cla32_fa18_18_and0 | s_csamul_cla32_fa18_18_and1;
  assign s_csamul_cla32_and19_18 = a[19] & b[18];
  assign s_csamul_cla32_fa19_18_xor0 = s_csamul_cla32_and19_18 ^ s_csamul_cla32_fa20_17_xor1;
  assign s_csamul_cla32_fa19_18_and0 = s_csamul_cla32_and19_18 & s_csamul_cla32_fa20_17_xor1;
  assign s_csamul_cla32_fa19_18_xor1 = s_csamul_cla32_fa19_18_xor0 ^ s_csamul_cla32_fa19_17_or0;
  assign s_csamul_cla32_fa19_18_and1 = s_csamul_cla32_fa19_18_xor0 & s_csamul_cla32_fa19_17_or0;
  assign s_csamul_cla32_fa19_18_or0 = s_csamul_cla32_fa19_18_and0 | s_csamul_cla32_fa19_18_and1;
  assign s_csamul_cla32_and20_18 = a[20] & b[18];
  assign s_csamul_cla32_fa20_18_xor0 = s_csamul_cla32_and20_18 ^ s_csamul_cla32_fa21_17_xor1;
  assign s_csamul_cla32_fa20_18_and0 = s_csamul_cla32_and20_18 & s_csamul_cla32_fa21_17_xor1;
  assign s_csamul_cla32_fa20_18_xor1 = s_csamul_cla32_fa20_18_xor0 ^ s_csamul_cla32_fa20_17_or0;
  assign s_csamul_cla32_fa20_18_and1 = s_csamul_cla32_fa20_18_xor0 & s_csamul_cla32_fa20_17_or0;
  assign s_csamul_cla32_fa20_18_or0 = s_csamul_cla32_fa20_18_and0 | s_csamul_cla32_fa20_18_and1;
  assign s_csamul_cla32_and21_18 = a[21] & b[18];
  assign s_csamul_cla32_fa21_18_xor0 = s_csamul_cla32_and21_18 ^ s_csamul_cla32_fa22_17_xor1;
  assign s_csamul_cla32_fa21_18_and0 = s_csamul_cla32_and21_18 & s_csamul_cla32_fa22_17_xor1;
  assign s_csamul_cla32_fa21_18_xor1 = s_csamul_cla32_fa21_18_xor0 ^ s_csamul_cla32_fa21_17_or0;
  assign s_csamul_cla32_fa21_18_and1 = s_csamul_cla32_fa21_18_xor0 & s_csamul_cla32_fa21_17_or0;
  assign s_csamul_cla32_fa21_18_or0 = s_csamul_cla32_fa21_18_and0 | s_csamul_cla32_fa21_18_and1;
  assign s_csamul_cla32_and22_18 = a[22] & b[18];
  assign s_csamul_cla32_fa22_18_xor0 = s_csamul_cla32_and22_18 ^ s_csamul_cla32_fa23_17_xor1;
  assign s_csamul_cla32_fa22_18_and0 = s_csamul_cla32_and22_18 & s_csamul_cla32_fa23_17_xor1;
  assign s_csamul_cla32_fa22_18_xor1 = s_csamul_cla32_fa22_18_xor0 ^ s_csamul_cla32_fa22_17_or0;
  assign s_csamul_cla32_fa22_18_and1 = s_csamul_cla32_fa22_18_xor0 & s_csamul_cla32_fa22_17_or0;
  assign s_csamul_cla32_fa22_18_or0 = s_csamul_cla32_fa22_18_and0 | s_csamul_cla32_fa22_18_and1;
  assign s_csamul_cla32_and23_18 = a[23] & b[18];
  assign s_csamul_cla32_fa23_18_xor0 = s_csamul_cla32_and23_18 ^ s_csamul_cla32_fa24_17_xor1;
  assign s_csamul_cla32_fa23_18_and0 = s_csamul_cla32_and23_18 & s_csamul_cla32_fa24_17_xor1;
  assign s_csamul_cla32_fa23_18_xor1 = s_csamul_cla32_fa23_18_xor0 ^ s_csamul_cla32_fa23_17_or0;
  assign s_csamul_cla32_fa23_18_and1 = s_csamul_cla32_fa23_18_xor0 & s_csamul_cla32_fa23_17_or0;
  assign s_csamul_cla32_fa23_18_or0 = s_csamul_cla32_fa23_18_and0 | s_csamul_cla32_fa23_18_and1;
  assign s_csamul_cla32_and24_18 = a[24] & b[18];
  assign s_csamul_cla32_fa24_18_xor0 = s_csamul_cla32_and24_18 ^ s_csamul_cla32_fa25_17_xor1;
  assign s_csamul_cla32_fa24_18_and0 = s_csamul_cla32_and24_18 & s_csamul_cla32_fa25_17_xor1;
  assign s_csamul_cla32_fa24_18_xor1 = s_csamul_cla32_fa24_18_xor0 ^ s_csamul_cla32_fa24_17_or0;
  assign s_csamul_cla32_fa24_18_and1 = s_csamul_cla32_fa24_18_xor0 & s_csamul_cla32_fa24_17_or0;
  assign s_csamul_cla32_fa24_18_or0 = s_csamul_cla32_fa24_18_and0 | s_csamul_cla32_fa24_18_and1;
  assign s_csamul_cla32_and25_18 = a[25] & b[18];
  assign s_csamul_cla32_fa25_18_xor0 = s_csamul_cla32_and25_18 ^ s_csamul_cla32_fa26_17_xor1;
  assign s_csamul_cla32_fa25_18_and0 = s_csamul_cla32_and25_18 & s_csamul_cla32_fa26_17_xor1;
  assign s_csamul_cla32_fa25_18_xor1 = s_csamul_cla32_fa25_18_xor0 ^ s_csamul_cla32_fa25_17_or0;
  assign s_csamul_cla32_fa25_18_and1 = s_csamul_cla32_fa25_18_xor0 & s_csamul_cla32_fa25_17_or0;
  assign s_csamul_cla32_fa25_18_or0 = s_csamul_cla32_fa25_18_and0 | s_csamul_cla32_fa25_18_and1;
  assign s_csamul_cla32_and26_18 = a[26] & b[18];
  assign s_csamul_cla32_fa26_18_xor0 = s_csamul_cla32_and26_18 ^ s_csamul_cla32_fa27_17_xor1;
  assign s_csamul_cla32_fa26_18_and0 = s_csamul_cla32_and26_18 & s_csamul_cla32_fa27_17_xor1;
  assign s_csamul_cla32_fa26_18_xor1 = s_csamul_cla32_fa26_18_xor0 ^ s_csamul_cla32_fa26_17_or0;
  assign s_csamul_cla32_fa26_18_and1 = s_csamul_cla32_fa26_18_xor0 & s_csamul_cla32_fa26_17_or0;
  assign s_csamul_cla32_fa26_18_or0 = s_csamul_cla32_fa26_18_and0 | s_csamul_cla32_fa26_18_and1;
  assign s_csamul_cla32_and27_18 = a[27] & b[18];
  assign s_csamul_cla32_fa27_18_xor0 = s_csamul_cla32_and27_18 ^ s_csamul_cla32_fa28_17_xor1;
  assign s_csamul_cla32_fa27_18_and0 = s_csamul_cla32_and27_18 & s_csamul_cla32_fa28_17_xor1;
  assign s_csamul_cla32_fa27_18_xor1 = s_csamul_cla32_fa27_18_xor0 ^ s_csamul_cla32_fa27_17_or0;
  assign s_csamul_cla32_fa27_18_and1 = s_csamul_cla32_fa27_18_xor0 & s_csamul_cla32_fa27_17_or0;
  assign s_csamul_cla32_fa27_18_or0 = s_csamul_cla32_fa27_18_and0 | s_csamul_cla32_fa27_18_and1;
  assign s_csamul_cla32_and28_18 = a[28] & b[18];
  assign s_csamul_cla32_fa28_18_xor0 = s_csamul_cla32_and28_18 ^ s_csamul_cla32_fa29_17_xor1;
  assign s_csamul_cla32_fa28_18_and0 = s_csamul_cla32_and28_18 & s_csamul_cla32_fa29_17_xor1;
  assign s_csamul_cla32_fa28_18_xor1 = s_csamul_cla32_fa28_18_xor0 ^ s_csamul_cla32_fa28_17_or0;
  assign s_csamul_cla32_fa28_18_and1 = s_csamul_cla32_fa28_18_xor0 & s_csamul_cla32_fa28_17_or0;
  assign s_csamul_cla32_fa28_18_or0 = s_csamul_cla32_fa28_18_and0 | s_csamul_cla32_fa28_18_and1;
  assign s_csamul_cla32_and29_18 = a[29] & b[18];
  assign s_csamul_cla32_fa29_18_xor0 = s_csamul_cla32_and29_18 ^ s_csamul_cla32_fa30_17_xor1;
  assign s_csamul_cla32_fa29_18_and0 = s_csamul_cla32_and29_18 & s_csamul_cla32_fa30_17_xor1;
  assign s_csamul_cla32_fa29_18_xor1 = s_csamul_cla32_fa29_18_xor0 ^ s_csamul_cla32_fa29_17_or0;
  assign s_csamul_cla32_fa29_18_and1 = s_csamul_cla32_fa29_18_xor0 & s_csamul_cla32_fa29_17_or0;
  assign s_csamul_cla32_fa29_18_or0 = s_csamul_cla32_fa29_18_and0 | s_csamul_cla32_fa29_18_and1;
  assign s_csamul_cla32_and30_18 = a[30] & b[18];
  assign s_csamul_cla32_fa30_18_xor0 = s_csamul_cla32_and30_18 ^ s_csamul_cla32_ha31_17_xor0;
  assign s_csamul_cla32_fa30_18_and0 = s_csamul_cla32_and30_18 & s_csamul_cla32_ha31_17_xor0;
  assign s_csamul_cla32_fa30_18_xor1 = s_csamul_cla32_fa30_18_xor0 ^ s_csamul_cla32_fa30_17_or0;
  assign s_csamul_cla32_fa30_18_and1 = s_csamul_cla32_fa30_18_xor0 & s_csamul_cla32_fa30_17_or0;
  assign s_csamul_cla32_fa30_18_or0 = s_csamul_cla32_fa30_18_and0 | s_csamul_cla32_fa30_18_and1;
  assign s_csamul_cla32_nand31_18 = ~(a[31] & b[18]);
  assign s_csamul_cla32_ha31_18_xor0 = s_csamul_cla32_nand31_18 ^ s_csamul_cla32_ha31_17_and0;
  assign s_csamul_cla32_ha31_18_and0 = s_csamul_cla32_nand31_18 & s_csamul_cla32_ha31_17_and0;
  assign s_csamul_cla32_and0_19 = a[0] & b[19];
  assign s_csamul_cla32_fa0_19_xor0 = s_csamul_cla32_and0_19 ^ s_csamul_cla32_fa1_18_xor1;
  assign s_csamul_cla32_fa0_19_and0 = s_csamul_cla32_and0_19 & s_csamul_cla32_fa1_18_xor1;
  assign s_csamul_cla32_fa0_19_xor1 = s_csamul_cla32_fa0_19_xor0 ^ s_csamul_cla32_fa0_18_or0;
  assign s_csamul_cla32_fa0_19_and1 = s_csamul_cla32_fa0_19_xor0 & s_csamul_cla32_fa0_18_or0;
  assign s_csamul_cla32_fa0_19_or0 = s_csamul_cla32_fa0_19_and0 | s_csamul_cla32_fa0_19_and1;
  assign s_csamul_cla32_and1_19 = a[1] & b[19];
  assign s_csamul_cla32_fa1_19_xor0 = s_csamul_cla32_and1_19 ^ s_csamul_cla32_fa2_18_xor1;
  assign s_csamul_cla32_fa1_19_and0 = s_csamul_cla32_and1_19 & s_csamul_cla32_fa2_18_xor1;
  assign s_csamul_cla32_fa1_19_xor1 = s_csamul_cla32_fa1_19_xor0 ^ s_csamul_cla32_fa1_18_or0;
  assign s_csamul_cla32_fa1_19_and1 = s_csamul_cla32_fa1_19_xor0 & s_csamul_cla32_fa1_18_or0;
  assign s_csamul_cla32_fa1_19_or0 = s_csamul_cla32_fa1_19_and0 | s_csamul_cla32_fa1_19_and1;
  assign s_csamul_cla32_and2_19 = a[2] & b[19];
  assign s_csamul_cla32_fa2_19_xor0 = s_csamul_cla32_and2_19 ^ s_csamul_cla32_fa3_18_xor1;
  assign s_csamul_cla32_fa2_19_and0 = s_csamul_cla32_and2_19 & s_csamul_cla32_fa3_18_xor1;
  assign s_csamul_cla32_fa2_19_xor1 = s_csamul_cla32_fa2_19_xor0 ^ s_csamul_cla32_fa2_18_or0;
  assign s_csamul_cla32_fa2_19_and1 = s_csamul_cla32_fa2_19_xor0 & s_csamul_cla32_fa2_18_or0;
  assign s_csamul_cla32_fa2_19_or0 = s_csamul_cla32_fa2_19_and0 | s_csamul_cla32_fa2_19_and1;
  assign s_csamul_cla32_and3_19 = a[3] & b[19];
  assign s_csamul_cla32_fa3_19_xor0 = s_csamul_cla32_and3_19 ^ s_csamul_cla32_fa4_18_xor1;
  assign s_csamul_cla32_fa3_19_and0 = s_csamul_cla32_and3_19 & s_csamul_cla32_fa4_18_xor1;
  assign s_csamul_cla32_fa3_19_xor1 = s_csamul_cla32_fa3_19_xor0 ^ s_csamul_cla32_fa3_18_or0;
  assign s_csamul_cla32_fa3_19_and1 = s_csamul_cla32_fa3_19_xor0 & s_csamul_cla32_fa3_18_or0;
  assign s_csamul_cla32_fa3_19_or0 = s_csamul_cla32_fa3_19_and0 | s_csamul_cla32_fa3_19_and1;
  assign s_csamul_cla32_and4_19 = a[4] & b[19];
  assign s_csamul_cla32_fa4_19_xor0 = s_csamul_cla32_and4_19 ^ s_csamul_cla32_fa5_18_xor1;
  assign s_csamul_cla32_fa4_19_and0 = s_csamul_cla32_and4_19 & s_csamul_cla32_fa5_18_xor1;
  assign s_csamul_cla32_fa4_19_xor1 = s_csamul_cla32_fa4_19_xor0 ^ s_csamul_cla32_fa4_18_or0;
  assign s_csamul_cla32_fa4_19_and1 = s_csamul_cla32_fa4_19_xor0 & s_csamul_cla32_fa4_18_or0;
  assign s_csamul_cla32_fa4_19_or0 = s_csamul_cla32_fa4_19_and0 | s_csamul_cla32_fa4_19_and1;
  assign s_csamul_cla32_and5_19 = a[5] & b[19];
  assign s_csamul_cla32_fa5_19_xor0 = s_csamul_cla32_and5_19 ^ s_csamul_cla32_fa6_18_xor1;
  assign s_csamul_cla32_fa5_19_and0 = s_csamul_cla32_and5_19 & s_csamul_cla32_fa6_18_xor1;
  assign s_csamul_cla32_fa5_19_xor1 = s_csamul_cla32_fa5_19_xor0 ^ s_csamul_cla32_fa5_18_or0;
  assign s_csamul_cla32_fa5_19_and1 = s_csamul_cla32_fa5_19_xor0 & s_csamul_cla32_fa5_18_or0;
  assign s_csamul_cla32_fa5_19_or0 = s_csamul_cla32_fa5_19_and0 | s_csamul_cla32_fa5_19_and1;
  assign s_csamul_cla32_and6_19 = a[6] & b[19];
  assign s_csamul_cla32_fa6_19_xor0 = s_csamul_cla32_and6_19 ^ s_csamul_cla32_fa7_18_xor1;
  assign s_csamul_cla32_fa6_19_and0 = s_csamul_cla32_and6_19 & s_csamul_cla32_fa7_18_xor1;
  assign s_csamul_cla32_fa6_19_xor1 = s_csamul_cla32_fa6_19_xor0 ^ s_csamul_cla32_fa6_18_or0;
  assign s_csamul_cla32_fa6_19_and1 = s_csamul_cla32_fa6_19_xor0 & s_csamul_cla32_fa6_18_or0;
  assign s_csamul_cla32_fa6_19_or0 = s_csamul_cla32_fa6_19_and0 | s_csamul_cla32_fa6_19_and1;
  assign s_csamul_cla32_and7_19 = a[7] & b[19];
  assign s_csamul_cla32_fa7_19_xor0 = s_csamul_cla32_and7_19 ^ s_csamul_cla32_fa8_18_xor1;
  assign s_csamul_cla32_fa7_19_and0 = s_csamul_cla32_and7_19 & s_csamul_cla32_fa8_18_xor1;
  assign s_csamul_cla32_fa7_19_xor1 = s_csamul_cla32_fa7_19_xor0 ^ s_csamul_cla32_fa7_18_or0;
  assign s_csamul_cla32_fa7_19_and1 = s_csamul_cla32_fa7_19_xor0 & s_csamul_cla32_fa7_18_or0;
  assign s_csamul_cla32_fa7_19_or0 = s_csamul_cla32_fa7_19_and0 | s_csamul_cla32_fa7_19_and1;
  assign s_csamul_cla32_and8_19 = a[8] & b[19];
  assign s_csamul_cla32_fa8_19_xor0 = s_csamul_cla32_and8_19 ^ s_csamul_cla32_fa9_18_xor1;
  assign s_csamul_cla32_fa8_19_and0 = s_csamul_cla32_and8_19 & s_csamul_cla32_fa9_18_xor1;
  assign s_csamul_cla32_fa8_19_xor1 = s_csamul_cla32_fa8_19_xor0 ^ s_csamul_cla32_fa8_18_or0;
  assign s_csamul_cla32_fa8_19_and1 = s_csamul_cla32_fa8_19_xor0 & s_csamul_cla32_fa8_18_or0;
  assign s_csamul_cla32_fa8_19_or0 = s_csamul_cla32_fa8_19_and0 | s_csamul_cla32_fa8_19_and1;
  assign s_csamul_cla32_and9_19 = a[9] & b[19];
  assign s_csamul_cla32_fa9_19_xor0 = s_csamul_cla32_and9_19 ^ s_csamul_cla32_fa10_18_xor1;
  assign s_csamul_cla32_fa9_19_and0 = s_csamul_cla32_and9_19 & s_csamul_cla32_fa10_18_xor1;
  assign s_csamul_cla32_fa9_19_xor1 = s_csamul_cla32_fa9_19_xor0 ^ s_csamul_cla32_fa9_18_or0;
  assign s_csamul_cla32_fa9_19_and1 = s_csamul_cla32_fa9_19_xor0 & s_csamul_cla32_fa9_18_or0;
  assign s_csamul_cla32_fa9_19_or0 = s_csamul_cla32_fa9_19_and0 | s_csamul_cla32_fa9_19_and1;
  assign s_csamul_cla32_and10_19 = a[10] & b[19];
  assign s_csamul_cla32_fa10_19_xor0 = s_csamul_cla32_and10_19 ^ s_csamul_cla32_fa11_18_xor1;
  assign s_csamul_cla32_fa10_19_and0 = s_csamul_cla32_and10_19 & s_csamul_cla32_fa11_18_xor1;
  assign s_csamul_cla32_fa10_19_xor1 = s_csamul_cla32_fa10_19_xor0 ^ s_csamul_cla32_fa10_18_or0;
  assign s_csamul_cla32_fa10_19_and1 = s_csamul_cla32_fa10_19_xor0 & s_csamul_cla32_fa10_18_or0;
  assign s_csamul_cla32_fa10_19_or0 = s_csamul_cla32_fa10_19_and0 | s_csamul_cla32_fa10_19_and1;
  assign s_csamul_cla32_and11_19 = a[11] & b[19];
  assign s_csamul_cla32_fa11_19_xor0 = s_csamul_cla32_and11_19 ^ s_csamul_cla32_fa12_18_xor1;
  assign s_csamul_cla32_fa11_19_and0 = s_csamul_cla32_and11_19 & s_csamul_cla32_fa12_18_xor1;
  assign s_csamul_cla32_fa11_19_xor1 = s_csamul_cla32_fa11_19_xor0 ^ s_csamul_cla32_fa11_18_or0;
  assign s_csamul_cla32_fa11_19_and1 = s_csamul_cla32_fa11_19_xor0 & s_csamul_cla32_fa11_18_or0;
  assign s_csamul_cla32_fa11_19_or0 = s_csamul_cla32_fa11_19_and0 | s_csamul_cla32_fa11_19_and1;
  assign s_csamul_cla32_and12_19 = a[12] & b[19];
  assign s_csamul_cla32_fa12_19_xor0 = s_csamul_cla32_and12_19 ^ s_csamul_cla32_fa13_18_xor1;
  assign s_csamul_cla32_fa12_19_and0 = s_csamul_cla32_and12_19 & s_csamul_cla32_fa13_18_xor1;
  assign s_csamul_cla32_fa12_19_xor1 = s_csamul_cla32_fa12_19_xor0 ^ s_csamul_cla32_fa12_18_or0;
  assign s_csamul_cla32_fa12_19_and1 = s_csamul_cla32_fa12_19_xor0 & s_csamul_cla32_fa12_18_or0;
  assign s_csamul_cla32_fa12_19_or0 = s_csamul_cla32_fa12_19_and0 | s_csamul_cla32_fa12_19_and1;
  assign s_csamul_cla32_and13_19 = a[13] & b[19];
  assign s_csamul_cla32_fa13_19_xor0 = s_csamul_cla32_and13_19 ^ s_csamul_cla32_fa14_18_xor1;
  assign s_csamul_cla32_fa13_19_and0 = s_csamul_cla32_and13_19 & s_csamul_cla32_fa14_18_xor1;
  assign s_csamul_cla32_fa13_19_xor1 = s_csamul_cla32_fa13_19_xor0 ^ s_csamul_cla32_fa13_18_or0;
  assign s_csamul_cla32_fa13_19_and1 = s_csamul_cla32_fa13_19_xor0 & s_csamul_cla32_fa13_18_or0;
  assign s_csamul_cla32_fa13_19_or0 = s_csamul_cla32_fa13_19_and0 | s_csamul_cla32_fa13_19_and1;
  assign s_csamul_cla32_and14_19 = a[14] & b[19];
  assign s_csamul_cla32_fa14_19_xor0 = s_csamul_cla32_and14_19 ^ s_csamul_cla32_fa15_18_xor1;
  assign s_csamul_cla32_fa14_19_and0 = s_csamul_cla32_and14_19 & s_csamul_cla32_fa15_18_xor1;
  assign s_csamul_cla32_fa14_19_xor1 = s_csamul_cla32_fa14_19_xor0 ^ s_csamul_cla32_fa14_18_or0;
  assign s_csamul_cla32_fa14_19_and1 = s_csamul_cla32_fa14_19_xor0 & s_csamul_cla32_fa14_18_or0;
  assign s_csamul_cla32_fa14_19_or0 = s_csamul_cla32_fa14_19_and0 | s_csamul_cla32_fa14_19_and1;
  assign s_csamul_cla32_and15_19 = a[15] & b[19];
  assign s_csamul_cla32_fa15_19_xor0 = s_csamul_cla32_and15_19 ^ s_csamul_cla32_fa16_18_xor1;
  assign s_csamul_cla32_fa15_19_and0 = s_csamul_cla32_and15_19 & s_csamul_cla32_fa16_18_xor1;
  assign s_csamul_cla32_fa15_19_xor1 = s_csamul_cla32_fa15_19_xor0 ^ s_csamul_cla32_fa15_18_or0;
  assign s_csamul_cla32_fa15_19_and1 = s_csamul_cla32_fa15_19_xor0 & s_csamul_cla32_fa15_18_or0;
  assign s_csamul_cla32_fa15_19_or0 = s_csamul_cla32_fa15_19_and0 | s_csamul_cla32_fa15_19_and1;
  assign s_csamul_cla32_and16_19 = a[16] & b[19];
  assign s_csamul_cla32_fa16_19_xor0 = s_csamul_cla32_and16_19 ^ s_csamul_cla32_fa17_18_xor1;
  assign s_csamul_cla32_fa16_19_and0 = s_csamul_cla32_and16_19 & s_csamul_cla32_fa17_18_xor1;
  assign s_csamul_cla32_fa16_19_xor1 = s_csamul_cla32_fa16_19_xor0 ^ s_csamul_cla32_fa16_18_or0;
  assign s_csamul_cla32_fa16_19_and1 = s_csamul_cla32_fa16_19_xor0 & s_csamul_cla32_fa16_18_or0;
  assign s_csamul_cla32_fa16_19_or0 = s_csamul_cla32_fa16_19_and0 | s_csamul_cla32_fa16_19_and1;
  assign s_csamul_cla32_and17_19 = a[17] & b[19];
  assign s_csamul_cla32_fa17_19_xor0 = s_csamul_cla32_and17_19 ^ s_csamul_cla32_fa18_18_xor1;
  assign s_csamul_cla32_fa17_19_and0 = s_csamul_cla32_and17_19 & s_csamul_cla32_fa18_18_xor1;
  assign s_csamul_cla32_fa17_19_xor1 = s_csamul_cla32_fa17_19_xor0 ^ s_csamul_cla32_fa17_18_or0;
  assign s_csamul_cla32_fa17_19_and1 = s_csamul_cla32_fa17_19_xor0 & s_csamul_cla32_fa17_18_or0;
  assign s_csamul_cla32_fa17_19_or0 = s_csamul_cla32_fa17_19_and0 | s_csamul_cla32_fa17_19_and1;
  assign s_csamul_cla32_and18_19 = a[18] & b[19];
  assign s_csamul_cla32_fa18_19_xor0 = s_csamul_cla32_and18_19 ^ s_csamul_cla32_fa19_18_xor1;
  assign s_csamul_cla32_fa18_19_and0 = s_csamul_cla32_and18_19 & s_csamul_cla32_fa19_18_xor1;
  assign s_csamul_cla32_fa18_19_xor1 = s_csamul_cla32_fa18_19_xor0 ^ s_csamul_cla32_fa18_18_or0;
  assign s_csamul_cla32_fa18_19_and1 = s_csamul_cla32_fa18_19_xor0 & s_csamul_cla32_fa18_18_or0;
  assign s_csamul_cla32_fa18_19_or0 = s_csamul_cla32_fa18_19_and0 | s_csamul_cla32_fa18_19_and1;
  assign s_csamul_cla32_and19_19 = a[19] & b[19];
  assign s_csamul_cla32_fa19_19_xor0 = s_csamul_cla32_and19_19 ^ s_csamul_cla32_fa20_18_xor1;
  assign s_csamul_cla32_fa19_19_and0 = s_csamul_cla32_and19_19 & s_csamul_cla32_fa20_18_xor1;
  assign s_csamul_cla32_fa19_19_xor1 = s_csamul_cla32_fa19_19_xor0 ^ s_csamul_cla32_fa19_18_or0;
  assign s_csamul_cla32_fa19_19_and1 = s_csamul_cla32_fa19_19_xor0 & s_csamul_cla32_fa19_18_or0;
  assign s_csamul_cla32_fa19_19_or0 = s_csamul_cla32_fa19_19_and0 | s_csamul_cla32_fa19_19_and1;
  assign s_csamul_cla32_and20_19 = a[20] & b[19];
  assign s_csamul_cla32_fa20_19_xor0 = s_csamul_cla32_and20_19 ^ s_csamul_cla32_fa21_18_xor1;
  assign s_csamul_cla32_fa20_19_and0 = s_csamul_cla32_and20_19 & s_csamul_cla32_fa21_18_xor1;
  assign s_csamul_cla32_fa20_19_xor1 = s_csamul_cla32_fa20_19_xor0 ^ s_csamul_cla32_fa20_18_or0;
  assign s_csamul_cla32_fa20_19_and1 = s_csamul_cla32_fa20_19_xor0 & s_csamul_cla32_fa20_18_or0;
  assign s_csamul_cla32_fa20_19_or0 = s_csamul_cla32_fa20_19_and0 | s_csamul_cla32_fa20_19_and1;
  assign s_csamul_cla32_and21_19 = a[21] & b[19];
  assign s_csamul_cla32_fa21_19_xor0 = s_csamul_cla32_and21_19 ^ s_csamul_cla32_fa22_18_xor1;
  assign s_csamul_cla32_fa21_19_and0 = s_csamul_cla32_and21_19 & s_csamul_cla32_fa22_18_xor1;
  assign s_csamul_cla32_fa21_19_xor1 = s_csamul_cla32_fa21_19_xor0 ^ s_csamul_cla32_fa21_18_or0;
  assign s_csamul_cla32_fa21_19_and1 = s_csamul_cla32_fa21_19_xor0 & s_csamul_cla32_fa21_18_or0;
  assign s_csamul_cla32_fa21_19_or0 = s_csamul_cla32_fa21_19_and0 | s_csamul_cla32_fa21_19_and1;
  assign s_csamul_cla32_and22_19 = a[22] & b[19];
  assign s_csamul_cla32_fa22_19_xor0 = s_csamul_cla32_and22_19 ^ s_csamul_cla32_fa23_18_xor1;
  assign s_csamul_cla32_fa22_19_and0 = s_csamul_cla32_and22_19 & s_csamul_cla32_fa23_18_xor1;
  assign s_csamul_cla32_fa22_19_xor1 = s_csamul_cla32_fa22_19_xor0 ^ s_csamul_cla32_fa22_18_or0;
  assign s_csamul_cla32_fa22_19_and1 = s_csamul_cla32_fa22_19_xor0 & s_csamul_cla32_fa22_18_or0;
  assign s_csamul_cla32_fa22_19_or0 = s_csamul_cla32_fa22_19_and0 | s_csamul_cla32_fa22_19_and1;
  assign s_csamul_cla32_and23_19 = a[23] & b[19];
  assign s_csamul_cla32_fa23_19_xor0 = s_csamul_cla32_and23_19 ^ s_csamul_cla32_fa24_18_xor1;
  assign s_csamul_cla32_fa23_19_and0 = s_csamul_cla32_and23_19 & s_csamul_cla32_fa24_18_xor1;
  assign s_csamul_cla32_fa23_19_xor1 = s_csamul_cla32_fa23_19_xor0 ^ s_csamul_cla32_fa23_18_or0;
  assign s_csamul_cla32_fa23_19_and1 = s_csamul_cla32_fa23_19_xor0 & s_csamul_cla32_fa23_18_or0;
  assign s_csamul_cla32_fa23_19_or0 = s_csamul_cla32_fa23_19_and0 | s_csamul_cla32_fa23_19_and1;
  assign s_csamul_cla32_and24_19 = a[24] & b[19];
  assign s_csamul_cla32_fa24_19_xor0 = s_csamul_cla32_and24_19 ^ s_csamul_cla32_fa25_18_xor1;
  assign s_csamul_cla32_fa24_19_and0 = s_csamul_cla32_and24_19 & s_csamul_cla32_fa25_18_xor1;
  assign s_csamul_cla32_fa24_19_xor1 = s_csamul_cla32_fa24_19_xor0 ^ s_csamul_cla32_fa24_18_or0;
  assign s_csamul_cla32_fa24_19_and1 = s_csamul_cla32_fa24_19_xor0 & s_csamul_cla32_fa24_18_or0;
  assign s_csamul_cla32_fa24_19_or0 = s_csamul_cla32_fa24_19_and0 | s_csamul_cla32_fa24_19_and1;
  assign s_csamul_cla32_and25_19 = a[25] & b[19];
  assign s_csamul_cla32_fa25_19_xor0 = s_csamul_cla32_and25_19 ^ s_csamul_cla32_fa26_18_xor1;
  assign s_csamul_cla32_fa25_19_and0 = s_csamul_cla32_and25_19 & s_csamul_cla32_fa26_18_xor1;
  assign s_csamul_cla32_fa25_19_xor1 = s_csamul_cla32_fa25_19_xor0 ^ s_csamul_cla32_fa25_18_or0;
  assign s_csamul_cla32_fa25_19_and1 = s_csamul_cla32_fa25_19_xor0 & s_csamul_cla32_fa25_18_or0;
  assign s_csamul_cla32_fa25_19_or0 = s_csamul_cla32_fa25_19_and0 | s_csamul_cla32_fa25_19_and1;
  assign s_csamul_cla32_and26_19 = a[26] & b[19];
  assign s_csamul_cla32_fa26_19_xor0 = s_csamul_cla32_and26_19 ^ s_csamul_cla32_fa27_18_xor1;
  assign s_csamul_cla32_fa26_19_and0 = s_csamul_cla32_and26_19 & s_csamul_cla32_fa27_18_xor1;
  assign s_csamul_cla32_fa26_19_xor1 = s_csamul_cla32_fa26_19_xor0 ^ s_csamul_cla32_fa26_18_or0;
  assign s_csamul_cla32_fa26_19_and1 = s_csamul_cla32_fa26_19_xor0 & s_csamul_cla32_fa26_18_or0;
  assign s_csamul_cla32_fa26_19_or0 = s_csamul_cla32_fa26_19_and0 | s_csamul_cla32_fa26_19_and1;
  assign s_csamul_cla32_and27_19 = a[27] & b[19];
  assign s_csamul_cla32_fa27_19_xor0 = s_csamul_cla32_and27_19 ^ s_csamul_cla32_fa28_18_xor1;
  assign s_csamul_cla32_fa27_19_and0 = s_csamul_cla32_and27_19 & s_csamul_cla32_fa28_18_xor1;
  assign s_csamul_cla32_fa27_19_xor1 = s_csamul_cla32_fa27_19_xor0 ^ s_csamul_cla32_fa27_18_or0;
  assign s_csamul_cla32_fa27_19_and1 = s_csamul_cla32_fa27_19_xor0 & s_csamul_cla32_fa27_18_or0;
  assign s_csamul_cla32_fa27_19_or0 = s_csamul_cla32_fa27_19_and0 | s_csamul_cla32_fa27_19_and1;
  assign s_csamul_cla32_and28_19 = a[28] & b[19];
  assign s_csamul_cla32_fa28_19_xor0 = s_csamul_cla32_and28_19 ^ s_csamul_cla32_fa29_18_xor1;
  assign s_csamul_cla32_fa28_19_and0 = s_csamul_cla32_and28_19 & s_csamul_cla32_fa29_18_xor1;
  assign s_csamul_cla32_fa28_19_xor1 = s_csamul_cla32_fa28_19_xor0 ^ s_csamul_cla32_fa28_18_or0;
  assign s_csamul_cla32_fa28_19_and1 = s_csamul_cla32_fa28_19_xor0 & s_csamul_cla32_fa28_18_or0;
  assign s_csamul_cla32_fa28_19_or0 = s_csamul_cla32_fa28_19_and0 | s_csamul_cla32_fa28_19_and1;
  assign s_csamul_cla32_and29_19 = a[29] & b[19];
  assign s_csamul_cla32_fa29_19_xor0 = s_csamul_cla32_and29_19 ^ s_csamul_cla32_fa30_18_xor1;
  assign s_csamul_cla32_fa29_19_and0 = s_csamul_cla32_and29_19 & s_csamul_cla32_fa30_18_xor1;
  assign s_csamul_cla32_fa29_19_xor1 = s_csamul_cla32_fa29_19_xor0 ^ s_csamul_cla32_fa29_18_or0;
  assign s_csamul_cla32_fa29_19_and1 = s_csamul_cla32_fa29_19_xor0 & s_csamul_cla32_fa29_18_or0;
  assign s_csamul_cla32_fa29_19_or0 = s_csamul_cla32_fa29_19_and0 | s_csamul_cla32_fa29_19_and1;
  assign s_csamul_cla32_and30_19 = a[30] & b[19];
  assign s_csamul_cla32_fa30_19_xor0 = s_csamul_cla32_and30_19 ^ s_csamul_cla32_ha31_18_xor0;
  assign s_csamul_cla32_fa30_19_and0 = s_csamul_cla32_and30_19 & s_csamul_cla32_ha31_18_xor0;
  assign s_csamul_cla32_fa30_19_xor1 = s_csamul_cla32_fa30_19_xor0 ^ s_csamul_cla32_fa30_18_or0;
  assign s_csamul_cla32_fa30_19_and1 = s_csamul_cla32_fa30_19_xor0 & s_csamul_cla32_fa30_18_or0;
  assign s_csamul_cla32_fa30_19_or0 = s_csamul_cla32_fa30_19_and0 | s_csamul_cla32_fa30_19_and1;
  assign s_csamul_cla32_nand31_19 = ~(a[31] & b[19]);
  assign s_csamul_cla32_ha31_19_xor0 = s_csamul_cla32_nand31_19 ^ s_csamul_cla32_ha31_18_and0;
  assign s_csamul_cla32_ha31_19_and0 = s_csamul_cla32_nand31_19 & s_csamul_cla32_ha31_18_and0;
  assign s_csamul_cla32_and0_20 = a[0] & b[20];
  assign s_csamul_cla32_fa0_20_xor0 = s_csamul_cla32_and0_20 ^ s_csamul_cla32_fa1_19_xor1;
  assign s_csamul_cla32_fa0_20_and0 = s_csamul_cla32_and0_20 & s_csamul_cla32_fa1_19_xor1;
  assign s_csamul_cla32_fa0_20_xor1 = s_csamul_cla32_fa0_20_xor0 ^ s_csamul_cla32_fa0_19_or0;
  assign s_csamul_cla32_fa0_20_and1 = s_csamul_cla32_fa0_20_xor0 & s_csamul_cla32_fa0_19_or0;
  assign s_csamul_cla32_fa0_20_or0 = s_csamul_cla32_fa0_20_and0 | s_csamul_cla32_fa0_20_and1;
  assign s_csamul_cla32_and1_20 = a[1] & b[20];
  assign s_csamul_cla32_fa1_20_xor0 = s_csamul_cla32_and1_20 ^ s_csamul_cla32_fa2_19_xor1;
  assign s_csamul_cla32_fa1_20_and0 = s_csamul_cla32_and1_20 & s_csamul_cla32_fa2_19_xor1;
  assign s_csamul_cla32_fa1_20_xor1 = s_csamul_cla32_fa1_20_xor0 ^ s_csamul_cla32_fa1_19_or0;
  assign s_csamul_cla32_fa1_20_and1 = s_csamul_cla32_fa1_20_xor0 & s_csamul_cla32_fa1_19_or0;
  assign s_csamul_cla32_fa1_20_or0 = s_csamul_cla32_fa1_20_and0 | s_csamul_cla32_fa1_20_and1;
  assign s_csamul_cla32_and2_20 = a[2] & b[20];
  assign s_csamul_cla32_fa2_20_xor0 = s_csamul_cla32_and2_20 ^ s_csamul_cla32_fa3_19_xor1;
  assign s_csamul_cla32_fa2_20_and0 = s_csamul_cla32_and2_20 & s_csamul_cla32_fa3_19_xor1;
  assign s_csamul_cla32_fa2_20_xor1 = s_csamul_cla32_fa2_20_xor0 ^ s_csamul_cla32_fa2_19_or0;
  assign s_csamul_cla32_fa2_20_and1 = s_csamul_cla32_fa2_20_xor0 & s_csamul_cla32_fa2_19_or0;
  assign s_csamul_cla32_fa2_20_or0 = s_csamul_cla32_fa2_20_and0 | s_csamul_cla32_fa2_20_and1;
  assign s_csamul_cla32_and3_20 = a[3] & b[20];
  assign s_csamul_cla32_fa3_20_xor0 = s_csamul_cla32_and3_20 ^ s_csamul_cla32_fa4_19_xor1;
  assign s_csamul_cla32_fa3_20_and0 = s_csamul_cla32_and3_20 & s_csamul_cla32_fa4_19_xor1;
  assign s_csamul_cla32_fa3_20_xor1 = s_csamul_cla32_fa3_20_xor0 ^ s_csamul_cla32_fa3_19_or0;
  assign s_csamul_cla32_fa3_20_and1 = s_csamul_cla32_fa3_20_xor0 & s_csamul_cla32_fa3_19_or0;
  assign s_csamul_cla32_fa3_20_or0 = s_csamul_cla32_fa3_20_and0 | s_csamul_cla32_fa3_20_and1;
  assign s_csamul_cla32_and4_20 = a[4] & b[20];
  assign s_csamul_cla32_fa4_20_xor0 = s_csamul_cla32_and4_20 ^ s_csamul_cla32_fa5_19_xor1;
  assign s_csamul_cla32_fa4_20_and0 = s_csamul_cla32_and4_20 & s_csamul_cla32_fa5_19_xor1;
  assign s_csamul_cla32_fa4_20_xor1 = s_csamul_cla32_fa4_20_xor0 ^ s_csamul_cla32_fa4_19_or0;
  assign s_csamul_cla32_fa4_20_and1 = s_csamul_cla32_fa4_20_xor0 & s_csamul_cla32_fa4_19_or0;
  assign s_csamul_cla32_fa4_20_or0 = s_csamul_cla32_fa4_20_and0 | s_csamul_cla32_fa4_20_and1;
  assign s_csamul_cla32_and5_20 = a[5] & b[20];
  assign s_csamul_cla32_fa5_20_xor0 = s_csamul_cla32_and5_20 ^ s_csamul_cla32_fa6_19_xor1;
  assign s_csamul_cla32_fa5_20_and0 = s_csamul_cla32_and5_20 & s_csamul_cla32_fa6_19_xor1;
  assign s_csamul_cla32_fa5_20_xor1 = s_csamul_cla32_fa5_20_xor0 ^ s_csamul_cla32_fa5_19_or0;
  assign s_csamul_cla32_fa5_20_and1 = s_csamul_cla32_fa5_20_xor0 & s_csamul_cla32_fa5_19_or0;
  assign s_csamul_cla32_fa5_20_or0 = s_csamul_cla32_fa5_20_and0 | s_csamul_cla32_fa5_20_and1;
  assign s_csamul_cla32_and6_20 = a[6] & b[20];
  assign s_csamul_cla32_fa6_20_xor0 = s_csamul_cla32_and6_20 ^ s_csamul_cla32_fa7_19_xor1;
  assign s_csamul_cla32_fa6_20_and0 = s_csamul_cla32_and6_20 & s_csamul_cla32_fa7_19_xor1;
  assign s_csamul_cla32_fa6_20_xor1 = s_csamul_cla32_fa6_20_xor0 ^ s_csamul_cla32_fa6_19_or0;
  assign s_csamul_cla32_fa6_20_and1 = s_csamul_cla32_fa6_20_xor0 & s_csamul_cla32_fa6_19_or0;
  assign s_csamul_cla32_fa6_20_or0 = s_csamul_cla32_fa6_20_and0 | s_csamul_cla32_fa6_20_and1;
  assign s_csamul_cla32_and7_20 = a[7] & b[20];
  assign s_csamul_cla32_fa7_20_xor0 = s_csamul_cla32_and7_20 ^ s_csamul_cla32_fa8_19_xor1;
  assign s_csamul_cla32_fa7_20_and0 = s_csamul_cla32_and7_20 & s_csamul_cla32_fa8_19_xor1;
  assign s_csamul_cla32_fa7_20_xor1 = s_csamul_cla32_fa7_20_xor0 ^ s_csamul_cla32_fa7_19_or0;
  assign s_csamul_cla32_fa7_20_and1 = s_csamul_cla32_fa7_20_xor0 & s_csamul_cla32_fa7_19_or0;
  assign s_csamul_cla32_fa7_20_or0 = s_csamul_cla32_fa7_20_and0 | s_csamul_cla32_fa7_20_and1;
  assign s_csamul_cla32_and8_20 = a[8] & b[20];
  assign s_csamul_cla32_fa8_20_xor0 = s_csamul_cla32_and8_20 ^ s_csamul_cla32_fa9_19_xor1;
  assign s_csamul_cla32_fa8_20_and0 = s_csamul_cla32_and8_20 & s_csamul_cla32_fa9_19_xor1;
  assign s_csamul_cla32_fa8_20_xor1 = s_csamul_cla32_fa8_20_xor0 ^ s_csamul_cla32_fa8_19_or0;
  assign s_csamul_cla32_fa8_20_and1 = s_csamul_cla32_fa8_20_xor0 & s_csamul_cla32_fa8_19_or0;
  assign s_csamul_cla32_fa8_20_or0 = s_csamul_cla32_fa8_20_and0 | s_csamul_cla32_fa8_20_and1;
  assign s_csamul_cla32_and9_20 = a[9] & b[20];
  assign s_csamul_cla32_fa9_20_xor0 = s_csamul_cla32_and9_20 ^ s_csamul_cla32_fa10_19_xor1;
  assign s_csamul_cla32_fa9_20_and0 = s_csamul_cla32_and9_20 & s_csamul_cla32_fa10_19_xor1;
  assign s_csamul_cla32_fa9_20_xor1 = s_csamul_cla32_fa9_20_xor0 ^ s_csamul_cla32_fa9_19_or0;
  assign s_csamul_cla32_fa9_20_and1 = s_csamul_cla32_fa9_20_xor0 & s_csamul_cla32_fa9_19_or0;
  assign s_csamul_cla32_fa9_20_or0 = s_csamul_cla32_fa9_20_and0 | s_csamul_cla32_fa9_20_and1;
  assign s_csamul_cla32_and10_20 = a[10] & b[20];
  assign s_csamul_cla32_fa10_20_xor0 = s_csamul_cla32_and10_20 ^ s_csamul_cla32_fa11_19_xor1;
  assign s_csamul_cla32_fa10_20_and0 = s_csamul_cla32_and10_20 & s_csamul_cla32_fa11_19_xor1;
  assign s_csamul_cla32_fa10_20_xor1 = s_csamul_cla32_fa10_20_xor0 ^ s_csamul_cla32_fa10_19_or0;
  assign s_csamul_cla32_fa10_20_and1 = s_csamul_cla32_fa10_20_xor0 & s_csamul_cla32_fa10_19_or0;
  assign s_csamul_cla32_fa10_20_or0 = s_csamul_cla32_fa10_20_and0 | s_csamul_cla32_fa10_20_and1;
  assign s_csamul_cla32_and11_20 = a[11] & b[20];
  assign s_csamul_cla32_fa11_20_xor0 = s_csamul_cla32_and11_20 ^ s_csamul_cla32_fa12_19_xor1;
  assign s_csamul_cla32_fa11_20_and0 = s_csamul_cla32_and11_20 & s_csamul_cla32_fa12_19_xor1;
  assign s_csamul_cla32_fa11_20_xor1 = s_csamul_cla32_fa11_20_xor0 ^ s_csamul_cla32_fa11_19_or0;
  assign s_csamul_cla32_fa11_20_and1 = s_csamul_cla32_fa11_20_xor0 & s_csamul_cla32_fa11_19_or0;
  assign s_csamul_cla32_fa11_20_or0 = s_csamul_cla32_fa11_20_and0 | s_csamul_cla32_fa11_20_and1;
  assign s_csamul_cla32_and12_20 = a[12] & b[20];
  assign s_csamul_cla32_fa12_20_xor0 = s_csamul_cla32_and12_20 ^ s_csamul_cla32_fa13_19_xor1;
  assign s_csamul_cla32_fa12_20_and0 = s_csamul_cla32_and12_20 & s_csamul_cla32_fa13_19_xor1;
  assign s_csamul_cla32_fa12_20_xor1 = s_csamul_cla32_fa12_20_xor0 ^ s_csamul_cla32_fa12_19_or0;
  assign s_csamul_cla32_fa12_20_and1 = s_csamul_cla32_fa12_20_xor0 & s_csamul_cla32_fa12_19_or0;
  assign s_csamul_cla32_fa12_20_or0 = s_csamul_cla32_fa12_20_and0 | s_csamul_cla32_fa12_20_and1;
  assign s_csamul_cla32_and13_20 = a[13] & b[20];
  assign s_csamul_cla32_fa13_20_xor0 = s_csamul_cla32_and13_20 ^ s_csamul_cla32_fa14_19_xor1;
  assign s_csamul_cla32_fa13_20_and0 = s_csamul_cla32_and13_20 & s_csamul_cla32_fa14_19_xor1;
  assign s_csamul_cla32_fa13_20_xor1 = s_csamul_cla32_fa13_20_xor0 ^ s_csamul_cla32_fa13_19_or0;
  assign s_csamul_cla32_fa13_20_and1 = s_csamul_cla32_fa13_20_xor0 & s_csamul_cla32_fa13_19_or0;
  assign s_csamul_cla32_fa13_20_or0 = s_csamul_cla32_fa13_20_and0 | s_csamul_cla32_fa13_20_and1;
  assign s_csamul_cla32_and14_20 = a[14] & b[20];
  assign s_csamul_cla32_fa14_20_xor0 = s_csamul_cla32_and14_20 ^ s_csamul_cla32_fa15_19_xor1;
  assign s_csamul_cla32_fa14_20_and0 = s_csamul_cla32_and14_20 & s_csamul_cla32_fa15_19_xor1;
  assign s_csamul_cla32_fa14_20_xor1 = s_csamul_cla32_fa14_20_xor0 ^ s_csamul_cla32_fa14_19_or0;
  assign s_csamul_cla32_fa14_20_and1 = s_csamul_cla32_fa14_20_xor0 & s_csamul_cla32_fa14_19_or0;
  assign s_csamul_cla32_fa14_20_or0 = s_csamul_cla32_fa14_20_and0 | s_csamul_cla32_fa14_20_and1;
  assign s_csamul_cla32_and15_20 = a[15] & b[20];
  assign s_csamul_cla32_fa15_20_xor0 = s_csamul_cla32_and15_20 ^ s_csamul_cla32_fa16_19_xor1;
  assign s_csamul_cla32_fa15_20_and0 = s_csamul_cla32_and15_20 & s_csamul_cla32_fa16_19_xor1;
  assign s_csamul_cla32_fa15_20_xor1 = s_csamul_cla32_fa15_20_xor0 ^ s_csamul_cla32_fa15_19_or0;
  assign s_csamul_cla32_fa15_20_and1 = s_csamul_cla32_fa15_20_xor0 & s_csamul_cla32_fa15_19_or0;
  assign s_csamul_cla32_fa15_20_or0 = s_csamul_cla32_fa15_20_and0 | s_csamul_cla32_fa15_20_and1;
  assign s_csamul_cla32_and16_20 = a[16] & b[20];
  assign s_csamul_cla32_fa16_20_xor0 = s_csamul_cla32_and16_20 ^ s_csamul_cla32_fa17_19_xor1;
  assign s_csamul_cla32_fa16_20_and0 = s_csamul_cla32_and16_20 & s_csamul_cla32_fa17_19_xor1;
  assign s_csamul_cla32_fa16_20_xor1 = s_csamul_cla32_fa16_20_xor0 ^ s_csamul_cla32_fa16_19_or0;
  assign s_csamul_cla32_fa16_20_and1 = s_csamul_cla32_fa16_20_xor0 & s_csamul_cla32_fa16_19_or0;
  assign s_csamul_cla32_fa16_20_or0 = s_csamul_cla32_fa16_20_and0 | s_csamul_cla32_fa16_20_and1;
  assign s_csamul_cla32_and17_20 = a[17] & b[20];
  assign s_csamul_cla32_fa17_20_xor0 = s_csamul_cla32_and17_20 ^ s_csamul_cla32_fa18_19_xor1;
  assign s_csamul_cla32_fa17_20_and0 = s_csamul_cla32_and17_20 & s_csamul_cla32_fa18_19_xor1;
  assign s_csamul_cla32_fa17_20_xor1 = s_csamul_cla32_fa17_20_xor0 ^ s_csamul_cla32_fa17_19_or0;
  assign s_csamul_cla32_fa17_20_and1 = s_csamul_cla32_fa17_20_xor0 & s_csamul_cla32_fa17_19_or0;
  assign s_csamul_cla32_fa17_20_or0 = s_csamul_cla32_fa17_20_and0 | s_csamul_cla32_fa17_20_and1;
  assign s_csamul_cla32_and18_20 = a[18] & b[20];
  assign s_csamul_cla32_fa18_20_xor0 = s_csamul_cla32_and18_20 ^ s_csamul_cla32_fa19_19_xor1;
  assign s_csamul_cla32_fa18_20_and0 = s_csamul_cla32_and18_20 & s_csamul_cla32_fa19_19_xor1;
  assign s_csamul_cla32_fa18_20_xor1 = s_csamul_cla32_fa18_20_xor0 ^ s_csamul_cla32_fa18_19_or0;
  assign s_csamul_cla32_fa18_20_and1 = s_csamul_cla32_fa18_20_xor0 & s_csamul_cla32_fa18_19_or0;
  assign s_csamul_cla32_fa18_20_or0 = s_csamul_cla32_fa18_20_and0 | s_csamul_cla32_fa18_20_and1;
  assign s_csamul_cla32_and19_20 = a[19] & b[20];
  assign s_csamul_cla32_fa19_20_xor0 = s_csamul_cla32_and19_20 ^ s_csamul_cla32_fa20_19_xor1;
  assign s_csamul_cla32_fa19_20_and0 = s_csamul_cla32_and19_20 & s_csamul_cla32_fa20_19_xor1;
  assign s_csamul_cla32_fa19_20_xor1 = s_csamul_cla32_fa19_20_xor0 ^ s_csamul_cla32_fa19_19_or0;
  assign s_csamul_cla32_fa19_20_and1 = s_csamul_cla32_fa19_20_xor0 & s_csamul_cla32_fa19_19_or0;
  assign s_csamul_cla32_fa19_20_or0 = s_csamul_cla32_fa19_20_and0 | s_csamul_cla32_fa19_20_and1;
  assign s_csamul_cla32_and20_20 = a[20] & b[20];
  assign s_csamul_cla32_fa20_20_xor0 = s_csamul_cla32_and20_20 ^ s_csamul_cla32_fa21_19_xor1;
  assign s_csamul_cla32_fa20_20_and0 = s_csamul_cla32_and20_20 & s_csamul_cla32_fa21_19_xor1;
  assign s_csamul_cla32_fa20_20_xor1 = s_csamul_cla32_fa20_20_xor0 ^ s_csamul_cla32_fa20_19_or0;
  assign s_csamul_cla32_fa20_20_and1 = s_csamul_cla32_fa20_20_xor0 & s_csamul_cla32_fa20_19_or0;
  assign s_csamul_cla32_fa20_20_or0 = s_csamul_cla32_fa20_20_and0 | s_csamul_cla32_fa20_20_and1;
  assign s_csamul_cla32_and21_20 = a[21] & b[20];
  assign s_csamul_cla32_fa21_20_xor0 = s_csamul_cla32_and21_20 ^ s_csamul_cla32_fa22_19_xor1;
  assign s_csamul_cla32_fa21_20_and0 = s_csamul_cla32_and21_20 & s_csamul_cla32_fa22_19_xor1;
  assign s_csamul_cla32_fa21_20_xor1 = s_csamul_cla32_fa21_20_xor0 ^ s_csamul_cla32_fa21_19_or0;
  assign s_csamul_cla32_fa21_20_and1 = s_csamul_cla32_fa21_20_xor0 & s_csamul_cla32_fa21_19_or0;
  assign s_csamul_cla32_fa21_20_or0 = s_csamul_cla32_fa21_20_and0 | s_csamul_cla32_fa21_20_and1;
  assign s_csamul_cla32_and22_20 = a[22] & b[20];
  assign s_csamul_cla32_fa22_20_xor0 = s_csamul_cla32_and22_20 ^ s_csamul_cla32_fa23_19_xor1;
  assign s_csamul_cla32_fa22_20_and0 = s_csamul_cla32_and22_20 & s_csamul_cla32_fa23_19_xor1;
  assign s_csamul_cla32_fa22_20_xor1 = s_csamul_cla32_fa22_20_xor0 ^ s_csamul_cla32_fa22_19_or0;
  assign s_csamul_cla32_fa22_20_and1 = s_csamul_cla32_fa22_20_xor0 & s_csamul_cla32_fa22_19_or0;
  assign s_csamul_cla32_fa22_20_or0 = s_csamul_cla32_fa22_20_and0 | s_csamul_cla32_fa22_20_and1;
  assign s_csamul_cla32_and23_20 = a[23] & b[20];
  assign s_csamul_cla32_fa23_20_xor0 = s_csamul_cla32_and23_20 ^ s_csamul_cla32_fa24_19_xor1;
  assign s_csamul_cla32_fa23_20_and0 = s_csamul_cla32_and23_20 & s_csamul_cla32_fa24_19_xor1;
  assign s_csamul_cla32_fa23_20_xor1 = s_csamul_cla32_fa23_20_xor0 ^ s_csamul_cla32_fa23_19_or0;
  assign s_csamul_cla32_fa23_20_and1 = s_csamul_cla32_fa23_20_xor0 & s_csamul_cla32_fa23_19_or0;
  assign s_csamul_cla32_fa23_20_or0 = s_csamul_cla32_fa23_20_and0 | s_csamul_cla32_fa23_20_and1;
  assign s_csamul_cla32_and24_20 = a[24] & b[20];
  assign s_csamul_cla32_fa24_20_xor0 = s_csamul_cla32_and24_20 ^ s_csamul_cla32_fa25_19_xor1;
  assign s_csamul_cla32_fa24_20_and0 = s_csamul_cla32_and24_20 & s_csamul_cla32_fa25_19_xor1;
  assign s_csamul_cla32_fa24_20_xor1 = s_csamul_cla32_fa24_20_xor0 ^ s_csamul_cla32_fa24_19_or0;
  assign s_csamul_cla32_fa24_20_and1 = s_csamul_cla32_fa24_20_xor0 & s_csamul_cla32_fa24_19_or0;
  assign s_csamul_cla32_fa24_20_or0 = s_csamul_cla32_fa24_20_and0 | s_csamul_cla32_fa24_20_and1;
  assign s_csamul_cla32_and25_20 = a[25] & b[20];
  assign s_csamul_cla32_fa25_20_xor0 = s_csamul_cla32_and25_20 ^ s_csamul_cla32_fa26_19_xor1;
  assign s_csamul_cla32_fa25_20_and0 = s_csamul_cla32_and25_20 & s_csamul_cla32_fa26_19_xor1;
  assign s_csamul_cla32_fa25_20_xor1 = s_csamul_cla32_fa25_20_xor0 ^ s_csamul_cla32_fa25_19_or0;
  assign s_csamul_cla32_fa25_20_and1 = s_csamul_cla32_fa25_20_xor0 & s_csamul_cla32_fa25_19_or0;
  assign s_csamul_cla32_fa25_20_or0 = s_csamul_cla32_fa25_20_and0 | s_csamul_cla32_fa25_20_and1;
  assign s_csamul_cla32_and26_20 = a[26] & b[20];
  assign s_csamul_cla32_fa26_20_xor0 = s_csamul_cla32_and26_20 ^ s_csamul_cla32_fa27_19_xor1;
  assign s_csamul_cla32_fa26_20_and0 = s_csamul_cla32_and26_20 & s_csamul_cla32_fa27_19_xor1;
  assign s_csamul_cla32_fa26_20_xor1 = s_csamul_cla32_fa26_20_xor0 ^ s_csamul_cla32_fa26_19_or0;
  assign s_csamul_cla32_fa26_20_and1 = s_csamul_cla32_fa26_20_xor0 & s_csamul_cla32_fa26_19_or0;
  assign s_csamul_cla32_fa26_20_or0 = s_csamul_cla32_fa26_20_and0 | s_csamul_cla32_fa26_20_and1;
  assign s_csamul_cla32_and27_20 = a[27] & b[20];
  assign s_csamul_cla32_fa27_20_xor0 = s_csamul_cla32_and27_20 ^ s_csamul_cla32_fa28_19_xor1;
  assign s_csamul_cla32_fa27_20_and0 = s_csamul_cla32_and27_20 & s_csamul_cla32_fa28_19_xor1;
  assign s_csamul_cla32_fa27_20_xor1 = s_csamul_cla32_fa27_20_xor0 ^ s_csamul_cla32_fa27_19_or0;
  assign s_csamul_cla32_fa27_20_and1 = s_csamul_cla32_fa27_20_xor0 & s_csamul_cla32_fa27_19_or0;
  assign s_csamul_cla32_fa27_20_or0 = s_csamul_cla32_fa27_20_and0 | s_csamul_cla32_fa27_20_and1;
  assign s_csamul_cla32_and28_20 = a[28] & b[20];
  assign s_csamul_cla32_fa28_20_xor0 = s_csamul_cla32_and28_20 ^ s_csamul_cla32_fa29_19_xor1;
  assign s_csamul_cla32_fa28_20_and0 = s_csamul_cla32_and28_20 & s_csamul_cla32_fa29_19_xor1;
  assign s_csamul_cla32_fa28_20_xor1 = s_csamul_cla32_fa28_20_xor0 ^ s_csamul_cla32_fa28_19_or0;
  assign s_csamul_cla32_fa28_20_and1 = s_csamul_cla32_fa28_20_xor0 & s_csamul_cla32_fa28_19_or0;
  assign s_csamul_cla32_fa28_20_or0 = s_csamul_cla32_fa28_20_and0 | s_csamul_cla32_fa28_20_and1;
  assign s_csamul_cla32_and29_20 = a[29] & b[20];
  assign s_csamul_cla32_fa29_20_xor0 = s_csamul_cla32_and29_20 ^ s_csamul_cla32_fa30_19_xor1;
  assign s_csamul_cla32_fa29_20_and0 = s_csamul_cla32_and29_20 & s_csamul_cla32_fa30_19_xor1;
  assign s_csamul_cla32_fa29_20_xor1 = s_csamul_cla32_fa29_20_xor0 ^ s_csamul_cla32_fa29_19_or0;
  assign s_csamul_cla32_fa29_20_and1 = s_csamul_cla32_fa29_20_xor0 & s_csamul_cla32_fa29_19_or0;
  assign s_csamul_cla32_fa29_20_or0 = s_csamul_cla32_fa29_20_and0 | s_csamul_cla32_fa29_20_and1;
  assign s_csamul_cla32_and30_20 = a[30] & b[20];
  assign s_csamul_cla32_fa30_20_xor0 = s_csamul_cla32_and30_20 ^ s_csamul_cla32_ha31_19_xor0;
  assign s_csamul_cla32_fa30_20_and0 = s_csamul_cla32_and30_20 & s_csamul_cla32_ha31_19_xor0;
  assign s_csamul_cla32_fa30_20_xor1 = s_csamul_cla32_fa30_20_xor0 ^ s_csamul_cla32_fa30_19_or0;
  assign s_csamul_cla32_fa30_20_and1 = s_csamul_cla32_fa30_20_xor0 & s_csamul_cla32_fa30_19_or0;
  assign s_csamul_cla32_fa30_20_or0 = s_csamul_cla32_fa30_20_and0 | s_csamul_cla32_fa30_20_and1;
  assign s_csamul_cla32_nand31_20 = ~(a[31] & b[20]);
  assign s_csamul_cla32_ha31_20_xor0 = s_csamul_cla32_nand31_20 ^ s_csamul_cla32_ha31_19_and0;
  assign s_csamul_cla32_ha31_20_and0 = s_csamul_cla32_nand31_20 & s_csamul_cla32_ha31_19_and0;
  assign s_csamul_cla32_and0_21 = a[0] & b[21];
  assign s_csamul_cla32_fa0_21_xor0 = s_csamul_cla32_and0_21 ^ s_csamul_cla32_fa1_20_xor1;
  assign s_csamul_cla32_fa0_21_and0 = s_csamul_cla32_and0_21 & s_csamul_cla32_fa1_20_xor1;
  assign s_csamul_cla32_fa0_21_xor1 = s_csamul_cla32_fa0_21_xor0 ^ s_csamul_cla32_fa0_20_or0;
  assign s_csamul_cla32_fa0_21_and1 = s_csamul_cla32_fa0_21_xor0 & s_csamul_cla32_fa0_20_or0;
  assign s_csamul_cla32_fa0_21_or0 = s_csamul_cla32_fa0_21_and0 | s_csamul_cla32_fa0_21_and1;
  assign s_csamul_cla32_and1_21 = a[1] & b[21];
  assign s_csamul_cla32_fa1_21_xor0 = s_csamul_cla32_and1_21 ^ s_csamul_cla32_fa2_20_xor1;
  assign s_csamul_cla32_fa1_21_and0 = s_csamul_cla32_and1_21 & s_csamul_cla32_fa2_20_xor1;
  assign s_csamul_cla32_fa1_21_xor1 = s_csamul_cla32_fa1_21_xor0 ^ s_csamul_cla32_fa1_20_or0;
  assign s_csamul_cla32_fa1_21_and1 = s_csamul_cla32_fa1_21_xor0 & s_csamul_cla32_fa1_20_or0;
  assign s_csamul_cla32_fa1_21_or0 = s_csamul_cla32_fa1_21_and0 | s_csamul_cla32_fa1_21_and1;
  assign s_csamul_cla32_and2_21 = a[2] & b[21];
  assign s_csamul_cla32_fa2_21_xor0 = s_csamul_cla32_and2_21 ^ s_csamul_cla32_fa3_20_xor1;
  assign s_csamul_cla32_fa2_21_and0 = s_csamul_cla32_and2_21 & s_csamul_cla32_fa3_20_xor1;
  assign s_csamul_cla32_fa2_21_xor1 = s_csamul_cla32_fa2_21_xor0 ^ s_csamul_cla32_fa2_20_or0;
  assign s_csamul_cla32_fa2_21_and1 = s_csamul_cla32_fa2_21_xor0 & s_csamul_cla32_fa2_20_or0;
  assign s_csamul_cla32_fa2_21_or0 = s_csamul_cla32_fa2_21_and0 | s_csamul_cla32_fa2_21_and1;
  assign s_csamul_cla32_and3_21 = a[3] & b[21];
  assign s_csamul_cla32_fa3_21_xor0 = s_csamul_cla32_and3_21 ^ s_csamul_cla32_fa4_20_xor1;
  assign s_csamul_cla32_fa3_21_and0 = s_csamul_cla32_and3_21 & s_csamul_cla32_fa4_20_xor1;
  assign s_csamul_cla32_fa3_21_xor1 = s_csamul_cla32_fa3_21_xor0 ^ s_csamul_cla32_fa3_20_or0;
  assign s_csamul_cla32_fa3_21_and1 = s_csamul_cla32_fa3_21_xor0 & s_csamul_cla32_fa3_20_or0;
  assign s_csamul_cla32_fa3_21_or0 = s_csamul_cla32_fa3_21_and0 | s_csamul_cla32_fa3_21_and1;
  assign s_csamul_cla32_and4_21 = a[4] & b[21];
  assign s_csamul_cla32_fa4_21_xor0 = s_csamul_cla32_and4_21 ^ s_csamul_cla32_fa5_20_xor1;
  assign s_csamul_cla32_fa4_21_and0 = s_csamul_cla32_and4_21 & s_csamul_cla32_fa5_20_xor1;
  assign s_csamul_cla32_fa4_21_xor1 = s_csamul_cla32_fa4_21_xor0 ^ s_csamul_cla32_fa4_20_or0;
  assign s_csamul_cla32_fa4_21_and1 = s_csamul_cla32_fa4_21_xor0 & s_csamul_cla32_fa4_20_or0;
  assign s_csamul_cla32_fa4_21_or0 = s_csamul_cla32_fa4_21_and0 | s_csamul_cla32_fa4_21_and1;
  assign s_csamul_cla32_and5_21 = a[5] & b[21];
  assign s_csamul_cla32_fa5_21_xor0 = s_csamul_cla32_and5_21 ^ s_csamul_cla32_fa6_20_xor1;
  assign s_csamul_cla32_fa5_21_and0 = s_csamul_cla32_and5_21 & s_csamul_cla32_fa6_20_xor1;
  assign s_csamul_cla32_fa5_21_xor1 = s_csamul_cla32_fa5_21_xor0 ^ s_csamul_cla32_fa5_20_or0;
  assign s_csamul_cla32_fa5_21_and1 = s_csamul_cla32_fa5_21_xor0 & s_csamul_cla32_fa5_20_or0;
  assign s_csamul_cla32_fa5_21_or0 = s_csamul_cla32_fa5_21_and0 | s_csamul_cla32_fa5_21_and1;
  assign s_csamul_cla32_and6_21 = a[6] & b[21];
  assign s_csamul_cla32_fa6_21_xor0 = s_csamul_cla32_and6_21 ^ s_csamul_cla32_fa7_20_xor1;
  assign s_csamul_cla32_fa6_21_and0 = s_csamul_cla32_and6_21 & s_csamul_cla32_fa7_20_xor1;
  assign s_csamul_cla32_fa6_21_xor1 = s_csamul_cla32_fa6_21_xor0 ^ s_csamul_cla32_fa6_20_or0;
  assign s_csamul_cla32_fa6_21_and1 = s_csamul_cla32_fa6_21_xor0 & s_csamul_cla32_fa6_20_or0;
  assign s_csamul_cla32_fa6_21_or0 = s_csamul_cla32_fa6_21_and0 | s_csamul_cla32_fa6_21_and1;
  assign s_csamul_cla32_and7_21 = a[7] & b[21];
  assign s_csamul_cla32_fa7_21_xor0 = s_csamul_cla32_and7_21 ^ s_csamul_cla32_fa8_20_xor1;
  assign s_csamul_cla32_fa7_21_and0 = s_csamul_cla32_and7_21 & s_csamul_cla32_fa8_20_xor1;
  assign s_csamul_cla32_fa7_21_xor1 = s_csamul_cla32_fa7_21_xor0 ^ s_csamul_cla32_fa7_20_or0;
  assign s_csamul_cla32_fa7_21_and1 = s_csamul_cla32_fa7_21_xor0 & s_csamul_cla32_fa7_20_or0;
  assign s_csamul_cla32_fa7_21_or0 = s_csamul_cla32_fa7_21_and0 | s_csamul_cla32_fa7_21_and1;
  assign s_csamul_cla32_and8_21 = a[8] & b[21];
  assign s_csamul_cla32_fa8_21_xor0 = s_csamul_cla32_and8_21 ^ s_csamul_cla32_fa9_20_xor1;
  assign s_csamul_cla32_fa8_21_and0 = s_csamul_cla32_and8_21 & s_csamul_cla32_fa9_20_xor1;
  assign s_csamul_cla32_fa8_21_xor1 = s_csamul_cla32_fa8_21_xor0 ^ s_csamul_cla32_fa8_20_or0;
  assign s_csamul_cla32_fa8_21_and1 = s_csamul_cla32_fa8_21_xor0 & s_csamul_cla32_fa8_20_or0;
  assign s_csamul_cla32_fa8_21_or0 = s_csamul_cla32_fa8_21_and0 | s_csamul_cla32_fa8_21_and1;
  assign s_csamul_cla32_and9_21 = a[9] & b[21];
  assign s_csamul_cla32_fa9_21_xor0 = s_csamul_cla32_and9_21 ^ s_csamul_cla32_fa10_20_xor1;
  assign s_csamul_cla32_fa9_21_and0 = s_csamul_cla32_and9_21 & s_csamul_cla32_fa10_20_xor1;
  assign s_csamul_cla32_fa9_21_xor1 = s_csamul_cla32_fa9_21_xor0 ^ s_csamul_cla32_fa9_20_or0;
  assign s_csamul_cla32_fa9_21_and1 = s_csamul_cla32_fa9_21_xor0 & s_csamul_cla32_fa9_20_or0;
  assign s_csamul_cla32_fa9_21_or0 = s_csamul_cla32_fa9_21_and0 | s_csamul_cla32_fa9_21_and1;
  assign s_csamul_cla32_and10_21 = a[10] & b[21];
  assign s_csamul_cla32_fa10_21_xor0 = s_csamul_cla32_and10_21 ^ s_csamul_cla32_fa11_20_xor1;
  assign s_csamul_cla32_fa10_21_and0 = s_csamul_cla32_and10_21 & s_csamul_cla32_fa11_20_xor1;
  assign s_csamul_cla32_fa10_21_xor1 = s_csamul_cla32_fa10_21_xor0 ^ s_csamul_cla32_fa10_20_or0;
  assign s_csamul_cla32_fa10_21_and1 = s_csamul_cla32_fa10_21_xor0 & s_csamul_cla32_fa10_20_or0;
  assign s_csamul_cla32_fa10_21_or0 = s_csamul_cla32_fa10_21_and0 | s_csamul_cla32_fa10_21_and1;
  assign s_csamul_cla32_and11_21 = a[11] & b[21];
  assign s_csamul_cla32_fa11_21_xor0 = s_csamul_cla32_and11_21 ^ s_csamul_cla32_fa12_20_xor1;
  assign s_csamul_cla32_fa11_21_and0 = s_csamul_cla32_and11_21 & s_csamul_cla32_fa12_20_xor1;
  assign s_csamul_cla32_fa11_21_xor1 = s_csamul_cla32_fa11_21_xor0 ^ s_csamul_cla32_fa11_20_or0;
  assign s_csamul_cla32_fa11_21_and1 = s_csamul_cla32_fa11_21_xor0 & s_csamul_cla32_fa11_20_or0;
  assign s_csamul_cla32_fa11_21_or0 = s_csamul_cla32_fa11_21_and0 | s_csamul_cla32_fa11_21_and1;
  assign s_csamul_cla32_and12_21 = a[12] & b[21];
  assign s_csamul_cla32_fa12_21_xor0 = s_csamul_cla32_and12_21 ^ s_csamul_cla32_fa13_20_xor1;
  assign s_csamul_cla32_fa12_21_and0 = s_csamul_cla32_and12_21 & s_csamul_cla32_fa13_20_xor1;
  assign s_csamul_cla32_fa12_21_xor1 = s_csamul_cla32_fa12_21_xor0 ^ s_csamul_cla32_fa12_20_or0;
  assign s_csamul_cla32_fa12_21_and1 = s_csamul_cla32_fa12_21_xor0 & s_csamul_cla32_fa12_20_or0;
  assign s_csamul_cla32_fa12_21_or0 = s_csamul_cla32_fa12_21_and0 | s_csamul_cla32_fa12_21_and1;
  assign s_csamul_cla32_and13_21 = a[13] & b[21];
  assign s_csamul_cla32_fa13_21_xor0 = s_csamul_cla32_and13_21 ^ s_csamul_cla32_fa14_20_xor1;
  assign s_csamul_cla32_fa13_21_and0 = s_csamul_cla32_and13_21 & s_csamul_cla32_fa14_20_xor1;
  assign s_csamul_cla32_fa13_21_xor1 = s_csamul_cla32_fa13_21_xor0 ^ s_csamul_cla32_fa13_20_or0;
  assign s_csamul_cla32_fa13_21_and1 = s_csamul_cla32_fa13_21_xor0 & s_csamul_cla32_fa13_20_or0;
  assign s_csamul_cla32_fa13_21_or0 = s_csamul_cla32_fa13_21_and0 | s_csamul_cla32_fa13_21_and1;
  assign s_csamul_cla32_and14_21 = a[14] & b[21];
  assign s_csamul_cla32_fa14_21_xor0 = s_csamul_cla32_and14_21 ^ s_csamul_cla32_fa15_20_xor1;
  assign s_csamul_cla32_fa14_21_and0 = s_csamul_cla32_and14_21 & s_csamul_cla32_fa15_20_xor1;
  assign s_csamul_cla32_fa14_21_xor1 = s_csamul_cla32_fa14_21_xor0 ^ s_csamul_cla32_fa14_20_or0;
  assign s_csamul_cla32_fa14_21_and1 = s_csamul_cla32_fa14_21_xor0 & s_csamul_cla32_fa14_20_or0;
  assign s_csamul_cla32_fa14_21_or0 = s_csamul_cla32_fa14_21_and0 | s_csamul_cla32_fa14_21_and1;
  assign s_csamul_cla32_and15_21 = a[15] & b[21];
  assign s_csamul_cla32_fa15_21_xor0 = s_csamul_cla32_and15_21 ^ s_csamul_cla32_fa16_20_xor1;
  assign s_csamul_cla32_fa15_21_and0 = s_csamul_cla32_and15_21 & s_csamul_cla32_fa16_20_xor1;
  assign s_csamul_cla32_fa15_21_xor1 = s_csamul_cla32_fa15_21_xor0 ^ s_csamul_cla32_fa15_20_or0;
  assign s_csamul_cla32_fa15_21_and1 = s_csamul_cla32_fa15_21_xor0 & s_csamul_cla32_fa15_20_or0;
  assign s_csamul_cla32_fa15_21_or0 = s_csamul_cla32_fa15_21_and0 | s_csamul_cla32_fa15_21_and1;
  assign s_csamul_cla32_and16_21 = a[16] & b[21];
  assign s_csamul_cla32_fa16_21_xor0 = s_csamul_cla32_and16_21 ^ s_csamul_cla32_fa17_20_xor1;
  assign s_csamul_cla32_fa16_21_and0 = s_csamul_cla32_and16_21 & s_csamul_cla32_fa17_20_xor1;
  assign s_csamul_cla32_fa16_21_xor1 = s_csamul_cla32_fa16_21_xor0 ^ s_csamul_cla32_fa16_20_or0;
  assign s_csamul_cla32_fa16_21_and1 = s_csamul_cla32_fa16_21_xor0 & s_csamul_cla32_fa16_20_or0;
  assign s_csamul_cla32_fa16_21_or0 = s_csamul_cla32_fa16_21_and0 | s_csamul_cla32_fa16_21_and1;
  assign s_csamul_cla32_and17_21 = a[17] & b[21];
  assign s_csamul_cla32_fa17_21_xor0 = s_csamul_cla32_and17_21 ^ s_csamul_cla32_fa18_20_xor1;
  assign s_csamul_cla32_fa17_21_and0 = s_csamul_cla32_and17_21 & s_csamul_cla32_fa18_20_xor1;
  assign s_csamul_cla32_fa17_21_xor1 = s_csamul_cla32_fa17_21_xor0 ^ s_csamul_cla32_fa17_20_or0;
  assign s_csamul_cla32_fa17_21_and1 = s_csamul_cla32_fa17_21_xor0 & s_csamul_cla32_fa17_20_or0;
  assign s_csamul_cla32_fa17_21_or0 = s_csamul_cla32_fa17_21_and0 | s_csamul_cla32_fa17_21_and1;
  assign s_csamul_cla32_and18_21 = a[18] & b[21];
  assign s_csamul_cla32_fa18_21_xor0 = s_csamul_cla32_and18_21 ^ s_csamul_cla32_fa19_20_xor1;
  assign s_csamul_cla32_fa18_21_and0 = s_csamul_cla32_and18_21 & s_csamul_cla32_fa19_20_xor1;
  assign s_csamul_cla32_fa18_21_xor1 = s_csamul_cla32_fa18_21_xor0 ^ s_csamul_cla32_fa18_20_or0;
  assign s_csamul_cla32_fa18_21_and1 = s_csamul_cla32_fa18_21_xor0 & s_csamul_cla32_fa18_20_or0;
  assign s_csamul_cla32_fa18_21_or0 = s_csamul_cla32_fa18_21_and0 | s_csamul_cla32_fa18_21_and1;
  assign s_csamul_cla32_and19_21 = a[19] & b[21];
  assign s_csamul_cla32_fa19_21_xor0 = s_csamul_cla32_and19_21 ^ s_csamul_cla32_fa20_20_xor1;
  assign s_csamul_cla32_fa19_21_and0 = s_csamul_cla32_and19_21 & s_csamul_cla32_fa20_20_xor1;
  assign s_csamul_cla32_fa19_21_xor1 = s_csamul_cla32_fa19_21_xor0 ^ s_csamul_cla32_fa19_20_or0;
  assign s_csamul_cla32_fa19_21_and1 = s_csamul_cla32_fa19_21_xor0 & s_csamul_cla32_fa19_20_or0;
  assign s_csamul_cla32_fa19_21_or0 = s_csamul_cla32_fa19_21_and0 | s_csamul_cla32_fa19_21_and1;
  assign s_csamul_cla32_and20_21 = a[20] & b[21];
  assign s_csamul_cla32_fa20_21_xor0 = s_csamul_cla32_and20_21 ^ s_csamul_cla32_fa21_20_xor1;
  assign s_csamul_cla32_fa20_21_and0 = s_csamul_cla32_and20_21 & s_csamul_cla32_fa21_20_xor1;
  assign s_csamul_cla32_fa20_21_xor1 = s_csamul_cla32_fa20_21_xor0 ^ s_csamul_cla32_fa20_20_or0;
  assign s_csamul_cla32_fa20_21_and1 = s_csamul_cla32_fa20_21_xor0 & s_csamul_cla32_fa20_20_or0;
  assign s_csamul_cla32_fa20_21_or0 = s_csamul_cla32_fa20_21_and0 | s_csamul_cla32_fa20_21_and1;
  assign s_csamul_cla32_and21_21 = a[21] & b[21];
  assign s_csamul_cla32_fa21_21_xor0 = s_csamul_cla32_and21_21 ^ s_csamul_cla32_fa22_20_xor1;
  assign s_csamul_cla32_fa21_21_and0 = s_csamul_cla32_and21_21 & s_csamul_cla32_fa22_20_xor1;
  assign s_csamul_cla32_fa21_21_xor1 = s_csamul_cla32_fa21_21_xor0 ^ s_csamul_cla32_fa21_20_or0;
  assign s_csamul_cla32_fa21_21_and1 = s_csamul_cla32_fa21_21_xor0 & s_csamul_cla32_fa21_20_or0;
  assign s_csamul_cla32_fa21_21_or0 = s_csamul_cla32_fa21_21_and0 | s_csamul_cla32_fa21_21_and1;
  assign s_csamul_cla32_and22_21 = a[22] & b[21];
  assign s_csamul_cla32_fa22_21_xor0 = s_csamul_cla32_and22_21 ^ s_csamul_cla32_fa23_20_xor1;
  assign s_csamul_cla32_fa22_21_and0 = s_csamul_cla32_and22_21 & s_csamul_cla32_fa23_20_xor1;
  assign s_csamul_cla32_fa22_21_xor1 = s_csamul_cla32_fa22_21_xor0 ^ s_csamul_cla32_fa22_20_or0;
  assign s_csamul_cla32_fa22_21_and1 = s_csamul_cla32_fa22_21_xor0 & s_csamul_cla32_fa22_20_or0;
  assign s_csamul_cla32_fa22_21_or0 = s_csamul_cla32_fa22_21_and0 | s_csamul_cla32_fa22_21_and1;
  assign s_csamul_cla32_and23_21 = a[23] & b[21];
  assign s_csamul_cla32_fa23_21_xor0 = s_csamul_cla32_and23_21 ^ s_csamul_cla32_fa24_20_xor1;
  assign s_csamul_cla32_fa23_21_and0 = s_csamul_cla32_and23_21 & s_csamul_cla32_fa24_20_xor1;
  assign s_csamul_cla32_fa23_21_xor1 = s_csamul_cla32_fa23_21_xor0 ^ s_csamul_cla32_fa23_20_or0;
  assign s_csamul_cla32_fa23_21_and1 = s_csamul_cla32_fa23_21_xor0 & s_csamul_cla32_fa23_20_or0;
  assign s_csamul_cla32_fa23_21_or0 = s_csamul_cla32_fa23_21_and0 | s_csamul_cla32_fa23_21_and1;
  assign s_csamul_cla32_and24_21 = a[24] & b[21];
  assign s_csamul_cla32_fa24_21_xor0 = s_csamul_cla32_and24_21 ^ s_csamul_cla32_fa25_20_xor1;
  assign s_csamul_cla32_fa24_21_and0 = s_csamul_cla32_and24_21 & s_csamul_cla32_fa25_20_xor1;
  assign s_csamul_cla32_fa24_21_xor1 = s_csamul_cla32_fa24_21_xor0 ^ s_csamul_cla32_fa24_20_or0;
  assign s_csamul_cla32_fa24_21_and1 = s_csamul_cla32_fa24_21_xor0 & s_csamul_cla32_fa24_20_or0;
  assign s_csamul_cla32_fa24_21_or0 = s_csamul_cla32_fa24_21_and0 | s_csamul_cla32_fa24_21_and1;
  assign s_csamul_cla32_and25_21 = a[25] & b[21];
  assign s_csamul_cla32_fa25_21_xor0 = s_csamul_cla32_and25_21 ^ s_csamul_cla32_fa26_20_xor1;
  assign s_csamul_cla32_fa25_21_and0 = s_csamul_cla32_and25_21 & s_csamul_cla32_fa26_20_xor1;
  assign s_csamul_cla32_fa25_21_xor1 = s_csamul_cla32_fa25_21_xor0 ^ s_csamul_cla32_fa25_20_or0;
  assign s_csamul_cla32_fa25_21_and1 = s_csamul_cla32_fa25_21_xor0 & s_csamul_cla32_fa25_20_or0;
  assign s_csamul_cla32_fa25_21_or0 = s_csamul_cla32_fa25_21_and0 | s_csamul_cla32_fa25_21_and1;
  assign s_csamul_cla32_and26_21 = a[26] & b[21];
  assign s_csamul_cla32_fa26_21_xor0 = s_csamul_cla32_and26_21 ^ s_csamul_cla32_fa27_20_xor1;
  assign s_csamul_cla32_fa26_21_and0 = s_csamul_cla32_and26_21 & s_csamul_cla32_fa27_20_xor1;
  assign s_csamul_cla32_fa26_21_xor1 = s_csamul_cla32_fa26_21_xor0 ^ s_csamul_cla32_fa26_20_or0;
  assign s_csamul_cla32_fa26_21_and1 = s_csamul_cla32_fa26_21_xor0 & s_csamul_cla32_fa26_20_or0;
  assign s_csamul_cla32_fa26_21_or0 = s_csamul_cla32_fa26_21_and0 | s_csamul_cla32_fa26_21_and1;
  assign s_csamul_cla32_and27_21 = a[27] & b[21];
  assign s_csamul_cla32_fa27_21_xor0 = s_csamul_cla32_and27_21 ^ s_csamul_cla32_fa28_20_xor1;
  assign s_csamul_cla32_fa27_21_and0 = s_csamul_cla32_and27_21 & s_csamul_cla32_fa28_20_xor1;
  assign s_csamul_cla32_fa27_21_xor1 = s_csamul_cla32_fa27_21_xor0 ^ s_csamul_cla32_fa27_20_or0;
  assign s_csamul_cla32_fa27_21_and1 = s_csamul_cla32_fa27_21_xor0 & s_csamul_cla32_fa27_20_or0;
  assign s_csamul_cla32_fa27_21_or0 = s_csamul_cla32_fa27_21_and0 | s_csamul_cla32_fa27_21_and1;
  assign s_csamul_cla32_and28_21 = a[28] & b[21];
  assign s_csamul_cla32_fa28_21_xor0 = s_csamul_cla32_and28_21 ^ s_csamul_cla32_fa29_20_xor1;
  assign s_csamul_cla32_fa28_21_and0 = s_csamul_cla32_and28_21 & s_csamul_cla32_fa29_20_xor1;
  assign s_csamul_cla32_fa28_21_xor1 = s_csamul_cla32_fa28_21_xor0 ^ s_csamul_cla32_fa28_20_or0;
  assign s_csamul_cla32_fa28_21_and1 = s_csamul_cla32_fa28_21_xor0 & s_csamul_cla32_fa28_20_or0;
  assign s_csamul_cla32_fa28_21_or0 = s_csamul_cla32_fa28_21_and0 | s_csamul_cla32_fa28_21_and1;
  assign s_csamul_cla32_and29_21 = a[29] & b[21];
  assign s_csamul_cla32_fa29_21_xor0 = s_csamul_cla32_and29_21 ^ s_csamul_cla32_fa30_20_xor1;
  assign s_csamul_cla32_fa29_21_and0 = s_csamul_cla32_and29_21 & s_csamul_cla32_fa30_20_xor1;
  assign s_csamul_cla32_fa29_21_xor1 = s_csamul_cla32_fa29_21_xor0 ^ s_csamul_cla32_fa29_20_or0;
  assign s_csamul_cla32_fa29_21_and1 = s_csamul_cla32_fa29_21_xor0 & s_csamul_cla32_fa29_20_or0;
  assign s_csamul_cla32_fa29_21_or0 = s_csamul_cla32_fa29_21_and0 | s_csamul_cla32_fa29_21_and1;
  assign s_csamul_cla32_and30_21 = a[30] & b[21];
  assign s_csamul_cla32_fa30_21_xor0 = s_csamul_cla32_and30_21 ^ s_csamul_cla32_ha31_20_xor0;
  assign s_csamul_cla32_fa30_21_and0 = s_csamul_cla32_and30_21 & s_csamul_cla32_ha31_20_xor0;
  assign s_csamul_cla32_fa30_21_xor1 = s_csamul_cla32_fa30_21_xor0 ^ s_csamul_cla32_fa30_20_or0;
  assign s_csamul_cla32_fa30_21_and1 = s_csamul_cla32_fa30_21_xor0 & s_csamul_cla32_fa30_20_or0;
  assign s_csamul_cla32_fa30_21_or0 = s_csamul_cla32_fa30_21_and0 | s_csamul_cla32_fa30_21_and1;
  assign s_csamul_cla32_nand31_21 = ~(a[31] & b[21]);
  assign s_csamul_cla32_ha31_21_xor0 = s_csamul_cla32_nand31_21 ^ s_csamul_cla32_ha31_20_and0;
  assign s_csamul_cla32_ha31_21_and0 = s_csamul_cla32_nand31_21 & s_csamul_cla32_ha31_20_and0;
  assign s_csamul_cla32_and0_22 = a[0] & b[22];
  assign s_csamul_cla32_fa0_22_xor0 = s_csamul_cla32_and0_22 ^ s_csamul_cla32_fa1_21_xor1;
  assign s_csamul_cla32_fa0_22_and0 = s_csamul_cla32_and0_22 & s_csamul_cla32_fa1_21_xor1;
  assign s_csamul_cla32_fa0_22_xor1 = s_csamul_cla32_fa0_22_xor0 ^ s_csamul_cla32_fa0_21_or0;
  assign s_csamul_cla32_fa0_22_and1 = s_csamul_cla32_fa0_22_xor0 & s_csamul_cla32_fa0_21_or0;
  assign s_csamul_cla32_fa0_22_or0 = s_csamul_cla32_fa0_22_and0 | s_csamul_cla32_fa0_22_and1;
  assign s_csamul_cla32_and1_22 = a[1] & b[22];
  assign s_csamul_cla32_fa1_22_xor0 = s_csamul_cla32_and1_22 ^ s_csamul_cla32_fa2_21_xor1;
  assign s_csamul_cla32_fa1_22_and0 = s_csamul_cla32_and1_22 & s_csamul_cla32_fa2_21_xor1;
  assign s_csamul_cla32_fa1_22_xor1 = s_csamul_cla32_fa1_22_xor0 ^ s_csamul_cla32_fa1_21_or0;
  assign s_csamul_cla32_fa1_22_and1 = s_csamul_cla32_fa1_22_xor0 & s_csamul_cla32_fa1_21_or0;
  assign s_csamul_cla32_fa1_22_or0 = s_csamul_cla32_fa1_22_and0 | s_csamul_cla32_fa1_22_and1;
  assign s_csamul_cla32_and2_22 = a[2] & b[22];
  assign s_csamul_cla32_fa2_22_xor0 = s_csamul_cla32_and2_22 ^ s_csamul_cla32_fa3_21_xor1;
  assign s_csamul_cla32_fa2_22_and0 = s_csamul_cla32_and2_22 & s_csamul_cla32_fa3_21_xor1;
  assign s_csamul_cla32_fa2_22_xor1 = s_csamul_cla32_fa2_22_xor0 ^ s_csamul_cla32_fa2_21_or0;
  assign s_csamul_cla32_fa2_22_and1 = s_csamul_cla32_fa2_22_xor0 & s_csamul_cla32_fa2_21_or0;
  assign s_csamul_cla32_fa2_22_or0 = s_csamul_cla32_fa2_22_and0 | s_csamul_cla32_fa2_22_and1;
  assign s_csamul_cla32_and3_22 = a[3] & b[22];
  assign s_csamul_cla32_fa3_22_xor0 = s_csamul_cla32_and3_22 ^ s_csamul_cla32_fa4_21_xor1;
  assign s_csamul_cla32_fa3_22_and0 = s_csamul_cla32_and3_22 & s_csamul_cla32_fa4_21_xor1;
  assign s_csamul_cla32_fa3_22_xor1 = s_csamul_cla32_fa3_22_xor0 ^ s_csamul_cla32_fa3_21_or0;
  assign s_csamul_cla32_fa3_22_and1 = s_csamul_cla32_fa3_22_xor0 & s_csamul_cla32_fa3_21_or0;
  assign s_csamul_cla32_fa3_22_or0 = s_csamul_cla32_fa3_22_and0 | s_csamul_cla32_fa3_22_and1;
  assign s_csamul_cla32_and4_22 = a[4] & b[22];
  assign s_csamul_cla32_fa4_22_xor0 = s_csamul_cla32_and4_22 ^ s_csamul_cla32_fa5_21_xor1;
  assign s_csamul_cla32_fa4_22_and0 = s_csamul_cla32_and4_22 & s_csamul_cla32_fa5_21_xor1;
  assign s_csamul_cla32_fa4_22_xor1 = s_csamul_cla32_fa4_22_xor0 ^ s_csamul_cla32_fa4_21_or0;
  assign s_csamul_cla32_fa4_22_and1 = s_csamul_cla32_fa4_22_xor0 & s_csamul_cla32_fa4_21_or0;
  assign s_csamul_cla32_fa4_22_or0 = s_csamul_cla32_fa4_22_and0 | s_csamul_cla32_fa4_22_and1;
  assign s_csamul_cla32_and5_22 = a[5] & b[22];
  assign s_csamul_cla32_fa5_22_xor0 = s_csamul_cla32_and5_22 ^ s_csamul_cla32_fa6_21_xor1;
  assign s_csamul_cla32_fa5_22_and0 = s_csamul_cla32_and5_22 & s_csamul_cla32_fa6_21_xor1;
  assign s_csamul_cla32_fa5_22_xor1 = s_csamul_cla32_fa5_22_xor0 ^ s_csamul_cla32_fa5_21_or0;
  assign s_csamul_cla32_fa5_22_and1 = s_csamul_cla32_fa5_22_xor0 & s_csamul_cla32_fa5_21_or0;
  assign s_csamul_cla32_fa5_22_or0 = s_csamul_cla32_fa5_22_and0 | s_csamul_cla32_fa5_22_and1;
  assign s_csamul_cla32_and6_22 = a[6] & b[22];
  assign s_csamul_cla32_fa6_22_xor0 = s_csamul_cla32_and6_22 ^ s_csamul_cla32_fa7_21_xor1;
  assign s_csamul_cla32_fa6_22_and0 = s_csamul_cla32_and6_22 & s_csamul_cla32_fa7_21_xor1;
  assign s_csamul_cla32_fa6_22_xor1 = s_csamul_cla32_fa6_22_xor0 ^ s_csamul_cla32_fa6_21_or0;
  assign s_csamul_cla32_fa6_22_and1 = s_csamul_cla32_fa6_22_xor0 & s_csamul_cla32_fa6_21_or0;
  assign s_csamul_cla32_fa6_22_or0 = s_csamul_cla32_fa6_22_and0 | s_csamul_cla32_fa6_22_and1;
  assign s_csamul_cla32_and7_22 = a[7] & b[22];
  assign s_csamul_cla32_fa7_22_xor0 = s_csamul_cla32_and7_22 ^ s_csamul_cla32_fa8_21_xor1;
  assign s_csamul_cla32_fa7_22_and0 = s_csamul_cla32_and7_22 & s_csamul_cla32_fa8_21_xor1;
  assign s_csamul_cla32_fa7_22_xor1 = s_csamul_cla32_fa7_22_xor0 ^ s_csamul_cla32_fa7_21_or0;
  assign s_csamul_cla32_fa7_22_and1 = s_csamul_cla32_fa7_22_xor0 & s_csamul_cla32_fa7_21_or0;
  assign s_csamul_cla32_fa7_22_or0 = s_csamul_cla32_fa7_22_and0 | s_csamul_cla32_fa7_22_and1;
  assign s_csamul_cla32_and8_22 = a[8] & b[22];
  assign s_csamul_cla32_fa8_22_xor0 = s_csamul_cla32_and8_22 ^ s_csamul_cla32_fa9_21_xor1;
  assign s_csamul_cla32_fa8_22_and0 = s_csamul_cla32_and8_22 & s_csamul_cla32_fa9_21_xor1;
  assign s_csamul_cla32_fa8_22_xor1 = s_csamul_cla32_fa8_22_xor0 ^ s_csamul_cla32_fa8_21_or0;
  assign s_csamul_cla32_fa8_22_and1 = s_csamul_cla32_fa8_22_xor0 & s_csamul_cla32_fa8_21_or0;
  assign s_csamul_cla32_fa8_22_or0 = s_csamul_cla32_fa8_22_and0 | s_csamul_cla32_fa8_22_and1;
  assign s_csamul_cla32_and9_22 = a[9] & b[22];
  assign s_csamul_cla32_fa9_22_xor0 = s_csamul_cla32_and9_22 ^ s_csamul_cla32_fa10_21_xor1;
  assign s_csamul_cla32_fa9_22_and0 = s_csamul_cla32_and9_22 & s_csamul_cla32_fa10_21_xor1;
  assign s_csamul_cla32_fa9_22_xor1 = s_csamul_cla32_fa9_22_xor0 ^ s_csamul_cla32_fa9_21_or0;
  assign s_csamul_cla32_fa9_22_and1 = s_csamul_cla32_fa9_22_xor0 & s_csamul_cla32_fa9_21_or0;
  assign s_csamul_cla32_fa9_22_or0 = s_csamul_cla32_fa9_22_and0 | s_csamul_cla32_fa9_22_and1;
  assign s_csamul_cla32_and10_22 = a[10] & b[22];
  assign s_csamul_cla32_fa10_22_xor0 = s_csamul_cla32_and10_22 ^ s_csamul_cla32_fa11_21_xor1;
  assign s_csamul_cla32_fa10_22_and0 = s_csamul_cla32_and10_22 & s_csamul_cla32_fa11_21_xor1;
  assign s_csamul_cla32_fa10_22_xor1 = s_csamul_cla32_fa10_22_xor0 ^ s_csamul_cla32_fa10_21_or0;
  assign s_csamul_cla32_fa10_22_and1 = s_csamul_cla32_fa10_22_xor0 & s_csamul_cla32_fa10_21_or0;
  assign s_csamul_cla32_fa10_22_or0 = s_csamul_cla32_fa10_22_and0 | s_csamul_cla32_fa10_22_and1;
  assign s_csamul_cla32_and11_22 = a[11] & b[22];
  assign s_csamul_cla32_fa11_22_xor0 = s_csamul_cla32_and11_22 ^ s_csamul_cla32_fa12_21_xor1;
  assign s_csamul_cla32_fa11_22_and0 = s_csamul_cla32_and11_22 & s_csamul_cla32_fa12_21_xor1;
  assign s_csamul_cla32_fa11_22_xor1 = s_csamul_cla32_fa11_22_xor0 ^ s_csamul_cla32_fa11_21_or0;
  assign s_csamul_cla32_fa11_22_and1 = s_csamul_cla32_fa11_22_xor0 & s_csamul_cla32_fa11_21_or0;
  assign s_csamul_cla32_fa11_22_or0 = s_csamul_cla32_fa11_22_and0 | s_csamul_cla32_fa11_22_and1;
  assign s_csamul_cla32_and12_22 = a[12] & b[22];
  assign s_csamul_cla32_fa12_22_xor0 = s_csamul_cla32_and12_22 ^ s_csamul_cla32_fa13_21_xor1;
  assign s_csamul_cla32_fa12_22_and0 = s_csamul_cla32_and12_22 & s_csamul_cla32_fa13_21_xor1;
  assign s_csamul_cla32_fa12_22_xor1 = s_csamul_cla32_fa12_22_xor0 ^ s_csamul_cla32_fa12_21_or0;
  assign s_csamul_cla32_fa12_22_and1 = s_csamul_cla32_fa12_22_xor0 & s_csamul_cla32_fa12_21_or0;
  assign s_csamul_cla32_fa12_22_or0 = s_csamul_cla32_fa12_22_and0 | s_csamul_cla32_fa12_22_and1;
  assign s_csamul_cla32_and13_22 = a[13] & b[22];
  assign s_csamul_cla32_fa13_22_xor0 = s_csamul_cla32_and13_22 ^ s_csamul_cla32_fa14_21_xor1;
  assign s_csamul_cla32_fa13_22_and0 = s_csamul_cla32_and13_22 & s_csamul_cla32_fa14_21_xor1;
  assign s_csamul_cla32_fa13_22_xor1 = s_csamul_cla32_fa13_22_xor0 ^ s_csamul_cla32_fa13_21_or0;
  assign s_csamul_cla32_fa13_22_and1 = s_csamul_cla32_fa13_22_xor0 & s_csamul_cla32_fa13_21_or0;
  assign s_csamul_cla32_fa13_22_or0 = s_csamul_cla32_fa13_22_and0 | s_csamul_cla32_fa13_22_and1;
  assign s_csamul_cla32_and14_22 = a[14] & b[22];
  assign s_csamul_cla32_fa14_22_xor0 = s_csamul_cla32_and14_22 ^ s_csamul_cla32_fa15_21_xor1;
  assign s_csamul_cla32_fa14_22_and0 = s_csamul_cla32_and14_22 & s_csamul_cla32_fa15_21_xor1;
  assign s_csamul_cla32_fa14_22_xor1 = s_csamul_cla32_fa14_22_xor0 ^ s_csamul_cla32_fa14_21_or0;
  assign s_csamul_cla32_fa14_22_and1 = s_csamul_cla32_fa14_22_xor0 & s_csamul_cla32_fa14_21_or0;
  assign s_csamul_cla32_fa14_22_or0 = s_csamul_cla32_fa14_22_and0 | s_csamul_cla32_fa14_22_and1;
  assign s_csamul_cla32_and15_22 = a[15] & b[22];
  assign s_csamul_cla32_fa15_22_xor0 = s_csamul_cla32_and15_22 ^ s_csamul_cla32_fa16_21_xor1;
  assign s_csamul_cla32_fa15_22_and0 = s_csamul_cla32_and15_22 & s_csamul_cla32_fa16_21_xor1;
  assign s_csamul_cla32_fa15_22_xor1 = s_csamul_cla32_fa15_22_xor0 ^ s_csamul_cla32_fa15_21_or0;
  assign s_csamul_cla32_fa15_22_and1 = s_csamul_cla32_fa15_22_xor0 & s_csamul_cla32_fa15_21_or0;
  assign s_csamul_cla32_fa15_22_or0 = s_csamul_cla32_fa15_22_and0 | s_csamul_cla32_fa15_22_and1;
  assign s_csamul_cla32_and16_22 = a[16] & b[22];
  assign s_csamul_cla32_fa16_22_xor0 = s_csamul_cla32_and16_22 ^ s_csamul_cla32_fa17_21_xor1;
  assign s_csamul_cla32_fa16_22_and0 = s_csamul_cla32_and16_22 & s_csamul_cla32_fa17_21_xor1;
  assign s_csamul_cla32_fa16_22_xor1 = s_csamul_cla32_fa16_22_xor0 ^ s_csamul_cla32_fa16_21_or0;
  assign s_csamul_cla32_fa16_22_and1 = s_csamul_cla32_fa16_22_xor0 & s_csamul_cla32_fa16_21_or0;
  assign s_csamul_cla32_fa16_22_or0 = s_csamul_cla32_fa16_22_and0 | s_csamul_cla32_fa16_22_and1;
  assign s_csamul_cla32_and17_22 = a[17] & b[22];
  assign s_csamul_cla32_fa17_22_xor0 = s_csamul_cla32_and17_22 ^ s_csamul_cla32_fa18_21_xor1;
  assign s_csamul_cla32_fa17_22_and0 = s_csamul_cla32_and17_22 & s_csamul_cla32_fa18_21_xor1;
  assign s_csamul_cla32_fa17_22_xor1 = s_csamul_cla32_fa17_22_xor0 ^ s_csamul_cla32_fa17_21_or0;
  assign s_csamul_cla32_fa17_22_and1 = s_csamul_cla32_fa17_22_xor0 & s_csamul_cla32_fa17_21_or0;
  assign s_csamul_cla32_fa17_22_or0 = s_csamul_cla32_fa17_22_and0 | s_csamul_cla32_fa17_22_and1;
  assign s_csamul_cla32_and18_22 = a[18] & b[22];
  assign s_csamul_cla32_fa18_22_xor0 = s_csamul_cla32_and18_22 ^ s_csamul_cla32_fa19_21_xor1;
  assign s_csamul_cla32_fa18_22_and0 = s_csamul_cla32_and18_22 & s_csamul_cla32_fa19_21_xor1;
  assign s_csamul_cla32_fa18_22_xor1 = s_csamul_cla32_fa18_22_xor0 ^ s_csamul_cla32_fa18_21_or0;
  assign s_csamul_cla32_fa18_22_and1 = s_csamul_cla32_fa18_22_xor0 & s_csamul_cla32_fa18_21_or0;
  assign s_csamul_cla32_fa18_22_or0 = s_csamul_cla32_fa18_22_and0 | s_csamul_cla32_fa18_22_and1;
  assign s_csamul_cla32_and19_22 = a[19] & b[22];
  assign s_csamul_cla32_fa19_22_xor0 = s_csamul_cla32_and19_22 ^ s_csamul_cla32_fa20_21_xor1;
  assign s_csamul_cla32_fa19_22_and0 = s_csamul_cla32_and19_22 & s_csamul_cla32_fa20_21_xor1;
  assign s_csamul_cla32_fa19_22_xor1 = s_csamul_cla32_fa19_22_xor0 ^ s_csamul_cla32_fa19_21_or0;
  assign s_csamul_cla32_fa19_22_and1 = s_csamul_cla32_fa19_22_xor0 & s_csamul_cla32_fa19_21_or0;
  assign s_csamul_cla32_fa19_22_or0 = s_csamul_cla32_fa19_22_and0 | s_csamul_cla32_fa19_22_and1;
  assign s_csamul_cla32_and20_22 = a[20] & b[22];
  assign s_csamul_cla32_fa20_22_xor0 = s_csamul_cla32_and20_22 ^ s_csamul_cla32_fa21_21_xor1;
  assign s_csamul_cla32_fa20_22_and0 = s_csamul_cla32_and20_22 & s_csamul_cla32_fa21_21_xor1;
  assign s_csamul_cla32_fa20_22_xor1 = s_csamul_cla32_fa20_22_xor0 ^ s_csamul_cla32_fa20_21_or0;
  assign s_csamul_cla32_fa20_22_and1 = s_csamul_cla32_fa20_22_xor0 & s_csamul_cla32_fa20_21_or0;
  assign s_csamul_cla32_fa20_22_or0 = s_csamul_cla32_fa20_22_and0 | s_csamul_cla32_fa20_22_and1;
  assign s_csamul_cla32_and21_22 = a[21] & b[22];
  assign s_csamul_cla32_fa21_22_xor0 = s_csamul_cla32_and21_22 ^ s_csamul_cla32_fa22_21_xor1;
  assign s_csamul_cla32_fa21_22_and0 = s_csamul_cla32_and21_22 & s_csamul_cla32_fa22_21_xor1;
  assign s_csamul_cla32_fa21_22_xor1 = s_csamul_cla32_fa21_22_xor0 ^ s_csamul_cla32_fa21_21_or0;
  assign s_csamul_cla32_fa21_22_and1 = s_csamul_cla32_fa21_22_xor0 & s_csamul_cla32_fa21_21_or0;
  assign s_csamul_cla32_fa21_22_or0 = s_csamul_cla32_fa21_22_and0 | s_csamul_cla32_fa21_22_and1;
  assign s_csamul_cla32_and22_22 = a[22] & b[22];
  assign s_csamul_cla32_fa22_22_xor0 = s_csamul_cla32_and22_22 ^ s_csamul_cla32_fa23_21_xor1;
  assign s_csamul_cla32_fa22_22_and0 = s_csamul_cla32_and22_22 & s_csamul_cla32_fa23_21_xor1;
  assign s_csamul_cla32_fa22_22_xor1 = s_csamul_cla32_fa22_22_xor0 ^ s_csamul_cla32_fa22_21_or0;
  assign s_csamul_cla32_fa22_22_and1 = s_csamul_cla32_fa22_22_xor0 & s_csamul_cla32_fa22_21_or0;
  assign s_csamul_cla32_fa22_22_or0 = s_csamul_cla32_fa22_22_and0 | s_csamul_cla32_fa22_22_and1;
  assign s_csamul_cla32_and23_22 = a[23] & b[22];
  assign s_csamul_cla32_fa23_22_xor0 = s_csamul_cla32_and23_22 ^ s_csamul_cla32_fa24_21_xor1;
  assign s_csamul_cla32_fa23_22_and0 = s_csamul_cla32_and23_22 & s_csamul_cla32_fa24_21_xor1;
  assign s_csamul_cla32_fa23_22_xor1 = s_csamul_cla32_fa23_22_xor0 ^ s_csamul_cla32_fa23_21_or0;
  assign s_csamul_cla32_fa23_22_and1 = s_csamul_cla32_fa23_22_xor0 & s_csamul_cla32_fa23_21_or0;
  assign s_csamul_cla32_fa23_22_or0 = s_csamul_cla32_fa23_22_and0 | s_csamul_cla32_fa23_22_and1;
  assign s_csamul_cla32_and24_22 = a[24] & b[22];
  assign s_csamul_cla32_fa24_22_xor0 = s_csamul_cla32_and24_22 ^ s_csamul_cla32_fa25_21_xor1;
  assign s_csamul_cla32_fa24_22_and0 = s_csamul_cla32_and24_22 & s_csamul_cla32_fa25_21_xor1;
  assign s_csamul_cla32_fa24_22_xor1 = s_csamul_cla32_fa24_22_xor0 ^ s_csamul_cla32_fa24_21_or0;
  assign s_csamul_cla32_fa24_22_and1 = s_csamul_cla32_fa24_22_xor0 & s_csamul_cla32_fa24_21_or0;
  assign s_csamul_cla32_fa24_22_or0 = s_csamul_cla32_fa24_22_and0 | s_csamul_cla32_fa24_22_and1;
  assign s_csamul_cla32_and25_22 = a[25] & b[22];
  assign s_csamul_cla32_fa25_22_xor0 = s_csamul_cla32_and25_22 ^ s_csamul_cla32_fa26_21_xor1;
  assign s_csamul_cla32_fa25_22_and0 = s_csamul_cla32_and25_22 & s_csamul_cla32_fa26_21_xor1;
  assign s_csamul_cla32_fa25_22_xor1 = s_csamul_cla32_fa25_22_xor0 ^ s_csamul_cla32_fa25_21_or0;
  assign s_csamul_cla32_fa25_22_and1 = s_csamul_cla32_fa25_22_xor0 & s_csamul_cla32_fa25_21_or0;
  assign s_csamul_cla32_fa25_22_or0 = s_csamul_cla32_fa25_22_and0 | s_csamul_cla32_fa25_22_and1;
  assign s_csamul_cla32_and26_22 = a[26] & b[22];
  assign s_csamul_cla32_fa26_22_xor0 = s_csamul_cla32_and26_22 ^ s_csamul_cla32_fa27_21_xor1;
  assign s_csamul_cla32_fa26_22_and0 = s_csamul_cla32_and26_22 & s_csamul_cla32_fa27_21_xor1;
  assign s_csamul_cla32_fa26_22_xor1 = s_csamul_cla32_fa26_22_xor0 ^ s_csamul_cla32_fa26_21_or0;
  assign s_csamul_cla32_fa26_22_and1 = s_csamul_cla32_fa26_22_xor0 & s_csamul_cla32_fa26_21_or0;
  assign s_csamul_cla32_fa26_22_or0 = s_csamul_cla32_fa26_22_and0 | s_csamul_cla32_fa26_22_and1;
  assign s_csamul_cla32_and27_22 = a[27] & b[22];
  assign s_csamul_cla32_fa27_22_xor0 = s_csamul_cla32_and27_22 ^ s_csamul_cla32_fa28_21_xor1;
  assign s_csamul_cla32_fa27_22_and0 = s_csamul_cla32_and27_22 & s_csamul_cla32_fa28_21_xor1;
  assign s_csamul_cla32_fa27_22_xor1 = s_csamul_cla32_fa27_22_xor0 ^ s_csamul_cla32_fa27_21_or0;
  assign s_csamul_cla32_fa27_22_and1 = s_csamul_cla32_fa27_22_xor0 & s_csamul_cla32_fa27_21_or0;
  assign s_csamul_cla32_fa27_22_or0 = s_csamul_cla32_fa27_22_and0 | s_csamul_cla32_fa27_22_and1;
  assign s_csamul_cla32_and28_22 = a[28] & b[22];
  assign s_csamul_cla32_fa28_22_xor0 = s_csamul_cla32_and28_22 ^ s_csamul_cla32_fa29_21_xor1;
  assign s_csamul_cla32_fa28_22_and0 = s_csamul_cla32_and28_22 & s_csamul_cla32_fa29_21_xor1;
  assign s_csamul_cla32_fa28_22_xor1 = s_csamul_cla32_fa28_22_xor0 ^ s_csamul_cla32_fa28_21_or0;
  assign s_csamul_cla32_fa28_22_and1 = s_csamul_cla32_fa28_22_xor0 & s_csamul_cla32_fa28_21_or0;
  assign s_csamul_cla32_fa28_22_or0 = s_csamul_cla32_fa28_22_and0 | s_csamul_cla32_fa28_22_and1;
  assign s_csamul_cla32_and29_22 = a[29] & b[22];
  assign s_csamul_cla32_fa29_22_xor0 = s_csamul_cla32_and29_22 ^ s_csamul_cla32_fa30_21_xor1;
  assign s_csamul_cla32_fa29_22_and0 = s_csamul_cla32_and29_22 & s_csamul_cla32_fa30_21_xor1;
  assign s_csamul_cla32_fa29_22_xor1 = s_csamul_cla32_fa29_22_xor0 ^ s_csamul_cla32_fa29_21_or0;
  assign s_csamul_cla32_fa29_22_and1 = s_csamul_cla32_fa29_22_xor0 & s_csamul_cla32_fa29_21_or0;
  assign s_csamul_cla32_fa29_22_or0 = s_csamul_cla32_fa29_22_and0 | s_csamul_cla32_fa29_22_and1;
  assign s_csamul_cla32_and30_22 = a[30] & b[22];
  assign s_csamul_cla32_fa30_22_xor0 = s_csamul_cla32_and30_22 ^ s_csamul_cla32_ha31_21_xor0;
  assign s_csamul_cla32_fa30_22_and0 = s_csamul_cla32_and30_22 & s_csamul_cla32_ha31_21_xor0;
  assign s_csamul_cla32_fa30_22_xor1 = s_csamul_cla32_fa30_22_xor0 ^ s_csamul_cla32_fa30_21_or0;
  assign s_csamul_cla32_fa30_22_and1 = s_csamul_cla32_fa30_22_xor0 & s_csamul_cla32_fa30_21_or0;
  assign s_csamul_cla32_fa30_22_or0 = s_csamul_cla32_fa30_22_and0 | s_csamul_cla32_fa30_22_and1;
  assign s_csamul_cla32_nand31_22 = ~(a[31] & b[22]);
  assign s_csamul_cla32_ha31_22_xor0 = s_csamul_cla32_nand31_22 ^ s_csamul_cla32_ha31_21_and0;
  assign s_csamul_cla32_ha31_22_and0 = s_csamul_cla32_nand31_22 & s_csamul_cla32_ha31_21_and0;
  assign s_csamul_cla32_and0_23 = a[0] & b[23];
  assign s_csamul_cla32_fa0_23_xor0 = s_csamul_cla32_and0_23 ^ s_csamul_cla32_fa1_22_xor1;
  assign s_csamul_cla32_fa0_23_and0 = s_csamul_cla32_and0_23 & s_csamul_cla32_fa1_22_xor1;
  assign s_csamul_cla32_fa0_23_xor1 = s_csamul_cla32_fa0_23_xor0 ^ s_csamul_cla32_fa0_22_or0;
  assign s_csamul_cla32_fa0_23_and1 = s_csamul_cla32_fa0_23_xor0 & s_csamul_cla32_fa0_22_or0;
  assign s_csamul_cla32_fa0_23_or0 = s_csamul_cla32_fa0_23_and0 | s_csamul_cla32_fa0_23_and1;
  assign s_csamul_cla32_and1_23 = a[1] & b[23];
  assign s_csamul_cla32_fa1_23_xor0 = s_csamul_cla32_and1_23 ^ s_csamul_cla32_fa2_22_xor1;
  assign s_csamul_cla32_fa1_23_and0 = s_csamul_cla32_and1_23 & s_csamul_cla32_fa2_22_xor1;
  assign s_csamul_cla32_fa1_23_xor1 = s_csamul_cla32_fa1_23_xor0 ^ s_csamul_cla32_fa1_22_or0;
  assign s_csamul_cla32_fa1_23_and1 = s_csamul_cla32_fa1_23_xor0 & s_csamul_cla32_fa1_22_or0;
  assign s_csamul_cla32_fa1_23_or0 = s_csamul_cla32_fa1_23_and0 | s_csamul_cla32_fa1_23_and1;
  assign s_csamul_cla32_and2_23 = a[2] & b[23];
  assign s_csamul_cla32_fa2_23_xor0 = s_csamul_cla32_and2_23 ^ s_csamul_cla32_fa3_22_xor1;
  assign s_csamul_cla32_fa2_23_and0 = s_csamul_cla32_and2_23 & s_csamul_cla32_fa3_22_xor1;
  assign s_csamul_cla32_fa2_23_xor1 = s_csamul_cla32_fa2_23_xor0 ^ s_csamul_cla32_fa2_22_or0;
  assign s_csamul_cla32_fa2_23_and1 = s_csamul_cla32_fa2_23_xor0 & s_csamul_cla32_fa2_22_or0;
  assign s_csamul_cla32_fa2_23_or0 = s_csamul_cla32_fa2_23_and0 | s_csamul_cla32_fa2_23_and1;
  assign s_csamul_cla32_and3_23 = a[3] & b[23];
  assign s_csamul_cla32_fa3_23_xor0 = s_csamul_cla32_and3_23 ^ s_csamul_cla32_fa4_22_xor1;
  assign s_csamul_cla32_fa3_23_and0 = s_csamul_cla32_and3_23 & s_csamul_cla32_fa4_22_xor1;
  assign s_csamul_cla32_fa3_23_xor1 = s_csamul_cla32_fa3_23_xor0 ^ s_csamul_cla32_fa3_22_or0;
  assign s_csamul_cla32_fa3_23_and1 = s_csamul_cla32_fa3_23_xor0 & s_csamul_cla32_fa3_22_or0;
  assign s_csamul_cla32_fa3_23_or0 = s_csamul_cla32_fa3_23_and0 | s_csamul_cla32_fa3_23_and1;
  assign s_csamul_cla32_and4_23 = a[4] & b[23];
  assign s_csamul_cla32_fa4_23_xor0 = s_csamul_cla32_and4_23 ^ s_csamul_cla32_fa5_22_xor1;
  assign s_csamul_cla32_fa4_23_and0 = s_csamul_cla32_and4_23 & s_csamul_cla32_fa5_22_xor1;
  assign s_csamul_cla32_fa4_23_xor1 = s_csamul_cla32_fa4_23_xor0 ^ s_csamul_cla32_fa4_22_or0;
  assign s_csamul_cla32_fa4_23_and1 = s_csamul_cla32_fa4_23_xor0 & s_csamul_cla32_fa4_22_or0;
  assign s_csamul_cla32_fa4_23_or0 = s_csamul_cla32_fa4_23_and0 | s_csamul_cla32_fa4_23_and1;
  assign s_csamul_cla32_and5_23 = a[5] & b[23];
  assign s_csamul_cla32_fa5_23_xor0 = s_csamul_cla32_and5_23 ^ s_csamul_cla32_fa6_22_xor1;
  assign s_csamul_cla32_fa5_23_and0 = s_csamul_cla32_and5_23 & s_csamul_cla32_fa6_22_xor1;
  assign s_csamul_cla32_fa5_23_xor1 = s_csamul_cla32_fa5_23_xor0 ^ s_csamul_cla32_fa5_22_or0;
  assign s_csamul_cla32_fa5_23_and1 = s_csamul_cla32_fa5_23_xor0 & s_csamul_cla32_fa5_22_or0;
  assign s_csamul_cla32_fa5_23_or0 = s_csamul_cla32_fa5_23_and0 | s_csamul_cla32_fa5_23_and1;
  assign s_csamul_cla32_and6_23 = a[6] & b[23];
  assign s_csamul_cla32_fa6_23_xor0 = s_csamul_cla32_and6_23 ^ s_csamul_cla32_fa7_22_xor1;
  assign s_csamul_cla32_fa6_23_and0 = s_csamul_cla32_and6_23 & s_csamul_cla32_fa7_22_xor1;
  assign s_csamul_cla32_fa6_23_xor1 = s_csamul_cla32_fa6_23_xor0 ^ s_csamul_cla32_fa6_22_or0;
  assign s_csamul_cla32_fa6_23_and1 = s_csamul_cla32_fa6_23_xor0 & s_csamul_cla32_fa6_22_or0;
  assign s_csamul_cla32_fa6_23_or0 = s_csamul_cla32_fa6_23_and0 | s_csamul_cla32_fa6_23_and1;
  assign s_csamul_cla32_and7_23 = a[7] & b[23];
  assign s_csamul_cla32_fa7_23_xor0 = s_csamul_cla32_and7_23 ^ s_csamul_cla32_fa8_22_xor1;
  assign s_csamul_cla32_fa7_23_and0 = s_csamul_cla32_and7_23 & s_csamul_cla32_fa8_22_xor1;
  assign s_csamul_cla32_fa7_23_xor1 = s_csamul_cla32_fa7_23_xor0 ^ s_csamul_cla32_fa7_22_or0;
  assign s_csamul_cla32_fa7_23_and1 = s_csamul_cla32_fa7_23_xor0 & s_csamul_cla32_fa7_22_or0;
  assign s_csamul_cla32_fa7_23_or0 = s_csamul_cla32_fa7_23_and0 | s_csamul_cla32_fa7_23_and1;
  assign s_csamul_cla32_and8_23 = a[8] & b[23];
  assign s_csamul_cla32_fa8_23_xor0 = s_csamul_cla32_and8_23 ^ s_csamul_cla32_fa9_22_xor1;
  assign s_csamul_cla32_fa8_23_and0 = s_csamul_cla32_and8_23 & s_csamul_cla32_fa9_22_xor1;
  assign s_csamul_cla32_fa8_23_xor1 = s_csamul_cla32_fa8_23_xor0 ^ s_csamul_cla32_fa8_22_or0;
  assign s_csamul_cla32_fa8_23_and1 = s_csamul_cla32_fa8_23_xor0 & s_csamul_cla32_fa8_22_or0;
  assign s_csamul_cla32_fa8_23_or0 = s_csamul_cla32_fa8_23_and0 | s_csamul_cla32_fa8_23_and1;
  assign s_csamul_cla32_and9_23 = a[9] & b[23];
  assign s_csamul_cla32_fa9_23_xor0 = s_csamul_cla32_and9_23 ^ s_csamul_cla32_fa10_22_xor1;
  assign s_csamul_cla32_fa9_23_and0 = s_csamul_cla32_and9_23 & s_csamul_cla32_fa10_22_xor1;
  assign s_csamul_cla32_fa9_23_xor1 = s_csamul_cla32_fa9_23_xor0 ^ s_csamul_cla32_fa9_22_or0;
  assign s_csamul_cla32_fa9_23_and1 = s_csamul_cla32_fa9_23_xor0 & s_csamul_cla32_fa9_22_or0;
  assign s_csamul_cla32_fa9_23_or0 = s_csamul_cla32_fa9_23_and0 | s_csamul_cla32_fa9_23_and1;
  assign s_csamul_cla32_and10_23 = a[10] & b[23];
  assign s_csamul_cla32_fa10_23_xor0 = s_csamul_cla32_and10_23 ^ s_csamul_cla32_fa11_22_xor1;
  assign s_csamul_cla32_fa10_23_and0 = s_csamul_cla32_and10_23 & s_csamul_cla32_fa11_22_xor1;
  assign s_csamul_cla32_fa10_23_xor1 = s_csamul_cla32_fa10_23_xor0 ^ s_csamul_cla32_fa10_22_or0;
  assign s_csamul_cla32_fa10_23_and1 = s_csamul_cla32_fa10_23_xor0 & s_csamul_cla32_fa10_22_or0;
  assign s_csamul_cla32_fa10_23_or0 = s_csamul_cla32_fa10_23_and0 | s_csamul_cla32_fa10_23_and1;
  assign s_csamul_cla32_and11_23 = a[11] & b[23];
  assign s_csamul_cla32_fa11_23_xor0 = s_csamul_cla32_and11_23 ^ s_csamul_cla32_fa12_22_xor1;
  assign s_csamul_cla32_fa11_23_and0 = s_csamul_cla32_and11_23 & s_csamul_cla32_fa12_22_xor1;
  assign s_csamul_cla32_fa11_23_xor1 = s_csamul_cla32_fa11_23_xor0 ^ s_csamul_cla32_fa11_22_or0;
  assign s_csamul_cla32_fa11_23_and1 = s_csamul_cla32_fa11_23_xor0 & s_csamul_cla32_fa11_22_or0;
  assign s_csamul_cla32_fa11_23_or0 = s_csamul_cla32_fa11_23_and0 | s_csamul_cla32_fa11_23_and1;
  assign s_csamul_cla32_and12_23 = a[12] & b[23];
  assign s_csamul_cla32_fa12_23_xor0 = s_csamul_cla32_and12_23 ^ s_csamul_cla32_fa13_22_xor1;
  assign s_csamul_cla32_fa12_23_and0 = s_csamul_cla32_and12_23 & s_csamul_cla32_fa13_22_xor1;
  assign s_csamul_cla32_fa12_23_xor1 = s_csamul_cla32_fa12_23_xor0 ^ s_csamul_cla32_fa12_22_or0;
  assign s_csamul_cla32_fa12_23_and1 = s_csamul_cla32_fa12_23_xor0 & s_csamul_cla32_fa12_22_or0;
  assign s_csamul_cla32_fa12_23_or0 = s_csamul_cla32_fa12_23_and0 | s_csamul_cla32_fa12_23_and1;
  assign s_csamul_cla32_and13_23 = a[13] & b[23];
  assign s_csamul_cla32_fa13_23_xor0 = s_csamul_cla32_and13_23 ^ s_csamul_cla32_fa14_22_xor1;
  assign s_csamul_cla32_fa13_23_and0 = s_csamul_cla32_and13_23 & s_csamul_cla32_fa14_22_xor1;
  assign s_csamul_cla32_fa13_23_xor1 = s_csamul_cla32_fa13_23_xor0 ^ s_csamul_cla32_fa13_22_or0;
  assign s_csamul_cla32_fa13_23_and1 = s_csamul_cla32_fa13_23_xor0 & s_csamul_cla32_fa13_22_or0;
  assign s_csamul_cla32_fa13_23_or0 = s_csamul_cla32_fa13_23_and0 | s_csamul_cla32_fa13_23_and1;
  assign s_csamul_cla32_and14_23 = a[14] & b[23];
  assign s_csamul_cla32_fa14_23_xor0 = s_csamul_cla32_and14_23 ^ s_csamul_cla32_fa15_22_xor1;
  assign s_csamul_cla32_fa14_23_and0 = s_csamul_cla32_and14_23 & s_csamul_cla32_fa15_22_xor1;
  assign s_csamul_cla32_fa14_23_xor1 = s_csamul_cla32_fa14_23_xor0 ^ s_csamul_cla32_fa14_22_or0;
  assign s_csamul_cla32_fa14_23_and1 = s_csamul_cla32_fa14_23_xor0 & s_csamul_cla32_fa14_22_or0;
  assign s_csamul_cla32_fa14_23_or0 = s_csamul_cla32_fa14_23_and0 | s_csamul_cla32_fa14_23_and1;
  assign s_csamul_cla32_and15_23 = a[15] & b[23];
  assign s_csamul_cla32_fa15_23_xor0 = s_csamul_cla32_and15_23 ^ s_csamul_cla32_fa16_22_xor1;
  assign s_csamul_cla32_fa15_23_and0 = s_csamul_cla32_and15_23 & s_csamul_cla32_fa16_22_xor1;
  assign s_csamul_cla32_fa15_23_xor1 = s_csamul_cla32_fa15_23_xor0 ^ s_csamul_cla32_fa15_22_or0;
  assign s_csamul_cla32_fa15_23_and1 = s_csamul_cla32_fa15_23_xor0 & s_csamul_cla32_fa15_22_or0;
  assign s_csamul_cla32_fa15_23_or0 = s_csamul_cla32_fa15_23_and0 | s_csamul_cla32_fa15_23_and1;
  assign s_csamul_cla32_and16_23 = a[16] & b[23];
  assign s_csamul_cla32_fa16_23_xor0 = s_csamul_cla32_and16_23 ^ s_csamul_cla32_fa17_22_xor1;
  assign s_csamul_cla32_fa16_23_and0 = s_csamul_cla32_and16_23 & s_csamul_cla32_fa17_22_xor1;
  assign s_csamul_cla32_fa16_23_xor1 = s_csamul_cla32_fa16_23_xor0 ^ s_csamul_cla32_fa16_22_or0;
  assign s_csamul_cla32_fa16_23_and1 = s_csamul_cla32_fa16_23_xor0 & s_csamul_cla32_fa16_22_or0;
  assign s_csamul_cla32_fa16_23_or0 = s_csamul_cla32_fa16_23_and0 | s_csamul_cla32_fa16_23_and1;
  assign s_csamul_cla32_and17_23 = a[17] & b[23];
  assign s_csamul_cla32_fa17_23_xor0 = s_csamul_cla32_and17_23 ^ s_csamul_cla32_fa18_22_xor1;
  assign s_csamul_cla32_fa17_23_and0 = s_csamul_cla32_and17_23 & s_csamul_cla32_fa18_22_xor1;
  assign s_csamul_cla32_fa17_23_xor1 = s_csamul_cla32_fa17_23_xor0 ^ s_csamul_cla32_fa17_22_or0;
  assign s_csamul_cla32_fa17_23_and1 = s_csamul_cla32_fa17_23_xor0 & s_csamul_cla32_fa17_22_or0;
  assign s_csamul_cla32_fa17_23_or0 = s_csamul_cla32_fa17_23_and0 | s_csamul_cla32_fa17_23_and1;
  assign s_csamul_cla32_and18_23 = a[18] & b[23];
  assign s_csamul_cla32_fa18_23_xor0 = s_csamul_cla32_and18_23 ^ s_csamul_cla32_fa19_22_xor1;
  assign s_csamul_cla32_fa18_23_and0 = s_csamul_cla32_and18_23 & s_csamul_cla32_fa19_22_xor1;
  assign s_csamul_cla32_fa18_23_xor1 = s_csamul_cla32_fa18_23_xor0 ^ s_csamul_cla32_fa18_22_or0;
  assign s_csamul_cla32_fa18_23_and1 = s_csamul_cla32_fa18_23_xor0 & s_csamul_cla32_fa18_22_or0;
  assign s_csamul_cla32_fa18_23_or0 = s_csamul_cla32_fa18_23_and0 | s_csamul_cla32_fa18_23_and1;
  assign s_csamul_cla32_and19_23 = a[19] & b[23];
  assign s_csamul_cla32_fa19_23_xor0 = s_csamul_cla32_and19_23 ^ s_csamul_cla32_fa20_22_xor1;
  assign s_csamul_cla32_fa19_23_and0 = s_csamul_cla32_and19_23 & s_csamul_cla32_fa20_22_xor1;
  assign s_csamul_cla32_fa19_23_xor1 = s_csamul_cla32_fa19_23_xor0 ^ s_csamul_cla32_fa19_22_or0;
  assign s_csamul_cla32_fa19_23_and1 = s_csamul_cla32_fa19_23_xor0 & s_csamul_cla32_fa19_22_or0;
  assign s_csamul_cla32_fa19_23_or0 = s_csamul_cla32_fa19_23_and0 | s_csamul_cla32_fa19_23_and1;
  assign s_csamul_cla32_and20_23 = a[20] & b[23];
  assign s_csamul_cla32_fa20_23_xor0 = s_csamul_cla32_and20_23 ^ s_csamul_cla32_fa21_22_xor1;
  assign s_csamul_cla32_fa20_23_and0 = s_csamul_cla32_and20_23 & s_csamul_cla32_fa21_22_xor1;
  assign s_csamul_cla32_fa20_23_xor1 = s_csamul_cla32_fa20_23_xor0 ^ s_csamul_cla32_fa20_22_or0;
  assign s_csamul_cla32_fa20_23_and1 = s_csamul_cla32_fa20_23_xor0 & s_csamul_cla32_fa20_22_or0;
  assign s_csamul_cla32_fa20_23_or0 = s_csamul_cla32_fa20_23_and0 | s_csamul_cla32_fa20_23_and1;
  assign s_csamul_cla32_and21_23 = a[21] & b[23];
  assign s_csamul_cla32_fa21_23_xor0 = s_csamul_cla32_and21_23 ^ s_csamul_cla32_fa22_22_xor1;
  assign s_csamul_cla32_fa21_23_and0 = s_csamul_cla32_and21_23 & s_csamul_cla32_fa22_22_xor1;
  assign s_csamul_cla32_fa21_23_xor1 = s_csamul_cla32_fa21_23_xor0 ^ s_csamul_cla32_fa21_22_or0;
  assign s_csamul_cla32_fa21_23_and1 = s_csamul_cla32_fa21_23_xor0 & s_csamul_cla32_fa21_22_or0;
  assign s_csamul_cla32_fa21_23_or0 = s_csamul_cla32_fa21_23_and0 | s_csamul_cla32_fa21_23_and1;
  assign s_csamul_cla32_and22_23 = a[22] & b[23];
  assign s_csamul_cla32_fa22_23_xor0 = s_csamul_cla32_and22_23 ^ s_csamul_cla32_fa23_22_xor1;
  assign s_csamul_cla32_fa22_23_and0 = s_csamul_cla32_and22_23 & s_csamul_cla32_fa23_22_xor1;
  assign s_csamul_cla32_fa22_23_xor1 = s_csamul_cla32_fa22_23_xor0 ^ s_csamul_cla32_fa22_22_or0;
  assign s_csamul_cla32_fa22_23_and1 = s_csamul_cla32_fa22_23_xor0 & s_csamul_cla32_fa22_22_or0;
  assign s_csamul_cla32_fa22_23_or0 = s_csamul_cla32_fa22_23_and0 | s_csamul_cla32_fa22_23_and1;
  assign s_csamul_cla32_and23_23 = a[23] & b[23];
  assign s_csamul_cla32_fa23_23_xor0 = s_csamul_cla32_and23_23 ^ s_csamul_cla32_fa24_22_xor1;
  assign s_csamul_cla32_fa23_23_and0 = s_csamul_cla32_and23_23 & s_csamul_cla32_fa24_22_xor1;
  assign s_csamul_cla32_fa23_23_xor1 = s_csamul_cla32_fa23_23_xor0 ^ s_csamul_cla32_fa23_22_or0;
  assign s_csamul_cla32_fa23_23_and1 = s_csamul_cla32_fa23_23_xor0 & s_csamul_cla32_fa23_22_or0;
  assign s_csamul_cla32_fa23_23_or0 = s_csamul_cla32_fa23_23_and0 | s_csamul_cla32_fa23_23_and1;
  assign s_csamul_cla32_and24_23 = a[24] & b[23];
  assign s_csamul_cla32_fa24_23_xor0 = s_csamul_cla32_and24_23 ^ s_csamul_cla32_fa25_22_xor1;
  assign s_csamul_cla32_fa24_23_and0 = s_csamul_cla32_and24_23 & s_csamul_cla32_fa25_22_xor1;
  assign s_csamul_cla32_fa24_23_xor1 = s_csamul_cla32_fa24_23_xor0 ^ s_csamul_cla32_fa24_22_or0;
  assign s_csamul_cla32_fa24_23_and1 = s_csamul_cla32_fa24_23_xor0 & s_csamul_cla32_fa24_22_or0;
  assign s_csamul_cla32_fa24_23_or0 = s_csamul_cla32_fa24_23_and0 | s_csamul_cla32_fa24_23_and1;
  assign s_csamul_cla32_and25_23 = a[25] & b[23];
  assign s_csamul_cla32_fa25_23_xor0 = s_csamul_cla32_and25_23 ^ s_csamul_cla32_fa26_22_xor1;
  assign s_csamul_cla32_fa25_23_and0 = s_csamul_cla32_and25_23 & s_csamul_cla32_fa26_22_xor1;
  assign s_csamul_cla32_fa25_23_xor1 = s_csamul_cla32_fa25_23_xor0 ^ s_csamul_cla32_fa25_22_or0;
  assign s_csamul_cla32_fa25_23_and1 = s_csamul_cla32_fa25_23_xor0 & s_csamul_cla32_fa25_22_or0;
  assign s_csamul_cla32_fa25_23_or0 = s_csamul_cla32_fa25_23_and0 | s_csamul_cla32_fa25_23_and1;
  assign s_csamul_cla32_and26_23 = a[26] & b[23];
  assign s_csamul_cla32_fa26_23_xor0 = s_csamul_cla32_and26_23 ^ s_csamul_cla32_fa27_22_xor1;
  assign s_csamul_cla32_fa26_23_and0 = s_csamul_cla32_and26_23 & s_csamul_cla32_fa27_22_xor1;
  assign s_csamul_cla32_fa26_23_xor1 = s_csamul_cla32_fa26_23_xor0 ^ s_csamul_cla32_fa26_22_or0;
  assign s_csamul_cla32_fa26_23_and1 = s_csamul_cla32_fa26_23_xor0 & s_csamul_cla32_fa26_22_or0;
  assign s_csamul_cla32_fa26_23_or0 = s_csamul_cla32_fa26_23_and0 | s_csamul_cla32_fa26_23_and1;
  assign s_csamul_cla32_and27_23 = a[27] & b[23];
  assign s_csamul_cla32_fa27_23_xor0 = s_csamul_cla32_and27_23 ^ s_csamul_cla32_fa28_22_xor1;
  assign s_csamul_cla32_fa27_23_and0 = s_csamul_cla32_and27_23 & s_csamul_cla32_fa28_22_xor1;
  assign s_csamul_cla32_fa27_23_xor1 = s_csamul_cla32_fa27_23_xor0 ^ s_csamul_cla32_fa27_22_or0;
  assign s_csamul_cla32_fa27_23_and1 = s_csamul_cla32_fa27_23_xor0 & s_csamul_cla32_fa27_22_or0;
  assign s_csamul_cla32_fa27_23_or0 = s_csamul_cla32_fa27_23_and0 | s_csamul_cla32_fa27_23_and1;
  assign s_csamul_cla32_and28_23 = a[28] & b[23];
  assign s_csamul_cla32_fa28_23_xor0 = s_csamul_cla32_and28_23 ^ s_csamul_cla32_fa29_22_xor1;
  assign s_csamul_cla32_fa28_23_and0 = s_csamul_cla32_and28_23 & s_csamul_cla32_fa29_22_xor1;
  assign s_csamul_cla32_fa28_23_xor1 = s_csamul_cla32_fa28_23_xor0 ^ s_csamul_cla32_fa28_22_or0;
  assign s_csamul_cla32_fa28_23_and1 = s_csamul_cla32_fa28_23_xor0 & s_csamul_cla32_fa28_22_or0;
  assign s_csamul_cla32_fa28_23_or0 = s_csamul_cla32_fa28_23_and0 | s_csamul_cla32_fa28_23_and1;
  assign s_csamul_cla32_and29_23 = a[29] & b[23];
  assign s_csamul_cla32_fa29_23_xor0 = s_csamul_cla32_and29_23 ^ s_csamul_cla32_fa30_22_xor1;
  assign s_csamul_cla32_fa29_23_and0 = s_csamul_cla32_and29_23 & s_csamul_cla32_fa30_22_xor1;
  assign s_csamul_cla32_fa29_23_xor1 = s_csamul_cla32_fa29_23_xor0 ^ s_csamul_cla32_fa29_22_or0;
  assign s_csamul_cla32_fa29_23_and1 = s_csamul_cla32_fa29_23_xor0 & s_csamul_cla32_fa29_22_or0;
  assign s_csamul_cla32_fa29_23_or0 = s_csamul_cla32_fa29_23_and0 | s_csamul_cla32_fa29_23_and1;
  assign s_csamul_cla32_and30_23 = a[30] & b[23];
  assign s_csamul_cla32_fa30_23_xor0 = s_csamul_cla32_and30_23 ^ s_csamul_cla32_ha31_22_xor0;
  assign s_csamul_cla32_fa30_23_and0 = s_csamul_cla32_and30_23 & s_csamul_cla32_ha31_22_xor0;
  assign s_csamul_cla32_fa30_23_xor1 = s_csamul_cla32_fa30_23_xor0 ^ s_csamul_cla32_fa30_22_or0;
  assign s_csamul_cla32_fa30_23_and1 = s_csamul_cla32_fa30_23_xor0 & s_csamul_cla32_fa30_22_or0;
  assign s_csamul_cla32_fa30_23_or0 = s_csamul_cla32_fa30_23_and0 | s_csamul_cla32_fa30_23_and1;
  assign s_csamul_cla32_nand31_23 = ~(a[31] & b[23]);
  assign s_csamul_cla32_ha31_23_xor0 = s_csamul_cla32_nand31_23 ^ s_csamul_cla32_ha31_22_and0;
  assign s_csamul_cla32_ha31_23_and0 = s_csamul_cla32_nand31_23 & s_csamul_cla32_ha31_22_and0;
  assign s_csamul_cla32_and0_24 = a[0] & b[24];
  assign s_csamul_cla32_fa0_24_xor0 = s_csamul_cla32_and0_24 ^ s_csamul_cla32_fa1_23_xor1;
  assign s_csamul_cla32_fa0_24_and0 = s_csamul_cla32_and0_24 & s_csamul_cla32_fa1_23_xor1;
  assign s_csamul_cla32_fa0_24_xor1 = s_csamul_cla32_fa0_24_xor0 ^ s_csamul_cla32_fa0_23_or0;
  assign s_csamul_cla32_fa0_24_and1 = s_csamul_cla32_fa0_24_xor0 & s_csamul_cla32_fa0_23_or0;
  assign s_csamul_cla32_fa0_24_or0 = s_csamul_cla32_fa0_24_and0 | s_csamul_cla32_fa0_24_and1;
  assign s_csamul_cla32_and1_24 = a[1] & b[24];
  assign s_csamul_cla32_fa1_24_xor0 = s_csamul_cla32_and1_24 ^ s_csamul_cla32_fa2_23_xor1;
  assign s_csamul_cla32_fa1_24_and0 = s_csamul_cla32_and1_24 & s_csamul_cla32_fa2_23_xor1;
  assign s_csamul_cla32_fa1_24_xor1 = s_csamul_cla32_fa1_24_xor0 ^ s_csamul_cla32_fa1_23_or0;
  assign s_csamul_cla32_fa1_24_and1 = s_csamul_cla32_fa1_24_xor0 & s_csamul_cla32_fa1_23_or0;
  assign s_csamul_cla32_fa1_24_or0 = s_csamul_cla32_fa1_24_and0 | s_csamul_cla32_fa1_24_and1;
  assign s_csamul_cla32_and2_24 = a[2] & b[24];
  assign s_csamul_cla32_fa2_24_xor0 = s_csamul_cla32_and2_24 ^ s_csamul_cla32_fa3_23_xor1;
  assign s_csamul_cla32_fa2_24_and0 = s_csamul_cla32_and2_24 & s_csamul_cla32_fa3_23_xor1;
  assign s_csamul_cla32_fa2_24_xor1 = s_csamul_cla32_fa2_24_xor0 ^ s_csamul_cla32_fa2_23_or0;
  assign s_csamul_cla32_fa2_24_and1 = s_csamul_cla32_fa2_24_xor0 & s_csamul_cla32_fa2_23_or0;
  assign s_csamul_cla32_fa2_24_or0 = s_csamul_cla32_fa2_24_and0 | s_csamul_cla32_fa2_24_and1;
  assign s_csamul_cla32_and3_24 = a[3] & b[24];
  assign s_csamul_cla32_fa3_24_xor0 = s_csamul_cla32_and3_24 ^ s_csamul_cla32_fa4_23_xor1;
  assign s_csamul_cla32_fa3_24_and0 = s_csamul_cla32_and3_24 & s_csamul_cla32_fa4_23_xor1;
  assign s_csamul_cla32_fa3_24_xor1 = s_csamul_cla32_fa3_24_xor0 ^ s_csamul_cla32_fa3_23_or0;
  assign s_csamul_cla32_fa3_24_and1 = s_csamul_cla32_fa3_24_xor0 & s_csamul_cla32_fa3_23_or0;
  assign s_csamul_cla32_fa3_24_or0 = s_csamul_cla32_fa3_24_and0 | s_csamul_cla32_fa3_24_and1;
  assign s_csamul_cla32_and4_24 = a[4] & b[24];
  assign s_csamul_cla32_fa4_24_xor0 = s_csamul_cla32_and4_24 ^ s_csamul_cla32_fa5_23_xor1;
  assign s_csamul_cla32_fa4_24_and0 = s_csamul_cla32_and4_24 & s_csamul_cla32_fa5_23_xor1;
  assign s_csamul_cla32_fa4_24_xor1 = s_csamul_cla32_fa4_24_xor0 ^ s_csamul_cla32_fa4_23_or0;
  assign s_csamul_cla32_fa4_24_and1 = s_csamul_cla32_fa4_24_xor0 & s_csamul_cla32_fa4_23_or0;
  assign s_csamul_cla32_fa4_24_or0 = s_csamul_cla32_fa4_24_and0 | s_csamul_cla32_fa4_24_and1;
  assign s_csamul_cla32_and5_24 = a[5] & b[24];
  assign s_csamul_cla32_fa5_24_xor0 = s_csamul_cla32_and5_24 ^ s_csamul_cla32_fa6_23_xor1;
  assign s_csamul_cla32_fa5_24_and0 = s_csamul_cla32_and5_24 & s_csamul_cla32_fa6_23_xor1;
  assign s_csamul_cla32_fa5_24_xor1 = s_csamul_cla32_fa5_24_xor0 ^ s_csamul_cla32_fa5_23_or0;
  assign s_csamul_cla32_fa5_24_and1 = s_csamul_cla32_fa5_24_xor0 & s_csamul_cla32_fa5_23_or0;
  assign s_csamul_cla32_fa5_24_or0 = s_csamul_cla32_fa5_24_and0 | s_csamul_cla32_fa5_24_and1;
  assign s_csamul_cla32_and6_24 = a[6] & b[24];
  assign s_csamul_cla32_fa6_24_xor0 = s_csamul_cla32_and6_24 ^ s_csamul_cla32_fa7_23_xor1;
  assign s_csamul_cla32_fa6_24_and0 = s_csamul_cla32_and6_24 & s_csamul_cla32_fa7_23_xor1;
  assign s_csamul_cla32_fa6_24_xor1 = s_csamul_cla32_fa6_24_xor0 ^ s_csamul_cla32_fa6_23_or0;
  assign s_csamul_cla32_fa6_24_and1 = s_csamul_cla32_fa6_24_xor0 & s_csamul_cla32_fa6_23_or0;
  assign s_csamul_cla32_fa6_24_or0 = s_csamul_cla32_fa6_24_and0 | s_csamul_cla32_fa6_24_and1;
  assign s_csamul_cla32_and7_24 = a[7] & b[24];
  assign s_csamul_cla32_fa7_24_xor0 = s_csamul_cla32_and7_24 ^ s_csamul_cla32_fa8_23_xor1;
  assign s_csamul_cla32_fa7_24_and0 = s_csamul_cla32_and7_24 & s_csamul_cla32_fa8_23_xor1;
  assign s_csamul_cla32_fa7_24_xor1 = s_csamul_cla32_fa7_24_xor0 ^ s_csamul_cla32_fa7_23_or0;
  assign s_csamul_cla32_fa7_24_and1 = s_csamul_cla32_fa7_24_xor0 & s_csamul_cla32_fa7_23_or0;
  assign s_csamul_cla32_fa7_24_or0 = s_csamul_cla32_fa7_24_and0 | s_csamul_cla32_fa7_24_and1;
  assign s_csamul_cla32_and8_24 = a[8] & b[24];
  assign s_csamul_cla32_fa8_24_xor0 = s_csamul_cla32_and8_24 ^ s_csamul_cla32_fa9_23_xor1;
  assign s_csamul_cla32_fa8_24_and0 = s_csamul_cla32_and8_24 & s_csamul_cla32_fa9_23_xor1;
  assign s_csamul_cla32_fa8_24_xor1 = s_csamul_cla32_fa8_24_xor0 ^ s_csamul_cla32_fa8_23_or0;
  assign s_csamul_cla32_fa8_24_and1 = s_csamul_cla32_fa8_24_xor0 & s_csamul_cla32_fa8_23_or0;
  assign s_csamul_cla32_fa8_24_or0 = s_csamul_cla32_fa8_24_and0 | s_csamul_cla32_fa8_24_and1;
  assign s_csamul_cla32_and9_24 = a[9] & b[24];
  assign s_csamul_cla32_fa9_24_xor0 = s_csamul_cla32_and9_24 ^ s_csamul_cla32_fa10_23_xor1;
  assign s_csamul_cla32_fa9_24_and0 = s_csamul_cla32_and9_24 & s_csamul_cla32_fa10_23_xor1;
  assign s_csamul_cla32_fa9_24_xor1 = s_csamul_cla32_fa9_24_xor0 ^ s_csamul_cla32_fa9_23_or0;
  assign s_csamul_cla32_fa9_24_and1 = s_csamul_cla32_fa9_24_xor0 & s_csamul_cla32_fa9_23_or0;
  assign s_csamul_cla32_fa9_24_or0 = s_csamul_cla32_fa9_24_and0 | s_csamul_cla32_fa9_24_and1;
  assign s_csamul_cla32_and10_24 = a[10] & b[24];
  assign s_csamul_cla32_fa10_24_xor0 = s_csamul_cla32_and10_24 ^ s_csamul_cla32_fa11_23_xor1;
  assign s_csamul_cla32_fa10_24_and0 = s_csamul_cla32_and10_24 & s_csamul_cla32_fa11_23_xor1;
  assign s_csamul_cla32_fa10_24_xor1 = s_csamul_cla32_fa10_24_xor0 ^ s_csamul_cla32_fa10_23_or0;
  assign s_csamul_cla32_fa10_24_and1 = s_csamul_cla32_fa10_24_xor0 & s_csamul_cla32_fa10_23_or0;
  assign s_csamul_cla32_fa10_24_or0 = s_csamul_cla32_fa10_24_and0 | s_csamul_cla32_fa10_24_and1;
  assign s_csamul_cla32_and11_24 = a[11] & b[24];
  assign s_csamul_cla32_fa11_24_xor0 = s_csamul_cla32_and11_24 ^ s_csamul_cla32_fa12_23_xor1;
  assign s_csamul_cla32_fa11_24_and0 = s_csamul_cla32_and11_24 & s_csamul_cla32_fa12_23_xor1;
  assign s_csamul_cla32_fa11_24_xor1 = s_csamul_cla32_fa11_24_xor0 ^ s_csamul_cla32_fa11_23_or0;
  assign s_csamul_cla32_fa11_24_and1 = s_csamul_cla32_fa11_24_xor0 & s_csamul_cla32_fa11_23_or0;
  assign s_csamul_cla32_fa11_24_or0 = s_csamul_cla32_fa11_24_and0 | s_csamul_cla32_fa11_24_and1;
  assign s_csamul_cla32_and12_24 = a[12] & b[24];
  assign s_csamul_cla32_fa12_24_xor0 = s_csamul_cla32_and12_24 ^ s_csamul_cla32_fa13_23_xor1;
  assign s_csamul_cla32_fa12_24_and0 = s_csamul_cla32_and12_24 & s_csamul_cla32_fa13_23_xor1;
  assign s_csamul_cla32_fa12_24_xor1 = s_csamul_cla32_fa12_24_xor0 ^ s_csamul_cla32_fa12_23_or0;
  assign s_csamul_cla32_fa12_24_and1 = s_csamul_cla32_fa12_24_xor0 & s_csamul_cla32_fa12_23_or0;
  assign s_csamul_cla32_fa12_24_or0 = s_csamul_cla32_fa12_24_and0 | s_csamul_cla32_fa12_24_and1;
  assign s_csamul_cla32_and13_24 = a[13] & b[24];
  assign s_csamul_cla32_fa13_24_xor0 = s_csamul_cla32_and13_24 ^ s_csamul_cla32_fa14_23_xor1;
  assign s_csamul_cla32_fa13_24_and0 = s_csamul_cla32_and13_24 & s_csamul_cla32_fa14_23_xor1;
  assign s_csamul_cla32_fa13_24_xor1 = s_csamul_cla32_fa13_24_xor0 ^ s_csamul_cla32_fa13_23_or0;
  assign s_csamul_cla32_fa13_24_and1 = s_csamul_cla32_fa13_24_xor0 & s_csamul_cla32_fa13_23_or0;
  assign s_csamul_cla32_fa13_24_or0 = s_csamul_cla32_fa13_24_and0 | s_csamul_cla32_fa13_24_and1;
  assign s_csamul_cla32_and14_24 = a[14] & b[24];
  assign s_csamul_cla32_fa14_24_xor0 = s_csamul_cla32_and14_24 ^ s_csamul_cla32_fa15_23_xor1;
  assign s_csamul_cla32_fa14_24_and0 = s_csamul_cla32_and14_24 & s_csamul_cla32_fa15_23_xor1;
  assign s_csamul_cla32_fa14_24_xor1 = s_csamul_cla32_fa14_24_xor0 ^ s_csamul_cla32_fa14_23_or0;
  assign s_csamul_cla32_fa14_24_and1 = s_csamul_cla32_fa14_24_xor0 & s_csamul_cla32_fa14_23_or0;
  assign s_csamul_cla32_fa14_24_or0 = s_csamul_cla32_fa14_24_and0 | s_csamul_cla32_fa14_24_and1;
  assign s_csamul_cla32_and15_24 = a[15] & b[24];
  assign s_csamul_cla32_fa15_24_xor0 = s_csamul_cla32_and15_24 ^ s_csamul_cla32_fa16_23_xor1;
  assign s_csamul_cla32_fa15_24_and0 = s_csamul_cla32_and15_24 & s_csamul_cla32_fa16_23_xor1;
  assign s_csamul_cla32_fa15_24_xor1 = s_csamul_cla32_fa15_24_xor0 ^ s_csamul_cla32_fa15_23_or0;
  assign s_csamul_cla32_fa15_24_and1 = s_csamul_cla32_fa15_24_xor0 & s_csamul_cla32_fa15_23_or0;
  assign s_csamul_cla32_fa15_24_or0 = s_csamul_cla32_fa15_24_and0 | s_csamul_cla32_fa15_24_and1;
  assign s_csamul_cla32_and16_24 = a[16] & b[24];
  assign s_csamul_cla32_fa16_24_xor0 = s_csamul_cla32_and16_24 ^ s_csamul_cla32_fa17_23_xor1;
  assign s_csamul_cla32_fa16_24_and0 = s_csamul_cla32_and16_24 & s_csamul_cla32_fa17_23_xor1;
  assign s_csamul_cla32_fa16_24_xor1 = s_csamul_cla32_fa16_24_xor0 ^ s_csamul_cla32_fa16_23_or0;
  assign s_csamul_cla32_fa16_24_and1 = s_csamul_cla32_fa16_24_xor0 & s_csamul_cla32_fa16_23_or0;
  assign s_csamul_cla32_fa16_24_or0 = s_csamul_cla32_fa16_24_and0 | s_csamul_cla32_fa16_24_and1;
  assign s_csamul_cla32_and17_24 = a[17] & b[24];
  assign s_csamul_cla32_fa17_24_xor0 = s_csamul_cla32_and17_24 ^ s_csamul_cla32_fa18_23_xor1;
  assign s_csamul_cla32_fa17_24_and0 = s_csamul_cla32_and17_24 & s_csamul_cla32_fa18_23_xor1;
  assign s_csamul_cla32_fa17_24_xor1 = s_csamul_cla32_fa17_24_xor0 ^ s_csamul_cla32_fa17_23_or0;
  assign s_csamul_cla32_fa17_24_and1 = s_csamul_cla32_fa17_24_xor0 & s_csamul_cla32_fa17_23_or0;
  assign s_csamul_cla32_fa17_24_or0 = s_csamul_cla32_fa17_24_and0 | s_csamul_cla32_fa17_24_and1;
  assign s_csamul_cla32_and18_24 = a[18] & b[24];
  assign s_csamul_cla32_fa18_24_xor0 = s_csamul_cla32_and18_24 ^ s_csamul_cla32_fa19_23_xor1;
  assign s_csamul_cla32_fa18_24_and0 = s_csamul_cla32_and18_24 & s_csamul_cla32_fa19_23_xor1;
  assign s_csamul_cla32_fa18_24_xor1 = s_csamul_cla32_fa18_24_xor0 ^ s_csamul_cla32_fa18_23_or0;
  assign s_csamul_cla32_fa18_24_and1 = s_csamul_cla32_fa18_24_xor0 & s_csamul_cla32_fa18_23_or0;
  assign s_csamul_cla32_fa18_24_or0 = s_csamul_cla32_fa18_24_and0 | s_csamul_cla32_fa18_24_and1;
  assign s_csamul_cla32_and19_24 = a[19] & b[24];
  assign s_csamul_cla32_fa19_24_xor0 = s_csamul_cla32_and19_24 ^ s_csamul_cla32_fa20_23_xor1;
  assign s_csamul_cla32_fa19_24_and0 = s_csamul_cla32_and19_24 & s_csamul_cla32_fa20_23_xor1;
  assign s_csamul_cla32_fa19_24_xor1 = s_csamul_cla32_fa19_24_xor0 ^ s_csamul_cla32_fa19_23_or0;
  assign s_csamul_cla32_fa19_24_and1 = s_csamul_cla32_fa19_24_xor0 & s_csamul_cla32_fa19_23_or0;
  assign s_csamul_cla32_fa19_24_or0 = s_csamul_cla32_fa19_24_and0 | s_csamul_cla32_fa19_24_and1;
  assign s_csamul_cla32_and20_24 = a[20] & b[24];
  assign s_csamul_cla32_fa20_24_xor0 = s_csamul_cla32_and20_24 ^ s_csamul_cla32_fa21_23_xor1;
  assign s_csamul_cla32_fa20_24_and0 = s_csamul_cla32_and20_24 & s_csamul_cla32_fa21_23_xor1;
  assign s_csamul_cla32_fa20_24_xor1 = s_csamul_cla32_fa20_24_xor0 ^ s_csamul_cla32_fa20_23_or0;
  assign s_csamul_cla32_fa20_24_and1 = s_csamul_cla32_fa20_24_xor0 & s_csamul_cla32_fa20_23_or0;
  assign s_csamul_cla32_fa20_24_or0 = s_csamul_cla32_fa20_24_and0 | s_csamul_cla32_fa20_24_and1;
  assign s_csamul_cla32_and21_24 = a[21] & b[24];
  assign s_csamul_cla32_fa21_24_xor0 = s_csamul_cla32_and21_24 ^ s_csamul_cla32_fa22_23_xor1;
  assign s_csamul_cla32_fa21_24_and0 = s_csamul_cla32_and21_24 & s_csamul_cla32_fa22_23_xor1;
  assign s_csamul_cla32_fa21_24_xor1 = s_csamul_cla32_fa21_24_xor0 ^ s_csamul_cla32_fa21_23_or0;
  assign s_csamul_cla32_fa21_24_and1 = s_csamul_cla32_fa21_24_xor0 & s_csamul_cla32_fa21_23_or0;
  assign s_csamul_cla32_fa21_24_or0 = s_csamul_cla32_fa21_24_and0 | s_csamul_cla32_fa21_24_and1;
  assign s_csamul_cla32_and22_24 = a[22] & b[24];
  assign s_csamul_cla32_fa22_24_xor0 = s_csamul_cla32_and22_24 ^ s_csamul_cla32_fa23_23_xor1;
  assign s_csamul_cla32_fa22_24_and0 = s_csamul_cla32_and22_24 & s_csamul_cla32_fa23_23_xor1;
  assign s_csamul_cla32_fa22_24_xor1 = s_csamul_cla32_fa22_24_xor0 ^ s_csamul_cla32_fa22_23_or0;
  assign s_csamul_cla32_fa22_24_and1 = s_csamul_cla32_fa22_24_xor0 & s_csamul_cla32_fa22_23_or0;
  assign s_csamul_cla32_fa22_24_or0 = s_csamul_cla32_fa22_24_and0 | s_csamul_cla32_fa22_24_and1;
  assign s_csamul_cla32_and23_24 = a[23] & b[24];
  assign s_csamul_cla32_fa23_24_xor0 = s_csamul_cla32_and23_24 ^ s_csamul_cla32_fa24_23_xor1;
  assign s_csamul_cla32_fa23_24_and0 = s_csamul_cla32_and23_24 & s_csamul_cla32_fa24_23_xor1;
  assign s_csamul_cla32_fa23_24_xor1 = s_csamul_cla32_fa23_24_xor0 ^ s_csamul_cla32_fa23_23_or0;
  assign s_csamul_cla32_fa23_24_and1 = s_csamul_cla32_fa23_24_xor0 & s_csamul_cla32_fa23_23_or0;
  assign s_csamul_cla32_fa23_24_or0 = s_csamul_cla32_fa23_24_and0 | s_csamul_cla32_fa23_24_and1;
  assign s_csamul_cla32_and24_24 = a[24] & b[24];
  assign s_csamul_cla32_fa24_24_xor0 = s_csamul_cla32_and24_24 ^ s_csamul_cla32_fa25_23_xor1;
  assign s_csamul_cla32_fa24_24_and0 = s_csamul_cla32_and24_24 & s_csamul_cla32_fa25_23_xor1;
  assign s_csamul_cla32_fa24_24_xor1 = s_csamul_cla32_fa24_24_xor0 ^ s_csamul_cla32_fa24_23_or0;
  assign s_csamul_cla32_fa24_24_and1 = s_csamul_cla32_fa24_24_xor0 & s_csamul_cla32_fa24_23_or0;
  assign s_csamul_cla32_fa24_24_or0 = s_csamul_cla32_fa24_24_and0 | s_csamul_cla32_fa24_24_and1;
  assign s_csamul_cla32_and25_24 = a[25] & b[24];
  assign s_csamul_cla32_fa25_24_xor0 = s_csamul_cla32_and25_24 ^ s_csamul_cla32_fa26_23_xor1;
  assign s_csamul_cla32_fa25_24_and0 = s_csamul_cla32_and25_24 & s_csamul_cla32_fa26_23_xor1;
  assign s_csamul_cla32_fa25_24_xor1 = s_csamul_cla32_fa25_24_xor0 ^ s_csamul_cla32_fa25_23_or0;
  assign s_csamul_cla32_fa25_24_and1 = s_csamul_cla32_fa25_24_xor0 & s_csamul_cla32_fa25_23_or0;
  assign s_csamul_cla32_fa25_24_or0 = s_csamul_cla32_fa25_24_and0 | s_csamul_cla32_fa25_24_and1;
  assign s_csamul_cla32_and26_24 = a[26] & b[24];
  assign s_csamul_cla32_fa26_24_xor0 = s_csamul_cla32_and26_24 ^ s_csamul_cla32_fa27_23_xor1;
  assign s_csamul_cla32_fa26_24_and0 = s_csamul_cla32_and26_24 & s_csamul_cla32_fa27_23_xor1;
  assign s_csamul_cla32_fa26_24_xor1 = s_csamul_cla32_fa26_24_xor0 ^ s_csamul_cla32_fa26_23_or0;
  assign s_csamul_cla32_fa26_24_and1 = s_csamul_cla32_fa26_24_xor0 & s_csamul_cla32_fa26_23_or0;
  assign s_csamul_cla32_fa26_24_or0 = s_csamul_cla32_fa26_24_and0 | s_csamul_cla32_fa26_24_and1;
  assign s_csamul_cla32_and27_24 = a[27] & b[24];
  assign s_csamul_cla32_fa27_24_xor0 = s_csamul_cla32_and27_24 ^ s_csamul_cla32_fa28_23_xor1;
  assign s_csamul_cla32_fa27_24_and0 = s_csamul_cla32_and27_24 & s_csamul_cla32_fa28_23_xor1;
  assign s_csamul_cla32_fa27_24_xor1 = s_csamul_cla32_fa27_24_xor0 ^ s_csamul_cla32_fa27_23_or0;
  assign s_csamul_cla32_fa27_24_and1 = s_csamul_cla32_fa27_24_xor0 & s_csamul_cla32_fa27_23_or0;
  assign s_csamul_cla32_fa27_24_or0 = s_csamul_cla32_fa27_24_and0 | s_csamul_cla32_fa27_24_and1;
  assign s_csamul_cla32_and28_24 = a[28] & b[24];
  assign s_csamul_cla32_fa28_24_xor0 = s_csamul_cla32_and28_24 ^ s_csamul_cla32_fa29_23_xor1;
  assign s_csamul_cla32_fa28_24_and0 = s_csamul_cla32_and28_24 & s_csamul_cla32_fa29_23_xor1;
  assign s_csamul_cla32_fa28_24_xor1 = s_csamul_cla32_fa28_24_xor0 ^ s_csamul_cla32_fa28_23_or0;
  assign s_csamul_cla32_fa28_24_and1 = s_csamul_cla32_fa28_24_xor0 & s_csamul_cla32_fa28_23_or0;
  assign s_csamul_cla32_fa28_24_or0 = s_csamul_cla32_fa28_24_and0 | s_csamul_cla32_fa28_24_and1;
  assign s_csamul_cla32_and29_24 = a[29] & b[24];
  assign s_csamul_cla32_fa29_24_xor0 = s_csamul_cla32_and29_24 ^ s_csamul_cla32_fa30_23_xor1;
  assign s_csamul_cla32_fa29_24_and0 = s_csamul_cla32_and29_24 & s_csamul_cla32_fa30_23_xor1;
  assign s_csamul_cla32_fa29_24_xor1 = s_csamul_cla32_fa29_24_xor0 ^ s_csamul_cla32_fa29_23_or0;
  assign s_csamul_cla32_fa29_24_and1 = s_csamul_cla32_fa29_24_xor0 & s_csamul_cla32_fa29_23_or0;
  assign s_csamul_cla32_fa29_24_or0 = s_csamul_cla32_fa29_24_and0 | s_csamul_cla32_fa29_24_and1;
  assign s_csamul_cla32_and30_24 = a[30] & b[24];
  assign s_csamul_cla32_fa30_24_xor0 = s_csamul_cla32_and30_24 ^ s_csamul_cla32_ha31_23_xor0;
  assign s_csamul_cla32_fa30_24_and0 = s_csamul_cla32_and30_24 & s_csamul_cla32_ha31_23_xor0;
  assign s_csamul_cla32_fa30_24_xor1 = s_csamul_cla32_fa30_24_xor0 ^ s_csamul_cla32_fa30_23_or0;
  assign s_csamul_cla32_fa30_24_and1 = s_csamul_cla32_fa30_24_xor0 & s_csamul_cla32_fa30_23_or0;
  assign s_csamul_cla32_fa30_24_or0 = s_csamul_cla32_fa30_24_and0 | s_csamul_cla32_fa30_24_and1;
  assign s_csamul_cla32_nand31_24 = ~(a[31] & b[24]);
  assign s_csamul_cla32_ha31_24_xor0 = s_csamul_cla32_nand31_24 ^ s_csamul_cla32_ha31_23_and0;
  assign s_csamul_cla32_ha31_24_and0 = s_csamul_cla32_nand31_24 & s_csamul_cla32_ha31_23_and0;
  assign s_csamul_cla32_and0_25 = a[0] & b[25];
  assign s_csamul_cla32_fa0_25_xor0 = s_csamul_cla32_and0_25 ^ s_csamul_cla32_fa1_24_xor1;
  assign s_csamul_cla32_fa0_25_and0 = s_csamul_cla32_and0_25 & s_csamul_cla32_fa1_24_xor1;
  assign s_csamul_cla32_fa0_25_xor1 = s_csamul_cla32_fa0_25_xor0 ^ s_csamul_cla32_fa0_24_or0;
  assign s_csamul_cla32_fa0_25_and1 = s_csamul_cla32_fa0_25_xor0 & s_csamul_cla32_fa0_24_or0;
  assign s_csamul_cla32_fa0_25_or0 = s_csamul_cla32_fa0_25_and0 | s_csamul_cla32_fa0_25_and1;
  assign s_csamul_cla32_and1_25 = a[1] & b[25];
  assign s_csamul_cla32_fa1_25_xor0 = s_csamul_cla32_and1_25 ^ s_csamul_cla32_fa2_24_xor1;
  assign s_csamul_cla32_fa1_25_and0 = s_csamul_cla32_and1_25 & s_csamul_cla32_fa2_24_xor1;
  assign s_csamul_cla32_fa1_25_xor1 = s_csamul_cla32_fa1_25_xor0 ^ s_csamul_cla32_fa1_24_or0;
  assign s_csamul_cla32_fa1_25_and1 = s_csamul_cla32_fa1_25_xor0 & s_csamul_cla32_fa1_24_or0;
  assign s_csamul_cla32_fa1_25_or0 = s_csamul_cla32_fa1_25_and0 | s_csamul_cla32_fa1_25_and1;
  assign s_csamul_cla32_and2_25 = a[2] & b[25];
  assign s_csamul_cla32_fa2_25_xor0 = s_csamul_cla32_and2_25 ^ s_csamul_cla32_fa3_24_xor1;
  assign s_csamul_cla32_fa2_25_and0 = s_csamul_cla32_and2_25 & s_csamul_cla32_fa3_24_xor1;
  assign s_csamul_cla32_fa2_25_xor1 = s_csamul_cla32_fa2_25_xor0 ^ s_csamul_cla32_fa2_24_or0;
  assign s_csamul_cla32_fa2_25_and1 = s_csamul_cla32_fa2_25_xor0 & s_csamul_cla32_fa2_24_or0;
  assign s_csamul_cla32_fa2_25_or0 = s_csamul_cla32_fa2_25_and0 | s_csamul_cla32_fa2_25_and1;
  assign s_csamul_cla32_and3_25 = a[3] & b[25];
  assign s_csamul_cla32_fa3_25_xor0 = s_csamul_cla32_and3_25 ^ s_csamul_cla32_fa4_24_xor1;
  assign s_csamul_cla32_fa3_25_and0 = s_csamul_cla32_and3_25 & s_csamul_cla32_fa4_24_xor1;
  assign s_csamul_cla32_fa3_25_xor1 = s_csamul_cla32_fa3_25_xor0 ^ s_csamul_cla32_fa3_24_or0;
  assign s_csamul_cla32_fa3_25_and1 = s_csamul_cla32_fa3_25_xor0 & s_csamul_cla32_fa3_24_or0;
  assign s_csamul_cla32_fa3_25_or0 = s_csamul_cla32_fa3_25_and0 | s_csamul_cla32_fa3_25_and1;
  assign s_csamul_cla32_and4_25 = a[4] & b[25];
  assign s_csamul_cla32_fa4_25_xor0 = s_csamul_cla32_and4_25 ^ s_csamul_cla32_fa5_24_xor1;
  assign s_csamul_cla32_fa4_25_and0 = s_csamul_cla32_and4_25 & s_csamul_cla32_fa5_24_xor1;
  assign s_csamul_cla32_fa4_25_xor1 = s_csamul_cla32_fa4_25_xor0 ^ s_csamul_cla32_fa4_24_or0;
  assign s_csamul_cla32_fa4_25_and1 = s_csamul_cla32_fa4_25_xor0 & s_csamul_cla32_fa4_24_or0;
  assign s_csamul_cla32_fa4_25_or0 = s_csamul_cla32_fa4_25_and0 | s_csamul_cla32_fa4_25_and1;
  assign s_csamul_cla32_and5_25 = a[5] & b[25];
  assign s_csamul_cla32_fa5_25_xor0 = s_csamul_cla32_and5_25 ^ s_csamul_cla32_fa6_24_xor1;
  assign s_csamul_cla32_fa5_25_and0 = s_csamul_cla32_and5_25 & s_csamul_cla32_fa6_24_xor1;
  assign s_csamul_cla32_fa5_25_xor1 = s_csamul_cla32_fa5_25_xor0 ^ s_csamul_cla32_fa5_24_or0;
  assign s_csamul_cla32_fa5_25_and1 = s_csamul_cla32_fa5_25_xor0 & s_csamul_cla32_fa5_24_or0;
  assign s_csamul_cla32_fa5_25_or0 = s_csamul_cla32_fa5_25_and0 | s_csamul_cla32_fa5_25_and1;
  assign s_csamul_cla32_and6_25 = a[6] & b[25];
  assign s_csamul_cla32_fa6_25_xor0 = s_csamul_cla32_and6_25 ^ s_csamul_cla32_fa7_24_xor1;
  assign s_csamul_cla32_fa6_25_and0 = s_csamul_cla32_and6_25 & s_csamul_cla32_fa7_24_xor1;
  assign s_csamul_cla32_fa6_25_xor1 = s_csamul_cla32_fa6_25_xor0 ^ s_csamul_cla32_fa6_24_or0;
  assign s_csamul_cla32_fa6_25_and1 = s_csamul_cla32_fa6_25_xor0 & s_csamul_cla32_fa6_24_or0;
  assign s_csamul_cla32_fa6_25_or0 = s_csamul_cla32_fa6_25_and0 | s_csamul_cla32_fa6_25_and1;
  assign s_csamul_cla32_and7_25 = a[7] & b[25];
  assign s_csamul_cla32_fa7_25_xor0 = s_csamul_cla32_and7_25 ^ s_csamul_cla32_fa8_24_xor1;
  assign s_csamul_cla32_fa7_25_and0 = s_csamul_cla32_and7_25 & s_csamul_cla32_fa8_24_xor1;
  assign s_csamul_cla32_fa7_25_xor1 = s_csamul_cla32_fa7_25_xor0 ^ s_csamul_cla32_fa7_24_or0;
  assign s_csamul_cla32_fa7_25_and1 = s_csamul_cla32_fa7_25_xor0 & s_csamul_cla32_fa7_24_or0;
  assign s_csamul_cla32_fa7_25_or0 = s_csamul_cla32_fa7_25_and0 | s_csamul_cla32_fa7_25_and1;
  assign s_csamul_cla32_and8_25 = a[8] & b[25];
  assign s_csamul_cla32_fa8_25_xor0 = s_csamul_cla32_and8_25 ^ s_csamul_cla32_fa9_24_xor1;
  assign s_csamul_cla32_fa8_25_and0 = s_csamul_cla32_and8_25 & s_csamul_cla32_fa9_24_xor1;
  assign s_csamul_cla32_fa8_25_xor1 = s_csamul_cla32_fa8_25_xor0 ^ s_csamul_cla32_fa8_24_or0;
  assign s_csamul_cla32_fa8_25_and1 = s_csamul_cla32_fa8_25_xor0 & s_csamul_cla32_fa8_24_or0;
  assign s_csamul_cla32_fa8_25_or0 = s_csamul_cla32_fa8_25_and0 | s_csamul_cla32_fa8_25_and1;
  assign s_csamul_cla32_and9_25 = a[9] & b[25];
  assign s_csamul_cla32_fa9_25_xor0 = s_csamul_cla32_and9_25 ^ s_csamul_cla32_fa10_24_xor1;
  assign s_csamul_cla32_fa9_25_and0 = s_csamul_cla32_and9_25 & s_csamul_cla32_fa10_24_xor1;
  assign s_csamul_cla32_fa9_25_xor1 = s_csamul_cla32_fa9_25_xor0 ^ s_csamul_cla32_fa9_24_or0;
  assign s_csamul_cla32_fa9_25_and1 = s_csamul_cla32_fa9_25_xor0 & s_csamul_cla32_fa9_24_or0;
  assign s_csamul_cla32_fa9_25_or0 = s_csamul_cla32_fa9_25_and0 | s_csamul_cla32_fa9_25_and1;
  assign s_csamul_cla32_and10_25 = a[10] & b[25];
  assign s_csamul_cla32_fa10_25_xor0 = s_csamul_cla32_and10_25 ^ s_csamul_cla32_fa11_24_xor1;
  assign s_csamul_cla32_fa10_25_and0 = s_csamul_cla32_and10_25 & s_csamul_cla32_fa11_24_xor1;
  assign s_csamul_cla32_fa10_25_xor1 = s_csamul_cla32_fa10_25_xor0 ^ s_csamul_cla32_fa10_24_or0;
  assign s_csamul_cla32_fa10_25_and1 = s_csamul_cla32_fa10_25_xor0 & s_csamul_cla32_fa10_24_or0;
  assign s_csamul_cla32_fa10_25_or0 = s_csamul_cla32_fa10_25_and0 | s_csamul_cla32_fa10_25_and1;
  assign s_csamul_cla32_and11_25 = a[11] & b[25];
  assign s_csamul_cla32_fa11_25_xor0 = s_csamul_cla32_and11_25 ^ s_csamul_cla32_fa12_24_xor1;
  assign s_csamul_cla32_fa11_25_and0 = s_csamul_cla32_and11_25 & s_csamul_cla32_fa12_24_xor1;
  assign s_csamul_cla32_fa11_25_xor1 = s_csamul_cla32_fa11_25_xor0 ^ s_csamul_cla32_fa11_24_or0;
  assign s_csamul_cla32_fa11_25_and1 = s_csamul_cla32_fa11_25_xor0 & s_csamul_cla32_fa11_24_or0;
  assign s_csamul_cla32_fa11_25_or0 = s_csamul_cla32_fa11_25_and0 | s_csamul_cla32_fa11_25_and1;
  assign s_csamul_cla32_and12_25 = a[12] & b[25];
  assign s_csamul_cla32_fa12_25_xor0 = s_csamul_cla32_and12_25 ^ s_csamul_cla32_fa13_24_xor1;
  assign s_csamul_cla32_fa12_25_and0 = s_csamul_cla32_and12_25 & s_csamul_cla32_fa13_24_xor1;
  assign s_csamul_cla32_fa12_25_xor1 = s_csamul_cla32_fa12_25_xor0 ^ s_csamul_cla32_fa12_24_or0;
  assign s_csamul_cla32_fa12_25_and1 = s_csamul_cla32_fa12_25_xor0 & s_csamul_cla32_fa12_24_or0;
  assign s_csamul_cla32_fa12_25_or0 = s_csamul_cla32_fa12_25_and0 | s_csamul_cla32_fa12_25_and1;
  assign s_csamul_cla32_and13_25 = a[13] & b[25];
  assign s_csamul_cla32_fa13_25_xor0 = s_csamul_cla32_and13_25 ^ s_csamul_cla32_fa14_24_xor1;
  assign s_csamul_cla32_fa13_25_and0 = s_csamul_cla32_and13_25 & s_csamul_cla32_fa14_24_xor1;
  assign s_csamul_cla32_fa13_25_xor1 = s_csamul_cla32_fa13_25_xor0 ^ s_csamul_cla32_fa13_24_or0;
  assign s_csamul_cla32_fa13_25_and1 = s_csamul_cla32_fa13_25_xor0 & s_csamul_cla32_fa13_24_or0;
  assign s_csamul_cla32_fa13_25_or0 = s_csamul_cla32_fa13_25_and0 | s_csamul_cla32_fa13_25_and1;
  assign s_csamul_cla32_and14_25 = a[14] & b[25];
  assign s_csamul_cla32_fa14_25_xor0 = s_csamul_cla32_and14_25 ^ s_csamul_cla32_fa15_24_xor1;
  assign s_csamul_cla32_fa14_25_and0 = s_csamul_cla32_and14_25 & s_csamul_cla32_fa15_24_xor1;
  assign s_csamul_cla32_fa14_25_xor1 = s_csamul_cla32_fa14_25_xor0 ^ s_csamul_cla32_fa14_24_or0;
  assign s_csamul_cla32_fa14_25_and1 = s_csamul_cla32_fa14_25_xor0 & s_csamul_cla32_fa14_24_or0;
  assign s_csamul_cla32_fa14_25_or0 = s_csamul_cla32_fa14_25_and0 | s_csamul_cla32_fa14_25_and1;
  assign s_csamul_cla32_and15_25 = a[15] & b[25];
  assign s_csamul_cla32_fa15_25_xor0 = s_csamul_cla32_and15_25 ^ s_csamul_cla32_fa16_24_xor1;
  assign s_csamul_cla32_fa15_25_and0 = s_csamul_cla32_and15_25 & s_csamul_cla32_fa16_24_xor1;
  assign s_csamul_cla32_fa15_25_xor1 = s_csamul_cla32_fa15_25_xor0 ^ s_csamul_cla32_fa15_24_or0;
  assign s_csamul_cla32_fa15_25_and1 = s_csamul_cla32_fa15_25_xor0 & s_csamul_cla32_fa15_24_or0;
  assign s_csamul_cla32_fa15_25_or0 = s_csamul_cla32_fa15_25_and0 | s_csamul_cla32_fa15_25_and1;
  assign s_csamul_cla32_and16_25 = a[16] & b[25];
  assign s_csamul_cla32_fa16_25_xor0 = s_csamul_cla32_and16_25 ^ s_csamul_cla32_fa17_24_xor1;
  assign s_csamul_cla32_fa16_25_and0 = s_csamul_cla32_and16_25 & s_csamul_cla32_fa17_24_xor1;
  assign s_csamul_cla32_fa16_25_xor1 = s_csamul_cla32_fa16_25_xor0 ^ s_csamul_cla32_fa16_24_or0;
  assign s_csamul_cla32_fa16_25_and1 = s_csamul_cla32_fa16_25_xor0 & s_csamul_cla32_fa16_24_or0;
  assign s_csamul_cla32_fa16_25_or0 = s_csamul_cla32_fa16_25_and0 | s_csamul_cla32_fa16_25_and1;
  assign s_csamul_cla32_and17_25 = a[17] & b[25];
  assign s_csamul_cla32_fa17_25_xor0 = s_csamul_cla32_and17_25 ^ s_csamul_cla32_fa18_24_xor1;
  assign s_csamul_cla32_fa17_25_and0 = s_csamul_cla32_and17_25 & s_csamul_cla32_fa18_24_xor1;
  assign s_csamul_cla32_fa17_25_xor1 = s_csamul_cla32_fa17_25_xor0 ^ s_csamul_cla32_fa17_24_or0;
  assign s_csamul_cla32_fa17_25_and1 = s_csamul_cla32_fa17_25_xor0 & s_csamul_cla32_fa17_24_or0;
  assign s_csamul_cla32_fa17_25_or0 = s_csamul_cla32_fa17_25_and0 | s_csamul_cla32_fa17_25_and1;
  assign s_csamul_cla32_and18_25 = a[18] & b[25];
  assign s_csamul_cla32_fa18_25_xor0 = s_csamul_cla32_and18_25 ^ s_csamul_cla32_fa19_24_xor1;
  assign s_csamul_cla32_fa18_25_and0 = s_csamul_cla32_and18_25 & s_csamul_cla32_fa19_24_xor1;
  assign s_csamul_cla32_fa18_25_xor1 = s_csamul_cla32_fa18_25_xor0 ^ s_csamul_cla32_fa18_24_or0;
  assign s_csamul_cla32_fa18_25_and1 = s_csamul_cla32_fa18_25_xor0 & s_csamul_cla32_fa18_24_or0;
  assign s_csamul_cla32_fa18_25_or0 = s_csamul_cla32_fa18_25_and0 | s_csamul_cla32_fa18_25_and1;
  assign s_csamul_cla32_and19_25 = a[19] & b[25];
  assign s_csamul_cla32_fa19_25_xor0 = s_csamul_cla32_and19_25 ^ s_csamul_cla32_fa20_24_xor1;
  assign s_csamul_cla32_fa19_25_and0 = s_csamul_cla32_and19_25 & s_csamul_cla32_fa20_24_xor1;
  assign s_csamul_cla32_fa19_25_xor1 = s_csamul_cla32_fa19_25_xor0 ^ s_csamul_cla32_fa19_24_or0;
  assign s_csamul_cla32_fa19_25_and1 = s_csamul_cla32_fa19_25_xor0 & s_csamul_cla32_fa19_24_or0;
  assign s_csamul_cla32_fa19_25_or0 = s_csamul_cla32_fa19_25_and0 | s_csamul_cla32_fa19_25_and1;
  assign s_csamul_cla32_and20_25 = a[20] & b[25];
  assign s_csamul_cla32_fa20_25_xor0 = s_csamul_cla32_and20_25 ^ s_csamul_cla32_fa21_24_xor1;
  assign s_csamul_cla32_fa20_25_and0 = s_csamul_cla32_and20_25 & s_csamul_cla32_fa21_24_xor1;
  assign s_csamul_cla32_fa20_25_xor1 = s_csamul_cla32_fa20_25_xor0 ^ s_csamul_cla32_fa20_24_or0;
  assign s_csamul_cla32_fa20_25_and1 = s_csamul_cla32_fa20_25_xor0 & s_csamul_cla32_fa20_24_or0;
  assign s_csamul_cla32_fa20_25_or0 = s_csamul_cla32_fa20_25_and0 | s_csamul_cla32_fa20_25_and1;
  assign s_csamul_cla32_and21_25 = a[21] & b[25];
  assign s_csamul_cla32_fa21_25_xor0 = s_csamul_cla32_and21_25 ^ s_csamul_cla32_fa22_24_xor1;
  assign s_csamul_cla32_fa21_25_and0 = s_csamul_cla32_and21_25 & s_csamul_cla32_fa22_24_xor1;
  assign s_csamul_cla32_fa21_25_xor1 = s_csamul_cla32_fa21_25_xor0 ^ s_csamul_cla32_fa21_24_or0;
  assign s_csamul_cla32_fa21_25_and1 = s_csamul_cla32_fa21_25_xor0 & s_csamul_cla32_fa21_24_or0;
  assign s_csamul_cla32_fa21_25_or0 = s_csamul_cla32_fa21_25_and0 | s_csamul_cla32_fa21_25_and1;
  assign s_csamul_cla32_and22_25 = a[22] & b[25];
  assign s_csamul_cla32_fa22_25_xor0 = s_csamul_cla32_and22_25 ^ s_csamul_cla32_fa23_24_xor1;
  assign s_csamul_cla32_fa22_25_and0 = s_csamul_cla32_and22_25 & s_csamul_cla32_fa23_24_xor1;
  assign s_csamul_cla32_fa22_25_xor1 = s_csamul_cla32_fa22_25_xor0 ^ s_csamul_cla32_fa22_24_or0;
  assign s_csamul_cla32_fa22_25_and1 = s_csamul_cla32_fa22_25_xor0 & s_csamul_cla32_fa22_24_or0;
  assign s_csamul_cla32_fa22_25_or0 = s_csamul_cla32_fa22_25_and0 | s_csamul_cla32_fa22_25_and1;
  assign s_csamul_cla32_and23_25 = a[23] & b[25];
  assign s_csamul_cla32_fa23_25_xor0 = s_csamul_cla32_and23_25 ^ s_csamul_cla32_fa24_24_xor1;
  assign s_csamul_cla32_fa23_25_and0 = s_csamul_cla32_and23_25 & s_csamul_cla32_fa24_24_xor1;
  assign s_csamul_cla32_fa23_25_xor1 = s_csamul_cla32_fa23_25_xor0 ^ s_csamul_cla32_fa23_24_or0;
  assign s_csamul_cla32_fa23_25_and1 = s_csamul_cla32_fa23_25_xor0 & s_csamul_cla32_fa23_24_or0;
  assign s_csamul_cla32_fa23_25_or0 = s_csamul_cla32_fa23_25_and0 | s_csamul_cla32_fa23_25_and1;
  assign s_csamul_cla32_and24_25 = a[24] & b[25];
  assign s_csamul_cla32_fa24_25_xor0 = s_csamul_cla32_and24_25 ^ s_csamul_cla32_fa25_24_xor1;
  assign s_csamul_cla32_fa24_25_and0 = s_csamul_cla32_and24_25 & s_csamul_cla32_fa25_24_xor1;
  assign s_csamul_cla32_fa24_25_xor1 = s_csamul_cla32_fa24_25_xor0 ^ s_csamul_cla32_fa24_24_or0;
  assign s_csamul_cla32_fa24_25_and1 = s_csamul_cla32_fa24_25_xor0 & s_csamul_cla32_fa24_24_or0;
  assign s_csamul_cla32_fa24_25_or0 = s_csamul_cla32_fa24_25_and0 | s_csamul_cla32_fa24_25_and1;
  assign s_csamul_cla32_and25_25 = a[25] & b[25];
  assign s_csamul_cla32_fa25_25_xor0 = s_csamul_cla32_and25_25 ^ s_csamul_cla32_fa26_24_xor1;
  assign s_csamul_cla32_fa25_25_and0 = s_csamul_cla32_and25_25 & s_csamul_cla32_fa26_24_xor1;
  assign s_csamul_cla32_fa25_25_xor1 = s_csamul_cla32_fa25_25_xor0 ^ s_csamul_cla32_fa25_24_or0;
  assign s_csamul_cla32_fa25_25_and1 = s_csamul_cla32_fa25_25_xor0 & s_csamul_cla32_fa25_24_or0;
  assign s_csamul_cla32_fa25_25_or0 = s_csamul_cla32_fa25_25_and0 | s_csamul_cla32_fa25_25_and1;
  assign s_csamul_cla32_and26_25 = a[26] & b[25];
  assign s_csamul_cla32_fa26_25_xor0 = s_csamul_cla32_and26_25 ^ s_csamul_cla32_fa27_24_xor1;
  assign s_csamul_cla32_fa26_25_and0 = s_csamul_cla32_and26_25 & s_csamul_cla32_fa27_24_xor1;
  assign s_csamul_cla32_fa26_25_xor1 = s_csamul_cla32_fa26_25_xor0 ^ s_csamul_cla32_fa26_24_or0;
  assign s_csamul_cla32_fa26_25_and1 = s_csamul_cla32_fa26_25_xor0 & s_csamul_cla32_fa26_24_or0;
  assign s_csamul_cla32_fa26_25_or0 = s_csamul_cla32_fa26_25_and0 | s_csamul_cla32_fa26_25_and1;
  assign s_csamul_cla32_and27_25 = a[27] & b[25];
  assign s_csamul_cla32_fa27_25_xor0 = s_csamul_cla32_and27_25 ^ s_csamul_cla32_fa28_24_xor1;
  assign s_csamul_cla32_fa27_25_and0 = s_csamul_cla32_and27_25 & s_csamul_cla32_fa28_24_xor1;
  assign s_csamul_cla32_fa27_25_xor1 = s_csamul_cla32_fa27_25_xor0 ^ s_csamul_cla32_fa27_24_or0;
  assign s_csamul_cla32_fa27_25_and1 = s_csamul_cla32_fa27_25_xor0 & s_csamul_cla32_fa27_24_or0;
  assign s_csamul_cla32_fa27_25_or0 = s_csamul_cla32_fa27_25_and0 | s_csamul_cla32_fa27_25_and1;
  assign s_csamul_cla32_and28_25 = a[28] & b[25];
  assign s_csamul_cla32_fa28_25_xor0 = s_csamul_cla32_and28_25 ^ s_csamul_cla32_fa29_24_xor1;
  assign s_csamul_cla32_fa28_25_and0 = s_csamul_cla32_and28_25 & s_csamul_cla32_fa29_24_xor1;
  assign s_csamul_cla32_fa28_25_xor1 = s_csamul_cla32_fa28_25_xor0 ^ s_csamul_cla32_fa28_24_or0;
  assign s_csamul_cla32_fa28_25_and1 = s_csamul_cla32_fa28_25_xor0 & s_csamul_cla32_fa28_24_or0;
  assign s_csamul_cla32_fa28_25_or0 = s_csamul_cla32_fa28_25_and0 | s_csamul_cla32_fa28_25_and1;
  assign s_csamul_cla32_and29_25 = a[29] & b[25];
  assign s_csamul_cla32_fa29_25_xor0 = s_csamul_cla32_and29_25 ^ s_csamul_cla32_fa30_24_xor1;
  assign s_csamul_cla32_fa29_25_and0 = s_csamul_cla32_and29_25 & s_csamul_cla32_fa30_24_xor1;
  assign s_csamul_cla32_fa29_25_xor1 = s_csamul_cla32_fa29_25_xor0 ^ s_csamul_cla32_fa29_24_or0;
  assign s_csamul_cla32_fa29_25_and1 = s_csamul_cla32_fa29_25_xor0 & s_csamul_cla32_fa29_24_or0;
  assign s_csamul_cla32_fa29_25_or0 = s_csamul_cla32_fa29_25_and0 | s_csamul_cla32_fa29_25_and1;
  assign s_csamul_cla32_and30_25 = a[30] & b[25];
  assign s_csamul_cla32_fa30_25_xor0 = s_csamul_cla32_and30_25 ^ s_csamul_cla32_ha31_24_xor0;
  assign s_csamul_cla32_fa30_25_and0 = s_csamul_cla32_and30_25 & s_csamul_cla32_ha31_24_xor0;
  assign s_csamul_cla32_fa30_25_xor1 = s_csamul_cla32_fa30_25_xor0 ^ s_csamul_cla32_fa30_24_or0;
  assign s_csamul_cla32_fa30_25_and1 = s_csamul_cla32_fa30_25_xor0 & s_csamul_cla32_fa30_24_or0;
  assign s_csamul_cla32_fa30_25_or0 = s_csamul_cla32_fa30_25_and0 | s_csamul_cla32_fa30_25_and1;
  assign s_csamul_cla32_nand31_25 = ~(a[31] & b[25]);
  assign s_csamul_cla32_ha31_25_xor0 = s_csamul_cla32_nand31_25 ^ s_csamul_cla32_ha31_24_and0;
  assign s_csamul_cla32_ha31_25_and0 = s_csamul_cla32_nand31_25 & s_csamul_cla32_ha31_24_and0;
  assign s_csamul_cla32_and0_26 = a[0] & b[26];
  assign s_csamul_cla32_fa0_26_xor0 = s_csamul_cla32_and0_26 ^ s_csamul_cla32_fa1_25_xor1;
  assign s_csamul_cla32_fa0_26_and0 = s_csamul_cla32_and0_26 & s_csamul_cla32_fa1_25_xor1;
  assign s_csamul_cla32_fa0_26_xor1 = s_csamul_cla32_fa0_26_xor0 ^ s_csamul_cla32_fa0_25_or0;
  assign s_csamul_cla32_fa0_26_and1 = s_csamul_cla32_fa0_26_xor0 & s_csamul_cla32_fa0_25_or0;
  assign s_csamul_cla32_fa0_26_or0 = s_csamul_cla32_fa0_26_and0 | s_csamul_cla32_fa0_26_and1;
  assign s_csamul_cla32_and1_26 = a[1] & b[26];
  assign s_csamul_cla32_fa1_26_xor0 = s_csamul_cla32_and1_26 ^ s_csamul_cla32_fa2_25_xor1;
  assign s_csamul_cla32_fa1_26_and0 = s_csamul_cla32_and1_26 & s_csamul_cla32_fa2_25_xor1;
  assign s_csamul_cla32_fa1_26_xor1 = s_csamul_cla32_fa1_26_xor0 ^ s_csamul_cla32_fa1_25_or0;
  assign s_csamul_cla32_fa1_26_and1 = s_csamul_cla32_fa1_26_xor0 & s_csamul_cla32_fa1_25_or0;
  assign s_csamul_cla32_fa1_26_or0 = s_csamul_cla32_fa1_26_and0 | s_csamul_cla32_fa1_26_and1;
  assign s_csamul_cla32_and2_26 = a[2] & b[26];
  assign s_csamul_cla32_fa2_26_xor0 = s_csamul_cla32_and2_26 ^ s_csamul_cla32_fa3_25_xor1;
  assign s_csamul_cla32_fa2_26_and0 = s_csamul_cla32_and2_26 & s_csamul_cla32_fa3_25_xor1;
  assign s_csamul_cla32_fa2_26_xor1 = s_csamul_cla32_fa2_26_xor0 ^ s_csamul_cla32_fa2_25_or0;
  assign s_csamul_cla32_fa2_26_and1 = s_csamul_cla32_fa2_26_xor0 & s_csamul_cla32_fa2_25_or0;
  assign s_csamul_cla32_fa2_26_or0 = s_csamul_cla32_fa2_26_and0 | s_csamul_cla32_fa2_26_and1;
  assign s_csamul_cla32_and3_26 = a[3] & b[26];
  assign s_csamul_cla32_fa3_26_xor0 = s_csamul_cla32_and3_26 ^ s_csamul_cla32_fa4_25_xor1;
  assign s_csamul_cla32_fa3_26_and0 = s_csamul_cla32_and3_26 & s_csamul_cla32_fa4_25_xor1;
  assign s_csamul_cla32_fa3_26_xor1 = s_csamul_cla32_fa3_26_xor0 ^ s_csamul_cla32_fa3_25_or0;
  assign s_csamul_cla32_fa3_26_and1 = s_csamul_cla32_fa3_26_xor0 & s_csamul_cla32_fa3_25_or0;
  assign s_csamul_cla32_fa3_26_or0 = s_csamul_cla32_fa3_26_and0 | s_csamul_cla32_fa3_26_and1;
  assign s_csamul_cla32_and4_26 = a[4] & b[26];
  assign s_csamul_cla32_fa4_26_xor0 = s_csamul_cla32_and4_26 ^ s_csamul_cla32_fa5_25_xor1;
  assign s_csamul_cla32_fa4_26_and0 = s_csamul_cla32_and4_26 & s_csamul_cla32_fa5_25_xor1;
  assign s_csamul_cla32_fa4_26_xor1 = s_csamul_cla32_fa4_26_xor0 ^ s_csamul_cla32_fa4_25_or0;
  assign s_csamul_cla32_fa4_26_and1 = s_csamul_cla32_fa4_26_xor0 & s_csamul_cla32_fa4_25_or0;
  assign s_csamul_cla32_fa4_26_or0 = s_csamul_cla32_fa4_26_and0 | s_csamul_cla32_fa4_26_and1;
  assign s_csamul_cla32_and5_26 = a[5] & b[26];
  assign s_csamul_cla32_fa5_26_xor0 = s_csamul_cla32_and5_26 ^ s_csamul_cla32_fa6_25_xor1;
  assign s_csamul_cla32_fa5_26_and0 = s_csamul_cla32_and5_26 & s_csamul_cla32_fa6_25_xor1;
  assign s_csamul_cla32_fa5_26_xor1 = s_csamul_cla32_fa5_26_xor0 ^ s_csamul_cla32_fa5_25_or0;
  assign s_csamul_cla32_fa5_26_and1 = s_csamul_cla32_fa5_26_xor0 & s_csamul_cla32_fa5_25_or0;
  assign s_csamul_cla32_fa5_26_or0 = s_csamul_cla32_fa5_26_and0 | s_csamul_cla32_fa5_26_and1;
  assign s_csamul_cla32_and6_26 = a[6] & b[26];
  assign s_csamul_cla32_fa6_26_xor0 = s_csamul_cla32_and6_26 ^ s_csamul_cla32_fa7_25_xor1;
  assign s_csamul_cla32_fa6_26_and0 = s_csamul_cla32_and6_26 & s_csamul_cla32_fa7_25_xor1;
  assign s_csamul_cla32_fa6_26_xor1 = s_csamul_cla32_fa6_26_xor0 ^ s_csamul_cla32_fa6_25_or0;
  assign s_csamul_cla32_fa6_26_and1 = s_csamul_cla32_fa6_26_xor0 & s_csamul_cla32_fa6_25_or0;
  assign s_csamul_cla32_fa6_26_or0 = s_csamul_cla32_fa6_26_and0 | s_csamul_cla32_fa6_26_and1;
  assign s_csamul_cla32_and7_26 = a[7] & b[26];
  assign s_csamul_cla32_fa7_26_xor0 = s_csamul_cla32_and7_26 ^ s_csamul_cla32_fa8_25_xor1;
  assign s_csamul_cla32_fa7_26_and0 = s_csamul_cla32_and7_26 & s_csamul_cla32_fa8_25_xor1;
  assign s_csamul_cla32_fa7_26_xor1 = s_csamul_cla32_fa7_26_xor0 ^ s_csamul_cla32_fa7_25_or0;
  assign s_csamul_cla32_fa7_26_and1 = s_csamul_cla32_fa7_26_xor0 & s_csamul_cla32_fa7_25_or0;
  assign s_csamul_cla32_fa7_26_or0 = s_csamul_cla32_fa7_26_and0 | s_csamul_cla32_fa7_26_and1;
  assign s_csamul_cla32_and8_26 = a[8] & b[26];
  assign s_csamul_cla32_fa8_26_xor0 = s_csamul_cla32_and8_26 ^ s_csamul_cla32_fa9_25_xor1;
  assign s_csamul_cla32_fa8_26_and0 = s_csamul_cla32_and8_26 & s_csamul_cla32_fa9_25_xor1;
  assign s_csamul_cla32_fa8_26_xor1 = s_csamul_cla32_fa8_26_xor0 ^ s_csamul_cla32_fa8_25_or0;
  assign s_csamul_cla32_fa8_26_and1 = s_csamul_cla32_fa8_26_xor0 & s_csamul_cla32_fa8_25_or0;
  assign s_csamul_cla32_fa8_26_or0 = s_csamul_cla32_fa8_26_and0 | s_csamul_cla32_fa8_26_and1;
  assign s_csamul_cla32_and9_26 = a[9] & b[26];
  assign s_csamul_cla32_fa9_26_xor0 = s_csamul_cla32_and9_26 ^ s_csamul_cla32_fa10_25_xor1;
  assign s_csamul_cla32_fa9_26_and0 = s_csamul_cla32_and9_26 & s_csamul_cla32_fa10_25_xor1;
  assign s_csamul_cla32_fa9_26_xor1 = s_csamul_cla32_fa9_26_xor0 ^ s_csamul_cla32_fa9_25_or0;
  assign s_csamul_cla32_fa9_26_and1 = s_csamul_cla32_fa9_26_xor0 & s_csamul_cla32_fa9_25_or0;
  assign s_csamul_cla32_fa9_26_or0 = s_csamul_cla32_fa9_26_and0 | s_csamul_cla32_fa9_26_and1;
  assign s_csamul_cla32_and10_26 = a[10] & b[26];
  assign s_csamul_cla32_fa10_26_xor0 = s_csamul_cla32_and10_26 ^ s_csamul_cla32_fa11_25_xor1;
  assign s_csamul_cla32_fa10_26_and0 = s_csamul_cla32_and10_26 & s_csamul_cla32_fa11_25_xor1;
  assign s_csamul_cla32_fa10_26_xor1 = s_csamul_cla32_fa10_26_xor0 ^ s_csamul_cla32_fa10_25_or0;
  assign s_csamul_cla32_fa10_26_and1 = s_csamul_cla32_fa10_26_xor0 & s_csamul_cla32_fa10_25_or0;
  assign s_csamul_cla32_fa10_26_or0 = s_csamul_cla32_fa10_26_and0 | s_csamul_cla32_fa10_26_and1;
  assign s_csamul_cla32_and11_26 = a[11] & b[26];
  assign s_csamul_cla32_fa11_26_xor0 = s_csamul_cla32_and11_26 ^ s_csamul_cla32_fa12_25_xor1;
  assign s_csamul_cla32_fa11_26_and0 = s_csamul_cla32_and11_26 & s_csamul_cla32_fa12_25_xor1;
  assign s_csamul_cla32_fa11_26_xor1 = s_csamul_cla32_fa11_26_xor0 ^ s_csamul_cla32_fa11_25_or0;
  assign s_csamul_cla32_fa11_26_and1 = s_csamul_cla32_fa11_26_xor0 & s_csamul_cla32_fa11_25_or0;
  assign s_csamul_cla32_fa11_26_or0 = s_csamul_cla32_fa11_26_and0 | s_csamul_cla32_fa11_26_and1;
  assign s_csamul_cla32_and12_26 = a[12] & b[26];
  assign s_csamul_cla32_fa12_26_xor0 = s_csamul_cla32_and12_26 ^ s_csamul_cla32_fa13_25_xor1;
  assign s_csamul_cla32_fa12_26_and0 = s_csamul_cla32_and12_26 & s_csamul_cla32_fa13_25_xor1;
  assign s_csamul_cla32_fa12_26_xor1 = s_csamul_cla32_fa12_26_xor0 ^ s_csamul_cla32_fa12_25_or0;
  assign s_csamul_cla32_fa12_26_and1 = s_csamul_cla32_fa12_26_xor0 & s_csamul_cla32_fa12_25_or0;
  assign s_csamul_cla32_fa12_26_or0 = s_csamul_cla32_fa12_26_and0 | s_csamul_cla32_fa12_26_and1;
  assign s_csamul_cla32_and13_26 = a[13] & b[26];
  assign s_csamul_cla32_fa13_26_xor0 = s_csamul_cla32_and13_26 ^ s_csamul_cla32_fa14_25_xor1;
  assign s_csamul_cla32_fa13_26_and0 = s_csamul_cla32_and13_26 & s_csamul_cla32_fa14_25_xor1;
  assign s_csamul_cla32_fa13_26_xor1 = s_csamul_cla32_fa13_26_xor0 ^ s_csamul_cla32_fa13_25_or0;
  assign s_csamul_cla32_fa13_26_and1 = s_csamul_cla32_fa13_26_xor0 & s_csamul_cla32_fa13_25_or0;
  assign s_csamul_cla32_fa13_26_or0 = s_csamul_cla32_fa13_26_and0 | s_csamul_cla32_fa13_26_and1;
  assign s_csamul_cla32_and14_26 = a[14] & b[26];
  assign s_csamul_cla32_fa14_26_xor0 = s_csamul_cla32_and14_26 ^ s_csamul_cla32_fa15_25_xor1;
  assign s_csamul_cla32_fa14_26_and0 = s_csamul_cla32_and14_26 & s_csamul_cla32_fa15_25_xor1;
  assign s_csamul_cla32_fa14_26_xor1 = s_csamul_cla32_fa14_26_xor0 ^ s_csamul_cla32_fa14_25_or0;
  assign s_csamul_cla32_fa14_26_and1 = s_csamul_cla32_fa14_26_xor0 & s_csamul_cla32_fa14_25_or0;
  assign s_csamul_cla32_fa14_26_or0 = s_csamul_cla32_fa14_26_and0 | s_csamul_cla32_fa14_26_and1;
  assign s_csamul_cla32_and15_26 = a[15] & b[26];
  assign s_csamul_cla32_fa15_26_xor0 = s_csamul_cla32_and15_26 ^ s_csamul_cla32_fa16_25_xor1;
  assign s_csamul_cla32_fa15_26_and0 = s_csamul_cla32_and15_26 & s_csamul_cla32_fa16_25_xor1;
  assign s_csamul_cla32_fa15_26_xor1 = s_csamul_cla32_fa15_26_xor0 ^ s_csamul_cla32_fa15_25_or0;
  assign s_csamul_cla32_fa15_26_and1 = s_csamul_cla32_fa15_26_xor0 & s_csamul_cla32_fa15_25_or0;
  assign s_csamul_cla32_fa15_26_or0 = s_csamul_cla32_fa15_26_and0 | s_csamul_cla32_fa15_26_and1;
  assign s_csamul_cla32_and16_26 = a[16] & b[26];
  assign s_csamul_cla32_fa16_26_xor0 = s_csamul_cla32_and16_26 ^ s_csamul_cla32_fa17_25_xor1;
  assign s_csamul_cla32_fa16_26_and0 = s_csamul_cla32_and16_26 & s_csamul_cla32_fa17_25_xor1;
  assign s_csamul_cla32_fa16_26_xor1 = s_csamul_cla32_fa16_26_xor0 ^ s_csamul_cla32_fa16_25_or0;
  assign s_csamul_cla32_fa16_26_and1 = s_csamul_cla32_fa16_26_xor0 & s_csamul_cla32_fa16_25_or0;
  assign s_csamul_cla32_fa16_26_or0 = s_csamul_cla32_fa16_26_and0 | s_csamul_cla32_fa16_26_and1;
  assign s_csamul_cla32_and17_26 = a[17] & b[26];
  assign s_csamul_cla32_fa17_26_xor0 = s_csamul_cla32_and17_26 ^ s_csamul_cla32_fa18_25_xor1;
  assign s_csamul_cla32_fa17_26_and0 = s_csamul_cla32_and17_26 & s_csamul_cla32_fa18_25_xor1;
  assign s_csamul_cla32_fa17_26_xor1 = s_csamul_cla32_fa17_26_xor0 ^ s_csamul_cla32_fa17_25_or0;
  assign s_csamul_cla32_fa17_26_and1 = s_csamul_cla32_fa17_26_xor0 & s_csamul_cla32_fa17_25_or0;
  assign s_csamul_cla32_fa17_26_or0 = s_csamul_cla32_fa17_26_and0 | s_csamul_cla32_fa17_26_and1;
  assign s_csamul_cla32_and18_26 = a[18] & b[26];
  assign s_csamul_cla32_fa18_26_xor0 = s_csamul_cla32_and18_26 ^ s_csamul_cla32_fa19_25_xor1;
  assign s_csamul_cla32_fa18_26_and0 = s_csamul_cla32_and18_26 & s_csamul_cla32_fa19_25_xor1;
  assign s_csamul_cla32_fa18_26_xor1 = s_csamul_cla32_fa18_26_xor0 ^ s_csamul_cla32_fa18_25_or0;
  assign s_csamul_cla32_fa18_26_and1 = s_csamul_cla32_fa18_26_xor0 & s_csamul_cla32_fa18_25_or0;
  assign s_csamul_cla32_fa18_26_or0 = s_csamul_cla32_fa18_26_and0 | s_csamul_cla32_fa18_26_and1;
  assign s_csamul_cla32_and19_26 = a[19] & b[26];
  assign s_csamul_cla32_fa19_26_xor0 = s_csamul_cla32_and19_26 ^ s_csamul_cla32_fa20_25_xor1;
  assign s_csamul_cla32_fa19_26_and0 = s_csamul_cla32_and19_26 & s_csamul_cla32_fa20_25_xor1;
  assign s_csamul_cla32_fa19_26_xor1 = s_csamul_cla32_fa19_26_xor0 ^ s_csamul_cla32_fa19_25_or0;
  assign s_csamul_cla32_fa19_26_and1 = s_csamul_cla32_fa19_26_xor0 & s_csamul_cla32_fa19_25_or0;
  assign s_csamul_cla32_fa19_26_or0 = s_csamul_cla32_fa19_26_and0 | s_csamul_cla32_fa19_26_and1;
  assign s_csamul_cla32_and20_26 = a[20] & b[26];
  assign s_csamul_cla32_fa20_26_xor0 = s_csamul_cla32_and20_26 ^ s_csamul_cla32_fa21_25_xor1;
  assign s_csamul_cla32_fa20_26_and0 = s_csamul_cla32_and20_26 & s_csamul_cla32_fa21_25_xor1;
  assign s_csamul_cla32_fa20_26_xor1 = s_csamul_cla32_fa20_26_xor0 ^ s_csamul_cla32_fa20_25_or0;
  assign s_csamul_cla32_fa20_26_and1 = s_csamul_cla32_fa20_26_xor0 & s_csamul_cla32_fa20_25_or0;
  assign s_csamul_cla32_fa20_26_or0 = s_csamul_cla32_fa20_26_and0 | s_csamul_cla32_fa20_26_and1;
  assign s_csamul_cla32_and21_26 = a[21] & b[26];
  assign s_csamul_cla32_fa21_26_xor0 = s_csamul_cla32_and21_26 ^ s_csamul_cla32_fa22_25_xor1;
  assign s_csamul_cla32_fa21_26_and0 = s_csamul_cla32_and21_26 & s_csamul_cla32_fa22_25_xor1;
  assign s_csamul_cla32_fa21_26_xor1 = s_csamul_cla32_fa21_26_xor0 ^ s_csamul_cla32_fa21_25_or0;
  assign s_csamul_cla32_fa21_26_and1 = s_csamul_cla32_fa21_26_xor0 & s_csamul_cla32_fa21_25_or0;
  assign s_csamul_cla32_fa21_26_or0 = s_csamul_cla32_fa21_26_and0 | s_csamul_cla32_fa21_26_and1;
  assign s_csamul_cla32_and22_26 = a[22] & b[26];
  assign s_csamul_cla32_fa22_26_xor0 = s_csamul_cla32_and22_26 ^ s_csamul_cla32_fa23_25_xor1;
  assign s_csamul_cla32_fa22_26_and0 = s_csamul_cla32_and22_26 & s_csamul_cla32_fa23_25_xor1;
  assign s_csamul_cla32_fa22_26_xor1 = s_csamul_cla32_fa22_26_xor0 ^ s_csamul_cla32_fa22_25_or0;
  assign s_csamul_cla32_fa22_26_and1 = s_csamul_cla32_fa22_26_xor0 & s_csamul_cla32_fa22_25_or0;
  assign s_csamul_cla32_fa22_26_or0 = s_csamul_cla32_fa22_26_and0 | s_csamul_cla32_fa22_26_and1;
  assign s_csamul_cla32_and23_26 = a[23] & b[26];
  assign s_csamul_cla32_fa23_26_xor0 = s_csamul_cla32_and23_26 ^ s_csamul_cla32_fa24_25_xor1;
  assign s_csamul_cla32_fa23_26_and0 = s_csamul_cla32_and23_26 & s_csamul_cla32_fa24_25_xor1;
  assign s_csamul_cla32_fa23_26_xor1 = s_csamul_cla32_fa23_26_xor0 ^ s_csamul_cla32_fa23_25_or0;
  assign s_csamul_cla32_fa23_26_and1 = s_csamul_cla32_fa23_26_xor0 & s_csamul_cla32_fa23_25_or0;
  assign s_csamul_cla32_fa23_26_or0 = s_csamul_cla32_fa23_26_and0 | s_csamul_cla32_fa23_26_and1;
  assign s_csamul_cla32_and24_26 = a[24] & b[26];
  assign s_csamul_cla32_fa24_26_xor0 = s_csamul_cla32_and24_26 ^ s_csamul_cla32_fa25_25_xor1;
  assign s_csamul_cla32_fa24_26_and0 = s_csamul_cla32_and24_26 & s_csamul_cla32_fa25_25_xor1;
  assign s_csamul_cla32_fa24_26_xor1 = s_csamul_cla32_fa24_26_xor0 ^ s_csamul_cla32_fa24_25_or0;
  assign s_csamul_cla32_fa24_26_and1 = s_csamul_cla32_fa24_26_xor0 & s_csamul_cla32_fa24_25_or0;
  assign s_csamul_cla32_fa24_26_or0 = s_csamul_cla32_fa24_26_and0 | s_csamul_cla32_fa24_26_and1;
  assign s_csamul_cla32_and25_26 = a[25] & b[26];
  assign s_csamul_cla32_fa25_26_xor0 = s_csamul_cla32_and25_26 ^ s_csamul_cla32_fa26_25_xor1;
  assign s_csamul_cla32_fa25_26_and0 = s_csamul_cla32_and25_26 & s_csamul_cla32_fa26_25_xor1;
  assign s_csamul_cla32_fa25_26_xor1 = s_csamul_cla32_fa25_26_xor0 ^ s_csamul_cla32_fa25_25_or0;
  assign s_csamul_cla32_fa25_26_and1 = s_csamul_cla32_fa25_26_xor0 & s_csamul_cla32_fa25_25_or0;
  assign s_csamul_cla32_fa25_26_or0 = s_csamul_cla32_fa25_26_and0 | s_csamul_cla32_fa25_26_and1;
  assign s_csamul_cla32_and26_26 = a[26] & b[26];
  assign s_csamul_cla32_fa26_26_xor0 = s_csamul_cla32_and26_26 ^ s_csamul_cla32_fa27_25_xor1;
  assign s_csamul_cla32_fa26_26_and0 = s_csamul_cla32_and26_26 & s_csamul_cla32_fa27_25_xor1;
  assign s_csamul_cla32_fa26_26_xor1 = s_csamul_cla32_fa26_26_xor0 ^ s_csamul_cla32_fa26_25_or0;
  assign s_csamul_cla32_fa26_26_and1 = s_csamul_cla32_fa26_26_xor0 & s_csamul_cla32_fa26_25_or0;
  assign s_csamul_cla32_fa26_26_or0 = s_csamul_cla32_fa26_26_and0 | s_csamul_cla32_fa26_26_and1;
  assign s_csamul_cla32_and27_26 = a[27] & b[26];
  assign s_csamul_cla32_fa27_26_xor0 = s_csamul_cla32_and27_26 ^ s_csamul_cla32_fa28_25_xor1;
  assign s_csamul_cla32_fa27_26_and0 = s_csamul_cla32_and27_26 & s_csamul_cla32_fa28_25_xor1;
  assign s_csamul_cla32_fa27_26_xor1 = s_csamul_cla32_fa27_26_xor0 ^ s_csamul_cla32_fa27_25_or0;
  assign s_csamul_cla32_fa27_26_and1 = s_csamul_cla32_fa27_26_xor0 & s_csamul_cla32_fa27_25_or0;
  assign s_csamul_cla32_fa27_26_or0 = s_csamul_cla32_fa27_26_and0 | s_csamul_cla32_fa27_26_and1;
  assign s_csamul_cla32_and28_26 = a[28] & b[26];
  assign s_csamul_cla32_fa28_26_xor0 = s_csamul_cla32_and28_26 ^ s_csamul_cla32_fa29_25_xor1;
  assign s_csamul_cla32_fa28_26_and0 = s_csamul_cla32_and28_26 & s_csamul_cla32_fa29_25_xor1;
  assign s_csamul_cla32_fa28_26_xor1 = s_csamul_cla32_fa28_26_xor0 ^ s_csamul_cla32_fa28_25_or0;
  assign s_csamul_cla32_fa28_26_and1 = s_csamul_cla32_fa28_26_xor0 & s_csamul_cla32_fa28_25_or0;
  assign s_csamul_cla32_fa28_26_or0 = s_csamul_cla32_fa28_26_and0 | s_csamul_cla32_fa28_26_and1;
  assign s_csamul_cla32_and29_26 = a[29] & b[26];
  assign s_csamul_cla32_fa29_26_xor0 = s_csamul_cla32_and29_26 ^ s_csamul_cla32_fa30_25_xor1;
  assign s_csamul_cla32_fa29_26_and0 = s_csamul_cla32_and29_26 & s_csamul_cla32_fa30_25_xor1;
  assign s_csamul_cla32_fa29_26_xor1 = s_csamul_cla32_fa29_26_xor0 ^ s_csamul_cla32_fa29_25_or0;
  assign s_csamul_cla32_fa29_26_and1 = s_csamul_cla32_fa29_26_xor0 & s_csamul_cla32_fa29_25_or0;
  assign s_csamul_cla32_fa29_26_or0 = s_csamul_cla32_fa29_26_and0 | s_csamul_cla32_fa29_26_and1;
  assign s_csamul_cla32_and30_26 = a[30] & b[26];
  assign s_csamul_cla32_fa30_26_xor0 = s_csamul_cla32_and30_26 ^ s_csamul_cla32_ha31_25_xor0;
  assign s_csamul_cla32_fa30_26_and0 = s_csamul_cla32_and30_26 & s_csamul_cla32_ha31_25_xor0;
  assign s_csamul_cla32_fa30_26_xor1 = s_csamul_cla32_fa30_26_xor0 ^ s_csamul_cla32_fa30_25_or0;
  assign s_csamul_cla32_fa30_26_and1 = s_csamul_cla32_fa30_26_xor0 & s_csamul_cla32_fa30_25_or0;
  assign s_csamul_cla32_fa30_26_or0 = s_csamul_cla32_fa30_26_and0 | s_csamul_cla32_fa30_26_and1;
  assign s_csamul_cla32_nand31_26 = ~(a[31] & b[26]);
  assign s_csamul_cla32_ha31_26_xor0 = s_csamul_cla32_nand31_26 ^ s_csamul_cla32_ha31_25_and0;
  assign s_csamul_cla32_ha31_26_and0 = s_csamul_cla32_nand31_26 & s_csamul_cla32_ha31_25_and0;
  assign s_csamul_cla32_and0_27 = a[0] & b[27];
  assign s_csamul_cla32_fa0_27_xor0 = s_csamul_cla32_and0_27 ^ s_csamul_cla32_fa1_26_xor1;
  assign s_csamul_cla32_fa0_27_and0 = s_csamul_cla32_and0_27 & s_csamul_cla32_fa1_26_xor1;
  assign s_csamul_cla32_fa0_27_xor1 = s_csamul_cla32_fa0_27_xor0 ^ s_csamul_cla32_fa0_26_or0;
  assign s_csamul_cla32_fa0_27_and1 = s_csamul_cla32_fa0_27_xor0 & s_csamul_cla32_fa0_26_or0;
  assign s_csamul_cla32_fa0_27_or0 = s_csamul_cla32_fa0_27_and0 | s_csamul_cla32_fa0_27_and1;
  assign s_csamul_cla32_and1_27 = a[1] & b[27];
  assign s_csamul_cla32_fa1_27_xor0 = s_csamul_cla32_and1_27 ^ s_csamul_cla32_fa2_26_xor1;
  assign s_csamul_cla32_fa1_27_and0 = s_csamul_cla32_and1_27 & s_csamul_cla32_fa2_26_xor1;
  assign s_csamul_cla32_fa1_27_xor1 = s_csamul_cla32_fa1_27_xor0 ^ s_csamul_cla32_fa1_26_or0;
  assign s_csamul_cla32_fa1_27_and1 = s_csamul_cla32_fa1_27_xor0 & s_csamul_cla32_fa1_26_or0;
  assign s_csamul_cla32_fa1_27_or0 = s_csamul_cla32_fa1_27_and0 | s_csamul_cla32_fa1_27_and1;
  assign s_csamul_cla32_and2_27 = a[2] & b[27];
  assign s_csamul_cla32_fa2_27_xor0 = s_csamul_cla32_and2_27 ^ s_csamul_cla32_fa3_26_xor1;
  assign s_csamul_cla32_fa2_27_and0 = s_csamul_cla32_and2_27 & s_csamul_cla32_fa3_26_xor1;
  assign s_csamul_cla32_fa2_27_xor1 = s_csamul_cla32_fa2_27_xor0 ^ s_csamul_cla32_fa2_26_or0;
  assign s_csamul_cla32_fa2_27_and1 = s_csamul_cla32_fa2_27_xor0 & s_csamul_cla32_fa2_26_or0;
  assign s_csamul_cla32_fa2_27_or0 = s_csamul_cla32_fa2_27_and0 | s_csamul_cla32_fa2_27_and1;
  assign s_csamul_cla32_and3_27 = a[3] & b[27];
  assign s_csamul_cla32_fa3_27_xor0 = s_csamul_cla32_and3_27 ^ s_csamul_cla32_fa4_26_xor1;
  assign s_csamul_cla32_fa3_27_and0 = s_csamul_cla32_and3_27 & s_csamul_cla32_fa4_26_xor1;
  assign s_csamul_cla32_fa3_27_xor1 = s_csamul_cla32_fa3_27_xor0 ^ s_csamul_cla32_fa3_26_or0;
  assign s_csamul_cla32_fa3_27_and1 = s_csamul_cla32_fa3_27_xor0 & s_csamul_cla32_fa3_26_or0;
  assign s_csamul_cla32_fa3_27_or0 = s_csamul_cla32_fa3_27_and0 | s_csamul_cla32_fa3_27_and1;
  assign s_csamul_cla32_and4_27 = a[4] & b[27];
  assign s_csamul_cla32_fa4_27_xor0 = s_csamul_cla32_and4_27 ^ s_csamul_cla32_fa5_26_xor1;
  assign s_csamul_cla32_fa4_27_and0 = s_csamul_cla32_and4_27 & s_csamul_cla32_fa5_26_xor1;
  assign s_csamul_cla32_fa4_27_xor1 = s_csamul_cla32_fa4_27_xor0 ^ s_csamul_cla32_fa4_26_or0;
  assign s_csamul_cla32_fa4_27_and1 = s_csamul_cla32_fa4_27_xor0 & s_csamul_cla32_fa4_26_or0;
  assign s_csamul_cla32_fa4_27_or0 = s_csamul_cla32_fa4_27_and0 | s_csamul_cla32_fa4_27_and1;
  assign s_csamul_cla32_and5_27 = a[5] & b[27];
  assign s_csamul_cla32_fa5_27_xor0 = s_csamul_cla32_and5_27 ^ s_csamul_cla32_fa6_26_xor1;
  assign s_csamul_cla32_fa5_27_and0 = s_csamul_cla32_and5_27 & s_csamul_cla32_fa6_26_xor1;
  assign s_csamul_cla32_fa5_27_xor1 = s_csamul_cla32_fa5_27_xor0 ^ s_csamul_cla32_fa5_26_or0;
  assign s_csamul_cla32_fa5_27_and1 = s_csamul_cla32_fa5_27_xor0 & s_csamul_cla32_fa5_26_or0;
  assign s_csamul_cla32_fa5_27_or0 = s_csamul_cla32_fa5_27_and0 | s_csamul_cla32_fa5_27_and1;
  assign s_csamul_cla32_and6_27 = a[6] & b[27];
  assign s_csamul_cla32_fa6_27_xor0 = s_csamul_cla32_and6_27 ^ s_csamul_cla32_fa7_26_xor1;
  assign s_csamul_cla32_fa6_27_and0 = s_csamul_cla32_and6_27 & s_csamul_cla32_fa7_26_xor1;
  assign s_csamul_cla32_fa6_27_xor1 = s_csamul_cla32_fa6_27_xor0 ^ s_csamul_cla32_fa6_26_or0;
  assign s_csamul_cla32_fa6_27_and1 = s_csamul_cla32_fa6_27_xor0 & s_csamul_cla32_fa6_26_or0;
  assign s_csamul_cla32_fa6_27_or0 = s_csamul_cla32_fa6_27_and0 | s_csamul_cla32_fa6_27_and1;
  assign s_csamul_cla32_and7_27 = a[7] & b[27];
  assign s_csamul_cla32_fa7_27_xor0 = s_csamul_cla32_and7_27 ^ s_csamul_cla32_fa8_26_xor1;
  assign s_csamul_cla32_fa7_27_and0 = s_csamul_cla32_and7_27 & s_csamul_cla32_fa8_26_xor1;
  assign s_csamul_cla32_fa7_27_xor1 = s_csamul_cla32_fa7_27_xor0 ^ s_csamul_cla32_fa7_26_or0;
  assign s_csamul_cla32_fa7_27_and1 = s_csamul_cla32_fa7_27_xor0 & s_csamul_cla32_fa7_26_or0;
  assign s_csamul_cla32_fa7_27_or0 = s_csamul_cla32_fa7_27_and0 | s_csamul_cla32_fa7_27_and1;
  assign s_csamul_cla32_and8_27 = a[8] & b[27];
  assign s_csamul_cla32_fa8_27_xor0 = s_csamul_cla32_and8_27 ^ s_csamul_cla32_fa9_26_xor1;
  assign s_csamul_cla32_fa8_27_and0 = s_csamul_cla32_and8_27 & s_csamul_cla32_fa9_26_xor1;
  assign s_csamul_cla32_fa8_27_xor1 = s_csamul_cla32_fa8_27_xor0 ^ s_csamul_cla32_fa8_26_or0;
  assign s_csamul_cla32_fa8_27_and1 = s_csamul_cla32_fa8_27_xor0 & s_csamul_cla32_fa8_26_or0;
  assign s_csamul_cla32_fa8_27_or0 = s_csamul_cla32_fa8_27_and0 | s_csamul_cla32_fa8_27_and1;
  assign s_csamul_cla32_and9_27 = a[9] & b[27];
  assign s_csamul_cla32_fa9_27_xor0 = s_csamul_cla32_and9_27 ^ s_csamul_cla32_fa10_26_xor1;
  assign s_csamul_cla32_fa9_27_and0 = s_csamul_cla32_and9_27 & s_csamul_cla32_fa10_26_xor1;
  assign s_csamul_cla32_fa9_27_xor1 = s_csamul_cla32_fa9_27_xor0 ^ s_csamul_cla32_fa9_26_or0;
  assign s_csamul_cla32_fa9_27_and1 = s_csamul_cla32_fa9_27_xor0 & s_csamul_cla32_fa9_26_or0;
  assign s_csamul_cla32_fa9_27_or0 = s_csamul_cla32_fa9_27_and0 | s_csamul_cla32_fa9_27_and1;
  assign s_csamul_cla32_and10_27 = a[10] & b[27];
  assign s_csamul_cla32_fa10_27_xor0 = s_csamul_cla32_and10_27 ^ s_csamul_cla32_fa11_26_xor1;
  assign s_csamul_cla32_fa10_27_and0 = s_csamul_cla32_and10_27 & s_csamul_cla32_fa11_26_xor1;
  assign s_csamul_cla32_fa10_27_xor1 = s_csamul_cla32_fa10_27_xor0 ^ s_csamul_cla32_fa10_26_or0;
  assign s_csamul_cla32_fa10_27_and1 = s_csamul_cla32_fa10_27_xor0 & s_csamul_cla32_fa10_26_or0;
  assign s_csamul_cla32_fa10_27_or0 = s_csamul_cla32_fa10_27_and0 | s_csamul_cla32_fa10_27_and1;
  assign s_csamul_cla32_and11_27 = a[11] & b[27];
  assign s_csamul_cla32_fa11_27_xor0 = s_csamul_cla32_and11_27 ^ s_csamul_cla32_fa12_26_xor1;
  assign s_csamul_cla32_fa11_27_and0 = s_csamul_cla32_and11_27 & s_csamul_cla32_fa12_26_xor1;
  assign s_csamul_cla32_fa11_27_xor1 = s_csamul_cla32_fa11_27_xor0 ^ s_csamul_cla32_fa11_26_or0;
  assign s_csamul_cla32_fa11_27_and1 = s_csamul_cla32_fa11_27_xor0 & s_csamul_cla32_fa11_26_or0;
  assign s_csamul_cla32_fa11_27_or0 = s_csamul_cla32_fa11_27_and0 | s_csamul_cla32_fa11_27_and1;
  assign s_csamul_cla32_and12_27 = a[12] & b[27];
  assign s_csamul_cla32_fa12_27_xor0 = s_csamul_cla32_and12_27 ^ s_csamul_cla32_fa13_26_xor1;
  assign s_csamul_cla32_fa12_27_and0 = s_csamul_cla32_and12_27 & s_csamul_cla32_fa13_26_xor1;
  assign s_csamul_cla32_fa12_27_xor1 = s_csamul_cla32_fa12_27_xor0 ^ s_csamul_cla32_fa12_26_or0;
  assign s_csamul_cla32_fa12_27_and1 = s_csamul_cla32_fa12_27_xor0 & s_csamul_cla32_fa12_26_or0;
  assign s_csamul_cla32_fa12_27_or0 = s_csamul_cla32_fa12_27_and0 | s_csamul_cla32_fa12_27_and1;
  assign s_csamul_cla32_and13_27 = a[13] & b[27];
  assign s_csamul_cla32_fa13_27_xor0 = s_csamul_cla32_and13_27 ^ s_csamul_cla32_fa14_26_xor1;
  assign s_csamul_cla32_fa13_27_and0 = s_csamul_cla32_and13_27 & s_csamul_cla32_fa14_26_xor1;
  assign s_csamul_cla32_fa13_27_xor1 = s_csamul_cla32_fa13_27_xor0 ^ s_csamul_cla32_fa13_26_or0;
  assign s_csamul_cla32_fa13_27_and1 = s_csamul_cla32_fa13_27_xor0 & s_csamul_cla32_fa13_26_or0;
  assign s_csamul_cla32_fa13_27_or0 = s_csamul_cla32_fa13_27_and0 | s_csamul_cla32_fa13_27_and1;
  assign s_csamul_cla32_and14_27 = a[14] & b[27];
  assign s_csamul_cla32_fa14_27_xor0 = s_csamul_cla32_and14_27 ^ s_csamul_cla32_fa15_26_xor1;
  assign s_csamul_cla32_fa14_27_and0 = s_csamul_cla32_and14_27 & s_csamul_cla32_fa15_26_xor1;
  assign s_csamul_cla32_fa14_27_xor1 = s_csamul_cla32_fa14_27_xor0 ^ s_csamul_cla32_fa14_26_or0;
  assign s_csamul_cla32_fa14_27_and1 = s_csamul_cla32_fa14_27_xor0 & s_csamul_cla32_fa14_26_or0;
  assign s_csamul_cla32_fa14_27_or0 = s_csamul_cla32_fa14_27_and0 | s_csamul_cla32_fa14_27_and1;
  assign s_csamul_cla32_and15_27 = a[15] & b[27];
  assign s_csamul_cla32_fa15_27_xor0 = s_csamul_cla32_and15_27 ^ s_csamul_cla32_fa16_26_xor1;
  assign s_csamul_cla32_fa15_27_and0 = s_csamul_cla32_and15_27 & s_csamul_cla32_fa16_26_xor1;
  assign s_csamul_cla32_fa15_27_xor1 = s_csamul_cla32_fa15_27_xor0 ^ s_csamul_cla32_fa15_26_or0;
  assign s_csamul_cla32_fa15_27_and1 = s_csamul_cla32_fa15_27_xor0 & s_csamul_cla32_fa15_26_or0;
  assign s_csamul_cla32_fa15_27_or0 = s_csamul_cla32_fa15_27_and0 | s_csamul_cla32_fa15_27_and1;
  assign s_csamul_cla32_and16_27 = a[16] & b[27];
  assign s_csamul_cla32_fa16_27_xor0 = s_csamul_cla32_and16_27 ^ s_csamul_cla32_fa17_26_xor1;
  assign s_csamul_cla32_fa16_27_and0 = s_csamul_cla32_and16_27 & s_csamul_cla32_fa17_26_xor1;
  assign s_csamul_cla32_fa16_27_xor1 = s_csamul_cla32_fa16_27_xor0 ^ s_csamul_cla32_fa16_26_or0;
  assign s_csamul_cla32_fa16_27_and1 = s_csamul_cla32_fa16_27_xor0 & s_csamul_cla32_fa16_26_or0;
  assign s_csamul_cla32_fa16_27_or0 = s_csamul_cla32_fa16_27_and0 | s_csamul_cla32_fa16_27_and1;
  assign s_csamul_cla32_and17_27 = a[17] & b[27];
  assign s_csamul_cla32_fa17_27_xor0 = s_csamul_cla32_and17_27 ^ s_csamul_cla32_fa18_26_xor1;
  assign s_csamul_cla32_fa17_27_and0 = s_csamul_cla32_and17_27 & s_csamul_cla32_fa18_26_xor1;
  assign s_csamul_cla32_fa17_27_xor1 = s_csamul_cla32_fa17_27_xor0 ^ s_csamul_cla32_fa17_26_or0;
  assign s_csamul_cla32_fa17_27_and1 = s_csamul_cla32_fa17_27_xor0 & s_csamul_cla32_fa17_26_or0;
  assign s_csamul_cla32_fa17_27_or0 = s_csamul_cla32_fa17_27_and0 | s_csamul_cla32_fa17_27_and1;
  assign s_csamul_cla32_and18_27 = a[18] & b[27];
  assign s_csamul_cla32_fa18_27_xor0 = s_csamul_cla32_and18_27 ^ s_csamul_cla32_fa19_26_xor1;
  assign s_csamul_cla32_fa18_27_and0 = s_csamul_cla32_and18_27 & s_csamul_cla32_fa19_26_xor1;
  assign s_csamul_cla32_fa18_27_xor1 = s_csamul_cla32_fa18_27_xor0 ^ s_csamul_cla32_fa18_26_or0;
  assign s_csamul_cla32_fa18_27_and1 = s_csamul_cla32_fa18_27_xor0 & s_csamul_cla32_fa18_26_or0;
  assign s_csamul_cla32_fa18_27_or0 = s_csamul_cla32_fa18_27_and0 | s_csamul_cla32_fa18_27_and1;
  assign s_csamul_cla32_and19_27 = a[19] & b[27];
  assign s_csamul_cla32_fa19_27_xor0 = s_csamul_cla32_and19_27 ^ s_csamul_cla32_fa20_26_xor1;
  assign s_csamul_cla32_fa19_27_and0 = s_csamul_cla32_and19_27 & s_csamul_cla32_fa20_26_xor1;
  assign s_csamul_cla32_fa19_27_xor1 = s_csamul_cla32_fa19_27_xor0 ^ s_csamul_cla32_fa19_26_or0;
  assign s_csamul_cla32_fa19_27_and1 = s_csamul_cla32_fa19_27_xor0 & s_csamul_cla32_fa19_26_or0;
  assign s_csamul_cla32_fa19_27_or0 = s_csamul_cla32_fa19_27_and0 | s_csamul_cla32_fa19_27_and1;
  assign s_csamul_cla32_and20_27 = a[20] & b[27];
  assign s_csamul_cla32_fa20_27_xor0 = s_csamul_cla32_and20_27 ^ s_csamul_cla32_fa21_26_xor1;
  assign s_csamul_cla32_fa20_27_and0 = s_csamul_cla32_and20_27 & s_csamul_cla32_fa21_26_xor1;
  assign s_csamul_cla32_fa20_27_xor1 = s_csamul_cla32_fa20_27_xor0 ^ s_csamul_cla32_fa20_26_or0;
  assign s_csamul_cla32_fa20_27_and1 = s_csamul_cla32_fa20_27_xor0 & s_csamul_cla32_fa20_26_or0;
  assign s_csamul_cla32_fa20_27_or0 = s_csamul_cla32_fa20_27_and0 | s_csamul_cla32_fa20_27_and1;
  assign s_csamul_cla32_and21_27 = a[21] & b[27];
  assign s_csamul_cla32_fa21_27_xor0 = s_csamul_cla32_and21_27 ^ s_csamul_cla32_fa22_26_xor1;
  assign s_csamul_cla32_fa21_27_and0 = s_csamul_cla32_and21_27 & s_csamul_cla32_fa22_26_xor1;
  assign s_csamul_cla32_fa21_27_xor1 = s_csamul_cla32_fa21_27_xor0 ^ s_csamul_cla32_fa21_26_or0;
  assign s_csamul_cla32_fa21_27_and1 = s_csamul_cla32_fa21_27_xor0 & s_csamul_cla32_fa21_26_or0;
  assign s_csamul_cla32_fa21_27_or0 = s_csamul_cla32_fa21_27_and0 | s_csamul_cla32_fa21_27_and1;
  assign s_csamul_cla32_and22_27 = a[22] & b[27];
  assign s_csamul_cla32_fa22_27_xor0 = s_csamul_cla32_and22_27 ^ s_csamul_cla32_fa23_26_xor1;
  assign s_csamul_cla32_fa22_27_and0 = s_csamul_cla32_and22_27 & s_csamul_cla32_fa23_26_xor1;
  assign s_csamul_cla32_fa22_27_xor1 = s_csamul_cla32_fa22_27_xor0 ^ s_csamul_cla32_fa22_26_or0;
  assign s_csamul_cla32_fa22_27_and1 = s_csamul_cla32_fa22_27_xor0 & s_csamul_cla32_fa22_26_or0;
  assign s_csamul_cla32_fa22_27_or0 = s_csamul_cla32_fa22_27_and0 | s_csamul_cla32_fa22_27_and1;
  assign s_csamul_cla32_and23_27 = a[23] & b[27];
  assign s_csamul_cla32_fa23_27_xor0 = s_csamul_cla32_and23_27 ^ s_csamul_cla32_fa24_26_xor1;
  assign s_csamul_cla32_fa23_27_and0 = s_csamul_cla32_and23_27 & s_csamul_cla32_fa24_26_xor1;
  assign s_csamul_cla32_fa23_27_xor1 = s_csamul_cla32_fa23_27_xor0 ^ s_csamul_cla32_fa23_26_or0;
  assign s_csamul_cla32_fa23_27_and1 = s_csamul_cla32_fa23_27_xor0 & s_csamul_cla32_fa23_26_or0;
  assign s_csamul_cla32_fa23_27_or0 = s_csamul_cla32_fa23_27_and0 | s_csamul_cla32_fa23_27_and1;
  assign s_csamul_cla32_and24_27 = a[24] & b[27];
  assign s_csamul_cla32_fa24_27_xor0 = s_csamul_cla32_and24_27 ^ s_csamul_cla32_fa25_26_xor1;
  assign s_csamul_cla32_fa24_27_and0 = s_csamul_cla32_and24_27 & s_csamul_cla32_fa25_26_xor1;
  assign s_csamul_cla32_fa24_27_xor1 = s_csamul_cla32_fa24_27_xor0 ^ s_csamul_cla32_fa24_26_or0;
  assign s_csamul_cla32_fa24_27_and1 = s_csamul_cla32_fa24_27_xor0 & s_csamul_cla32_fa24_26_or0;
  assign s_csamul_cla32_fa24_27_or0 = s_csamul_cla32_fa24_27_and0 | s_csamul_cla32_fa24_27_and1;
  assign s_csamul_cla32_and25_27 = a[25] & b[27];
  assign s_csamul_cla32_fa25_27_xor0 = s_csamul_cla32_and25_27 ^ s_csamul_cla32_fa26_26_xor1;
  assign s_csamul_cla32_fa25_27_and0 = s_csamul_cla32_and25_27 & s_csamul_cla32_fa26_26_xor1;
  assign s_csamul_cla32_fa25_27_xor1 = s_csamul_cla32_fa25_27_xor0 ^ s_csamul_cla32_fa25_26_or0;
  assign s_csamul_cla32_fa25_27_and1 = s_csamul_cla32_fa25_27_xor0 & s_csamul_cla32_fa25_26_or0;
  assign s_csamul_cla32_fa25_27_or0 = s_csamul_cla32_fa25_27_and0 | s_csamul_cla32_fa25_27_and1;
  assign s_csamul_cla32_and26_27 = a[26] & b[27];
  assign s_csamul_cla32_fa26_27_xor0 = s_csamul_cla32_and26_27 ^ s_csamul_cla32_fa27_26_xor1;
  assign s_csamul_cla32_fa26_27_and0 = s_csamul_cla32_and26_27 & s_csamul_cla32_fa27_26_xor1;
  assign s_csamul_cla32_fa26_27_xor1 = s_csamul_cla32_fa26_27_xor0 ^ s_csamul_cla32_fa26_26_or0;
  assign s_csamul_cla32_fa26_27_and1 = s_csamul_cla32_fa26_27_xor0 & s_csamul_cla32_fa26_26_or0;
  assign s_csamul_cla32_fa26_27_or0 = s_csamul_cla32_fa26_27_and0 | s_csamul_cla32_fa26_27_and1;
  assign s_csamul_cla32_and27_27 = a[27] & b[27];
  assign s_csamul_cla32_fa27_27_xor0 = s_csamul_cla32_and27_27 ^ s_csamul_cla32_fa28_26_xor1;
  assign s_csamul_cla32_fa27_27_and0 = s_csamul_cla32_and27_27 & s_csamul_cla32_fa28_26_xor1;
  assign s_csamul_cla32_fa27_27_xor1 = s_csamul_cla32_fa27_27_xor0 ^ s_csamul_cla32_fa27_26_or0;
  assign s_csamul_cla32_fa27_27_and1 = s_csamul_cla32_fa27_27_xor0 & s_csamul_cla32_fa27_26_or0;
  assign s_csamul_cla32_fa27_27_or0 = s_csamul_cla32_fa27_27_and0 | s_csamul_cla32_fa27_27_and1;
  assign s_csamul_cla32_and28_27 = a[28] & b[27];
  assign s_csamul_cla32_fa28_27_xor0 = s_csamul_cla32_and28_27 ^ s_csamul_cla32_fa29_26_xor1;
  assign s_csamul_cla32_fa28_27_and0 = s_csamul_cla32_and28_27 & s_csamul_cla32_fa29_26_xor1;
  assign s_csamul_cla32_fa28_27_xor1 = s_csamul_cla32_fa28_27_xor0 ^ s_csamul_cla32_fa28_26_or0;
  assign s_csamul_cla32_fa28_27_and1 = s_csamul_cla32_fa28_27_xor0 & s_csamul_cla32_fa28_26_or0;
  assign s_csamul_cla32_fa28_27_or0 = s_csamul_cla32_fa28_27_and0 | s_csamul_cla32_fa28_27_and1;
  assign s_csamul_cla32_and29_27 = a[29] & b[27];
  assign s_csamul_cla32_fa29_27_xor0 = s_csamul_cla32_and29_27 ^ s_csamul_cla32_fa30_26_xor1;
  assign s_csamul_cla32_fa29_27_and0 = s_csamul_cla32_and29_27 & s_csamul_cla32_fa30_26_xor1;
  assign s_csamul_cla32_fa29_27_xor1 = s_csamul_cla32_fa29_27_xor0 ^ s_csamul_cla32_fa29_26_or0;
  assign s_csamul_cla32_fa29_27_and1 = s_csamul_cla32_fa29_27_xor0 & s_csamul_cla32_fa29_26_or0;
  assign s_csamul_cla32_fa29_27_or0 = s_csamul_cla32_fa29_27_and0 | s_csamul_cla32_fa29_27_and1;
  assign s_csamul_cla32_and30_27 = a[30] & b[27];
  assign s_csamul_cla32_fa30_27_xor0 = s_csamul_cla32_and30_27 ^ s_csamul_cla32_ha31_26_xor0;
  assign s_csamul_cla32_fa30_27_and0 = s_csamul_cla32_and30_27 & s_csamul_cla32_ha31_26_xor0;
  assign s_csamul_cla32_fa30_27_xor1 = s_csamul_cla32_fa30_27_xor0 ^ s_csamul_cla32_fa30_26_or0;
  assign s_csamul_cla32_fa30_27_and1 = s_csamul_cla32_fa30_27_xor0 & s_csamul_cla32_fa30_26_or0;
  assign s_csamul_cla32_fa30_27_or0 = s_csamul_cla32_fa30_27_and0 | s_csamul_cla32_fa30_27_and1;
  assign s_csamul_cla32_nand31_27 = ~(a[31] & b[27]);
  assign s_csamul_cla32_ha31_27_xor0 = s_csamul_cla32_nand31_27 ^ s_csamul_cla32_ha31_26_and0;
  assign s_csamul_cla32_ha31_27_and0 = s_csamul_cla32_nand31_27 & s_csamul_cla32_ha31_26_and0;
  assign s_csamul_cla32_and0_28 = a[0] & b[28];
  assign s_csamul_cla32_fa0_28_xor0 = s_csamul_cla32_and0_28 ^ s_csamul_cla32_fa1_27_xor1;
  assign s_csamul_cla32_fa0_28_and0 = s_csamul_cla32_and0_28 & s_csamul_cla32_fa1_27_xor1;
  assign s_csamul_cla32_fa0_28_xor1 = s_csamul_cla32_fa0_28_xor0 ^ s_csamul_cla32_fa0_27_or0;
  assign s_csamul_cla32_fa0_28_and1 = s_csamul_cla32_fa0_28_xor0 & s_csamul_cla32_fa0_27_or0;
  assign s_csamul_cla32_fa0_28_or0 = s_csamul_cla32_fa0_28_and0 | s_csamul_cla32_fa0_28_and1;
  assign s_csamul_cla32_and1_28 = a[1] & b[28];
  assign s_csamul_cla32_fa1_28_xor0 = s_csamul_cla32_and1_28 ^ s_csamul_cla32_fa2_27_xor1;
  assign s_csamul_cla32_fa1_28_and0 = s_csamul_cla32_and1_28 & s_csamul_cla32_fa2_27_xor1;
  assign s_csamul_cla32_fa1_28_xor1 = s_csamul_cla32_fa1_28_xor0 ^ s_csamul_cla32_fa1_27_or0;
  assign s_csamul_cla32_fa1_28_and1 = s_csamul_cla32_fa1_28_xor0 & s_csamul_cla32_fa1_27_or0;
  assign s_csamul_cla32_fa1_28_or0 = s_csamul_cla32_fa1_28_and0 | s_csamul_cla32_fa1_28_and1;
  assign s_csamul_cla32_and2_28 = a[2] & b[28];
  assign s_csamul_cla32_fa2_28_xor0 = s_csamul_cla32_and2_28 ^ s_csamul_cla32_fa3_27_xor1;
  assign s_csamul_cla32_fa2_28_and0 = s_csamul_cla32_and2_28 & s_csamul_cla32_fa3_27_xor1;
  assign s_csamul_cla32_fa2_28_xor1 = s_csamul_cla32_fa2_28_xor0 ^ s_csamul_cla32_fa2_27_or0;
  assign s_csamul_cla32_fa2_28_and1 = s_csamul_cla32_fa2_28_xor0 & s_csamul_cla32_fa2_27_or0;
  assign s_csamul_cla32_fa2_28_or0 = s_csamul_cla32_fa2_28_and0 | s_csamul_cla32_fa2_28_and1;
  assign s_csamul_cla32_and3_28 = a[3] & b[28];
  assign s_csamul_cla32_fa3_28_xor0 = s_csamul_cla32_and3_28 ^ s_csamul_cla32_fa4_27_xor1;
  assign s_csamul_cla32_fa3_28_and0 = s_csamul_cla32_and3_28 & s_csamul_cla32_fa4_27_xor1;
  assign s_csamul_cla32_fa3_28_xor1 = s_csamul_cla32_fa3_28_xor0 ^ s_csamul_cla32_fa3_27_or0;
  assign s_csamul_cla32_fa3_28_and1 = s_csamul_cla32_fa3_28_xor0 & s_csamul_cla32_fa3_27_or0;
  assign s_csamul_cla32_fa3_28_or0 = s_csamul_cla32_fa3_28_and0 | s_csamul_cla32_fa3_28_and1;
  assign s_csamul_cla32_and4_28 = a[4] & b[28];
  assign s_csamul_cla32_fa4_28_xor0 = s_csamul_cla32_and4_28 ^ s_csamul_cla32_fa5_27_xor1;
  assign s_csamul_cla32_fa4_28_and0 = s_csamul_cla32_and4_28 & s_csamul_cla32_fa5_27_xor1;
  assign s_csamul_cla32_fa4_28_xor1 = s_csamul_cla32_fa4_28_xor0 ^ s_csamul_cla32_fa4_27_or0;
  assign s_csamul_cla32_fa4_28_and1 = s_csamul_cla32_fa4_28_xor0 & s_csamul_cla32_fa4_27_or0;
  assign s_csamul_cla32_fa4_28_or0 = s_csamul_cla32_fa4_28_and0 | s_csamul_cla32_fa4_28_and1;
  assign s_csamul_cla32_and5_28 = a[5] & b[28];
  assign s_csamul_cla32_fa5_28_xor0 = s_csamul_cla32_and5_28 ^ s_csamul_cla32_fa6_27_xor1;
  assign s_csamul_cla32_fa5_28_and0 = s_csamul_cla32_and5_28 & s_csamul_cla32_fa6_27_xor1;
  assign s_csamul_cla32_fa5_28_xor1 = s_csamul_cla32_fa5_28_xor0 ^ s_csamul_cla32_fa5_27_or0;
  assign s_csamul_cla32_fa5_28_and1 = s_csamul_cla32_fa5_28_xor0 & s_csamul_cla32_fa5_27_or0;
  assign s_csamul_cla32_fa5_28_or0 = s_csamul_cla32_fa5_28_and0 | s_csamul_cla32_fa5_28_and1;
  assign s_csamul_cla32_and6_28 = a[6] & b[28];
  assign s_csamul_cla32_fa6_28_xor0 = s_csamul_cla32_and6_28 ^ s_csamul_cla32_fa7_27_xor1;
  assign s_csamul_cla32_fa6_28_and0 = s_csamul_cla32_and6_28 & s_csamul_cla32_fa7_27_xor1;
  assign s_csamul_cla32_fa6_28_xor1 = s_csamul_cla32_fa6_28_xor0 ^ s_csamul_cla32_fa6_27_or0;
  assign s_csamul_cla32_fa6_28_and1 = s_csamul_cla32_fa6_28_xor0 & s_csamul_cla32_fa6_27_or0;
  assign s_csamul_cla32_fa6_28_or0 = s_csamul_cla32_fa6_28_and0 | s_csamul_cla32_fa6_28_and1;
  assign s_csamul_cla32_and7_28 = a[7] & b[28];
  assign s_csamul_cla32_fa7_28_xor0 = s_csamul_cla32_and7_28 ^ s_csamul_cla32_fa8_27_xor1;
  assign s_csamul_cla32_fa7_28_and0 = s_csamul_cla32_and7_28 & s_csamul_cla32_fa8_27_xor1;
  assign s_csamul_cla32_fa7_28_xor1 = s_csamul_cla32_fa7_28_xor0 ^ s_csamul_cla32_fa7_27_or0;
  assign s_csamul_cla32_fa7_28_and1 = s_csamul_cla32_fa7_28_xor0 & s_csamul_cla32_fa7_27_or0;
  assign s_csamul_cla32_fa7_28_or0 = s_csamul_cla32_fa7_28_and0 | s_csamul_cla32_fa7_28_and1;
  assign s_csamul_cla32_and8_28 = a[8] & b[28];
  assign s_csamul_cla32_fa8_28_xor0 = s_csamul_cla32_and8_28 ^ s_csamul_cla32_fa9_27_xor1;
  assign s_csamul_cla32_fa8_28_and0 = s_csamul_cla32_and8_28 & s_csamul_cla32_fa9_27_xor1;
  assign s_csamul_cla32_fa8_28_xor1 = s_csamul_cla32_fa8_28_xor0 ^ s_csamul_cla32_fa8_27_or0;
  assign s_csamul_cla32_fa8_28_and1 = s_csamul_cla32_fa8_28_xor0 & s_csamul_cla32_fa8_27_or0;
  assign s_csamul_cla32_fa8_28_or0 = s_csamul_cla32_fa8_28_and0 | s_csamul_cla32_fa8_28_and1;
  assign s_csamul_cla32_and9_28 = a[9] & b[28];
  assign s_csamul_cla32_fa9_28_xor0 = s_csamul_cla32_and9_28 ^ s_csamul_cla32_fa10_27_xor1;
  assign s_csamul_cla32_fa9_28_and0 = s_csamul_cla32_and9_28 & s_csamul_cla32_fa10_27_xor1;
  assign s_csamul_cla32_fa9_28_xor1 = s_csamul_cla32_fa9_28_xor0 ^ s_csamul_cla32_fa9_27_or0;
  assign s_csamul_cla32_fa9_28_and1 = s_csamul_cla32_fa9_28_xor0 & s_csamul_cla32_fa9_27_or0;
  assign s_csamul_cla32_fa9_28_or0 = s_csamul_cla32_fa9_28_and0 | s_csamul_cla32_fa9_28_and1;
  assign s_csamul_cla32_and10_28 = a[10] & b[28];
  assign s_csamul_cla32_fa10_28_xor0 = s_csamul_cla32_and10_28 ^ s_csamul_cla32_fa11_27_xor1;
  assign s_csamul_cla32_fa10_28_and0 = s_csamul_cla32_and10_28 & s_csamul_cla32_fa11_27_xor1;
  assign s_csamul_cla32_fa10_28_xor1 = s_csamul_cla32_fa10_28_xor0 ^ s_csamul_cla32_fa10_27_or0;
  assign s_csamul_cla32_fa10_28_and1 = s_csamul_cla32_fa10_28_xor0 & s_csamul_cla32_fa10_27_or0;
  assign s_csamul_cla32_fa10_28_or0 = s_csamul_cla32_fa10_28_and0 | s_csamul_cla32_fa10_28_and1;
  assign s_csamul_cla32_and11_28 = a[11] & b[28];
  assign s_csamul_cla32_fa11_28_xor0 = s_csamul_cla32_and11_28 ^ s_csamul_cla32_fa12_27_xor1;
  assign s_csamul_cla32_fa11_28_and0 = s_csamul_cla32_and11_28 & s_csamul_cla32_fa12_27_xor1;
  assign s_csamul_cla32_fa11_28_xor1 = s_csamul_cla32_fa11_28_xor0 ^ s_csamul_cla32_fa11_27_or0;
  assign s_csamul_cla32_fa11_28_and1 = s_csamul_cla32_fa11_28_xor0 & s_csamul_cla32_fa11_27_or0;
  assign s_csamul_cla32_fa11_28_or0 = s_csamul_cla32_fa11_28_and0 | s_csamul_cla32_fa11_28_and1;
  assign s_csamul_cla32_and12_28 = a[12] & b[28];
  assign s_csamul_cla32_fa12_28_xor0 = s_csamul_cla32_and12_28 ^ s_csamul_cla32_fa13_27_xor1;
  assign s_csamul_cla32_fa12_28_and0 = s_csamul_cla32_and12_28 & s_csamul_cla32_fa13_27_xor1;
  assign s_csamul_cla32_fa12_28_xor1 = s_csamul_cla32_fa12_28_xor0 ^ s_csamul_cla32_fa12_27_or0;
  assign s_csamul_cla32_fa12_28_and1 = s_csamul_cla32_fa12_28_xor0 & s_csamul_cla32_fa12_27_or0;
  assign s_csamul_cla32_fa12_28_or0 = s_csamul_cla32_fa12_28_and0 | s_csamul_cla32_fa12_28_and1;
  assign s_csamul_cla32_and13_28 = a[13] & b[28];
  assign s_csamul_cla32_fa13_28_xor0 = s_csamul_cla32_and13_28 ^ s_csamul_cla32_fa14_27_xor1;
  assign s_csamul_cla32_fa13_28_and0 = s_csamul_cla32_and13_28 & s_csamul_cla32_fa14_27_xor1;
  assign s_csamul_cla32_fa13_28_xor1 = s_csamul_cla32_fa13_28_xor0 ^ s_csamul_cla32_fa13_27_or0;
  assign s_csamul_cla32_fa13_28_and1 = s_csamul_cla32_fa13_28_xor0 & s_csamul_cla32_fa13_27_or0;
  assign s_csamul_cla32_fa13_28_or0 = s_csamul_cla32_fa13_28_and0 | s_csamul_cla32_fa13_28_and1;
  assign s_csamul_cla32_and14_28 = a[14] & b[28];
  assign s_csamul_cla32_fa14_28_xor0 = s_csamul_cla32_and14_28 ^ s_csamul_cla32_fa15_27_xor1;
  assign s_csamul_cla32_fa14_28_and0 = s_csamul_cla32_and14_28 & s_csamul_cla32_fa15_27_xor1;
  assign s_csamul_cla32_fa14_28_xor1 = s_csamul_cla32_fa14_28_xor0 ^ s_csamul_cla32_fa14_27_or0;
  assign s_csamul_cla32_fa14_28_and1 = s_csamul_cla32_fa14_28_xor0 & s_csamul_cla32_fa14_27_or0;
  assign s_csamul_cla32_fa14_28_or0 = s_csamul_cla32_fa14_28_and0 | s_csamul_cla32_fa14_28_and1;
  assign s_csamul_cla32_and15_28 = a[15] & b[28];
  assign s_csamul_cla32_fa15_28_xor0 = s_csamul_cla32_and15_28 ^ s_csamul_cla32_fa16_27_xor1;
  assign s_csamul_cla32_fa15_28_and0 = s_csamul_cla32_and15_28 & s_csamul_cla32_fa16_27_xor1;
  assign s_csamul_cla32_fa15_28_xor1 = s_csamul_cla32_fa15_28_xor0 ^ s_csamul_cla32_fa15_27_or0;
  assign s_csamul_cla32_fa15_28_and1 = s_csamul_cla32_fa15_28_xor0 & s_csamul_cla32_fa15_27_or0;
  assign s_csamul_cla32_fa15_28_or0 = s_csamul_cla32_fa15_28_and0 | s_csamul_cla32_fa15_28_and1;
  assign s_csamul_cla32_and16_28 = a[16] & b[28];
  assign s_csamul_cla32_fa16_28_xor0 = s_csamul_cla32_and16_28 ^ s_csamul_cla32_fa17_27_xor1;
  assign s_csamul_cla32_fa16_28_and0 = s_csamul_cla32_and16_28 & s_csamul_cla32_fa17_27_xor1;
  assign s_csamul_cla32_fa16_28_xor1 = s_csamul_cla32_fa16_28_xor0 ^ s_csamul_cla32_fa16_27_or0;
  assign s_csamul_cla32_fa16_28_and1 = s_csamul_cla32_fa16_28_xor0 & s_csamul_cla32_fa16_27_or0;
  assign s_csamul_cla32_fa16_28_or0 = s_csamul_cla32_fa16_28_and0 | s_csamul_cla32_fa16_28_and1;
  assign s_csamul_cla32_and17_28 = a[17] & b[28];
  assign s_csamul_cla32_fa17_28_xor0 = s_csamul_cla32_and17_28 ^ s_csamul_cla32_fa18_27_xor1;
  assign s_csamul_cla32_fa17_28_and0 = s_csamul_cla32_and17_28 & s_csamul_cla32_fa18_27_xor1;
  assign s_csamul_cla32_fa17_28_xor1 = s_csamul_cla32_fa17_28_xor0 ^ s_csamul_cla32_fa17_27_or0;
  assign s_csamul_cla32_fa17_28_and1 = s_csamul_cla32_fa17_28_xor0 & s_csamul_cla32_fa17_27_or0;
  assign s_csamul_cla32_fa17_28_or0 = s_csamul_cla32_fa17_28_and0 | s_csamul_cla32_fa17_28_and1;
  assign s_csamul_cla32_and18_28 = a[18] & b[28];
  assign s_csamul_cla32_fa18_28_xor0 = s_csamul_cla32_and18_28 ^ s_csamul_cla32_fa19_27_xor1;
  assign s_csamul_cla32_fa18_28_and0 = s_csamul_cla32_and18_28 & s_csamul_cla32_fa19_27_xor1;
  assign s_csamul_cla32_fa18_28_xor1 = s_csamul_cla32_fa18_28_xor0 ^ s_csamul_cla32_fa18_27_or0;
  assign s_csamul_cla32_fa18_28_and1 = s_csamul_cla32_fa18_28_xor0 & s_csamul_cla32_fa18_27_or0;
  assign s_csamul_cla32_fa18_28_or0 = s_csamul_cla32_fa18_28_and0 | s_csamul_cla32_fa18_28_and1;
  assign s_csamul_cla32_and19_28 = a[19] & b[28];
  assign s_csamul_cla32_fa19_28_xor0 = s_csamul_cla32_and19_28 ^ s_csamul_cla32_fa20_27_xor1;
  assign s_csamul_cla32_fa19_28_and0 = s_csamul_cla32_and19_28 & s_csamul_cla32_fa20_27_xor1;
  assign s_csamul_cla32_fa19_28_xor1 = s_csamul_cla32_fa19_28_xor0 ^ s_csamul_cla32_fa19_27_or0;
  assign s_csamul_cla32_fa19_28_and1 = s_csamul_cla32_fa19_28_xor0 & s_csamul_cla32_fa19_27_or0;
  assign s_csamul_cla32_fa19_28_or0 = s_csamul_cla32_fa19_28_and0 | s_csamul_cla32_fa19_28_and1;
  assign s_csamul_cla32_and20_28 = a[20] & b[28];
  assign s_csamul_cla32_fa20_28_xor0 = s_csamul_cla32_and20_28 ^ s_csamul_cla32_fa21_27_xor1;
  assign s_csamul_cla32_fa20_28_and0 = s_csamul_cla32_and20_28 & s_csamul_cla32_fa21_27_xor1;
  assign s_csamul_cla32_fa20_28_xor1 = s_csamul_cla32_fa20_28_xor0 ^ s_csamul_cla32_fa20_27_or0;
  assign s_csamul_cla32_fa20_28_and1 = s_csamul_cla32_fa20_28_xor0 & s_csamul_cla32_fa20_27_or0;
  assign s_csamul_cla32_fa20_28_or0 = s_csamul_cla32_fa20_28_and0 | s_csamul_cla32_fa20_28_and1;
  assign s_csamul_cla32_and21_28 = a[21] & b[28];
  assign s_csamul_cla32_fa21_28_xor0 = s_csamul_cla32_and21_28 ^ s_csamul_cla32_fa22_27_xor1;
  assign s_csamul_cla32_fa21_28_and0 = s_csamul_cla32_and21_28 & s_csamul_cla32_fa22_27_xor1;
  assign s_csamul_cla32_fa21_28_xor1 = s_csamul_cla32_fa21_28_xor0 ^ s_csamul_cla32_fa21_27_or0;
  assign s_csamul_cla32_fa21_28_and1 = s_csamul_cla32_fa21_28_xor0 & s_csamul_cla32_fa21_27_or0;
  assign s_csamul_cla32_fa21_28_or0 = s_csamul_cla32_fa21_28_and0 | s_csamul_cla32_fa21_28_and1;
  assign s_csamul_cla32_and22_28 = a[22] & b[28];
  assign s_csamul_cla32_fa22_28_xor0 = s_csamul_cla32_and22_28 ^ s_csamul_cla32_fa23_27_xor1;
  assign s_csamul_cla32_fa22_28_and0 = s_csamul_cla32_and22_28 & s_csamul_cla32_fa23_27_xor1;
  assign s_csamul_cla32_fa22_28_xor1 = s_csamul_cla32_fa22_28_xor0 ^ s_csamul_cla32_fa22_27_or0;
  assign s_csamul_cla32_fa22_28_and1 = s_csamul_cla32_fa22_28_xor0 & s_csamul_cla32_fa22_27_or0;
  assign s_csamul_cla32_fa22_28_or0 = s_csamul_cla32_fa22_28_and0 | s_csamul_cla32_fa22_28_and1;
  assign s_csamul_cla32_and23_28 = a[23] & b[28];
  assign s_csamul_cla32_fa23_28_xor0 = s_csamul_cla32_and23_28 ^ s_csamul_cla32_fa24_27_xor1;
  assign s_csamul_cla32_fa23_28_and0 = s_csamul_cla32_and23_28 & s_csamul_cla32_fa24_27_xor1;
  assign s_csamul_cla32_fa23_28_xor1 = s_csamul_cla32_fa23_28_xor0 ^ s_csamul_cla32_fa23_27_or0;
  assign s_csamul_cla32_fa23_28_and1 = s_csamul_cla32_fa23_28_xor0 & s_csamul_cla32_fa23_27_or0;
  assign s_csamul_cla32_fa23_28_or0 = s_csamul_cla32_fa23_28_and0 | s_csamul_cla32_fa23_28_and1;
  assign s_csamul_cla32_and24_28 = a[24] & b[28];
  assign s_csamul_cla32_fa24_28_xor0 = s_csamul_cla32_and24_28 ^ s_csamul_cla32_fa25_27_xor1;
  assign s_csamul_cla32_fa24_28_and0 = s_csamul_cla32_and24_28 & s_csamul_cla32_fa25_27_xor1;
  assign s_csamul_cla32_fa24_28_xor1 = s_csamul_cla32_fa24_28_xor0 ^ s_csamul_cla32_fa24_27_or0;
  assign s_csamul_cla32_fa24_28_and1 = s_csamul_cla32_fa24_28_xor0 & s_csamul_cla32_fa24_27_or0;
  assign s_csamul_cla32_fa24_28_or0 = s_csamul_cla32_fa24_28_and0 | s_csamul_cla32_fa24_28_and1;
  assign s_csamul_cla32_and25_28 = a[25] & b[28];
  assign s_csamul_cla32_fa25_28_xor0 = s_csamul_cla32_and25_28 ^ s_csamul_cla32_fa26_27_xor1;
  assign s_csamul_cla32_fa25_28_and0 = s_csamul_cla32_and25_28 & s_csamul_cla32_fa26_27_xor1;
  assign s_csamul_cla32_fa25_28_xor1 = s_csamul_cla32_fa25_28_xor0 ^ s_csamul_cla32_fa25_27_or0;
  assign s_csamul_cla32_fa25_28_and1 = s_csamul_cla32_fa25_28_xor0 & s_csamul_cla32_fa25_27_or0;
  assign s_csamul_cla32_fa25_28_or0 = s_csamul_cla32_fa25_28_and0 | s_csamul_cla32_fa25_28_and1;
  assign s_csamul_cla32_and26_28 = a[26] & b[28];
  assign s_csamul_cla32_fa26_28_xor0 = s_csamul_cla32_and26_28 ^ s_csamul_cla32_fa27_27_xor1;
  assign s_csamul_cla32_fa26_28_and0 = s_csamul_cla32_and26_28 & s_csamul_cla32_fa27_27_xor1;
  assign s_csamul_cla32_fa26_28_xor1 = s_csamul_cla32_fa26_28_xor0 ^ s_csamul_cla32_fa26_27_or0;
  assign s_csamul_cla32_fa26_28_and1 = s_csamul_cla32_fa26_28_xor0 & s_csamul_cla32_fa26_27_or0;
  assign s_csamul_cla32_fa26_28_or0 = s_csamul_cla32_fa26_28_and0 | s_csamul_cla32_fa26_28_and1;
  assign s_csamul_cla32_and27_28 = a[27] & b[28];
  assign s_csamul_cla32_fa27_28_xor0 = s_csamul_cla32_and27_28 ^ s_csamul_cla32_fa28_27_xor1;
  assign s_csamul_cla32_fa27_28_and0 = s_csamul_cla32_and27_28 & s_csamul_cla32_fa28_27_xor1;
  assign s_csamul_cla32_fa27_28_xor1 = s_csamul_cla32_fa27_28_xor0 ^ s_csamul_cla32_fa27_27_or0;
  assign s_csamul_cla32_fa27_28_and1 = s_csamul_cla32_fa27_28_xor0 & s_csamul_cla32_fa27_27_or0;
  assign s_csamul_cla32_fa27_28_or0 = s_csamul_cla32_fa27_28_and0 | s_csamul_cla32_fa27_28_and1;
  assign s_csamul_cla32_and28_28 = a[28] & b[28];
  assign s_csamul_cla32_fa28_28_xor0 = s_csamul_cla32_and28_28 ^ s_csamul_cla32_fa29_27_xor1;
  assign s_csamul_cla32_fa28_28_and0 = s_csamul_cla32_and28_28 & s_csamul_cla32_fa29_27_xor1;
  assign s_csamul_cla32_fa28_28_xor1 = s_csamul_cla32_fa28_28_xor0 ^ s_csamul_cla32_fa28_27_or0;
  assign s_csamul_cla32_fa28_28_and1 = s_csamul_cla32_fa28_28_xor0 & s_csamul_cla32_fa28_27_or0;
  assign s_csamul_cla32_fa28_28_or0 = s_csamul_cla32_fa28_28_and0 | s_csamul_cla32_fa28_28_and1;
  assign s_csamul_cla32_and29_28 = a[29] & b[28];
  assign s_csamul_cla32_fa29_28_xor0 = s_csamul_cla32_and29_28 ^ s_csamul_cla32_fa30_27_xor1;
  assign s_csamul_cla32_fa29_28_and0 = s_csamul_cla32_and29_28 & s_csamul_cla32_fa30_27_xor1;
  assign s_csamul_cla32_fa29_28_xor1 = s_csamul_cla32_fa29_28_xor0 ^ s_csamul_cla32_fa29_27_or0;
  assign s_csamul_cla32_fa29_28_and1 = s_csamul_cla32_fa29_28_xor0 & s_csamul_cla32_fa29_27_or0;
  assign s_csamul_cla32_fa29_28_or0 = s_csamul_cla32_fa29_28_and0 | s_csamul_cla32_fa29_28_and1;
  assign s_csamul_cla32_and30_28 = a[30] & b[28];
  assign s_csamul_cla32_fa30_28_xor0 = s_csamul_cla32_and30_28 ^ s_csamul_cla32_ha31_27_xor0;
  assign s_csamul_cla32_fa30_28_and0 = s_csamul_cla32_and30_28 & s_csamul_cla32_ha31_27_xor0;
  assign s_csamul_cla32_fa30_28_xor1 = s_csamul_cla32_fa30_28_xor0 ^ s_csamul_cla32_fa30_27_or0;
  assign s_csamul_cla32_fa30_28_and1 = s_csamul_cla32_fa30_28_xor0 & s_csamul_cla32_fa30_27_or0;
  assign s_csamul_cla32_fa30_28_or0 = s_csamul_cla32_fa30_28_and0 | s_csamul_cla32_fa30_28_and1;
  assign s_csamul_cla32_nand31_28 = ~(a[31] & b[28]);
  assign s_csamul_cla32_ha31_28_xor0 = s_csamul_cla32_nand31_28 ^ s_csamul_cla32_ha31_27_and0;
  assign s_csamul_cla32_ha31_28_and0 = s_csamul_cla32_nand31_28 & s_csamul_cla32_ha31_27_and0;
  assign s_csamul_cla32_and0_29 = a[0] & b[29];
  assign s_csamul_cla32_fa0_29_xor0 = s_csamul_cla32_and0_29 ^ s_csamul_cla32_fa1_28_xor1;
  assign s_csamul_cla32_fa0_29_and0 = s_csamul_cla32_and0_29 & s_csamul_cla32_fa1_28_xor1;
  assign s_csamul_cla32_fa0_29_xor1 = s_csamul_cla32_fa0_29_xor0 ^ s_csamul_cla32_fa0_28_or0;
  assign s_csamul_cla32_fa0_29_and1 = s_csamul_cla32_fa0_29_xor0 & s_csamul_cla32_fa0_28_or0;
  assign s_csamul_cla32_fa0_29_or0 = s_csamul_cla32_fa0_29_and0 | s_csamul_cla32_fa0_29_and1;
  assign s_csamul_cla32_and1_29 = a[1] & b[29];
  assign s_csamul_cla32_fa1_29_xor0 = s_csamul_cla32_and1_29 ^ s_csamul_cla32_fa2_28_xor1;
  assign s_csamul_cla32_fa1_29_and0 = s_csamul_cla32_and1_29 & s_csamul_cla32_fa2_28_xor1;
  assign s_csamul_cla32_fa1_29_xor1 = s_csamul_cla32_fa1_29_xor0 ^ s_csamul_cla32_fa1_28_or0;
  assign s_csamul_cla32_fa1_29_and1 = s_csamul_cla32_fa1_29_xor0 & s_csamul_cla32_fa1_28_or0;
  assign s_csamul_cla32_fa1_29_or0 = s_csamul_cla32_fa1_29_and0 | s_csamul_cla32_fa1_29_and1;
  assign s_csamul_cla32_and2_29 = a[2] & b[29];
  assign s_csamul_cla32_fa2_29_xor0 = s_csamul_cla32_and2_29 ^ s_csamul_cla32_fa3_28_xor1;
  assign s_csamul_cla32_fa2_29_and0 = s_csamul_cla32_and2_29 & s_csamul_cla32_fa3_28_xor1;
  assign s_csamul_cla32_fa2_29_xor1 = s_csamul_cla32_fa2_29_xor0 ^ s_csamul_cla32_fa2_28_or0;
  assign s_csamul_cla32_fa2_29_and1 = s_csamul_cla32_fa2_29_xor0 & s_csamul_cla32_fa2_28_or0;
  assign s_csamul_cla32_fa2_29_or0 = s_csamul_cla32_fa2_29_and0 | s_csamul_cla32_fa2_29_and1;
  assign s_csamul_cla32_and3_29 = a[3] & b[29];
  assign s_csamul_cla32_fa3_29_xor0 = s_csamul_cla32_and3_29 ^ s_csamul_cla32_fa4_28_xor1;
  assign s_csamul_cla32_fa3_29_and0 = s_csamul_cla32_and3_29 & s_csamul_cla32_fa4_28_xor1;
  assign s_csamul_cla32_fa3_29_xor1 = s_csamul_cla32_fa3_29_xor0 ^ s_csamul_cla32_fa3_28_or0;
  assign s_csamul_cla32_fa3_29_and1 = s_csamul_cla32_fa3_29_xor0 & s_csamul_cla32_fa3_28_or0;
  assign s_csamul_cla32_fa3_29_or0 = s_csamul_cla32_fa3_29_and0 | s_csamul_cla32_fa3_29_and1;
  assign s_csamul_cla32_and4_29 = a[4] & b[29];
  assign s_csamul_cla32_fa4_29_xor0 = s_csamul_cla32_and4_29 ^ s_csamul_cla32_fa5_28_xor1;
  assign s_csamul_cla32_fa4_29_and0 = s_csamul_cla32_and4_29 & s_csamul_cla32_fa5_28_xor1;
  assign s_csamul_cla32_fa4_29_xor1 = s_csamul_cla32_fa4_29_xor0 ^ s_csamul_cla32_fa4_28_or0;
  assign s_csamul_cla32_fa4_29_and1 = s_csamul_cla32_fa4_29_xor0 & s_csamul_cla32_fa4_28_or0;
  assign s_csamul_cla32_fa4_29_or0 = s_csamul_cla32_fa4_29_and0 | s_csamul_cla32_fa4_29_and1;
  assign s_csamul_cla32_and5_29 = a[5] & b[29];
  assign s_csamul_cla32_fa5_29_xor0 = s_csamul_cla32_and5_29 ^ s_csamul_cla32_fa6_28_xor1;
  assign s_csamul_cla32_fa5_29_and0 = s_csamul_cla32_and5_29 & s_csamul_cla32_fa6_28_xor1;
  assign s_csamul_cla32_fa5_29_xor1 = s_csamul_cla32_fa5_29_xor0 ^ s_csamul_cla32_fa5_28_or0;
  assign s_csamul_cla32_fa5_29_and1 = s_csamul_cla32_fa5_29_xor0 & s_csamul_cla32_fa5_28_or0;
  assign s_csamul_cla32_fa5_29_or0 = s_csamul_cla32_fa5_29_and0 | s_csamul_cla32_fa5_29_and1;
  assign s_csamul_cla32_and6_29 = a[6] & b[29];
  assign s_csamul_cla32_fa6_29_xor0 = s_csamul_cla32_and6_29 ^ s_csamul_cla32_fa7_28_xor1;
  assign s_csamul_cla32_fa6_29_and0 = s_csamul_cla32_and6_29 & s_csamul_cla32_fa7_28_xor1;
  assign s_csamul_cla32_fa6_29_xor1 = s_csamul_cla32_fa6_29_xor0 ^ s_csamul_cla32_fa6_28_or0;
  assign s_csamul_cla32_fa6_29_and1 = s_csamul_cla32_fa6_29_xor0 & s_csamul_cla32_fa6_28_or0;
  assign s_csamul_cla32_fa6_29_or0 = s_csamul_cla32_fa6_29_and0 | s_csamul_cla32_fa6_29_and1;
  assign s_csamul_cla32_and7_29 = a[7] & b[29];
  assign s_csamul_cla32_fa7_29_xor0 = s_csamul_cla32_and7_29 ^ s_csamul_cla32_fa8_28_xor1;
  assign s_csamul_cla32_fa7_29_and0 = s_csamul_cla32_and7_29 & s_csamul_cla32_fa8_28_xor1;
  assign s_csamul_cla32_fa7_29_xor1 = s_csamul_cla32_fa7_29_xor0 ^ s_csamul_cla32_fa7_28_or0;
  assign s_csamul_cla32_fa7_29_and1 = s_csamul_cla32_fa7_29_xor0 & s_csamul_cla32_fa7_28_or0;
  assign s_csamul_cla32_fa7_29_or0 = s_csamul_cla32_fa7_29_and0 | s_csamul_cla32_fa7_29_and1;
  assign s_csamul_cla32_and8_29 = a[8] & b[29];
  assign s_csamul_cla32_fa8_29_xor0 = s_csamul_cla32_and8_29 ^ s_csamul_cla32_fa9_28_xor1;
  assign s_csamul_cla32_fa8_29_and0 = s_csamul_cla32_and8_29 & s_csamul_cla32_fa9_28_xor1;
  assign s_csamul_cla32_fa8_29_xor1 = s_csamul_cla32_fa8_29_xor0 ^ s_csamul_cla32_fa8_28_or0;
  assign s_csamul_cla32_fa8_29_and1 = s_csamul_cla32_fa8_29_xor0 & s_csamul_cla32_fa8_28_or0;
  assign s_csamul_cla32_fa8_29_or0 = s_csamul_cla32_fa8_29_and0 | s_csamul_cla32_fa8_29_and1;
  assign s_csamul_cla32_and9_29 = a[9] & b[29];
  assign s_csamul_cla32_fa9_29_xor0 = s_csamul_cla32_and9_29 ^ s_csamul_cla32_fa10_28_xor1;
  assign s_csamul_cla32_fa9_29_and0 = s_csamul_cla32_and9_29 & s_csamul_cla32_fa10_28_xor1;
  assign s_csamul_cla32_fa9_29_xor1 = s_csamul_cla32_fa9_29_xor0 ^ s_csamul_cla32_fa9_28_or0;
  assign s_csamul_cla32_fa9_29_and1 = s_csamul_cla32_fa9_29_xor0 & s_csamul_cla32_fa9_28_or0;
  assign s_csamul_cla32_fa9_29_or0 = s_csamul_cla32_fa9_29_and0 | s_csamul_cla32_fa9_29_and1;
  assign s_csamul_cla32_and10_29 = a[10] & b[29];
  assign s_csamul_cla32_fa10_29_xor0 = s_csamul_cla32_and10_29 ^ s_csamul_cla32_fa11_28_xor1;
  assign s_csamul_cla32_fa10_29_and0 = s_csamul_cla32_and10_29 & s_csamul_cla32_fa11_28_xor1;
  assign s_csamul_cla32_fa10_29_xor1 = s_csamul_cla32_fa10_29_xor0 ^ s_csamul_cla32_fa10_28_or0;
  assign s_csamul_cla32_fa10_29_and1 = s_csamul_cla32_fa10_29_xor0 & s_csamul_cla32_fa10_28_or0;
  assign s_csamul_cla32_fa10_29_or0 = s_csamul_cla32_fa10_29_and0 | s_csamul_cla32_fa10_29_and1;
  assign s_csamul_cla32_and11_29 = a[11] & b[29];
  assign s_csamul_cla32_fa11_29_xor0 = s_csamul_cla32_and11_29 ^ s_csamul_cla32_fa12_28_xor1;
  assign s_csamul_cla32_fa11_29_and0 = s_csamul_cla32_and11_29 & s_csamul_cla32_fa12_28_xor1;
  assign s_csamul_cla32_fa11_29_xor1 = s_csamul_cla32_fa11_29_xor0 ^ s_csamul_cla32_fa11_28_or0;
  assign s_csamul_cla32_fa11_29_and1 = s_csamul_cla32_fa11_29_xor0 & s_csamul_cla32_fa11_28_or0;
  assign s_csamul_cla32_fa11_29_or0 = s_csamul_cla32_fa11_29_and0 | s_csamul_cla32_fa11_29_and1;
  assign s_csamul_cla32_and12_29 = a[12] & b[29];
  assign s_csamul_cla32_fa12_29_xor0 = s_csamul_cla32_and12_29 ^ s_csamul_cla32_fa13_28_xor1;
  assign s_csamul_cla32_fa12_29_and0 = s_csamul_cla32_and12_29 & s_csamul_cla32_fa13_28_xor1;
  assign s_csamul_cla32_fa12_29_xor1 = s_csamul_cla32_fa12_29_xor0 ^ s_csamul_cla32_fa12_28_or0;
  assign s_csamul_cla32_fa12_29_and1 = s_csamul_cla32_fa12_29_xor0 & s_csamul_cla32_fa12_28_or0;
  assign s_csamul_cla32_fa12_29_or0 = s_csamul_cla32_fa12_29_and0 | s_csamul_cla32_fa12_29_and1;
  assign s_csamul_cla32_and13_29 = a[13] & b[29];
  assign s_csamul_cla32_fa13_29_xor0 = s_csamul_cla32_and13_29 ^ s_csamul_cla32_fa14_28_xor1;
  assign s_csamul_cla32_fa13_29_and0 = s_csamul_cla32_and13_29 & s_csamul_cla32_fa14_28_xor1;
  assign s_csamul_cla32_fa13_29_xor1 = s_csamul_cla32_fa13_29_xor0 ^ s_csamul_cla32_fa13_28_or0;
  assign s_csamul_cla32_fa13_29_and1 = s_csamul_cla32_fa13_29_xor0 & s_csamul_cla32_fa13_28_or0;
  assign s_csamul_cla32_fa13_29_or0 = s_csamul_cla32_fa13_29_and0 | s_csamul_cla32_fa13_29_and1;
  assign s_csamul_cla32_and14_29 = a[14] & b[29];
  assign s_csamul_cla32_fa14_29_xor0 = s_csamul_cla32_and14_29 ^ s_csamul_cla32_fa15_28_xor1;
  assign s_csamul_cla32_fa14_29_and0 = s_csamul_cla32_and14_29 & s_csamul_cla32_fa15_28_xor1;
  assign s_csamul_cla32_fa14_29_xor1 = s_csamul_cla32_fa14_29_xor0 ^ s_csamul_cla32_fa14_28_or0;
  assign s_csamul_cla32_fa14_29_and1 = s_csamul_cla32_fa14_29_xor0 & s_csamul_cla32_fa14_28_or0;
  assign s_csamul_cla32_fa14_29_or0 = s_csamul_cla32_fa14_29_and0 | s_csamul_cla32_fa14_29_and1;
  assign s_csamul_cla32_and15_29 = a[15] & b[29];
  assign s_csamul_cla32_fa15_29_xor0 = s_csamul_cla32_and15_29 ^ s_csamul_cla32_fa16_28_xor1;
  assign s_csamul_cla32_fa15_29_and0 = s_csamul_cla32_and15_29 & s_csamul_cla32_fa16_28_xor1;
  assign s_csamul_cla32_fa15_29_xor1 = s_csamul_cla32_fa15_29_xor0 ^ s_csamul_cla32_fa15_28_or0;
  assign s_csamul_cla32_fa15_29_and1 = s_csamul_cla32_fa15_29_xor0 & s_csamul_cla32_fa15_28_or0;
  assign s_csamul_cla32_fa15_29_or0 = s_csamul_cla32_fa15_29_and0 | s_csamul_cla32_fa15_29_and1;
  assign s_csamul_cla32_and16_29 = a[16] & b[29];
  assign s_csamul_cla32_fa16_29_xor0 = s_csamul_cla32_and16_29 ^ s_csamul_cla32_fa17_28_xor1;
  assign s_csamul_cla32_fa16_29_and0 = s_csamul_cla32_and16_29 & s_csamul_cla32_fa17_28_xor1;
  assign s_csamul_cla32_fa16_29_xor1 = s_csamul_cla32_fa16_29_xor0 ^ s_csamul_cla32_fa16_28_or0;
  assign s_csamul_cla32_fa16_29_and1 = s_csamul_cla32_fa16_29_xor0 & s_csamul_cla32_fa16_28_or0;
  assign s_csamul_cla32_fa16_29_or0 = s_csamul_cla32_fa16_29_and0 | s_csamul_cla32_fa16_29_and1;
  assign s_csamul_cla32_and17_29 = a[17] & b[29];
  assign s_csamul_cla32_fa17_29_xor0 = s_csamul_cla32_and17_29 ^ s_csamul_cla32_fa18_28_xor1;
  assign s_csamul_cla32_fa17_29_and0 = s_csamul_cla32_and17_29 & s_csamul_cla32_fa18_28_xor1;
  assign s_csamul_cla32_fa17_29_xor1 = s_csamul_cla32_fa17_29_xor0 ^ s_csamul_cla32_fa17_28_or0;
  assign s_csamul_cla32_fa17_29_and1 = s_csamul_cla32_fa17_29_xor0 & s_csamul_cla32_fa17_28_or0;
  assign s_csamul_cla32_fa17_29_or0 = s_csamul_cla32_fa17_29_and0 | s_csamul_cla32_fa17_29_and1;
  assign s_csamul_cla32_and18_29 = a[18] & b[29];
  assign s_csamul_cla32_fa18_29_xor0 = s_csamul_cla32_and18_29 ^ s_csamul_cla32_fa19_28_xor1;
  assign s_csamul_cla32_fa18_29_and0 = s_csamul_cla32_and18_29 & s_csamul_cla32_fa19_28_xor1;
  assign s_csamul_cla32_fa18_29_xor1 = s_csamul_cla32_fa18_29_xor0 ^ s_csamul_cla32_fa18_28_or0;
  assign s_csamul_cla32_fa18_29_and1 = s_csamul_cla32_fa18_29_xor0 & s_csamul_cla32_fa18_28_or0;
  assign s_csamul_cla32_fa18_29_or0 = s_csamul_cla32_fa18_29_and0 | s_csamul_cla32_fa18_29_and1;
  assign s_csamul_cla32_and19_29 = a[19] & b[29];
  assign s_csamul_cla32_fa19_29_xor0 = s_csamul_cla32_and19_29 ^ s_csamul_cla32_fa20_28_xor1;
  assign s_csamul_cla32_fa19_29_and0 = s_csamul_cla32_and19_29 & s_csamul_cla32_fa20_28_xor1;
  assign s_csamul_cla32_fa19_29_xor1 = s_csamul_cla32_fa19_29_xor0 ^ s_csamul_cla32_fa19_28_or0;
  assign s_csamul_cla32_fa19_29_and1 = s_csamul_cla32_fa19_29_xor0 & s_csamul_cla32_fa19_28_or0;
  assign s_csamul_cla32_fa19_29_or0 = s_csamul_cla32_fa19_29_and0 | s_csamul_cla32_fa19_29_and1;
  assign s_csamul_cla32_and20_29 = a[20] & b[29];
  assign s_csamul_cla32_fa20_29_xor0 = s_csamul_cla32_and20_29 ^ s_csamul_cla32_fa21_28_xor1;
  assign s_csamul_cla32_fa20_29_and0 = s_csamul_cla32_and20_29 & s_csamul_cla32_fa21_28_xor1;
  assign s_csamul_cla32_fa20_29_xor1 = s_csamul_cla32_fa20_29_xor0 ^ s_csamul_cla32_fa20_28_or0;
  assign s_csamul_cla32_fa20_29_and1 = s_csamul_cla32_fa20_29_xor0 & s_csamul_cla32_fa20_28_or0;
  assign s_csamul_cla32_fa20_29_or0 = s_csamul_cla32_fa20_29_and0 | s_csamul_cla32_fa20_29_and1;
  assign s_csamul_cla32_and21_29 = a[21] & b[29];
  assign s_csamul_cla32_fa21_29_xor0 = s_csamul_cla32_and21_29 ^ s_csamul_cla32_fa22_28_xor1;
  assign s_csamul_cla32_fa21_29_and0 = s_csamul_cla32_and21_29 & s_csamul_cla32_fa22_28_xor1;
  assign s_csamul_cla32_fa21_29_xor1 = s_csamul_cla32_fa21_29_xor0 ^ s_csamul_cla32_fa21_28_or0;
  assign s_csamul_cla32_fa21_29_and1 = s_csamul_cla32_fa21_29_xor0 & s_csamul_cla32_fa21_28_or0;
  assign s_csamul_cla32_fa21_29_or0 = s_csamul_cla32_fa21_29_and0 | s_csamul_cla32_fa21_29_and1;
  assign s_csamul_cla32_and22_29 = a[22] & b[29];
  assign s_csamul_cla32_fa22_29_xor0 = s_csamul_cla32_and22_29 ^ s_csamul_cla32_fa23_28_xor1;
  assign s_csamul_cla32_fa22_29_and0 = s_csamul_cla32_and22_29 & s_csamul_cla32_fa23_28_xor1;
  assign s_csamul_cla32_fa22_29_xor1 = s_csamul_cla32_fa22_29_xor0 ^ s_csamul_cla32_fa22_28_or0;
  assign s_csamul_cla32_fa22_29_and1 = s_csamul_cla32_fa22_29_xor0 & s_csamul_cla32_fa22_28_or0;
  assign s_csamul_cla32_fa22_29_or0 = s_csamul_cla32_fa22_29_and0 | s_csamul_cla32_fa22_29_and1;
  assign s_csamul_cla32_and23_29 = a[23] & b[29];
  assign s_csamul_cla32_fa23_29_xor0 = s_csamul_cla32_and23_29 ^ s_csamul_cla32_fa24_28_xor1;
  assign s_csamul_cla32_fa23_29_and0 = s_csamul_cla32_and23_29 & s_csamul_cla32_fa24_28_xor1;
  assign s_csamul_cla32_fa23_29_xor1 = s_csamul_cla32_fa23_29_xor0 ^ s_csamul_cla32_fa23_28_or0;
  assign s_csamul_cla32_fa23_29_and1 = s_csamul_cla32_fa23_29_xor0 & s_csamul_cla32_fa23_28_or0;
  assign s_csamul_cla32_fa23_29_or0 = s_csamul_cla32_fa23_29_and0 | s_csamul_cla32_fa23_29_and1;
  assign s_csamul_cla32_and24_29 = a[24] & b[29];
  assign s_csamul_cla32_fa24_29_xor0 = s_csamul_cla32_and24_29 ^ s_csamul_cla32_fa25_28_xor1;
  assign s_csamul_cla32_fa24_29_and0 = s_csamul_cla32_and24_29 & s_csamul_cla32_fa25_28_xor1;
  assign s_csamul_cla32_fa24_29_xor1 = s_csamul_cla32_fa24_29_xor0 ^ s_csamul_cla32_fa24_28_or0;
  assign s_csamul_cla32_fa24_29_and1 = s_csamul_cla32_fa24_29_xor0 & s_csamul_cla32_fa24_28_or0;
  assign s_csamul_cla32_fa24_29_or0 = s_csamul_cla32_fa24_29_and0 | s_csamul_cla32_fa24_29_and1;
  assign s_csamul_cla32_and25_29 = a[25] & b[29];
  assign s_csamul_cla32_fa25_29_xor0 = s_csamul_cla32_and25_29 ^ s_csamul_cla32_fa26_28_xor1;
  assign s_csamul_cla32_fa25_29_and0 = s_csamul_cla32_and25_29 & s_csamul_cla32_fa26_28_xor1;
  assign s_csamul_cla32_fa25_29_xor1 = s_csamul_cla32_fa25_29_xor0 ^ s_csamul_cla32_fa25_28_or0;
  assign s_csamul_cla32_fa25_29_and1 = s_csamul_cla32_fa25_29_xor0 & s_csamul_cla32_fa25_28_or0;
  assign s_csamul_cla32_fa25_29_or0 = s_csamul_cla32_fa25_29_and0 | s_csamul_cla32_fa25_29_and1;
  assign s_csamul_cla32_and26_29 = a[26] & b[29];
  assign s_csamul_cla32_fa26_29_xor0 = s_csamul_cla32_and26_29 ^ s_csamul_cla32_fa27_28_xor1;
  assign s_csamul_cla32_fa26_29_and0 = s_csamul_cla32_and26_29 & s_csamul_cla32_fa27_28_xor1;
  assign s_csamul_cla32_fa26_29_xor1 = s_csamul_cla32_fa26_29_xor0 ^ s_csamul_cla32_fa26_28_or0;
  assign s_csamul_cla32_fa26_29_and1 = s_csamul_cla32_fa26_29_xor0 & s_csamul_cla32_fa26_28_or0;
  assign s_csamul_cla32_fa26_29_or0 = s_csamul_cla32_fa26_29_and0 | s_csamul_cla32_fa26_29_and1;
  assign s_csamul_cla32_and27_29 = a[27] & b[29];
  assign s_csamul_cla32_fa27_29_xor0 = s_csamul_cla32_and27_29 ^ s_csamul_cla32_fa28_28_xor1;
  assign s_csamul_cla32_fa27_29_and0 = s_csamul_cla32_and27_29 & s_csamul_cla32_fa28_28_xor1;
  assign s_csamul_cla32_fa27_29_xor1 = s_csamul_cla32_fa27_29_xor0 ^ s_csamul_cla32_fa27_28_or0;
  assign s_csamul_cla32_fa27_29_and1 = s_csamul_cla32_fa27_29_xor0 & s_csamul_cla32_fa27_28_or0;
  assign s_csamul_cla32_fa27_29_or0 = s_csamul_cla32_fa27_29_and0 | s_csamul_cla32_fa27_29_and1;
  assign s_csamul_cla32_and28_29 = a[28] & b[29];
  assign s_csamul_cla32_fa28_29_xor0 = s_csamul_cla32_and28_29 ^ s_csamul_cla32_fa29_28_xor1;
  assign s_csamul_cla32_fa28_29_and0 = s_csamul_cla32_and28_29 & s_csamul_cla32_fa29_28_xor1;
  assign s_csamul_cla32_fa28_29_xor1 = s_csamul_cla32_fa28_29_xor0 ^ s_csamul_cla32_fa28_28_or0;
  assign s_csamul_cla32_fa28_29_and1 = s_csamul_cla32_fa28_29_xor0 & s_csamul_cla32_fa28_28_or0;
  assign s_csamul_cla32_fa28_29_or0 = s_csamul_cla32_fa28_29_and0 | s_csamul_cla32_fa28_29_and1;
  assign s_csamul_cla32_and29_29 = a[29] & b[29];
  assign s_csamul_cla32_fa29_29_xor0 = s_csamul_cla32_and29_29 ^ s_csamul_cla32_fa30_28_xor1;
  assign s_csamul_cla32_fa29_29_and0 = s_csamul_cla32_and29_29 & s_csamul_cla32_fa30_28_xor1;
  assign s_csamul_cla32_fa29_29_xor1 = s_csamul_cla32_fa29_29_xor0 ^ s_csamul_cla32_fa29_28_or0;
  assign s_csamul_cla32_fa29_29_and1 = s_csamul_cla32_fa29_29_xor0 & s_csamul_cla32_fa29_28_or0;
  assign s_csamul_cla32_fa29_29_or0 = s_csamul_cla32_fa29_29_and0 | s_csamul_cla32_fa29_29_and1;
  assign s_csamul_cla32_and30_29 = a[30] & b[29];
  assign s_csamul_cla32_fa30_29_xor0 = s_csamul_cla32_and30_29 ^ s_csamul_cla32_ha31_28_xor0;
  assign s_csamul_cla32_fa30_29_and0 = s_csamul_cla32_and30_29 & s_csamul_cla32_ha31_28_xor0;
  assign s_csamul_cla32_fa30_29_xor1 = s_csamul_cla32_fa30_29_xor0 ^ s_csamul_cla32_fa30_28_or0;
  assign s_csamul_cla32_fa30_29_and1 = s_csamul_cla32_fa30_29_xor0 & s_csamul_cla32_fa30_28_or0;
  assign s_csamul_cla32_fa30_29_or0 = s_csamul_cla32_fa30_29_and0 | s_csamul_cla32_fa30_29_and1;
  assign s_csamul_cla32_nand31_29 = ~(a[31] & b[29]);
  assign s_csamul_cla32_ha31_29_xor0 = s_csamul_cla32_nand31_29 ^ s_csamul_cla32_ha31_28_and0;
  assign s_csamul_cla32_ha31_29_and0 = s_csamul_cla32_nand31_29 & s_csamul_cla32_ha31_28_and0;
  assign s_csamul_cla32_and0_30 = a[0] & b[30];
  assign s_csamul_cla32_fa0_30_xor0 = s_csamul_cla32_and0_30 ^ s_csamul_cla32_fa1_29_xor1;
  assign s_csamul_cla32_fa0_30_and0 = s_csamul_cla32_and0_30 & s_csamul_cla32_fa1_29_xor1;
  assign s_csamul_cla32_fa0_30_xor1 = s_csamul_cla32_fa0_30_xor0 ^ s_csamul_cla32_fa0_29_or0;
  assign s_csamul_cla32_fa0_30_and1 = s_csamul_cla32_fa0_30_xor0 & s_csamul_cla32_fa0_29_or0;
  assign s_csamul_cla32_fa0_30_or0 = s_csamul_cla32_fa0_30_and0 | s_csamul_cla32_fa0_30_and1;
  assign s_csamul_cla32_and1_30 = a[1] & b[30];
  assign s_csamul_cla32_fa1_30_xor0 = s_csamul_cla32_and1_30 ^ s_csamul_cla32_fa2_29_xor1;
  assign s_csamul_cla32_fa1_30_and0 = s_csamul_cla32_and1_30 & s_csamul_cla32_fa2_29_xor1;
  assign s_csamul_cla32_fa1_30_xor1 = s_csamul_cla32_fa1_30_xor0 ^ s_csamul_cla32_fa1_29_or0;
  assign s_csamul_cla32_fa1_30_and1 = s_csamul_cla32_fa1_30_xor0 & s_csamul_cla32_fa1_29_or0;
  assign s_csamul_cla32_fa1_30_or0 = s_csamul_cla32_fa1_30_and0 | s_csamul_cla32_fa1_30_and1;
  assign s_csamul_cla32_and2_30 = a[2] & b[30];
  assign s_csamul_cla32_fa2_30_xor0 = s_csamul_cla32_and2_30 ^ s_csamul_cla32_fa3_29_xor1;
  assign s_csamul_cla32_fa2_30_and0 = s_csamul_cla32_and2_30 & s_csamul_cla32_fa3_29_xor1;
  assign s_csamul_cla32_fa2_30_xor1 = s_csamul_cla32_fa2_30_xor0 ^ s_csamul_cla32_fa2_29_or0;
  assign s_csamul_cla32_fa2_30_and1 = s_csamul_cla32_fa2_30_xor0 & s_csamul_cla32_fa2_29_or0;
  assign s_csamul_cla32_fa2_30_or0 = s_csamul_cla32_fa2_30_and0 | s_csamul_cla32_fa2_30_and1;
  assign s_csamul_cla32_and3_30 = a[3] & b[30];
  assign s_csamul_cla32_fa3_30_xor0 = s_csamul_cla32_and3_30 ^ s_csamul_cla32_fa4_29_xor1;
  assign s_csamul_cla32_fa3_30_and0 = s_csamul_cla32_and3_30 & s_csamul_cla32_fa4_29_xor1;
  assign s_csamul_cla32_fa3_30_xor1 = s_csamul_cla32_fa3_30_xor0 ^ s_csamul_cla32_fa3_29_or0;
  assign s_csamul_cla32_fa3_30_and1 = s_csamul_cla32_fa3_30_xor0 & s_csamul_cla32_fa3_29_or0;
  assign s_csamul_cla32_fa3_30_or0 = s_csamul_cla32_fa3_30_and0 | s_csamul_cla32_fa3_30_and1;
  assign s_csamul_cla32_and4_30 = a[4] & b[30];
  assign s_csamul_cla32_fa4_30_xor0 = s_csamul_cla32_and4_30 ^ s_csamul_cla32_fa5_29_xor1;
  assign s_csamul_cla32_fa4_30_and0 = s_csamul_cla32_and4_30 & s_csamul_cla32_fa5_29_xor1;
  assign s_csamul_cla32_fa4_30_xor1 = s_csamul_cla32_fa4_30_xor0 ^ s_csamul_cla32_fa4_29_or0;
  assign s_csamul_cla32_fa4_30_and1 = s_csamul_cla32_fa4_30_xor0 & s_csamul_cla32_fa4_29_or0;
  assign s_csamul_cla32_fa4_30_or0 = s_csamul_cla32_fa4_30_and0 | s_csamul_cla32_fa4_30_and1;
  assign s_csamul_cla32_and5_30 = a[5] & b[30];
  assign s_csamul_cla32_fa5_30_xor0 = s_csamul_cla32_and5_30 ^ s_csamul_cla32_fa6_29_xor1;
  assign s_csamul_cla32_fa5_30_and0 = s_csamul_cla32_and5_30 & s_csamul_cla32_fa6_29_xor1;
  assign s_csamul_cla32_fa5_30_xor1 = s_csamul_cla32_fa5_30_xor0 ^ s_csamul_cla32_fa5_29_or0;
  assign s_csamul_cla32_fa5_30_and1 = s_csamul_cla32_fa5_30_xor0 & s_csamul_cla32_fa5_29_or0;
  assign s_csamul_cla32_fa5_30_or0 = s_csamul_cla32_fa5_30_and0 | s_csamul_cla32_fa5_30_and1;
  assign s_csamul_cla32_and6_30 = a[6] & b[30];
  assign s_csamul_cla32_fa6_30_xor0 = s_csamul_cla32_and6_30 ^ s_csamul_cla32_fa7_29_xor1;
  assign s_csamul_cla32_fa6_30_and0 = s_csamul_cla32_and6_30 & s_csamul_cla32_fa7_29_xor1;
  assign s_csamul_cla32_fa6_30_xor1 = s_csamul_cla32_fa6_30_xor0 ^ s_csamul_cla32_fa6_29_or0;
  assign s_csamul_cla32_fa6_30_and1 = s_csamul_cla32_fa6_30_xor0 & s_csamul_cla32_fa6_29_or0;
  assign s_csamul_cla32_fa6_30_or0 = s_csamul_cla32_fa6_30_and0 | s_csamul_cla32_fa6_30_and1;
  assign s_csamul_cla32_and7_30 = a[7] & b[30];
  assign s_csamul_cla32_fa7_30_xor0 = s_csamul_cla32_and7_30 ^ s_csamul_cla32_fa8_29_xor1;
  assign s_csamul_cla32_fa7_30_and0 = s_csamul_cla32_and7_30 & s_csamul_cla32_fa8_29_xor1;
  assign s_csamul_cla32_fa7_30_xor1 = s_csamul_cla32_fa7_30_xor0 ^ s_csamul_cla32_fa7_29_or0;
  assign s_csamul_cla32_fa7_30_and1 = s_csamul_cla32_fa7_30_xor0 & s_csamul_cla32_fa7_29_or0;
  assign s_csamul_cla32_fa7_30_or0 = s_csamul_cla32_fa7_30_and0 | s_csamul_cla32_fa7_30_and1;
  assign s_csamul_cla32_and8_30 = a[8] & b[30];
  assign s_csamul_cla32_fa8_30_xor0 = s_csamul_cla32_and8_30 ^ s_csamul_cla32_fa9_29_xor1;
  assign s_csamul_cla32_fa8_30_and0 = s_csamul_cla32_and8_30 & s_csamul_cla32_fa9_29_xor1;
  assign s_csamul_cla32_fa8_30_xor1 = s_csamul_cla32_fa8_30_xor0 ^ s_csamul_cla32_fa8_29_or0;
  assign s_csamul_cla32_fa8_30_and1 = s_csamul_cla32_fa8_30_xor0 & s_csamul_cla32_fa8_29_or0;
  assign s_csamul_cla32_fa8_30_or0 = s_csamul_cla32_fa8_30_and0 | s_csamul_cla32_fa8_30_and1;
  assign s_csamul_cla32_and9_30 = a[9] & b[30];
  assign s_csamul_cla32_fa9_30_xor0 = s_csamul_cla32_and9_30 ^ s_csamul_cla32_fa10_29_xor1;
  assign s_csamul_cla32_fa9_30_and0 = s_csamul_cla32_and9_30 & s_csamul_cla32_fa10_29_xor1;
  assign s_csamul_cla32_fa9_30_xor1 = s_csamul_cla32_fa9_30_xor0 ^ s_csamul_cla32_fa9_29_or0;
  assign s_csamul_cla32_fa9_30_and1 = s_csamul_cla32_fa9_30_xor0 & s_csamul_cla32_fa9_29_or0;
  assign s_csamul_cla32_fa9_30_or0 = s_csamul_cla32_fa9_30_and0 | s_csamul_cla32_fa9_30_and1;
  assign s_csamul_cla32_and10_30 = a[10] & b[30];
  assign s_csamul_cla32_fa10_30_xor0 = s_csamul_cla32_and10_30 ^ s_csamul_cla32_fa11_29_xor1;
  assign s_csamul_cla32_fa10_30_and0 = s_csamul_cla32_and10_30 & s_csamul_cla32_fa11_29_xor1;
  assign s_csamul_cla32_fa10_30_xor1 = s_csamul_cla32_fa10_30_xor0 ^ s_csamul_cla32_fa10_29_or0;
  assign s_csamul_cla32_fa10_30_and1 = s_csamul_cla32_fa10_30_xor0 & s_csamul_cla32_fa10_29_or0;
  assign s_csamul_cla32_fa10_30_or0 = s_csamul_cla32_fa10_30_and0 | s_csamul_cla32_fa10_30_and1;
  assign s_csamul_cla32_and11_30 = a[11] & b[30];
  assign s_csamul_cla32_fa11_30_xor0 = s_csamul_cla32_and11_30 ^ s_csamul_cla32_fa12_29_xor1;
  assign s_csamul_cla32_fa11_30_and0 = s_csamul_cla32_and11_30 & s_csamul_cla32_fa12_29_xor1;
  assign s_csamul_cla32_fa11_30_xor1 = s_csamul_cla32_fa11_30_xor0 ^ s_csamul_cla32_fa11_29_or0;
  assign s_csamul_cla32_fa11_30_and1 = s_csamul_cla32_fa11_30_xor0 & s_csamul_cla32_fa11_29_or0;
  assign s_csamul_cla32_fa11_30_or0 = s_csamul_cla32_fa11_30_and0 | s_csamul_cla32_fa11_30_and1;
  assign s_csamul_cla32_and12_30 = a[12] & b[30];
  assign s_csamul_cla32_fa12_30_xor0 = s_csamul_cla32_and12_30 ^ s_csamul_cla32_fa13_29_xor1;
  assign s_csamul_cla32_fa12_30_and0 = s_csamul_cla32_and12_30 & s_csamul_cla32_fa13_29_xor1;
  assign s_csamul_cla32_fa12_30_xor1 = s_csamul_cla32_fa12_30_xor0 ^ s_csamul_cla32_fa12_29_or0;
  assign s_csamul_cla32_fa12_30_and1 = s_csamul_cla32_fa12_30_xor0 & s_csamul_cla32_fa12_29_or0;
  assign s_csamul_cla32_fa12_30_or0 = s_csamul_cla32_fa12_30_and0 | s_csamul_cla32_fa12_30_and1;
  assign s_csamul_cla32_and13_30 = a[13] & b[30];
  assign s_csamul_cla32_fa13_30_xor0 = s_csamul_cla32_and13_30 ^ s_csamul_cla32_fa14_29_xor1;
  assign s_csamul_cla32_fa13_30_and0 = s_csamul_cla32_and13_30 & s_csamul_cla32_fa14_29_xor1;
  assign s_csamul_cla32_fa13_30_xor1 = s_csamul_cla32_fa13_30_xor0 ^ s_csamul_cla32_fa13_29_or0;
  assign s_csamul_cla32_fa13_30_and1 = s_csamul_cla32_fa13_30_xor0 & s_csamul_cla32_fa13_29_or0;
  assign s_csamul_cla32_fa13_30_or0 = s_csamul_cla32_fa13_30_and0 | s_csamul_cla32_fa13_30_and1;
  assign s_csamul_cla32_and14_30 = a[14] & b[30];
  assign s_csamul_cla32_fa14_30_xor0 = s_csamul_cla32_and14_30 ^ s_csamul_cla32_fa15_29_xor1;
  assign s_csamul_cla32_fa14_30_and0 = s_csamul_cla32_and14_30 & s_csamul_cla32_fa15_29_xor1;
  assign s_csamul_cla32_fa14_30_xor1 = s_csamul_cla32_fa14_30_xor0 ^ s_csamul_cla32_fa14_29_or0;
  assign s_csamul_cla32_fa14_30_and1 = s_csamul_cla32_fa14_30_xor0 & s_csamul_cla32_fa14_29_or0;
  assign s_csamul_cla32_fa14_30_or0 = s_csamul_cla32_fa14_30_and0 | s_csamul_cla32_fa14_30_and1;
  assign s_csamul_cla32_and15_30 = a[15] & b[30];
  assign s_csamul_cla32_fa15_30_xor0 = s_csamul_cla32_and15_30 ^ s_csamul_cla32_fa16_29_xor1;
  assign s_csamul_cla32_fa15_30_and0 = s_csamul_cla32_and15_30 & s_csamul_cla32_fa16_29_xor1;
  assign s_csamul_cla32_fa15_30_xor1 = s_csamul_cla32_fa15_30_xor0 ^ s_csamul_cla32_fa15_29_or0;
  assign s_csamul_cla32_fa15_30_and1 = s_csamul_cla32_fa15_30_xor0 & s_csamul_cla32_fa15_29_or0;
  assign s_csamul_cla32_fa15_30_or0 = s_csamul_cla32_fa15_30_and0 | s_csamul_cla32_fa15_30_and1;
  assign s_csamul_cla32_and16_30 = a[16] & b[30];
  assign s_csamul_cla32_fa16_30_xor0 = s_csamul_cla32_and16_30 ^ s_csamul_cla32_fa17_29_xor1;
  assign s_csamul_cla32_fa16_30_and0 = s_csamul_cla32_and16_30 & s_csamul_cla32_fa17_29_xor1;
  assign s_csamul_cla32_fa16_30_xor1 = s_csamul_cla32_fa16_30_xor0 ^ s_csamul_cla32_fa16_29_or0;
  assign s_csamul_cla32_fa16_30_and1 = s_csamul_cla32_fa16_30_xor0 & s_csamul_cla32_fa16_29_or0;
  assign s_csamul_cla32_fa16_30_or0 = s_csamul_cla32_fa16_30_and0 | s_csamul_cla32_fa16_30_and1;
  assign s_csamul_cla32_and17_30 = a[17] & b[30];
  assign s_csamul_cla32_fa17_30_xor0 = s_csamul_cla32_and17_30 ^ s_csamul_cla32_fa18_29_xor1;
  assign s_csamul_cla32_fa17_30_and0 = s_csamul_cla32_and17_30 & s_csamul_cla32_fa18_29_xor1;
  assign s_csamul_cla32_fa17_30_xor1 = s_csamul_cla32_fa17_30_xor0 ^ s_csamul_cla32_fa17_29_or0;
  assign s_csamul_cla32_fa17_30_and1 = s_csamul_cla32_fa17_30_xor0 & s_csamul_cla32_fa17_29_or0;
  assign s_csamul_cla32_fa17_30_or0 = s_csamul_cla32_fa17_30_and0 | s_csamul_cla32_fa17_30_and1;
  assign s_csamul_cla32_and18_30 = a[18] & b[30];
  assign s_csamul_cla32_fa18_30_xor0 = s_csamul_cla32_and18_30 ^ s_csamul_cla32_fa19_29_xor1;
  assign s_csamul_cla32_fa18_30_and0 = s_csamul_cla32_and18_30 & s_csamul_cla32_fa19_29_xor1;
  assign s_csamul_cla32_fa18_30_xor1 = s_csamul_cla32_fa18_30_xor0 ^ s_csamul_cla32_fa18_29_or0;
  assign s_csamul_cla32_fa18_30_and1 = s_csamul_cla32_fa18_30_xor0 & s_csamul_cla32_fa18_29_or0;
  assign s_csamul_cla32_fa18_30_or0 = s_csamul_cla32_fa18_30_and0 | s_csamul_cla32_fa18_30_and1;
  assign s_csamul_cla32_and19_30 = a[19] & b[30];
  assign s_csamul_cla32_fa19_30_xor0 = s_csamul_cla32_and19_30 ^ s_csamul_cla32_fa20_29_xor1;
  assign s_csamul_cla32_fa19_30_and0 = s_csamul_cla32_and19_30 & s_csamul_cla32_fa20_29_xor1;
  assign s_csamul_cla32_fa19_30_xor1 = s_csamul_cla32_fa19_30_xor0 ^ s_csamul_cla32_fa19_29_or0;
  assign s_csamul_cla32_fa19_30_and1 = s_csamul_cla32_fa19_30_xor0 & s_csamul_cla32_fa19_29_or0;
  assign s_csamul_cla32_fa19_30_or0 = s_csamul_cla32_fa19_30_and0 | s_csamul_cla32_fa19_30_and1;
  assign s_csamul_cla32_and20_30 = a[20] & b[30];
  assign s_csamul_cla32_fa20_30_xor0 = s_csamul_cla32_and20_30 ^ s_csamul_cla32_fa21_29_xor1;
  assign s_csamul_cla32_fa20_30_and0 = s_csamul_cla32_and20_30 & s_csamul_cla32_fa21_29_xor1;
  assign s_csamul_cla32_fa20_30_xor1 = s_csamul_cla32_fa20_30_xor0 ^ s_csamul_cla32_fa20_29_or0;
  assign s_csamul_cla32_fa20_30_and1 = s_csamul_cla32_fa20_30_xor0 & s_csamul_cla32_fa20_29_or0;
  assign s_csamul_cla32_fa20_30_or0 = s_csamul_cla32_fa20_30_and0 | s_csamul_cla32_fa20_30_and1;
  assign s_csamul_cla32_and21_30 = a[21] & b[30];
  assign s_csamul_cla32_fa21_30_xor0 = s_csamul_cla32_and21_30 ^ s_csamul_cla32_fa22_29_xor1;
  assign s_csamul_cla32_fa21_30_and0 = s_csamul_cla32_and21_30 & s_csamul_cla32_fa22_29_xor1;
  assign s_csamul_cla32_fa21_30_xor1 = s_csamul_cla32_fa21_30_xor0 ^ s_csamul_cla32_fa21_29_or0;
  assign s_csamul_cla32_fa21_30_and1 = s_csamul_cla32_fa21_30_xor0 & s_csamul_cla32_fa21_29_or0;
  assign s_csamul_cla32_fa21_30_or0 = s_csamul_cla32_fa21_30_and0 | s_csamul_cla32_fa21_30_and1;
  assign s_csamul_cla32_and22_30 = a[22] & b[30];
  assign s_csamul_cla32_fa22_30_xor0 = s_csamul_cla32_and22_30 ^ s_csamul_cla32_fa23_29_xor1;
  assign s_csamul_cla32_fa22_30_and0 = s_csamul_cla32_and22_30 & s_csamul_cla32_fa23_29_xor1;
  assign s_csamul_cla32_fa22_30_xor1 = s_csamul_cla32_fa22_30_xor0 ^ s_csamul_cla32_fa22_29_or0;
  assign s_csamul_cla32_fa22_30_and1 = s_csamul_cla32_fa22_30_xor0 & s_csamul_cla32_fa22_29_or0;
  assign s_csamul_cla32_fa22_30_or0 = s_csamul_cla32_fa22_30_and0 | s_csamul_cla32_fa22_30_and1;
  assign s_csamul_cla32_and23_30 = a[23] & b[30];
  assign s_csamul_cla32_fa23_30_xor0 = s_csamul_cla32_and23_30 ^ s_csamul_cla32_fa24_29_xor1;
  assign s_csamul_cla32_fa23_30_and0 = s_csamul_cla32_and23_30 & s_csamul_cla32_fa24_29_xor1;
  assign s_csamul_cla32_fa23_30_xor1 = s_csamul_cla32_fa23_30_xor0 ^ s_csamul_cla32_fa23_29_or0;
  assign s_csamul_cla32_fa23_30_and1 = s_csamul_cla32_fa23_30_xor0 & s_csamul_cla32_fa23_29_or0;
  assign s_csamul_cla32_fa23_30_or0 = s_csamul_cla32_fa23_30_and0 | s_csamul_cla32_fa23_30_and1;
  assign s_csamul_cla32_and24_30 = a[24] & b[30];
  assign s_csamul_cla32_fa24_30_xor0 = s_csamul_cla32_and24_30 ^ s_csamul_cla32_fa25_29_xor1;
  assign s_csamul_cla32_fa24_30_and0 = s_csamul_cla32_and24_30 & s_csamul_cla32_fa25_29_xor1;
  assign s_csamul_cla32_fa24_30_xor1 = s_csamul_cla32_fa24_30_xor0 ^ s_csamul_cla32_fa24_29_or0;
  assign s_csamul_cla32_fa24_30_and1 = s_csamul_cla32_fa24_30_xor0 & s_csamul_cla32_fa24_29_or0;
  assign s_csamul_cla32_fa24_30_or0 = s_csamul_cla32_fa24_30_and0 | s_csamul_cla32_fa24_30_and1;
  assign s_csamul_cla32_and25_30 = a[25] & b[30];
  assign s_csamul_cla32_fa25_30_xor0 = s_csamul_cla32_and25_30 ^ s_csamul_cla32_fa26_29_xor1;
  assign s_csamul_cla32_fa25_30_and0 = s_csamul_cla32_and25_30 & s_csamul_cla32_fa26_29_xor1;
  assign s_csamul_cla32_fa25_30_xor1 = s_csamul_cla32_fa25_30_xor0 ^ s_csamul_cla32_fa25_29_or0;
  assign s_csamul_cla32_fa25_30_and1 = s_csamul_cla32_fa25_30_xor0 & s_csamul_cla32_fa25_29_or0;
  assign s_csamul_cla32_fa25_30_or0 = s_csamul_cla32_fa25_30_and0 | s_csamul_cla32_fa25_30_and1;
  assign s_csamul_cla32_and26_30 = a[26] & b[30];
  assign s_csamul_cla32_fa26_30_xor0 = s_csamul_cla32_and26_30 ^ s_csamul_cla32_fa27_29_xor1;
  assign s_csamul_cla32_fa26_30_and0 = s_csamul_cla32_and26_30 & s_csamul_cla32_fa27_29_xor1;
  assign s_csamul_cla32_fa26_30_xor1 = s_csamul_cla32_fa26_30_xor0 ^ s_csamul_cla32_fa26_29_or0;
  assign s_csamul_cla32_fa26_30_and1 = s_csamul_cla32_fa26_30_xor0 & s_csamul_cla32_fa26_29_or0;
  assign s_csamul_cla32_fa26_30_or0 = s_csamul_cla32_fa26_30_and0 | s_csamul_cla32_fa26_30_and1;
  assign s_csamul_cla32_and27_30 = a[27] & b[30];
  assign s_csamul_cla32_fa27_30_xor0 = s_csamul_cla32_and27_30 ^ s_csamul_cla32_fa28_29_xor1;
  assign s_csamul_cla32_fa27_30_and0 = s_csamul_cla32_and27_30 & s_csamul_cla32_fa28_29_xor1;
  assign s_csamul_cla32_fa27_30_xor1 = s_csamul_cla32_fa27_30_xor0 ^ s_csamul_cla32_fa27_29_or0;
  assign s_csamul_cla32_fa27_30_and1 = s_csamul_cla32_fa27_30_xor0 & s_csamul_cla32_fa27_29_or0;
  assign s_csamul_cla32_fa27_30_or0 = s_csamul_cla32_fa27_30_and0 | s_csamul_cla32_fa27_30_and1;
  assign s_csamul_cla32_and28_30 = a[28] & b[30];
  assign s_csamul_cla32_fa28_30_xor0 = s_csamul_cla32_and28_30 ^ s_csamul_cla32_fa29_29_xor1;
  assign s_csamul_cla32_fa28_30_and0 = s_csamul_cla32_and28_30 & s_csamul_cla32_fa29_29_xor1;
  assign s_csamul_cla32_fa28_30_xor1 = s_csamul_cla32_fa28_30_xor0 ^ s_csamul_cla32_fa28_29_or0;
  assign s_csamul_cla32_fa28_30_and1 = s_csamul_cla32_fa28_30_xor0 & s_csamul_cla32_fa28_29_or0;
  assign s_csamul_cla32_fa28_30_or0 = s_csamul_cla32_fa28_30_and0 | s_csamul_cla32_fa28_30_and1;
  assign s_csamul_cla32_and29_30 = a[29] & b[30];
  assign s_csamul_cla32_fa29_30_xor0 = s_csamul_cla32_and29_30 ^ s_csamul_cla32_fa30_29_xor1;
  assign s_csamul_cla32_fa29_30_and0 = s_csamul_cla32_and29_30 & s_csamul_cla32_fa30_29_xor1;
  assign s_csamul_cla32_fa29_30_xor1 = s_csamul_cla32_fa29_30_xor0 ^ s_csamul_cla32_fa29_29_or0;
  assign s_csamul_cla32_fa29_30_and1 = s_csamul_cla32_fa29_30_xor0 & s_csamul_cla32_fa29_29_or0;
  assign s_csamul_cla32_fa29_30_or0 = s_csamul_cla32_fa29_30_and0 | s_csamul_cla32_fa29_30_and1;
  assign s_csamul_cla32_and30_30 = a[30] & b[30];
  assign s_csamul_cla32_fa30_30_xor0 = s_csamul_cla32_and30_30 ^ s_csamul_cla32_ha31_29_xor0;
  assign s_csamul_cla32_fa30_30_and0 = s_csamul_cla32_and30_30 & s_csamul_cla32_ha31_29_xor0;
  assign s_csamul_cla32_fa30_30_xor1 = s_csamul_cla32_fa30_30_xor0 ^ s_csamul_cla32_fa30_29_or0;
  assign s_csamul_cla32_fa30_30_and1 = s_csamul_cla32_fa30_30_xor0 & s_csamul_cla32_fa30_29_or0;
  assign s_csamul_cla32_fa30_30_or0 = s_csamul_cla32_fa30_30_and0 | s_csamul_cla32_fa30_30_and1;
  assign s_csamul_cla32_nand31_30 = ~(a[31] & b[30]);
  assign s_csamul_cla32_ha31_30_xor0 = s_csamul_cla32_nand31_30 ^ s_csamul_cla32_ha31_29_and0;
  assign s_csamul_cla32_ha31_30_and0 = s_csamul_cla32_nand31_30 & s_csamul_cla32_ha31_29_and0;
  assign s_csamul_cla32_nand0_31 = ~(a[0] & b[31]);
  assign s_csamul_cla32_fa0_31_xor0 = s_csamul_cla32_nand0_31 ^ s_csamul_cla32_fa1_30_xor1;
  assign s_csamul_cla32_fa0_31_and0 = s_csamul_cla32_nand0_31 & s_csamul_cla32_fa1_30_xor1;
  assign s_csamul_cla32_fa0_31_xor1 = s_csamul_cla32_fa0_31_xor0 ^ s_csamul_cla32_fa0_30_or0;
  assign s_csamul_cla32_fa0_31_and1 = s_csamul_cla32_fa0_31_xor0 & s_csamul_cla32_fa0_30_or0;
  assign s_csamul_cla32_fa0_31_or0 = s_csamul_cla32_fa0_31_and0 | s_csamul_cla32_fa0_31_and1;
  assign s_csamul_cla32_nand1_31 = ~(a[1] & b[31]);
  assign s_csamul_cla32_fa1_31_xor0 = s_csamul_cla32_nand1_31 ^ s_csamul_cla32_fa2_30_xor1;
  assign s_csamul_cla32_fa1_31_and0 = s_csamul_cla32_nand1_31 & s_csamul_cla32_fa2_30_xor1;
  assign s_csamul_cla32_fa1_31_xor1 = s_csamul_cla32_fa1_31_xor0 ^ s_csamul_cla32_fa1_30_or0;
  assign s_csamul_cla32_fa1_31_and1 = s_csamul_cla32_fa1_31_xor0 & s_csamul_cla32_fa1_30_or0;
  assign s_csamul_cla32_fa1_31_or0 = s_csamul_cla32_fa1_31_and0 | s_csamul_cla32_fa1_31_and1;
  assign s_csamul_cla32_nand2_31 = ~(a[2] & b[31]);
  assign s_csamul_cla32_fa2_31_xor0 = s_csamul_cla32_nand2_31 ^ s_csamul_cla32_fa3_30_xor1;
  assign s_csamul_cla32_fa2_31_and0 = s_csamul_cla32_nand2_31 & s_csamul_cla32_fa3_30_xor1;
  assign s_csamul_cla32_fa2_31_xor1 = s_csamul_cla32_fa2_31_xor0 ^ s_csamul_cla32_fa2_30_or0;
  assign s_csamul_cla32_fa2_31_and1 = s_csamul_cla32_fa2_31_xor0 & s_csamul_cla32_fa2_30_or0;
  assign s_csamul_cla32_fa2_31_or0 = s_csamul_cla32_fa2_31_and0 | s_csamul_cla32_fa2_31_and1;
  assign s_csamul_cla32_nand3_31 = ~(a[3] & b[31]);
  assign s_csamul_cla32_fa3_31_xor0 = s_csamul_cla32_nand3_31 ^ s_csamul_cla32_fa4_30_xor1;
  assign s_csamul_cla32_fa3_31_and0 = s_csamul_cla32_nand3_31 & s_csamul_cla32_fa4_30_xor1;
  assign s_csamul_cla32_fa3_31_xor1 = s_csamul_cla32_fa3_31_xor0 ^ s_csamul_cla32_fa3_30_or0;
  assign s_csamul_cla32_fa3_31_and1 = s_csamul_cla32_fa3_31_xor0 & s_csamul_cla32_fa3_30_or0;
  assign s_csamul_cla32_fa3_31_or0 = s_csamul_cla32_fa3_31_and0 | s_csamul_cla32_fa3_31_and1;
  assign s_csamul_cla32_nand4_31 = ~(a[4] & b[31]);
  assign s_csamul_cla32_fa4_31_xor0 = s_csamul_cla32_nand4_31 ^ s_csamul_cla32_fa5_30_xor1;
  assign s_csamul_cla32_fa4_31_and0 = s_csamul_cla32_nand4_31 & s_csamul_cla32_fa5_30_xor1;
  assign s_csamul_cla32_fa4_31_xor1 = s_csamul_cla32_fa4_31_xor0 ^ s_csamul_cla32_fa4_30_or0;
  assign s_csamul_cla32_fa4_31_and1 = s_csamul_cla32_fa4_31_xor0 & s_csamul_cla32_fa4_30_or0;
  assign s_csamul_cla32_fa4_31_or0 = s_csamul_cla32_fa4_31_and0 | s_csamul_cla32_fa4_31_and1;
  assign s_csamul_cla32_nand5_31 = ~(a[5] & b[31]);
  assign s_csamul_cla32_fa5_31_xor0 = s_csamul_cla32_nand5_31 ^ s_csamul_cla32_fa6_30_xor1;
  assign s_csamul_cla32_fa5_31_and0 = s_csamul_cla32_nand5_31 & s_csamul_cla32_fa6_30_xor1;
  assign s_csamul_cla32_fa5_31_xor1 = s_csamul_cla32_fa5_31_xor0 ^ s_csamul_cla32_fa5_30_or0;
  assign s_csamul_cla32_fa5_31_and1 = s_csamul_cla32_fa5_31_xor0 & s_csamul_cla32_fa5_30_or0;
  assign s_csamul_cla32_fa5_31_or0 = s_csamul_cla32_fa5_31_and0 | s_csamul_cla32_fa5_31_and1;
  assign s_csamul_cla32_nand6_31 = ~(a[6] & b[31]);
  assign s_csamul_cla32_fa6_31_xor0 = s_csamul_cla32_nand6_31 ^ s_csamul_cla32_fa7_30_xor1;
  assign s_csamul_cla32_fa6_31_and0 = s_csamul_cla32_nand6_31 & s_csamul_cla32_fa7_30_xor1;
  assign s_csamul_cla32_fa6_31_xor1 = s_csamul_cla32_fa6_31_xor0 ^ s_csamul_cla32_fa6_30_or0;
  assign s_csamul_cla32_fa6_31_and1 = s_csamul_cla32_fa6_31_xor0 & s_csamul_cla32_fa6_30_or0;
  assign s_csamul_cla32_fa6_31_or0 = s_csamul_cla32_fa6_31_and0 | s_csamul_cla32_fa6_31_and1;
  assign s_csamul_cla32_nand7_31 = ~(a[7] & b[31]);
  assign s_csamul_cla32_fa7_31_xor0 = s_csamul_cla32_nand7_31 ^ s_csamul_cla32_fa8_30_xor1;
  assign s_csamul_cla32_fa7_31_and0 = s_csamul_cla32_nand7_31 & s_csamul_cla32_fa8_30_xor1;
  assign s_csamul_cla32_fa7_31_xor1 = s_csamul_cla32_fa7_31_xor0 ^ s_csamul_cla32_fa7_30_or0;
  assign s_csamul_cla32_fa7_31_and1 = s_csamul_cla32_fa7_31_xor0 & s_csamul_cla32_fa7_30_or0;
  assign s_csamul_cla32_fa7_31_or0 = s_csamul_cla32_fa7_31_and0 | s_csamul_cla32_fa7_31_and1;
  assign s_csamul_cla32_nand8_31 = ~(a[8] & b[31]);
  assign s_csamul_cla32_fa8_31_xor0 = s_csamul_cla32_nand8_31 ^ s_csamul_cla32_fa9_30_xor1;
  assign s_csamul_cla32_fa8_31_and0 = s_csamul_cla32_nand8_31 & s_csamul_cla32_fa9_30_xor1;
  assign s_csamul_cla32_fa8_31_xor1 = s_csamul_cla32_fa8_31_xor0 ^ s_csamul_cla32_fa8_30_or0;
  assign s_csamul_cla32_fa8_31_and1 = s_csamul_cla32_fa8_31_xor0 & s_csamul_cla32_fa8_30_or0;
  assign s_csamul_cla32_fa8_31_or0 = s_csamul_cla32_fa8_31_and0 | s_csamul_cla32_fa8_31_and1;
  assign s_csamul_cla32_nand9_31 = ~(a[9] & b[31]);
  assign s_csamul_cla32_fa9_31_xor0 = s_csamul_cla32_nand9_31 ^ s_csamul_cla32_fa10_30_xor1;
  assign s_csamul_cla32_fa9_31_and0 = s_csamul_cla32_nand9_31 & s_csamul_cla32_fa10_30_xor1;
  assign s_csamul_cla32_fa9_31_xor1 = s_csamul_cla32_fa9_31_xor0 ^ s_csamul_cla32_fa9_30_or0;
  assign s_csamul_cla32_fa9_31_and1 = s_csamul_cla32_fa9_31_xor0 & s_csamul_cla32_fa9_30_or0;
  assign s_csamul_cla32_fa9_31_or0 = s_csamul_cla32_fa9_31_and0 | s_csamul_cla32_fa9_31_and1;
  assign s_csamul_cla32_nand10_31 = ~(a[10] & b[31]);
  assign s_csamul_cla32_fa10_31_xor0 = s_csamul_cla32_nand10_31 ^ s_csamul_cla32_fa11_30_xor1;
  assign s_csamul_cla32_fa10_31_and0 = s_csamul_cla32_nand10_31 & s_csamul_cla32_fa11_30_xor1;
  assign s_csamul_cla32_fa10_31_xor1 = s_csamul_cla32_fa10_31_xor0 ^ s_csamul_cla32_fa10_30_or0;
  assign s_csamul_cla32_fa10_31_and1 = s_csamul_cla32_fa10_31_xor0 & s_csamul_cla32_fa10_30_or0;
  assign s_csamul_cla32_fa10_31_or0 = s_csamul_cla32_fa10_31_and0 | s_csamul_cla32_fa10_31_and1;
  assign s_csamul_cla32_nand11_31 = ~(a[11] & b[31]);
  assign s_csamul_cla32_fa11_31_xor0 = s_csamul_cla32_nand11_31 ^ s_csamul_cla32_fa12_30_xor1;
  assign s_csamul_cla32_fa11_31_and0 = s_csamul_cla32_nand11_31 & s_csamul_cla32_fa12_30_xor1;
  assign s_csamul_cla32_fa11_31_xor1 = s_csamul_cla32_fa11_31_xor0 ^ s_csamul_cla32_fa11_30_or0;
  assign s_csamul_cla32_fa11_31_and1 = s_csamul_cla32_fa11_31_xor0 & s_csamul_cla32_fa11_30_or0;
  assign s_csamul_cla32_fa11_31_or0 = s_csamul_cla32_fa11_31_and0 | s_csamul_cla32_fa11_31_and1;
  assign s_csamul_cla32_nand12_31 = ~(a[12] & b[31]);
  assign s_csamul_cla32_fa12_31_xor0 = s_csamul_cla32_nand12_31 ^ s_csamul_cla32_fa13_30_xor1;
  assign s_csamul_cla32_fa12_31_and0 = s_csamul_cla32_nand12_31 & s_csamul_cla32_fa13_30_xor1;
  assign s_csamul_cla32_fa12_31_xor1 = s_csamul_cla32_fa12_31_xor0 ^ s_csamul_cla32_fa12_30_or0;
  assign s_csamul_cla32_fa12_31_and1 = s_csamul_cla32_fa12_31_xor0 & s_csamul_cla32_fa12_30_or0;
  assign s_csamul_cla32_fa12_31_or0 = s_csamul_cla32_fa12_31_and0 | s_csamul_cla32_fa12_31_and1;
  assign s_csamul_cla32_nand13_31 = ~(a[13] & b[31]);
  assign s_csamul_cla32_fa13_31_xor0 = s_csamul_cla32_nand13_31 ^ s_csamul_cla32_fa14_30_xor1;
  assign s_csamul_cla32_fa13_31_and0 = s_csamul_cla32_nand13_31 & s_csamul_cla32_fa14_30_xor1;
  assign s_csamul_cla32_fa13_31_xor1 = s_csamul_cla32_fa13_31_xor0 ^ s_csamul_cla32_fa13_30_or0;
  assign s_csamul_cla32_fa13_31_and1 = s_csamul_cla32_fa13_31_xor0 & s_csamul_cla32_fa13_30_or0;
  assign s_csamul_cla32_fa13_31_or0 = s_csamul_cla32_fa13_31_and0 | s_csamul_cla32_fa13_31_and1;
  assign s_csamul_cla32_nand14_31 = ~(a[14] & b[31]);
  assign s_csamul_cla32_fa14_31_xor0 = s_csamul_cla32_nand14_31 ^ s_csamul_cla32_fa15_30_xor1;
  assign s_csamul_cla32_fa14_31_and0 = s_csamul_cla32_nand14_31 & s_csamul_cla32_fa15_30_xor1;
  assign s_csamul_cla32_fa14_31_xor1 = s_csamul_cla32_fa14_31_xor0 ^ s_csamul_cla32_fa14_30_or0;
  assign s_csamul_cla32_fa14_31_and1 = s_csamul_cla32_fa14_31_xor0 & s_csamul_cla32_fa14_30_or0;
  assign s_csamul_cla32_fa14_31_or0 = s_csamul_cla32_fa14_31_and0 | s_csamul_cla32_fa14_31_and1;
  assign s_csamul_cla32_nand15_31 = ~(a[15] & b[31]);
  assign s_csamul_cla32_fa15_31_xor0 = s_csamul_cla32_nand15_31 ^ s_csamul_cla32_fa16_30_xor1;
  assign s_csamul_cla32_fa15_31_and0 = s_csamul_cla32_nand15_31 & s_csamul_cla32_fa16_30_xor1;
  assign s_csamul_cla32_fa15_31_xor1 = s_csamul_cla32_fa15_31_xor0 ^ s_csamul_cla32_fa15_30_or0;
  assign s_csamul_cla32_fa15_31_and1 = s_csamul_cla32_fa15_31_xor0 & s_csamul_cla32_fa15_30_or0;
  assign s_csamul_cla32_fa15_31_or0 = s_csamul_cla32_fa15_31_and0 | s_csamul_cla32_fa15_31_and1;
  assign s_csamul_cla32_nand16_31 = ~(a[16] & b[31]);
  assign s_csamul_cla32_fa16_31_xor0 = s_csamul_cla32_nand16_31 ^ s_csamul_cla32_fa17_30_xor1;
  assign s_csamul_cla32_fa16_31_and0 = s_csamul_cla32_nand16_31 & s_csamul_cla32_fa17_30_xor1;
  assign s_csamul_cla32_fa16_31_xor1 = s_csamul_cla32_fa16_31_xor0 ^ s_csamul_cla32_fa16_30_or0;
  assign s_csamul_cla32_fa16_31_and1 = s_csamul_cla32_fa16_31_xor0 & s_csamul_cla32_fa16_30_or0;
  assign s_csamul_cla32_fa16_31_or0 = s_csamul_cla32_fa16_31_and0 | s_csamul_cla32_fa16_31_and1;
  assign s_csamul_cla32_nand17_31 = ~(a[17] & b[31]);
  assign s_csamul_cla32_fa17_31_xor0 = s_csamul_cla32_nand17_31 ^ s_csamul_cla32_fa18_30_xor1;
  assign s_csamul_cla32_fa17_31_and0 = s_csamul_cla32_nand17_31 & s_csamul_cla32_fa18_30_xor1;
  assign s_csamul_cla32_fa17_31_xor1 = s_csamul_cla32_fa17_31_xor0 ^ s_csamul_cla32_fa17_30_or0;
  assign s_csamul_cla32_fa17_31_and1 = s_csamul_cla32_fa17_31_xor0 & s_csamul_cla32_fa17_30_or0;
  assign s_csamul_cla32_fa17_31_or0 = s_csamul_cla32_fa17_31_and0 | s_csamul_cla32_fa17_31_and1;
  assign s_csamul_cla32_nand18_31 = ~(a[18] & b[31]);
  assign s_csamul_cla32_fa18_31_xor0 = s_csamul_cla32_nand18_31 ^ s_csamul_cla32_fa19_30_xor1;
  assign s_csamul_cla32_fa18_31_and0 = s_csamul_cla32_nand18_31 & s_csamul_cla32_fa19_30_xor1;
  assign s_csamul_cla32_fa18_31_xor1 = s_csamul_cla32_fa18_31_xor0 ^ s_csamul_cla32_fa18_30_or0;
  assign s_csamul_cla32_fa18_31_and1 = s_csamul_cla32_fa18_31_xor0 & s_csamul_cla32_fa18_30_or0;
  assign s_csamul_cla32_fa18_31_or0 = s_csamul_cla32_fa18_31_and0 | s_csamul_cla32_fa18_31_and1;
  assign s_csamul_cla32_nand19_31 = ~(a[19] & b[31]);
  assign s_csamul_cla32_fa19_31_xor0 = s_csamul_cla32_nand19_31 ^ s_csamul_cla32_fa20_30_xor1;
  assign s_csamul_cla32_fa19_31_and0 = s_csamul_cla32_nand19_31 & s_csamul_cla32_fa20_30_xor1;
  assign s_csamul_cla32_fa19_31_xor1 = s_csamul_cla32_fa19_31_xor0 ^ s_csamul_cla32_fa19_30_or0;
  assign s_csamul_cla32_fa19_31_and1 = s_csamul_cla32_fa19_31_xor0 & s_csamul_cla32_fa19_30_or0;
  assign s_csamul_cla32_fa19_31_or0 = s_csamul_cla32_fa19_31_and0 | s_csamul_cla32_fa19_31_and1;
  assign s_csamul_cla32_nand20_31 = ~(a[20] & b[31]);
  assign s_csamul_cla32_fa20_31_xor0 = s_csamul_cla32_nand20_31 ^ s_csamul_cla32_fa21_30_xor1;
  assign s_csamul_cla32_fa20_31_and0 = s_csamul_cla32_nand20_31 & s_csamul_cla32_fa21_30_xor1;
  assign s_csamul_cla32_fa20_31_xor1 = s_csamul_cla32_fa20_31_xor0 ^ s_csamul_cla32_fa20_30_or0;
  assign s_csamul_cla32_fa20_31_and1 = s_csamul_cla32_fa20_31_xor0 & s_csamul_cla32_fa20_30_or0;
  assign s_csamul_cla32_fa20_31_or0 = s_csamul_cla32_fa20_31_and0 | s_csamul_cla32_fa20_31_and1;
  assign s_csamul_cla32_nand21_31 = ~(a[21] & b[31]);
  assign s_csamul_cla32_fa21_31_xor0 = s_csamul_cla32_nand21_31 ^ s_csamul_cla32_fa22_30_xor1;
  assign s_csamul_cla32_fa21_31_and0 = s_csamul_cla32_nand21_31 & s_csamul_cla32_fa22_30_xor1;
  assign s_csamul_cla32_fa21_31_xor1 = s_csamul_cla32_fa21_31_xor0 ^ s_csamul_cla32_fa21_30_or0;
  assign s_csamul_cla32_fa21_31_and1 = s_csamul_cla32_fa21_31_xor0 & s_csamul_cla32_fa21_30_or0;
  assign s_csamul_cla32_fa21_31_or0 = s_csamul_cla32_fa21_31_and0 | s_csamul_cla32_fa21_31_and1;
  assign s_csamul_cla32_nand22_31 = ~(a[22] & b[31]);
  assign s_csamul_cla32_fa22_31_xor0 = s_csamul_cla32_nand22_31 ^ s_csamul_cla32_fa23_30_xor1;
  assign s_csamul_cla32_fa22_31_and0 = s_csamul_cla32_nand22_31 & s_csamul_cla32_fa23_30_xor1;
  assign s_csamul_cla32_fa22_31_xor1 = s_csamul_cla32_fa22_31_xor0 ^ s_csamul_cla32_fa22_30_or0;
  assign s_csamul_cla32_fa22_31_and1 = s_csamul_cla32_fa22_31_xor0 & s_csamul_cla32_fa22_30_or0;
  assign s_csamul_cla32_fa22_31_or0 = s_csamul_cla32_fa22_31_and0 | s_csamul_cla32_fa22_31_and1;
  assign s_csamul_cla32_nand23_31 = ~(a[23] & b[31]);
  assign s_csamul_cla32_fa23_31_xor0 = s_csamul_cla32_nand23_31 ^ s_csamul_cla32_fa24_30_xor1;
  assign s_csamul_cla32_fa23_31_and0 = s_csamul_cla32_nand23_31 & s_csamul_cla32_fa24_30_xor1;
  assign s_csamul_cla32_fa23_31_xor1 = s_csamul_cla32_fa23_31_xor0 ^ s_csamul_cla32_fa23_30_or0;
  assign s_csamul_cla32_fa23_31_and1 = s_csamul_cla32_fa23_31_xor0 & s_csamul_cla32_fa23_30_or0;
  assign s_csamul_cla32_fa23_31_or0 = s_csamul_cla32_fa23_31_and0 | s_csamul_cla32_fa23_31_and1;
  assign s_csamul_cla32_nand24_31 = ~(a[24] & b[31]);
  assign s_csamul_cla32_fa24_31_xor0 = s_csamul_cla32_nand24_31 ^ s_csamul_cla32_fa25_30_xor1;
  assign s_csamul_cla32_fa24_31_and0 = s_csamul_cla32_nand24_31 & s_csamul_cla32_fa25_30_xor1;
  assign s_csamul_cla32_fa24_31_xor1 = s_csamul_cla32_fa24_31_xor0 ^ s_csamul_cla32_fa24_30_or0;
  assign s_csamul_cla32_fa24_31_and1 = s_csamul_cla32_fa24_31_xor0 & s_csamul_cla32_fa24_30_or0;
  assign s_csamul_cla32_fa24_31_or0 = s_csamul_cla32_fa24_31_and0 | s_csamul_cla32_fa24_31_and1;
  assign s_csamul_cla32_nand25_31 = ~(a[25] & b[31]);
  assign s_csamul_cla32_fa25_31_xor0 = s_csamul_cla32_nand25_31 ^ s_csamul_cla32_fa26_30_xor1;
  assign s_csamul_cla32_fa25_31_and0 = s_csamul_cla32_nand25_31 & s_csamul_cla32_fa26_30_xor1;
  assign s_csamul_cla32_fa25_31_xor1 = s_csamul_cla32_fa25_31_xor0 ^ s_csamul_cla32_fa25_30_or0;
  assign s_csamul_cla32_fa25_31_and1 = s_csamul_cla32_fa25_31_xor0 & s_csamul_cla32_fa25_30_or0;
  assign s_csamul_cla32_fa25_31_or0 = s_csamul_cla32_fa25_31_and0 | s_csamul_cla32_fa25_31_and1;
  assign s_csamul_cla32_nand26_31 = ~(a[26] & b[31]);
  assign s_csamul_cla32_fa26_31_xor0 = s_csamul_cla32_nand26_31 ^ s_csamul_cla32_fa27_30_xor1;
  assign s_csamul_cla32_fa26_31_and0 = s_csamul_cla32_nand26_31 & s_csamul_cla32_fa27_30_xor1;
  assign s_csamul_cla32_fa26_31_xor1 = s_csamul_cla32_fa26_31_xor0 ^ s_csamul_cla32_fa26_30_or0;
  assign s_csamul_cla32_fa26_31_and1 = s_csamul_cla32_fa26_31_xor0 & s_csamul_cla32_fa26_30_or0;
  assign s_csamul_cla32_fa26_31_or0 = s_csamul_cla32_fa26_31_and0 | s_csamul_cla32_fa26_31_and1;
  assign s_csamul_cla32_nand27_31 = ~(a[27] & b[31]);
  assign s_csamul_cla32_fa27_31_xor0 = s_csamul_cla32_nand27_31 ^ s_csamul_cla32_fa28_30_xor1;
  assign s_csamul_cla32_fa27_31_and0 = s_csamul_cla32_nand27_31 & s_csamul_cla32_fa28_30_xor1;
  assign s_csamul_cla32_fa27_31_xor1 = s_csamul_cla32_fa27_31_xor0 ^ s_csamul_cla32_fa27_30_or0;
  assign s_csamul_cla32_fa27_31_and1 = s_csamul_cla32_fa27_31_xor0 & s_csamul_cla32_fa27_30_or0;
  assign s_csamul_cla32_fa27_31_or0 = s_csamul_cla32_fa27_31_and0 | s_csamul_cla32_fa27_31_and1;
  assign s_csamul_cla32_nand28_31 = ~(a[28] & b[31]);
  assign s_csamul_cla32_fa28_31_xor0 = s_csamul_cla32_nand28_31 ^ s_csamul_cla32_fa29_30_xor1;
  assign s_csamul_cla32_fa28_31_and0 = s_csamul_cla32_nand28_31 & s_csamul_cla32_fa29_30_xor1;
  assign s_csamul_cla32_fa28_31_xor1 = s_csamul_cla32_fa28_31_xor0 ^ s_csamul_cla32_fa28_30_or0;
  assign s_csamul_cla32_fa28_31_and1 = s_csamul_cla32_fa28_31_xor0 & s_csamul_cla32_fa28_30_or0;
  assign s_csamul_cla32_fa28_31_or0 = s_csamul_cla32_fa28_31_and0 | s_csamul_cla32_fa28_31_and1;
  assign s_csamul_cla32_nand29_31 = ~(a[29] & b[31]);
  assign s_csamul_cla32_fa29_31_xor0 = s_csamul_cla32_nand29_31 ^ s_csamul_cla32_fa30_30_xor1;
  assign s_csamul_cla32_fa29_31_and0 = s_csamul_cla32_nand29_31 & s_csamul_cla32_fa30_30_xor1;
  assign s_csamul_cla32_fa29_31_xor1 = s_csamul_cla32_fa29_31_xor0 ^ s_csamul_cla32_fa29_30_or0;
  assign s_csamul_cla32_fa29_31_and1 = s_csamul_cla32_fa29_31_xor0 & s_csamul_cla32_fa29_30_or0;
  assign s_csamul_cla32_fa29_31_or0 = s_csamul_cla32_fa29_31_and0 | s_csamul_cla32_fa29_31_and1;
  assign s_csamul_cla32_nand30_31 = ~(a[30] & b[31]);
  assign s_csamul_cla32_fa30_31_xor0 = s_csamul_cla32_nand30_31 ^ s_csamul_cla32_ha31_30_xor0;
  assign s_csamul_cla32_fa30_31_and0 = s_csamul_cla32_nand30_31 & s_csamul_cla32_ha31_30_xor0;
  assign s_csamul_cla32_fa30_31_xor1 = s_csamul_cla32_fa30_31_xor0 ^ s_csamul_cla32_fa30_30_or0;
  assign s_csamul_cla32_fa30_31_and1 = s_csamul_cla32_fa30_31_xor0 & s_csamul_cla32_fa30_30_or0;
  assign s_csamul_cla32_fa30_31_or0 = s_csamul_cla32_fa30_31_and0 | s_csamul_cla32_fa30_31_and1;
  assign s_csamul_cla32_and31_31 = a[31] & b[31];
  assign s_csamul_cla32_ha31_31_xor0 = s_csamul_cla32_and31_31 ^ s_csamul_cla32_ha31_30_and0;
  assign s_csamul_cla32_ha31_31_and0 = s_csamul_cla32_and31_31 & s_csamul_cla32_ha31_30_and0;
  assign s_csamul_cla32_u_cla32_pg_logic0_or0 = s_csamul_cla32_fa1_31_xor1 | s_csamul_cla32_fa0_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic0_and0 = s_csamul_cla32_fa1_31_xor1 & s_csamul_cla32_fa0_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic0_xor0 = s_csamul_cla32_fa1_31_xor1 ^ s_csamul_cla32_fa0_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic1_or0 = s_csamul_cla32_fa2_31_xor1 | s_csamul_cla32_fa1_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic1_and0 = s_csamul_cla32_fa2_31_xor1 & s_csamul_cla32_fa1_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic1_xor0 = s_csamul_cla32_fa2_31_xor1 ^ s_csamul_cla32_fa1_31_or0;
  assign s_csamul_cla32_u_cla32_xor1 = s_csamul_cla32_u_cla32_pg_logic1_xor0 ^ s_csamul_cla32_u_cla32_pg_logic0_and0;
  assign s_csamul_cla32_u_cla32_and0 = s_csamul_cla32_u_cla32_pg_logic0_and0 & s_csamul_cla32_u_cla32_pg_logic1_or0;
  assign s_csamul_cla32_u_cla32_or0 = s_csamul_cla32_u_cla32_pg_logic1_and0 | s_csamul_cla32_u_cla32_and0;
  assign s_csamul_cla32_u_cla32_pg_logic2_or0 = s_csamul_cla32_fa3_31_xor1 | s_csamul_cla32_fa2_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic2_and0 = s_csamul_cla32_fa3_31_xor1 & s_csamul_cla32_fa2_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic2_xor0 = s_csamul_cla32_fa3_31_xor1 ^ s_csamul_cla32_fa2_31_or0;
  assign s_csamul_cla32_u_cla32_xor2 = s_csamul_cla32_u_cla32_pg_logic2_xor0 ^ s_csamul_cla32_u_cla32_or0;
  assign s_csamul_cla32_u_cla32_and1 = s_csamul_cla32_u_cla32_pg_logic2_or0 & s_csamul_cla32_u_cla32_pg_logic0_or0;
  assign s_csamul_cla32_u_cla32_and2 = s_csamul_cla32_u_cla32_pg_logic0_and0 & s_csamul_cla32_u_cla32_pg_logic2_or0;
  assign s_csamul_cla32_u_cla32_and3 = s_csamul_cla32_u_cla32_and2 & s_csamul_cla32_u_cla32_pg_logic1_or0;
  assign s_csamul_cla32_u_cla32_and4 = s_csamul_cla32_u_cla32_pg_logic1_and0 & s_csamul_cla32_u_cla32_pg_logic2_or0;
  assign s_csamul_cla32_u_cla32_or1 = s_csamul_cla32_u_cla32_and3 | s_csamul_cla32_u_cla32_and4;
  assign s_csamul_cla32_u_cla32_or2 = s_csamul_cla32_u_cla32_pg_logic2_and0 | s_csamul_cla32_u_cla32_or1;
  assign s_csamul_cla32_u_cla32_pg_logic3_or0 = s_csamul_cla32_fa4_31_xor1 | s_csamul_cla32_fa3_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic3_and0 = s_csamul_cla32_fa4_31_xor1 & s_csamul_cla32_fa3_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic3_xor0 = s_csamul_cla32_fa4_31_xor1 ^ s_csamul_cla32_fa3_31_or0;
  assign s_csamul_cla32_u_cla32_xor3 = s_csamul_cla32_u_cla32_pg_logic3_xor0 ^ s_csamul_cla32_u_cla32_or2;
  assign s_csamul_cla32_u_cla32_and5 = s_csamul_cla32_u_cla32_pg_logic3_or0 & s_csamul_cla32_u_cla32_pg_logic1_or0;
  assign s_csamul_cla32_u_cla32_and6 = s_csamul_cla32_u_cla32_pg_logic0_and0 & s_csamul_cla32_u_cla32_pg_logic2_or0;
  assign s_csamul_cla32_u_cla32_and7 = s_csamul_cla32_u_cla32_pg_logic3_or0 & s_csamul_cla32_u_cla32_pg_logic1_or0;
  assign s_csamul_cla32_u_cla32_and8 = s_csamul_cla32_u_cla32_and6 & s_csamul_cla32_u_cla32_and7;
  assign s_csamul_cla32_u_cla32_and9 = s_csamul_cla32_u_cla32_pg_logic1_and0 & s_csamul_cla32_u_cla32_pg_logic3_or0;
  assign s_csamul_cla32_u_cla32_and10 = s_csamul_cla32_u_cla32_and9 & s_csamul_cla32_u_cla32_pg_logic2_or0;
  assign s_csamul_cla32_u_cla32_and11 = s_csamul_cla32_u_cla32_pg_logic2_and0 & s_csamul_cla32_u_cla32_pg_logic3_or0;
  assign s_csamul_cla32_u_cla32_or3 = s_csamul_cla32_u_cla32_and8 | s_csamul_cla32_u_cla32_and11;
  assign s_csamul_cla32_u_cla32_or4 = s_csamul_cla32_u_cla32_and10 | s_csamul_cla32_u_cla32_or3;
  assign s_csamul_cla32_u_cla32_or5 = s_csamul_cla32_u_cla32_pg_logic3_and0 | s_csamul_cla32_u_cla32_or4;
  assign s_csamul_cla32_u_cla32_pg_logic4_or0 = s_csamul_cla32_fa5_31_xor1 | s_csamul_cla32_fa4_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic4_and0 = s_csamul_cla32_fa5_31_xor1 & s_csamul_cla32_fa4_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic4_xor0 = s_csamul_cla32_fa5_31_xor1 ^ s_csamul_cla32_fa4_31_or0;
  assign s_csamul_cla32_u_cla32_xor4 = s_csamul_cla32_u_cla32_pg_logic4_xor0 ^ s_csamul_cla32_u_cla32_or5;
  assign s_csamul_cla32_u_cla32_and12 = s_csamul_cla32_u_cla32_or5 & s_csamul_cla32_u_cla32_pg_logic4_or0;
  assign s_csamul_cla32_u_cla32_or6 = s_csamul_cla32_u_cla32_pg_logic4_and0 | s_csamul_cla32_u_cla32_and12;
  assign s_csamul_cla32_u_cla32_pg_logic5_or0 = s_csamul_cla32_fa6_31_xor1 | s_csamul_cla32_fa5_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic5_and0 = s_csamul_cla32_fa6_31_xor1 & s_csamul_cla32_fa5_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic5_xor0 = s_csamul_cla32_fa6_31_xor1 ^ s_csamul_cla32_fa5_31_or0;
  assign s_csamul_cla32_u_cla32_xor5 = s_csamul_cla32_u_cla32_pg_logic5_xor0 ^ s_csamul_cla32_u_cla32_or6;
  assign s_csamul_cla32_u_cla32_and13 = s_csamul_cla32_u_cla32_or5 & s_csamul_cla32_u_cla32_pg_logic5_or0;
  assign s_csamul_cla32_u_cla32_and14 = s_csamul_cla32_u_cla32_and13 & s_csamul_cla32_u_cla32_pg_logic4_or0;
  assign s_csamul_cla32_u_cla32_and15 = s_csamul_cla32_u_cla32_pg_logic4_and0 & s_csamul_cla32_u_cla32_pg_logic5_or0;
  assign s_csamul_cla32_u_cla32_or7 = s_csamul_cla32_u_cla32_and14 | s_csamul_cla32_u_cla32_and15;
  assign s_csamul_cla32_u_cla32_or8 = s_csamul_cla32_u_cla32_pg_logic5_and0 | s_csamul_cla32_u_cla32_or7;
  assign s_csamul_cla32_u_cla32_pg_logic6_or0 = s_csamul_cla32_fa7_31_xor1 | s_csamul_cla32_fa6_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic6_and0 = s_csamul_cla32_fa7_31_xor1 & s_csamul_cla32_fa6_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic6_xor0 = s_csamul_cla32_fa7_31_xor1 ^ s_csamul_cla32_fa6_31_or0;
  assign s_csamul_cla32_u_cla32_xor6 = s_csamul_cla32_u_cla32_pg_logic6_xor0 ^ s_csamul_cla32_u_cla32_or8;
  assign s_csamul_cla32_u_cla32_and16 = s_csamul_cla32_u_cla32_or5 & s_csamul_cla32_u_cla32_pg_logic5_or0;
  assign s_csamul_cla32_u_cla32_and17 = s_csamul_cla32_u_cla32_pg_logic6_or0 & s_csamul_cla32_u_cla32_pg_logic4_or0;
  assign s_csamul_cla32_u_cla32_and18 = s_csamul_cla32_u_cla32_and16 & s_csamul_cla32_u_cla32_and17;
  assign s_csamul_cla32_u_cla32_and19 = s_csamul_cla32_u_cla32_pg_logic4_and0 & s_csamul_cla32_u_cla32_pg_logic6_or0;
  assign s_csamul_cla32_u_cla32_and20 = s_csamul_cla32_u_cla32_and19 & s_csamul_cla32_u_cla32_pg_logic5_or0;
  assign s_csamul_cla32_u_cla32_and21 = s_csamul_cla32_u_cla32_pg_logic5_and0 & s_csamul_cla32_u_cla32_pg_logic6_or0;
  assign s_csamul_cla32_u_cla32_or9 = s_csamul_cla32_u_cla32_and18 | s_csamul_cla32_u_cla32_and20;
  assign s_csamul_cla32_u_cla32_or10 = s_csamul_cla32_u_cla32_or9 | s_csamul_cla32_u_cla32_and21;
  assign s_csamul_cla32_u_cla32_or11 = s_csamul_cla32_u_cla32_pg_logic6_and0 | s_csamul_cla32_u_cla32_or10;
  assign s_csamul_cla32_u_cla32_pg_logic7_or0 = s_csamul_cla32_fa8_31_xor1 | s_csamul_cla32_fa7_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic7_and0 = s_csamul_cla32_fa8_31_xor1 & s_csamul_cla32_fa7_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic7_xor0 = s_csamul_cla32_fa8_31_xor1 ^ s_csamul_cla32_fa7_31_or0;
  assign s_csamul_cla32_u_cla32_xor7 = s_csamul_cla32_u_cla32_pg_logic7_xor0 ^ s_csamul_cla32_u_cla32_or11;
  assign s_csamul_cla32_u_cla32_and22 = s_csamul_cla32_u_cla32_or5 & s_csamul_cla32_u_cla32_pg_logic6_or0;
  assign s_csamul_cla32_u_cla32_and23 = s_csamul_cla32_u_cla32_pg_logic7_or0 & s_csamul_cla32_u_cla32_pg_logic5_or0;
  assign s_csamul_cla32_u_cla32_and24 = s_csamul_cla32_u_cla32_and22 & s_csamul_cla32_u_cla32_and23;
  assign s_csamul_cla32_u_cla32_and25 = s_csamul_cla32_u_cla32_and24 & s_csamul_cla32_u_cla32_pg_logic4_or0;
  assign s_csamul_cla32_u_cla32_and26 = s_csamul_cla32_u_cla32_pg_logic4_and0 & s_csamul_cla32_u_cla32_pg_logic6_or0;
  assign s_csamul_cla32_u_cla32_and27 = s_csamul_cla32_u_cla32_pg_logic7_or0 & s_csamul_cla32_u_cla32_pg_logic5_or0;
  assign s_csamul_cla32_u_cla32_and28 = s_csamul_cla32_u_cla32_and26 & s_csamul_cla32_u_cla32_and27;
  assign s_csamul_cla32_u_cla32_and29 = s_csamul_cla32_u_cla32_pg_logic5_and0 & s_csamul_cla32_u_cla32_pg_logic7_or0;
  assign s_csamul_cla32_u_cla32_and30 = s_csamul_cla32_u_cla32_and29 & s_csamul_cla32_u_cla32_pg_logic6_or0;
  assign s_csamul_cla32_u_cla32_and31 = s_csamul_cla32_u_cla32_pg_logic6_and0 & s_csamul_cla32_u_cla32_pg_logic7_or0;
  assign s_csamul_cla32_u_cla32_or12 = s_csamul_cla32_u_cla32_and25 | s_csamul_cla32_u_cla32_and30;
  assign s_csamul_cla32_u_cla32_or13 = s_csamul_cla32_u_cla32_and28 | s_csamul_cla32_u_cla32_and31;
  assign s_csamul_cla32_u_cla32_or14 = s_csamul_cla32_u_cla32_or12 | s_csamul_cla32_u_cla32_or13;
  assign s_csamul_cla32_u_cla32_or15 = s_csamul_cla32_u_cla32_pg_logic7_and0 | s_csamul_cla32_u_cla32_or14;
  assign s_csamul_cla32_u_cla32_pg_logic8_or0 = s_csamul_cla32_fa9_31_xor1 | s_csamul_cla32_fa8_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic8_and0 = s_csamul_cla32_fa9_31_xor1 & s_csamul_cla32_fa8_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic8_xor0 = s_csamul_cla32_fa9_31_xor1 ^ s_csamul_cla32_fa8_31_or0;
  assign s_csamul_cla32_u_cla32_xor8 = s_csamul_cla32_u_cla32_pg_logic8_xor0 ^ s_csamul_cla32_u_cla32_or15;
  assign s_csamul_cla32_u_cla32_and32 = s_csamul_cla32_u_cla32_or15 & s_csamul_cla32_u_cla32_pg_logic8_or0;
  assign s_csamul_cla32_u_cla32_or16 = s_csamul_cla32_u_cla32_pg_logic8_and0 | s_csamul_cla32_u_cla32_and32;
  assign s_csamul_cla32_u_cla32_pg_logic9_or0 = s_csamul_cla32_fa10_31_xor1 | s_csamul_cla32_fa9_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic9_and0 = s_csamul_cla32_fa10_31_xor1 & s_csamul_cla32_fa9_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic9_xor0 = s_csamul_cla32_fa10_31_xor1 ^ s_csamul_cla32_fa9_31_or0;
  assign s_csamul_cla32_u_cla32_xor9 = s_csamul_cla32_u_cla32_pg_logic9_xor0 ^ s_csamul_cla32_u_cla32_or16;
  assign s_csamul_cla32_u_cla32_and33 = s_csamul_cla32_u_cla32_or15 & s_csamul_cla32_u_cla32_pg_logic9_or0;
  assign s_csamul_cla32_u_cla32_and34 = s_csamul_cla32_u_cla32_and33 & s_csamul_cla32_u_cla32_pg_logic8_or0;
  assign s_csamul_cla32_u_cla32_and35 = s_csamul_cla32_u_cla32_pg_logic8_and0 & s_csamul_cla32_u_cla32_pg_logic9_or0;
  assign s_csamul_cla32_u_cla32_or17 = s_csamul_cla32_u_cla32_and34 | s_csamul_cla32_u_cla32_and35;
  assign s_csamul_cla32_u_cla32_or18 = s_csamul_cla32_u_cla32_pg_logic9_and0 | s_csamul_cla32_u_cla32_or17;
  assign s_csamul_cla32_u_cla32_pg_logic10_or0 = s_csamul_cla32_fa11_31_xor1 | s_csamul_cla32_fa10_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic10_and0 = s_csamul_cla32_fa11_31_xor1 & s_csamul_cla32_fa10_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic10_xor0 = s_csamul_cla32_fa11_31_xor1 ^ s_csamul_cla32_fa10_31_or0;
  assign s_csamul_cla32_u_cla32_xor10 = s_csamul_cla32_u_cla32_pg_logic10_xor0 ^ s_csamul_cla32_u_cla32_or18;
  assign s_csamul_cla32_u_cla32_and36 = s_csamul_cla32_u_cla32_or15 & s_csamul_cla32_u_cla32_pg_logic9_or0;
  assign s_csamul_cla32_u_cla32_and37 = s_csamul_cla32_u_cla32_pg_logic10_or0 & s_csamul_cla32_u_cla32_pg_logic8_or0;
  assign s_csamul_cla32_u_cla32_and38 = s_csamul_cla32_u_cla32_and36 & s_csamul_cla32_u_cla32_and37;
  assign s_csamul_cla32_u_cla32_and39 = s_csamul_cla32_u_cla32_pg_logic8_and0 & s_csamul_cla32_u_cla32_pg_logic10_or0;
  assign s_csamul_cla32_u_cla32_and40 = s_csamul_cla32_u_cla32_and39 & s_csamul_cla32_u_cla32_pg_logic9_or0;
  assign s_csamul_cla32_u_cla32_and41 = s_csamul_cla32_u_cla32_pg_logic9_and0 & s_csamul_cla32_u_cla32_pg_logic10_or0;
  assign s_csamul_cla32_u_cla32_or19 = s_csamul_cla32_u_cla32_and38 | s_csamul_cla32_u_cla32_and40;
  assign s_csamul_cla32_u_cla32_or20 = s_csamul_cla32_u_cla32_or19 | s_csamul_cla32_u_cla32_and41;
  assign s_csamul_cla32_u_cla32_or21 = s_csamul_cla32_u_cla32_pg_logic10_and0 | s_csamul_cla32_u_cla32_or20;
  assign s_csamul_cla32_u_cla32_pg_logic11_or0 = s_csamul_cla32_fa12_31_xor1 | s_csamul_cla32_fa11_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic11_and0 = s_csamul_cla32_fa12_31_xor1 & s_csamul_cla32_fa11_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic11_xor0 = s_csamul_cla32_fa12_31_xor1 ^ s_csamul_cla32_fa11_31_or0;
  assign s_csamul_cla32_u_cla32_xor11 = s_csamul_cla32_u_cla32_pg_logic11_xor0 ^ s_csamul_cla32_u_cla32_or21;
  assign s_csamul_cla32_u_cla32_and42 = s_csamul_cla32_u_cla32_or15 & s_csamul_cla32_u_cla32_pg_logic10_or0;
  assign s_csamul_cla32_u_cla32_and43 = s_csamul_cla32_u_cla32_pg_logic11_or0 & s_csamul_cla32_u_cla32_pg_logic9_or0;
  assign s_csamul_cla32_u_cla32_and44 = s_csamul_cla32_u_cla32_and42 & s_csamul_cla32_u_cla32_and43;
  assign s_csamul_cla32_u_cla32_and45 = s_csamul_cla32_u_cla32_and44 & s_csamul_cla32_u_cla32_pg_logic8_or0;
  assign s_csamul_cla32_u_cla32_and46 = s_csamul_cla32_u_cla32_pg_logic8_and0 & s_csamul_cla32_u_cla32_pg_logic10_or0;
  assign s_csamul_cla32_u_cla32_and47 = s_csamul_cla32_u_cla32_pg_logic11_or0 & s_csamul_cla32_u_cla32_pg_logic9_or0;
  assign s_csamul_cla32_u_cla32_and48 = s_csamul_cla32_u_cla32_and46 & s_csamul_cla32_u_cla32_and47;
  assign s_csamul_cla32_u_cla32_and49 = s_csamul_cla32_u_cla32_pg_logic9_and0 & s_csamul_cla32_u_cla32_pg_logic11_or0;
  assign s_csamul_cla32_u_cla32_and50 = s_csamul_cla32_u_cla32_and49 & s_csamul_cla32_u_cla32_pg_logic10_or0;
  assign s_csamul_cla32_u_cla32_and51 = s_csamul_cla32_u_cla32_pg_logic10_and0 & s_csamul_cla32_u_cla32_pg_logic11_or0;
  assign s_csamul_cla32_u_cla32_or22 = s_csamul_cla32_u_cla32_and45 | s_csamul_cla32_u_cla32_and50;
  assign s_csamul_cla32_u_cla32_or23 = s_csamul_cla32_u_cla32_and48 | s_csamul_cla32_u_cla32_and51;
  assign s_csamul_cla32_u_cla32_or24 = s_csamul_cla32_u_cla32_or22 | s_csamul_cla32_u_cla32_or23;
  assign s_csamul_cla32_u_cla32_or25 = s_csamul_cla32_u_cla32_pg_logic11_and0 | s_csamul_cla32_u_cla32_or24;
  assign s_csamul_cla32_u_cla32_pg_logic12_or0 = s_csamul_cla32_fa13_31_xor1 | s_csamul_cla32_fa12_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic12_and0 = s_csamul_cla32_fa13_31_xor1 & s_csamul_cla32_fa12_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic12_xor0 = s_csamul_cla32_fa13_31_xor1 ^ s_csamul_cla32_fa12_31_or0;
  assign s_csamul_cla32_u_cla32_xor12 = s_csamul_cla32_u_cla32_pg_logic12_xor0 ^ s_csamul_cla32_u_cla32_or25;
  assign s_csamul_cla32_u_cla32_and52 = s_csamul_cla32_u_cla32_or25 & s_csamul_cla32_u_cla32_pg_logic12_or0;
  assign s_csamul_cla32_u_cla32_or26 = s_csamul_cla32_u_cla32_pg_logic12_and0 | s_csamul_cla32_u_cla32_and52;
  assign s_csamul_cla32_u_cla32_pg_logic13_or0 = s_csamul_cla32_fa14_31_xor1 | s_csamul_cla32_fa13_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic13_and0 = s_csamul_cla32_fa14_31_xor1 & s_csamul_cla32_fa13_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic13_xor0 = s_csamul_cla32_fa14_31_xor1 ^ s_csamul_cla32_fa13_31_or0;
  assign s_csamul_cla32_u_cla32_xor13 = s_csamul_cla32_u_cla32_pg_logic13_xor0 ^ s_csamul_cla32_u_cla32_or26;
  assign s_csamul_cla32_u_cla32_and53 = s_csamul_cla32_u_cla32_or25 & s_csamul_cla32_u_cla32_pg_logic13_or0;
  assign s_csamul_cla32_u_cla32_and54 = s_csamul_cla32_u_cla32_and53 & s_csamul_cla32_u_cla32_pg_logic12_or0;
  assign s_csamul_cla32_u_cla32_and55 = s_csamul_cla32_u_cla32_pg_logic12_and0 & s_csamul_cla32_u_cla32_pg_logic13_or0;
  assign s_csamul_cla32_u_cla32_or27 = s_csamul_cla32_u_cla32_and54 | s_csamul_cla32_u_cla32_and55;
  assign s_csamul_cla32_u_cla32_or28 = s_csamul_cla32_u_cla32_pg_logic13_and0 | s_csamul_cla32_u_cla32_or27;
  assign s_csamul_cla32_u_cla32_pg_logic14_or0 = s_csamul_cla32_fa15_31_xor1 | s_csamul_cla32_fa14_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic14_and0 = s_csamul_cla32_fa15_31_xor1 & s_csamul_cla32_fa14_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic14_xor0 = s_csamul_cla32_fa15_31_xor1 ^ s_csamul_cla32_fa14_31_or0;
  assign s_csamul_cla32_u_cla32_xor14 = s_csamul_cla32_u_cla32_pg_logic14_xor0 ^ s_csamul_cla32_u_cla32_or28;
  assign s_csamul_cla32_u_cla32_and56 = s_csamul_cla32_u_cla32_or25 & s_csamul_cla32_u_cla32_pg_logic13_or0;
  assign s_csamul_cla32_u_cla32_and57 = s_csamul_cla32_u_cla32_pg_logic14_or0 & s_csamul_cla32_u_cla32_pg_logic12_or0;
  assign s_csamul_cla32_u_cla32_and58 = s_csamul_cla32_u_cla32_and56 & s_csamul_cla32_u_cla32_and57;
  assign s_csamul_cla32_u_cla32_and59 = s_csamul_cla32_u_cla32_pg_logic12_and0 & s_csamul_cla32_u_cla32_pg_logic14_or0;
  assign s_csamul_cla32_u_cla32_and60 = s_csamul_cla32_u_cla32_and59 & s_csamul_cla32_u_cla32_pg_logic13_or0;
  assign s_csamul_cla32_u_cla32_and61 = s_csamul_cla32_u_cla32_pg_logic13_and0 & s_csamul_cla32_u_cla32_pg_logic14_or0;
  assign s_csamul_cla32_u_cla32_or29 = s_csamul_cla32_u_cla32_and58 | s_csamul_cla32_u_cla32_and60;
  assign s_csamul_cla32_u_cla32_or30 = s_csamul_cla32_u_cla32_or29 | s_csamul_cla32_u_cla32_and61;
  assign s_csamul_cla32_u_cla32_or31 = s_csamul_cla32_u_cla32_pg_logic14_and0 | s_csamul_cla32_u_cla32_or30;
  assign s_csamul_cla32_u_cla32_pg_logic15_or0 = s_csamul_cla32_fa16_31_xor1 | s_csamul_cla32_fa15_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic15_and0 = s_csamul_cla32_fa16_31_xor1 & s_csamul_cla32_fa15_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic15_xor0 = s_csamul_cla32_fa16_31_xor1 ^ s_csamul_cla32_fa15_31_or0;
  assign s_csamul_cla32_u_cla32_xor15 = s_csamul_cla32_u_cla32_pg_logic15_xor0 ^ s_csamul_cla32_u_cla32_or31;
  assign s_csamul_cla32_u_cla32_and62 = s_csamul_cla32_u_cla32_or25 & s_csamul_cla32_u_cla32_pg_logic14_or0;
  assign s_csamul_cla32_u_cla32_and63 = s_csamul_cla32_u_cla32_pg_logic15_or0 & s_csamul_cla32_u_cla32_pg_logic13_or0;
  assign s_csamul_cla32_u_cla32_and64 = s_csamul_cla32_u_cla32_and62 & s_csamul_cla32_u_cla32_and63;
  assign s_csamul_cla32_u_cla32_and65 = s_csamul_cla32_u_cla32_and64 & s_csamul_cla32_u_cla32_pg_logic12_or0;
  assign s_csamul_cla32_u_cla32_and66 = s_csamul_cla32_u_cla32_pg_logic12_and0 & s_csamul_cla32_u_cla32_pg_logic14_or0;
  assign s_csamul_cla32_u_cla32_and67 = s_csamul_cla32_u_cla32_pg_logic15_or0 & s_csamul_cla32_u_cla32_pg_logic13_or0;
  assign s_csamul_cla32_u_cla32_and68 = s_csamul_cla32_u_cla32_and66 & s_csamul_cla32_u_cla32_and67;
  assign s_csamul_cla32_u_cla32_and69 = s_csamul_cla32_u_cla32_pg_logic13_and0 & s_csamul_cla32_u_cla32_pg_logic15_or0;
  assign s_csamul_cla32_u_cla32_and70 = s_csamul_cla32_u_cla32_and69 & s_csamul_cla32_u_cla32_pg_logic14_or0;
  assign s_csamul_cla32_u_cla32_and71 = s_csamul_cla32_u_cla32_pg_logic14_and0 & s_csamul_cla32_u_cla32_pg_logic15_or0;
  assign s_csamul_cla32_u_cla32_or32 = s_csamul_cla32_u_cla32_and65 | s_csamul_cla32_u_cla32_and70;
  assign s_csamul_cla32_u_cla32_or33 = s_csamul_cla32_u_cla32_and68 | s_csamul_cla32_u_cla32_and71;
  assign s_csamul_cla32_u_cla32_or34 = s_csamul_cla32_u_cla32_or32 | s_csamul_cla32_u_cla32_or33;
  assign s_csamul_cla32_u_cla32_or35 = s_csamul_cla32_u_cla32_pg_logic15_and0 | s_csamul_cla32_u_cla32_or34;
  assign s_csamul_cla32_u_cla32_pg_logic16_or0 = s_csamul_cla32_fa17_31_xor1 | s_csamul_cla32_fa16_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic16_and0 = s_csamul_cla32_fa17_31_xor1 & s_csamul_cla32_fa16_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic16_xor0 = s_csamul_cla32_fa17_31_xor1 ^ s_csamul_cla32_fa16_31_or0;
  assign s_csamul_cla32_u_cla32_xor16 = s_csamul_cla32_u_cla32_pg_logic16_xor0 ^ s_csamul_cla32_u_cla32_or35;
  assign s_csamul_cla32_u_cla32_and72 = s_csamul_cla32_u_cla32_or35 & s_csamul_cla32_u_cla32_pg_logic16_or0;
  assign s_csamul_cla32_u_cla32_or36 = s_csamul_cla32_u_cla32_pg_logic16_and0 | s_csamul_cla32_u_cla32_and72;
  assign s_csamul_cla32_u_cla32_pg_logic17_or0 = s_csamul_cla32_fa18_31_xor1 | s_csamul_cla32_fa17_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic17_and0 = s_csamul_cla32_fa18_31_xor1 & s_csamul_cla32_fa17_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic17_xor0 = s_csamul_cla32_fa18_31_xor1 ^ s_csamul_cla32_fa17_31_or0;
  assign s_csamul_cla32_u_cla32_xor17 = s_csamul_cla32_u_cla32_pg_logic17_xor0 ^ s_csamul_cla32_u_cla32_or36;
  assign s_csamul_cla32_u_cla32_and73 = s_csamul_cla32_u_cla32_or35 & s_csamul_cla32_u_cla32_pg_logic17_or0;
  assign s_csamul_cla32_u_cla32_and74 = s_csamul_cla32_u_cla32_and73 & s_csamul_cla32_u_cla32_pg_logic16_or0;
  assign s_csamul_cla32_u_cla32_and75 = s_csamul_cla32_u_cla32_pg_logic16_and0 & s_csamul_cla32_u_cla32_pg_logic17_or0;
  assign s_csamul_cla32_u_cla32_or37 = s_csamul_cla32_u_cla32_and74 | s_csamul_cla32_u_cla32_and75;
  assign s_csamul_cla32_u_cla32_or38 = s_csamul_cla32_u_cla32_pg_logic17_and0 | s_csamul_cla32_u_cla32_or37;
  assign s_csamul_cla32_u_cla32_pg_logic18_or0 = s_csamul_cla32_fa19_31_xor1 | s_csamul_cla32_fa18_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic18_and0 = s_csamul_cla32_fa19_31_xor1 & s_csamul_cla32_fa18_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic18_xor0 = s_csamul_cla32_fa19_31_xor1 ^ s_csamul_cla32_fa18_31_or0;
  assign s_csamul_cla32_u_cla32_xor18 = s_csamul_cla32_u_cla32_pg_logic18_xor0 ^ s_csamul_cla32_u_cla32_or38;
  assign s_csamul_cla32_u_cla32_and76 = s_csamul_cla32_u_cla32_or35 & s_csamul_cla32_u_cla32_pg_logic17_or0;
  assign s_csamul_cla32_u_cla32_and77 = s_csamul_cla32_u_cla32_pg_logic18_or0 & s_csamul_cla32_u_cla32_pg_logic16_or0;
  assign s_csamul_cla32_u_cla32_and78 = s_csamul_cla32_u_cla32_and76 & s_csamul_cla32_u_cla32_and77;
  assign s_csamul_cla32_u_cla32_and79 = s_csamul_cla32_u_cla32_pg_logic16_and0 & s_csamul_cla32_u_cla32_pg_logic18_or0;
  assign s_csamul_cla32_u_cla32_and80 = s_csamul_cla32_u_cla32_and79 & s_csamul_cla32_u_cla32_pg_logic17_or0;
  assign s_csamul_cla32_u_cla32_and81 = s_csamul_cla32_u_cla32_pg_logic17_and0 & s_csamul_cla32_u_cla32_pg_logic18_or0;
  assign s_csamul_cla32_u_cla32_or39 = s_csamul_cla32_u_cla32_and78 | s_csamul_cla32_u_cla32_and80;
  assign s_csamul_cla32_u_cla32_or40 = s_csamul_cla32_u_cla32_or39 | s_csamul_cla32_u_cla32_and81;
  assign s_csamul_cla32_u_cla32_or41 = s_csamul_cla32_u_cla32_pg_logic18_and0 | s_csamul_cla32_u_cla32_or40;
  assign s_csamul_cla32_u_cla32_pg_logic19_or0 = s_csamul_cla32_fa20_31_xor1 | s_csamul_cla32_fa19_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic19_and0 = s_csamul_cla32_fa20_31_xor1 & s_csamul_cla32_fa19_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic19_xor0 = s_csamul_cla32_fa20_31_xor1 ^ s_csamul_cla32_fa19_31_or0;
  assign s_csamul_cla32_u_cla32_xor19 = s_csamul_cla32_u_cla32_pg_logic19_xor0 ^ s_csamul_cla32_u_cla32_or41;
  assign s_csamul_cla32_u_cla32_and82 = s_csamul_cla32_u_cla32_or35 & s_csamul_cla32_u_cla32_pg_logic18_or0;
  assign s_csamul_cla32_u_cla32_and83 = s_csamul_cla32_u_cla32_pg_logic19_or0 & s_csamul_cla32_u_cla32_pg_logic17_or0;
  assign s_csamul_cla32_u_cla32_and84 = s_csamul_cla32_u_cla32_and82 & s_csamul_cla32_u_cla32_and83;
  assign s_csamul_cla32_u_cla32_and85 = s_csamul_cla32_u_cla32_and84 & s_csamul_cla32_u_cla32_pg_logic16_or0;
  assign s_csamul_cla32_u_cla32_and86 = s_csamul_cla32_u_cla32_pg_logic16_and0 & s_csamul_cla32_u_cla32_pg_logic18_or0;
  assign s_csamul_cla32_u_cla32_and87 = s_csamul_cla32_u_cla32_pg_logic19_or0 & s_csamul_cla32_u_cla32_pg_logic17_or0;
  assign s_csamul_cla32_u_cla32_and88 = s_csamul_cla32_u_cla32_and86 & s_csamul_cla32_u_cla32_and87;
  assign s_csamul_cla32_u_cla32_and89 = s_csamul_cla32_u_cla32_pg_logic17_and0 & s_csamul_cla32_u_cla32_pg_logic19_or0;
  assign s_csamul_cla32_u_cla32_and90 = s_csamul_cla32_u_cla32_and89 & s_csamul_cla32_u_cla32_pg_logic18_or0;
  assign s_csamul_cla32_u_cla32_and91 = s_csamul_cla32_u_cla32_pg_logic18_and0 & s_csamul_cla32_u_cla32_pg_logic19_or0;
  assign s_csamul_cla32_u_cla32_or42 = s_csamul_cla32_u_cla32_and85 | s_csamul_cla32_u_cla32_and90;
  assign s_csamul_cla32_u_cla32_or43 = s_csamul_cla32_u_cla32_and88 | s_csamul_cla32_u_cla32_and91;
  assign s_csamul_cla32_u_cla32_or44 = s_csamul_cla32_u_cla32_or42 | s_csamul_cla32_u_cla32_or43;
  assign s_csamul_cla32_u_cla32_or45 = s_csamul_cla32_u_cla32_pg_logic19_and0 | s_csamul_cla32_u_cla32_or44;
  assign s_csamul_cla32_u_cla32_pg_logic20_or0 = s_csamul_cla32_fa21_31_xor1 | s_csamul_cla32_fa20_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic20_and0 = s_csamul_cla32_fa21_31_xor1 & s_csamul_cla32_fa20_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic20_xor0 = s_csamul_cla32_fa21_31_xor1 ^ s_csamul_cla32_fa20_31_or0;
  assign s_csamul_cla32_u_cla32_xor20 = s_csamul_cla32_u_cla32_pg_logic20_xor0 ^ s_csamul_cla32_u_cla32_or45;
  assign s_csamul_cla32_u_cla32_and92 = s_csamul_cla32_u_cla32_or45 & s_csamul_cla32_u_cla32_pg_logic20_or0;
  assign s_csamul_cla32_u_cla32_or46 = s_csamul_cla32_u_cla32_pg_logic20_and0 | s_csamul_cla32_u_cla32_and92;
  assign s_csamul_cla32_u_cla32_pg_logic21_or0 = s_csamul_cla32_fa22_31_xor1 | s_csamul_cla32_fa21_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic21_and0 = s_csamul_cla32_fa22_31_xor1 & s_csamul_cla32_fa21_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic21_xor0 = s_csamul_cla32_fa22_31_xor1 ^ s_csamul_cla32_fa21_31_or0;
  assign s_csamul_cla32_u_cla32_xor21 = s_csamul_cla32_u_cla32_pg_logic21_xor0 ^ s_csamul_cla32_u_cla32_or46;
  assign s_csamul_cla32_u_cla32_and93 = s_csamul_cla32_u_cla32_or45 & s_csamul_cla32_u_cla32_pg_logic21_or0;
  assign s_csamul_cla32_u_cla32_and94 = s_csamul_cla32_u_cla32_and93 & s_csamul_cla32_u_cla32_pg_logic20_or0;
  assign s_csamul_cla32_u_cla32_and95 = s_csamul_cla32_u_cla32_pg_logic20_and0 & s_csamul_cla32_u_cla32_pg_logic21_or0;
  assign s_csamul_cla32_u_cla32_or47 = s_csamul_cla32_u_cla32_and94 | s_csamul_cla32_u_cla32_and95;
  assign s_csamul_cla32_u_cla32_or48 = s_csamul_cla32_u_cla32_pg_logic21_and0 | s_csamul_cla32_u_cla32_or47;
  assign s_csamul_cla32_u_cla32_pg_logic22_or0 = s_csamul_cla32_fa23_31_xor1 | s_csamul_cla32_fa22_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic22_and0 = s_csamul_cla32_fa23_31_xor1 & s_csamul_cla32_fa22_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic22_xor0 = s_csamul_cla32_fa23_31_xor1 ^ s_csamul_cla32_fa22_31_or0;
  assign s_csamul_cla32_u_cla32_xor22 = s_csamul_cla32_u_cla32_pg_logic22_xor0 ^ s_csamul_cla32_u_cla32_or48;
  assign s_csamul_cla32_u_cla32_and96 = s_csamul_cla32_u_cla32_or45 & s_csamul_cla32_u_cla32_pg_logic21_or0;
  assign s_csamul_cla32_u_cla32_and97 = s_csamul_cla32_u_cla32_pg_logic22_or0 & s_csamul_cla32_u_cla32_pg_logic20_or0;
  assign s_csamul_cla32_u_cla32_and98 = s_csamul_cla32_u_cla32_and96 & s_csamul_cla32_u_cla32_and97;
  assign s_csamul_cla32_u_cla32_and99 = s_csamul_cla32_u_cla32_pg_logic20_and0 & s_csamul_cla32_u_cla32_pg_logic22_or0;
  assign s_csamul_cla32_u_cla32_and100 = s_csamul_cla32_u_cla32_and99 & s_csamul_cla32_u_cla32_pg_logic21_or0;
  assign s_csamul_cla32_u_cla32_and101 = s_csamul_cla32_u_cla32_pg_logic21_and0 & s_csamul_cla32_u_cla32_pg_logic22_or0;
  assign s_csamul_cla32_u_cla32_or49 = s_csamul_cla32_u_cla32_and98 | s_csamul_cla32_u_cla32_and100;
  assign s_csamul_cla32_u_cla32_or50 = s_csamul_cla32_u_cla32_or49 | s_csamul_cla32_u_cla32_and101;
  assign s_csamul_cla32_u_cla32_or51 = s_csamul_cla32_u_cla32_pg_logic22_and0 | s_csamul_cla32_u_cla32_or50;
  assign s_csamul_cla32_u_cla32_pg_logic23_or0 = s_csamul_cla32_fa24_31_xor1 | s_csamul_cla32_fa23_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic23_and0 = s_csamul_cla32_fa24_31_xor1 & s_csamul_cla32_fa23_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic23_xor0 = s_csamul_cla32_fa24_31_xor1 ^ s_csamul_cla32_fa23_31_or0;
  assign s_csamul_cla32_u_cla32_xor23 = s_csamul_cla32_u_cla32_pg_logic23_xor0 ^ s_csamul_cla32_u_cla32_or51;
  assign s_csamul_cla32_u_cla32_and102 = s_csamul_cla32_u_cla32_or45 & s_csamul_cla32_u_cla32_pg_logic22_or0;
  assign s_csamul_cla32_u_cla32_and103 = s_csamul_cla32_u_cla32_pg_logic23_or0 & s_csamul_cla32_u_cla32_pg_logic21_or0;
  assign s_csamul_cla32_u_cla32_and104 = s_csamul_cla32_u_cla32_and102 & s_csamul_cla32_u_cla32_and103;
  assign s_csamul_cla32_u_cla32_and105 = s_csamul_cla32_u_cla32_and104 & s_csamul_cla32_u_cla32_pg_logic20_or0;
  assign s_csamul_cla32_u_cla32_and106 = s_csamul_cla32_u_cla32_pg_logic20_and0 & s_csamul_cla32_u_cla32_pg_logic22_or0;
  assign s_csamul_cla32_u_cla32_and107 = s_csamul_cla32_u_cla32_pg_logic23_or0 & s_csamul_cla32_u_cla32_pg_logic21_or0;
  assign s_csamul_cla32_u_cla32_and108 = s_csamul_cla32_u_cla32_and106 & s_csamul_cla32_u_cla32_and107;
  assign s_csamul_cla32_u_cla32_and109 = s_csamul_cla32_u_cla32_pg_logic21_and0 & s_csamul_cla32_u_cla32_pg_logic23_or0;
  assign s_csamul_cla32_u_cla32_and110 = s_csamul_cla32_u_cla32_and109 & s_csamul_cla32_u_cla32_pg_logic22_or0;
  assign s_csamul_cla32_u_cla32_and111 = s_csamul_cla32_u_cla32_pg_logic22_and0 & s_csamul_cla32_u_cla32_pg_logic23_or0;
  assign s_csamul_cla32_u_cla32_or52 = s_csamul_cla32_u_cla32_and105 | s_csamul_cla32_u_cla32_and110;
  assign s_csamul_cla32_u_cla32_or53 = s_csamul_cla32_u_cla32_and108 | s_csamul_cla32_u_cla32_and111;
  assign s_csamul_cla32_u_cla32_or54 = s_csamul_cla32_u_cla32_or52 | s_csamul_cla32_u_cla32_or53;
  assign s_csamul_cla32_u_cla32_or55 = s_csamul_cla32_u_cla32_pg_logic23_and0 | s_csamul_cla32_u_cla32_or54;
  assign s_csamul_cla32_u_cla32_pg_logic24_or0 = s_csamul_cla32_fa25_31_xor1 | s_csamul_cla32_fa24_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic24_and0 = s_csamul_cla32_fa25_31_xor1 & s_csamul_cla32_fa24_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic24_xor0 = s_csamul_cla32_fa25_31_xor1 ^ s_csamul_cla32_fa24_31_or0;
  assign s_csamul_cla32_u_cla32_xor24 = s_csamul_cla32_u_cla32_pg_logic24_xor0 ^ s_csamul_cla32_u_cla32_or55;
  assign s_csamul_cla32_u_cla32_and112 = s_csamul_cla32_u_cla32_or55 & s_csamul_cla32_u_cla32_pg_logic24_or0;
  assign s_csamul_cla32_u_cla32_or56 = s_csamul_cla32_u_cla32_pg_logic24_and0 | s_csamul_cla32_u_cla32_and112;
  assign s_csamul_cla32_u_cla32_pg_logic25_or0 = s_csamul_cla32_fa26_31_xor1 | s_csamul_cla32_fa25_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic25_and0 = s_csamul_cla32_fa26_31_xor1 & s_csamul_cla32_fa25_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic25_xor0 = s_csamul_cla32_fa26_31_xor1 ^ s_csamul_cla32_fa25_31_or0;
  assign s_csamul_cla32_u_cla32_xor25 = s_csamul_cla32_u_cla32_pg_logic25_xor0 ^ s_csamul_cla32_u_cla32_or56;
  assign s_csamul_cla32_u_cla32_and113 = s_csamul_cla32_u_cla32_or55 & s_csamul_cla32_u_cla32_pg_logic25_or0;
  assign s_csamul_cla32_u_cla32_and114 = s_csamul_cla32_u_cla32_and113 & s_csamul_cla32_u_cla32_pg_logic24_or0;
  assign s_csamul_cla32_u_cla32_and115 = s_csamul_cla32_u_cla32_pg_logic24_and0 & s_csamul_cla32_u_cla32_pg_logic25_or0;
  assign s_csamul_cla32_u_cla32_or57 = s_csamul_cla32_u_cla32_and114 | s_csamul_cla32_u_cla32_and115;
  assign s_csamul_cla32_u_cla32_or58 = s_csamul_cla32_u_cla32_pg_logic25_and0 | s_csamul_cla32_u_cla32_or57;
  assign s_csamul_cla32_u_cla32_pg_logic26_or0 = s_csamul_cla32_fa27_31_xor1 | s_csamul_cla32_fa26_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic26_and0 = s_csamul_cla32_fa27_31_xor1 & s_csamul_cla32_fa26_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic26_xor0 = s_csamul_cla32_fa27_31_xor1 ^ s_csamul_cla32_fa26_31_or0;
  assign s_csamul_cla32_u_cla32_xor26 = s_csamul_cla32_u_cla32_pg_logic26_xor0 ^ s_csamul_cla32_u_cla32_or58;
  assign s_csamul_cla32_u_cla32_and116 = s_csamul_cla32_u_cla32_or55 & s_csamul_cla32_u_cla32_pg_logic25_or0;
  assign s_csamul_cla32_u_cla32_and117 = s_csamul_cla32_u_cla32_pg_logic26_or0 & s_csamul_cla32_u_cla32_pg_logic24_or0;
  assign s_csamul_cla32_u_cla32_and118 = s_csamul_cla32_u_cla32_and116 & s_csamul_cla32_u_cla32_and117;
  assign s_csamul_cla32_u_cla32_and119 = s_csamul_cla32_u_cla32_pg_logic24_and0 & s_csamul_cla32_u_cla32_pg_logic26_or0;
  assign s_csamul_cla32_u_cla32_and120 = s_csamul_cla32_u_cla32_and119 & s_csamul_cla32_u_cla32_pg_logic25_or0;
  assign s_csamul_cla32_u_cla32_and121 = s_csamul_cla32_u_cla32_pg_logic25_and0 & s_csamul_cla32_u_cla32_pg_logic26_or0;
  assign s_csamul_cla32_u_cla32_or59 = s_csamul_cla32_u_cla32_and118 | s_csamul_cla32_u_cla32_and120;
  assign s_csamul_cla32_u_cla32_or60 = s_csamul_cla32_u_cla32_or59 | s_csamul_cla32_u_cla32_and121;
  assign s_csamul_cla32_u_cla32_or61 = s_csamul_cla32_u_cla32_pg_logic26_and0 | s_csamul_cla32_u_cla32_or60;
  assign s_csamul_cla32_u_cla32_pg_logic27_or0 = s_csamul_cla32_fa28_31_xor1 | s_csamul_cla32_fa27_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic27_and0 = s_csamul_cla32_fa28_31_xor1 & s_csamul_cla32_fa27_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic27_xor0 = s_csamul_cla32_fa28_31_xor1 ^ s_csamul_cla32_fa27_31_or0;
  assign s_csamul_cla32_u_cla32_xor27 = s_csamul_cla32_u_cla32_pg_logic27_xor0 ^ s_csamul_cla32_u_cla32_or61;
  assign s_csamul_cla32_u_cla32_and122 = s_csamul_cla32_u_cla32_or55 & s_csamul_cla32_u_cla32_pg_logic26_or0;
  assign s_csamul_cla32_u_cla32_and123 = s_csamul_cla32_u_cla32_pg_logic27_or0 & s_csamul_cla32_u_cla32_pg_logic25_or0;
  assign s_csamul_cla32_u_cla32_and124 = s_csamul_cla32_u_cla32_and122 & s_csamul_cla32_u_cla32_and123;
  assign s_csamul_cla32_u_cla32_and125 = s_csamul_cla32_u_cla32_and124 & s_csamul_cla32_u_cla32_pg_logic24_or0;
  assign s_csamul_cla32_u_cla32_and126 = s_csamul_cla32_u_cla32_pg_logic24_and0 & s_csamul_cla32_u_cla32_pg_logic26_or0;
  assign s_csamul_cla32_u_cla32_and127 = s_csamul_cla32_u_cla32_pg_logic27_or0 & s_csamul_cla32_u_cla32_pg_logic25_or0;
  assign s_csamul_cla32_u_cla32_and128 = s_csamul_cla32_u_cla32_and126 & s_csamul_cla32_u_cla32_and127;
  assign s_csamul_cla32_u_cla32_and129 = s_csamul_cla32_u_cla32_pg_logic25_and0 & s_csamul_cla32_u_cla32_pg_logic27_or0;
  assign s_csamul_cla32_u_cla32_and130 = s_csamul_cla32_u_cla32_and129 & s_csamul_cla32_u_cla32_pg_logic26_or0;
  assign s_csamul_cla32_u_cla32_and131 = s_csamul_cla32_u_cla32_pg_logic26_and0 & s_csamul_cla32_u_cla32_pg_logic27_or0;
  assign s_csamul_cla32_u_cla32_or62 = s_csamul_cla32_u_cla32_and125 | s_csamul_cla32_u_cla32_and130;
  assign s_csamul_cla32_u_cla32_or63 = s_csamul_cla32_u_cla32_and128 | s_csamul_cla32_u_cla32_and131;
  assign s_csamul_cla32_u_cla32_or64 = s_csamul_cla32_u_cla32_or62 | s_csamul_cla32_u_cla32_or63;
  assign s_csamul_cla32_u_cla32_or65 = s_csamul_cla32_u_cla32_pg_logic27_and0 | s_csamul_cla32_u_cla32_or64;
  assign s_csamul_cla32_u_cla32_pg_logic28_or0 = s_csamul_cla32_fa29_31_xor1 | s_csamul_cla32_fa28_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic28_and0 = s_csamul_cla32_fa29_31_xor1 & s_csamul_cla32_fa28_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic28_xor0 = s_csamul_cla32_fa29_31_xor1 ^ s_csamul_cla32_fa28_31_or0;
  assign s_csamul_cla32_u_cla32_xor28 = s_csamul_cla32_u_cla32_pg_logic28_xor0 ^ s_csamul_cla32_u_cla32_or65;
  assign s_csamul_cla32_u_cla32_and132 = s_csamul_cla32_u_cla32_or65 & s_csamul_cla32_u_cla32_pg_logic28_or0;
  assign s_csamul_cla32_u_cla32_or66 = s_csamul_cla32_u_cla32_pg_logic28_and0 | s_csamul_cla32_u_cla32_and132;
  assign s_csamul_cla32_u_cla32_pg_logic29_or0 = s_csamul_cla32_fa30_31_xor1 | s_csamul_cla32_fa29_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic29_and0 = s_csamul_cla32_fa30_31_xor1 & s_csamul_cla32_fa29_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic29_xor0 = s_csamul_cla32_fa30_31_xor1 ^ s_csamul_cla32_fa29_31_or0;
  assign s_csamul_cla32_u_cla32_xor29 = s_csamul_cla32_u_cla32_pg_logic29_xor0 ^ s_csamul_cla32_u_cla32_or66;
  assign s_csamul_cla32_u_cla32_and133 = s_csamul_cla32_u_cla32_or65 & s_csamul_cla32_u_cla32_pg_logic29_or0;
  assign s_csamul_cla32_u_cla32_and134 = s_csamul_cla32_u_cla32_and133 & s_csamul_cla32_u_cla32_pg_logic28_or0;
  assign s_csamul_cla32_u_cla32_and135 = s_csamul_cla32_u_cla32_pg_logic28_and0 & s_csamul_cla32_u_cla32_pg_logic29_or0;
  assign s_csamul_cla32_u_cla32_or67 = s_csamul_cla32_u_cla32_and134 | s_csamul_cla32_u_cla32_and135;
  assign s_csamul_cla32_u_cla32_or68 = s_csamul_cla32_u_cla32_pg_logic29_and0 | s_csamul_cla32_u_cla32_or67;
  assign s_csamul_cla32_u_cla32_pg_logic30_or0 = s_csamul_cla32_ha31_31_xor0 | s_csamul_cla32_fa30_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic30_and0 = s_csamul_cla32_ha31_31_xor0 & s_csamul_cla32_fa30_31_or0;
  assign s_csamul_cla32_u_cla32_pg_logic30_xor0 = s_csamul_cla32_ha31_31_xor0 ^ s_csamul_cla32_fa30_31_or0;
  assign s_csamul_cla32_u_cla32_xor30 = s_csamul_cla32_u_cla32_pg_logic30_xor0 ^ s_csamul_cla32_u_cla32_or68;
  assign s_csamul_cla32_u_cla32_and136 = s_csamul_cla32_u_cla32_or65 & s_csamul_cla32_u_cla32_pg_logic29_or0;
  assign s_csamul_cla32_u_cla32_and137 = s_csamul_cla32_u_cla32_pg_logic30_or0 & s_csamul_cla32_u_cla32_pg_logic28_or0;
  assign s_csamul_cla32_u_cla32_and138 = s_csamul_cla32_u_cla32_and136 & s_csamul_cla32_u_cla32_and137;
  assign s_csamul_cla32_u_cla32_and139 = s_csamul_cla32_u_cla32_pg_logic28_and0 & s_csamul_cla32_u_cla32_pg_logic30_or0;
  assign s_csamul_cla32_u_cla32_and140 = s_csamul_cla32_u_cla32_and139 & s_csamul_cla32_u_cla32_pg_logic29_or0;
  assign s_csamul_cla32_u_cla32_and141 = s_csamul_cla32_u_cla32_pg_logic29_and0 & s_csamul_cla32_u_cla32_pg_logic30_or0;
  assign s_csamul_cla32_u_cla32_or69 = s_csamul_cla32_u_cla32_and138 | s_csamul_cla32_u_cla32_and140;
  assign s_csamul_cla32_u_cla32_or70 = s_csamul_cla32_u_cla32_or69 | s_csamul_cla32_u_cla32_and141;
  assign s_csamul_cla32_u_cla32_or71 = s_csamul_cla32_u_cla32_pg_logic30_and0 | s_csamul_cla32_u_cla32_or70;
  assign s_csamul_cla32_u_cla32_pg_logic31_xor0 = ~s_csamul_cla32_ha31_31_and0;
  assign s_csamul_cla32_u_cla32_xor31 = s_csamul_cla32_u_cla32_pg_logic31_xor0 ^ s_csamul_cla32_u_cla32_or71;
  assign s_csamul_cla32_u_cla32_and142 = s_csamul_cla32_u_cla32_or65 & s_csamul_cla32_u_cla32_pg_logic30_or0;
  assign s_csamul_cla32_u_cla32_and143 = s_csamul_cla32_u_cla32_and142 & s_csamul_cla32_u_cla32_pg_logic29_or0;
  assign s_csamul_cla32_u_cla32_and144 = s_csamul_cla32_u_cla32_and143 & s_csamul_cla32_u_cla32_pg_logic28_or0;
  assign s_csamul_cla32_u_cla32_and145 = s_csamul_cla32_u_cla32_pg_logic28_and0 & s_csamul_cla32_u_cla32_pg_logic30_or0;
  assign s_csamul_cla32_u_cla32_and146 = s_csamul_cla32_u_cla32_and145 & s_csamul_cla32_u_cla32_pg_logic29_or0;
  assign s_csamul_cla32_u_cla32_and147 = s_csamul_cla32_u_cla32_pg_logic29_and0 & s_csamul_cla32_u_cla32_pg_logic30_or0;
  assign s_csamul_cla32_u_cla32_or72 = s_csamul_cla32_u_cla32_and144 | s_csamul_cla32_u_cla32_and147;
  assign s_csamul_cla32_u_cla32_or73 = s_csamul_cla32_u_cla32_and146 | s_csamul_cla32_u_cla32_pg_logic30_and0;
  assign s_csamul_cla32_u_cla32_or74 = s_csamul_cla32_u_cla32_or72 | s_csamul_cla32_u_cla32_or73;
  assign s_csamul_cla32_u_cla32_or75 = s_csamul_cla32_ha31_31_and0 | s_csamul_cla32_u_cla32_or74;

  assign s_csamul_cla32_out[0] = s_csamul_cla32_and0_0;
  assign s_csamul_cla32_out[1] = s_csamul_cla32_ha0_1_xor0;
  assign s_csamul_cla32_out[2] = s_csamul_cla32_fa0_2_xor1;
  assign s_csamul_cla32_out[3] = s_csamul_cla32_fa0_3_xor1;
  assign s_csamul_cla32_out[4] = s_csamul_cla32_fa0_4_xor1;
  assign s_csamul_cla32_out[5] = s_csamul_cla32_fa0_5_xor1;
  assign s_csamul_cla32_out[6] = s_csamul_cla32_fa0_6_xor1;
  assign s_csamul_cla32_out[7] = s_csamul_cla32_fa0_7_xor1;
  assign s_csamul_cla32_out[8] = s_csamul_cla32_fa0_8_xor1;
  assign s_csamul_cla32_out[9] = s_csamul_cla32_fa0_9_xor1;
  assign s_csamul_cla32_out[10] = s_csamul_cla32_fa0_10_xor1;
  assign s_csamul_cla32_out[11] = s_csamul_cla32_fa0_11_xor1;
  assign s_csamul_cla32_out[12] = s_csamul_cla32_fa0_12_xor1;
  assign s_csamul_cla32_out[13] = s_csamul_cla32_fa0_13_xor1;
  assign s_csamul_cla32_out[14] = s_csamul_cla32_fa0_14_xor1;
  assign s_csamul_cla32_out[15] = s_csamul_cla32_fa0_15_xor1;
  assign s_csamul_cla32_out[16] = s_csamul_cla32_fa0_16_xor1;
  assign s_csamul_cla32_out[17] = s_csamul_cla32_fa0_17_xor1;
  assign s_csamul_cla32_out[18] = s_csamul_cla32_fa0_18_xor1;
  assign s_csamul_cla32_out[19] = s_csamul_cla32_fa0_19_xor1;
  assign s_csamul_cla32_out[20] = s_csamul_cla32_fa0_20_xor1;
  assign s_csamul_cla32_out[21] = s_csamul_cla32_fa0_21_xor1;
  assign s_csamul_cla32_out[22] = s_csamul_cla32_fa0_22_xor1;
  assign s_csamul_cla32_out[23] = s_csamul_cla32_fa0_23_xor1;
  assign s_csamul_cla32_out[24] = s_csamul_cla32_fa0_24_xor1;
  assign s_csamul_cla32_out[25] = s_csamul_cla32_fa0_25_xor1;
  assign s_csamul_cla32_out[26] = s_csamul_cla32_fa0_26_xor1;
  assign s_csamul_cla32_out[27] = s_csamul_cla32_fa0_27_xor1;
  assign s_csamul_cla32_out[28] = s_csamul_cla32_fa0_28_xor1;
  assign s_csamul_cla32_out[29] = s_csamul_cla32_fa0_29_xor1;
  assign s_csamul_cla32_out[30] = s_csamul_cla32_fa0_30_xor1;
  assign s_csamul_cla32_out[31] = s_csamul_cla32_fa0_31_xor1;
  assign s_csamul_cla32_out[32] = s_csamul_cla32_u_cla32_pg_logic0_xor0;
  assign s_csamul_cla32_out[33] = s_csamul_cla32_u_cla32_xor1;
  assign s_csamul_cla32_out[34] = s_csamul_cla32_u_cla32_xor2;
  assign s_csamul_cla32_out[35] = s_csamul_cla32_u_cla32_xor3;
  assign s_csamul_cla32_out[36] = s_csamul_cla32_u_cla32_xor4;
  assign s_csamul_cla32_out[37] = s_csamul_cla32_u_cla32_xor5;
  assign s_csamul_cla32_out[38] = s_csamul_cla32_u_cla32_xor6;
  assign s_csamul_cla32_out[39] = s_csamul_cla32_u_cla32_xor7;
  assign s_csamul_cla32_out[40] = s_csamul_cla32_u_cla32_xor8;
  assign s_csamul_cla32_out[41] = s_csamul_cla32_u_cla32_xor9;
  assign s_csamul_cla32_out[42] = s_csamul_cla32_u_cla32_xor10;
  assign s_csamul_cla32_out[43] = s_csamul_cla32_u_cla32_xor11;
  assign s_csamul_cla32_out[44] = s_csamul_cla32_u_cla32_xor12;
  assign s_csamul_cla32_out[45] = s_csamul_cla32_u_cla32_xor13;
  assign s_csamul_cla32_out[46] = s_csamul_cla32_u_cla32_xor14;
  assign s_csamul_cla32_out[47] = s_csamul_cla32_u_cla32_xor15;
  assign s_csamul_cla32_out[48] = s_csamul_cla32_u_cla32_xor16;
  assign s_csamul_cla32_out[49] = s_csamul_cla32_u_cla32_xor17;
  assign s_csamul_cla32_out[50] = s_csamul_cla32_u_cla32_xor18;
  assign s_csamul_cla32_out[51] = s_csamul_cla32_u_cla32_xor19;
  assign s_csamul_cla32_out[52] = s_csamul_cla32_u_cla32_xor20;
  assign s_csamul_cla32_out[53] = s_csamul_cla32_u_cla32_xor21;
  assign s_csamul_cla32_out[54] = s_csamul_cla32_u_cla32_xor22;
  assign s_csamul_cla32_out[55] = s_csamul_cla32_u_cla32_xor23;
  assign s_csamul_cla32_out[56] = s_csamul_cla32_u_cla32_xor24;
  assign s_csamul_cla32_out[57] = s_csamul_cla32_u_cla32_xor25;
  assign s_csamul_cla32_out[58] = s_csamul_cla32_u_cla32_xor26;
  assign s_csamul_cla32_out[59] = s_csamul_cla32_u_cla32_xor27;
  assign s_csamul_cla32_out[60] = s_csamul_cla32_u_cla32_xor28;
  assign s_csamul_cla32_out[61] = s_csamul_cla32_u_cla32_xor29;
  assign s_csamul_cla32_out[62] = s_csamul_cla32_u_cla32_xor30;
  assign s_csamul_cla32_out[63] = s_csamul_cla32_u_cla32_xor31;
endmodule