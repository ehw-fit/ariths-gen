module u_cla24(input [23:0] a, input [23:0] b, output [24:0] u_cla24_out);
  wire u_cla24_pg_logic0_or0;
  wire u_cla24_pg_logic0_and0;
  wire u_cla24_pg_logic0_xor0;
  wire u_cla24_pg_logic1_or0;
  wire u_cla24_pg_logic1_and0;
  wire u_cla24_pg_logic1_xor0;
  wire u_cla24_xor1;
  wire u_cla24_and0;
  wire u_cla24_or0;
  wire u_cla24_pg_logic2_or0;
  wire u_cla24_pg_logic2_and0;
  wire u_cla24_pg_logic2_xor0;
  wire u_cla24_xor2;
  wire u_cla24_and1;
  wire u_cla24_and2;
  wire u_cla24_and3;
  wire u_cla24_and4;
  wire u_cla24_or1;
  wire u_cla24_or2;
  wire u_cla24_pg_logic3_or0;
  wire u_cla24_pg_logic3_and0;
  wire u_cla24_pg_logic3_xor0;
  wire u_cla24_xor3;
  wire u_cla24_and5;
  wire u_cla24_and6;
  wire u_cla24_and7;
  wire u_cla24_and8;
  wire u_cla24_and9;
  wire u_cla24_and10;
  wire u_cla24_and11;
  wire u_cla24_or3;
  wire u_cla24_or4;
  wire u_cla24_or5;
  wire u_cla24_pg_logic4_or0;
  wire u_cla24_pg_logic4_and0;
  wire u_cla24_pg_logic4_xor0;
  wire u_cla24_xor4;
  wire u_cla24_and12;
  wire u_cla24_or6;
  wire u_cla24_pg_logic5_or0;
  wire u_cla24_pg_logic5_and0;
  wire u_cla24_pg_logic5_xor0;
  wire u_cla24_xor5;
  wire u_cla24_and13;
  wire u_cla24_and14;
  wire u_cla24_and15;
  wire u_cla24_or7;
  wire u_cla24_or8;
  wire u_cla24_pg_logic6_or0;
  wire u_cla24_pg_logic6_and0;
  wire u_cla24_pg_logic6_xor0;
  wire u_cla24_xor6;
  wire u_cla24_and16;
  wire u_cla24_and17;
  wire u_cla24_and18;
  wire u_cla24_and19;
  wire u_cla24_and20;
  wire u_cla24_and21;
  wire u_cla24_or9;
  wire u_cla24_or10;
  wire u_cla24_or11;
  wire u_cla24_pg_logic7_or0;
  wire u_cla24_pg_logic7_and0;
  wire u_cla24_pg_logic7_xor0;
  wire u_cla24_xor7;
  wire u_cla24_and22;
  wire u_cla24_and23;
  wire u_cla24_and24;
  wire u_cla24_and25;
  wire u_cla24_and26;
  wire u_cla24_and27;
  wire u_cla24_and28;
  wire u_cla24_and29;
  wire u_cla24_and30;
  wire u_cla24_and31;
  wire u_cla24_or12;
  wire u_cla24_or13;
  wire u_cla24_or14;
  wire u_cla24_or15;
  wire u_cla24_pg_logic8_or0;
  wire u_cla24_pg_logic8_and0;
  wire u_cla24_pg_logic8_xor0;
  wire u_cla24_xor8;
  wire u_cla24_and32;
  wire u_cla24_or16;
  wire u_cla24_pg_logic9_or0;
  wire u_cla24_pg_logic9_and0;
  wire u_cla24_pg_logic9_xor0;
  wire u_cla24_xor9;
  wire u_cla24_and33;
  wire u_cla24_and34;
  wire u_cla24_and35;
  wire u_cla24_or17;
  wire u_cla24_or18;
  wire u_cla24_pg_logic10_or0;
  wire u_cla24_pg_logic10_and0;
  wire u_cla24_pg_logic10_xor0;
  wire u_cla24_xor10;
  wire u_cla24_and36;
  wire u_cla24_and37;
  wire u_cla24_and38;
  wire u_cla24_and39;
  wire u_cla24_and40;
  wire u_cla24_and41;
  wire u_cla24_or19;
  wire u_cla24_or20;
  wire u_cla24_or21;
  wire u_cla24_pg_logic11_or0;
  wire u_cla24_pg_logic11_and0;
  wire u_cla24_pg_logic11_xor0;
  wire u_cla24_xor11;
  wire u_cla24_and42;
  wire u_cla24_and43;
  wire u_cla24_and44;
  wire u_cla24_and45;
  wire u_cla24_and46;
  wire u_cla24_and47;
  wire u_cla24_and48;
  wire u_cla24_and49;
  wire u_cla24_and50;
  wire u_cla24_and51;
  wire u_cla24_or22;
  wire u_cla24_or23;
  wire u_cla24_or24;
  wire u_cla24_or25;
  wire u_cla24_pg_logic12_or0;
  wire u_cla24_pg_logic12_and0;
  wire u_cla24_pg_logic12_xor0;
  wire u_cla24_xor12;
  wire u_cla24_and52;
  wire u_cla24_or26;
  wire u_cla24_pg_logic13_or0;
  wire u_cla24_pg_logic13_and0;
  wire u_cla24_pg_logic13_xor0;
  wire u_cla24_xor13;
  wire u_cla24_and53;
  wire u_cla24_and54;
  wire u_cla24_and55;
  wire u_cla24_or27;
  wire u_cla24_or28;
  wire u_cla24_pg_logic14_or0;
  wire u_cla24_pg_logic14_and0;
  wire u_cla24_pg_logic14_xor0;
  wire u_cla24_xor14;
  wire u_cla24_and56;
  wire u_cla24_and57;
  wire u_cla24_and58;
  wire u_cla24_and59;
  wire u_cla24_and60;
  wire u_cla24_and61;
  wire u_cla24_or29;
  wire u_cla24_or30;
  wire u_cla24_or31;
  wire u_cla24_pg_logic15_or0;
  wire u_cla24_pg_logic15_and0;
  wire u_cla24_pg_logic15_xor0;
  wire u_cla24_xor15;
  wire u_cla24_and62;
  wire u_cla24_and63;
  wire u_cla24_and64;
  wire u_cla24_and65;
  wire u_cla24_and66;
  wire u_cla24_and67;
  wire u_cla24_and68;
  wire u_cla24_and69;
  wire u_cla24_and70;
  wire u_cla24_and71;
  wire u_cla24_or32;
  wire u_cla24_or33;
  wire u_cla24_or34;
  wire u_cla24_or35;
  wire u_cla24_pg_logic16_or0;
  wire u_cla24_pg_logic16_and0;
  wire u_cla24_pg_logic16_xor0;
  wire u_cla24_xor16;
  wire u_cla24_and72;
  wire u_cla24_or36;
  wire u_cla24_pg_logic17_or0;
  wire u_cla24_pg_logic17_and0;
  wire u_cla24_pg_logic17_xor0;
  wire u_cla24_xor17;
  wire u_cla24_and73;
  wire u_cla24_and74;
  wire u_cla24_and75;
  wire u_cla24_or37;
  wire u_cla24_or38;
  wire u_cla24_pg_logic18_or0;
  wire u_cla24_pg_logic18_and0;
  wire u_cla24_pg_logic18_xor0;
  wire u_cla24_xor18;
  wire u_cla24_and76;
  wire u_cla24_and77;
  wire u_cla24_and78;
  wire u_cla24_and79;
  wire u_cla24_and80;
  wire u_cla24_and81;
  wire u_cla24_or39;
  wire u_cla24_or40;
  wire u_cla24_or41;
  wire u_cla24_pg_logic19_or0;
  wire u_cla24_pg_logic19_and0;
  wire u_cla24_pg_logic19_xor0;
  wire u_cla24_xor19;
  wire u_cla24_and82;
  wire u_cla24_and83;
  wire u_cla24_and84;
  wire u_cla24_and85;
  wire u_cla24_and86;
  wire u_cla24_and87;
  wire u_cla24_and88;
  wire u_cla24_and89;
  wire u_cla24_and90;
  wire u_cla24_and91;
  wire u_cla24_or42;
  wire u_cla24_or43;
  wire u_cla24_or44;
  wire u_cla24_or45;
  wire u_cla24_pg_logic20_or0;
  wire u_cla24_pg_logic20_and0;
  wire u_cla24_pg_logic20_xor0;
  wire u_cla24_xor20;
  wire u_cla24_and92;
  wire u_cla24_or46;
  wire u_cla24_pg_logic21_or0;
  wire u_cla24_pg_logic21_and0;
  wire u_cla24_pg_logic21_xor0;
  wire u_cla24_xor21;
  wire u_cla24_and93;
  wire u_cla24_and94;
  wire u_cla24_and95;
  wire u_cla24_or47;
  wire u_cla24_or48;
  wire u_cla24_pg_logic22_or0;
  wire u_cla24_pg_logic22_and0;
  wire u_cla24_pg_logic22_xor0;
  wire u_cla24_xor22;
  wire u_cla24_and96;
  wire u_cla24_and97;
  wire u_cla24_and98;
  wire u_cla24_and99;
  wire u_cla24_and100;
  wire u_cla24_and101;
  wire u_cla24_or49;
  wire u_cla24_or50;
  wire u_cla24_or51;
  wire u_cla24_pg_logic23_or0;
  wire u_cla24_pg_logic23_and0;
  wire u_cla24_pg_logic23_xor0;
  wire u_cla24_xor23;
  wire u_cla24_and102;
  wire u_cla24_and103;
  wire u_cla24_and104;
  wire u_cla24_and105;
  wire u_cla24_and106;
  wire u_cla24_and107;
  wire u_cla24_and108;
  wire u_cla24_and109;
  wire u_cla24_and110;
  wire u_cla24_and111;
  wire u_cla24_or52;
  wire u_cla24_or53;
  wire u_cla24_or54;
  wire u_cla24_or55;

  assign u_cla24_pg_logic0_or0 = a[0] | b[0];
  assign u_cla24_pg_logic0_and0 = a[0] & b[0];
  assign u_cla24_pg_logic0_xor0 = a[0] ^ b[0];
  assign u_cla24_pg_logic1_or0 = a[1] | b[1];
  assign u_cla24_pg_logic1_and0 = a[1] & b[1];
  assign u_cla24_pg_logic1_xor0 = a[1] ^ b[1];
  assign u_cla24_xor1 = u_cla24_pg_logic1_xor0 ^ u_cla24_pg_logic0_and0;
  assign u_cla24_and0 = u_cla24_pg_logic0_and0 & u_cla24_pg_logic1_or0;
  assign u_cla24_or0 = u_cla24_pg_logic1_and0 | u_cla24_and0;
  assign u_cla24_pg_logic2_or0 = a[2] | b[2];
  assign u_cla24_pg_logic2_and0 = a[2] & b[2];
  assign u_cla24_pg_logic2_xor0 = a[2] ^ b[2];
  assign u_cla24_xor2 = u_cla24_pg_logic2_xor0 ^ u_cla24_or0;
  assign u_cla24_and1 = u_cla24_pg_logic2_or0 & u_cla24_pg_logic0_or0;
  assign u_cla24_and2 = u_cla24_pg_logic0_and0 & u_cla24_pg_logic2_or0;
  assign u_cla24_and3 = u_cla24_and2 & u_cla24_pg_logic1_or0;
  assign u_cla24_and4 = u_cla24_pg_logic1_and0 & u_cla24_pg_logic2_or0;
  assign u_cla24_or1 = u_cla24_and3 | u_cla24_and4;
  assign u_cla24_or2 = u_cla24_pg_logic2_and0 | u_cla24_or1;
  assign u_cla24_pg_logic3_or0 = a[3] | b[3];
  assign u_cla24_pg_logic3_and0 = a[3] & b[3];
  assign u_cla24_pg_logic3_xor0 = a[3] ^ b[3];
  assign u_cla24_xor3 = u_cla24_pg_logic3_xor0 ^ u_cla24_or2;
  assign u_cla24_and5 = u_cla24_pg_logic3_or0 & u_cla24_pg_logic1_or0;
  assign u_cla24_and6 = u_cla24_pg_logic0_and0 & u_cla24_pg_logic2_or0;
  assign u_cla24_and7 = u_cla24_pg_logic3_or0 & u_cla24_pg_logic1_or0;
  assign u_cla24_and8 = u_cla24_and6 & u_cla24_and7;
  assign u_cla24_and9 = u_cla24_pg_logic1_and0 & u_cla24_pg_logic3_or0;
  assign u_cla24_and10 = u_cla24_and9 & u_cla24_pg_logic2_or0;
  assign u_cla24_and11 = u_cla24_pg_logic2_and0 & u_cla24_pg_logic3_or0;
  assign u_cla24_or3 = u_cla24_and8 | u_cla24_and11;
  assign u_cla24_or4 = u_cla24_and10 | u_cla24_or3;
  assign u_cla24_or5 = u_cla24_pg_logic3_and0 | u_cla24_or4;
  assign u_cla24_pg_logic4_or0 = a[4] | b[4];
  assign u_cla24_pg_logic4_and0 = a[4] & b[4];
  assign u_cla24_pg_logic4_xor0 = a[4] ^ b[4];
  assign u_cla24_xor4 = u_cla24_pg_logic4_xor0 ^ u_cla24_or5;
  assign u_cla24_and12 = u_cla24_or5 & u_cla24_pg_logic4_or0;
  assign u_cla24_or6 = u_cla24_pg_logic4_and0 | u_cla24_and12;
  assign u_cla24_pg_logic5_or0 = a[5] | b[5];
  assign u_cla24_pg_logic5_and0 = a[5] & b[5];
  assign u_cla24_pg_logic5_xor0 = a[5] ^ b[5];
  assign u_cla24_xor5 = u_cla24_pg_logic5_xor0 ^ u_cla24_or6;
  assign u_cla24_and13 = u_cla24_or5 & u_cla24_pg_logic5_or0;
  assign u_cla24_and14 = u_cla24_and13 & u_cla24_pg_logic4_or0;
  assign u_cla24_and15 = u_cla24_pg_logic4_and0 & u_cla24_pg_logic5_or0;
  assign u_cla24_or7 = u_cla24_and14 | u_cla24_and15;
  assign u_cla24_or8 = u_cla24_pg_logic5_and0 | u_cla24_or7;
  assign u_cla24_pg_logic6_or0 = a[6] | b[6];
  assign u_cla24_pg_logic6_and0 = a[6] & b[6];
  assign u_cla24_pg_logic6_xor0 = a[6] ^ b[6];
  assign u_cla24_xor6 = u_cla24_pg_logic6_xor0 ^ u_cla24_or8;
  assign u_cla24_and16 = u_cla24_or5 & u_cla24_pg_logic5_or0;
  assign u_cla24_and17 = u_cla24_pg_logic6_or0 & u_cla24_pg_logic4_or0;
  assign u_cla24_and18 = u_cla24_and16 & u_cla24_and17;
  assign u_cla24_and19 = u_cla24_pg_logic4_and0 & u_cla24_pg_logic6_or0;
  assign u_cla24_and20 = u_cla24_and19 & u_cla24_pg_logic5_or0;
  assign u_cla24_and21 = u_cla24_pg_logic5_and0 & u_cla24_pg_logic6_or0;
  assign u_cla24_or9 = u_cla24_and18 | u_cla24_and20;
  assign u_cla24_or10 = u_cla24_or9 | u_cla24_and21;
  assign u_cla24_or11 = u_cla24_pg_logic6_and0 | u_cla24_or10;
  assign u_cla24_pg_logic7_or0 = a[7] | b[7];
  assign u_cla24_pg_logic7_and0 = a[7] & b[7];
  assign u_cla24_pg_logic7_xor0 = a[7] ^ b[7];
  assign u_cla24_xor7 = u_cla24_pg_logic7_xor0 ^ u_cla24_or11;
  assign u_cla24_and22 = u_cla24_or5 & u_cla24_pg_logic6_or0;
  assign u_cla24_and23 = u_cla24_pg_logic7_or0 & u_cla24_pg_logic5_or0;
  assign u_cla24_and24 = u_cla24_and22 & u_cla24_and23;
  assign u_cla24_and25 = u_cla24_and24 & u_cla24_pg_logic4_or0;
  assign u_cla24_and26 = u_cla24_pg_logic4_and0 & u_cla24_pg_logic6_or0;
  assign u_cla24_and27 = u_cla24_pg_logic7_or0 & u_cla24_pg_logic5_or0;
  assign u_cla24_and28 = u_cla24_and26 & u_cla24_and27;
  assign u_cla24_and29 = u_cla24_pg_logic5_and0 & u_cla24_pg_logic7_or0;
  assign u_cla24_and30 = u_cla24_and29 & u_cla24_pg_logic6_or0;
  assign u_cla24_and31 = u_cla24_pg_logic6_and0 & u_cla24_pg_logic7_or0;
  assign u_cla24_or12 = u_cla24_and25 | u_cla24_and30;
  assign u_cla24_or13 = u_cla24_and28 | u_cla24_and31;
  assign u_cla24_or14 = u_cla24_or12 | u_cla24_or13;
  assign u_cla24_or15 = u_cla24_pg_logic7_and0 | u_cla24_or14;
  assign u_cla24_pg_logic8_or0 = a[8] | b[8];
  assign u_cla24_pg_logic8_and0 = a[8] & b[8];
  assign u_cla24_pg_logic8_xor0 = a[8] ^ b[8];
  assign u_cla24_xor8 = u_cla24_pg_logic8_xor0 ^ u_cla24_or15;
  assign u_cla24_and32 = u_cla24_or15 & u_cla24_pg_logic8_or0;
  assign u_cla24_or16 = u_cla24_pg_logic8_and0 | u_cla24_and32;
  assign u_cla24_pg_logic9_or0 = a[9] | b[9];
  assign u_cla24_pg_logic9_and0 = a[9] & b[9];
  assign u_cla24_pg_logic9_xor0 = a[9] ^ b[9];
  assign u_cla24_xor9 = u_cla24_pg_logic9_xor0 ^ u_cla24_or16;
  assign u_cla24_and33 = u_cla24_or15 & u_cla24_pg_logic9_or0;
  assign u_cla24_and34 = u_cla24_and33 & u_cla24_pg_logic8_or0;
  assign u_cla24_and35 = u_cla24_pg_logic8_and0 & u_cla24_pg_logic9_or0;
  assign u_cla24_or17 = u_cla24_and34 | u_cla24_and35;
  assign u_cla24_or18 = u_cla24_pg_logic9_and0 | u_cla24_or17;
  assign u_cla24_pg_logic10_or0 = a[10] | b[10];
  assign u_cla24_pg_logic10_and0 = a[10] & b[10];
  assign u_cla24_pg_logic10_xor0 = a[10] ^ b[10];
  assign u_cla24_xor10 = u_cla24_pg_logic10_xor0 ^ u_cla24_or18;
  assign u_cla24_and36 = u_cla24_or15 & u_cla24_pg_logic9_or0;
  assign u_cla24_and37 = u_cla24_pg_logic10_or0 & u_cla24_pg_logic8_or0;
  assign u_cla24_and38 = u_cla24_and36 & u_cla24_and37;
  assign u_cla24_and39 = u_cla24_pg_logic8_and0 & u_cla24_pg_logic10_or0;
  assign u_cla24_and40 = u_cla24_and39 & u_cla24_pg_logic9_or0;
  assign u_cla24_and41 = u_cla24_pg_logic9_and0 & u_cla24_pg_logic10_or0;
  assign u_cla24_or19 = u_cla24_and38 | u_cla24_and40;
  assign u_cla24_or20 = u_cla24_or19 | u_cla24_and41;
  assign u_cla24_or21 = u_cla24_pg_logic10_and0 | u_cla24_or20;
  assign u_cla24_pg_logic11_or0 = a[11] | b[11];
  assign u_cla24_pg_logic11_and0 = a[11] & b[11];
  assign u_cla24_pg_logic11_xor0 = a[11] ^ b[11];
  assign u_cla24_xor11 = u_cla24_pg_logic11_xor0 ^ u_cla24_or21;
  assign u_cla24_and42 = u_cla24_or15 & u_cla24_pg_logic10_or0;
  assign u_cla24_and43 = u_cla24_pg_logic11_or0 & u_cla24_pg_logic9_or0;
  assign u_cla24_and44 = u_cla24_and42 & u_cla24_and43;
  assign u_cla24_and45 = u_cla24_and44 & u_cla24_pg_logic8_or0;
  assign u_cla24_and46 = u_cla24_pg_logic8_and0 & u_cla24_pg_logic10_or0;
  assign u_cla24_and47 = u_cla24_pg_logic11_or0 & u_cla24_pg_logic9_or0;
  assign u_cla24_and48 = u_cla24_and46 & u_cla24_and47;
  assign u_cla24_and49 = u_cla24_pg_logic9_and0 & u_cla24_pg_logic11_or0;
  assign u_cla24_and50 = u_cla24_and49 & u_cla24_pg_logic10_or0;
  assign u_cla24_and51 = u_cla24_pg_logic10_and0 & u_cla24_pg_logic11_or0;
  assign u_cla24_or22 = u_cla24_and45 | u_cla24_and50;
  assign u_cla24_or23 = u_cla24_and48 | u_cla24_and51;
  assign u_cla24_or24 = u_cla24_or22 | u_cla24_or23;
  assign u_cla24_or25 = u_cla24_pg_logic11_and0 | u_cla24_or24;
  assign u_cla24_pg_logic12_or0 = a[12] | b[12];
  assign u_cla24_pg_logic12_and0 = a[12] & b[12];
  assign u_cla24_pg_logic12_xor0 = a[12] ^ b[12];
  assign u_cla24_xor12 = u_cla24_pg_logic12_xor0 ^ u_cla24_or25;
  assign u_cla24_and52 = u_cla24_or25 & u_cla24_pg_logic12_or0;
  assign u_cla24_or26 = u_cla24_pg_logic12_and0 | u_cla24_and52;
  assign u_cla24_pg_logic13_or0 = a[13] | b[13];
  assign u_cla24_pg_logic13_and0 = a[13] & b[13];
  assign u_cla24_pg_logic13_xor0 = a[13] ^ b[13];
  assign u_cla24_xor13 = u_cla24_pg_logic13_xor0 ^ u_cla24_or26;
  assign u_cla24_and53 = u_cla24_or25 & u_cla24_pg_logic13_or0;
  assign u_cla24_and54 = u_cla24_and53 & u_cla24_pg_logic12_or0;
  assign u_cla24_and55 = u_cla24_pg_logic12_and0 & u_cla24_pg_logic13_or0;
  assign u_cla24_or27 = u_cla24_and54 | u_cla24_and55;
  assign u_cla24_or28 = u_cla24_pg_logic13_and0 | u_cla24_or27;
  assign u_cla24_pg_logic14_or0 = a[14] | b[14];
  assign u_cla24_pg_logic14_and0 = a[14] & b[14];
  assign u_cla24_pg_logic14_xor0 = a[14] ^ b[14];
  assign u_cla24_xor14 = u_cla24_pg_logic14_xor0 ^ u_cla24_or28;
  assign u_cla24_and56 = u_cla24_or25 & u_cla24_pg_logic13_or0;
  assign u_cla24_and57 = u_cla24_pg_logic14_or0 & u_cla24_pg_logic12_or0;
  assign u_cla24_and58 = u_cla24_and56 & u_cla24_and57;
  assign u_cla24_and59 = u_cla24_pg_logic12_and0 & u_cla24_pg_logic14_or0;
  assign u_cla24_and60 = u_cla24_and59 & u_cla24_pg_logic13_or0;
  assign u_cla24_and61 = u_cla24_pg_logic13_and0 & u_cla24_pg_logic14_or0;
  assign u_cla24_or29 = u_cla24_and58 | u_cla24_and60;
  assign u_cla24_or30 = u_cla24_or29 | u_cla24_and61;
  assign u_cla24_or31 = u_cla24_pg_logic14_and0 | u_cla24_or30;
  assign u_cla24_pg_logic15_or0 = a[15] | b[15];
  assign u_cla24_pg_logic15_and0 = a[15] & b[15];
  assign u_cla24_pg_logic15_xor0 = a[15] ^ b[15];
  assign u_cla24_xor15 = u_cla24_pg_logic15_xor0 ^ u_cla24_or31;
  assign u_cla24_and62 = u_cla24_or25 & u_cla24_pg_logic14_or0;
  assign u_cla24_and63 = u_cla24_pg_logic15_or0 & u_cla24_pg_logic13_or0;
  assign u_cla24_and64 = u_cla24_and62 & u_cla24_and63;
  assign u_cla24_and65 = u_cla24_and64 & u_cla24_pg_logic12_or0;
  assign u_cla24_and66 = u_cla24_pg_logic12_and0 & u_cla24_pg_logic14_or0;
  assign u_cla24_and67 = u_cla24_pg_logic15_or0 & u_cla24_pg_logic13_or0;
  assign u_cla24_and68 = u_cla24_and66 & u_cla24_and67;
  assign u_cla24_and69 = u_cla24_pg_logic13_and0 & u_cla24_pg_logic15_or0;
  assign u_cla24_and70 = u_cla24_and69 & u_cla24_pg_logic14_or0;
  assign u_cla24_and71 = u_cla24_pg_logic14_and0 & u_cla24_pg_logic15_or0;
  assign u_cla24_or32 = u_cla24_and65 | u_cla24_and70;
  assign u_cla24_or33 = u_cla24_and68 | u_cla24_and71;
  assign u_cla24_or34 = u_cla24_or32 | u_cla24_or33;
  assign u_cla24_or35 = u_cla24_pg_logic15_and0 | u_cla24_or34;
  assign u_cla24_pg_logic16_or0 = a[16] | b[16];
  assign u_cla24_pg_logic16_and0 = a[16] & b[16];
  assign u_cla24_pg_logic16_xor0 = a[16] ^ b[16];
  assign u_cla24_xor16 = u_cla24_pg_logic16_xor0 ^ u_cla24_or35;
  assign u_cla24_and72 = u_cla24_or35 & u_cla24_pg_logic16_or0;
  assign u_cla24_or36 = u_cla24_pg_logic16_and0 | u_cla24_and72;
  assign u_cla24_pg_logic17_or0 = a[17] | b[17];
  assign u_cla24_pg_logic17_and0 = a[17] & b[17];
  assign u_cla24_pg_logic17_xor0 = a[17] ^ b[17];
  assign u_cla24_xor17 = u_cla24_pg_logic17_xor0 ^ u_cla24_or36;
  assign u_cla24_and73 = u_cla24_or35 & u_cla24_pg_logic17_or0;
  assign u_cla24_and74 = u_cla24_and73 & u_cla24_pg_logic16_or0;
  assign u_cla24_and75 = u_cla24_pg_logic16_and0 & u_cla24_pg_logic17_or0;
  assign u_cla24_or37 = u_cla24_and74 | u_cla24_and75;
  assign u_cla24_or38 = u_cla24_pg_logic17_and0 | u_cla24_or37;
  assign u_cla24_pg_logic18_or0 = a[18] | b[18];
  assign u_cla24_pg_logic18_and0 = a[18] & b[18];
  assign u_cla24_pg_logic18_xor0 = a[18] ^ b[18];
  assign u_cla24_xor18 = u_cla24_pg_logic18_xor0 ^ u_cla24_or38;
  assign u_cla24_and76 = u_cla24_or35 & u_cla24_pg_logic17_or0;
  assign u_cla24_and77 = u_cla24_pg_logic18_or0 & u_cla24_pg_logic16_or0;
  assign u_cla24_and78 = u_cla24_and76 & u_cla24_and77;
  assign u_cla24_and79 = u_cla24_pg_logic16_and0 & u_cla24_pg_logic18_or0;
  assign u_cla24_and80 = u_cla24_and79 & u_cla24_pg_logic17_or0;
  assign u_cla24_and81 = u_cla24_pg_logic17_and0 & u_cla24_pg_logic18_or0;
  assign u_cla24_or39 = u_cla24_and78 | u_cla24_and80;
  assign u_cla24_or40 = u_cla24_or39 | u_cla24_and81;
  assign u_cla24_or41 = u_cla24_pg_logic18_and0 | u_cla24_or40;
  assign u_cla24_pg_logic19_or0 = a[19] | b[19];
  assign u_cla24_pg_logic19_and0 = a[19] & b[19];
  assign u_cla24_pg_logic19_xor0 = a[19] ^ b[19];
  assign u_cla24_xor19 = u_cla24_pg_logic19_xor0 ^ u_cla24_or41;
  assign u_cla24_and82 = u_cla24_or35 & u_cla24_pg_logic18_or0;
  assign u_cla24_and83 = u_cla24_pg_logic19_or0 & u_cla24_pg_logic17_or0;
  assign u_cla24_and84 = u_cla24_and82 & u_cla24_and83;
  assign u_cla24_and85 = u_cla24_and84 & u_cla24_pg_logic16_or0;
  assign u_cla24_and86 = u_cla24_pg_logic16_and0 & u_cla24_pg_logic18_or0;
  assign u_cla24_and87 = u_cla24_pg_logic19_or0 & u_cla24_pg_logic17_or0;
  assign u_cla24_and88 = u_cla24_and86 & u_cla24_and87;
  assign u_cla24_and89 = u_cla24_pg_logic17_and0 & u_cla24_pg_logic19_or0;
  assign u_cla24_and90 = u_cla24_and89 & u_cla24_pg_logic18_or0;
  assign u_cla24_and91 = u_cla24_pg_logic18_and0 & u_cla24_pg_logic19_or0;
  assign u_cla24_or42 = u_cla24_and85 | u_cla24_and90;
  assign u_cla24_or43 = u_cla24_and88 | u_cla24_and91;
  assign u_cla24_or44 = u_cla24_or42 | u_cla24_or43;
  assign u_cla24_or45 = u_cla24_pg_logic19_and0 | u_cla24_or44;
  assign u_cla24_pg_logic20_or0 = a[20] | b[20];
  assign u_cla24_pg_logic20_and0 = a[20] & b[20];
  assign u_cla24_pg_logic20_xor0 = a[20] ^ b[20];
  assign u_cla24_xor20 = u_cla24_pg_logic20_xor0 ^ u_cla24_or45;
  assign u_cla24_and92 = u_cla24_or45 & u_cla24_pg_logic20_or0;
  assign u_cla24_or46 = u_cla24_pg_logic20_and0 | u_cla24_and92;
  assign u_cla24_pg_logic21_or0 = a[21] | b[21];
  assign u_cla24_pg_logic21_and0 = a[21] & b[21];
  assign u_cla24_pg_logic21_xor0 = a[21] ^ b[21];
  assign u_cla24_xor21 = u_cla24_pg_logic21_xor0 ^ u_cla24_or46;
  assign u_cla24_and93 = u_cla24_or45 & u_cla24_pg_logic21_or0;
  assign u_cla24_and94 = u_cla24_and93 & u_cla24_pg_logic20_or0;
  assign u_cla24_and95 = u_cla24_pg_logic20_and0 & u_cla24_pg_logic21_or0;
  assign u_cla24_or47 = u_cla24_and94 | u_cla24_and95;
  assign u_cla24_or48 = u_cla24_pg_logic21_and0 | u_cla24_or47;
  assign u_cla24_pg_logic22_or0 = a[22] | b[22];
  assign u_cla24_pg_logic22_and0 = a[22] & b[22];
  assign u_cla24_pg_logic22_xor0 = a[22] ^ b[22];
  assign u_cla24_xor22 = u_cla24_pg_logic22_xor0 ^ u_cla24_or48;
  assign u_cla24_and96 = u_cla24_or45 & u_cla24_pg_logic21_or0;
  assign u_cla24_and97 = u_cla24_pg_logic22_or0 & u_cla24_pg_logic20_or0;
  assign u_cla24_and98 = u_cla24_and96 & u_cla24_and97;
  assign u_cla24_and99 = u_cla24_pg_logic20_and0 & u_cla24_pg_logic22_or0;
  assign u_cla24_and100 = u_cla24_and99 & u_cla24_pg_logic21_or0;
  assign u_cla24_and101 = u_cla24_pg_logic21_and0 & u_cla24_pg_logic22_or0;
  assign u_cla24_or49 = u_cla24_and98 | u_cla24_and100;
  assign u_cla24_or50 = u_cla24_or49 | u_cla24_and101;
  assign u_cla24_or51 = u_cla24_pg_logic22_and0 | u_cla24_or50;
  assign u_cla24_pg_logic23_or0 = a[23] | b[23];
  assign u_cla24_pg_logic23_and0 = a[23] & b[23];
  assign u_cla24_pg_logic23_xor0 = a[23] ^ b[23];
  assign u_cla24_xor23 = u_cla24_pg_logic23_xor0 ^ u_cla24_or51;
  assign u_cla24_and102 = u_cla24_or45 & u_cla24_pg_logic22_or0;
  assign u_cla24_and103 = u_cla24_pg_logic23_or0 & u_cla24_pg_logic21_or0;
  assign u_cla24_and104 = u_cla24_and102 & u_cla24_and103;
  assign u_cla24_and105 = u_cla24_and104 & u_cla24_pg_logic20_or0;
  assign u_cla24_and106 = u_cla24_pg_logic20_and0 & u_cla24_pg_logic22_or0;
  assign u_cla24_and107 = u_cla24_pg_logic23_or0 & u_cla24_pg_logic21_or0;
  assign u_cla24_and108 = u_cla24_and106 & u_cla24_and107;
  assign u_cla24_and109 = u_cla24_pg_logic21_and0 & u_cla24_pg_logic23_or0;
  assign u_cla24_and110 = u_cla24_and109 & u_cla24_pg_logic22_or0;
  assign u_cla24_and111 = u_cla24_pg_logic22_and0 & u_cla24_pg_logic23_or0;
  assign u_cla24_or52 = u_cla24_and105 | u_cla24_and110;
  assign u_cla24_or53 = u_cla24_and108 | u_cla24_and111;
  assign u_cla24_or54 = u_cla24_or52 | u_cla24_or53;
  assign u_cla24_or55 = u_cla24_pg_logic23_and0 | u_cla24_or54;

  assign u_cla24_out[0] = u_cla24_pg_logic0_xor0;
  assign u_cla24_out[1] = u_cla24_xor1;
  assign u_cla24_out[2] = u_cla24_xor2;
  assign u_cla24_out[3] = u_cla24_xor3;
  assign u_cla24_out[4] = u_cla24_xor4;
  assign u_cla24_out[5] = u_cla24_xor5;
  assign u_cla24_out[6] = u_cla24_xor6;
  assign u_cla24_out[7] = u_cla24_xor7;
  assign u_cla24_out[8] = u_cla24_xor8;
  assign u_cla24_out[9] = u_cla24_xor9;
  assign u_cla24_out[10] = u_cla24_xor10;
  assign u_cla24_out[11] = u_cla24_xor11;
  assign u_cla24_out[12] = u_cla24_xor12;
  assign u_cla24_out[13] = u_cla24_xor13;
  assign u_cla24_out[14] = u_cla24_xor14;
  assign u_cla24_out[15] = u_cla24_xor15;
  assign u_cla24_out[16] = u_cla24_xor16;
  assign u_cla24_out[17] = u_cla24_xor17;
  assign u_cla24_out[18] = u_cla24_xor18;
  assign u_cla24_out[19] = u_cla24_xor19;
  assign u_cla24_out[20] = u_cla24_xor20;
  assign u_cla24_out[21] = u_cla24_xor21;
  assign u_cla24_out[22] = u_cla24_xor22;
  assign u_cla24_out[23] = u_cla24_xor23;
  assign u_cla24_out[24] = u_cla24_or55;
endmodule