module u_pg_rca8(input [7:0] a, input [7:0] b, output [8:0] u_pg_rca8_out);
  wire u_pg_rca8_pg_fa0_xor0;
  wire u_pg_rca8_pg_fa0_and0;
  wire u_pg_rca8_pg_fa1_xor0;
  wire u_pg_rca8_pg_fa1_and0;
  wire u_pg_rca8_pg_fa1_xor1;
  wire u_pg_rca8_and1;
  wire u_pg_rca8_or1;
  wire u_pg_rca8_pg_fa2_xor0;
  wire u_pg_rca8_pg_fa2_and0;
  wire u_pg_rca8_pg_fa2_xor1;
  wire u_pg_rca8_and2;
  wire u_pg_rca8_or2;
  wire u_pg_rca8_pg_fa3_xor0;
  wire u_pg_rca8_pg_fa3_and0;
  wire u_pg_rca8_pg_fa3_xor1;
  wire u_pg_rca8_and3;
  wire u_pg_rca8_or3;
  wire u_pg_rca8_pg_fa4_xor0;
  wire u_pg_rca8_pg_fa4_and0;
  wire u_pg_rca8_pg_fa4_xor1;
  wire u_pg_rca8_and4;
  wire u_pg_rca8_or4;
  wire u_pg_rca8_pg_fa5_xor0;
  wire u_pg_rca8_pg_fa5_and0;
  wire u_pg_rca8_pg_fa5_xor1;
  wire u_pg_rca8_and5;
  wire u_pg_rca8_or5;
  wire u_pg_rca8_pg_fa6_xor0;
  wire u_pg_rca8_pg_fa6_and0;
  wire u_pg_rca8_pg_fa6_xor1;
  wire u_pg_rca8_and6;
  wire u_pg_rca8_or6;
  wire u_pg_rca8_pg_fa7_xor0;
  wire u_pg_rca8_pg_fa7_and0;
  wire u_pg_rca8_pg_fa7_xor1;
  wire u_pg_rca8_and7;
  wire u_pg_rca8_or7;

  assign u_pg_rca8_pg_fa0_xor0 = a[0] ^ b[0];
  assign u_pg_rca8_pg_fa0_and0 = a[0] & b[0];
  assign u_pg_rca8_pg_fa1_xor0 = a[1] ^ b[1];
  assign u_pg_rca8_pg_fa1_and0 = a[1] & b[1];
  assign u_pg_rca8_pg_fa1_xor1 = u_pg_rca8_pg_fa1_xor0 ^ u_pg_rca8_pg_fa0_and0;
  assign u_pg_rca8_and1 = u_pg_rca8_pg_fa0_and0 & u_pg_rca8_pg_fa1_xor0;
  assign u_pg_rca8_or1 = u_pg_rca8_and1 | u_pg_rca8_pg_fa1_and0;
  assign u_pg_rca8_pg_fa2_xor0 = a[2] ^ b[2];
  assign u_pg_rca8_pg_fa2_and0 = a[2] & b[2];
  assign u_pg_rca8_pg_fa2_xor1 = u_pg_rca8_pg_fa2_xor0 ^ u_pg_rca8_or1;
  assign u_pg_rca8_and2 = u_pg_rca8_or1 & u_pg_rca8_pg_fa2_xor0;
  assign u_pg_rca8_or2 = u_pg_rca8_and2 | u_pg_rca8_pg_fa2_and0;
  assign u_pg_rca8_pg_fa3_xor0 = a[3] ^ b[3];
  assign u_pg_rca8_pg_fa3_and0 = a[3] & b[3];
  assign u_pg_rca8_pg_fa3_xor1 = u_pg_rca8_pg_fa3_xor0 ^ u_pg_rca8_or2;
  assign u_pg_rca8_and3 = u_pg_rca8_or2 & u_pg_rca8_pg_fa3_xor0;
  assign u_pg_rca8_or3 = u_pg_rca8_and3 | u_pg_rca8_pg_fa3_and0;
  assign u_pg_rca8_pg_fa4_xor0 = a[4] ^ b[4];
  assign u_pg_rca8_pg_fa4_and0 = a[4] & b[4];
  assign u_pg_rca8_pg_fa4_xor1 = u_pg_rca8_pg_fa4_xor0 ^ u_pg_rca8_or3;
  assign u_pg_rca8_and4 = u_pg_rca8_or3 & u_pg_rca8_pg_fa4_xor0;
  assign u_pg_rca8_or4 = u_pg_rca8_and4 | u_pg_rca8_pg_fa4_and0;
  assign u_pg_rca8_pg_fa5_xor0 = a[5] ^ b[5];
  assign u_pg_rca8_pg_fa5_and0 = a[5] & b[5];
  assign u_pg_rca8_pg_fa5_xor1 = u_pg_rca8_pg_fa5_xor0 ^ u_pg_rca8_or4;
  assign u_pg_rca8_and5 = u_pg_rca8_or4 & u_pg_rca8_pg_fa5_xor0;
  assign u_pg_rca8_or5 = u_pg_rca8_and5 | u_pg_rca8_pg_fa5_and0;
  assign u_pg_rca8_pg_fa6_xor0 = a[6] ^ b[6];
  assign u_pg_rca8_pg_fa6_and0 = a[6] & b[6];
  assign u_pg_rca8_pg_fa6_xor1 = u_pg_rca8_pg_fa6_xor0 ^ u_pg_rca8_or5;
  assign u_pg_rca8_and6 = u_pg_rca8_or5 & u_pg_rca8_pg_fa6_xor0;
  assign u_pg_rca8_or6 = u_pg_rca8_and6 | u_pg_rca8_pg_fa6_and0;
  assign u_pg_rca8_pg_fa7_xor0 = a[7] ^ b[7];
  assign u_pg_rca8_pg_fa7_and0 = a[7] & b[7];
  assign u_pg_rca8_pg_fa7_xor1 = u_pg_rca8_pg_fa7_xor0 ^ u_pg_rca8_or6;
  assign u_pg_rca8_and7 = u_pg_rca8_or6 & u_pg_rca8_pg_fa7_xor0;
  assign u_pg_rca8_or7 = u_pg_rca8_and7 | u_pg_rca8_pg_fa7_and0;

  assign u_pg_rca8_out[0] = u_pg_rca8_pg_fa0_xor0;
  assign u_pg_rca8_out[1] = u_pg_rca8_pg_fa1_xor1;
  assign u_pg_rca8_out[2] = u_pg_rca8_pg_fa2_xor1;
  assign u_pg_rca8_out[3] = u_pg_rca8_pg_fa3_xor1;
  assign u_pg_rca8_out[4] = u_pg_rca8_pg_fa4_xor1;
  assign u_pg_rca8_out[5] = u_pg_rca8_pg_fa5_xor1;
  assign u_pg_rca8_out[6] = u_pg_rca8_pg_fa6_xor1;
  assign u_pg_rca8_out[7] = u_pg_rca8_pg_fa7_xor1;
  assign u_pg_rca8_out[8] = u_pg_rca8_or7;
endmodule