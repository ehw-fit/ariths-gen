module f_u_dadda_pg_rca16(input [15:0] a, input [15:0] b, output [31:0] out);
  wire a_0;
  wire a_1;
  wire a_2;
  wire a_3;
  wire a_4;
  wire a_5;
  wire a_6;
  wire a_7;
  wire a_8;
  wire a_9;
  wire a_10;
  wire a_11;
  wire a_12;
  wire a_13;
  wire a_14;
  wire a_15;
  wire b_0;
  wire b_1;
  wire b_2;
  wire b_3;
  wire b_4;
  wire b_5;
  wire b_6;
  wire b_7;
  wire b_8;
  wire b_9;
  wire b_10;
  wire b_11;
  wire b_12;
  wire b_13;
  wire b_14;
  wire b_15;
  wire f_u_dadda_pg_rca16_and_13_0_a_13;
  wire f_u_dadda_pg_rca16_and_13_0_b_0;
  wire f_u_dadda_pg_rca16_and_13_0_y0;
  wire f_u_dadda_pg_rca16_and_12_1_a_12;
  wire f_u_dadda_pg_rca16_and_12_1_b_1;
  wire f_u_dadda_pg_rca16_and_12_1_y0;
  wire f_u_dadda_pg_rca16_ha0_f_u_dadda_pg_rca16_and_13_0_y0;
  wire f_u_dadda_pg_rca16_ha0_f_u_dadda_pg_rca16_and_12_1_y0;
  wire f_u_dadda_pg_rca16_ha0_y0;
  wire f_u_dadda_pg_rca16_ha0_y1;
  wire f_u_dadda_pg_rca16_and_14_0_a_14;
  wire f_u_dadda_pg_rca16_and_14_0_b_0;
  wire f_u_dadda_pg_rca16_and_14_0_y0;
  wire f_u_dadda_pg_rca16_and_13_1_a_13;
  wire f_u_dadda_pg_rca16_and_13_1_b_1;
  wire f_u_dadda_pg_rca16_and_13_1_y0;
  wire f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_ha0_y1;
  wire f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_and_14_0_y0;
  wire f_u_dadda_pg_rca16_fa0_y0;
  wire f_u_dadda_pg_rca16_fa0_y1;
  wire f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_and_13_1_y0;
  wire f_u_dadda_pg_rca16_fa0_y2;
  wire f_u_dadda_pg_rca16_fa0_y3;
  wire f_u_dadda_pg_rca16_fa0_y4;
  wire f_u_dadda_pg_rca16_and_12_2_a_12;
  wire f_u_dadda_pg_rca16_and_12_2_b_2;
  wire f_u_dadda_pg_rca16_and_12_2_y0;
  wire f_u_dadda_pg_rca16_and_11_3_a_11;
  wire f_u_dadda_pg_rca16_and_11_3_b_3;
  wire f_u_dadda_pg_rca16_and_11_3_y0;
  wire f_u_dadda_pg_rca16_ha1_f_u_dadda_pg_rca16_and_12_2_y0;
  wire f_u_dadda_pg_rca16_ha1_f_u_dadda_pg_rca16_and_11_3_y0;
  wire f_u_dadda_pg_rca16_ha1_y0;
  wire f_u_dadda_pg_rca16_ha1_y1;
  wire f_u_dadda_pg_rca16_and_15_0_a_15;
  wire f_u_dadda_pg_rca16_and_15_0_b_0;
  wire f_u_dadda_pg_rca16_and_15_0_y0;
  wire f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_ha1_y1;
  wire f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_fa0_y4;
  wire f_u_dadda_pg_rca16_fa1_y0;
  wire f_u_dadda_pg_rca16_fa1_y1;
  wire f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_and_15_0_y0;
  wire f_u_dadda_pg_rca16_fa1_y2;
  wire f_u_dadda_pg_rca16_fa1_y3;
  wire f_u_dadda_pg_rca16_fa1_y4;
  wire f_u_dadda_pg_rca16_and_14_1_a_14;
  wire f_u_dadda_pg_rca16_and_14_1_b_1;
  wire f_u_dadda_pg_rca16_and_14_1_y0;
  wire f_u_dadda_pg_rca16_and_13_2_a_13;
  wire f_u_dadda_pg_rca16_and_13_2_b_2;
  wire f_u_dadda_pg_rca16_and_13_2_y0;
  wire f_u_dadda_pg_rca16_and_12_3_a_12;
  wire f_u_dadda_pg_rca16_and_12_3_b_3;
  wire f_u_dadda_pg_rca16_and_12_3_y0;
  wire f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_14_1_y0;
  wire f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_13_2_y0;
  wire f_u_dadda_pg_rca16_fa2_y0;
  wire f_u_dadda_pg_rca16_fa2_y1;
  wire f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_12_3_y0;
  wire f_u_dadda_pg_rca16_fa2_y2;
  wire f_u_dadda_pg_rca16_fa2_y3;
  wire f_u_dadda_pg_rca16_fa2_y4;
  wire f_u_dadda_pg_rca16_and_11_4_a_11;
  wire f_u_dadda_pg_rca16_and_11_4_b_4;
  wire f_u_dadda_pg_rca16_and_11_4_y0;
  wire f_u_dadda_pg_rca16_and_10_5_a_10;
  wire f_u_dadda_pg_rca16_and_10_5_b_5;
  wire f_u_dadda_pg_rca16_and_10_5_y0;
  wire f_u_dadda_pg_rca16_ha2_f_u_dadda_pg_rca16_and_11_4_y0;
  wire f_u_dadda_pg_rca16_ha2_f_u_dadda_pg_rca16_and_10_5_y0;
  wire f_u_dadda_pg_rca16_ha2_y0;
  wire f_u_dadda_pg_rca16_ha2_y1;
  wire f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_ha2_y1;
  wire f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_fa2_y4;
  wire f_u_dadda_pg_rca16_fa3_y0;
  wire f_u_dadda_pg_rca16_fa3_y1;
  wire f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_fa1_y4;
  wire f_u_dadda_pg_rca16_fa3_y2;
  wire f_u_dadda_pg_rca16_fa3_y3;
  wire f_u_dadda_pg_rca16_fa3_y4;
  wire f_u_dadda_pg_rca16_and_15_1_a_15;
  wire f_u_dadda_pg_rca16_and_15_1_b_1;
  wire f_u_dadda_pg_rca16_and_15_1_y0;
  wire f_u_dadda_pg_rca16_and_14_2_a_14;
  wire f_u_dadda_pg_rca16_and_14_2_b_2;
  wire f_u_dadda_pg_rca16_and_14_2_y0;
  wire f_u_dadda_pg_rca16_and_13_3_a_13;
  wire f_u_dadda_pg_rca16_and_13_3_b_3;
  wire f_u_dadda_pg_rca16_and_13_3_y0;
  wire f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_15_1_y0;
  wire f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_14_2_y0;
  wire f_u_dadda_pg_rca16_fa4_y0;
  wire f_u_dadda_pg_rca16_fa4_y1;
  wire f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_13_3_y0;
  wire f_u_dadda_pg_rca16_fa4_y2;
  wire f_u_dadda_pg_rca16_fa4_y3;
  wire f_u_dadda_pg_rca16_fa4_y4;
  wire f_u_dadda_pg_rca16_and_12_4_a_12;
  wire f_u_dadda_pg_rca16_and_12_4_b_4;
  wire f_u_dadda_pg_rca16_and_12_4_y0;
  wire f_u_dadda_pg_rca16_and_11_5_a_11;
  wire f_u_dadda_pg_rca16_and_11_5_b_5;
  wire f_u_dadda_pg_rca16_and_11_5_y0;
  wire f_u_dadda_pg_rca16_ha3_f_u_dadda_pg_rca16_and_12_4_y0;
  wire f_u_dadda_pg_rca16_ha3_f_u_dadda_pg_rca16_and_11_5_y0;
  wire f_u_dadda_pg_rca16_ha3_y0;
  wire f_u_dadda_pg_rca16_ha3_y1;
  wire f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_ha3_y1;
  wire f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_fa4_y4;
  wire f_u_dadda_pg_rca16_fa5_y0;
  wire f_u_dadda_pg_rca16_fa5_y1;
  wire f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_fa3_y4;
  wire f_u_dadda_pg_rca16_fa5_y2;
  wire f_u_dadda_pg_rca16_fa5_y3;
  wire f_u_dadda_pg_rca16_fa5_y4;
  wire f_u_dadda_pg_rca16_and_15_2_a_15;
  wire f_u_dadda_pg_rca16_and_15_2_b_2;
  wire f_u_dadda_pg_rca16_and_15_2_y0;
  wire f_u_dadda_pg_rca16_and_14_3_a_14;
  wire f_u_dadda_pg_rca16_and_14_3_b_3;
  wire f_u_dadda_pg_rca16_and_14_3_y0;
  wire f_u_dadda_pg_rca16_and_13_4_a_13;
  wire f_u_dadda_pg_rca16_and_13_4_b_4;
  wire f_u_dadda_pg_rca16_and_13_4_y0;
  wire f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_15_2_y0;
  wire f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_14_3_y0;
  wire f_u_dadda_pg_rca16_fa6_y0;
  wire f_u_dadda_pg_rca16_fa6_y1;
  wire f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_13_4_y0;
  wire f_u_dadda_pg_rca16_fa6_y2;
  wire f_u_dadda_pg_rca16_fa6_y3;
  wire f_u_dadda_pg_rca16_fa6_y4;
  wire f_u_dadda_pg_rca16_and_15_3_a_15;
  wire f_u_dadda_pg_rca16_and_15_3_b_3;
  wire f_u_dadda_pg_rca16_and_15_3_y0;
  wire f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_fa6_y4;
  wire f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_fa5_y4;
  wire f_u_dadda_pg_rca16_fa7_y0;
  wire f_u_dadda_pg_rca16_fa7_y1;
  wire f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_and_15_3_y0;
  wire f_u_dadda_pg_rca16_fa7_y2;
  wire f_u_dadda_pg_rca16_fa7_y3;
  wire f_u_dadda_pg_rca16_fa7_y4;
  wire f_u_dadda_pg_rca16_and_4_0_a_4;
  wire f_u_dadda_pg_rca16_and_4_0_b_0;
  wire f_u_dadda_pg_rca16_and_4_0_y0;
  wire f_u_dadda_pg_rca16_and_3_1_a_3;
  wire f_u_dadda_pg_rca16_and_3_1_b_1;
  wire f_u_dadda_pg_rca16_and_3_1_y0;
  wire f_u_dadda_pg_rca16_ha4_f_u_dadda_pg_rca16_and_4_0_y0;
  wire f_u_dadda_pg_rca16_ha4_f_u_dadda_pg_rca16_and_3_1_y0;
  wire f_u_dadda_pg_rca16_ha4_y0;
  wire f_u_dadda_pg_rca16_ha4_y1;
  wire f_u_dadda_pg_rca16_and_5_0_a_5;
  wire f_u_dadda_pg_rca16_and_5_0_b_0;
  wire f_u_dadda_pg_rca16_and_5_0_y0;
  wire f_u_dadda_pg_rca16_and_4_1_a_4;
  wire f_u_dadda_pg_rca16_and_4_1_b_1;
  wire f_u_dadda_pg_rca16_and_4_1_y0;
  wire f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_ha4_y1;
  wire f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_and_5_0_y0;
  wire f_u_dadda_pg_rca16_fa8_y0;
  wire f_u_dadda_pg_rca16_fa8_y1;
  wire f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_and_4_1_y0;
  wire f_u_dadda_pg_rca16_fa8_y2;
  wire f_u_dadda_pg_rca16_fa8_y3;
  wire f_u_dadda_pg_rca16_fa8_y4;
  wire f_u_dadda_pg_rca16_and_3_2_a_3;
  wire f_u_dadda_pg_rca16_and_3_2_b_2;
  wire f_u_dadda_pg_rca16_and_3_2_y0;
  wire f_u_dadda_pg_rca16_and_2_3_a_2;
  wire f_u_dadda_pg_rca16_and_2_3_b_3;
  wire f_u_dadda_pg_rca16_and_2_3_y0;
  wire f_u_dadda_pg_rca16_ha5_f_u_dadda_pg_rca16_and_3_2_y0;
  wire f_u_dadda_pg_rca16_ha5_f_u_dadda_pg_rca16_and_2_3_y0;
  wire f_u_dadda_pg_rca16_ha5_y0;
  wire f_u_dadda_pg_rca16_ha5_y1;
  wire f_u_dadda_pg_rca16_and_6_0_a_6;
  wire f_u_dadda_pg_rca16_and_6_0_b_0;
  wire f_u_dadda_pg_rca16_and_6_0_y0;
  wire f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_ha5_y1;
  wire f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_fa8_y4;
  wire f_u_dadda_pg_rca16_fa9_y0;
  wire f_u_dadda_pg_rca16_fa9_y1;
  wire f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_and_6_0_y0;
  wire f_u_dadda_pg_rca16_fa9_y2;
  wire f_u_dadda_pg_rca16_fa9_y3;
  wire f_u_dadda_pg_rca16_fa9_y4;
  wire f_u_dadda_pg_rca16_and_5_1_a_5;
  wire f_u_dadda_pg_rca16_and_5_1_b_1;
  wire f_u_dadda_pg_rca16_and_5_1_y0;
  wire f_u_dadda_pg_rca16_and_4_2_a_4;
  wire f_u_dadda_pg_rca16_and_4_2_b_2;
  wire f_u_dadda_pg_rca16_and_4_2_y0;
  wire f_u_dadda_pg_rca16_and_3_3_a_3;
  wire f_u_dadda_pg_rca16_and_3_3_b_3;
  wire f_u_dadda_pg_rca16_and_3_3_y0;
  wire f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_5_1_y0;
  wire f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_4_2_y0;
  wire f_u_dadda_pg_rca16_fa10_y0;
  wire f_u_dadda_pg_rca16_fa10_y1;
  wire f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_3_3_y0;
  wire f_u_dadda_pg_rca16_fa10_y2;
  wire f_u_dadda_pg_rca16_fa10_y3;
  wire f_u_dadda_pg_rca16_fa10_y4;
  wire f_u_dadda_pg_rca16_and_2_4_a_2;
  wire f_u_dadda_pg_rca16_and_2_4_b_4;
  wire f_u_dadda_pg_rca16_and_2_4_y0;
  wire f_u_dadda_pg_rca16_and_1_5_a_1;
  wire f_u_dadda_pg_rca16_and_1_5_b_5;
  wire f_u_dadda_pg_rca16_and_1_5_y0;
  wire f_u_dadda_pg_rca16_ha6_f_u_dadda_pg_rca16_and_2_4_y0;
  wire f_u_dadda_pg_rca16_ha6_f_u_dadda_pg_rca16_and_1_5_y0;
  wire f_u_dadda_pg_rca16_ha6_y0;
  wire f_u_dadda_pg_rca16_ha6_y1;
  wire f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_ha6_y1;
  wire f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_fa10_y4;
  wire f_u_dadda_pg_rca16_fa11_y0;
  wire f_u_dadda_pg_rca16_fa11_y1;
  wire f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_fa9_y4;
  wire f_u_dadda_pg_rca16_fa11_y2;
  wire f_u_dadda_pg_rca16_fa11_y3;
  wire f_u_dadda_pg_rca16_fa11_y4;
  wire f_u_dadda_pg_rca16_and_7_0_a_7;
  wire f_u_dadda_pg_rca16_and_7_0_b_0;
  wire f_u_dadda_pg_rca16_and_7_0_y0;
  wire f_u_dadda_pg_rca16_and_6_1_a_6;
  wire f_u_dadda_pg_rca16_and_6_1_b_1;
  wire f_u_dadda_pg_rca16_and_6_1_y0;
  wire f_u_dadda_pg_rca16_and_5_2_a_5;
  wire f_u_dadda_pg_rca16_and_5_2_b_2;
  wire f_u_dadda_pg_rca16_and_5_2_y0;
  wire f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_7_0_y0;
  wire f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_6_1_y0;
  wire f_u_dadda_pg_rca16_fa12_y0;
  wire f_u_dadda_pg_rca16_fa12_y1;
  wire f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_5_2_y0;
  wire f_u_dadda_pg_rca16_fa12_y2;
  wire f_u_dadda_pg_rca16_fa12_y3;
  wire f_u_dadda_pg_rca16_fa12_y4;
  wire f_u_dadda_pg_rca16_and_4_3_a_4;
  wire f_u_dadda_pg_rca16_and_4_3_b_3;
  wire f_u_dadda_pg_rca16_and_4_3_y0;
  wire f_u_dadda_pg_rca16_and_3_4_a_3;
  wire f_u_dadda_pg_rca16_and_3_4_b_4;
  wire f_u_dadda_pg_rca16_and_3_4_y0;
  wire f_u_dadda_pg_rca16_and_2_5_a_2;
  wire f_u_dadda_pg_rca16_and_2_5_b_5;
  wire f_u_dadda_pg_rca16_and_2_5_y0;
  wire f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_4_3_y0;
  wire f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_3_4_y0;
  wire f_u_dadda_pg_rca16_fa13_y0;
  wire f_u_dadda_pg_rca16_fa13_y1;
  wire f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_2_5_y0;
  wire f_u_dadda_pg_rca16_fa13_y2;
  wire f_u_dadda_pg_rca16_fa13_y3;
  wire f_u_dadda_pg_rca16_fa13_y4;
  wire f_u_dadda_pg_rca16_and_1_6_a_1;
  wire f_u_dadda_pg_rca16_and_1_6_b_6;
  wire f_u_dadda_pg_rca16_and_1_6_y0;
  wire f_u_dadda_pg_rca16_and_0_7_a_0;
  wire f_u_dadda_pg_rca16_and_0_7_b_7;
  wire f_u_dadda_pg_rca16_and_0_7_y0;
  wire f_u_dadda_pg_rca16_ha7_f_u_dadda_pg_rca16_and_1_6_y0;
  wire f_u_dadda_pg_rca16_ha7_f_u_dadda_pg_rca16_and_0_7_y0;
  wire f_u_dadda_pg_rca16_ha7_y0;
  wire f_u_dadda_pg_rca16_ha7_y1;
  wire f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_ha7_y1;
  wire f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_fa13_y4;
  wire f_u_dadda_pg_rca16_fa14_y0;
  wire f_u_dadda_pg_rca16_fa14_y1;
  wire f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_fa12_y4;
  wire f_u_dadda_pg_rca16_fa14_y2;
  wire f_u_dadda_pg_rca16_fa14_y3;
  wire f_u_dadda_pg_rca16_fa14_y4;
  wire f_u_dadda_pg_rca16_and_8_0_a_8;
  wire f_u_dadda_pg_rca16_and_8_0_b_0;
  wire f_u_dadda_pg_rca16_and_8_0_y0;
  wire f_u_dadda_pg_rca16_and_7_1_a_7;
  wire f_u_dadda_pg_rca16_and_7_1_b_1;
  wire f_u_dadda_pg_rca16_and_7_1_y0;
  wire f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_fa11_y4;
  wire f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_and_8_0_y0;
  wire f_u_dadda_pg_rca16_fa15_y0;
  wire f_u_dadda_pg_rca16_fa15_y1;
  wire f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_and_7_1_y0;
  wire f_u_dadda_pg_rca16_fa15_y2;
  wire f_u_dadda_pg_rca16_fa15_y3;
  wire f_u_dadda_pg_rca16_fa15_y4;
  wire f_u_dadda_pg_rca16_and_6_2_a_6;
  wire f_u_dadda_pg_rca16_and_6_2_b_2;
  wire f_u_dadda_pg_rca16_and_6_2_y0;
  wire f_u_dadda_pg_rca16_and_5_3_a_5;
  wire f_u_dadda_pg_rca16_and_5_3_b_3;
  wire f_u_dadda_pg_rca16_and_5_3_y0;
  wire f_u_dadda_pg_rca16_and_4_4_a_4;
  wire f_u_dadda_pg_rca16_and_4_4_b_4;
  wire f_u_dadda_pg_rca16_and_4_4_y0;
  wire f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_6_2_y0;
  wire f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_5_3_y0;
  wire f_u_dadda_pg_rca16_fa16_y0;
  wire f_u_dadda_pg_rca16_fa16_y1;
  wire f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_4_4_y0;
  wire f_u_dadda_pg_rca16_fa16_y2;
  wire f_u_dadda_pg_rca16_fa16_y3;
  wire f_u_dadda_pg_rca16_fa16_y4;
  wire f_u_dadda_pg_rca16_and_3_5_a_3;
  wire f_u_dadda_pg_rca16_and_3_5_b_5;
  wire f_u_dadda_pg_rca16_and_3_5_y0;
  wire f_u_dadda_pg_rca16_and_2_6_a_2;
  wire f_u_dadda_pg_rca16_and_2_6_b_6;
  wire f_u_dadda_pg_rca16_and_2_6_y0;
  wire f_u_dadda_pg_rca16_and_1_7_a_1;
  wire f_u_dadda_pg_rca16_and_1_7_b_7;
  wire f_u_dadda_pg_rca16_and_1_7_y0;
  wire f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_3_5_y0;
  wire f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_2_6_y0;
  wire f_u_dadda_pg_rca16_fa17_y0;
  wire f_u_dadda_pg_rca16_fa17_y1;
  wire f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_1_7_y0;
  wire f_u_dadda_pg_rca16_fa17_y2;
  wire f_u_dadda_pg_rca16_fa17_y3;
  wire f_u_dadda_pg_rca16_fa17_y4;
  wire f_u_dadda_pg_rca16_and_0_8_a_0;
  wire f_u_dadda_pg_rca16_and_0_8_b_8;
  wire f_u_dadda_pg_rca16_and_0_8_y0;
  wire f_u_dadda_pg_rca16_ha8_f_u_dadda_pg_rca16_and_0_8_y0;
  wire f_u_dadda_pg_rca16_ha8_f_u_dadda_pg_rca16_fa14_y2;
  wire f_u_dadda_pg_rca16_ha8_y0;
  wire f_u_dadda_pg_rca16_ha8_y1;
  wire f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_ha8_y1;
  wire f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_fa17_y4;
  wire f_u_dadda_pg_rca16_fa18_y0;
  wire f_u_dadda_pg_rca16_fa18_y1;
  wire f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_fa16_y4;
  wire f_u_dadda_pg_rca16_fa18_y2;
  wire f_u_dadda_pg_rca16_fa18_y3;
  wire f_u_dadda_pg_rca16_fa18_y4;
  wire f_u_dadda_pg_rca16_and_9_0_a_9;
  wire f_u_dadda_pg_rca16_and_9_0_b_0;
  wire f_u_dadda_pg_rca16_and_9_0_y0;
  wire f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_fa15_y4;
  wire f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_fa14_y4;
  wire f_u_dadda_pg_rca16_fa19_y0;
  wire f_u_dadda_pg_rca16_fa19_y1;
  wire f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_and_9_0_y0;
  wire f_u_dadda_pg_rca16_fa19_y2;
  wire f_u_dadda_pg_rca16_fa19_y3;
  wire f_u_dadda_pg_rca16_fa19_y4;
  wire f_u_dadda_pg_rca16_and_8_1_a_8;
  wire f_u_dadda_pg_rca16_and_8_1_b_1;
  wire f_u_dadda_pg_rca16_and_8_1_y0;
  wire f_u_dadda_pg_rca16_and_7_2_a_7;
  wire f_u_dadda_pg_rca16_and_7_2_b_2;
  wire f_u_dadda_pg_rca16_and_7_2_y0;
  wire f_u_dadda_pg_rca16_and_6_3_a_6;
  wire f_u_dadda_pg_rca16_and_6_3_b_3;
  wire f_u_dadda_pg_rca16_and_6_3_y0;
  wire f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_8_1_y0;
  wire f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_7_2_y0;
  wire f_u_dadda_pg_rca16_fa20_y0;
  wire f_u_dadda_pg_rca16_fa20_y1;
  wire f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_6_3_y0;
  wire f_u_dadda_pg_rca16_fa20_y2;
  wire f_u_dadda_pg_rca16_fa20_y3;
  wire f_u_dadda_pg_rca16_fa20_y4;
  wire f_u_dadda_pg_rca16_and_5_4_a_5;
  wire f_u_dadda_pg_rca16_and_5_4_b_4;
  wire f_u_dadda_pg_rca16_and_5_4_y0;
  wire f_u_dadda_pg_rca16_and_4_5_a_4;
  wire f_u_dadda_pg_rca16_and_4_5_b_5;
  wire f_u_dadda_pg_rca16_and_4_5_y0;
  wire f_u_dadda_pg_rca16_and_3_6_a_3;
  wire f_u_dadda_pg_rca16_and_3_6_b_6;
  wire f_u_dadda_pg_rca16_and_3_6_y0;
  wire f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_5_4_y0;
  wire f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_4_5_y0;
  wire f_u_dadda_pg_rca16_fa21_y0;
  wire f_u_dadda_pg_rca16_fa21_y1;
  wire f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_3_6_y0;
  wire f_u_dadda_pg_rca16_fa21_y2;
  wire f_u_dadda_pg_rca16_fa21_y3;
  wire f_u_dadda_pg_rca16_fa21_y4;
  wire f_u_dadda_pg_rca16_and_2_7_a_2;
  wire f_u_dadda_pg_rca16_and_2_7_b_7;
  wire f_u_dadda_pg_rca16_and_2_7_y0;
  wire f_u_dadda_pg_rca16_and_1_8_a_1;
  wire f_u_dadda_pg_rca16_and_1_8_b_8;
  wire f_u_dadda_pg_rca16_and_1_8_y0;
  wire f_u_dadda_pg_rca16_and_0_9_a_0;
  wire f_u_dadda_pg_rca16_and_0_9_b_9;
  wire f_u_dadda_pg_rca16_and_0_9_y0;
  wire f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_2_7_y0;
  wire f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_1_8_y0;
  wire f_u_dadda_pg_rca16_fa22_y0;
  wire f_u_dadda_pg_rca16_fa22_y1;
  wire f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_0_9_y0;
  wire f_u_dadda_pg_rca16_fa22_y2;
  wire f_u_dadda_pg_rca16_fa22_y3;
  wire f_u_dadda_pg_rca16_fa22_y4;
  wire f_u_dadda_pg_rca16_ha9_f_u_dadda_pg_rca16_fa18_y2;
  wire f_u_dadda_pg_rca16_ha9_f_u_dadda_pg_rca16_fa19_y2;
  wire f_u_dadda_pg_rca16_ha9_y0;
  wire f_u_dadda_pg_rca16_ha9_y1;
  wire f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_ha9_y1;
  wire f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_fa22_y4;
  wire f_u_dadda_pg_rca16_fa23_y0;
  wire f_u_dadda_pg_rca16_fa23_y1;
  wire f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_fa21_y4;
  wire f_u_dadda_pg_rca16_fa23_y2;
  wire f_u_dadda_pg_rca16_fa23_y3;
  wire f_u_dadda_pg_rca16_fa23_y4;
  wire f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa20_y4;
  wire f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa19_y4;
  wire f_u_dadda_pg_rca16_fa24_y0;
  wire f_u_dadda_pg_rca16_fa24_y1;
  wire f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa18_y4;
  wire f_u_dadda_pg_rca16_fa24_y2;
  wire f_u_dadda_pg_rca16_fa24_y3;
  wire f_u_dadda_pg_rca16_fa24_y4;
  wire f_u_dadda_pg_rca16_and_10_0_a_10;
  wire f_u_dadda_pg_rca16_and_10_0_b_0;
  wire f_u_dadda_pg_rca16_and_10_0_y0;
  wire f_u_dadda_pg_rca16_and_9_1_a_9;
  wire f_u_dadda_pg_rca16_and_9_1_b_1;
  wire f_u_dadda_pg_rca16_and_9_1_y0;
  wire f_u_dadda_pg_rca16_and_8_2_a_8;
  wire f_u_dadda_pg_rca16_and_8_2_b_2;
  wire f_u_dadda_pg_rca16_and_8_2_y0;
  wire f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_10_0_y0;
  wire f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_9_1_y0;
  wire f_u_dadda_pg_rca16_fa25_y0;
  wire f_u_dadda_pg_rca16_fa25_y1;
  wire f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_8_2_y0;
  wire f_u_dadda_pg_rca16_fa25_y2;
  wire f_u_dadda_pg_rca16_fa25_y3;
  wire f_u_dadda_pg_rca16_fa25_y4;
  wire f_u_dadda_pg_rca16_and_7_3_a_7;
  wire f_u_dadda_pg_rca16_and_7_3_b_3;
  wire f_u_dadda_pg_rca16_and_7_3_y0;
  wire f_u_dadda_pg_rca16_and_6_4_a_6;
  wire f_u_dadda_pg_rca16_and_6_4_b_4;
  wire f_u_dadda_pg_rca16_and_6_4_y0;
  wire f_u_dadda_pg_rca16_and_5_5_a_5;
  wire f_u_dadda_pg_rca16_and_5_5_b_5;
  wire f_u_dadda_pg_rca16_and_5_5_y0;
  wire f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_7_3_y0;
  wire f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_6_4_y0;
  wire f_u_dadda_pg_rca16_fa26_y0;
  wire f_u_dadda_pg_rca16_fa26_y1;
  wire f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_5_5_y0;
  wire f_u_dadda_pg_rca16_fa26_y2;
  wire f_u_dadda_pg_rca16_fa26_y3;
  wire f_u_dadda_pg_rca16_fa26_y4;
  wire f_u_dadda_pg_rca16_and_4_6_a_4;
  wire f_u_dadda_pg_rca16_and_4_6_b_6;
  wire f_u_dadda_pg_rca16_and_4_6_y0;
  wire f_u_dadda_pg_rca16_and_3_7_a_3;
  wire f_u_dadda_pg_rca16_and_3_7_b_7;
  wire f_u_dadda_pg_rca16_and_3_7_y0;
  wire f_u_dadda_pg_rca16_and_2_8_a_2;
  wire f_u_dadda_pg_rca16_and_2_8_b_8;
  wire f_u_dadda_pg_rca16_and_2_8_y0;
  wire f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_4_6_y0;
  wire f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_3_7_y0;
  wire f_u_dadda_pg_rca16_fa27_y0;
  wire f_u_dadda_pg_rca16_fa27_y1;
  wire f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_2_8_y0;
  wire f_u_dadda_pg_rca16_fa27_y2;
  wire f_u_dadda_pg_rca16_fa27_y3;
  wire f_u_dadda_pg_rca16_fa27_y4;
  wire f_u_dadda_pg_rca16_and_1_9_a_1;
  wire f_u_dadda_pg_rca16_and_1_9_b_9;
  wire f_u_dadda_pg_rca16_and_1_9_y0;
  wire f_u_dadda_pg_rca16_and_0_10_a_0;
  wire f_u_dadda_pg_rca16_and_0_10_b_10;
  wire f_u_dadda_pg_rca16_and_0_10_y0;
  wire f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_and_1_9_y0;
  wire f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_and_0_10_y0;
  wire f_u_dadda_pg_rca16_fa28_y0;
  wire f_u_dadda_pg_rca16_fa28_y1;
  wire f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_fa23_y2;
  wire f_u_dadda_pg_rca16_fa28_y2;
  wire f_u_dadda_pg_rca16_fa28_y3;
  wire f_u_dadda_pg_rca16_fa28_y4;
  wire f_u_dadda_pg_rca16_ha10_f_u_dadda_pg_rca16_fa24_y2;
  wire f_u_dadda_pg_rca16_ha10_f_u_dadda_pg_rca16_fa25_y2;
  wire f_u_dadda_pg_rca16_ha10_y0;
  wire f_u_dadda_pg_rca16_ha10_y1;
  wire f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_ha10_y1;
  wire f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_fa28_y4;
  wire f_u_dadda_pg_rca16_fa29_y0;
  wire f_u_dadda_pg_rca16_fa29_y1;
  wire f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_fa27_y4;
  wire f_u_dadda_pg_rca16_fa29_y2;
  wire f_u_dadda_pg_rca16_fa29_y3;
  wire f_u_dadda_pg_rca16_fa29_y4;
  wire f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa26_y4;
  wire f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa25_y4;
  wire f_u_dadda_pg_rca16_fa30_y0;
  wire f_u_dadda_pg_rca16_fa30_y1;
  wire f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa24_y4;
  wire f_u_dadda_pg_rca16_fa30_y2;
  wire f_u_dadda_pg_rca16_fa30_y3;
  wire f_u_dadda_pg_rca16_fa30_y4;
  wire f_u_dadda_pg_rca16_and_11_0_a_11;
  wire f_u_dadda_pg_rca16_and_11_0_b_0;
  wire f_u_dadda_pg_rca16_and_11_0_y0;
  wire f_u_dadda_pg_rca16_and_10_1_a_10;
  wire f_u_dadda_pg_rca16_and_10_1_b_1;
  wire f_u_dadda_pg_rca16_and_10_1_y0;
  wire f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_fa23_y4;
  wire f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_and_11_0_y0;
  wire f_u_dadda_pg_rca16_fa31_y0;
  wire f_u_dadda_pg_rca16_fa31_y1;
  wire f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_and_10_1_y0;
  wire f_u_dadda_pg_rca16_fa31_y2;
  wire f_u_dadda_pg_rca16_fa31_y3;
  wire f_u_dadda_pg_rca16_fa31_y4;
  wire f_u_dadda_pg_rca16_and_9_2_a_9;
  wire f_u_dadda_pg_rca16_and_9_2_b_2;
  wire f_u_dadda_pg_rca16_and_9_2_y0;
  wire f_u_dadda_pg_rca16_and_8_3_a_8;
  wire f_u_dadda_pg_rca16_and_8_3_b_3;
  wire f_u_dadda_pg_rca16_and_8_3_y0;
  wire f_u_dadda_pg_rca16_and_7_4_a_7;
  wire f_u_dadda_pg_rca16_and_7_4_b_4;
  wire f_u_dadda_pg_rca16_and_7_4_y0;
  wire f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_9_2_y0;
  wire f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_8_3_y0;
  wire f_u_dadda_pg_rca16_fa32_y0;
  wire f_u_dadda_pg_rca16_fa32_y1;
  wire f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_7_4_y0;
  wire f_u_dadda_pg_rca16_fa32_y2;
  wire f_u_dadda_pg_rca16_fa32_y3;
  wire f_u_dadda_pg_rca16_fa32_y4;
  wire f_u_dadda_pg_rca16_and_6_5_a_6;
  wire f_u_dadda_pg_rca16_and_6_5_b_5;
  wire f_u_dadda_pg_rca16_and_6_5_y0;
  wire f_u_dadda_pg_rca16_and_5_6_a_5;
  wire f_u_dadda_pg_rca16_and_5_6_b_6;
  wire f_u_dadda_pg_rca16_and_5_6_y0;
  wire f_u_dadda_pg_rca16_and_4_7_a_4;
  wire f_u_dadda_pg_rca16_and_4_7_b_7;
  wire f_u_dadda_pg_rca16_and_4_7_y0;
  wire f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_6_5_y0;
  wire f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_5_6_y0;
  wire f_u_dadda_pg_rca16_fa33_y0;
  wire f_u_dadda_pg_rca16_fa33_y1;
  wire f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_4_7_y0;
  wire f_u_dadda_pg_rca16_fa33_y2;
  wire f_u_dadda_pg_rca16_fa33_y3;
  wire f_u_dadda_pg_rca16_fa33_y4;
  wire f_u_dadda_pg_rca16_and_3_8_a_3;
  wire f_u_dadda_pg_rca16_and_3_8_b_8;
  wire f_u_dadda_pg_rca16_and_3_8_y0;
  wire f_u_dadda_pg_rca16_and_2_9_a_2;
  wire f_u_dadda_pg_rca16_and_2_9_b_9;
  wire f_u_dadda_pg_rca16_and_2_9_y0;
  wire f_u_dadda_pg_rca16_and_1_10_a_1;
  wire f_u_dadda_pg_rca16_and_1_10_b_10;
  wire f_u_dadda_pg_rca16_and_1_10_y0;
  wire f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_3_8_y0;
  wire f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_2_9_y0;
  wire f_u_dadda_pg_rca16_fa34_y0;
  wire f_u_dadda_pg_rca16_fa34_y1;
  wire f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_1_10_y0;
  wire f_u_dadda_pg_rca16_fa34_y2;
  wire f_u_dadda_pg_rca16_fa34_y3;
  wire f_u_dadda_pg_rca16_fa34_y4;
  wire f_u_dadda_pg_rca16_and_0_11_a_0;
  wire f_u_dadda_pg_rca16_and_0_11_b_11;
  wire f_u_dadda_pg_rca16_and_0_11_y0;
  wire f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_and_0_11_y0;
  wire f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_fa29_y2;
  wire f_u_dadda_pg_rca16_fa35_y0;
  wire f_u_dadda_pg_rca16_fa35_y1;
  wire f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_fa30_y2;
  wire f_u_dadda_pg_rca16_fa35_y2;
  wire f_u_dadda_pg_rca16_fa35_y3;
  wire f_u_dadda_pg_rca16_fa35_y4;
  wire f_u_dadda_pg_rca16_ha11_f_u_dadda_pg_rca16_fa31_y2;
  wire f_u_dadda_pg_rca16_ha11_f_u_dadda_pg_rca16_fa32_y2;
  wire f_u_dadda_pg_rca16_ha11_y0;
  wire f_u_dadda_pg_rca16_ha11_y1;
  wire f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_ha11_y1;
  wire f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_fa35_y4;
  wire f_u_dadda_pg_rca16_fa36_y0;
  wire f_u_dadda_pg_rca16_fa36_y1;
  wire f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_fa34_y4;
  wire f_u_dadda_pg_rca16_fa36_y2;
  wire f_u_dadda_pg_rca16_fa36_y3;
  wire f_u_dadda_pg_rca16_fa36_y4;
  wire f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa33_y4;
  wire f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa32_y4;
  wire f_u_dadda_pg_rca16_fa37_y0;
  wire f_u_dadda_pg_rca16_fa37_y1;
  wire f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa31_y4;
  wire f_u_dadda_pg_rca16_fa37_y2;
  wire f_u_dadda_pg_rca16_fa37_y3;
  wire f_u_dadda_pg_rca16_fa37_y4;
  wire f_u_dadda_pg_rca16_and_12_0_a_12;
  wire f_u_dadda_pg_rca16_and_12_0_b_0;
  wire f_u_dadda_pg_rca16_and_12_0_y0;
  wire f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_fa30_y4;
  wire f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_fa29_y4;
  wire f_u_dadda_pg_rca16_fa38_y0;
  wire f_u_dadda_pg_rca16_fa38_y1;
  wire f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_and_12_0_y0;
  wire f_u_dadda_pg_rca16_fa38_y2;
  wire f_u_dadda_pg_rca16_fa38_y3;
  wire f_u_dadda_pg_rca16_fa38_y4;
  wire f_u_dadda_pg_rca16_and_11_1_a_11;
  wire f_u_dadda_pg_rca16_and_11_1_b_1;
  wire f_u_dadda_pg_rca16_and_11_1_y0;
  wire f_u_dadda_pg_rca16_and_10_2_a_10;
  wire f_u_dadda_pg_rca16_and_10_2_b_2;
  wire f_u_dadda_pg_rca16_and_10_2_y0;
  wire f_u_dadda_pg_rca16_and_9_3_a_9;
  wire f_u_dadda_pg_rca16_and_9_3_b_3;
  wire f_u_dadda_pg_rca16_and_9_3_y0;
  wire f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_11_1_y0;
  wire f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_10_2_y0;
  wire f_u_dadda_pg_rca16_fa39_y0;
  wire f_u_dadda_pg_rca16_fa39_y1;
  wire f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_9_3_y0;
  wire f_u_dadda_pg_rca16_fa39_y2;
  wire f_u_dadda_pg_rca16_fa39_y3;
  wire f_u_dadda_pg_rca16_fa39_y4;
  wire f_u_dadda_pg_rca16_and_8_4_a_8;
  wire f_u_dadda_pg_rca16_and_8_4_b_4;
  wire f_u_dadda_pg_rca16_and_8_4_y0;
  wire f_u_dadda_pg_rca16_and_7_5_a_7;
  wire f_u_dadda_pg_rca16_and_7_5_b_5;
  wire f_u_dadda_pg_rca16_and_7_5_y0;
  wire f_u_dadda_pg_rca16_and_6_6_a_6;
  wire f_u_dadda_pg_rca16_and_6_6_b_6;
  wire f_u_dadda_pg_rca16_and_6_6_y0;
  wire f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_8_4_y0;
  wire f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_7_5_y0;
  wire f_u_dadda_pg_rca16_fa40_y0;
  wire f_u_dadda_pg_rca16_fa40_y1;
  wire f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_6_6_y0;
  wire f_u_dadda_pg_rca16_fa40_y2;
  wire f_u_dadda_pg_rca16_fa40_y3;
  wire f_u_dadda_pg_rca16_fa40_y4;
  wire f_u_dadda_pg_rca16_and_5_7_a_5;
  wire f_u_dadda_pg_rca16_and_5_7_b_7;
  wire f_u_dadda_pg_rca16_and_5_7_y0;
  wire f_u_dadda_pg_rca16_and_4_8_a_4;
  wire f_u_dadda_pg_rca16_and_4_8_b_8;
  wire f_u_dadda_pg_rca16_and_4_8_y0;
  wire f_u_dadda_pg_rca16_and_3_9_a_3;
  wire f_u_dadda_pg_rca16_and_3_9_b_9;
  wire f_u_dadda_pg_rca16_and_3_9_y0;
  wire f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_5_7_y0;
  wire f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_4_8_y0;
  wire f_u_dadda_pg_rca16_fa41_y0;
  wire f_u_dadda_pg_rca16_fa41_y1;
  wire f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_3_9_y0;
  wire f_u_dadda_pg_rca16_fa41_y2;
  wire f_u_dadda_pg_rca16_fa41_y3;
  wire f_u_dadda_pg_rca16_fa41_y4;
  wire f_u_dadda_pg_rca16_and_2_10_a_2;
  wire f_u_dadda_pg_rca16_and_2_10_b_10;
  wire f_u_dadda_pg_rca16_and_2_10_y0;
  wire f_u_dadda_pg_rca16_and_1_11_a_1;
  wire f_u_dadda_pg_rca16_and_1_11_b_11;
  wire f_u_dadda_pg_rca16_and_1_11_y0;
  wire f_u_dadda_pg_rca16_and_0_12_a_0;
  wire f_u_dadda_pg_rca16_and_0_12_b_12;
  wire f_u_dadda_pg_rca16_and_0_12_y0;
  wire f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_2_10_y0;
  wire f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_1_11_y0;
  wire f_u_dadda_pg_rca16_fa42_y0;
  wire f_u_dadda_pg_rca16_fa42_y1;
  wire f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_0_12_y0;
  wire f_u_dadda_pg_rca16_fa42_y2;
  wire f_u_dadda_pg_rca16_fa42_y3;
  wire f_u_dadda_pg_rca16_fa42_y4;
  wire f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa36_y2;
  wire f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa37_y2;
  wire f_u_dadda_pg_rca16_fa43_y0;
  wire f_u_dadda_pg_rca16_fa43_y1;
  wire f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa38_y2;
  wire f_u_dadda_pg_rca16_fa43_y2;
  wire f_u_dadda_pg_rca16_fa43_y3;
  wire f_u_dadda_pg_rca16_fa43_y4;
  wire f_u_dadda_pg_rca16_ha12_f_u_dadda_pg_rca16_fa39_y2;
  wire f_u_dadda_pg_rca16_ha12_f_u_dadda_pg_rca16_fa40_y2;
  wire f_u_dadda_pg_rca16_ha12_y0;
  wire f_u_dadda_pg_rca16_ha12_y1;
  wire f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_ha12_y1;
  wire f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_fa43_y4;
  wire f_u_dadda_pg_rca16_fa44_y0;
  wire f_u_dadda_pg_rca16_fa44_y1;
  wire f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_fa42_y4;
  wire f_u_dadda_pg_rca16_fa44_y2;
  wire f_u_dadda_pg_rca16_fa44_y3;
  wire f_u_dadda_pg_rca16_fa44_y4;
  wire f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa41_y4;
  wire f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa40_y4;
  wire f_u_dadda_pg_rca16_fa45_y0;
  wire f_u_dadda_pg_rca16_fa45_y1;
  wire f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa39_y4;
  wire f_u_dadda_pg_rca16_fa45_y2;
  wire f_u_dadda_pg_rca16_fa45_y3;
  wire f_u_dadda_pg_rca16_fa45_y4;
  wire f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa38_y4;
  wire f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa37_y4;
  wire f_u_dadda_pg_rca16_fa46_y0;
  wire f_u_dadda_pg_rca16_fa46_y1;
  wire f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa36_y4;
  wire f_u_dadda_pg_rca16_fa46_y2;
  wire f_u_dadda_pg_rca16_fa46_y3;
  wire f_u_dadda_pg_rca16_fa46_y4;
  wire f_u_dadda_pg_rca16_and_11_2_a_11;
  wire f_u_dadda_pg_rca16_and_11_2_b_2;
  wire f_u_dadda_pg_rca16_and_11_2_y0;
  wire f_u_dadda_pg_rca16_and_10_3_a_10;
  wire f_u_dadda_pg_rca16_and_10_3_b_3;
  wire f_u_dadda_pg_rca16_and_10_3_y0;
  wire f_u_dadda_pg_rca16_and_9_4_a_9;
  wire f_u_dadda_pg_rca16_and_9_4_b_4;
  wire f_u_dadda_pg_rca16_and_9_4_y0;
  wire f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_11_2_y0;
  wire f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_10_3_y0;
  wire f_u_dadda_pg_rca16_fa47_y0;
  wire f_u_dadda_pg_rca16_fa47_y1;
  wire f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_9_4_y0;
  wire f_u_dadda_pg_rca16_fa47_y2;
  wire f_u_dadda_pg_rca16_fa47_y3;
  wire f_u_dadda_pg_rca16_fa47_y4;
  wire f_u_dadda_pg_rca16_and_8_5_a_8;
  wire f_u_dadda_pg_rca16_and_8_5_b_5;
  wire f_u_dadda_pg_rca16_and_8_5_y0;
  wire f_u_dadda_pg_rca16_and_7_6_a_7;
  wire f_u_dadda_pg_rca16_and_7_6_b_6;
  wire f_u_dadda_pg_rca16_and_7_6_y0;
  wire f_u_dadda_pg_rca16_and_6_7_a_6;
  wire f_u_dadda_pg_rca16_and_6_7_b_7;
  wire f_u_dadda_pg_rca16_and_6_7_y0;
  wire f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_8_5_y0;
  wire f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_7_6_y0;
  wire f_u_dadda_pg_rca16_fa48_y0;
  wire f_u_dadda_pg_rca16_fa48_y1;
  wire f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_6_7_y0;
  wire f_u_dadda_pg_rca16_fa48_y2;
  wire f_u_dadda_pg_rca16_fa48_y3;
  wire f_u_dadda_pg_rca16_fa48_y4;
  wire f_u_dadda_pg_rca16_and_5_8_a_5;
  wire f_u_dadda_pg_rca16_and_5_8_b_8;
  wire f_u_dadda_pg_rca16_and_5_8_y0;
  wire f_u_dadda_pg_rca16_and_4_9_a_4;
  wire f_u_dadda_pg_rca16_and_4_9_b_9;
  wire f_u_dadda_pg_rca16_and_4_9_y0;
  wire f_u_dadda_pg_rca16_and_3_10_a_3;
  wire f_u_dadda_pg_rca16_and_3_10_b_10;
  wire f_u_dadda_pg_rca16_and_3_10_y0;
  wire f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_5_8_y0;
  wire f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_4_9_y0;
  wire f_u_dadda_pg_rca16_fa49_y0;
  wire f_u_dadda_pg_rca16_fa49_y1;
  wire f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_3_10_y0;
  wire f_u_dadda_pg_rca16_fa49_y2;
  wire f_u_dadda_pg_rca16_fa49_y3;
  wire f_u_dadda_pg_rca16_fa49_y4;
  wire f_u_dadda_pg_rca16_and_2_11_a_2;
  wire f_u_dadda_pg_rca16_and_2_11_b_11;
  wire f_u_dadda_pg_rca16_and_2_11_y0;
  wire f_u_dadda_pg_rca16_and_1_12_a_1;
  wire f_u_dadda_pg_rca16_and_1_12_b_12;
  wire f_u_dadda_pg_rca16_and_1_12_y0;
  wire f_u_dadda_pg_rca16_and_0_13_a_0;
  wire f_u_dadda_pg_rca16_and_0_13_b_13;
  wire f_u_dadda_pg_rca16_and_0_13_y0;
  wire f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_2_11_y0;
  wire f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_1_12_y0;
  wire f_u_dadda_pg_rca16_fa50_y0;
  wire f_u_dadda_pg_rca16_fa50_y1;
  wire f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_0_13_y0;
  wire f_u_dadda_pg_rca16_fa50_y2;
  wire f_u_dadda_pg_rca16_fa50_y3;
  wire f_u_dadda_pg_rca16_fa50_y4;
  wire f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_ha0_y0;
  wire f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_fa44_y2;
  wire f_u_dadda_pg_rca16_fa51_y0;
  wire f_u_dadda_pg_rca16_fa51_y1;
  wire f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_fa45_y2;
  wire f_u_dadda_pg_rca16_fa51_y2;
  wire f_u_dadda_pg_rca16_fa51_y3;
  wire f_u_dadda_pg_rca16_fa51_y4;
  wire f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa46_y2;
  wire f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa47_y2;
  wire f_u_dadda_pg_rca16_fa52_y0;
  wire f_u_dadda_pg_rca16_fa52_y1;
  wire f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa48_y2;
  wire f_u_dadda_pg_rca16_fa52_y2;
  wire f_u_dadda_pg_rca16_fa52_y3;
  wire f_u_dadda_pg_rca16_fa52_y4;
  wire f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa52_y4;
  wire f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa51_y4;
  wire f_u_dadda_pg_rca16_fa53_y0;
  wire f_u_dadda_pg_rca16_fa53_y1;
  wire f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa50_y4;
  wire f_u_dadda_pg_rca16_fa53_y2;
  wire f_u_dadda_pg_rca16_fa53_y3;
  wire f_u_dadda_pg_rca16_fa53_y4;
  wire f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa49_y4;
  wire f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa48_y4;
  wire f_u_dadda_pg_rca16_fa54_y0;
  wire f_u_dadda_pg_rca16_fa54_y1;
  wire f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa47_y4;
  wire f_u_dadda_pg_rca16_fa54_y2;
  wire f_u_dadda_pg_rca16_fa54_y3;
  wire f_u_dadda_pg_rca16_fa54_y4;
  wire f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa46_y4;
  wire f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa45_y4;
  wire f_u_dadda_pg_rca16_fa55_y0;
  wire f_u_dadda_pg_rca16_fa55_y1;
  wire f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa44_y4;
  wire f_u_dadda_pg_rca16_fa55_y2;
  wire f_u_dadda_pg_rca16_fa55_y3;
  wire f_u_dadda_pg_rca16_fa55_y4;
  wire f_u_dadda_pg_rca16_and_10_4_a_10;
  wire f_u_dadda_pg_rca16_and_10_4_b_4;
  wire f_u_dadda_pg_rca16_and_10_4_y0;
  wire f_u_dadda_pg_rca16_and_9_5_a_9;
  wire f_u_dadda_pg_rca16_and_9_5_b_5;
  wire f_u_dadda_pg_rca16_and_9_5_y0;
  wire f_u_dadda_pg_rca16_and_8_6_a_8;
  wire f_u_dadda_pg_rca16_and_8_6_b_6;
  wire f_u_dadda_pg_rca16_and_8_6_y0;
  wire f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_10_4_y0;
  wire f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_9_5_y0;
  wire f_u_dadda_pg_rca16_fa56_y0;
  wire f_u_dadda_pg_rca16_fa56_y1;
  wire f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_8_6_y0;
  wire f_u_dadda_pg_rca16_fa56_y2;
  wire f_u_dadda_pg_rca16_fa56_y3;
  wire f_u_dadda_pg_rca16_fa56_y4;
  wire f_u_dadda_pg_rca16_and_7_7_a_7;
  wire f_u_dadda_pg_rca16_and_7_7_b_7;
  wire f_u_dadda_pg_rca16_and_7_7_y0;
  wire f_u_dadda_pg_rca16_and_6_8_a_6;
  wire f_u_dadda_pg_rca16_and_6_8_b_8;
  wire f_u_dadda_pg_rca16_and_6_8_y0;
  wire f_u_dadda_pg_rca16_and_5_9_a_5;
  wire f_u_dadda_pg_rca16_and_5_9_b_9;
  wire f_u_dadda_pg_rca16_and_5_9_y0;
  wire f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_7_7_y0;
  wire f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_6_8_y0;
  wire f_u_dadda_pg_rca16_fa57_y0;
  wire f_u_dadda_pg_rca16_fa57_y1;
  wire f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_5_9_y0;
  wire f_u_dadda_pg_rca16_fa57_y2;
  wire f_u_dadda_pg_rca16_fa57_y3;
  wire f_u_dadda_pg_rca16_fa57_y4;
  wire f_u_dadda_pg_rca16_and_4_10_a_4;
  wire f_u_dadda_pg_rca16_and_4_10_b_10;
  wire f_u_dadda_pg_rca16_and_4_10_y0;
  wire f_u_dadda_pg_rca16_and_3_11_a_3;
  wire f_u_dadda_pg_rca16_and_3_11_b_11;
  wire f_u_dadda_pg_rca16_and_3_11_y0;
  wire f_u_dadda_pg_rca16_and_2_12_a_2;
  wire f_u_dadda_pg_rca16_and_2_12_b_12;
  wire f_u_dadda_pg_rca16_and_2_12_y0;
  wire f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_4_10_y0;
  wire f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_3_11_y0;
  wire f_u_dadda_pg_rca16_fa58_y0;
  wire f_u_dadda_pg_rca16_fa58_y1;
  wire f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_2_12_y0;
  wire f_u_dadda_pg_rca16_fa58_y2;
  wire f_u_dadda_pg_rca16_fa58_y3;
  wire f_u_dadda_pg_rca16_fa58_y4;
  wire f_u_dadda_pg_rca16_and_1_13_a_1;
  wire f_u_dadda_pg_rca16_and_1_13_b_13;
  wire f_u_dadda_pg_rca16_and_1_13_y0;
  wire f_u_dadda_pg_rca16_and_0_14_a_0;
  wire f_u_dadda_pg_rca16_and_0_14_b_14;
  wire f_u_dadda_pg_rca16_and_0_14_y0;
  wire f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_and_1_13_y0;
  wire f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_and_0_14_y0;
  wire f_u_dadda_pg_rca16_fa59_y0;
  wire f_u_dadda_pg_rca16_fa59_y1;
  wire f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_fa0_y2;
  wire f_u_dadda_pg_rca16_fa59_y2;
  wire f_u_dadda_pg_rca16_fa59_y3;
  wire f_u_dadda_pg_rca16_fa59_y4;
  wire f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_ha1_y0;
  wire f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_fa53_y2;
  wire f_u_dadda_pg_rca16_fa60_y0;
  wire f_u_dadda_pg_rca16_fa60_y1;
  wire f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_fa54_y2;
  wire f_u_dadda_pg_rca16_fa60_y2;
  wire f_u_dadda_pg_rca16_fa60_y3;
  wire f_u_dadda_pg_rca16_fa60_y4;
  wire f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa55_y2;
  wire f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa56_y2;
  wire f_u_dadda_pg_rca16_fa61_y0;
  wire f_u_dadda_pg_rca16_fa61_y1;
  wire f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa57_y2;
  wire f_u_dadda_pg_rca16_fa61_y2;
  wire f_u_dadda_pg_rca16_fa61_y3;
  wire f_u_dadda_pg_rca16_fa61_y4;
  wire f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa61_y4;
  wire f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa60_y4;
  wire f_u_dadda_pg_rca16_fa62_y0;
  wire f_u_dadda_pg_rca16_fa62_y1;
  wire f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa59_y4;
  wire f_u_dadda_pg_rca16_fa62_y2;
  wire f_u_dadda_pg_rca16_fa62_y3;
  wire f_u_dadda_pg_rca16_fa62_y4;
  wire f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa58_y4;
  wire f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa57_y4;
  wire f_u_dadda_pg_rca16_fa63_y0;
  wire f_u_dadda_pg_rca16_fa63_y1;
  wire f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa56_y4;
  wire f_u_dadda_pg_rca16_fa63_y2;
  wire f_u_dadda_pg_rca16_fa63_y3;
  wire f_u_dadda_pg_rca16_fa63_y4;
  wire f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa55_y4;
  wire f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa54_y4;
  wire f_u_dadda_pg_rca16_fa64_y0;
  wire f_u_dadda_pg_rca16_fa64_y1;
  wire f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa53_y4;
  wire f_u_dadda_pg_rca16_fa64_y2;
  wire f_u_dadda_pg_rca16_fa64_y3;
  wire f_u_dadda_pg_rca16_fa64_y4;
  wire f_u_dadda_pg_rca16_and_9_6_a_9;
  wire f_u_dadda_pg_rca16_and_9_6_b_6;
  wire f_u_dadda_pg_rca16_and_9_6_y0;
  wire f_u_dadda_pg_rca16_and_8_7_a_8;
  wire f_u_dadda_pg_rca16_and_8_7_b_7;
  wire f_u_dadda_pg_rca16_and_8_7_y0;
  wire f_u_dadda_pg_rca16_and_7_8_a_7;
  wire f_u_dadda_pg_rca16_and_7_8_b_8;
  wire f_u_dadda_pg_rca16_and_7_8_y0;
  wire f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_9_6_y0;
  wire f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_8_7_y0;
  wire f_u_dadda_pg_rca16_fa65_y0;
  wire f_u_dadda_pg_rca16_fa65_y1;
  wire f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_7_8_y0;
  wire f_u_dadda_pg_rca16_fa65_y2;
  wire f_u_dadda_pg_rca16_fa65_y3;
  wire f_u_dadda_pg_rca16_fa65_y4;
  wire f_u_dadda_pg_rca16_and_6_9_a_6;
  wire f_u_dadda_pg_rca16_and_6_9_b_9;
  wire f_u_dadda_pg_rca16_and_6_9_y0;
  wire f_u_dadda_pg_rca16_and_5_10_a_5;
  wire f_u_dadda_pg_rca16_and_5_10_b_10;
  wire f_u_dadda_pg_rca16_and_5_10_y0;
  wire f_u_dadda_pg_rca16_and_4_11_a_4;
  wire f_u_dadda_pg_rca16_and_4_11_b_11;
  wire f_u_dadda_pg_rca16_and_4_11_y0;
  wire f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_6_9_y0;
  wire f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_5_10_y0;
  wire f_u_dadda_pg_rca16_fa66_y0;
  wire f_u_dadda_pg_rca16_fa66_y1;
  wire f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_4_11_y0;
  wire f_u_dadda_pg_rca16_fa66_y2;
  wire f_u_dadda_pg_rca16_fa66_y3;
  wire f_u_dadda_pg_rca16_fa66_y4;
  wire f_u_dadda_pg_rca16_and_3_12_a_3;
  wire f_u_dadda_pg_rca16_and_3_12_b_12;
  wire f_u_dadda_pg_rca16_and_3_12_y0;
  wire f_u_dadda_pg_rca16_and_2_13_a_2;
  wire f_u_dadda_pg_rca16_and_2_13_b_13;
  wire f_u_dadda_pg_rca16_and_2_13_y0;
  wire f_u_dadda_pg_rca16_and_1_14_a_1;
  wire f_u_dadda_pg_rca16_and_1_14_b_14;
  wire f_u_dadda_pg_rca16_and_1_14_y0;
  wire f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_3_12_y0;
  wire f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_2_13_y0;
  wire f_u_dadda_pg_rca16_fa67_y0;
  wire f_u_dadda_pg_rca16_fa67_y1;
  wire f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_1_14_y0;
  wire f_u_dadda_pg_rca16_fa67_y2;
  wire f_u_dadda_pg_rca16_fa67_y3;
  wire f_u_dadda_pg_rca16_fa67_y4;
  wire f_u_dadda_pg_rca16_and_0_15_a_0;
  wire f_u_dadda_pg_rca16_and_0_15_b_15;
  wire f_u_dadda_pg_rca16_and_0_15_y0;
  wire f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_and_0_15_y0;
  wire f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_fa1_y2;
  wire f_u_dadda_pg_rca16_fa68_y0;
  wire f_u_dadda_pg_rca16_fa68_y1;
  wire f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_fa2_y2;
  wire f_u_dadda_pg_rca16_fa68_y2;
  wire f_u_dadda_pg_rca16_fa68_y3;
  wire f_u_dadda_pg_rca16_fa68_y4;
  wire f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_ha2_y0;
  wire f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_fa62_y2;
  wire f_u_dadda_pg_rca16_fa69_y0;
  wire f_u_dadda_pg_rca16_fa69_y1;
  wire f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_fa63_y2;
  wire f_u_dadda_pg_rca16_fa69_y2;
  wire f_u_dadda_pg_rca16_fa69_y3;
  wire f_u_dadda_pg_rca16_fa69_y4;
  wire f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa64_y2;
  wire f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa65_y2;
  wire f_u_dadda_pg_rca16_fa70_y0;
  wire f_u_dadda_pg_rca16_fa70_y1;
  wire f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa66_y2;
  wire f_u_dadda_pg_rca16_fa70_y2;
  wire f_u_dadda_pg_rca16_fa70_y3;
  wire f_u_dadda_pg_rca16_fa70_y4;
  wire f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa70_y4;
  wire f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa69_y4;
  wire f_u_dadda_pg_rca16_fa71_y0;
  wire f_u_dadda_pg_rca16_fa71_y1;
  wire f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa68_y4;
  wire f_u_dadda_pg_rca16_fa71_y2;
  wire f_u_dadda_pg_rca16_fa71_y3;
  wire f_u_dadda_pg_rca16_fa71_y4;
  wire f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa67_y4;
  wire f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa66_y4;
  wire f_u_dadda_pg_rca16_fa72_y0;
  wire f_u_dadda_pg_rca16_fa72_y1;
  wire f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa65_y4;
  wire f_u_dadda_pg_rca16_fa72_y2;
  wire f_u_dadda_pg_rca16_fa72_y3;
  wire f_u_dadda_pg_rca16_fa72_y4;
  wire f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa64_y4;
  wire f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa63_y4;
  wire f_u_dadda_pg_rca16_fa73_y0;
  wire f_u_dadda_pg_rca16_fa73_y1;
  wire f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa62_y4;
  wire f_u_dadda_pg_rca16_fa73_y2;
  wire f_u_dadda_pg_rca16_fa73_y3;
  wire f_u_dadda_pg_rca16_fa73_y4;
  wire f_u_dadda_pg_rca16_and_10_6_a_10;
  wire f_u_dadda_pg_rca16_and_10_6_b_6;
  wire f_u_dadda_pg_rca16_and_10_6_y0;
  wire f_u_dadda_pg_rca16_and_9_7_a_9;
  wire f_u_dadda_pg_rca16_and_9_7_b_7;
  wire f_u_dadda_pg_rca16_and_9_7_y0;
  wire f_u_dadda_pg_rca16_and_8_8_a_8;
  wire f_u_dadda_pg_rca16_and_8_8_b_8;
  wire f_u_dadda_pg_rca16_and_8_8_y0;
  wire f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_10_6_y0;
  wire f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_9_7_y0;
  wire f_u_dadda_pg_rca16_fa74_y0;
  wire f_u_dadda_pg_rca16_fa74_y1;
  wire f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_8_8_y0;
  wire f_u_dadda_pg_rca16_fa74_y2;
  wire f_u_dadda_pg_rca16_fa74_y3;
  wire f_u_dadda_pg_rca16_fa74_y4;
  wire f_u_dadda_pg_rca16_and_7_9_a_7;
  wire f_u_dadda_pg_rca16_and_7_9_b_9;
  wire f_u_dadda_pg_rca16_and_7_9_y0;
  wire f_u_dadda_pg_rca16_and_6_10_a_6;
  wire f_u_dadda_pg_rca16_and_6_10_b_10;
  wire f_u_dadda_pg_rca16_and_6_10_y0;
  wire f_u_dadda_pg_rca16_and_5_11_a_5;
  wire f_u_dadda_pg_rca16_and_5_11_b_11;
  wire f_u_dadda_pg_rca16_and_5_11_y0;
  wire f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_7_9_y0;
  wire f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_6_10_y0;
  wire f_u_dadda_pg_rca16_fa75_y0;
  wire f_u_dadda_pg_rca16_fa75_y1;
  wire f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_5_11_y0;
  wire f_u_dadda_pg_rca16_fa75_y2;
  wire f_u_dadda_pg_rca16_fa75_y3;
  wire f_u_dadda_pg_rca16_fa75_y4;
  wire f_u_dadda_pg_rca16_and_4_12_a_4;
  wire f_u_dadda_pg_rca16_and_4_12_b_12;
  wire f_u_dadda_pg_rca16_and_4_12_y0;
  wire f_u_dadda_pg_rca16_and_3_13_a_3;
  wire f_u_dadda_pg_rca16_and_3_13_b_13;
  wire f_u_dadda_pg_rca16_and_3_13_y0;
  wire f_u_dadda_pg_rca16_and_2_14_a_2;
  wire f_u_dadda_pg_rca16_and_2_14_b_14;
  wire f_u_dadda_pg_rca16_and_2_14_y0;
  wire f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_4_12_y0;
  wire f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_3_13_y0;
  wire f_u_dadda_pg_rca16_fa76_y0;
  wire f_u_dadda_pg_rca16_fa76_y1;
  wire f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_2_14_y0;
  wire f_u_dadda_pg_rca16_fa76_y2;
  wire f_u_dadda_pg_rca16_fa76_y3;
  wire f_u_dadda_pg_rca16_fa76_y4;
  wire f_u_dadda_pg_rca16_and_1_15_a_1;
  wire f_u_dadda_pg_rca16_and_1_15_b_15;
  wire f_u_dadda_pg_rca16_and_1_15_y0;
  wire f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_and_1_15_y0;
  wire f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_fa3_y2;
  wire f_u_dadda_pg_rca16_fa77_y0;
  wire f_u_dadda_pg_rca16_fa77_y1;
  wire f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_fa4_y2;
  wire f_u_dadda_pg_rca16_fa77_y2;
  wire f_u_dadda_pg_rca16_fa77_y3;
  wire f_u_dadda_pg_rca16_fa77_y4;
  wire f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_ha3_y0;
  wire f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_fa71_y2;
  wire f_u_dadda_pg_rca16_fa78_y0;
  wire f_u_dadda_pg_rca16_fa78_y1;
  wire f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_fa72_y2;
  wire f_u_dadda_pg_rca16_fa78_y2;
  wire f_u_dadda_pg_rca16_fa78_y3;
  wire f_u_dadda_pg_rca16_fa78_y4;
  wire f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa73_y2;
  wire f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa74_y2;
  wire f_u_dadda_pg_rca16_fa79_y0;
  wire f_u_dadda_pg_rca16_fa79_y1;
  wire f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa75_y2;
  wire f_u_dadda_pg_rca16_fa79_y2;
  wire f_u_dadda_pg_rca16_fa79_y3;
  wire f_u_dadda_pg_rca16_fa79_y4;
  wire f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa79_y4;
  wire f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa78_y4;
  wire f_u_dadda_pg_rca16_fa80_y0;
  wire f_u_dadda_pg_rca16_fa80_y1;
  wire f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa77_y4;
  wire f_u_dadda_pg_rca16_fa80_y2;
  wire f_u_dadda_pg_rca16_fa80_y3;
  wire f_u_dadda_pg_rca16_fa80_y4;
  wire f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa76_y4;
  wire f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa75_y4;
  wire f_u_dadda_pg_rca16_fa81_y0;
  wire f_u_dadda_pg_rca16_fa81_y1;
  wire f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa74_y4;
  wire f_u_dadda_pg_rca16_fa81_y2;
  wire f_u_dadda_pg_rca16_fa81_y3;
  wire f_u_dadda_pg_rca16_fa81_y4;
  wire f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa73_y4;
  wire f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa72_y4;
  wire f_u_dadda_pg_rca16_fa82_y0;
  wire f_u_dadda_pg_rca16_fa82_y1;
  wire f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa71_y4;
  wire f_u_dadda_pg_rca16_fa82_y2;
  wire f_u_dadda_pg_rca16_fa82_y3;
  wire f_u_dadda_pg_rca16_fa82_y4;
  wire f_u_dadda_pg_rca16_and_12_5_a_12;
  wire f_u_dadda_pg_rca16_and_12_5_b_5;
  wire f_u_dadda_pg_rca16_and_12_5_y0;
  wire f_u_dadda_pg_rca16_and_11_6_a_11;
  wire f_u_dadda_pg_rca16_and_11_6_b_6;
  wire f_u_dadda_pg_rca16_and_11_6_y0;
  wire f_u_dadda_pg_rca16_and_10_7_a_10;
  wire f_u_dadda_pg_rca16_and_10_7_b_7;
  wire f_u_dadda_pg_rca16_and_10_7_y0;
  wire f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_12_5_y0;
  wire f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_11_6_y0;
  wire f_u_dadda_pg_rca16_fa83_y0;
  wire f_u_dadda_pg_rca16_fa83_y1;
  wire f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_10_7_y0;
  wire f_u_dadda_pg_rca16_fa83_y2;
  wire f_u_dadda_pg_rca16_fa83_y3;
  wire f_u_dadda_pg_rca16_fa83_y4;
  wire f_u_dadda_pg_rca16_and_9_8_a_9;
  wire f_u_dadda_pg_rca16_and_9_8_b_8;
  wire f_u_dadda_pg_rca16_and_9_8_y0;
  wire f_u_dadda_pg_rca16_and_8_9_a_8;
  wire f_u_dadda_pg_rca16_and_8_9_b_9;
  wire f_u_dadda_pg_rca16_and_8_9_y0;
  wire f_u_dadda_pg_rca16_and_7_10_a_7;
  wire f_u_dadda_pg_rca16_and_7_10_b_10;
  wire f_u_dadda_pg_rca16_and_7_10_y0;
  wire f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_9_8_y0;
  wire f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_8_9_y0;
  wire f_u_dadda_pg_rca16_fa84_y0;
  wire f_u_dadda_pg_rca16_fa84_y1;
  wire f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_7_10_y0;
  wire f_u_dadda_pg_rca16_fa84_y2;
  wire f_u_dadda_pg_rca16_fa84_y3;
  wire f_u_dadda_pg_rca16_fa84_y4;
  wire f_u_dadda_pg_rca16_and_6_11_a_6;
  wire f_u_dadda_pg_rca16_and_6_11_b_11;
  wire f_u_dadda_pg_rca16_and_6_11_y0;
  wire f_u_dadda_pg_rca16_and_5_12_a_5;
  wire f_u_dadda_pg_rca16_and_5_12_b_12;
  wire f_u_dadda_pg_rca16_and_5_12_y0;
  wire f_u_dadda_pg_rca16_and_4_13_a_4;
  wire f_u_dadda_pg_rca16_and_4_13_b_13;
  wire f_u_dadda_pg_rca16_and_4_13_y0;
  wire f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_6_11_y0;
  wire f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_5_12_y0;
  wire f_u_dadda_pg_rca16_fa85_y0;
  wire f_u_dadda_pg_rca16_fa85_y1;
  wire f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_4_13_y0;
  wire f_u_dadda_pg_rca16_fa85_y2;
  wire f_u_dadda_pg_rca16_fa85_y3;
  wire f_u_dadda_pg_rca16_fa85_y4;
  wire f_u_dadda_pg_rca16_and_3_14_a_3;
  wire f_u_dadda_pg_rca16_and_3_14_b_14;
  wire f_u_dadda_pg_rca16_and_3_14_y0;
  wire f_u_dadda_pg_rca16_and_2_15_a_2;
  wire f_u_dadda_pg_rca16_and_2_15_b_15;
  wire f_u_dadda_pg_rca16_and_2_15_y0;
  wire f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_and_3_14_y0;
  wire f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_and_2_15_y0;
  wire f_u_dadda_pg_rca16_fa86_y0;
  wire f_u_dadda_pg_rca16_fa86_y1;
  wire f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_fa5_y2;
  wire f_u_dadda_pg_rca16_fa86_y2;
  wire f_u_dadda_pg_rca16_fa86_y3;
  wire f_u_dadda_pg_rca16_fa86_y4;
  wire f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa6_y2;
  wire f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa80_y2;
  wire f_u_dadda_pg_rca16_fa87_y0;
  wire f_u_dadda_pg_rca16_fa87_y1;
  wire f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa81_y2;
  wire f_u_dadda_pg_rca16_fa87_y2;
  wire f_u_dadda_pg_rca16_fa87_y3;
  wire f_u_dadda_pg_rca16_fa87_y4;
  wire f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa82_y2;
  wire f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa83_y2;
  wire f_u_dadda_pg_rca16_fa88_y0;
  wire f_u_dadda_pg_rca16_fa88_y1;
  wire f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa84_y2;
  wire f_u_dadda_pg_rca16_fa88_y2;
  wire f_u_dadda_pg_rca16_fa88_y3;
  wire f_u_dadda_pg_rca16_fa88_y4;
  wire f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa88_y4;
  wire f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa87_y4;
  wire f_u_dadda_pg_rca16_fa89_y0;
  wire f_u_dadda_pg_rca16_fa89_y1;
  wire f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa86_y4;
  wire f_u_dadda_pg_rca16_fa89_y2;
  wire f_u_dadda_pg_rca16_fa89_y3;
  wire f_u_dadda_pg_rca16_fa89_y4;
  wire f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa85_y4;
  wire f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa84_y4;
  wire f_u_dadda_pg_rca16_fa90_y0;
  wire f_u_dadda_pg_rca16_fa90_y1;
  wire f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa83_y4;
  wire f_u_dadda_pg_rca16_fa90_y2;
  wire f_u_dadda_pg_rca16_fa90_y3;
  wire f_u_dadda_pg_rca16_fa90_y4;
  wire f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa82_y4;
  wire f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa81_y4;
  wire f_u_dadda_pg_rca16_fa91_y0;
  wire f_u_dadda_pg_rca16_fa91_y1;
  wire f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa80_y4;
  wire f_u_dadda_pg_rca16_fa91_y2;
  wire f_u_dadda_pg_rca16_fa91_y3;
  wire f_u_dadda_pg_rca16_fa91_y4;
  wire f_u_dadda_pg_rca16_and_14_4_a_14;
  wire f_u_dadda_pg_rca16_and_14_4_b_4;
  wire f_u_dadda_pg_rca16_and_14_4_y0;
  wire f_u_dadda_pg_rca16_and_13_5_a_13;
  wire f_u_dadda_pg_rca16_and_13_5_b_5;
  wire f_u_dadda_pg_rca16_and_13_5_y0;
  wire f_u_dadda_pg_rca16_and_12_6_a_12;
  wire f_u_dadda_pg_rca16_and_12_6_b_6;
  wire f_u_dadda_pg_rca16_and_12_6_y0;
  wire f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_14_4_y0;
  wire f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_13_5_y0;
  wire f_u_dadda_pg_rca16_fa92_y0;
  wire f_u_dadda_pg_rca16_fa92_y1;
  wire f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_12_6_y0;
  wire f_u_dadda_pg_rca16_fa92_y2;
  wire f_u_dadda_pg_rca16_fa92_y3;
  wire f_u_dadda_pg_rca16_fa92_y4;
  wire f_u_dadda_pg_rca16_and_11_7_a_11;
  wire f_u_dadda_pg_rca16_and_11_7_b_7;
  wire f_u_dadda_pg_rca16_and_11_7_y0;
  wire f_u_dadda_pg_rca16_and_10_8_a_10;
  wire f_u_dadda_pg_rca16_and_10_8_b_8;
  wire f_u_dadda_pg_rca16_and_10_8_y0;
  wire f_u_dadda_pg_rca16_and_9_9_a_9;
  wire f_u_dadda_pg_rca16_and_9_9_b_9;
  wire f_u_dadda_pg_rca16_and_9_9_y0;
  wire f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_11_7_y0;
  wire f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_10_8_y0;
  wire f_u_dadda_pg_rca16_fa93_y0;
  wire f_u_dadda_pg_rca16_fa93_y1;
  wire f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_9_9_y0;
  wire f_u_dadda_pg_rca16_fa93_y2;
  wire f_u_dadda_pg_rca16_fa93_y3;
  wire f_u_dadda_pg_rca16_fa93_y4;
  wire f_u_dadda_pg_rca16_and_8_10_a_8;
  wire f_u_dadda_pg_rca16_and_8_10_b_10;
  wire f_u_dadda_pg_rca16_and_8_10_y0;
  wire f_u_dadda_pg_rca16_and_7_11_a_7;
  wire f_u_dadda_pg_rca16_and_7_11_b_11;
  wire f_u_dadda_pg_rca16_and_7_11_y0;
  wire f_u_dadda_pg_rca16_and_6_12_a_6;
  wire f_u_dadda_pg_rca16_and_6_12_b_12;
  wire f_u_dadda_pg_rca16_and_6_12_y0;
  wire f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_8_10_y0;
  wire f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_7_11_y0;
  wire f_u_dadda_pg_rca16_fa94_y0;
  wire f_u_dadda_pg_rca16_fa94_y1;
  wire f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_6_12_y0;
  wire f_u_dadda_pg_rca16_fa94_y2;
  wire f_u_dadda_pg_rca16_fa94_y3;
  wire f_u_dadda_pg_rca16_fa94_y4;
  wire f_u_dadda_pg_rca16_and_5_13_a_5;
  wire f_u_dadda_pg_rca16_and_5_13_b_13;
  wire f_u_dadda_pg_rca16_and_5_13_y0;
  wire f_u_dadda_pg_rca16_and_4_14_a_4;
  wire f_u_dadda_pg_rca16_and_4_14_b_14;
  wire f_u_dadda_pg_rca16_and_4_14_y0;
  wire f_u_dadda_pg_rca16_and_3_15_a_3;
  wire f_u_dadda_pg_rca16_and_3_15_b_15;
  wire f_u_dadda_pg_rca16_and_3_15_y0;
  wire f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_5_13_y0;
  wire f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_4_14_y0;
  wire f_u_dadda_pg_rca16_fa95_y0;
  wire f_u_dadda_pg_rca16_fa95_y1;
  wire f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_3_15_y0;
  wire f_u_dadda_pg_rca16_fa95_y2;
  wire f_u_dadda_pg_rca16_fa95_y3;
  wire f_u_dadda_pg_rca16_fa95_y4;
  wire f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa7_y2;
  wire f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa89_y2;
  wire f_u_dadda_pg_rca16_fa96_y0;
  wire f_u_dadda_pg_rca16_fa96_y1;
  wire f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa90_y2;
  wire f_u_dadda_pg_rca16_fa96_y2;
  wire f_u_dadda_pg_rca16_fa96_y3;
  wire f_u_dadda_pg_rca16_fa96_y4;
  wire f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa91_y2;
  wire f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa92_y2;
  wire f_u_dadda_pg_rca16_fa97_y0;
  wire f_u_dadda_pg_rca16_fa97_y1;
  wire f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa93_y2;
  wire f_u_dadda_pg_rca16_fa97_y2;
  wire f_u_dadda_pg_rca16_fa97_y3;
  wire f_u_dadda_pg_rca16_fa97_y4;
  wire f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa97_y4;
  wire f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa96_y4;
  wire f_u_dadda_pg_rca16_fa98_y0;
  wire f_u_dadda_pg_rca16_fa98_y1;
  wire f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa95_y4;
  wire f_u_dadda_pg_rca16_fa98_y2;
  wire f_u_dadda_pg_rca16_fa98_y3;
  wire f_u_dadda_pg_rca16_fa98_y4;
  wire f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa94_y4;
  wire f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa93_y4;
  wire f_u_dadda_pg_rca16_fa99_y0;
  wire f_u_dadda_pg_rca16_fa99_y1;
  wire f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa92_y4;
  wire f_u_dadda_pg_rca16_fa99_y2;
  wire f_u_dadda_pg_rca16_fa99_y3;
  wire f_u_dadda_pg_rca16_fa99_y4;
  wire f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa91_y4;
  wire f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa90_y4;
  wire f_u_dadda_pg_rca16_fa100_y0;
  wire f_u_dadda_pg_rca16_fa100_y1;
  wire f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa89_y4;
  wire f_u_dadda_pg_rca16_fa100_y2;
  wire f_u_dadda_pg_rca16_fa100_y3;
  wire f_u_dadda_pg_rca16_fa100_y4;
  wire f_u_dadda_pg_rca16_and_15_4_a_15;
  wire f_u_dadda_pg_rca16_and_15_4_b_4;
  wire f_u_dadda_pg_rca16_and_15_4_y0;
  wire f_u_dadda_pg_rca16_and_14_5_a_14;
  wire f_u_dadda_pg_rca16_and_14_5_b_5;
  wire f_u_dadda_pg_rca16_and_14_5_y0;
  wire f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_fa7_y4;
  wire f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_and_15_4_y0;
  wire f_u_dadda_pg_rca16_fa101_y0;
  wire f_u_dadda_pg_rca16_fa101_y1;
  wire f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_and_14_5_y0;
  wire f_u_dadda_pg_rca16_fa101_y2;
  wire f_u_dadda_pg_rca16_fa101_y3;
  wire f_u_dadda_pg_rca16_fa101_y4;
  wire f_u_dadda_pg_rca16_and_13_6_a_13;
  wire f_u_dadda_pg_rca16_and_13_6_b_6;
  wire f_u_dadda_pg_rca16_and_13_6_y0;
  wire f_u_dadda_pg_rca16_and_12_7_a_12;
  wire f_u_dadda_pg_rca16_and_12_7_b_7;
  wire f_u_dadda_pg_rca16_and_12_7_y0;
  wire f_u_dadda_pg_rca16_and_11_8_a_11;
  wire f_u_dadda_pg_rca16_and_11_8_b_8;
  wire f_u_dadda_pg_rca16_and_11_8_y0;
  wire f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_13_6_y0;
  wire f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_12_7_y0;
  wire f_u_dadda_pg_rca16_fa102_y0;
  wire f_u_dadda_pg_rca16_fa102_y1;
  wire f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_11_8_y0;
  wire f_u_dadda_pg_rca16_fa102_y2;
  wire f_u_dadda_pg_rca16_fa102_y3;
  wire f_u_dadda_pg_rca16_fa102_y4;
  wire f_u_dadda_pg_rca16_and_10_9_a_10;
  wire f_u_dadda_pg_rca16_and_10_9_b_9;
  wire f_u_dadda_pg_rca16_and_10_9_y0;
  wire f_u_dadda_pg_rca16_and_9_10_a_9;
  wire f_u_dadda_pg_rca16_and_9_10_b_10;
  wire f_u_dadda_pg_rca16_and_9_10_y0;
  wire f_u_dadda_pg_rca16_and_8_11_a_8;
  wire f_u_dadda_pg_rca16_and_8_11_b_11;
  wire f_u_dadda_pg_rca16_and_8_11_y0;
  wire f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_10_9_y0;
  wire f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_9_10_y0;
  wire f_u_dadda_pg_rca16_fa103_y0;
  wire f_u_dadda_pg_rca16_fa103_y1;
  wire f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_8_11_y0;
  wire f_u_dadda_pg_rca16_fa103_y2;
  wire f_u_dadda_pg_rca16_fa103_y3;
  wire f_u_dadda_pg_rca16_fa103_y4;
  wire f_u_dadda_pg_rca16_and_7_12_a_7;
  wire f_u_dadda_pg_rca16_and_7_12_b_12;
  wire f_u_dadda_pg_rca16_and_7_12_y0;
  wire f_u_dadda_pg_rca16_and_6_13_a_6;
  wire f_u_dadda_pg_rca16_and_6_13_b_13;
  wire f_u_dadda_pg_rca16_and_6_13_y0;
  wire f_u_dadda_pg_rca16_and_5_14_a_5;
  wire f_u_dadda_pg_rca16_and_5_14_b_14;
  wire f_u_dadda_pg_rca16_and_5_14_y0;
  wire f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_7_12_y0;
  wire f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_6_13_y0;
  wire f_u_dadda_pg_rca16_fa104_y0;
  wire f_u_dadda_pg_rca16_fa104_y1;
  wire f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_5_14_y0;
  wire f_u_dadda_pg_rca16_fa104_y2;
  wire f_u_dadda_pg_rca16_fa104_y3;
  wire f_u_dadda_pg_rca16_fa104_y4;
  wire f_u_dadda_pg_rca16_and_4_15_a_4;
  wire f_u_dadda_pg_rca16_and_4_15_b_15;
  wire f_u_dadda_pg_rca16_and_4_15_y0;
  wire f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_and_4_15_y0;
  wire f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_fa98_y2;
  wire f_u_dadda_pg_rca16_fa105_y0;
  wire f_u_dadda_pg_rca16_fa105_y1;
  wire f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_fa99_y2;
  wire f_u_dadda_pg_rca16_fa105_y2;
  wire f_u_dadda_pg_rca16_fa105_y3;
  wire f_u_dadda_pg_rca16_fa105_y4;
  wire f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa100_y2;
  wire f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa101_y2;
  wire f_u_dadda_pg_rca16_fa106_y0;
  wire f_u_dadda_pg_rca16_fa106_y1;
  wire f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa102_y2;
  wire f_u_dadda_pg_rca16_fa106_y2;
  wire f_u_dadda_pg_rca16_fa106_y3;
  wire f_u_dadda_pg_rca16_fa106_y4;
  wire f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa106_y4;
  wire f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa105_y4;
  wire f_u_dadda_pg_rca16_fa107_y0;
  wire f_u_dadda_pg_rca16_fa107_y1;
  wire f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa104_y4;
  wire f_u_dadda_pg_rca16_fa107_y2;
  wire f_u_dadda_pg_rca16_fa107_y3;
  wire f_u_dadda_pg_rca16_fa107_y4;
  wire f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa103_y4;
  wire f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa102_y4;
  wire f_u_dadda_pg_rca16_fa108_y0;
  wire f_u_dadda_pg_rca16_fa108_y1;
  wire f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa101_y4;
  wire f_u_dadda_pg_rca16_fa108_y2;
  wire f_u_dadda_pg_rca16_fa108_y3;
  wire f_u_dadda_pg_rca16_fa108_y4;
  wire f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa100_y4;
  wire f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa99_y4;
  wire f_u_dadda_pg_rca16_fa109_y0;
  wire f_u_dadda_pg_rca16_fa109_y1;
  wire f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa98_y4;
  wire f_u_dadda_pg_rca16_fa109_y2;
  wire f_u_dadda_pg_rca16_fa109_y3;
  wire f_u_dadda_pg_rca16_fa109_y4;
  wire f_u_dadda_pg_rca16_and_15_5_a_15;
  wire f_u_dadda_pg_rca16_and_15_5_b_5;
  wire f_u_dadda_pg_rca16_and_15_5_y0;
  wire f_u_dadda_pg_rca16_and_14_6_a_14;
  wire f_u_dadda_pg_rca16_and_14_6_b_6;
  wire f_u_dadda_pg_rca16_and_14_6_y0;
  wire f_u_dadda_pg_rca16_and_13_7_a_13;
  wire f_u_dadda_pg_rca16_and_13_7_b_7;
  wire f_u_dadda_pg_rca16_and_13_7_y0;
  wire f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_15_5_y0;
  wire f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_14_6_y0;
  wire f_u_dadda_pg_rca16_fa110_y0;
  wire f_u_dadda_pg_rca16_fa110_y1;
  wire f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_13_7_y0;
  wire f_u_dadda_pg_rca16_fa110_y2;
  wire f_u_dadda_pg_rca16_fa110_y3;
  wire f_u_dadda_pg_rca16_fa110_y4;
  wire f_u_dadda_pg_rca16_and_12_8_a_12;
  wire f_u_dadda_pg_rca16_and_12_8_b_8;
  wire f_u_dadda_pg_rca16_and_12_8_y0;
  wire f_u_dadda_pg_rca16_and_11_9_a_11;
  wire f_u_dadda_pg_rca16_and_11_9_b_9;
  wire f_u_dadda_pg_rca16_and_11_9_y0;
  wire f_u_dadda_pg_rca16_and_10_10_a_10;
  wire f_u_dadda_pg_rca16_and_10_10_b_10;
  wire f_u_dadda_pg_rca16_and_10_10_y0;
  wire f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_12_8_y0;
  wire f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_11_9_y0;
  wire f_u_dadda_pg_rca16_fa111_y0;
  wire f_u_dadda_pg_rca16_fa111_y1;
  wire f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_10_10_y0;
  wire f_u_dadda_pg_rca16_fa111_y2;
  wire f_u_dadda_pg_rca16_fa111_y3;
  wire f_u_dadda_pg_rca16_fa111_y4;
  wire f_u_dadda_pg_rca16_and_9_11_a_9;
  wire f_u_dadda_pg_rca16_and_9_11_b_11;
  wire f_u_dadda_pg_rca16_and_9_11_y0;
  wire f_u_dadda_pg_rca16_and_8_12_a_8;
  wire f_u_dadda_pg_rca16_and_8_12_b_12;
  wire f_u_dadda_pg_rca16_and_8_12_y0;
  wire f_u_dadda_pg_rca16_and_7_13_a_7;
  wire f_u_dadda_pg_rca16_and_7_13_b_13;
  wire f_u_dadda_pg_rca16_and_7_13_y0;
  wire f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_9_11_y0;
  wire f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_8_12_y0;
  wire f_u_dadda_pg_rca16_fa112_y0;
  wire f_u_dadda_pg_rca16_fa112_y1;
  wire f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_7_13_y0;
  wire f_u_dadda_pg_rca16_fa112_y2;
  wire f_u_dadda_pg_rca16_fa112_y3;
  wire f_u_dadda_pg_rca16_fa112_y4;
  wire f_u_dadda_pg_rca16_and_6_14_a_6;
  wire f_u_dadda_pg_rca16_and_6_14_b_14;
  wire f_u_dadda_pg_rca16_and_6_14_y0;
  wire f_u_dadda_pg_rca16_and_5_15_a_5;
  wire f_u_dadda_pg_rca16_and_5_15_b_15;
  wire f_u_dadda_pg_rca16_and_5_15_y0;
  wire f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_and_6_14_y0;
  wire f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_and_5_15_y0;
  wire f_u_dadda_pg_rca16_fa113_y0;
  wire f_u_dadda_pg_rca16_fa113_y1;
  wire f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_fa107_y2;
  wire f_u_dadda_pg_rca16_fa113_y2;
  wire f_u_dadda_pg_rca16_fa113_y3;
  wire f_u_dadda_pg_rca16_fa113_y4;
  wire f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa108_y2;
  wire f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa109_y2;
  wire f_u_dadda_pg_rca16_fa114_y0;
  wire f_u_dadda_pg_rca16_fa114_y1;
  wire f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa110_y2;
  wire f_u_dadda_pg_rca16_fa114_y2;
  wire f_u_dadda_pg_rca16_fa114_y3;
  wire f_u_dadda_pg_rca16_fa114_y4;
  wire f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa114_y4;
  wire f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa113_y4;
  wire f_u_dadda_pg_rca16_fa115_y0;
  wire f_u_dadda_pg_rca16_fa115_y1;
  wire f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa112_y4;
  wire f_u_dadda_pg_rca16_fa115_y2;
  wire f_u_dadda_pg_rca16_fa115_y3;
  wire f_u_dadda_pg_rca16_fa115_y4;
  wire f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa111_y4;
  wire f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa110_y4;
  wire f_u_dadda_pg_rca16_fa116_y0;
  wire f_u_dadda_pg_rca16_fa116_y1;
  wire f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa109_y4;
  wire f_u_dadda_pg_rca16_fa116_y2;
  wire f_u_dadda_pg_rca16_fa116_y3;
  wire f_u_dadda_pg_rca16_fa116_y4;
  wire f_u_dadda_pg_rca16_and_15_6_a_15;
  wire f_u_dadda_pg_rca16_and_15_6_b_6;
  wire f_u_dadda_pg_rca16_and_15_6_y0;
  wire f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_fa108_y4;
  wire f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_fa107_y4;
  wire f_u_dadda_pg_rca16_fa117_y0;
  wire f_u_dadda_pg_rca16_fa117_y1;
  wire f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_and_15_6_y0;
  wire f_u_dadda_pg_rca16_fa117_y2;
  wire f_u_dadda_pg_rca16_fa117_y3;
  wire f_u_dadda_pg_rca16_fa117_y4;
  wire f_u_dadda_pg_rca16_and_14_7_a_14;
  wire f_u_dadda_pg_rca16_and_14_7_b_7;
  wire f_u_dadda_pg_rca16_and_14_7_y0;
  wire f_u_dadda_pg_rca16_and_13_8_a_13;
  wire f_u_dadda_pg_rca16_and_13_8_b_8;
  wire f_u_dadda_pg_rca16_and_13_8_y0;
  wire f_u_dadda_pg_rca16_and_12_9_a_12;
  wire f_u_dadda_pg_rca16_and_12_9_b_9;
  wire f_u_dadda_pg_rca16_and_12_9_y0;
  wire f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_14_7_y0;
  wire f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_13_8_y0;
  wire f_u_dadda_pg_rca16_fa118_y0;
  wire f_u_dadda_pg_rca16_fa118_y1;
  wire f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_12_9_y0;
  wire f_u_dadda_pg_rca16_fa118_y2;
  wire f_u_dadda_pg_rca16_fa118_y3;
  wire f_u_dadda_pg_rca16_fa118_y4;
  wire f_u_dadda_pg_rca16_and_11_10_a_11;
  wire f_u_dadda_pg_rca16_and_11_10_b_10;
  wire f_u_dadda_pg_rca16_and_11_10_y0;
  wire f_u_dadda_pg_rca16_and_10_11_a_10;
  wire f_u_dadda_pg_rca16_and_10_11_b_11;
  wire f_u_dadda_pg_rca16_and_10_11_y0;
  wire f_u_dadda_pg_rca16_and_9_12_a_9;
  wire f_u_dadda_pg_rca16_and_9_12_b_12;
  wire f_u_dadda_pg_rca16_and_9_12_y0;
  wire f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_11_10_y0;
  wire f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_10_11_y0;
  wire f_u_dadda_pg_rca16_fa119_y0;
  wire f_u_dadda_pg_rca16_fa119_y1;
  wire f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_9_12_y0;
  wire f_u_dadda_pg_rca16_fa119_y2;
  wire f_u_dadda_pg_rca16_fa119_y3;
  wire f_u_dadda_pg_rca16_fa119_y4;
  wire f_u_dadda_pg_rca16_and_8_13_a_8;
  wire f_u_dadda_pg_rca16_and_8_13_b_13;
  wire f_u_dadda_pg_rca16_and_8_13_y0;
  wire f_u_dadda_pg_rca16_and_7_14_a_7;
  wire f_u_dadda_pg_rca16_and_7_14_b_14;
  wire f_u_dadda_pg_rca16_and_7_14_y0;
  wire f_u_dadda_pg_rca16_and_6_15_a_6;
  wire f_u_dadda_pg_rca16_and_6_15_b_15;
  wire f_u_dadda_pg_rca16_and_6_15_y0;
  wire f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_8_13_y0;
  wire f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_7_14_y0;
  wire f_u_dadda_pg_rca16_fa120_y0;
  wire f_u_dadda_pg_rca16_fa120_y1;
  wire f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_6_15_y0;
  wire f_u_dadda_pg_rca16_fa120_y2;
  wire f_u_dadda_pg_rca16_fa120_y3;
  wire f_u_dadda_pg_rca16_fa120_y4;
  wire f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa115_y2;
  wire f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa116_y2;
  wire f_u_dadda_pg_rca16_fa121_y0;
  wire f_u_dadda_pg_rca16_fa121_y1;
  wire f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa117_y2;
  wire f_u_dadda_pg_rca16_fa121_y2;
  wire f_u_dadda_pg_rca16_fa121_y3;
  wire f_u_dadda_pg_rca16_fa121_y4;
  wire f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa121_y4;
  wire f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa120_y4;
  wire f_u_dadda_pg_rca16_fa122_y0;
  wire f_u_dadda_pg_rca16_fa122_y1;
  wire f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa119_y4;
  wire f_u_dadda_pg_rca16_fa122_y2;
  wire f_u_dadda_pg_rca16_fa122_y3;
  wire f_u_dadda_pg_rca16_fa122_y4;
  wire f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa118_y4;
  wire f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa117_y4;
  wire f_u_dadda_pg_rca16_fa123_y0;
  wire f_u_dadda_pg_rca16_fa123_y1;
  wire f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa116_y4;
  wire f_u_dadda_pg_rca16_fa123_y2;
  wire f_u_dadda_pg_rca16_fa123_y3;
  wire f_u_dadda_pg_rca16_fa123_y4;
  wire f_u_dadda_pg_rca16_and_15_7_a_15;
  wire f_u_dadda_pg_rca16_and_15_7_b_7;
  wire f_u_dadda_pg_rca16_and_15_7_y0;
  wire f_u_dadda_pg_rca16_and_14_8_a_14;
  wire f_u_dadda_pg_rca16_and_14_8_b_8;
  wire f_u_dadda_pg_rca16_and_14_8_y0;
  wire f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_fa115_y4;
  wire f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_and_15_7_y0;
  wire f_u_dadda_pg_rca16_fa124_y0;
  wire f_u_dadda_pg_rca16_fa124_y1;
  wire f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_and_14_8_y0;
  wire f_u_dadda_pg_rca16_fa124_y2;
  wire f_u_dadda_pg_rca16_fa124_y3;
  wire f_u_dadda_pg_rca16_fa124_y4;
  wire f_u_dadda_pg_rca16_and_13_9_a_13;
  wire f_u_dadda_pg_rca16_and_13_9_b_9;
  wire f_u_dadda_pg_rca16_and_13_9_y0;
  wire f_u_dadda_pg_rca16_and_12_10_a_12;
  wire f_u_dadda_pg_rca16_and_12_10_b_10;
  wire f_u_dadda_pg_rca16_and_12_10_y0;
  wire f_u_dadda_pg_rca16_and_11_11_a_11;
  wire f_u_dadda_pg_rca16_and_11_11_b_11;
  wire f_u_dadda_pg_rca16_and_11_11_y0;
  wire f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_13_9_y0;
  wire f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_12_10_y0;
  wire f_u_dadda_pg_rca16_fa125_y0;
  wire f_u_dadda_pg_rca16_fa125_y1;
  wire f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_11_11_y0;
  wire f_u_dadda_pg_rca16_fa125_y2;
  wire f_u_dadda_pg_rca16_fa125_y3;
  wire f_u_dadda_pg_rca16_fa125_y4;
  wire f_u_dadda_pg_rca16_and_10_12_a_10;
  wire f_u_dadda_pg_rca16_and_10_12_b_12;
  wire f_u_dadda_pg_rca16_and_10_12_y0;
  wire f_u_dadda_pg_rca16_and_9_13_a_9;
  wire f_u_dadda_pg_rca16_and_9_13_b_13;
  wire f_u_dadda_pg_rca16_and_9_13_y0;
  wire f_u_dadda_pg_rca16_and_8_14_a_8;
  wire f_u_dadda_pg_rca16_and_8_14_b_14;
  wire f_u_dadda_pg_rca16_and_8_14_y0;
  wire f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_10_12_y0;
  wire f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_9_13_y0;
  wire f_u_dadda_pg_rca16_fa126_y0;
  wire f_u_dadda_pg_rca16_fa126_y1;
  wire f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_8_14_y0;
  wire f_u_dadda_pg_rca16_fa126_y2;
  wire f_u_dadda_pg_rca16_fa126_y3;
  wire f_u_dadda_pg_rca16_fa126_y4;
  wire f_u_dadda_pg_rca16_and_7_15_a_7;
  wire f_u_dadda_pg_rca16_and_7_15_b_15;
  wire f_u_dadda_pg_rca16_and_7_15_y0;
  wire f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_and_7_15_y0;
  wire f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_fa122_y2;
  wire f_u_dadda_pg_rca16_fa127_y0;
  wire f_u_dadda_pg_rca16_fa127_y1;
  wire f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_fa123_y2;
  wire f_u_dadda_pg_rca16_fa127_y2;
  wire f_u_dadda_pg_rca16_fa127_y3;
  wire f_u_dadda_pg_rca16_fa127_y4;
  wire f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa127_y4;
  wire f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa126_y4;
  wire f_u_dadda_pg_rca16_fa128_y0;
  wire f_u_dadda_pg_rca16_fa128_y1;
  wire f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa125_y4;
  wire f_u_dadda_pg_rca16_fa128_y2;
  wire f_u_dadda_pg_rca16_fa128_y3;
  wire f_u_dadda_pg_rca16_fa128_y4;
  wire f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa124_y4;
  wire f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa123_y4;
  wire f_u_dadda_pg_rca16_fa129_y0;
  wire f_u_dadda_pg_rca16_fa129_y1;
  wire f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa122_y4;
  wire f_u_dadda_pg_rca16_fa129_y2;
  wire f_u_dadda_pg_rca16_fa129_y3;
  wire f_u_dadda_pg_rca16_fa129_y4;
  wire f_u_dadda_pg_rca16_and_15_8_a_15;
  wire f_u_dadda_pg_rca16_and_15_8_b_8;
  wire f_u_dadda_pg_rca16_and_15_8_y0;
  wire f_u_dadda_pg_rca16_and_14_9_a_14;
  wire f_u_dadda_pg_rca16_and_14_9_b_9;
  wire f_u_dadda_pg_rca16_and_14_9_y0;
  wire f_u_dadda_pg_rca16_and_13_10_a_13;
  wire f_u_dadda_pg_rca16_and_13_10_b_10;
  wire f_u_dadda_pg_rca16_and_13_10_y0;
  wire f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_15_8_y0;
  wire f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_14_9_y0;
  wire f_u_dadda_pg_rca16_fa130_y0;
  wire f_u_dadda_pg_rca16_fa130_y1;
  wire f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_13_10_y0;
  wire f_u_dadda_pg_rca16_fa130_y2;
  wire f_u_dadda_pg_rca16_fa130_y3;
  wire f_u_dadda_pg_rca16_fa130_y4;
  wire f_u_dadda_pg_rca16_and_12_11_a_12;
  wire f_u_dadda_pg_rca16_and_12_11_b_11;
  wire f_u_dadda_pg_rca16_and_12_11_y0;
  wire f_u_dadda_pg_rca16_and_11_12_a_11;
  wire f_u_dadda_pg_rca16_and_11_12_b_12;
  wire f_u_dadda_pg_rca16_and_11_12_y0;
  wire f_u_dadda_pg_rca16_and_10_13_a_10;
  wire f_u_dadda_pg_rca16_and_10_13_b_13;
  wire f_u_dadda_pg_rca16_and_10_13_y0;
  wire f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_12_11_y0;
  wire f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_11_12_y0;
  wire f_u_dadda_pg_rca16_fa131_y0;
  wire f_u_dadda_pg_rca16_fa131_y1;
  wire f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_10_13_y0;
  wire f_u_dadda_pg_rca16_fa131_y2;
  wire f_u_dadda_pg_rca16_fa131_y3;
  wire f_u_dadda_pg_rca16_fa131_y4;
  wire f_u_dadda_pg_rca16_and_9_14_a_9;
  wire f_u_dadda_pg_rca16_and_9_14_b_14;
  wire f_u_dadda_pg_rca16_and_9_14_y0;
  wire f_u_dadda_pg_rca16_and_8_15_a_8;
  wire f_u_dadda_pg_rca16_and_8_15_b_15;
  wire f_u_dadda_pg_rca16_and_8_15_y0;
  wire f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_and_9_14_y0;
  wire f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_and_8_15_y0;
  wire f_u_dadda_pg_rca16_fa132_y0;
  wire f_u_dadda_pg_rca16_fa132_y1;
  wire f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_fa128_y2;
  wire f_u_dadda_pg_rca16_fa132_y2;
  wire f_u_dadda_pg_rca16_fa132_y3;
  wire f_u_dadda_pg_rca16_fa132_y4;
  wire f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa132_y4;
  wire f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa131_y4;
  wire f_u_dadda_pg_rca16_fa133_y0;
  wire f_u_dadda_pg_rca16_fa133_y1;
  wire f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa130_y4;
  wire f_u_dadda_pg_rca16_fa133_y2;
  wire f_u_dadda_pg_rca16_fa133_y3;
  wire f_u_dadda_pg_rca16_fa133_y4;
  wire f_u_dadda_pg_rca16_and_15_9_a_15;
  wire f_u_dadda_pg_rca16_and_15_9_b_9;
  wire f_u_dadda_pg_rca16_and_15_9_y0;
  wire f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_fa129_y4;
  wire f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_fa128_y4;
  wire f_u_dadda_pg_rca16_fa134_y0;
  wire f_u_dadda_pg_rca16_fa134_y1;
  wire f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_and_15_9_y0;
  wire f_u_dadda_pg_rca16_fa134_y2;
  wire f_u_dadda_pg_rca16_fa134_y3;
  wire f_u_dadda_pg_rca16_fa134_y4;
  wire f_u_dadda_pg_rca16_and_14_10_a_14;
  wire f_u_dadda_pg_rca16_and_14_10_b_10;
  wire f_u_dadda_pg_rca16_and_14_10_y0;
  wire f_u_dadda_pg_rca16_and_13_11_a_13;
  wire f_u_dadda_pg_rca16_and_13_11_b_11;
  wire f_u_dadda_pg_rca16_and_13_11_y0;
  wire f_u_dadda_pg_rca16_and_12_12_a_12;
  wire f_u_dadda_pg_rca16_and_12_12_b_12;
  wire f_u_dadda_pg_rca16_and_12_12_y0;
  wire f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_14_10_y0;
  wire f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_13_11_y0;
  wire f_u_dadda_pg_rca16_fa135_y0;
  wire f_u_dadda_pg_rca16_fa135_y1;
  wire f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_12_12_y0;
  wire f_u_dadda_pg_rca16_fa135_y2;
  wire f_u_dadda_pg_rca16_fa135_y3;
  wire f_u_dadda_pg_rca16_fa135_y4;
  wire f_u_dadda_pg_rca16_and_11_13_a_11;
  wire f_u_dadda_pg_rca16_and_11_13_b_13;
  wire f_u_dadda_pg_rca16_and_11_13_y0;
  wire f_u_dadda_pg_rca16_and_10_14_a_10;
  wire f_u_dadda_pg_rca16_and_10_14_b_14;
  wire f_u_dadda_pg_rca16_and_10_14_y0;
  wire f_u_dadda_pg_rca16_and_9_15_a_9;
  wire f_u_dadda_pg_rca16_and_9_15_b_15;
  wire f_u_dadda_pg_rca16_and_9_15_y0;
  wire f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_11_13_y0;
  wire f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_10_14_y0;
  wire f_u_dadda_pg_rca16_fa136_y0;
  wire f_u_dadda_pg_rca16_fa136_y1;
  wire f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_9_15_y0;
  wire f_u_dadda_pg_rca16_fa136_y2;
  wire f_u_dadda_pg_rca16_fa136_y3;
  wire f_u_dadda_pg_rca16_fa136_y4;
  wire f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa136_y4;
  wire f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa135_y4;
  wire f_u_dadda_pg_rca16_fa137_y0;
  wire f_u_dadda_pg_rca16_fa137_y1;
  wire f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa134_y4;
  wire f_u_dadda_pg_rca16_fa137_y2;
  wire f_u_dadda_pg_rca16_fa137_y3;
  wire f_u_dadda_pg_rca16_fa137_y4;
  wire f_u_dadda_pg_rca16_and_15_10_a_15;
  wire f_u_dadda_pg_rca16_and_15_10_b_10;
  wire f_u_dadda_pg_rca16_and_15_10_y0;
  wire f_u_dadda_pg_rca16_and_14_11_a_14;
  wire f_u_dadda_pg_rca16_and_14_11_b_11;
  wire f_u_dadda_pg_rca16_and_14_11_y0;
  wire f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_fa133_y4;
  wire f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_and_15_10_y0;
  wire f_u_dadda_pg_rca16_fa138_y0;
  wire f_u_dadda_pg_rca16_fa138_y1;
  wire f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_and_14_11_y0;
  wire f_u_dadda_pg_rca16_fa138_y2;
  wire f_u_dadda_pg_rca16_fa138_y3;
  wire f_u_dadda_pg_rca16_fa138_y4;
  wire f_u_dadda_pg_rca16_and_13_12_a_13;
  wire f_u_dadda_pg_rca16_and_13_12_b_12;
  wire f_u_dadda_pg_rca16_and_13_12_y0;
  wire f_u_dadda_pg_rca16_and_12_13_a_12;
  wire f_u_dadda_pg_rca16_and_12_13_b_13;
  wire f_u_dadda_pg_rca16_and_12_13_y0;
  wire f_u_dadda_pg_rca16_and_11_14_a_11;
  wire f_u_dadda_pg_rca16_and_11_14_b_14;
  wire f_u_dadda_pg_rca16_and_11_14_y0;
  wire f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_13_12_y0;
  wire f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_12_13_y0;
  wire f_u_dadda_pg_rca16_fa139_y0;
  wire f_u_dadda_pg_rca16_fa139_y1;
  wire f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_11_14_y0;
  wire f_u_dadda_pg_rca16_fa139_y2;
  wire f_u_dadda_pg_rca16_fa139_y3;
  wire f_u_dadda_pg_rca16_fa139_y4;
  wire f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa139_y4;
  wire f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa138_y4;
  wire f_u_dadda_pg_rca16_fa140_y0;
  wire f_u_dadda_pg_rca16_fa140_y1;
  wire f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa137_y4;
  wire f_u_dadda_pg_rca16_fa140_y2;
  wire f_u_dadda_pg_rca16_fa140_y3;
  wire f_u_dadda_pg_rca16_fa140_y4;
  wire f_u_dadda_pg_rca16_and_15_11_a_15;
  wire f_u_dadda_pg_rca16_and_15_11_b_11;
  wire f_u_dadda_pg_rca16_and_15_11_y0;
  wire f_u_dadda_pg_rca16_and_14_12_a_14;
  wire f_u_dadda_pg_rca16_and_14_12_b_12;
  wire f_u_dadda_pg_rca16_and_14_12_y0;
  wire f_u_dadda_pg_rca16_and_13_13_a_13;
  wire f_u_dadda_pg_rca16_and_13_13_b_13;
  wire f_u_dadda_pg_rca16_and_13_13_y0;
  wire f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_15_11_y0;
  wire f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_14_12_y0;
  wire f_u_dadda_pg_rca16_fa141_y0;
  wire f_u_dadda_pg_rca16_fa141_y1;
  wire f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_13_13_y0;
  wire f_u_dadda_pg_rca16_fa141_y2;
  wire f_u_dadda_pg_rca16_fa141_y3;
  wire f_u_dadda_pg_rca16_fa141_y4;
  wire f_u_dadda_pg_rca16_and_15_12_a_15;
  wire f_u_dadda_pg_rca16_and_15_12_b_12;
  wire f_u_dadda_pg_rca16_and_15_12_y0;
  wire f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_fa141_y4;
  wire f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_fa140_y4;
  wire f_u_dadda_pg_rca16_fa142_y0;
  wire f_u_dadda_pg_rca16_fa142_y1;
  wire f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_and_15_12_y0;
  wire f_u_dadda_pg_rca16_fa142_y2;
  wire f_u_dadda_pg_rca16_fa142_y3;
  wire f_u_dadda_pg_rca16_fa142_y4;
  wire f_u_dadda_pg_rca16_and_3_0_a_3;
  wire f_u_dadda_pg_rca16_and_3_0_b_0;
  wire f_u_dadda_pg_rca16_and_3_0_y0;
  wire f_u_dadda_pg_rca16_and_2_1_a_2;
  wire f_u_dadda_pg_rca16_and_2_1_b_1;
  wire f_u_dadda_pg_rca16_and_2_1_y0;
  wire f_u_dadda_pg_rca16_ha13_f_u_dadda_pg_rca16_and_3_0_y0;
  wire f_u_dadda_pg_rca16_ha13_f_u_dadda_pg_rca16_and_2_1_y0;
  wire f_u_dadda_pg_rca16_ha13_y0;
  wire f_u_dadda_pg_rca16_ha13_y1;
  wire f_u_dadda_pg_rca16_and_2_2_a_2;
  wire f_u_dadda_pg_rca16_and_2_2_b_2;
  wire f_u_dadda_pg_rca16_and_2_2_y0;
  wire f_u_dadda_pg_rca16_and_1_3_a_1;
  wire f_u_dadda_pg_rca16_and_1_3_b_3;
  wire f_u_dadda_pg_rca16_and_1_3_y0;
  wire f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_ha13_y1;
  wire f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_and_2_2_y0;
  wire f_u_dadda_pg_rca16_fa143_y0;
  wire f_u_dadda_pg_rca16_fa143_y1;
  wire f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_and_1_3_y0;
  wire f_u_dadda_pg_rca16_fa143_y2;
  wire f_u_dadda_pg_rca16_fa143_y3;
  wire f_u_dadda_pg_rca16_fa143_y4;
  wire f_u_dadda_pg_rca16_and_1_4_a_1;
  wire f_u_dadda_pg_rca16_and_1_4_b_4;
  wire f_u_dadda_pg_rca16_and_1_4_y0;
  wire f_u_dadda_pg_rca16_and_0_5_a_0;
  wire f_u_dadda_pg_rca16_and_0_5_b_5;
  wire f_u_dadda_pg_rca16_and_0_5_y0;
  wire f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_fa143_y4;
  wire f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_and_1_4_y0;
  wire f_u_dadda_pg_rca16_fa144_y0;
  wire f_u_dadda_pg_rca16_fa144_y1;
  wire f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_and_0_5_y0;
  wire f_u_dadda_pg_rca16_fa144_y2;
  wire f_u_dadda_pg_rca16_fa144_y3;
  wire f_u_dadda_pg_rca16_fa144_y4;
  wire f_u_dadda_pg_rca16_and_0_6_a_0;
  wire f_u_dadda_pg_rca16_and_0_6_b_6;
  wire f_u_dadda_pg_rca16_and_0_6_y0;
  wire f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_fa144_y4;
  wire f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_and_0_6_y0;
  wire f_u_dadda_pg_rca16_fa145_y0;
  wire f_u_dadda_pg_rca16_fa145_y1;
  wire f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_fa9_y2;
  wire f_u_dadda_pg_rca16_fa145_y2;
  wire f_u_dadda_pg_rca16_fa145_y3;
  wire f_u_dadda_pg_rca16_fa145_y4;
  wire f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa145_y4;
  wire f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa11_y2;
  wire f_u_dadda_pg_rca16_fa146_y0;
  wire f_u_dadda_pg_rca16_fa146_y1;
  wire f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa12_y2;
  wire f_u_dadda_pg_rca16_fa146_y2;
  wire f_u_dadda_pg_rca16_fa146_y3;
  wire f_u_dadda_pg_rca16_fa146_y4;
  wire f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa146_y4;
  wire f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa15_y2;
  wire f_u_dadda_pg_rca16_fa147_y0;
  wire f_u_dadda_pg_rca16_fa147_y1;
  wire f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa16_y2;
  wire f_u_dadda_pg_rca16_fa147_y2;
  wire f_u_dadda_pg_rca16_fa147_y3;
  wire f_u_dadda_pg_rca16_fa147_y4;
  wire f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa147_y4;
  wire f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa20_y2;
  wire f_u_dadda_pg_rca16_fa148_y0;
  wire f_u_dadda_pg_rca16_fa148_y1;
  wire f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa21_y2;
  wire f_u_dadda_pg_rca16_fa148_y2;
  wire f_u_dadda_pg_rca16_fa148_y3;
  wire f_u_dadda_pg_rca16_fa148_y4;
  wire f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa148_y4;
  wire f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa26_y2;
  wire f_u_dadda_pg_rca16_fa149_y0;
  wire f_u_dadda_pg_rca16_fa149_y1;
  wire f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa27_y2;
  wire f_u_dadda_pg_rca16_fa149_y2;
  wire f_u_dadda_pg_rca16_fa149_y3;
  wire f_u_dadda_pg_rca16_fa149_y4;
  wire f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa149_y4;
  wire f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa33_y2;
  wire f_u_dadda_pg_rca16_fa150_y0;
  wire f_u_dadda_pg_rca16_fa150_y1;
  wire f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa34_y2;
  wire f_u_dadda_pg_rca16_fa150_y2;
  wire f_u_dadda_pg_rca16_fa150_y3;
  wire f_u_dadda_pg_rca16_fa150_y4;
  wire f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa150_y4;
  wire f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa41_y2;
  wire f_u_dadda_pg_rca16_fa151_y0;
  wire f_u_dadda_pg_rca16_fa151_y1;
  wire f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa42_y2;
  wire f_u_dadda_pg_rca16_fa151_y2;
  wire f_u_dadda_pg_rca16_fa151_y3;
  wire f_u_dadda_pg_rca16_fa151_y4;
  wire f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa151_y4;
  wire f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa49_y2;
  wire f_u_dadda_pg_rca16_fa152_y0;
  wire f_u_dadda_pg_rca16_fa152_y1;
  wire f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa50_y2;
  wire f_u_dadda_pg_rca16_fa152_y2;
  wire f_u_dadda_pg_rca16_fa152_y3;
  wire f_u_dadda_pg_rca16_fa152_y4;
  wire f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa152_y4;
  wire f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa58_y2;
  wire f_u_dadda_pg_rca16_fa153_y0;
  wire f_u_dadda_pg_rca16_fa153_y1;
  wire f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa59_y2;
  wire f_u_dadda_pg_rca16_fa153_y2;
  wire f_u_dadda_pg_rca16_fa153_y3;
  wire f_u_dadda_pg_rca16_fa153_y4;
  wire f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa153_y4;
  wire f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa67_y2;
  wire f_u_dadda_pg_rca16_fa154_y0;
  wire f_u_dadda_pg_rca16_fa154_y1;
  wire f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa68_y2;
  wire f_u_dadda_pg_rca16_fa154_y2;
  wire f_u_dadda_pg_rca16_fa154_y3;
  wire f_u_dadda_pg_rca16_fa154_y4;
  wire f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa154_y4;
  wire f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa76_y2;
  wire f_u_dadda_pg_rca16_fa155_y0;
  wire f_u_dadda_pg_rca16_fa155_y1;
  wire f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa77_y2;
  wire f_u_dadda_pg_rca16_fa155_y2;
  wire f_u_dadda_pg_rca16_fa155_y3;
  wire f_u_dadda_pg_rca16_fa155_y4;
  wire f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa155_y4;
  wire f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa85_y2;
  wire f_u_dadda_pg_rca16_fa156_y0;
  wire f_u_dadda_pg_rca16_fa156_y1;
  wire f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa86_y2;
  wire f_u_dadda_pg_rca16_fa156_y2;
  wire f_u_dadda_pg_rca16_fa156_y3;
  wire f_u_dadda_pg_rca16_fa156_y4;
  wire f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa156_y4;
  wire f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa94_y2;
  wire f_u_dadda_pg_rca16_fa157_y0;
  wire f_u_dadda_pg_rca16_fa157_y1;
  wire f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa95_y2;
  wire f_u_dadda_pg_rca16_fa157_y2;
  wire f_u_dadda_pg_rca16_fa157_y3;
  wire f_u_dadda_pg_rca16_fa157_y4;
  wire f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa157_y4;
  wire f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa103_y2;
  wire f_u_dadda_pg_rca16_fa158_y0;
  wire f_u_dadda_pg_rca16_fa158_y1;
  wire f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa104_y2;
  wire f_u_dadda_pg_rca16_fa158_y2;
  wire f_u_dadda_pg_rca16_fa158_y3;
  wire f_u_dadda_pg_rca16_fa158_y4;
  wire f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa158_y4;
  wire f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa111_y2;
  wire f_u_dadda_pg_rca16_fa159_y0;
  wire f_u_dadda_pg_rca16_fa159_y1;
  wire f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa112_y2;
  wire f_u_dadda_pg_rca16_fa159_y2;
  wire f_u_dadda_pg_rca16_fa159_y3;
  wire f_u_dadda_pg_rca16_fa159_y4;
  wire f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa159_y4;
  wire f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa118_y2;
  wire f_u_dadda_pg_rca16_fa160_y0;
  wire f_u_dadda_pg_rca16_fa160_y1;
  wire f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa119_y2;
  wire f_u_dadda_pg_rca16_fa160_y2;
  wire f_u_dadda_pg_rca16_fa160_y3;
  wire f_u_dadda_pg_rca16_fa160_y4;
  wire f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa160_y4;
  wire f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa124_y2;
  wire f_u_dadda_pg_rca16_fa161_y0;
  wire f_u_dadda_pg_rca16_fa161_y1;
  wire f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa125_y2;
  wire f_u_dadda_pg_rca16_fa161_y2;
  wire f_u_dadda_pg_rca16_fa161_y3;
  wire f_u_dadda_pg_rca16_fa161_y4;
  wire f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa161_y4;
  wire f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa129_y2;
  wire f_u_dadda_pg_rca16_fa162_y0;
  wire f_u_dadda_pg_rca16_fa162_y1;
  wire f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa130_y2;
  wire f_u_dadda_pg_rca16_fa162_y2;
  wire f_u_dadda_pg_rca16_fa162_y3;
  wire f_u_dadda_pg_rca16_fa162_y4;
  wire f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa162_y4;
  wire f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa133_y2;
  wire f_u_dadda_pg_rca16_fa163_y0;
  wire f_u_dadda_pg_rca16_fa163_y1;
  wire f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa134_y2;
  wire f_u_dadda_pg_rca16_fa163_y2;
  wire f_u_dadda_pg_rca16_fa163_y3;
  wire f_u_dadda_pg_rca16_fa163_y4;
  wire f_u_dadda_pg_rca16_and_10_15_a_10;
  wire f_u_dadda_pg_rca16_and_10_15_b_15;
  wire f_u_dadda_pg_rca16_and_10_15_y0;
  wire f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_fa163_y4;
  wire f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_and_10_15_y0;
  wire f_u_dadda_pg_rca16_fa164_y0;
  wire f_u_dadda_pg_rca16_fa164_y1;
  wire f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_fa137_y2;
  wire f_u_dadda_pg_rca16_fa164_y2;
  wire f_u_dadda_pg_rca16_fa164_y3;
  wire f_u_dadda_pg_rca16_fa164_y4;
  wire f_u_dadda_pg_rca16_and_12_14_a_12;
  wire f_u_dadda_pg_rca16_and_12_14_b_14;
  wire f_u_dadda_pg_rca16_and_12_14_y0;
  wire f_u_dadda_pg_rca16_and_11_15_a_11;
  wire f_u_dadda_pg_rca16_and_11_15_b_15;
  wire f_u_dadda_pg_rca16_and_11_15_y0;
  wire f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_fa164_y4;
  wire f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_and_12_14_y0;
  wire f_u_dadda_pg_rca16_fa165_y0;
  wire f_u_dadda_pg_rca16_fa165_y1;
  wire f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_and_11_15_y0;
  wire f_u_dadda_pg_rca16_fa165_y2;
  wire f_u_dadda_pg_rca16_fa165_y3;
  wire f_u_dadda_pg_rca16_fa165_y4;
  wire f_u_dadda_pg_rca16_and_14_13_a_14;
  wire f_u_dadda_pg_rca16_and_14_13_b_13;
  wire f_u_dadda_pg_rca16_and_14_13_y0;
  wire f_u_dadda_pg_rca16_and_13_14_a_13;
  wire f_u_dadda_pg_rca16_and_13_14_b_14;
  wire f_u_dadda_pg_rca16_and_13_14_y0;
  wire f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_fa165_y4;
  wire f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_and_14_13_y0;
  wire f_u_dadda_pg_rca16_fa166_y0;
  wire f_u_dadda_pg_rca16_fa166_y1;
  wire f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_and_13_14_y0;
  wire f_u_dadda_pg_rca16_fa166_y2;
  wire f_u_dadda_pg_rca16_fa166_y3;
  wire f_u_dadda_pg_rca16_fa166_y4;
  wire f_u_dadda_pg_rca16_and_15_13_a_15;
  wire f_u_dadda_pg_rca16_and_15_13_b_13;
  wire f_u_dadda_pg_rca16_and_15_13_y0;
  wire f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_fa166_y4;
  wire f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_fa142_y4;
  wire f_u_dadda_pg_rca16_fa167_y0;
  wire f_u_dadda_pg_rca16_fa167_y1;
  wire f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_and_15_13_y0;
  wire f_u_dadda_pg_rca16_fa167_y2;
  wire f_u_dadda_pg_rca16_fa167_y3;
  wire f_u_dadda_pg_rca16_fa167_y4;
  wire f_u_dadda_pg_rca16_and_2_0_a_2;
  wire f_u_dadda_pg_rca16_and_2_0_b_0;
  wire f_u_dadda_pg_rca16_and_2_0_y0;
  wire f_u_dadda_pg_rca16_and_1_1_a_1;
  wire f_u_dadda_pg_rca16_and_1_1_b_1;
  wire f_u_dadda_pg_rca16_and_1_1_y0;
  wire f_u_dadda_pg_rca16_ha14_f_u_dadda_pg_rca16_and_2_0_y0;
  wire f_u_dadda_pg_rca16_ha14_f_u_dadda_pg_rca16_and_1_1_y0;
  wire f_u_dadda_pg_rca16_ha14_y0;
  wire f_u_dadda_pg_rca16_ha14_y1;
  wire f_u_dadda_pg_rca16_and_1_2_a_1;
  wire f_u_dadda_pg_rca16_and_1_2_b_2;
  wire f_u_dadda_pg_rca16_and_1_2_y0;
  wire f_u_dadda_pg_rca16_and_0_3_a_0;
  wire f_u_dadda_pg_rca16_and_0_3_b_3;
  wire f_u_dadda_pg_rca16_and_0_3_y0;
  wire f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_ha14_y1;
  wire f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_and_1_2_y0;
  wire f_u_dadda_pg_rca16_fa168_y0;
  wire f_u_dadda_pg_rca16_fa168_y1;
  wire f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_and_0_3_y0;
  wire f_u_dadda_pg_rca16_fa168_y2;
  wire f_u_dadda_pg_rca16_fa168_y3;
  wire f_u_dadda_pg_rca16_fa168_y4;
  wire f_u_dadda_pg_rca16_and_0_4_a_0;
  wire f_u_dadda_pg_rca16_and_0_4_b_4;
  wire f_u_dadda_pg_rca16_and_0_4_y0;
  wire f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_fa168_y4;
  wire f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_and_0_4_y0;
  wire f_u_dadda_pg_rca16_fa169_y0;
  wire f_u_dadda_pg_rca16_fa169_y1;
  wire f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_ha4_y0;
  wire f_u_dadda_pg_rca16_fa169_y2;
  wire f_u_dadda_pg_rca16_fa169_y3;
  wire f_u_dadda_pg_rca16_fa169_y4;
  wire f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_fa169_y4;
  wire f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_fa8_y2;
  wire f_u_dadda_pg_rca16_fa170_y0;
  wire f_u_dadda_pg_rca16_fa170_y1;
  wire f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_ha5_y0;
  wire f_u_dadda_pg_rca16_fa170_y2;
  wire f_u_dadda_pg_rca16_fa170_y3;
  wire f_u_dadda_pg_rca16_fa170_y4;
  wire f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_fa170_y4;
  wire f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_fa10_y2;
  wire f_u_dadda_pg_rca16_fa171_y0;
  wire f_u_dadda_pg_rca16_fa171_y1;
  wire f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_ha6_y0;
  wire f_u_dadda_pg_rca16_fa171_y2;
  wire f_u_dadda_pg_rca16_fa171_y3;
  wire f_u_dadda_pg_rca16_fa171_y4;
  wire f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_fa171_y4;
  wire f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_fa13_y2;
  wire f_u_dadda_pg_rca16_fa172_y0;
  wire f_u_dadda_pg_rca16_fa172_y1;
  wire f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_ha7_y0;
  wire f_u_dadda_pg_rca16_fa172_y2;
  wire f_u_dadda_pg_rca16_fa172_y3;
  wire f_u_dadda_pg_rca16_fa172_y4;
  wire f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_fa172_y4;
  wire f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_fa17_y2;
  wire f_u_dadda_pg_rca16_fa173_y0;
  wire f_u_dadda_pg_rca16_fa173_y1;
  wire f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_ha8_y0;
  wire f_u_dadda_pg_rca16_fa173_y2;
  wire f_u_dadda_pg_rca16_fa173_y3;
  wire f_u_dadda_pg_rca16_fa173_y4;
  wire f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_fa173_y4;
  wire f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_fa22_y2;
  wire f_u_dadda_pg_rca16_fa174_y0;
  wire f_u_dadda_pg_rca16_fa174_y1;
  wire f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_ha9_y0;
  wire f_u_dadda_pg_rca16_fa174_y2;
  wire f_u_dadda_pg_rca16_fa174_y3;
  wire f_u_dadda_pg_rca16_fa174_y4;
  wire f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_fa174_y4;
  wire f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_fa28_y2;
  wire f_u_dadda_pg_rca16_fa175_y0;
  wire f_u_dadda_pg_rca16_fa175_y1;
  wire f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_ha10_y0;
  wire f_u_dadda_pg_rca16_fa175_y2;
  wire f_u_dadda_pg_rca16_fa175_y3;
  wire f_u_dadda_pg_rca16_fa175_y4;
  wire f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_fa175_y4;
  wire f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_fa35_y2;
  wire f_u_dadda_pg_rca16_fa176_y0;
  wire f_u_dadda_pg_rca16_fa176_y1;
  wire f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_ha11_y0;
  wire f_u_dadda_pg_rca16_fa176_y2;
  wire f_u_dadda_pg_rca16_fa176_y3;
  wire f_u_dadda_pg_rca16_fa176_y4;
  wire f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_fa176_y4;
  wire f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_fa43_y2;
  wire f_u_dadda_pg_rca16_fa177_y0;
  wire f_u_dadda_pg_rca16_fa177_y1;
  wire f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_ha12_y0;
  wire f_u_dadda_pg_rca16_fa177_y2;
  wire f_u_dadda_pg_rca16_fa177_y3;
  wire f_u_dadda_pg_rca16_fa177_y4;
  wire f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa177_y4;
  wire f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa51_y2;
  wire f_u_dadda_pg_rca16_fa178_y0;
  wire f_u_dadda_pg_rca16_fa178_y1;
  wire f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa52_y2;
  wire f_u_dadda_pg_rca16_fa178_y2;
  wire f_u_dadda_pg_rca16_fa178_y3;
  wire f_u_dadda_pg_rca16_fa178_y4;
  wire f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa178_y4;
  wire f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa60_y2;
  wire f_u_dadda_pg_rca16_fa179_y0;
  wire f_u_dadda_pg_rca16_fa179_y1;
  wire f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa61_y2;
  wire f_u_dadda_pg_rca16_fa179_y2;
  wire f_u_dadda_pg_rca16_fa179_y3;
  wire f_u_dadda_pg_rca16_fa179_y4;
  wire f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa179_y4;
  wire f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa69_y2;
  wire f_u_dadda_pg_rca16_fa180_y0;
  wire f_u_dadda_pg_rca16_fa180_y1;
  wire f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa70_y2;
  wire f_u_dadda_pg_rca16_fa180_y2;
  wire f_u_dadda_pg_rca16_fa180_y3;
  wire f_u_dadda_pg_rca16_fa180_y4;
  wire f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa180_y4;
  wire f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa78_y2;
  wire f_u_dadda_pg_rca16_fa181_y0;
  wire f_u_dadda_pg_rca16_fa181_y1;
  wire f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa79_y2;
  wire f_u_dadda_pg_rca16_fa181_y2;
  wire f_u_dadda_pg_rca16_fa181_y3;
  wire f_u_dadda_pg_rca16_fa181_y4;
  wire f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa181_y4;
  wire f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa87_y2;
  wire f_u_dadda_pg_rca16_fa182_y0;
  wire f_u_dadda_pg_rca16_fa182_y1;
  wire f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa88_y2;
  wire f_u_dadda_pg_rca16_fa182_y2;
  wire f_u_dadda_pg_rca16_fa182_y3;
  wire f_u_dadda_pg_rca16_fa182_y4;
  wire f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa182_y4;
  wire f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa96_y2;
  wire f_u_dadda_pg_rca16_fa183_y0;
  wire f_u_dadda_pg_rca16_fa183_y1;
  wire f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa97_y2;
  wire f_u_dadda_pg_rca16_fa183_y2;
  wire f_u_dadda_pg_rca16_fa183_y3;
  wire f_u_dadda_pg_rca16_fa183_y4;
  wire f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa183_y4;
  wire f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa105_y2;
  wire f_u_dadda_pg_rca16_fa184_y0;
  wire f_u_dadda_pg_rca16_fa184_y1;
  wire f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa106_y2;
  wire f_u_dadda_pg_rca16_fa184_y2;
  wire f_u_dadda_pg_rca16_fa184_y3;
  wire f_u_dadda_pg_rca16_fa184_y4;
  wire f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa184_y4;
  wire f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa113_y2;
  wire f_u_dadda_pg_rca16_fa185_y0;
  wire f_u_dadda_pg_rca16_fa185_y1;
  wire f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa114_y2;
  wire f_u_dadda_pg_rca16_fa185_y2;
  wire f_u_dadda_pg_rca16_fa185_y3;
  wire f_u_dadda_pg_rca16_fa185_y4;
  wire f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa185_y4;
  wire f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa120_y2;
  wire f_u_dadda_pg_rca16_fa186_y0;
  wire f_u_dadda_pg_rca16_fa186_y1;
  wire f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa121_y2;
  wire f_u_dadda_pg_rca16_fa186_y2;
  wire f_u_dadda_pg_rca16_fa186_y3;
  wire f_u_dadda_pg_rca16_fa186_y4;
  wire f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa186_y4;
  wire f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa126_y2;
  wire f_u_dadda_pg_rca16_fa187_y0;
  wire f_u_dadda_pg_rca16_fa187_y1;
  wire f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa127_y2;
  wire f_u_dadda_pg_rca16_fa187_y2;
  wire f_u_dadda_pg_rca16_fa187_y3;
  wire f_u_dadda_pg_rca16_fa187_y4;
  wire f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa187_y4;
  wire f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa131_y2;
  wire f_u_dadda_pg_rca16_fa188_y0;
  wire f_u_dadda_pg_rca16_fa188_y1;
  wire f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa132_y2;
  wire f_u_dadda_pg_rca16_fa188_y2;
  wire f_u_dadda_pg_rca16_fa188_y3;
  wire f_u_dadda_pg_rca16_fa188_y4;
  wire f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa188_y4;
  wire f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa135_y2;
  wire f_u_dadda_pg_rca16_fa189_y0;
  wire f_u_dadda_pg_rca16_fa189_y1;
  wire f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa136_y2;
  wire f_u_dadda_pg_rca16_fa189_y2;
  wire f_u_dadda_pg_rca16_fa189_y3;
  wire f_u_dadda_pg_rca16_fa189_y4;
  wire f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa189_y4;
  wire f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa138_y2;
  wire f_u_dadda_pg_rca16_fa190_y0;
  wire f_u_dadda_pg_rca16_fa190_y1;
  wire f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa139_y2;
  wire f_u_dadda_pg_rca16_fa190_y2;
  wire f_u_dadda_pg_rca16_fa190_y3;
  wire f_u_dadda_pg_rca16_fa190_y4;
  wire f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa190_y4;
  wire f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa140_y2;
  wire f_u_dadda_pg_rca16_fa191_y0;
  wire f_u_dadda_pg_rca16_fa191_y1;
  wire f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa141_y2;
  wire f_u_dadda_pg_rca16_fa191_y2;
  wire f_u_dadda_pg_rca16_fa191_y3;
  wire f_u_dadda_pg_rca16_fa191_y4;
  wire f_u_dadda_pg_rca16_and_12_15_a_12;
  wire f_u_dadda_pg_rca16_and_12_15_b_15;
  wire f_u_dadda_pg_rca16_and_12_15_y0;
  wire f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_fa191_y4;
  wire f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_and_12_15_y0;
  wire f_u_dadda_pg_rca16_fa192_y0;
  wire f_u_dadda_pg_rca16_fa192_y1;
  wire f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_fa142_y2;
  wire f_u_dadda_pg_rca16_fa192_y2;
  wire f_u_dadda_pg_rca16_fa192_y3;
  wire f_u_dadda_pg_rca16_fa192_y4;
  wire f_u_dadda_pg_rca16_and_14_14_a_14;
  wire f_u_dadda_pg_rca16_and_14_14_b_14;
  wire f_u_dadda_pg_rca16_and_14_14_y0;
  wire f_u_dadda_pg_rca16_and_13_15_a_13;
  wire f_u_dadda_pg_rca16_and_13_15_b_15;
  wire f_u_dadda_pg_rca16_and_13_15_y0;
  wire f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_fa192_y4;
  wire f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_and_14_14_y0;
  wire f_u_dadda_pg_rca16_fa193_y0;
  wire f_u_dadda_pg_rca16_fa193_y1;
  wire f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_and_13_15_y0;
  wire f_u_dadda_pg_rca16_fa193_y2;
  wire f_u_dadda_pg_rca16_fa193_y3;
  wire f_u_dadda_pg_rca16_fa193_y4;
  wire f_u_dadda_pg_rca16_and_15_14_a_15;
  wire f_u_dadda_pg_rca16_and_15_14_b_14;
  wire f_u_dadda_pg_rca16_and_15_14_y0;
  wire f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_fa193_y4;
  wire f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_fa167_y4;
  wire f_u_dadda_pg_rca16_fa194_y0;
  wire f_u_dadda_pg_rca16_fa194_y1;
  wire f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_and_15_14_y0;
  wire f_u_dadda_pg_rca16_fa194_y2;
  wire f_u_dadda_pg_rca16_fa194_y3;
  wire f_u_dadda_pg_rca16_fa194_y4;
  wire f_u_dadda_pg_rca16_and_0_0_a_0;
  wire f_u_dadda_pg_rca16_and_0_0_b_0;
  wire f_u_dadda_pg_rca16_and_0_0_y0;
  wire f_u_dadda_pg_rca16_and_1_0_a_1;
  wire f_u_dadda_pg_rca16_and_1_0_b_0;
  wire f_u_dadda_pg_rca16_and_1_0_y0;
  wire f_u_dadda_pg_rca16_and_0_2_a_0;
  wire f_u_dadda_pg_rca16_and_0_2_b_2;
  wire f_u_dadda_pg_rca16_and_0_2_y0;
  wire f_u_dadda_pg_rca16_and_14_15_a_14;
  wire f_u_dadda_pg_rca16_and_14_15_b_15;
  wire f_u_dadda_pg_rca16_and_14_15_y0;
  wire f_u_dadda_pg_rca16_and_0_1_a_0;
  wire f_u_dadda_pg_rca16_and_0_1_b_1;
  wire f_u_dadda_pg_rca16_and_0_1_y0;
  wire f_u_dadda_pg_rca16_and_15_15_a_15;
  wire f_u_dadda_pg_rca16_and_15_15_b_15;
  wire f_u_dadda_pg_rca16_and_15_15_y0;
  wire constant_wire_value_0_f_u_dadda_pg_rca16_and_1_0_y0;
  wire constant_wire_value_0_f_u_dadda_pg_rca16_and_0_1_y0;
  wire constant_wire_value_0_y0;
  wire constant_wire_value_0_y1;
  wire constant_wire_0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa0_f_u_dadda_pg_rca16_and_1_0_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa0_f_u_dadda_pg_rca16_and_0_1_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa0_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa0_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa0_constant_wire_0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa0_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and0_constant_wire_0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and0_f_u_dadda_pg_rca16_u_pg_rca30_fa0_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and0_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or0_f_u_dadda_pg_rca16_u_pg_rca30_and0_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or0_f_u_dadda_pg_rca16_u_pg_rca30_fa0_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or0_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_and_0_2_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_ha14_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa1_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa1_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_u_pg_rca30_or0_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa1_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and1_f_u_dadda_pg_rca16_u_pg_rca30_or0_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and1_f_u_dadda_pg_rca16_u_pg_rca30_fa1_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and1_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or1_f_u_dadda_pg_rca16_u_pg_rca30_and1_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or1_f_u_dadda_pg_rca16_u_pg_rca30_fa1_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or1_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_ha13_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_fa168_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa2_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa2_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_u_pg_rca30_or1_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa2_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and2_f_u_dadda_pg_rca16_u_pg_rca30_or1_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and2_f_u_dadda_pg_rca16_u_pg_rca30_fa2_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and2_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or2_f_u_dadda_pg_rca16_u_pg_rca30_and2_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or2_f_u_dadda_pg_rca16_u_pg_rca30_fa2_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or2_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_fa143_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_fa169_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa3_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa3_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_u_pg_rca30_or2_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa3_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and3_f_u_dadda_pg_rca16_u_pg_rca30_or2_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and3_f_u_dadda_pg_rca16_u_pg_rca30_fa3_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and3_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or3_f_u_dadda_pg_rca16_u_pg_rca30_and3_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or3_f_u_dadda_pg_rca16_u_pg_rca30_fa3_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or3_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_fa144_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_fa170_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa4_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa4_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_u_pg_rca30_or3_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa4_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and4_f_u_dadda_pg_rca16_u_pg_rca30_or3_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and4_f_u_dadda_pg_rca16_u_pg_rca30_fa4_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and4_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or4_f_u_dadda_pg_rca16_u_pg_rca30_and4_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or4_f_u_dadda_pg_rca16_u_pg_rca30_fa4_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or4_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_fa145_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_fa171_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa5_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa5_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_u_pg_rca30_or4_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa5_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and5_f_u_dadda_pg_rca16_u_pg_rca30_or4_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and5_f_u_dadda_pg_rca16_u_pg_rca30_fa5_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and5_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or5_f_u_dadda_pg_rca16_u_pg_rca30_and5_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or5_f_u_dadda_pg_rca16_u_pg_rca30_fa5_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or5_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_fa146_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_fa172_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa6_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa6_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_u_pg_rca30_or5_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa6_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and6_f_u_dadda_pg_rca16_u_pg_rca30_or5_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and6_f_u_dadda_pg_rca16_u_pg_rca30_fa6_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and6_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or6_f_u_dadda_pg_rca16_u_pg_rca30_and6_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or6_f_u_dadda_pg_rca16_u_pg_rca30_fa6_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or6_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_fa147_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_fa173_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa7_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa7_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_u_pg_rca30_or6_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa7_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and7_f_u_dadda_pg_rca16_u_pg_rca30_or6_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and7_f_u_dadda_pg_rca16_u_pg_rca30_fa7_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and7_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or7_f_u_dadda_pg_rca16_u_pg_rca30_and7_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or7_f_u_dadda_pg_rca16_u_pg_rca30_fa7_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or7_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_fa148_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_fa174_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa8_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa8_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_u_pg_rca30_or7_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa8_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and8_f_u_dadda_pg_rca16_u_pg_rca30_or7_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and8_f_u_dadda_pg_rca16_u_pg_rca30_fa8_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and8_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or8_f_u_dadda_pg_rca16_u_pg_rca30_and8_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or8_f_u_dadda_pg_rca16_u_pg_rca30_fa8_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or8_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_fa149_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_fa175_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa9_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa9_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_u_pg_rca30_or8_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa9_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and9_f_u_dadda_pg_rca16_u_pg_rca30_or8_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and9_f_u_dadda_pg_rca16_u_pg_rca30_fa9_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and9_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or9_f_u_dadda_pg_rca16_u_pg_rca30_and9_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or9_f_u_dadda_pg_rca16_u_pg_rca30_fa9_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or9_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_fa150_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_fa176_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa10_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa10_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_u_pg_rca30_or9_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa10_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and10_f_u_dadda_pg_rca16_u_pg_rca30_or9_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and10_f_u_dadda_pg_rca16_u_pg_rca30_fa10_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and10_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or10_f_u_dadda_pg_rca16_u_pg_rca30_and10_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or10_f_u_dadda_pg_rca16_u_pg_rca30_fa10_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or10_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_fa151_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_fa177_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa11_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa11_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_u_pg_rca30_or10_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa11_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and11_f_u_dadda_pg_rca16_u_pg_rca30_or10_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and11_f_u_dadda_pg_rca16_u_pg_rca30_fa11_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and11_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or11_f_u_dadda_pg_rca16_u_pg_rca30_and11_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or11_f_u_dadda_pg_rca16_u_pg_rca30_fa11_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or11_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_fa152_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_fa178_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa12_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa12_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_u_pg_rca30_or11_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa12_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and12_f_u_dadda_pg_rca16_u_pg_rca30_or11_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and12_f_u_dadda_pg_rca16_u_pg_rca30_fa12_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and12_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or12_f_u_dadda_pg_rca16_u_pg_rca30_and12_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or12_f_u_dadda_pg_rca16_u_pg_rca30_fa12_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or12_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_fa153_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_fa179_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa13_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa13_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_u_pg_rca30_or12_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa13_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and13_f_u_dadda_pg_rca16_u_pg_rca30_or12_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and13_f_u_dadda_pg_rca16_u_pg_rca30_fa13_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and13_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or13_f_u_dadda_pg_rca16_u_pg_rca30_and13_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or13_f_u_dadda_pg_rca16_u_pg_rca30_fa13_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or13_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_fa154_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_fa180_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa14_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa14_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_u_pg_rca30_or13_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa14_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and14_f_u_dadda_pg_rca16_u_pg_rca30_or13_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and14_f_u_dadda_pg_rca16_u_pg_rca30_fa14_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and14_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or14_f_u_dadda_pg_rca16_u_pg_rca30_and14_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or14_f_u_dadda_pg_rca16_u_pg_rca30_fa14_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or14_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_fa155_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_fa181_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa15_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_u_pg_rca30_or14_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa15_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and15_f_u_dadda_pg_rca16_u_pg_rca30_or14_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and15_f_u_dadda_pg_rca16_u_pg_rca30_fa15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or15_f_u_dadda_pg_rca16_u_pg_rca30_and15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or15_f_u_dadda_pg_rca16_u_pg_rca30_fa15_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_fa156_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_fa182_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa16_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa16_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_u_pg_rca30_or15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa16_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and16_f_u_dadda_pg_rca16_u_pg_rca30_or15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and16_f_u_dadda_pg_rca16_u_pg_rca30_fa16_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and16_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or16_f_u_dadda_pg_rca16_u_pg_rca30_and16_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or16_f_u_dadda_pg_rca16_u_pg_rca30_fa16_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or16_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_fa157_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_fa183_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa17_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa17_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_u_pg_rca30_or16_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa17_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and17_f_u_dadda_pg_rca16_u_pg_rca30_or16_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and17_f_u_dadda_pg_rca16_u_pg_rca30_fa17_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and17_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or17_f_u_dadda_pg_rca16_u_pg_rca30_and17_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or17_f_u_dadda_pg_rca16_u_pg_rca30_fa17_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or17_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_fa158_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_fa184_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa18_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa18_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_u_pg_rca30_or17_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa18_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and18_f_u_dadda_pg_rca16_u_pg_rca30_or17_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and18_f_u_dadda_pg_rca16_u_pg_rca30_fa18_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and18_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or18_f_u_dadda_pg_rca16_u_pg_rca30_and18_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or18_f_u_dadda_pg_rca16_u_pg_rca30_fa18_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or18_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_fa159_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_fa185_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa19_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa19_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_u_pg_rca30_or18_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa19_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and19_f_u_dadda_pg_rca16_u_pg_rca30_or18_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and19_f_u_dadda_pg_rca16_u_pg_rca30_fa19_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and19_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or19_f_u_dadda_pg_rca16_u_pg_rca30_and19_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or19_f_u_dadda_pg_rca16_u_pg_rca30_fa19_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or19_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_fa160_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_fa186_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa20_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa20_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_u_pg_rca30_or19_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa20_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and20_f_u_dadda_pg_rca16_u_pg_rca30_or19_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and20_f_u_dadda_pg_rca16_u_pg_rca30_fa20_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and20_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or20_f_u_dadda_pg_rca16_u_pg_rca30_and20_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or20_f_u_dadda_pg_rca16_u_pg_rca30_fa20_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or20_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_fa161_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_fa187_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa21_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa21_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_u_pg_rca30_or20_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa21_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and21_f_u_dadda_pg_rca16_u_pg_rca30_or20_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and21_f_u_dadda_pg_rca16_u_pg_rca30_fa21_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and21_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or21_f_u_dadda_pg_rca16_u_pg_rca30_and21_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or21_f_u_dadda_pg_rca16_u_pg_rca30_fa21_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or21_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_fa162_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_fa188_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa22_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa22_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_u_pg_rca30_or21_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa22_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and22_f_u_dadda_pg_rca16_u_pg_rca30_or21_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and22_f_u_dadda_pg_rca16_u_pg_rca30_fa22_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and22_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or22_f_u_dadda_pg_rca16_u_pg_rca30_and22_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or22_f_u_dadda_pg_rca16_u_pg_rca30_fa22_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or22_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_fa163_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_fa189_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa23_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa23_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_u_pg_rca30_or22_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa23_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and23_f_u_dadda_pg_rca16_u_pg_rca30_or22_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and23_f_u_dadda_pg_rca16_u_pg_rca30_fa23_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and23_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or23_f_u_dadda_pg_rca16_u_pg_rca30_and23_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or23_f_u_dadda_pg_rca16_u_pg_rca30_fa23_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or23_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_fa164_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_fa190_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa24_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa24_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_u_pg_rca30_or23_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa24_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and24_f_u_dadda_pg_rca16_u_pg_rca30_or23_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and24_f_u_dadda_pg_rca16_u_pg_rca30_fa24_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and24_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or24_f_u_dadda_pg_rca16_u_pg_rca30_and24_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or24_f_u_dadda_pg_rca16_u_pg_rca30_fa24_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or24_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_fa165_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_fa191_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa25_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa25_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_u_pg_rca30_or24_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa25_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and25_f_u_dadda_pg_rca16_u_pg_rca30_or24_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and25_f_u_dadda_pg_rca16_u_pg_rca30_fa25_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and25_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or25_f_u_dadda_pg_rca16_u_pg_rca30_and25_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or25_f_u_dadda_pg_rca16_u_pg_rca30_fa25_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or25_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_fa166_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_fa192_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa26_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa26_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_u_pg_rca30_or25_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa26_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and26_f_u_dadda_pg_rca16_u_pg_rca30_or25_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and26_f_u_dadda_pg_rca16_u_pg_rca30_fa26_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and26_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or26_f_u_dadda_pg_rca16_u_pg_rca30_and26_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or26_f_u_dadda_pg_rca16_u_pg_rca30_fa26_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or26_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_fa167_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_fa193_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa27_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa27_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_u_pg_rca30_or26_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa27_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and27_f_u_dadda_pg_rca16_u_pg_rca30_or26_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and27_f_u_dadda_pg_rca16_u_pg_rca30_fa27_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and27_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or27_f_u_dadda_pg_rca16_u_pg_rca30_and27_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or27_f_u_dadda_pg_rca16_u_pg_rca30_fa27_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or27_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_and_14_15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_fa194_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa28_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa28_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_u_pg_rca30_or27_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa28_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and28_f_u_dadda_pg_rca16_u_pg_rca30_or27_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and28_f_u_dadda_pg_rca16_u_pg_rca30_fa28_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and28_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or28_f_u_dadda_pg_rca16_u_pg_rca30_and28_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or28_f_u_dadda_pg_rca16_u_pg_rca30_fa28_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or28_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_fa194_y4;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_and_15_15_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa29_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa29_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_u_pg_rca30_or28_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_fa29_y2;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and29_f_u_dadda_pg_rca16_u_pg_rca30_or28_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and29_f_u_dadda_pg_rca16_u_pg_rca30_fa29_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_and29_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or29_f_u_dadda_pg_rca16_u_pg_rca30_and29_y0;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or29_f_u_dadda_pg_rca16_u_pg_rca30_fa29_y1;
  wire f_u_dadda_pg_rca16_u_pg_rca30_or29_y0;

  assign a_0 = a[0];
  assign a_1 = a[1];
  assign a_2 = a[2];
  assign a_3 = a[3];
  assign a_4 = a[4];
  assign a_5 = a[5];
  assign a_6 = a[6];
  assign a_7 = a[7];
  assign a_8 = a[8];
  assign a_9 = a[9];
  assign a_10 = a[10];
  assign a_11 = a[11];
  assign a_12 = a[12];
  assign a_13 = a[13];
  assign a_14 = a[14];
  assign a_15 = a[15];
  assign b_0 = b[0];
  assign b_1 = b[1];
  assign b_2 = b[2];
  assign b_3 = b[3];
  assign b_4 = b[4];
  assign b_5 = b[5];
  assign b_6 = b[6];
  assign b_7 = b[7];
  assign b_8 = b[8];
  assign b_9 = b[9];
  assign b_10 = b[10];
  assign b_11 = b[11];
  assign b_12 = b[12];
  assign b_13 = b[13];
  assign b_14 = b[14];
  assign b_15 = b[15];
  assign f_u_dadda_pg_rca16_and_13_0_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_13_0_y0 = f_u_dadda_pg_rca16_and_13_0_a_13 & f_u_dadda_pg_rca16_and_13_0_b_0;
  assign f_u_dadda_pg_rca16_and_12_1_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_12_1_y0 = f_u_dadda_pg_rca16_and_12_1_a_12 & f_u_dadda_pg_rca16_and_12_1_b_1;
  assign f_u_dadda_pg_rca16_ha0_f_u_dadda_pg_rca16_and_13_0_y0 = f_u_dadda_pg_rca16_and_13_0_y0;
  assign f_u_dadda_pg_rca16_ha0_f_u_dadda_pg_rca16_and_12_1_y0 = f_u_dadda_pg_rca16_and_12_1_y0;
  assign f_u_dadda_pg_rca16_ha0_y0 = f_u_dadda_pg_rca16_ha0_f_u_dadda_pg_rca16_and_13_0_y0 ^ f_u_dadda_pg_rca16_ha0_f_u_dadda_pg_rca16_and_12_1_y0;
  assign f_u_dadda_pg_rca16_ha0_y1 = f_u_dadda_pg_rca16_ha0_f_u_dadda_pg_rca16_and_13_0_y0 & f_u_dadda_pg_rca16_ha0_f_u_dadda_pg_rca16_and_12_1_y0;
  assign f_u_dadda_pg_rca16_and_14_0_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_14_0_y0 = f_u_dadda_pg_rca16_and_14_0_a_14 & f_u_dadda_pg_rca16_and_14_0_b_0;
  assign f_u_dadda_pg_rca16_and_13_1_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_13_1_y0 = f_u_dadda_pg_rca16_and_13_1_a_13 & f_u_dadda_pg_rca16_and_13_1_b_1;
  assign f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_ha0_y1 = f_u_dadda_pg_rca16_ha0_y1;
  assign f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_and_14_0_y0 = f_u_dadda_pg_rca16_and_14_0_y0;
  assign f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_and_13_1_y0 = f_u_dadda_pg_rca16_and_13_1_y0;
  assign f_u_dadda_pg_rca16_fa0_y0 = f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_ha0_y1 ^ f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_and_14_0_y0;
  assign f_u_dadda_pg_rca16_fa0_y1 = f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_ha0_y1 & f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_and_14_0_y0;
  assign f_u_dadda_pg_rca16_fa0_y2 = f_u_dadda_pg_rca16_fa0_y0 ^ f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_and_13_1_y0;
  assign f_u_dadda_pg_rca16_fa0_y3 = f_u_dadda_pg_rca16_fa0_y0 & f_u_dadda_pg_rca16_fa0_f_u_dadda_pg_rca16_and_13_1_y0;
  assign f_u_dadda_pg_rca16_fa0_y4 = f_u_dadda_pg_rca16_fa0_y1 | f_u_dadda_pg_rca16_fa0_y3;
  assign f_u_dadda_pg_rca16_and_12_2_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_12_2_y0 = f_u_dadda_pg_rca16_and_12_2_a_12 & f_u_dadda_pg_rca16_and_12_2_b_2;
  assign f_u_dadda_pg_rca16_and_11_3_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_11_3_y0 = f_u_dadda_pg_rca16_and_11_3_a_11 & f_u_dadda_pg_rca16_and_11_3_b_3;
  assign f_u_dadda_pg_rca16_ha1_f_u_dadda_pg_rca16_and_12_2_y0 = f_u_dadda_pg_rca16_and_12_2_y0;
  assign f_u_dadda_pg_rca16_ha1_f_u_dadda_pg_rca16_and_11_3_y0 = f_u_dadda_pg_rca16_and_11_3_y0;
  assign f_u_dadda_pg_rca16_ha1_y0 = f_u_dadda_pg_rca16_ha1_f_u_dadda_pg_rca16_and_12_2_y0 ^ f_u_dadda_pg_rca16_ha1_f_u_dadda_pg_rca16_and_11_3_y0;
  assign f_u_dadda_pg_rca16_ha1_y1 = f_u_dadda_pg_rca16_ha1_f_u_dadda_pg_rca16_and_12_2_y0 & f_u_dadda_pg_rca16_ha1_f_u_dadda_pg_rca16_and_11_3_y0;
  assign f_u_dadda_pg_rca16_and_15_0_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_15_0_y0 = f_u_dadda_pg_rca16_and_15_0_a_15 & f_u_dadda_pg_rca16_and_15_0_b_0;
  assign f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_ha1_y1 = f_u_dadda_pg_rca16_ha1_y1;
  assign f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_fa0_y4 = f_u_dadda_pg_rca16_fa0_y4;
  assign f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_and_15_0_y0 = f_u_dadda_pg_rca16_and_15_0_y0;
  assign f_u_dadda_pg_rca16_fa1_y0 = f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_ha1_y1 ^ f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_fa0_y4;
  assign f_u_dadda_pg_rca16_fa1_y1 = f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_ha1_y1 & f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_fa0_y4;
  assign f_u_dadda_pg_rca16_fa1_y2 = f_u_dadda_pg_rca16_fa1_y0 ^ f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_and_15_0_y0;
  assign f_u_dadda_pg_rca16_fa1_y3 = f_u_dadda_pg_rca16_fa1_y0 & f_u_dadda_pg_rca16_fa1_f_u_dadda_pg_rca16_and_15_0_y0;
  assign f_u_dadda_pg_rca16_fa1_y4 = f_u_dadda_pg_rca16_fa1_y1 | f_u_dadda_pg_rca16_fa1_y3;
  assign f_u_dadda_pg_rca16_and_14_1_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_14_1_y0 = f_u_dadda_pg_rca16_and_14_1_a_14 & f_u_dadda_pg_rca16_and_14_1_b_1;
  assign f_u_dadda_pg_rca16_and_13_2_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_13_2_y0 = f_u_dadda_pg_rca16_and_13_2_a_13 & f_u_dadda_pg_rca16_and_13_2_b_2;
  assign f_u_dadda_pg_rca16_and_12_3_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_12_3_y0 = f_u_dadda_pg_rca16_and_12_3_a_12 & f_u_dadda_pg_rca16_and_12_3_b_3;
  assign f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_14_1_y0 = f_u_dadda_pg_rca16_and_14_1_y0;
  assign f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_13_2_y0 = f_u_dadda_pg_rca16_and_13_2_y0;
  assign f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_12_3_y0 = f_u_dadda_pg_rca16_and_12_3_y0;
  assign f_u_dadda_pg_rca16_fa2_y0 = f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_14_1_y0 ^ f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_13_2_y0;
  assign f_u_dadda_pg_rca16_fa2_y1 = f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_14_1_y0 & f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_13_2_y0;
  assign f_u_dadda_pg_rca16_fa2_y2 = f_u_dadda_pg_rca16_fa2_y0 ^ f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_12_3_y0;
  assign f_u_dadda_pg_rca16_fa2_y3 = f_u_dadda_pg_rca16_fa2_y0 & f_u_dadda_pg_rca16_fa2_f_u_dadda_pg_rca16_and_12_3_y0;
  assign f_u_dadda_pg_rca16_fa2_y4 = f_u_dadda_pg_rca16_fa2_y1 | f_u_dadda_pg_rca16_fa2_y3;
  assign f_u_dadda_pg_rca16_and_11_4_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_11_4_y0 = f_u_dadda_pg_rca16_and_11_4_a_11 & f_u_dadda_pg_rca16_and_11_4_b_4;
  assign f_u_dadda_pg_rca16_and_10_5_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_10_5_y0 = f_u_dadda_pg_rca16_and_10_5_a_10 & f_u_dadda_pg_rca16_and_10_5_b_5;
  assign f_u_dadda_pg_rca16_ha2_f_u_dadda_pg_rca16_and_11_4_y0 = f_u_dadda_pg_rca16_and_11_4_y0;
  assign f_u_dadda_pg_rca16_ha2_f_u_dadda_pg_rca16_and_10_5_y0 = f_u_dadda_pg_rca16_and_10_5_y0;
  assign f_u_dadda_pg_rca16_ha2_y0 = f_u_dadda_pg_rca16_ha2_f_u_dadda_pg_rca16_and_11_4_y0 ^ f_u_dadda_pg_rca16_ha2_f_u_dadda_pg_rca16_and_10_5_y0;
  assign f_u_dadda_pg_rca16_ha2_y1 = f_u_dadda_pg_rca16_ha2_f_u_dadda_pg_rca16_and_11_4_y0 & f_u_dadda_pg_rca16_ha2_f_u_dadda_pg_rca16_and_10_5_y0;
  assign f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_ha2_y1 = f_u_dadda_pg_rca16_ha2_y1;
  assign f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_fa2_y4 = f_u_dadda_pg_rca16_fa2_y4;
  assign f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_fa1_y4 = f_u_dadda_pg_rca16_fa1_y4;
  assign f_u_dadda_pg_rca16_fa3_y0 = f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_ha2_y1 ^ f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_fa2_y4;
  assign f_u_dadda_pg_rca16_fa3_y1 = f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_ha2_y1 & f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_fa2_y4;
  assign f_u_dadda_pg_rca16_fa3_y2 = f_u_dadda_pg_rca16_fa3_y0 ^ f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_fa1_y4;
  assign f_u_dadda_pg_rca16_fa3_y3 = f_u_dadda_pg_rca16_fa3_y0 & f_u_dadda_pg_rca16_fa3_f_u_dadda_pg_rca16_fa1_y4;
  assign f_u_dadda_pg_rca16_fa3_y4 = f_u_dadda_pg_rca16_fa3_y1 | f_u_dadda_pg_rca16_fa3_y3;
  assign f_u_dadda_pg_rca16_and_15_1_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_15_1_y0 = f_u_dadda_pg_rca16_and_15_1_a_15 & f_u_dadda_pg_rca16_and_15_1_b_1;
  assign f_u_dadda_pg_rca16_and_14_2_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_14_2_y0 = f_u_dadda_pg_rca16_and_14_2_a_14 & f_u_dadda_pg_rca16_and_14_2_b_2;
  assign f_u_dadda_pg_rca16_and_13_3_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_13_3_y0 = f_u_dadda_pg_rca16_and_13_3_a_13 & f_u_dadda_pg_rca16_and_13_3_b_3;
  assign f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_15_1_y0 = f_u_dadda_pg_rca16_and_15_1_y0;
  assign f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_14_2_y0 = f_u_dadda_pg_rca16_and_14_2_y0;
  assign f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_13_3_y0 = f_u_dadda_pg_rca16_and_13_3_y0;
  assign f_u_dadda_pg_rca16_fa4_y0 = f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_15_1_y0 ^ f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_14_2_y0;
  assign f_u_dadda_pg_rca16_fa4_y1 = f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_15_1_y0 & f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_14_2_y0;
  assign f_u_dadda_pg_rca16_fa4_y2 = f_u_dadda_pg_rca16_fa4_y0 ^ f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_13_3_y0;
  assign f_u_dadda_pg_rca16_fa4_y3 = f_u_dadda_pg_rca16_fa4_y0 & f_u_dadda_pg_rca16_fa4_f_u_dadda_pg_rca16_and_13_3_y0;
  assign f_u_dadda_pg_rca16_fa4_y4 = f_u_dadda_pg_rca16_fa4_y1 | f_u_dadda_pg_rca16_fa4_y3;
  assign f_u_dadda_pg_rca16_and_12_4_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_12_4_y0 = f_u_dadda_pg_rca16_and_12_4_a_12 & f_u_dadda_pg_rca16_and_12_4_b_4;
  assign f_u_dadda_pg_rca16_and_11_5_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_11_5_y0 = f_u_dadda_pg_rca16_and_11_5_a_11 & f_u_dadda_pg_rca16_and_11_5_b_5;
  assign f_u_dadda_pg_rca16_ha3_f_u_dadda_pg_rca16_and_12_4_y0 = f_u_dadda_pg_rca16_and_12_4_y0;
  assign f_u_dadda_pg_rca16_ha3_f_u_dadda_pg_rca16_and_11_5_y0 = f_u_dadda_pg_rca16_and_11_5_y0;
  assign f_u_dadda_pg_rca16_ha3_y0 = f_u_dadda_pg_rca16_ha3_f_u_dadda_pg_rca16_and_12_4_y0 ^ f_u_dadda_pg_rca16_ha3_f_u_dadda_pg_rca16_and_11_5_y0;
  assign f_u_dadda_pg_rca16_ha3_y1 = f_u_dadda_pg_rca16_ha3_f_u_dadda_pg_rca16_and_12_4_y0 & f_u_dadda_pg_rca16_ha3_f_u_dadda_pg_rca16_and_11_5_y0;
  assign f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_ha3_y1 = f_u_dadda_pg_rca16_ha3_y1;
  assign f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_fa4_y4 = f_u_dadda_pg_rca16_fa4_y4;
  assign f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_fa3_y4 = f_u_dadda_pg_rca16_fa3_y4;
  assign f_u_dadda_pg_rca16_fa5_y0 = f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_ha3_y1 ^ f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_fa4_y4;
  assign f_u_dadda_pg_rca16_fa5_y1 = f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_ha3_y1 & f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_fa4_y4;
  assign f_u_dadda_pg_rca16_fa5_y2 = f_u_dadda_pg_rca16_fa5_y0 ^ f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_fa3_y4;
  assign f_u_dadda_pg_rca16_fa5_y3 = f_u_dadda_pg_rca16_fa5_y0 & f_u_dadda_pg_rca16_fa5_f_u_dadda_pg_rca16_fa3_y4;
  assign f_u_dadda_pg_rca16_fa5_y4 = f_u_dadda_pg_rca16_fa5_y1 | f_u_dadda_pg_rca16_fa5_y3;
  assign f_u_dadda_pg_rca16_and_15_2_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_15_2_y0 = f_u_dadda_pg_rca16_and_15_2_a_15 & f_u_dadda_pg_rca16_and_15_2_b_2;
  assign f_u_dadda_pg_rca16_and_14_3_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_14_3_y0 = f_u_dadda_pg_rca16_and_14_3_a_14 & f_u_dadda_pg_rca16_and_14_3_b_3;
  assign f_u_dadda_pg_rca16_and_13_4_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_13_4_y0 = f_u_dadda_pg_rca16_and_13_4_a_13 & f_u_dadda_pg_rca16_and_13_4_b_4;
  assign f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_15_2_y0 = f_u_dadda_pg_rca16_and_15_2_y0;
  assign f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_14_3_y0 = f_u_dadda_pg_rca16_and_14_3_y0;
  assign f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_13_4_y0 = f_u_dadda_pg_rca16_and_13_4_y0;
  assign f_u_dadda_pg_rca16_fa6_y0 = f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_15_2_y0 ^ f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_14_3_y0;
  assign f_u_dadda_pg_rca16_fa6_y1 = f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_15_2_y0 & f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_14_3_y0;
  assign f_u_dadda_pg_rca16_fa6_y2 = f_u_dadda_pg_rca16_fa6_y0 ^ f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_13_4_y0;
  assign f_u_dadda_pg_rca16_fa6_y3 = f_u_dadda_pg_rca16_fa6_y0 & f_u_dadda_pg_rca16_fa6_f_u_dadda_pg_rca16_and_13_4_y0;
  assign f_u_dadda_pg_rca16_fa6_y4 = f_u_dadda_pg_rca16_fa6_y1 | f_u_dadda_pg_rca16_fa6_y3;
  assign f_u_dadda_pg_rca16_and_15_3_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_15_3_y0 = f_u_dadda_pg_rca16_and_15_3_a_15 & f_u_dadda_pg_rca16_and_15_3_b_3;
  assign f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_fa6_y4 = f_u_dadda_pg_rca16_fa6_y4;
  assign f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_fa5_y4 = f_u_dadda_pg_rca16_fa5_y4;
  assign f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_and_15_3_y0 = f_u_dadda_pg_rca16_and_15_3_y0;
  assign f_u_dadda_pg_rca16_fa7_y0 = f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_fa6_y4 ^ f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_fa5_y4;
  assign f_u_dadda_pg_rca16_fa7_y1 = f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_fa6_y4 & f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_fa5_y4;
  assign f_u_dadda_pg_rca16_fa7_y2 = f_u_dadda_pg_rca16_fa7_y0 ^ f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_and_15_3_y0;
  assign f_u_dadda_pg_rca16_fa7_y3 = f_u_dadda_pg_rca16_fa7_y0 & f_u_dadda_pg_rca16_fa7_f_u_dadda_pg_rca16_and_15_3_y0;
  assign f_u_dadda_pg_rca16_fa7_y4 = f_u_dadda_pg_rca16_fa7_y1 | f_u_dadda_pg_rca16_fa7_y3;
  assign f_u_dadda_pg_rca16_and_4_0_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_4_0_y0 = f_u_dadda_pg_rca16_and_4_0_a_4 & f_u_dadda_pg_rca16_and_4_0_b_0;
  assign f_u_dadda_pg_rca16_and_3_1_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_3_1_y0 = f_u_dadda_pg_rca16_and_3_1_a_3 & f_u_dadda_pg_rca16_and_3_1_b_1;
  assign f_u_dadda_pg_rca16_ha4_f_u_dadda_pg_rca16_and_4_0_y0 = f_u_dadda_pg_rca16_and_4_0_y0;
  assign f_u_dadda_pg_rca16_ha4_f_u_dadda_pg_rca16_and_3_1_y0 = f_u_dadda_pg_rca16_and_3_1_y0;
  assign f_u_dadda_pg_rca16_ha4_y0 = f_u_dadda_pg_rca16_ha4_f_u_dadda_pg_rca16_and_4_0_y0 ^ f_u_dadda_pg_rca16_ha4_f_u_dadda_pg_rca16_and_3_1_y0;
  assign f_u_dadda_pg_rca16_ha4_y1 = f_u_dadda_pg_rca16_ha4_f_u_dadda_pg_rca16_and_4_0_y0 & f_u_dadda_pg_rca16_ha4_f_u_dadda_pg_rca16_and_3_1_y0;
  assign f_u_dadda_pg_rca16_and_5_0_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_5_0_y0 = f_u_dadda_pg_rca16_and_5_0_a_5 & f_u_dadda_pg_rca16_and_5_0_b_0;
  assign f_u_dadda_pg_rca16_and_4_1_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_4_1_y0 = f_u_dadda_pg_rca16_and_4_1_a_4 & f_u_dadda_pg_rca16_and_4_1_b_1;
  assign f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_ha4_y1 = f_u_dadda_pg_rca16_ha4_y1;
  assign f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_and_5_0_y0 = f_u_dadda_pg_rca16_and_5_0_y0;
  assign f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_and_4_1_y0 = f_u_dadda_pg_rca16_and_4_1_y0;
  assign f_u_dadda_pg_rca16_fa8_y0 = f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_ha4_y1 ^ f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_and_5_0_y0;
  assign f_u_dadda_pg_rca16_fa8_y1 = f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_ha4_y1 & f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_and_5_0_y0;
  assign f_u_dadda_pg_rca16_fa8_y2 = f_u_dadda_pg_rca16_fa8_y0 ^ f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_and_4_1_y0;
  assign f_u_dadda_pg_rca16_fa8_y3 = f_u_dadda_pg_rca16_fa8_y0 & f_u_dadda_pg_rca16_fa8_f_u_dadda_pg_rca16_and_4_1_y0;
  assign f_u_dadda_pg_rca16_fa8_y4 = f_u_dadda_pg_rca16_fa8_y1 | f_u_dadda_pg_rca16_fa8_y3;
  assign f_u_dadda_pg_rca16_and_3_2_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_3_2_y0 = f_u_dadda_pg_rca16_and_3_2_a_3 & f_u_dadda_pg_rca16_and_3_2_b_2;
  assign f_u_dadda_pg_rca16_and_2_3_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_2_3_y0 = f_u_dadda_pg_rca16_and_2_3_a_2 & f_u_dadda_pg_rca16_and_2_3_b_3;
  assign f_u_dadda_pg_rca16_ha5_f_u_dadda_pg_rca16_and_3_2_y0 = f_u_dadda_pg_rca16_and_3_2_y0;
  assign f_u_dadda_pg_rca16_ha5_f_u_dadda_pg_rca16_and_2_3_y0 = f_u_dadda_pg_rca16_and_2_3_y0;
  assign f_u_dadda_pg_rca16_ha5_y0 = f_u_dadda_pg_rca16_ha5_f_u_dadda_pg_rca16_and_3_2_y0 ^ f_u_dadda_pg_rca16_ha5_f_u_dadda_pg_rca16_and_2_3_y0;
  assign f_u_dadda_pg_rca16_ha5_y1 = f_u_dadda_pg_rca16_ha5_f_u_dadda_pg_rca16_and_3_2_y0 & f_u_dadda_pg_rca16_ha5_f_u_dadda_pg_rca16_and_2_3_y0;
  assign f_u_dadda_pg_rca16_and_6_0_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_6_0_y0 = f_u_dadda_pg_rca16_and_6_0_a_6 & f_u_dadda_pg_rca16_and_6_0_b_0;
  assign f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_ha5_y1 = f_u_dadda_pg_rca16_ha5_y1;
  assign f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_fa8_y4 = f_u_dadda_pg_rca16_fa8_y4;
  assign f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_and_6_0_y0 = f_u_dadda_pg_rca16_and_6_0_y0;
  assign f_u_dadda_pg_rca16_fa9_y0 = f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_ha5_y1 ^ f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_fa8_y4;
  assign f_u_dadda_pg_rca16_fa9_y1 = f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_ha5_y1 & f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_fa8_y4;
  assign f_u_dadda_pg_rca16_fa9_y2 = f_u_dadda_pg_rca16_fa9_y0 ^ f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_and_6_0_y0;
  assign f_u_dadda_pg_rca16_fa9_y3 = f_u_dadda_pg_rca16_fa9_y0 & f_u_dadda_pg_rca16_fa9_f_u_dadda_pg_rca16_and_6_0_y0;
  assign f_u_dadda_pg_rca16_fa9_y4 = f_u_dadda_pg_rca16_fa9_y1 | f_u_dadda_pg_rca16_fa9_y3;
  assign f_u_dadda_pg_rca16_and_5_1_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_5_1_y0 = f_u_dadda_pg_rca16_and_5_1_a_5 & f_u_dadda_pg_rca16_and_5_1_b_1;
  assign f_u_dadda_pg_rca16_and_4_2_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_4_2_y0 = f_u_dadda_pg_rca16_and_4_2_a_4 & f_u_dadda_pg_rca16_and_4_2_b_2;
  assign f_u_dadda_pg_rca16_and_3_3_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_3_3_y0 = f_u_dadda_pg_rca16_and_3_3_a_3 & f_u_dadda_pg_rca16_and_3_3_b_3;
  assign f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_5_1_y0 = f_u_dadda_pg_rca16_and_5_1_y0;
  assign f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_4_2_y0 = f_u_dadda_pg_rca16_and_4_2_y0;
  assign f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_3_3_y0 = f_u_dadda_pg_rca16_and_3_3_y0;
  assign f_u_dadda_pg_rca16_fa10_y0 = f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_5_1_y0 ^ f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_4_2_y0;
  assign f_u_dadda_pg_rca16_fa10_y1 = f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_5_1_y0 & f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_4_2_y0;
  assign f_u_dadda_pg_rca16_fa10_y2 = f_u_dadda_pg_rca16_fa10_y0 ^ f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_3_3_y0;
  assign f_u_dadda_pg_rca16_fa10_y3 = f_u_dadda_pg_rca16_fa10_y0 & f_u_dadda_pg_rca16_fa10_f_u_dadda_pg_rca16_and_3_3_y0;
  assign f_u_dadda_pg_rca16_fa10_y4 = f_u_dadda_pg_rca16_fa10_y1 | f_u_dadda_pg_rca16_fa10_y3;
  assign f_u_dadda_pg_rca16_and_2_4_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_2_4_y0 = f_u_dadda_pg_rca16_and_2_4_a_2 & f_u_dadda_pg_rca16_and_2_4_b_4;
  assign f_u_dadda_pg_rca16_and_1_5_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_1_5_y0 = f_u_dadda_pg_rca16_and_1_5_a_1 & f_u_dadda_pg_rca16_and_1_5_b_5;
  assign f_u_dadda_pg_rca16_ha6_f_u_dadda_pg_rca16_and_2_4_y0 = f_u_dadda_pg_rca16_and_2_4_y0;
  assign f_u_dadda_pg_rca16_ha6_f_u_dadda_pg_rca16_and_1_5_y0 = f_u_dadda_pg_rca16_and_1_5_y0;
  assign f_u_dadda_pg_rca16_ha6_y0 = f_u_dadda_pg_rca16_ha6_f_u_dadda_pg_rca16_and_2_4_y0 ^ f_u_dadda_pg_rca16_ha6_f_u_dadda_pg_rca16_and_1_5_y0;
  assign f_u_dadda_pg_rca16_ha6_y1 = f_u_dadda_pg_rca16_ha6_f_u_dadda_pg_rca16_and_2_4_y0 & f_u_dadda_pg_rca16_ha6_f_u_dadda_pg_rca16_and_1_5_y0;
  assign f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_ha6_y1 = f_u_dadda_pg_rca16_ha6_y1;
  assign f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_fa10_y4 = f_u_dadda_pg_rca16_fa10_y4;
  assign f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_fa9_y4 = f_u_dadda_pg_rca16_fa9_y4;
  assign f_u_dadda_pg_rca16_fa11_y0 = f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_ha6_y1 ^ f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_fa10_y4;
  assign f_u_dadda_pg_rca16_fa11_y1 = f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_ha6_y1 & f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_fa10_y4;
  assign f_u_dadda_pg_rca16_fa11_y2 = f_u_dadda_pg_rca16_fa11_y0 ^ f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_fa9_y4;
  assign f_u_dadda_pg_rca16_fa11_y3 = f_u_dadda_pg_rca16_fa11_y0 & f_u_dadda_pg_rca16_fa11_f_u_dadda_pg_rca16_fa9_y4;
  assign f_u_dadda_pg_rca16_fa11_y4 = f_u_dadda_pg_rca16_fa11_y1 | f_u_dadda_pg_rca16_fa11_y3;
  assign f_u_dadda_pg_rca16_and_7_0_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_7_0_y0 = f_u_dadda_pg_rca16_and_7_0_a_7 & f_u_dadda_pg_rca16_and_7_0_b_0;
  assign f_u_dadda_pg_rca16_and_6_1_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_6_1_y0 = f_u_dadda_pg_rca16_and_6_1_a_6 & f_u_dadda_pg_rca16_and_6_1_b_1;
  assign f_u_dadda_pg_rca16_and_5_2_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_5_2_y0 = f_u_dadda_pg_rca16_and_5_2_a_5 & f_u_dadda_pg_rca16_and_5_2_b_2;
  assign f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_7_0_y0 = f_u_dadda_pg_rca16_and_7_0_y0;
  assign f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_6_1_y0 = f_u_dadda_pg_rca16_and_6_1_y0;
  assign f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_5_2_y0 = f_u_dadda_pg_rca16_and_5_2_y0;
  assign f_u_dadda_pg_rca16_fa12_y0 = f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_7_0_y0 ^ f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_6_1_y0;
  assign f_u_dadda_pg_rca16_fa12_y1 = f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_7_0_y0 & f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_6_1_y0;
  assign f_u_dadda_pg_rca16_fa12_y2 = f_u_dadda_pg_rca16_fa12_y0 ^ f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_5_2_y0;
  assign f_u_dadda_pg_rca16_fa12_y3 = f_u_dadda_pg_rca16_fa12_y0 & f_u_dadda_pg_rca16_fa12_f_u_dadda_pg_rca16_and_5_2_y0;
  assign f_u_dadda_pg_rca16_fa12_y4 = f_u_dadda_pg_rca16_fa12_y1 | f_u_dadda_pg_rca16_fa12_y3;
  assign f_u_dadda_pg_rca16_and_4_3_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_4_3_y0 = f_u_dadda_pg_rca16_and_4_3_a_4 & f_u_dadda_pg_rca16_and_4_3_b_3;
  assign f_u_dadda_pg_rca16_and_3_4_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_3_4_y0 = f_u_dadda_pg_rca16_and_3_4_a_3 & f_u_dadda_pg_rca16_and_3_4_b_4;
  assign f_u_dadda_pg_rca16_and_2_5_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_2_5_y0 = f_u_dadda_pg_rca16_and_2_5_a_2 & f_u_dadda_pg_rca16_and_2_5_b_5;
  assign f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_4_3_y0 = f_u_dadda_pg_rca16_and_4_3_y0;
  assign f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_3_4_y0 = f_u_dadda_pg_rca16_and_3_4_y0;
  assign f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_2_5_y0 = f_u_dadda_pg_rca16_and_2_5_y0;
  assign f_u_dadda_pg_rca16_fa13_y0 = f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_4_3_y0 ^ f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_3_4_y0;
  assign f_u_dadda_pg_rca16_fa13_y1 = f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_4_3_y0 & f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_3_4_y0;
  assign f_u_dadda_pg_rca16_fa13_y2 = f_u_dadda_pg_rca16_fa13_y0 ^ f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_2_5_y0;
  assign f_u_dadda_pg_rca16_fa13_y3 = f_u_dadda_pg_rca16_fa13_y0 & f_u_dadda_pg_rca16_fa13_f_u_dadda_pg_rca16_and_2_5_y0;
  assign f_u_dadda_pg_rca16_fa13_y4 = f_u_dadda_pg_rca16_fa13_y1 | f_u_dadda_pg_rca16_fa13_y3;
  assign f_u_dadda_pg_rca16_and_1_6_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_1_6_y0 = f_u_dadda_pg_rca16_and_1_6_a_1 & f_u_dadda_pg_rca16_and_1_6_b_6;
  assign f_u_dadda_pg_rca16_and_0_7_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_0_7_y0 = f_u_dadda_pg_rca16_and_0_7_a_0 & f_u_dadda_pg_rca16_and_0_7_b_7;
  assign f_u_dadda_pg_rca16_ha7_f_u_dadda_pg_rca16_and_1_6_y0 = f_u_dadda_pg_rca16_and_1_6_y0;
  assign f_u_dadda_pg_rca16_ha7_f_u_dadda_pg_rca16_and_0_7_y0 = f_u_dadda_pg_rca16_and_0_7_y0;
  assign f_u_dadda_pg_rca16_ha7_y0 = f_u_dadda_pg_rca16_ha7_f_u_dadda_pg_rca16_and_1_6_y0 ^ f_u_dadda_pg_rca16_ha7_f_u_dadda_pg_rca16_and_0_7_y0;
  assign f_u_dadda_pg_rca16_ha7_y1 = f_u_dadda_pg_rca16_ha7_f_u_dadda_pg_rca16_and_1_6_y0 & f_u_dadda_pg_rca16_ha7_f_u_dadda_pg_rca16_and_0_7_y0;
  assign f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_ha7_y1 = f_u_dadda_pg_rca16_ha7_y1;
  assign f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_fa13_y4 = f_u_dadda_pg_rca16_fa13_y4;
  assign f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_fa12_y4 = f_u_dadda_pg_rca16_fa12_y4;
  assign f_u_dadda_pg_rca16_fa14_y0 = f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_ha7_y1 ^ f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_fa13_y4;
  assign f_u_dadda_pg_rca16_fa14_y1 = f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_ha7_y1 & f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_fa13_y4;
  assign f_u_dadda_pg_rca16_fa14_y2 = f_u_dadda_pg_rca16_fa14_y0 ^ f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_fa12_y4;
  assign f_u_dadda_pg_rca16_fa14_y3 = f_u_dadda_pg_rca16_fa14_y0 & f_u_dadda_pg_rca16_fa14_f_u_dadda_pg_rca16_fa12_y4;
  assign f_u_dadda_pg_rca16_fa14_y4 = f_u_dadda_pg_rca16_fa14_y1 | f_u_dadda_pg_rca16_fa14_y3;
  assign f_u_dadda_pg_rca16_and_8_0_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_8_0_y0 = f_u_dadda_pg_rca16_and_8_0_a_8 & f_u_dadda_pg_rca16_and_8_0_b_0;
  assign f_u_dadda_pg_rca16_and_7_1_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_7_1_y0 = f_u_dadda_pg_rca16_and_7_1_a_7 & f_u_dadda_pg_rca16_and_7_1_b_1;
  assign f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_fa11_y4 = f_u_dadda_pg_rca16_fa11_y4;
  assign f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_and_8_0_y0 = f_u_dadda_pg_rca16_and_8_0_y0;
  assign f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_and_7_1_y0 = f_u_dadda_pg_rca16_and_7_1_y0;
  assign f_u_dadda_pg_rca16_fa15_y0 = f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_fa11_y4 ^ f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_and_8_0_y0;
  assign f_u_dadda_pg_rca16_fa15_y1 = f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_fa11_y4 & f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_and_8_0_y0;
  assign f_u_dadda_pg_rca16_fa15_y2 = f_u_dadda_pg_rca16_fa15_y0 ^ f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_and_7_1_y0;
  assign f_u_dadda_pg_rca16_fa15_y3 = f_u_dadda_pg_rca16_fa15_y0 & f_u_dadda_pg_rca16_fa15_f_u_dadda_pg_rca16_and_7_1_y0;
  assign f_u_dadda_pg_rca16_fa15_y4 = f_u_dadda_pg_rca16_fa15_y1 | f_u_dadda_pg_rca16_fa15_y3;
  assign f_u_dadda_pg_rca16_and_6_2_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_6_2_y0 = f_u_dadda_pg_rca16_and_6_2_a_6 & f_u_dadda_pg_rca16_and_6_2_b_2;
  assign f_u_dadda_pg_rca16_and_5_3_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_5_3_y0 = f_u_dadda_pg_rca16_and_5_3_a_5 & f_u_dadda_pg_rca16_and_5_3_b_3;
  assign f_u_dadda_pg_rca16_and_4_4_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_4_4_y0 = f_u_dadda_pg_rca16_and_4_4_a_4 & f_u_dadda_pg_rca16_and_4_4_b_4;
  assign f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_6_2_y0 = f_u_dadda_pg_rca16_and_6_2_y0;
  assign f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_5_3_y0 = f_u_dadda_pg_rca16_and_5_3_y0;
  assign f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_4_4_y0 = f_u_dadda_pg_rca16_and_4_4_y0;
  assign f_u_dadda_pg_rca16_fa16_y0 = f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_6_2_y0 ^ f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_5_3_y0;
  assign f_u_dadda_pg_rca16_fa16_y1 = f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_6_2_y0 & f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_5_3_y0;
  assign f_u_dadda_pg_rca16_fa16_y2 = f_u_dadda_pg_rca16_fa16_y0 ^ f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_4_4_y0;
  assign f_u_dadda_pg_rca16_fa16_y3 = f_u_dadda_pg_rca16_fa16_y0 & f_u_dadda_pg_rca16_fa16_f_u_dadda_pg_rca16_and_4_4_y0;
  assign f_u_dadda_pg_rca16_fa16_y4 = f_u_dadda_pg_rca16_fa16_y1 | f_u_dadda_pg_rca16_fa16_y3;
  assign f_u_dadda_pg_rca16_and_3_5_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_3_5_y0 = f_u_dadda_pg_rca16_and_3_5_a_3 & f_u_dadda_pg_rca16_and_3_5_b_5;
  assign f_u_dadda_pg_rca16_and_2_6_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_2_6_y0 = f_u_dadda_pg_rca16_and_2_6_a_2 & f_u_dadda_pg_rca16_and_2_6_b_6;
  assign f_u_dadda_pg_rca16_and_1_7_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_1_7_y0 = f_u_dadda_pg_rca16_and_1_7_a_1 & f_u_dadda_pg_rca16_and_1_7_b_7;
  assign f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_3_5_y0 = f_u_dadda_pg_rca16_and_3_5_y0;
  assign f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_2_6_y0 = f_u_dadda_pg_rca16_and_2_6_y0;
  assign f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_1_7_y0 = f_u_dadda_pg_rca16_and_1_7_y0;
  assign f_u_dadda_pg_rca16_fa17_y0 = f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_3_5_y0 ^ f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_2_6_y0;
  assign f_u_dadda_pg_rca16_fa17_y1 = f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_3_5_y0 & f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_2_6_y0;
  assign f_u_dadda_pg_rca16_fa17_y2 = f_u_dadda_pg_rca16_fa17_y0 ^ f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_1_7_y0;
  assign f_u_dadda_pg_rca16_fa17_y3 = f_u_dadda_pg_rca16_fa17_y0 & f_u_dadda_pg_rca16_fa17_f_u_dadda_pg_rca16_and_1_7_y0;
  assign f_u_dadda_pg_rca16_fa17_y4 = f_u_dadda_pg_rca16_fa17_y1 | f_u_dadda_pg_rca16_fa17_y3;
  assign f_u_dadda_pg_rca16_and_0_8_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_0_8_y0 = f_u_dadda_pg_rca16_and_0_8_a_0 & f_u_dadda_pg_rca16_and_0_8_b_8;
  assign f_u_dadda_pg_rca16_ha8_f_u_dadda_pg_rca16_and_0_8_y0 = f_u_dadda_pg_rca16_and_0_8_y0;
  assign f_u_dadda_pg_rca16_ha8_f_u_dadda_pg_rca16_fa14_y2 = f_u_dadda_pg_rca16_fa14_y2;
  assign f_u_dadda_pg_rca16_ha8_y0 = f_u_dadda_pg_rca16_ha8_f_u_dadda_pg_rca16_and_0_8_y0 ^ f_u_dadda_pg_rca16_ha8_f_u_dadda_pg_rca16_fa14_y2;
  assign f_u_dadda_pg_rca16_ha8_y1 = f_u_dadda_pg_rca16_ha8_f_u_dadda_pg_rca16_and_0_8_y0 & f_u_dadda_pg_rca16_ha8_f_u_dadda_pg_rca16_fa14_y2;
  assign f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_ha8_y1 = f_u_dadda_pg_rca16_ha8_y1;
  assign f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_fa17_y4 = f_u_dadda_pg_rca16_fa17_y4;
  assign f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_fa16_y4 = f_u_dadda_pg_rca16_fa16_y4;
  assign f_u_dadda_pg_rca16_fa18_y0 = f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_ha8_y1 ^ f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_fa17_y4;
  assign f_u_dadda_pg_rca16_fa18_y1 = f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_ha8_y1 & f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_fa17_y4;
  assign f_u_dadda_pg_rca16_fa18_y2 = f_u_dadda_pg_rca16_fa18_y0 ^ f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_fa16_y4;
  assign f_u_dadda_pg_rca16_fa18_y3 = f_u_dadda_pg_rca16_fa18_y0 & f_u_dadda_pg_rca16_fa18_f_u_dadda_pg_rca16_fa16_y4;
  assign f_u_dadda_pg_rca16_fa18_y4 = f_u_dadda_pg_rca16_fa18_y1 | f_u_dadda_pg_rca16_fa18_y3;
  assign f_u_dadda_pg_rca16_and_9_0_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_9_0_y0 = f_u_dadda_pg_rca16_and_9_0_a_9 & f_u_dadda_pg_rca16_and_9_0_b_0;
  assign f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_fa15_y4 = f_u_dadda_pg_rca16_fa15_y4;
  assign f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_fa14_y4 = f_u_dadda_pg_rca16_fa14_y4;
  assign f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_and_9_0_y0 = f_u_dadda_pg_rca16_and_9_0_y0;
  assign f_u_dadda_pg_rca16_fa19_y0 = f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_fa15_y4 ^ f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_fa14_y4;
  assign f_u_dadda_pg_rca16_fa19_y1 = f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_fa15_y4 & f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_fa14_y4;
  assign f_u_dadda_pg_rca16_fa19_y2 = f_u_dadda_pg_rca16_fa19_y0 ^ f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_and_9_0_y0;
  assign f_u_dadda_pg_rca16_fa19_y3 = f_u_dadda_pg_rca16_fa19_y0 & f_u_dadda_pg_rca16_fa19_f_u_dadda_pg_rca16_and_9_0_y0;
  assign f_u_dadda_pg_rca16_fa19_y4 = f_u_dadda_pg_rca16_fa19_y1 | f_u_dadda_pg_rca16_fa19_y3;
  assign f_u_dadda_pg_rca16_and_8_1_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_8_1_y0 = f_u_dadda_pg_rca16_and_8_1_a_8 & f_u_dadda_pg_rca16_and_8_1_b_1;
  assign f_u_dadda_pg_rca16_and_7_2_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_7_2_y0 = f_u_dadda_pg_rca16_and_7_2_a_7 & f_u_dadda_pg_rca16_and_7_2_b_2;
  assign f_u_dadda_pg_rca16_and_6_3_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_6_3_y0 = f_u_dadda_pg_rca16_and_6_3_a_6 & f_u_dadda_pg_rca16_and_6_3_b_3;
  assign f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_8_1_y0 = f_u_dadda_pg_rca16_and_8_1_y0;
  assign f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_7_2_y0 = f_u_dadda_pg_rca16_and_7_2_y0;
  assign f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_6_3_y0 = f_u_dadda_pg_rca16_and_6_3_y0;
  assign f_u_dadda_pg_rca16_fa20_y0 = f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_8_1_y0 ^ f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_7_2_y0;
  assign f_u_dadda_pg_rca16_fa20_y1 = f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_8_1_y0 & f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_7_2_y0;
  assign f_u_dadda_pg_rca16_fa20_y2 = f_u_dadda_pg_rca16_fa20_y0 ^ f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_6_3_y0;
  assign f_u_dadda_pg_rca16_fa20_y3 = f_u_dadda_pg_rca16_fa20_y0 & f_u_dadda_pg_rca16_fa20_f_u_dadda_pg_rca16_and_6_3_y0;
  assign f_u_dadda_pg_rca16_fa20_y4 = f_u_dadda_pg_rca16_fa20_y1 | f_u_dadda_pg_rca16_fa20_y3;
  assign f_u_dadda_pg_rca16_and_5_4_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_5_4_y0 = f_u_dadda_pg_rca16_and_5_4_a_5 & f_u_dadda_pg_rca16_and_5_4_b_4;
  assign f_u_dadda_pg_rca16_and_4_5_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_4_5_y0 = f_u_dadda_pg_rca16_and_4_5_a_4 & f_u_dadda_pg_rca16_and_4_5_b_5;
  assign f_u_dadda_pg_rca16_and_3_6_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_3_6_y0 = f_u_dadda_pg_rca16_and_3_6_a_3 & f_u_dadda_pg_rca16_and_3_6_b_6;
  assign f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_5_4_y0 = f_u_dadda_pg_rca16_and_5_4_y0;
  assign f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_4_5_y0 = f_u_dadda_pg_rca16_and_4_5_y0;
  assign f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_3_6_y0 = f_u_dadda_pg_rca16_and_3_6_y0;
  assign f_u_dadda_pg_rca16_fa21_y0 = f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_5_4_y0 ^ f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_4_5_y0;
  assign f_u_dadda_pg_rca16_fa21_y1 = f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_5_4_y0 & f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_4_5_y0;
  assign f_u_dadda_pg_rca16_fa21_y2 = f_u_dadda_pg_rca16_fa21_y0 ^ f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_3_6_y0;
  assign f_u_dadda_pg_rca16_fa21_y3 = f_u_dadda_pg_rca16_fa21_y0 & f_u_dadda_pg_rca16_fa21_f_u_dadda_pg_rca16_and_3_6_y0;
  assign f_u_dadda_pg_rca16_fa21_y4 = f_u_dadda_pg_rca16_fa21_y1 | f_u_dadda_pg_rca16_fa21_y3;
  assign f_u_dadda_pg_rca16_and_2_7_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_2_7_y0 = f_u_dadda_pg_rca16_and_2_7_a_2 & f_u_dadda_pg_rca16_and_2_7_b_7;
  assign f_u_dadda_pg_rca16_and_1_8_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_1_8_y0 = f_u_dadda_pg_rca16_and_1_8_a_1 & f_u_dadda_pg_rca16_and_1_8_b_8;
  assign f_u_dadda_pg_rca16_and_0_9_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_0_9_y0 = f_u_dadda_pg_rca16_and_0_9_a_0 & f_u_dadda_pg_rca16_and_0_9_b_9;
  assign f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_2_7_y0 = f_u_dadda_pg_rca16_and_2_7_y0;
  assign f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_1_8_y0 = f_u_dadda_pg_rca16_and_1_8_y0;
  assign f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_0_9_y0 = f_u_dadda_pg_rca16_and_0_9_y0;
  assign f_u_dadda_pg_rca16_fa22_y0 = f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_2_7_y0 ^ f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_1_8_y0;
  assign f_u_dadda_pg_rca16_fa22_y1 = f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_2_7_y0 & f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_1_8_y0;
  assign f_u_dadda_pg_rca16_fa22_y2 = f_u_dadda_pg_rca16_fa22_y0 ^ f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_0_9_y0;
  assign f_u_dadda_pg_rca16_fa22_y3 = f_u_dadda_pg_rca16_fa22_y0 & f_u_dadda_pg_rca16_fa22_f_u_dadda_pg_rca16_and_0_9_y0;
  assign f_u_dadda_pg_rca16_fa22_y4 = f_u_dadda_pg_rca16_fa22_y1 | f_u_dadda_pg_rca16_fa22_y3;
  assign f_u_dadda_pg_rca16_ha9_f_u_dadda_pg_rca16_fa18_y2 = f_u_dadda_pg_rca16_fa18_y2;
  assign f_u_dadda_pg_rca16_ha9_f_u_dadda_pg_rca16_fa19_y2 = f_u_dadda_pg_rca16_fa19_y2;
  assign f_u_dadda_pg_rca16_ha9_y0 = f_u_dadda_pg_rca16_ha9_f_u_dadda_pg_rca16_fa18_y2 ^ f_u_dadda_pg_rca16_ha9_f_u_dadda_pg_rca16_fa19_y2;
  assign f_u_dadda_pg_rca16_ha9_y1 = f_u_dadda_pg_rca16_ha9_f_u_dadda_pg_rca16_fa18_y2 & f_u_dadda_pg_rca16_ha9_f_u_dadda_pg_rca16_fa19_y2;
  assign f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_ha9_y1 = f_u_dadda_pg_rca16_ha9_y1;
  assign f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_fa22_y4 = f_u_dadda_pg_rca16_fa22_y4;
  assign f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_fa21_y4 = f_u_dadda_pg_rca16_fa21_y4;
  assign f_u_dadda_pg_rca16_fa23_y0 = f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_ha9_y1 ^ f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_fa22_y4;
  assign f_u_dadda_pg_rca16_fa23_y1 = f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_ha9_y1 & f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_fa22_y4;
  assign f_u_dadda_pg_rca16_fa23_y2 = f_u_dadda_pg_rca16_fa23_y0 ^ f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_fa21_y4;
  assign f_u_dadda_pg_rca16_fa23_y3 = f_u_dadda_pg_rca16_fa23_y0 & f_u_dadda_pg_rca16_fa23_f_u_dadda_pg_rca16_fa21_y4;
  assign f_u_dadda_pg_rca16_fa23_y4 = f_u_dadda_pg_rca16_fa23_y1 | f_u_dadda_pg_rca16_fa23_y3;
  assign f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa20_y4 = f_u_dadda_pg_rca16_fa20_y4;
  assign f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa19_y4 = f_u_dadda_pg_rca16_fa19_y4;
  assign f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa18_y4 = f_u_dadda_pg_rca16_fa18_y4;
  assign f_u_dadda_pg_rca16_fa24_y0 = f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa20_y4 ^ f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa19_y4;
  assign f_u_dadda_pg_rca16_fa24_y1 = f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa20_y4 & f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa19_y4;
  assign f_u_dadda_pg_rca16_fa24_y2 = f_u_dadda_pg_rca16_fa24_y0 ^ f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa18_y4;
  assign f_u_dadda_pg_rca16_fa24_y3 = f_u_dadda_pg_rca16_fa24_y0 & f_u_dadda_pg_rca16_fa24_f_u_dadda_pg_rca16_fa18_y4;
  assign f_u_dadda_pg_rca16_fa24_y4 = f_u_dadda_pg_rca16_fa24_y1 | f_u_dadda_pg_rca16_fa24_y3;
  assign f_u_dadda_pg_rca16_and_10_0_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_10_0_y0 = f_u_dadda_pg_rca16_and_10_0_a_10 & f_u_dadda_pg_rca16_and_10_0_b_0;
  assign f_u_dadda_pg_rca16_and_9_1_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_9_1_y0 = f_u_dadda_pg_rca16_and_9_1_a_9 & f_u_dadda_pg_rca16_and_9_1_b_1;
  assign f_u_dadda_pg_rca16_and_8_2_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_8_2_y0 = f_u_dadda_pg_rca16_and_8_2_a_8 & f_u_dadda_pg_rca16_and_8_2_b_2;
  assign f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_10_0_y0 = f_u_dadda_pg_rca16_and_10_0_y0;
  assign f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_9_1_y0 = f_u_dadda_pg_rca16_and_9_1_y0;
  assign f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_8_2_y0 = f_u_dadda_pg_rca16_and_8_2_y0;
  assign f_u_dadda_pg_rca16_fa25_y0 = f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_10_0_y0 ^ f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_9_1_y0;
  assign f_u_dadda_pg_rca16_fa25_y1 = f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_10_0_y0 & f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_9_1_y0;
  assign f_u_dadda_pg_rca16_fa25_y2 = f_u_dadda_pg_rca16_fa25_y0 ^ f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_8_2_y0;
  assign f_u_dadda_pg_rca16_fa25_y3 = f_u_dadda_pg_rca16_fa25_y0 & f_u_dadda_pg_rca16_fa25_f_u_dadda_pg_rca16_and_8_2_y0;
  assign f_u_dadda_pg_rca16_fa25_y4 = f_u_dadda_pg_rca16_fa25_y1 | f_u_dadda_pg_rca16_fa25_y3;
  assign f_u_dadda_pg_rca16_and_7_3_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_7_3_y0 = f_u_dadda_pg_rca16_and_7_3_a_7 & f_u_dadda_pg_rca16_and_7_3_b_3;
  assign f_u_dadda_pg_rca16_and_6_4_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_6_4_y0 = f_u_dadda_pg_rca16_and_6_4_a_6 & f_u_dadda_pg_rca16_and_6_4_b_4;
  assign f_u_dadda_pg_rca16_and_5_5_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_5_5_y0 = f_u_dadda_pg_rca16_and_5_5_a_5 & f_u_dadda_pg_rca16_and_5_5_b_5;
  assign f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_7_3_y0 = f_u_dadda_pg_rca16_and_7_3_y0;
  assign f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_6_4_y0 = f_u_dadda_pg_rca16_and_6_4_y0;
  assign f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_5_5_y0 = f_u_dadda_pg_rca16_and_5_5_y0;
  assign f_u_dadda_pg_rca16_fa26_y0 = f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_7_3_y0 ^ f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_6_4_y0;
  assign f_u_dadda_pg_rca16_fa26_y1 = f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_7_3_y0 & f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_6_4_y0;
  assign f_u_dadda_pg_rca16_fa26_y2 = f_u_dadda_pg_rca16_fa26_y0 ^ f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_5_5_y0;
  assign f_u_dadda_pg_rca16_fa26_y3 = f_u_dadda_pg_rca16_fa26_y0 & f_u_dadda_pg_rca16_fa26_f_u_dadda_pg_rca16_and_5_5_y0;
  assign f_u_dadda_pg_rca16_fa26_y4 = f_u_dadda_pg_rca16_fa26_y1 | f_u_dadda_pg_rca16_fa26_y3;
  assign f_u_dadda_pg_rca16_and_4_6_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_4_6_y0 = f_u_dadda_pg_rca16_and_4_6_a_4 & f_u_dadda_pg_rca16_and_4_6_b_6;
  assign f_u_dadda_pg_rca16_and_3_7_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_3_7_y0 = f_u_dadda_pg_rca16_and_3_7_a_3 & f_u_dadda_pg_rca16_and_3_7_b_7;
  assign f_u_dadda_pg_rca16_and_2_8_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_2_8_y0 = f_u_dadda_pg_rca16_and_2_8_a_2 & f_u_dadda_pg_rca16_and_2_8_b_8;
  assign f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_4_6_y0 = f_u_dadda_pg_rca16_and_4_6_y0;
  assign f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_3_7_y0 = f_u_dadda_pg_rca16_and_3_7_y0;
  assign f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_2_8_y0 = f_u_dadda_pg_rca16_and_2_8_y0;
  assign f_u_dadda_pg_rca16_fa27_y0 = f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_4_6_y0 ^ f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_3_7_y0;
  assign f_u_dadda_pg_rca16_fa27_y1 = f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_4_6_y0 & f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_3_7_y0;
  assign f_u_dadda_pg_rca16_fa27_y2 = f_u_dadda_pg_rca16_fa27_y0 ^ f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_2_8_y0;
  assign f_u_dadda_pg_rca16_fa27_y3 = f_u_dadda_pg_rca16_fa27_y0 & f_u_dadda_pg_rca16_fa27_f_u_dadda_pg_rca16_and_2_8_y0;
  assign f_u_dadda_pg_rca16_fa27_y4 = f_u_dadda_pg_rca16_fa27_y1 | f_u_dadda_pg_rca16_fa27_y3;
  assign f_u_dadda_pg_rca16_and_1_9_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_1_9_y0 = f_u_dadda_pg_rca16_and_1_9_a_1 & f_u_dadda_pg_rca16_and_1_9_b_9;
  assign f_u_dadda_pg_rca16_and_0_10_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_0_10_y0 = f_u_dadda_pg_rca16_and_0_10_a_0 & f_u_dadda_pg_rca16_and_0_10_b_10;
  assign f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_and_1_9_y0 = f_u_dadda_pg_rca16_and_1_9_y0;
  assign f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_and_0_10_y0 = f_u_dadda_pg_rca16_and_0_10_y0;
  assign f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_fa23_y2 = f_u_dadda_pg_rca16_fa23_y2;
  assign f_u_dadda_pg_rca16_fa28_y0 = f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_and_1_9_y0 ^ f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_and_0_10_y0;
  assign f_u_dadda_pg_rca16_fa28_y1 = f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_and_1_9_y0 & f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_and_0_10_y0;
  assign f_u_dadda_pg_rca16_fa28_y2 = f_u_dadda_pg_rca16_fa28_y0 ^ f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_fa23_y2;
  assign f_u_dadda_pg_rca16_fa28_y3 = f_u_dadda_pg_rca16_fa28_y0 & f_u_dadda_pg_rca16_fa28_f_u_dadda_pg_rca16_fa23_y2;
  assign f_u_dadda_pg_rca16_fa28_y4 = f_u_dadda_pg_rca16_fa28_y1 | f_u_dadda_pg_rca16_fa28_y3;
  assign f_u_dadda_pg_rca16_ha10_f_u_dadda_pg_rca16_fa24_y2 = f_u_dadda_pg_rca16_fa24_y2;
  assign f_u_dadda_pg_rca16_ha10_f_u_dadda_pg_rca16_fa25_y2 = f_u_dadda_pg_rca16_fa25_y2;
  assign f_u_dadda_pg_rca16_ha10_y0 = f_u_dadda_pg_rca16_ha10_f_u_dadda_pg_rca16_fa24_y2 ^ f_u_dadda_pg_rca16_ha10_f_u_dadda_pg_rca16_fa25_y2;
  assign f_u_dadda_pg_rca16_ha10_y1 = f_u_dadda_pg_rca16_ha10_f_u_dadda_pg_rca16_fa24_y2 & f_u_dadda_pg_rca16_ha10_f_u_dadda_pg_rca16_fa25_y2;
  assign f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_ha10_y1 = f_u_dadda_pg_rca16_ha10_y1;
  assign f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_fa28_y4 = f_u_dadda_pg_rca16_fa28_y4;
  assign f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_fa27_y4 = f_u_dadda_pg_rca16_fa27_y4;
  assign f_u_dadda_pg_rca16_fa29_y0 = f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_ha10_y1 ^ f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_fa28_y4;
  assign f_u_dadda_pg_rca16_fa29_y1 = f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_ha10_y1 & f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_fa28_y4;
  assign f_u_dadda_pg_rca16_fa29_y2 = f_u_dadda_pg_rca16_fa29_y0 ^ f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_fa27_y4;
  assign f_u_dadda_pg_rca16_fa29_y3 = f_u_dadda_pg_rca16_fa29_y0 & f_u_dadda_pg_rca16_fa29_f_u_dadda_pg_rca16_fa27_y4;
  assign f_u_dadda_pg_rca16_fa29_y4 = f_u_dadda_pg_rca16_fa29_y1 | f_u_dadda_pg_rca16_fa29_y3;
  assign f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa26_y4 = f_u_dadda_pg_rca16_fa26_y4;
  assign f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa25_y4 = f_u_dadda_pg_rca16_fa25_y4;
  assign f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa24_y4 = f_u_dadda_pg_rca16_fa24_y4;
  assign f_u_dadda_pg_rca16_fa30_y0 = f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa26_y4 ^ f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa25_y4;
  assign f_u_dadda_pg_rca16_fa30_y1 = f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa26_y4 & f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa25_y4;
  assign f_u_dadda_pg_rca16_fa30_y2 = f_u_dadda_pg_rca16_fa30_y0 ^ f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa24_y4;
  assign f_u_dadda_pg_rca16_fa30_y3 = f_u_dadda_pg_rca16_fa30_y0 & f_u_dadda_pg_rca16_fa30_f_u_dadda_pg_rca16_fa24_y4;
  assign f_u_dadda_pg_rca16_fa30_y4 = f_u_dadda_pg_rca16_fa30_y1 | f_u_dadda_pg_rca16_fa30_y3;
  assign f_u_dadda_pg_rca16_and_11_0_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_11_0_y0 = f_u_dadda_pg_rca16_and_11_0_a_11 & f_u_dadda_pg_rca16_and_11_0_b_0;
  assign f_u_dadda_pg_rca16_and_10_1_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_10_1_y0 = f_u_dadda_pg_rca16_and_10_1_a_10 & f_u_dadda_pg_rca16_and_10_1_b_1;
  assign f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_fa23_y4 = f_u_dadda_pg_rca16_fa23_y4;
  assign f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_and_11_0_y0 = f_u_dadda_pg_rca16_and_11_0_y0;
  assign f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_and_10_1_y0 = f_u_dadda_pg_rca16_and_10_1_y0;
  assign f_u_dadda_pg_rca16_fa31_y0 = f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_fa23_y4 ^ f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_and_11_0_y0;
  assign f_u_dadda_pg_rca16_fa31_y1 = f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_fa23_y4 & f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_and_11_0_y0;
  assign f_u_dadda_pg_rca16_fa31_y2 = f_u_dadda_pg_rca16_fa31_y0 ^ f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_and_10_1_y0;
  assign f_u_dadda_pg_rca16_fa31_y3 = f_u_dadda_pg_rca16_fa31_y0 & f_u_dadda_pg_rca16_fa31_f_u_dadda_pg_rca16_and_10_1_y0;
  assign f_u_dadda_pg_rca16_fa31_y4 = f_u_dadda_pg_rca16_fa31_y1 | f_u_dadda_pg_rca16_fa31_y3;
  assign f_u_dadda_pg_rca16_and_9_2_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_9_2_y0 = f_u_dadda_pg_rca16_and_9_2_a_9 & f_u_dadda_pg_rca16_and_9_2_b_2;
  assign f_u_dadda_pg_rca16_and_8_3_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_8_3_y0 = f_u_dadda_pg_rca16_and_8_3_a_8 & f_u_dadda_pg_rca16_and_8_3_b_3;
  assign f_u_dadda_pg_rca16_and_7_4_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_7_4_y0 = f_u_dadda_pg_rca16_and_7_4_a_7 & f_u_dadda_pg_rca16_and_7_4_b_4;
  assign f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_9_2_y0 = f_u_dadda_pg_rca16_and_9_2_y0;
  assign f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_8_3_y0 = f_u_dadda_pg_rca16_and_8_3_y0;
  assign f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_7_4_y0 = f_u_dadda_pg_rca16_and_7_4_y0;
  assign f_u_dadda_pg_rca16_fa32_y0 = f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_9_2_y0 ^ f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_8_3_y0;
  assign f_u_dadda_pg_rca16_fa32_y1 = f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_9_2_y0 & f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_8_3_y0;
  assign f_u_dadda_pg_rca16_fa32_y2 = f_u_dadda_pg_rca16_fa32_y0 ^ f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_7_4_y0;
  assign f_u_dadda_pg_rca16_fa32_y3 = f_u_dadda_pg_rca16_fa32_y0 & f_u_dadda_pg_rca16_fa32_f_u_dadda_pg_rca16_and_7_4_y0;
  assign f_u_dadda_pg_rca16_fa32_y4 = f_u_dadda_pg_rca16_fa32_y1 | f_u_dadda_pg_rca16_fa32_y3;
  assign f_u_dadda_pg_rca16_and_6_5_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_6_5_y0 = f_u_dadda_pg_rca16_and_6_5_a_6 & f_u_dadda_pg_rca16_and_6_5_b_5;
  assign f_u_dadda_pg_rca16_and_5_6_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_5_6_y0 = f_u_dadda_pg_rca16_and_5_6_a_5 & f_u_dadda_pg_rca16_and_5_6_b_6;
  assign f_u_dadda_pg_rca16_and_4_7_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_4_7_y0 = f_u_dadda_pg_rca16_and_4_7_a_4 & f_u_dadda_pg_rca16_and_4_7_b_7;
  assign f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_6_5_y0 = f_u_dadda_pg_rca16_and_6_5_y0;
  assign f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_5_6_y0 = f_u_dadda_pg_rca16_and_5_6_y0;
  assign f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_4_7_y0 = f_u_dadda_pg_rca16_and_4_7_y0;
  assign f_u_dadda_pg_rca16_fa33_y0 = f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_6_5_y0 ^ f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_5_6_y0;
  assign f_u_dadda_pg_rca16_fa33_y1 = f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_6_5_y0 & f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_5_6_y0;
  assign f_u_dadda_pg_rca16_fa33_y2 = f_u_dadda_pg_rca16_fa33_y0 ^ f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_4_7_y0;
  assign f_u_dadda_pg_rca16_fa33_y3 = f_u_dadda_pg_rca16_fa33_y0 & f_u_dadda_pg_rca16_fa33_f_u_dadda_pg_rca16_and_4_7_y0;
  assign f_u_dadda_pg_rca16_fa33_y4 = f_u_dadda_pg_rca16_fa33_y1 | f_u_dadda_pg_rca16_fa33_y3;
  assign f_u_dadda_pg_rca16_and_3_8_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_3_8_y0 = f_u_dadda_pg_rca16_and_3_8_a_3 & f_u_dadda_pg_rca16_and_3_8_b_8;
  assign f_u_dadda_pg_rca16_and_2_9_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_2_9_y0 = f_u_dadda_pg_rca16_and_2_9_a_2 & f_u_dadda_pg_rca16_and_2_9_b_9;
  assign f_u_dadda_pg_rca16_and_1_10_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_1_10_y0 = f_u_dadda_pg_rca16_and_1_10_a_1 & f_u_dadda_pg_rca16_and_1_10_b_10;
  assign f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_3_8_y0 = f_u_dadda_pg_rca16_and_3_8_y0;
  assign f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_2_9_y0 = f_u_dadda_pg_rca16_and_2_9_y0;
  assign f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_1_10_y0 = f_u_dadda_pg_rca16_and_1_10_y0;
  assign f_u_dadda_pg_rca16_fa34_y0 = f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_3_8_y0 ^ f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_2_9_y0;
  assign f_u_dadda_pg_rca16_fa34_y1 = f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_3_8_y0 & f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_2_9_y0;
  assign f_u_dadda_pg_rca16_fa34_y2 = f_u_dadda_pg_rca16_fa34_y0 ^ f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_1_10_y0;
  assign f_u_dadda_pg_rca16_fa34_y3 = f_u_dadda_pg_rca16_fa34_y0 & f_u_dadda_pg_rca16_fa34_f_u_dadda_pg_rca16_and_1_10_y0;
  assign f_u_dadda_pg_rca16_fa34_y4 = f_u_dadda_pg_rca16_fa34_y1 | f_u_dadda_pg_rca16_fa34_y3;
  assign f_u_dadda_pg_rca16_and_0_11_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_0_11_y0 = f_u_dadda_pg_rca16_and_0_11_a_0 & f_u_dadda_pg_rca16_and_0_11_b_11;
  assign f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_and_0_11_y0 = f_u_dadda_pg_rca16_and_0_11_y0;
  assign f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_fa29_y2 = f_u_dadda_pg_rca16_fa29_y2;
  assign f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_fa30_y2 = f_u_dadda_pg_rca16_fa30_y2;
  assign f_u_dadda_pg_rca16_fa35_y0 = f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_and_0_11_y0 ^ f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_fa29_y2;
  assign f_u_dadda_pg_rca16_fa35_y1 = f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_and_0_11_y0 & f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_fa29_y2;
  assign f_u_dadda_pg_rca16_fa35_y2 = f_u_dadda_pg_rca16_fa35_y0 ^ f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_fa30_y2;
  assign f_u_dadda_pg_rca16_fa35_y3 = f_u_dadda_pg_rca16_fa35_y0 & f_u_dadda_pg_rca16_fa35_f_u_dadda_pg_rca16_fa30_y2;
  assign f_u_dadda_pg_rca16_fa35_y4 = f_u_dadda_pg_rca16_fa35_y1 | f_u_dadda_pg_rca16_fa35_y3;
  assign f_u_dadda_pg_rca16_ha11_f_u_dadda_pg_rca16_fa31_y2 = f_u_dadda_pg_rca16_fa31_y2;
  assign f_u_dadda_pg_rca16_ha11_f_u_dadda_pg_rca16_fa32_y2 = f_u_dadda_pg_rca16_fa32_y2;
  assign f_u_dadda_pg_rca16_ha11_y0 = f_u_dadda_pg_rca16_ha11_f_u_dadda_pg_rca16_fa31_y2 ^ f_u_dadda_pg_rca16_ha11_f_u_dadda_pg_rca16_fa32_y2;
  assign f_u_dadda_pg_rca16_ha11_y1 = f_u_dadda_pg_rca16_ha11_f_u_dadda_pg_rca16_fa31_y2 & f_u_dadda_pg_rca16_ha11_f_u_dadda_pg_rca16_fa32_y2;
  assign f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_ha11_y1 = f_u_dadda_pg_rca16_ha11_y1;
  assign f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_fa35_y4 = f_u_dadda_pg_rca16_fa35_y4;
  assign f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_fa34_y4 = f_u_dadda_pg_rca16_fa34_y4;
  assign f_u_dadda_pg_rca16_fa36_y0 = f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_ha11_y1 ^ f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_fa35_y4;
  assign f_u_dadda_pg_rca16_fa36_y1 = f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_ha11_y1 & f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_fa35_y4;
  assign f_u_dadda_pg_rca16_fa36_y2 = f_u_dadda_pg_rca16_fa36_y0 ^ f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_fa34_y4;
  assign f_u_dadda_pg_rca16_fa36_y3 = f_u_dadda_pg_rca16_fa36_y0 & f_u_dadda_pg_rca16_fa36_f_u_dadda_pg_rca16_fa34_y4;
  assign f_u_dadda_pg_rca16_fa36_y4 = f_u_dadda_pg_rca16_fa36_y1 | f_u_dadda_pg_rca16_fa36_y3;
  assign f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa33_y4 = f_u_dadda_pg_rca16_fa33_y4;
  assign f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa32_y4 = f_u_dadda_pg_rca16_fa32_y4;
  assign f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa31_y4 = f_u_dadda_pg_rca16_fa31_y4;
  assign f_u_dadda_pg_rca16_fa37_y0 = f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa33_y4 ^ f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa32_y4;
  assign f_u_dadda_pg_rca16_fa37_y1 = f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa33_y4 & f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa32_y4;
  assign f_u_dadda_pg_rca16_fa37_y2 = f_u_dadda_pg_rca16_fa37_y0 ^ f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa31_y4;
  assign f_u_dadda_pg_rca16_fa37_y3 = f_u_dadda_pg_rca16_fa37_y0 & f_u_dadda_pg_rca16_fa37_f_u_dadda_pg_rca16_fa31_y4;
  assign f_u_dadda_pg_rca16_fa37_y4 = f_u_dadda_pg_rca16_fa37_y1 | f_u_dadda_pg_rca16_fa37_y3;
  assign f_u_dadda_pg_rca16_and_12_0_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_12_0_y0 = f_u_dadda_pg_rca16_and_12_0_a_12 & f_u_dadda_pg_rca16_and_12_0_b_0;
  assign f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_fa30_y4 = f_u_dadda_pg_rca16_fa30_y4;
  assign f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_fa29_y4 = f_u_dadda_pg_rca16_fa29_y4;
  assign f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_and_12_0_y0 = f_u_dadda_pg_rca16_and_12_0_y0;
  assign f_u_dadda_pg_rca16_fa38_y0 = f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_fa30_y4 ^ f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_fa29_y4;
  assign f_u_dadda_pg_rca16_fa38_y1 = f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_fa30_y4 & f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_fa29_y4;
  assign f_u_dadda_pg_rca16_fa38_y2 = f_u_dadda_pg_rca16_fa38_y0 ^ f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_and_12_0_y0;
  assign f_u_dadda_pg_rca16_fa38_y3 = f_u_dadda_pg_rca16_fa38_y0 & f_u_dadda_pg_rca16_fa38_f_u_dadda_pg_rca16_and_12_0_y0;
  assign f_u_dadda_pg_rca16_fa38_y4 = f_u_dadda_pg_rca16_fa38_y1 | f_u_dadda_pg_rca16_fa38_y3;
  assign f_u_dadda_pg_rca16_and_11_1_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_11_1_y0 = f_u_dadda_pg_rca16_and_11_1_a_11 & f_u_dadda_pg_rca16_and_11_1_b_1;
  assign f_u_dadda_pg_rca16_and_10_2_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_10_2_y0 = f_u_dadda_pg_rca16_and_10_2_a_10 & f_u_dadda_pg_rca16_and_10_2_b_2;
  assign f_u_dadda_pg_rca16_and_9_3_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_9_3_y0 = f_u_dadda_pg_rca16_and_9_3_a_9 & f_u_dadda_pg_rca16_and_9_3_b_3;
  assign f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_11_1_y0 = f_u_dadda_pg_rca16_and_11_1_y0;
  assign f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_10_2_y0 = f_u_dadda_pg_rca16_and_10_2_y0;
  assign f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_9_3_y0 = f_u_dadda_pg_rca16_and_9_3_y0;
  assign f_u_dadda_pg_rca16_fa39_y0 = f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_11_1_y0 ^ f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_10_2_y0;
  assign f_u_dadda_pg_rca16_fa39_y1 = f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_11_1_y0 & f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_10_2_y0;
  assign f_u_dadda_pg_rca16_fa39_y2 = f_u_dadda_pg_rca16_fa39_y0 ^ f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_9_3_y0;
  assign f_u_dadda_pg_rca16_fa39_y3 = f_u_dadda_pg_rca16_fa39_y0 & f_u_dadda_pg_rca16_fa39_f_u_dadda_pg_rca16_and_9_3_y0;
  assign f_u_dadda_pg_rca16_fa39_y4 = f_u_dadda_pg_rca16_fa39_y1 | f_u_dadda_pg_rca16_fa39_y3;
  assign f_u_dadda_pg_rca16_and_8_4_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_8_4_y0 = f_u_dadda_pg_rca16_and_8_4_a_8 & f_u_dadda_pg_rca16_and_8_4_b_4;
  assign f_u_dadda_pg_rca16_and_7_5_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_7_5_y0 = f_u_dadda_pg_rca16_and_7_5_a_7 & f_u_dadda_pg_rca16_and_7_5_b_5;
  assign f_u_dadda_pg_rca16_and_6_6_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_6_6_y0 = f_u_dadda_pg_rca16_and_6_6_a_6 & f_u_dadda_pg_rca16_and_6_6_b_6;
  assign f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_8_4_y0 = f_u_dadda_pg_rca16_and_8_4_y0;
  assign f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_7_5_y0 = f_u_dadda_pg_rca16_and_7_5_y0;
  assign f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_6_6_y0 = f_u_dadda_pg_rca16_and_6_6_y0;
  assign f_u_dadda_pg_rca16_fa40_y0 = f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_8_4_y0 ^ f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_7_5_y0;
  assign f_u_dadda_pg_rca16_fa40_y1 = f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_8_4_y0 & f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_7_5_y0;
  assign f_u_dadda_pg_rca16_fa40_y2 = f_u_dadda_pg_rca16_fa40_y0 ^ f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_6_6_y0;
  assign f_u_dadda_pg_rca16_fa40_y3 = f_u_dadda_pg_rca16_fa40_y0 & f_u_dadda_pg_rca16_fa40_f_u_dadda_pg_rca16_and_6_6_y0;
  assign f_u_dadda_pg_rca16_fa40_y4 = f_u_dadda_pg_rca16_fa40_y1 | f_u_dadda_pg_rca16_fa40_y3;
  assign f_u_dadda_pg_rca16_and_5_7_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_5_7_y0 = f_u_dadda_pg_rca16_and_5_7_a_5 & f_u_dadda_pg_rca16_and_5_7_b_7;
  assign f_u_dadda_pg_rca16_and_4_8_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_4_8_y0 = f_u_dadda_pg_rca16_and_4_8_a_4 & f_u_dadda_pg_rca16_and_4_8_b_8;
  assign f_u_dadda_pg_rca16_and_3_9_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_3_9_y0 = f_u_dadda_pg_rca16_and_3_9_a_3 & f_u_dadda_pg_rca16_and_3_9_b_9;
  assign f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_5_7_y0 = f_u_dadda_pg_rca16_and_5_7_y0;
  assign f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_4_8_y0 = f_u_dadda_pg_rca16_and_4_8_y0;
  assign f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_3_9_y0 = f_u_dadda_pg_rca16_and_3_9_y0;
  assign f_u_dadda_pg_rca16_fa41_y0 = f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_5_7_y0 ^ f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_4_8_y0;
  assign f_u_dadda_pg_rca16_fa41_y1 = f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_5_7_y0 & f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_4_8_y0;
  assign f_u_dadda_pg_rca16_fa41_y2 = f_u_dadda_pg_rca16_fa41_y0 ^ f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_3_9_y0;
  assign f_u_dadda_pg_rca16_fa41_y3 = f_u_dadda_pg_rca16_fa41_y0 & f_u_dadda_pg_rca16_fa41_f_u_dadda_pg_rca16_and_3_9_y0;
  assign f_u_dadda_pg_rca16_fa41_y4 = f_u_dadda_pg_rca16_fa41_y1 | f_u_dadda_pg_rca16_fa41_y3;
  assign f_u_dadda_pg_rca16_and_2_10_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_2_10_y0 = f_u_dadda_pg_rca16_and_2_10_a_2 & f_u_dadda_pg_rca16_and_2_10_b_10;
  assign f_u_dadda_pg_rca16_and_1_11_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_1_11_y0 = f_u_dadda_pg_rca16_and_1_11_a_1 & f_u_dadda_pg_rca16_and_1_11_b_11;
  assign f_u_dadda_pg_rca16_and_0_12_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_0_12_y0 = f_u_dadda_pg_rca16_and_0_12_a_0 & f_u_dadda_pg_rca16_and_0_12_b_12;
  assign f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_2_10_y0 = f_u_dadda_pg_rca16_and_2_10_y0;
  assign f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_1_11_y0 = f_u_dadda_pg_rca16_and_1_11_y0;
  assign f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_0_12_y0 = f_u_dadda_pg_rca16_and_0_12_y0;
  assign f_u_dadda_pg_rca16_fa42_y0 = f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_2_10_y0 ^ f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_1_11_y0;
  assign f_u_dadda_pg_rca16_fa42_y1 = f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_2_10_y0 & f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_1_11_y0;
  assign f_u_dadda_pg_rca16_fa42_y2 = f_u_dadda_pg_rca16_fa42_y0 ^ f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_0_12_y0;
  assign f_u_dadda_pg_rca16_fa42_y3 = f_u_dadda_pg_rca16_fa42_y0 & f_u_dadda_pg_rca16_fa42_f_u_dadda_pg_rca16_and_0_12_y0;
  assign f_u_dadda_pg_rca16_fa42_y4 = f_u_dadda_pg_rca16_fa42_y1 | f_u_dadda_pg_rca16_fa42_y3;
  assign f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa36_y2 = f_u_dadda_pg_rca16_fa36_y2;
  assign f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa37_y2 = f_u_dadda_pg_rca16_fa37_y2;
  assign f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa38_y2 = f_u_dadda_pg_rca16_fa38_y2;
  assign f_u_dadda_pg_rca16_fa43_y0 = f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa36_y2 ^ f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa37_y2;
  assign f_u_dadda_pg_rca16_fa43_y1 = f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa36_y2 & f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa37_y2;
  assign f_u_dadda_pg_rca16_fa43_y2 = f_u_dadda_pg_rca16_fa43_y0 ^ f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa38_y2;
  assign f_u_dadda_pg_rca16_fa43_y3 = f_u_dadda_pg_rca16_fa43_y0 & f_u_dadda_pg_rca16_fa43_f_u_dadda_pg_rca16_fa38_y2;
  assign f_u_dadda_pg_rca16_fa43_y4 = f_u_dadda_pg_rca16_fa43_y1 | f_u_dadda_pg_rca16_fa43_y3;
  assign f_u_dadda_pg_rca16_ha12_f_u_dadda_pg_rca16_fa39_y2 = f_u_dadda_pg_rca16_fa39_y2;
  assign f_u_dadda_pg_rca16_ha12_f_u_dadda_pg_rca16_fa40_y2 = f_u_dadda_pg_rca16_fa40_y2;
  assign f_u_dadda_pg_rca16_ha12_y0 = f_u_dadda_pg_rca16_ha12_f_u_dadda_pg_rca16_fa39_y2 ^ f_u_dadda_pg_rca16_ha12_f_u_dadda_pg_rca16_fa40_y2;
  assign f_u_dadda_pg_rca16_ha12_y1 = f_u_dadda_pg_rca16_ha12_f_u_dadda_pg_rca16_fa39_y2 & f_u_dadda_pg_rca16_ha12_f_u_dadda_pg_rca16_fa40_y2;
  assign f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_ha12_y1 = f_u_dadda_pg_rca16_ha12_y1;
  assign f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_fa43_y4 = f_u_dadda_pg_rca16_fa43_y4;
  assign f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_fa42_y4 = f_u_dadda_pg_rca16_fa42_y4;
  assign f_u_dadda_pg_rca16_fa44_y0 = f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_ha12_y1 ^ f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_fa43_y4;
  assign f_u_dadda_pg_rca16_fa44_y1 = f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_ha12_y1 & f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_fa43_y4;
  assign f_u_dadda_pg_rca16_fa44_y2 = f_u_dadda_pg_rca16_fa44_y0 ^ f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_fa42_y4;
  assign f_u_dadda_pg_rca16_fa44_y3 = f_u_dadda_pg_rca16_fa44_y0 & f_u_dadda_pg_rca16_fa44_f_u_dadda_pg_rca16_fa42_y4;
  assign f_u_dadda_pg_rca16_fa44_y4 = f_u_dadda_pg_rca16_fa44_y1 | f_u_dadda_pg_rca16_fa44_y3;
  assign f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa41_y4 = f_u_dadda_pg_rca16_fa41_y4;
  assign f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa40_y4 = f_u_dadda_pg_rca16_fa40_y4;
  assign f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa39_y4 = f_u_dadda_pg_rca16_fa39_y4;
  assign f_u_dadda_pg_rca16_fa45_y0 = f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa41_y4 ^ f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa40_y4;
  assign f_u_dadda_pg_rca16_fa45_y1 = f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa41_y4 & f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa40_y4;
  assign f_u_dadda_pg_rca16_fa45_y2 = f_u_dadda_pg_rca16_fa45_y0 ^ f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa39_y4;
  assign f_u_dadda_pg_rca16_fa45_y3 = f_u_dadda_pg_rca16_fa45_y0 & f_u_dadda_pg_rca16_fa45_f_u_dadda_pg_rca16_fa39_y4;
  assign f_u_dadda_pg_rca16_fa45_y4 = f_u_dadda_pg_rca16_fa45_y1 | f_u_dadda_pg_rca16_fa45_y3;
  assign f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa38_y4 = f_u_dadda_pg_rca16_fa38_y4;
  assign f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa37_y4 = f_u_dadda_pg_rca16_fa37_y4;
  assign f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa36_y4 = f_u_dadda_pg_rca16_fa36_y4;
  assign f_u_dadda_pg_rca16_fa46_y0 = f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa38_y4 ^ f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa37_y4;
  assign f_u_dadda_pg_rca16_fa46_y1 = f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa38_y4 & f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa37_y4;
  assign f_u_dadda_pg_rca16_fa46_y2 = f_u_dadda_pg_rca16_fa46_y0 ^ f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa36_y4;
  assign f_u_dadda_pg_rca16_fa46_y3 = f_u_dadda_pg_rca16_fa46_y0 & f_u_dadda_pg_rca16_fa46_f_u_dadda_pg_rca16_fa36_y4;
  assign f_u_dadda_pg_rca16_fa46_y4 = f_u_dadda_pg_rca16_fa46_y1 | f_u_dadda_pg_rca16_fa46_y3;
  assign f_u_dadda_pg_rca16_and_11_2_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_11_2_y0 = f_u_dadda_pg_rca16_and_11_2_a_11 & f_u_dadda_pg_rca16_and_11_2_b_2;
  assign f_u_dadda_pg_rca16_and_10_3_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_10_3_y0 = f_u_dadda_pg_rca16_and_10_3_a_10 & f_u_dadda_pg_rca16_and_10_3_b_3;
  assign f_u_dadda_pg_rca16_and_9_4_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_9_4_y0 = f_u_dadda_pg_rca16_and_9_4_a_9 & f_u_dadda_pg_rca16_and_9_4_b_4;
  assign f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_11_2_y0 = f_u_dadda_pg_rca16_and_11_2_y0;
  assign f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_10_3_y0 = f_u_dadda_pg_rca16_and_10_3_y0;
  assign f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_9_4_y0 = f_u_dadda_pg_rca16_and_9_4_y0;
  assign f_u_dadda_pg_rca16_fa47_y0 = f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_11_2_y0 ^ f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_10_3_y0;
  assign f_u_dadda_pg_rca16_fa47_y1 = f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_11_2_y0 & f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_10_3_y0;
  assign f_u_dadda_pg_rca16_fa47_y2 = f_u_dadda_pg_rca16_fa47_y0 ^ f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_9_4_y0;
  assign f_u_dadda_pg_rca16_fa47_y3 = f_u_dadda_pg_rca16_fa47_y0 & f_u_dadda_pg_rca16_fa47_f_u_dadda_pg_rca16_and_9_4_y0;
  assign f_u_dadda_pg_rca16_fa47_y4 = f_u_dadda_pg_rca16_fa47_y1 | f_u_dadda_pg_rca16_fa47_y3;
  assign f_u_dadda_pg_rca16_and_8_5_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_8_5_y0 = f_u_dadda_pg_rca16_and_8_5_a_8 & f_u_dadda_pg_rca16_and_8_5_b_5;
  assign f_u_dadda_pg_rca16_and_7_6_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_7_6_y0 = f_u_dadda_pg_rca16_and_7_6_a_7 & f_u_dadda_pg_rca16_and_7_6_b_6;
  assign f_u_dadda_pg_rca16_and_6_7_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_6_7_y0 = f_u_dadda_pg_rca16_and_6_7_a_6 & f_u_dadda_pg_rca16_and_6_7_b_7;
  assign f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_8_5_y0 = f_u_dadda_pg_rca16_and_8_5_y0;
  assign f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_7_6_y0 = f_u_dadda_pg_rca16_and_7_6_y0;
  assign f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_6_7_y0 = f_u_dadda_pg_rca16_and_6_7_y0;
  assign f_u_dadda_pg_rca16_fa48_y0 = f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_8_5_y0 ^ f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_7_6_y0;
  assign f_u_dadda_pg_rca16_fa48_y1 = f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_8_5_y0 & f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_7_6_y0;
  assign f_u_dadda_pg_rca16_fa48_y2 = f_u_dadda_pg_rca16_fa48_y0 ^ f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_6_7_y0;
  assign f_u_dadda_pg_rca16_fa48_y3 = f_u_dadda_pg_rca16_fa48_y0 & f_u_dadda_pg_rca16_fa48_f_u_dadda_pg_rca16_and_6_7_y0;
  assign f_u_dadda_pg_rca16_fa48_y4 = f_u_dadda_pg_rca16_fa48_y1 | f_u_dadda_pg_rca16_fa48_y3;
  assign f_u_dadda_pg_rca16_and_5_8_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_5_8_y0 = f_u_dadda_pg_rca16_and_5_8_a_5 & f_u_dadda_pg_rca16_and_5_8_b_8;
  assign f_u_dadda_pg_rca16_and_4_9_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_4_9_y0 = f_u_dadda_pg_rca16_and_4_9_a_4 & f_u_dadda_pg_rca16_and_4_9_b_9;
  assign f_u_dadda_pg_rca16_and_3_10_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_3_10_y0 = f_u_dadda_pg_rca16_and_3_10_a_3 & f_u_dadda_pg_rca16_and_3_10_b_10;
  assign f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_5_8_y0 = f_u_dadda_pg_rca16_and_5_8_y0;
  assign f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_4_9_y0 = f_u_dadda_pg_rca16_and_4_9_y0;
  assign f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_3_10_y0 = f_u_dadda_pg_rca16_and_3_10_y0;
  assign f_u_dadda_pg_rca16_fa49_y0 = f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_5_8_y0 ^ f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_4_9_y0;
  assign f_u_dadda_pg_rca16_fa49_y1 = f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_5_8_y0 & f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_4_9_y0;
  assign f_u_dadda_pg_rca16_fa49_y2 = f_u_dadda_pg_rca16_fa49_y0 ^ f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_3_10_y0;
  assign f_u_dadda_pg_rca16_fa49_y3 = f_u_dadda_pg_rca16_fa49_y0 & f_u_dadda_pg_rca16_fa49_f_u_dadda_pg_rca16_and_3_10_y0;
  assign f_u_dadda_pg_rca16_fa49_y4 = f_u_dadda_pg_rca16_fa49_y1 | f_u_dadda_pg_rca16_fa49_y3;
  assign f_u_dadda_pg_rca16_and_2_11_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_2_11_y0 = f_u_dadda_pg_rca16_and_2_11_a_2 & f_u_dadda_pg_rca16_and_2_11_b_11;
  assign f_u_dadda_pg_rca16_and_1_12_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_1_12_y0 = f_u_dadda_pg_rca16_and_1_12_a_1 & f_u_dadda_pg_rca16_and_1_12_b_12;
  assign f_u_dadda_pg_rca16_and_0_13_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_0_13_y0 = f_u_dadda_pg_rca16_and_0_13_a_0 & f_u_dadda_pg_rca16_and_0_13_b_13;
  assign f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_2_11_y0 = f_u_dadda_pg_rca16_and_2_11_y0;
  assign f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_1_12_y0 = f_u_dadda_pg_rca16_and_1_12_y0;
  assign f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_0_13_y0 = f_u_dadda_pg_rca16_and_0_13_y0;
  assign f_u_dadda_pg_rca16_fa50_y0 = f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_2_11_y0 ^ f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_1_12_y0;
  assign f_u_dadda_pg_rca16_fa50_y1 = f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_2_11_y0 & f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_1_12_y0;
  assign f_u_dadda_pg_rca16_fa50_y2 = f_u_dadda_pg_rca16_fa50_y0 ^ f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_0_13_y0;
  assign f_u_dadda_pg_rca16_fa50_y3 = f_u_dadda_pg_rca16_fa50_y0 & f_u_dadda_pg_rca16_fa50_f_u_dadda_pg_rca16_and_0_13_y0;
  assign f_u_dadda_pg_rca16_fa50_y4 = f_u_dadda_pg_rca16_fa50_y1 | f_u_dadda_pg_rca16_fa50_y3;
  assign f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_ha0_y0 = f_u_dadda_pg_rca16_ha0_y0;
  assign f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_fa44_y2 = f_u_dadda_pg_rca16_fa44_y2;
  assign f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_fa45_y2 = f_u_dadda_pg_rca16_fa45_y2;
  assign f_u_dadda_pg_rca16_fa51_y0 = f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_ha0_y0 ^ f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_fa44_y2;
  assign f_u_dadda_pg_rca16_fa51_y1 = f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_ha0_y0 & f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_fa44_y2;
  assign f_u_dadda_pg_rca16_fa51_y2 = f_u_dadda_pg_rca16_fa51_y0 ^ f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_fa45_y2;
  assign f_u_dadda_pg_rca16_fa51_y3 = f_u_dadda_pg_rca16_fa51_y0 & f_u_dadda_pg_rca16_fa51_f_u_dadda_pg_rca16_fa45_y2;
  assign f_u_dadda_pg_rca16_fa51_y4 = f_u_dadda_pg_rca16_fa51_y1 | f_u_dadda_pg_rca16_fa51_y3;
  assign f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa46_y2 = f_u_dadda_pg_rca16_fa46_y2;
  assign f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa47_y2 = f_u_dadda_pg_rca16_fa47_y2;
  assign f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa48_y2 = f_u_dadda_pg_rca16_fa48_y2;
  assign f_u_dadda_pg_rca16_fa52_y0 = f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa46_y2 ^ f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa47_y2;
  assign f_u_dadda_pg_rca16_fa52_y1 = f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa46_y2 & f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa47_y2;
  assign f_u_dadda_pg_rca16_fa52_y2 = f_u_dadda_pg_rca16_fa52_y0 ^ f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa48_y2;
  assign f_u_dadda_pg_rca16_fa52_y3 = f_u_dadda_pg_rca16_fa52_y0 & f_u_dadda_pg_rca16_fa52_f_u_dadda_pg_rca16_fa48_y2;
  assign f_u_dadda_pg_rca16_fa52_y4 = f_u_dadda_pg_rca16_fa52_y1 | f_u_dadda_pg_rca16_fa52_y3;
  assign f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa52_y4 = f_u_dadda_pg_rca16_fa52_y4;
  assign f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa51_y4 = f_u_dadda_pg_rca16_fa51_y4;
  assign f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa50_y4 = f_u_dadda_pg_rca16_fa50_y4;
  assign f_u_dadda_pg_rca16_fa53_y0 = f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa52_y4 ^ f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa51_y4;
  assign f_u_dadda_pg_rca16_fa53_y1 = f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa52_y4 & f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa51_y4;
  assign f_u_dadda_pg_rca16_fa53_y2 = f_u_dadda_pg_rca16_fa53_y0 ^ f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa50_y4;
  assign f_u_dadda_pg_rca16_fa53_y3 = f_u_dadda_pg_rca16_fa53_y0 & f_u_dadda_pg_rca16_fa53_f_u_dadda_pg_rca16_fa50_y4;
  assign f_u_dadda_pg_rca16_fa53_y4 = f_u_dadda_pg_rca16_fa53_y1 | f_u_dadda_pg_rca16_fa53_y3;
  assign f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa49_y4 = f_u_dadda_pg_rca16_fa49_y4;
  assign f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa48_y4 = f_u_dadda_pg_rca16_fa48_y4;
  assign f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa47_y4 = f_u_dadda_pg_rca16_fa47_y4;
  assign f_u_dadda_pg_rca16_fa54_y0 = f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa49_y4 ^ f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa48_y4;
  assign f_u_dadda_pg_rca16_fa54_y1 = f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa49_y4 & f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa48_y4;
  assign f_u_dadda_pg_rca16_fa54_y2 = f_u_dadda_pg_rca16_fa54_y0 ^ f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa47_y4;
  assign f_u_dadda_pg_rca16_fa54_y3 = f_u_dadda_pg_rca16_fa54_y0 & f_u_dadda_pg_rca16_fa54_f_u_dadda_pg_rca16_fa47_y4;
  assign f_u_dadda_pg_rca16_fa54_y4 = f_u_dadda_pg_rca16_fa54_y1 | f_u_dadda_pg_rca16_fa54_y3;
  assign f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa46_y4 = f_u_dadda_pg_rca16_fa46_y4;
  assign f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa45_y4 = f_u_dadda_pg_rca16_fa45_y4;
  assign f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa44_y4 = f_u_dadda_pg_rca16_fa44_y4;
  assign f_u_dadda_pg_rca16_fa55_y0 = f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa46_y4 ^ f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa45_y4;
  assign f_u_dadda_pg_rca16_fa55_y1 = f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa46_y4 & f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa45_y4;
  assign f_u_dadda_pg_rca16_fa55_y2 = f_u_dadda_pg_rca16_fa55_y0 ^ f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa44_y4;
  assign f_u_dadda_pg_rca16_fa55_y3 = f_u_dadda_pg_rca16_fa55_y0 & f_u_dadda_pg_rca16_fa55_f_u_dadda_pg_rca16_fa44_y4;
  assign f_u_dadda_pg_rca16_fa55_y4 = f_u_dadda_pg_rca16_fa55_y1 | f_u_dadda_pg_rca16_fa55_y3;
  assign f_u_dadda_pg_rca16_and_10_4_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_10_4_y0 = f_u_dadda_pg_rca16_and_10_4_a_10 & f_u_dadda_pg_rca16_and_10_4_b_4;
  assign f_u_dadda_pg_rca16_and_9_5_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_9_5_y0 = f_u_dadda_pg_rca16_and_9_5_a_9 & f_u_dadda_pg_rca16_and_9_5_b_5;
  assign f_u_dadda_pg_rca16_and_8_6_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_8_6_y0 = f_u_dadda_pg_rca16_and_8_6_a_8 & f_u_dadda_pg_rca16_and_8_6_b_6;
  assign f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_10_4_y0 = f_u_dadda_pg_rca16_and_10_4_y0;
  assign f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_9_5_y0 = f_u_dadda_pg_rca16_and_9_5_y0;
  assign f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_8_6_y0 = f_u_dadda_pg_rca16_and_8_6_y0;
  assign f_u_dadda_pg_rca16_fa56_y0 = f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_10_4_y0 ^ f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_9_5_y0;
  assign f_u_dadda_pg_rca16_fa56_y1 = f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_10_4_y0 & f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_9_5_y0;
  assign f_u_dadda_pg_rca16_fa56_y2 = f_u_dadda_pg_rca16_fa56_y0 ^ f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_8_6_y0;
  assign f_u_dadda_pg_rca16_fa56_y3 = f_u_dadda_pg_rca16_fa56_y0 & f_u_dadda_pg_rca16_fa56_f_u_dadda_pg_rca16_and_8_6_y0;
  assign f_u_dadda_pg_rca16_fa56_y4 = f_u_dadda_pg_rca16_fa56_y1 | f_u_dadda_pg_rca16_fa56_y3;
  assign f_u_dadda_pg_rca16_and_7_7_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_7_7_y0 = f_u_dadda_pg_rca16_and_7_7_a_7 & f_u_dadda_pg_rca16_and_7_7_b_7;
  assign f_u_dadda_pg_rca16_and_6_8_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_6_8_y0 = f_u_dadda_pg_rca16_and_6_8_a_6 & f_u_dadda_pg_rca16_and_6_8_b_8;
  assign f_u_dadda_pg_rca16_and_5_9_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_5_9_y0 = f_u_dadda_pg_rca16_and_5_9_a_5 & f_u_dadda_pg_rca16_and_5_9_b_9;
  assign f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_7_7_y0 = f_u_dadda_pg_rca16_and_7_7_y0;
  assign f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_6_8_y0 = f_u_dadda_pg_rca16_and_6_8_y0;
  assign f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_5_9_y0 = f_u_dadda_pg_rca16_and_5_9_y0;
  assign f_u_dadda_pg_rca16_fa57_y0 = f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_7_7_y0 ^ f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_6_8_y0;
  assign f_u_dadda_pg_rca16_fa57_y1 = f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_7_7_y0 & f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_6_8_y0;
  assign f_u_dadda_pg_rca16_fa57_y2 = f_u_dadda_pg_rca16_fa57_y0 ^ f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_5_9_y0;
  assign f_u_dadda_pg_rca16_fa57_y3 = f_u_dadda_pg_rca16_fa57_y0 & f_u_dadda_pg_rca16_fa57_f_u_dadda_pg_rca16_and_5_9_y0;
  assign f_u_dadda_pg_rca16_fa57_y4 = f_u_dadda_pg_rca16_fa57_y1 | f_u_dadda_pg_rca16_fa57_y3;
  assign f_u_dadda_pg_rca16_and_4_10_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_4_10_y0 = f_u_dadda_pg_rca16_and_4_10_a_4 & f_u_dadda_pg_rca16_and_4_10_b_10;
  assign f_u_dadda_pg_rca16_and_3_11_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_3_11_y0 = f_u_dadda_pg_rca16_and_3_11_a_3 & f_u_dadda_pg_rca16_and_3_11_b_11;
  assign f_u_dadda_pg_rca16_and_2_12_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_2_12_y0 = f_u_dadda_pg_rca16_and_2_12_a_2 & f_u_dadda_pg_rca16_and_2_12_b_12;
  assign f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_4_10_y0 = f_u_dadda_pg_rca16_and_4_10_y0;
  assign f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_3_11_y0 = f_u_dadda_pg_rca16_and_3_11_y0;
  assign f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_2_12_y0 = f_u_dadda_pg_rca16_and_2_12_y0;
  assign f_u_dadda_pg_rca16_fa58_y0 = f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_4_10_y0 ^ f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_3_11_y0;
  assign f_u_dadda_pg_rca16_fa58_y1 = f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_4_10_y0 & f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_3_11_y0;
  assign f_u_dadda_pg_rca16_fa58_y2 = f_u_dadda_pg_rca16_fa58_y0 ^ f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_2_12_y0;
  assign f_u_dadda_pg_rca16_fa58_y3 = f_u_dadda_pg_rca16_fa58_y0 & f_u_dadda_pg_rca16_fa58_f_u_dadda_pg_rca16_and_2_12_y0;
  assign f_u_dadda_pg_rca16_fa58_y4 = f_u_dadda_pg_rca16_fa58_y1 | f_u_dadda_pg_rca16_fa58_y3;
  assign f_u_dadda_pg_rca16_and_1_13_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_1_13_y0 = f_u_dadda_pg_rca16_and_1_13_a_1 & f_u_dadda_pg_rca16_and_1_13_b_13;
  assign f_u_dadda_pg_rca16_and_0_14_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_0_14_y0 = f_u_dadda_pg_rca16_and_0_14_a_0 & f_u_dadda_pg_rca16_and_0_14_b_14;
  assign f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_and_1_13_y0 = f_u_dadda_pg_rca16_and_1_13_y0;
  assign f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_and_0_14_y0 = f_u_dadda_pg_rca16_and_0_14_y0;
  assign f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_fa0_y2 = f_u_dadda_pg_rca16_fa0_y2;
  assign f_u_dadda_pg_rca16_fa59_y0 = f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_and_1_13_y0 ^ f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_and_0_14_y0;
  assign f_u_dadda_pg_rca16_fa59_y1 = f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_and_1_13_y0 & f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_and_0_14_y0;
  assign f_u_dadda_pg_rca16_fa59_y2 = f_u_dadda_pg_rca16_fa59_y0 ^ f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_fa0_y2;
  assign f_u_dadda_pg_rca16_fa59_y3 = f_u_dadda_pg_rca16_fa59_y0 & f_u_dadda_pg_rca16_fa59_f_u_dadda_pg_rca16_fa0_y2;
  assign f_u_dadda_pg_rca16_fa59_y4 = f_u_dadda_pg_rca16_fa59_y1 | f_u_dadda_pg_rca16_fa59_y3;
  assign f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_ha1_y0 = f_u_dadda_pg_rca16_ha1_y0;
  assign f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_fa53_y2 = f_u_dadda_pg_rca16_fa53_y2;
  assign f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_fa54_y2 = f_u_dadda_pg_rca16_fa54_y2;
  assign f_u_dadda_pg_rca16_fa60_y0 = f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_ha1_y0 ^ f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_fa53_y2;
  assign f_u_dadda_pg_rca16_fa60_y1 = f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_ha1_y0 & f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_fa53_y2;
  assign f_u_dadda_pg_rca16_fa60_y2 = f_u_dadda_pg_rca16_fa60_y0 ^ f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_fa54_y2;
  assign f_u_dadda_pg_rca16_fa60_y3 = f_u_dadda_pg_rca16_fa60_y0 & f_u_dadda_pg_rca16_fa60_f_u_dadda_pg_rca16_fa54_y2;
  assign f_u_dadda_pg_rca16_fa60_y4 = f_u_dadda_pg_rca16_fa60_y1 | f_u_dadda_pg_rca16_fa60_y3;
  assign f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa55_y2 = f_u_dadda_pg_rca16_fa55_y2;
  assign f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa56_y2 = f_u_dadda_pg_rca16_fa56_y2;
  assign f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa57_y2 = f_u_dadda_pg_rca16_fa57_y2;
  assign f_u_dadda_pg_rca16_fa61_y0 = f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa55_y2 ^ f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa56_y2;
  assign f_u_dadda_pg_rca16_fa61_y1 = f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa55_y2 & f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa56_y2;
  assign f_u_dadda_pg_rca16_fa61_y2 = f_u_dadda_pg_rca16_fa61_y0 ^ f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa57_y2;
  assign f_u_dadda_pg_rca16_fa61_y3 = f_u_dadda_pg_rca16_fa61_y0 & f_u_dadda_pg_rca16_fa61_f_u_dadda_pg_rca16_fa57_y2;
  assign f_u_dadda_pg_rca16_fa61_y4 = f_u_dadda_pg_rca16_fa61_y1 | f_u_dadda_pg_rca16_fa61_y3;
  assign f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa61_y4 = f_u_dadda_pg_rca16_fa61_y4;
  assign f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa60_y4 = f_u_dadda_pg_rca16_fa60_y4;
  assign f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa59_y4 = f_u_dadda_pg_rca16_fa59_y4;
  assign f_u_dadda_pg_rca16_fa62_y0 = f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa61_y4 ^ f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa60_y4;
  assign f_u_dadda_pg_rca16_fa62_y1 = f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa61_y4 & f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa60_y4;
  assign f_u_dadda_pg_rca16_fa62_y2 = f_u_dadda_pg_rca16_fa62_y0 ^ f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa59_y4;
  assign f_u_dadda_pg_rca16_fa62_y3 = f_u_dadda_pg_rca16_fa62_y0 & f_u_dadda_pg_rca16_fa62_f_u_dadda_pg_rca16_fa59_y4;
  assign f_u_dadda_pg_rca16_fa62_y4 = f_u_dadda_pg_rca16_fa62_y1 | f_u_dadda_pg_rca16_fa62_y3;
  assign f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa58_y4 = f_u_dadda_pg_rca16_fa58_y4;
  assign f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa57_y4 = f_u_dadda_pg_rca16_fa57_y4;
  assign f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa56_y4 = f_u_dadda_pg_rca16_fa56_y4;
  assign f_u_dadda_pg_rca16_fa63_y0 = f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa58_y4 ^ f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa57_y4;
  assign f_u_dadda_pg_rca16_fa63_y1 = f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa58_y4 & f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa57_y4;
  assign f_u_dadda_pg_rca16_fa63_y2 = f_u_dadda_pg_rca16_fa63_y0 ^ f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa56_y4;
  assign f_u_dadda_pg_rca16_fa63_y3 = f_u_dadda_pg_rca16_fa63_y0 & f_u_dadda_pg_rca16_fa63_f_u_dadda_pg_rca16_fa56_y4;
  assign f_u_dadda_pg_rca16_fa63_y4 = f_u_dadda_pg_rca16_fa63_y1 | f_u_dadda_pg_rca16_fa63_y3;
  assign f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa55_y4 = f_u_dadda_pg_rca16_fa55_y4;
  assign f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa54_y4 = f_u_dadda_pg_rca16_fa54_y4;
  assign f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa53_y4 = f_u_dadda_pg_rca16_fa53_y4;
  assign f_u_dadda_pg_rca16_fa64_y0 = f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa55_y4 ^ f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa54_y4;
  assign f_u_dadda_pg_rca16_fa64_y1 = f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa55_y4 & f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa54_y4;
  assign f_u_dadda_pg_rca16_fa64_y2 = f_u_dadda_pg_rca16_fa64_y0 ^ f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa53_y4;
  assign f_u_dadda_pg_rca16_fa64_y3 = f_u_dadda_pg_rca16_fa64_y0 & f_u_dadda_pg_rca16_fa64_f_u_dadda_pg_rca16_fa53_y4;
  assign f_u_dadda_pg_rca16_fa64_y4 = f_u_dadda_pg_rca16_fa64_y1 | f_u_dadda_pg_rca16_fa64_y3;
  assign f_u_dadda_pg_rca16_and_9_6_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_9_6_y0 = f_u_dadda_pg_rca16_and_9_6_a_9 & f_u_dadda_pg_rca16_and_9_6_b_6;
  assign f_u_dadda_pg_rca16_and_8_7_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_8_7_y0 = f_u_dadda_pg_rca16_and_8_7_a_8 & f_u_dadda_pg_rca16_and_8_7_b_7;
  assign f_u_dadda_pg_rca16_and_7_8_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_7_8_y0 = f_u_dadda_pg_rca16_and_7_8_a_7 & f_u_dadda_pg_rca16_and_7_8_b_8;
  assign f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_9_6_y0 = f_u_dadda_pg_rca16_and_9_6_y0;
  assign f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_8_7_y0 = f_u_dadda_pg_rca16_and_8_7_y0;
  assign f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_7_8_y0 = f_u_dadda_pg_rca16_and_7_8_y0;
  assign f_u_dadda_pg_rca16_fa65_y0 = f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_9_6_y0 ^ f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_8_7_y0;
  assign f_u_dadda_pg_rca16_fa65_y1 = f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_9_6_y0 & f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_8_7_y0;
  assign f_u_dadda_pg_rca16_fa65_y2 = f_u_dadda_pg_rca16_fa65_y0 ^ f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_7_8_y0;
  assign f_u_dadda_pg_rca16_fa65_y3 = f_u_dadda_pg_rca16_fa65_y0 & f_u_dadda_pg_rca16_fa65_f_u_dadda_pg_rca16_and_7_8_y0;
  assign f_u_dadda_pg_rca16_fa65_y4 = f_u_dadda_pg_rca16_fa65_y1 | f_u_dadda_pg_rca16_fa65_y3;
  assign f_u_dadda_pg_rca16_and_6_9_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_6_9_y0 = f_u_dadda_pg_rca16_and_6_9_a_6 & f_u_dadda_pg_rca16_and_6_9_b_9;
  assign f_u_dadda_pg_rca16_and_5_10_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_5_10_y0 = f_u_dadda_pg_rca16_and_5_10_a_5 & f_u_dadda_pg_rca16_and_5_10_b_10;
  assign f_u_dadda_pg_rca16_and_4_11_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_4_11_y0 = f_u_dadda_pg_rca16_and_4_11_a_4 & f_u_dadda_pg_rca16_and_4_11_b_11;
  assign f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_6_9_y0 = f_u_dadda_pg_rca16_and_6_9_y0;
  assign f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_5_10_y0 = f_u_dadda_pg_rca16_and_5_10_y0;
  assign f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_4_11_y0 = f_u_dadda_pg_rca16_and_4_11_y0;
  assign f_u_dadda_pg_rca16_fa66_y0 = f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_6_9_y0 ^ f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_5_10_y0;
  assign f_u_dadda_pg_rca16_fa66_y1 = f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_6_9_y0 & f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_5_10_y0;
  assign f_u_dadda_pg_rca16_fa66_y2 = f_u_dadda_pg_rca16_fa66_y0 ^ f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_4_11_y0;
  assign f_u_dadda_pg_rca16_fa66_y3 = f_u_dadda_pg_rca16_fa66_y0 & f_u_dadda_pg_rca16_fa66_f_u_dadda_pg_rca16_and_4_11_y0;
  assign f_u_dadda_pg_rca16_fa66_y4 = f_u_dadda_pg_rca16_fa66_y1 | f_u_dadda_pg_rca16_fa66_y3;
  assign f_u_dadda_pg_rca16_and_3_12_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_3_12_y0 = f_u_dadda_pg_rca16_and_3_12_a_3 & f_u_dadda_pg_rca16_and_3_12_b_12;
  assign f_u_dadda_pg_rca16_and_2_13_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_2_13_y0 = f_u_dadda_pg_rca16_and_2_13_a_2 & f_u_dadda_pg_rca16_and_2_13_b_13;
  assign f_u_dadda_pg_rca16_and_1_14_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_1_14_y0 = f_u_dadda_pg_rca16_and_1_14_a_1 & f_u_dadda_pg_rca16_and_1_14_b_14;
  assign f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_3_12_y0 = f_u_dadda_pg_rca16_and_3_12_y0;
  assign f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_2_13_y0 = f_u_dadda_pg_rca16_and_2_13_y0;
  assign f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_1_14_y0 = f_u_dadda_pg_rca16_and_1_14_y0;
  assign f_u_dadda_pg_rca16_fa67_y0 = f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_3_12_y0 ^ f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_2_13_y0;
  assign f_u_dadda_pg_rca16_fa67_y1 = f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_3_12_y0 & f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_2_13_y0;
  assign f_u_dadda_pg_rca16_fa67_y2 = f_u_dadda_pg_rca16_fa67_y0 ^ f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_1_14_y0;
  assign f_u_dadda_pg_rca16_fa67_y3 = f_u_dadda_pg_rca16_fa67_y0 & f_u_dadda_pg_rca16_fa67_f_u_dadda_pg_rca16_and_1_14_y0;
  assign f_u_dadda_pg_rca16_fa67_y4 = f_u_dadda_pg_rca16_fa67_y1 | f_u_dadda_pg_rca16_fa67_y3;
  assign f_u_dadda_pg_rca16_and_0_15_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_0_15_y0 = f_u_dadda_pg_rca16_and_0_15_a_0 & f_u_dadda_pg_rca16_and_0_15_b_15;
  assign f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_and_0_15_y0 = f_u_dadda_pg_rca16_and_0_15_y0;
  assign f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_fa1_y2 = f_u_dadda_pg_rca16_fa1_y2;
  assign f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_fa2_y2 = f_u_dadda_pg_rca16_fa2_y2;
  assign f_u_dadda_pg_rca16_fa68_y0 = f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_and_0_15_y0 ^ f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_fa1_y2;
  assign f_u_dadda_pg_rca16_fa68_y1 = f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_and_0_15_y0 & f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_fa1_y2;
  assign f_u_dadda_pg_rca16_fa68_y2 = f_u_dadda_pg_rca16_fa68_y0 ^ f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_fa2_y2;
  assign f_u_dadda_pg_rca16_fa68_y3 = f_u_dadda_pg_rca16_fa68_y0 & f_u_dadda_pg_rca16_fa68_f_u_dadda_pg_rca16_fa2_y2;
  assign f_u_dadda_pg_rca16_fa68_y4 = f_u_dadda_pg_rca16_fa68_y1 | f_u_dadda_pg_rca16_fa68_y3;
  assign f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_ha2_y0 = f_u_dadda_pg_rca16_ha2_y0;
  assign f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_fa62_y2 = f_u_dadda_pg_rca16_fa62_y2;
  assign f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_fa63_y2 = f_u_dadda_pg_rca16_fa63_y2;
  assign f_u_dadda_pg_rca16_fa69_y0 = f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_ha2_y0 ^ f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_fa62_y2;
  assign f_u_dadda_pg_rca16_fa69_y1 = f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_ha2_y0 & f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_fa62_y2;
  assign f_u_dadda_pg_rca16_fa69_y2 = f_u_dadda_pg_rca16_fa69_y0 ^ f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_fa63_y2;
  assign f_u_dadda_pg_rca16_fa69_y3 = f_u_dadda_pg_rca16_fa69_y0 & f_u_dadda_pg_rca16_fa69_f_u_dadda_pg_rca16_fa63_y2;
  assign f_u_dadda_pg_rca16_fa69_y4 = f_u_dadda_pg_rca16_fa69_y1 | f_u_dadda_pg_rca16_fa69_y3;
  assign f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa64_y2 = f_u_dadda_pg_rca16_fa64_y2;
  assign f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa65_y2 = f_u_dadda_pg_rca16_fa65_y2;
  assign f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa66_y2 = f_u_dadda_pg_rca16_fa66_y2;
  assign f_u_dadda_pg_rca16_fa70_y0 = f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa64_y2 ^ f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa65_y2;
  assign f_u_dadda_pg_rca16_fa70_y1 = f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa64_y2 & f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa65_y2;
  assign f_u_dadda_pg_rca16_fa70_y2 = f_u_dadda_pg_rca16_fa70_y0 ^ f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa66_y2;
  assign f_u_dadda_pg_rca16_fa70_y3 = f_u_dadda_pg_rca16_fa70_y0 & f_u_dadda_pg_rca16_fa70_f_u_dadda_pg_rca16_fa66_y2;
  assign f_u_dadda_pg_rca16_fa70_y4 = f_u_dadda_pg_rca16_fa70_y1 | f_u_dadda_pg_rca16_fa70_y3;
  assign f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa70_y4 = f_u_dadda_pg_rca16_fa70_y4;
  assign f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa69_y4 = f_u_dadda_pg_rca16_fa69_y4;
  assign f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa68_y4 = f_u_dadda_pg_rca16_fa68_y4;
  assign f_u_dadda_pg_rca16_fa71_y0 = f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa70_y4 ^ f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa69_y4;
  assign f_u_dadda_pg_rca16_fa71_y1 = f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa70_y4 & f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa69_y4;
  assign f_u_dadda_pg_rca16_fa71_y2 = f_u_dadda_pg_rca16_fa71_y0 ^ f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa68_y4;
  assign f_u_dadda_pg_rca16_fa71_y3 = f_u_dadda_pg_rca16_fa71_y0 & f_u_dadda_pg_rca16_fa71_f_u_dadda_pg_rca16_fa68_y4;
  assign f_u_dadda_pg_rca16_fa71_y4 = f_u_dadda_pg_rca16_fa71_y1 | f_u_dadda_pg_rca16_fa71_y3;
  assign f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa67_y4 = f_u_dadda_pg_rca16_fa67_y4;
  assign f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa66_y4 = f_u_dadda_pg_rca16_fa66_y4;
  assign f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa65_y4 = f_u_dadda_pg_rca16_fa65_y4;
  assign f_u_dadda_pg_rca16_fa72_y0 = f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa67_y4 ^ f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa66_y4;
  assign f_u_dadda_pg_rca16_fa72_y1 = f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa67_y4 & f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa66_y4;
  assign f_u_dadda_pg_rca16_fa72_y2 = f_u_dadda_pg_rca16_fa72_y0 ^ f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa65_y4;
  assign f_u_dadda_pg_rca16_fa72_y3 = f_u_dadda_pg_rca16_fa72_y0 & f_u_dadda_pg_rca16_fa72_f_u_dadda_pg_rca16_fa65_y4;
  assign f_u_dadda_pg_rca16_fa72_y4 = f_u_dadda_pg_rca16_fa72_y1 | f_u_dadda_pg_rca16_fa72_y3;
  assign f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa64_y4 = f_u_dadda_pg_rca16_fa64_y4;
  assign f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa63_y4 = f_u_dadda_pg_rca16_fa63_y4;
  assign f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa62_y4 = f_u_dadda_pg_rca16_fa62_y4;
  assign f_u_dadda_pg_rca16_fa73_y0 = f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa64_y4 ^ f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa63_y4;
  assign f_u_dadda_pg_rca16_fa73_y1 = f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa64_y4 & f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa63_y4;
  assign f_u_dadda_pg_rca16_fa73_y2 = f_u_dadda_pg_rca16_fa73_y0 ^ f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa62_y4;
  assign f_u_dadda_pg_rca16_fa73_y3 = f_u_dadda_pg_rca16_fa73_y0 & f_u_dadda_pg_rca16_fa73_f_u_dadda_pg_rca16_fa62_y4;
  assign f_u_dadda_pg_rca16_fa73_y4 = f_u_dadda_pg_rca16_fa73_y1 | f_u_dadda_pg_rca16_fa73_y3;
  assign f_u_dadda_pg_rca16_and_10_6_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_10_6_y0 = f_u_dadda_pg_rca16_and_10_6_a_10 & f_u_dadda_pg_rca16_and_10_6_b_6;
  assign f_u_dadda_pg_rca16_and_9_7_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_9_7_y0 = f_u_dadda_pg_rca16_and_9_7_a_9 & f_u_dadda_pg_rca16_and_9_7_b_7;
  assign f_u_dadda_pg_rca16_and_8_8_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_8_8_y0 = f_u_dadda_pg_rca16_and_8_8_a_8 & f_u_dadda_pg_rca16_and_8_8_b_8;
  assign f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_10_6_y0 = f_u_dadda_pg_rca16_and_10_6_y0;
  assign f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_9_7_y0 = f_u_dadda_pg_rca16_and_9_7_y0;
  assign f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_8_8_y0 = f_u_dadda_pg_rca16_and_8_8_y0;
  assign f_u_dadda_pg_rca16_fa74_y0 = f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_10_6_y0 ^ f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_9_7_y0;
  assign f_u_dadda_pg_rca16_fa74_y1 = f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_10_6_y0 & f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_9_7_y0;
  assign f_u_dadda_pg_rca16_fa74_y2 = f_u_dadda_pg_rca16_fa74_y0 ^ f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_8_8_y0;
  assign f_u_dadda_pg_rca16_fa74_y3 = f_u_dadda_pg_rca16_fa74_y0 & f_u_dadda_pg_rca16_fa74_f_u_dadda_pg_rca16_and_8_8_y0;
  assign f_u_dadda_pg_rca16_fa74_y4 = f_u_dadda_pg_rca16_fa74_y1 | f_u_dadda_pg_rca16_fa74_y3;
  assign f_u_dadda_pg_rca16_and_7_9_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_7_9_y0 = f_u_dadda_pg_rca16_and_7_9_a_7 & f_u_dadda_pg_rca16_and_7_9_b_9;
  assign f_u_dadda_pg_rca16_and_6_10_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_6_10_y0 = f_u_dadda_pg_rca16_and_6_10_a_6 & f_u_dadda_pg_rca16_and_6_10_b_10;
  assign f_u_dadda_pg_rca16_and_5_11_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_5_11_y0 = f_u_dadda_pg_rca16_and_5_11_a_5 & f_u_dadda_pg_rca16_and_5_11_b_11;
  assign f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_7_9_y0 = f_u_dadda_pg_rca16_and_7_9_y0;
  assign f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_6_10_y0 = f_u_dadda_pg_rca16_and_6_10_y0;
  assign f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_5_11_y0 = f_u_dadda_pg_rca16_and_5_11_y0;
  assign f_u_dadda_pg_rca16_fa75_y0 = f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_7_9_y0 ^ f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_6_10_y0;
  assign f_u_dadda_pg_rca16_fa75_y1 = f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_7_9_y0 & f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_6_10_y0;
  assign f_u_dadda_pg_rca16_fa75_y2 = f_u_dadda_pg_rca16_fa75_y0 ^ f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_5_11_y0;
  assign f_u_dadda_pg_rca16_fa75_y3 = f_u_dadda_pg_rca16_fa75_y0 & f_u_dadda_pg_rca16_fa75_f_u_dadda_pg_rca16_and_5_11_y0;
  assign f_u_dadda_pg_rca16_fa75_y4 = f_u_dadda_pg_rca16_fa75_y1 | f_u_dadda_pg_rca16_fa75_y3;
  assign f_u_dadda_pg_rca16_and_4_12_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_4_12_y0 = f_u_dadda_pg_rca16_and_4_12_a_4 & f_u_dadda_pg_rca16_and_4_12_b_12;
  assign f_u_dadda_pg_rca16_and_3_13_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_3_13_y0 = f_u_dadda_pg_rca16_and_3_13_a_3 & f_u_dadda_pg_rca16_and_3_13_b_13;
  assign f_u_dadda_pg_rca16_and_2_14_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_2_14_y0 = f_u_dadda_pg_rca16_and_2_14_a_2 & f_u_dadda_pg_rca16_and_2_14_b_14;
  assign f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_4_12_y0 = f_u_dadda_pg_rca16_and_4_12_y0;
  assign f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_3_13_y0 = f_u_dadda_pg_rca16_and_3_13_y0;
  assign f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_2_14_y0 = f_u_dadda_pg_rca16_and_2_14_y0;
  assign f_u_dadda_pg_rca16_fa76_y0 = f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_4_12_y0 ^ f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_3_13_y0;
  assign f_u_dadda_pg_rca16_fa76_y1 = f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_4_12_y0 & f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_3_13_y0;
  assign f_u_dadda_pg_rca16_fa76_y2 = f_u_dadda_pg_rca16_fa76_y0 ^ f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_2_14_y0;
  assign f_u_dadda_pg_rca16_fa76_y3 = f_u_dadda_pg_rca16_fa76_y0 & f_u_dadda_pg_rca16_fa76_f_u_dadda_pg_rca16_and_2_14_y0;
  assign f_u_dadda_pg_rca16_fa76_y4 = f_u_dadda_pg_rca16_fa76_y1 | f_u_dadda_pg_rca16_fa76_y3;
  assign f_u_dadda_pg_rca16_and_1_15_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_1_15_y0 = f_u_dadda_pg_rca16_and_1_15_a_1 & f_u_dadda_pg_rca16_and_1_15_b_15;
  assign f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_and_1_15_y0 = f_u_dadda_pg_rca16_and_1_15_y0;
  assign f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_fa3_y2 = f_u_dadda_pg_rca16_fa3_y2;
  assign f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_fa4_y2 = f_u_dadda_pg_rca16_fa4_y2;
  assign f_u_dadda_pg_rca16_fa77_y0 = f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_and_1_15_y0 ^ f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_fa3_y2;
  assign f_u_dadda_pg_rca16_fa77_y1 = f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_and_1_15_y0 & f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_fa3_y2;
  assign f_u_dadda_pg_rca16_fa77_y2 = f_u_dadda_pg_rca16_fa77_y0 ^ f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_fa4_y2;
  assign f_u_dadda_pg_rca16_fa77_y3 = f_u_dadda_pg_rca16_fa77_y0 & f_u_dadda_pg_rca16_fa77_f_u_dadda_pg_rca16_fa4_y2;
  assign f_u_dadda_pg_rca16_fa77_y4 = f_u_dadda_pg_rca16_fa77_y1 | f_u_dadda_pg_rca16_fa77_y3;
  assign f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_ha3_y0 = f_u_dadda_pg_rca16_ha3_y0;
  assign f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_fa71_y2 = f_u_dadda_pg_rca16_fa71_y2;
  assign f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_fa72_y2 = f_u_dadda_pg_rca16_fa72_y2;
  assign f_u_dadda_pg_rca16_fa78_y0 = f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_ha3_y0 ^ f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_fa71_y2;
  assign f_u_dadda_pg_rca16_fa78_y1 = f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_ha3_y0 & f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_fa71_y2;
  assign f_u_dadda_pg_rca16_fa78_y2 = f_u_dadda_pg_rca16_fa78_y0 ^ f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_fa72_y2;
  assign f_u_dadda_pg_rca16_fa78_y3 = f_u_dadda_pg_rca16_fa78_y0 & f_u_dadda_pg_rca16_fa78_f_u_dadda_pg_rca16_fa72_y2;
  assign f_u_dadda_pg_rca16_fa78_y4 = f_u_dadda_pg_rca16_fa78_y1 | f_u_dadda_pg_rca16_fa78_y3;
  assign f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa73_y2 = f_u_dadda_pg_rca16_fa73_y2;
  assign f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa74_y2 = f_u_dadda_pg_rca16_fa74_y2;
  assign f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa75_y2 = f_u_dadda_pg_rca16_fa75_y2;
  assign f_u_dadda_pg_rca16_fa79_y0 = f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa73_y2 ^ f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa74_y2;
  assign f_u_dadda_pg_rca16_fa79_y1 = f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa73_y2 & f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa74_y2;
  assign f_u_dadda_pg_rca16_fa79_y2 = f_u_dadda_pg_rca16_fa79_y0 ^ f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa75_y2;
  assign f_u_dadda_pg_rca16_fa79_y3 = f_u_dadda_pg_rca16_fa79_y0 & f_u_dadda_pg_rca16_fa79_f_u_dadda_pg_rca16_fa75_y2;
  assign f_u_dadda_pg_rca16_fa79_y4 = f_u_dadda_pg_rca16_fa79_y1 | f_u_dadda_pg_rca16_fa79_y3;
  assign f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa79_y4 = f_u_dadda_pg_rca16_fa79_y4;
  assign f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa78_y4 = f_u_dadda_pg_rca16_fa78_y4;
  assign f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa77_y4 = f_u_dadda_pg_rca16_fa77_y4;
  assign f_u_dadda_pg_rca16_fa80_y0 = f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa79_y4 ^ f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa78_y4;
  assign f_u_dadda_pg_rca16_fa80_y1 = f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa79_y4 & f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa78_y4;
  assign f_u_dadda_pg_rca16_fa80_y2 = f_u_dadda_pg_rca16_fa80_y0 ^ f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa77_y4;
  assign f_u_dadda_pg_rca16_fa80_y3 = f_u_dadda_pg_rca16_fa80_y0 & f_u_dadda_pg_rca16_fa80_f_u_dadda_pg_rca16_fa77_y4;
  assign f_u_dadda_pg_rca16_fa80_y4 = f_u_dadda_pg_rca16_fa80_y1 | f_u_dadda_pg_rca16_fa80_y3;
  assign f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa76_y4 = f_u_dadda_pg_rca16_fa76_y4;
  assign f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa75_y4 = f_u_dadda_pg_rca16_fa75_y4;
  assign f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa74_y4 = f_u_dadda_pg_rca16_fa74_y4;
  assign f_u_dadda_pg_rca16_fa81_y0 = f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa76_y4 ^ f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa75_y4;
  assign f_u_dadda_pg_rca16_fa81_y1 = f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa76_y4 & f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa75_y4;
  assign f_u_dadda_pg_rca16_fa81_y2 = f_u_dadda_pg_rca16_fa81_y0 ^ f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa74_y4;
  assign f_u_dadda_pg_rca16_fa81_y3 = f_u_dadda_pg_rca16_fa81_y0 & f_u_dadda_pg_rca16_fa81_f_u_dadda_pg_rca16_fa74_y4;
  assign f_u_dadda_pg_rca16_fa81_y4 = f_u_dadda_pg_rca16_fa81_y1 | f_u_dadda_pg_rca16_fa81_y3;
  assign f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa73_y4 = f_u_dadda_pg_rca16_fa73_y4;
  assign f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa72_y4 = f_u_dadda_pg_rca16_fa72_y4;
  assign f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa71_y4 = f_u_dadda_pg_rca16_fa71_y4;
  assign f_u_dadda_pg_rca16_fa82_y0 = f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa73_y4 ^ f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa72_y4;
  assign f_u_dadda_pg_rca16_fa82_y1 = f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa73_y4 & f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa72_y4;
  assign f_u_dadda_pg_rca16_fa82_y2 = f_u_dadda_pg_rca16_fa82_y0 ^ f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa71_y4;
  assign f_u_dadda_pg_rca16_fa82_y3 = f_u_dadda_pg_rca16_fa82_y0 & f_u_dadda_pg_rca16_fa82_f_u_dadda_pg_rca16_fa71_y4;
  assign f_u_dadda_pg_rca16_fa82_y4 = f_u_dadda_pg_rca16_fa82_y1 | f_u_dadda_pg_rca16_fa82_y3;
  assign f_u_dadda_pg_rca16_and_12_5_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_12_5_y0 = f_u_dadda_pg_rca16_and_12_5_a_12 & f_u_dadda_pg_rca16_and_12_5_b_5;
  assign f_u_dadda_pg_rca16_and_11_6_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_11_6_y0 = f_u_dadda_pg_rca16_and_11_6_a_11 & f_u_dadda_pg_rca16_and_11_6_b_6;
  assign f_u_dadda_pg_rca16_and_10_7_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_10_7_y0 = f_u_dadda_pg_rca16_and_10_7_a_10 & f_u_dadda_pg_rca16_and_10_7_b_7;
  assign f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_12_5_y0 = f_u_dadda_pg_rca16_and_12_5_y0;
  assign f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_11_6_y0 = f_u_dadda_pg_rca16_and_11_6_y0;
  assign f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_10_7_y0 = f_u_dadda_pg_rca16_and_10_7_y0;
  assign f_u_dadda_pg_rca16_fa83_y0 = f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_12_5_y0 ^ f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_11_6_y0;
  assign f_u_dadda_pg_rca16_fa83_y1 = f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_12_5_y0 & f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_11_6_y0;
  assign f_u_dadda_pg_rca16_fa83_y2 = f_u_dadda_pg_rca16_fa83_y0 ^ f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_10_7_y0;
  assign f_u_dadda_pg_rca16_fa83_y3 = f_u_dadda_pg_rca16_fa83_y0 & f_u_dadda_pg_rca16_fa83_f_u_dadda_pg_rca16_and_10_7_y0;
  assign f_u_dadda_pg_rca16_fa83_y4 = f_u_dadda_pg_rca16_fa83_y1 | f_u_dadda_pg_rca16_fa83_y3;
  assign f_u_dadda_pg_rca16_and_9_8_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_9_8_y0 = f_u_dadda_pg_rca16_and_9_8_a_9 & f_u_dadda_pg_rca16_and_9_8_b_8;
  assign f_u_dadda_pg_rca16_and_8_9_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_8_9_y0 = f_u_dadda_pg_rca16_and_8_9_a_8 & f_u_dadda_pg_rca16_and_8_9_b_9;
  assign f_u_dadda_pg_rca16_and_7_10_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_7_10_y0 = f_u_dadda_pg_rca16_and_7_10_a_7 & f_u_dadda_pg_rca16_and_7_10_b_10;
  assign f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_9_8_y0 = f_u_dadda_pg_rca16_and_9_8_y0;
  assign f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_8_9_y0 = f_u_dadda_pg_rca16_and_8_9_y0;
  assign f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_7_10_y0 = f_u_dadda_pg_rca16_and_7_10_y0;
  assign f_u_dadda_pg_rca16_fa84_y0 = f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_9_8_y0 ^ f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_8_9_y0;
  assign f_u_dadda_pg_rca16_fa84_y1 = f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_9_8_y0 & f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_8_9_y0;
  assign f_u_dadda_pg_rca16_fa84_y2 = f_u_dadda_pg_rca16_fa84_y0 ^ f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_7_10_y0;
  assign f_u_dadda_pg_rca16_fa84_y3 = f_u_dadda_pg_rca16_fa84_y0 & f_u_dadda_pg_rca16_fa84_f_u_dadda_pg_rca16_and_7_10_y0;
  assign f_u_dadda_pg_rca16_fa84_y4 = f_u_dadda_pg_rca16_fa84_y1 | f_u_dadda_pg_rca16_fa84_y3;
  assign f_u_dadda_pg_rca16_and_6_11_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_6_11_y0 = f_u_dadda_pg_rca16_and_6_11_a_6 & f_u_dadda_pg_rca16_and_6_11_b_11;
  assign f_u_dadda_pg_rca16_and_5_12_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_5_12_y0 = f_u_dadda_pg_rca16_and_5_12_a_5 & f_u_dadda_pg_rca16_and_5_12_b_12;
  assign f_u_dadda_pg_rca16_and_4_13_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_4_13_y0 = f_u_dadda_pg_rca16_and_4_13_a_4 & f_u_dadda_pg_rca16_and_4_13_b_13;
  assign f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_6_11_y0 = f_u_dadda_pg_rca16_and_6_11_y0;
  assign f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_5_12_y0 = f_u_dadda_pg_rca16_and_5_12_y0;
  assign f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_4_13_y0 = f_u_dadda_pg_rca16_and_4_13_y0;
  assign f_u_dadda_pg_rca16_fa85_y0 = f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_6_11_y0 ^ f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_5_12_y0;
  assign f_u_dadda_pg_rca16_fa85_y1 = f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_6_11_y0 & f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_5_12_y0;
  assign f_u_dadda_pg_rca16_fa85_y2 = f_u_dadda_pg_rca16_fa85_y0 ^ f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_4_13_y0;
  assign f_u_dadda_pg_rca16_fa85_y3 = f_u_dadda_pg_rca16_fa85_y0 & f_u_dadda_pg_rca16_fa85_f_u_dadda_pg_rca16_and_4_13_y0;
  assign f_u_dadda_pg_rca16_fa85_y4 = f_u_dadda_pg_rca16_fa85_y1 | f_u_dadda_pg_rca16_fa85_y3;
  assign f_u_dadda_pg_rca16_and_3_14_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_3_14_y0 = f_u_dadda_pg_rca16_and_3_14_a_3 & f_u_dadda_pg_rca16_and_3_14_b_14;
  assign f_u_dadda_pg_rca16_and_2_15_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_2_15_y0 = f_u_dadda_pg_rca16_and_2_15_a_2 & f_u_dadda_pg_rca16_and_2_15_b_15;
  assign f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_and_3_14_y0 = f_u_dadda_pg_rca16_and_3_14_y0;
  assign f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_and_2_15_y0 = f_u_dadda_pg_rca16_and_2_15_y0;
  assign f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_fa5_y2 = f_u_dadda_pg_rca16_fa5_y2;
  assign f_u_dadda_pg_rca16_fa86_y0 = f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_and_3_14_y0 ^ f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_and_2_15_y0;
  assign f_u_dadda_pg_rca16_fa86_y1 = f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_and_3_14_y0 & f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_and_2_15_y0;
  assign f_u_dadda_pg_rca16_fa86_y2 = f_u_dadda_pg_rca16_fa86_y0 ^ f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_fa5_y2;
  assign f_u_dadda_pg_rca16_fa86_y3 = f_u_dadda_pg_rca16_fa86_y0 & f_u_dadda_pg_rca16_fa86_f_u_dadda_pg_rca16_fa5_y2;
  assign f_u_dadda_pg_rca16_fa86_y4 = f_u_dadda_pg_rca16_fa86_y1 | f_u_dadda_pg_rca16_fa86_y3;
  assign f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa6_y2 = f_u_dadda_pg_rca16_fa6_y2;
  assign f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa80_y2 = f_u_dadda_pg_rca16_fa80_y2;
  assign f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa81_y2 = f_u_dadda_pg_rca16_fa81_y2;
  assign f_u_dadda_pg_rca16_fa87_y0 = f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa6_y2 ^ f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa80_y2;
  assign f_u_dadda_pg_rca16_fa87_y1 = f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa6_y2 & f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa80_y2;
  assign f_u_dadda_pg_rca16_fa87_y2 = f_u_dadda_pg_rca16_fa87_y0 ^ f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa81_y2;
  assign f_u_dadda_pg_rca16_fa87_y3 = f_u_dadda_pg_rca16_fa87_y0 & f_u_dadda_pg_rca16_fa87_f_u_dadda_pg_rca16_fa81_y2;
  assign f_u_dadda_pg_rca16_fa87_y4 = f_u_dadda_pg_rca16_fa87_y1 | f_u_dadda_pg_rca16_fa87_y3;
  assign f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa82_y2 = f_u_dadda_pg_rca16_fa82_y2;
  assign f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa83_y2 = f_u_dadda_pg_rca16_fa83_y2;
  assign f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa84_y2 = f_u_dadda_pg_rca16_fa84_y2;
  assign f_u_dadda_pg_rca16_fa88_y0 = f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa82_y2 ^ f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa83_y2;
  assign f_u_dadda_pg_rca16_fa88_y1 = f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa82_y2 & f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa83_y2;
  assign f_u_dadda_pg_rca16_fa88_y2 = f_u_dadda_pg_rca16_fa88_y0 ^ f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa84_y2;
  assign f_u_dadda_pg_rca16_fa88_y3 = f_u_dadda_pg_rca16_fa88_y0 & f_u_dadda_pg_rca16_fa88_f_u_dadda_pg_rca16_fa84_y2;
  assign f_u_dadda_pg_rca16_fa88_y4 = f_u_dadda_pg_rca16_fa88_y1 | f_u_dadda_pg_rca16_fa88_y3;
  assign f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa88_y4 = f_u_dadda_pg_rca16_fa88_y4;
  assign f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa87_y4 = f_u_dadda_pg_rca16_fa87_y4;
  assign f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa86_y4 = f_u_dadda_pg_rca16_fa86_y4;
  assign f_u_dadda_pg_rca16_fa89_y0 = f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa88_y4 ^ f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa87_y4;
  assign f_u_dadda_pg_rca16_fa89_y1 = f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa88_y4 & f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa87_y4;
  assign f_u_dadda_pg_rca16_fa89_y2 = f_u_dadda_pg_rca16_fa89_y0 ^ f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa86_y4;
  assign f_u_dadda_pg_rca16_fa89_y3 = f_u_dadda_pg_rca16_fa89_y0 & f_u_dadda_pg_rca16_fa89_f_u_dadda_pg_rca16_fa86_y4;
  assign f_u_dadda_pg_rca16_fa89_y4 = f_u_dadda_pg_rca16_fa89_y1 | f_u_dadda_pg_rca16_fa89_y3;
  assign f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa85_y4 = f_u_dadda_pg_rca16_fa85_y4;
  assign f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa84_y4 = f_u_dadda_pg_rca16_fa84_y4;
  assign f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa83_y4 = f_u_dadda_pg_rca16_fa83_y4;
  assign f_u_dadda_pg_rca16_fa90_y0 = f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa85_y4 ^ f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa84_y4;
  assign f_u_dadda_pg_rca16_fa90_y1 = f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa85_y4 & f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa84_y4;
  assign f_u_dadda_pg_rca16_fa90_y2 = f_u_dadda_pg_rca16_fa90_y0 ^ f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa83_y4;
  assign f_u_dadda_pg_rca16_fa90_y3 = f_u_dadda_pg_rca16_fa90_y0 & f_u_dadda_pg_rca16_fa90_f_u_dadda_pg_rca16_fa83_y4;
  assign f_u_dadda_pg_rca16_fa90_y4 = f_u_dadda_pg_rca16_fa90_y1 | f_u_dadda_pg_rca16_fa90_y3;
  assign f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa82_y4 = f_u_dadda_pg_rca16_fa82_y4;
  assign f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa81_y4 = f_u_dadda_pg_rca16_fa81_y4;
  assign f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa80_y4 = f_u_dadda_pg_rca16_fa80_y4;
  assign f_u_dadda_pg_rca16_fa91_y0 = f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa82_y4 ^ f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa81_y4;
  assign f_u_dadda_pg_rca16_fa91_y1 = f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa82_y4 & f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa81_y4;
  assign f_u_dadda_pg_rca16_fa91_y2 = f_u_dadda_pg_rca16_fa91_y0 ^ f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa80_y4;
  assign f_u_dadda_pg_rca16_fa91_y3 = f_u_dadda_pg_rca16_fa91_y0 & f_u_dadda_pg_rca16_fa91_f_u_dadda_pg_rca16_fa80_y4;
  assign f_u_dadda_pg_rca16_fa91_y4 = f_u_dadda_pg_rca16_fa91_y1 | f_u_dadda_pg_rca16_fa91_y3;
  assign f_u_dadda_pg_rca16_and_14_4_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_14_4_y0 = f_u_dadda_pg_rca16_and_14_4_a_14 & f_u_dadda_pg_rca16_and_14_4_b_4;
  assign f_u_dadda_pg_rca16_and_13_5_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_13_5_y0 = f_u_dadda_pg_rca16_and_13_5_a_13 & f_u_dadda_pg_rca16_and_13_5_b_5;
  assign f_u_dadda_pg_rca16_and_12_6_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_12_6_y0 = f_u_dadda_pg_rca16_and_12_6_a_12 & f_u_dadda_pg_rca16_and_12_6_b_6;
  assign f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_14_4_y0 = f_u_dadda_pg_rca16_and_14_4_y0;
  assign f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_13_5_y0 = f_u_dadda_pg_rca16_and_13_5_y0;
  assign f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_12_6_y0 = f_u_dadda_pg_rca16_and_12_6_y0;
  assign f_u_dadda_pg_rca16_fa92_y0 = f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_14_4_y0 ^ f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_13_5_y0;
  assign f_u_dadda_pg_rca16_fa92_y1 = f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_14_4_y0 & f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_13_5_y0;
  assign f_u_dadda_pg_rca16_fa92_y2 = f_u_dadda_pg_rca16_fa92_y0 ^ f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_12_6_y0;
  assign f_u_dadda_pg_rca16_fa92_y3 = f_u_dadda_pg_rca16_fa92_y0 & f_u_dadda_pg_rca16_fa92_f_u_dadda_pg_rca16_and_12_6_y0;
  assign f_u_dadda_pg_rca16_fa92_y4 = f_u_dadda_pg_rca16_fa92_y1 | f_u_dadda_pg_rca16_fa92_y3;
  assign f_u_dadda_pg_rca16_and_11_7_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_11_7_y0 = f_u_dadda_pg_rca16_and_11_7_a_11 & f_u_dadda_pg_rca16_and_11_7_b_7;
  assign f_u_dadda_pg_rca16_and_10_8_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_10_8_y0 = f_u_dadda_pg_rca16_and_10_8_a_10 & f_u_dadda_pg_rca16_and_10_8_b_8;
  assign f_u_dadda_pg_rca16_and_9_9_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_9_9_y0 = f_u_dadda_pg_rca16_and_9_9_a_9 & f_u_dadda_pg_rca16_and_9_9_b_9;
  assign f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_11_7_y0 = f_u_dadda_pg_rca16_and_11_7_y0;
  assign f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_10_8_y0 = f_u_dadda_pg_rca16_and_10_8_y0;
  assign f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_9_9_y0 = f_u_dadda_pg_rca16_and_9_9_y0;
  assign f_u_dadda_pg_rca16_fa93_y0 = f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_11_7_y0 ^ f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_10_8_y0;
  assign f_u_dadda_pg_rca16_fa93_y1 = f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_11_7_y0 & f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_10_8_y0;
  assign f_u_dadda_pg_rca16_fa93_y2 = f_u_dadda_pg_rca16_fa93_y0 ^ f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_9_9_y0;
  assign f_u_dadda_pg_rca16_fa93_y3 = f_u_dadda_pg_rca16_fa93_y0 & f_u_dadda_pg_rca16_fa93_f_u_dadda_pg_rca16_and_9_9_y0;
  assign f_u_dadda_pg_rca16_fa93_y4 = f_u_dadda_pg_rca16_fa93_y1 | f_u_dadda_pg_rca16_fa93_y3;
  assign f_u_dadda_pg_rca16_and_8_10_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_8_10_y0 = f_u_dadda_pg_rca16_and_8_10_a_8 & f_u_dadda_pg_rca16_and_8_10_b_10;
  assign f_u_dadda_pg_rca16_and_7_11_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_7_11_y0 = f_u_dadda_pg_rca16_and_7_11_a_7 & f_u_dadda_pg_rca16_and_7_11_b_11;
  assign f_u_dadda_pg_rca16_and_6_12_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_6_12_y0 = f_u_dadda_pg_rca16_and_6_12_a_6 & f_u_dadda_pg_rca16_and_6_12_b_12;
  assign f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_8_10_y0 = f_u_dadda_pg_rca16_and_8_10_y0;
  assign f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_7_11_y0 = f_u_dadda_pg_rca16_and_7_11_y0;
  assign f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_6_12_y0 = f_u_dadda_pg_rca16_and_6_12_y0;
  assign f_u_dadda_pg_rca16_fa94_y0 = f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_8_10_y0 ^ f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_7_11_y0;
  assign f_u_dadda_pg_rca16_fa94_y1 = f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_8_10_y0 & f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_7_11_y0;
  assign f_u_dadda_pg_rca16_fa94_y2 = f_u_dadda_pg_rca16_fa94_y0 ^ f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_6_12_y0;
  assign f_u_dadda_pg_rca16_fa94_y3 = f_u_dadda_pg_rca16_fa94_y0 & f_u_dadda_pg_rca16_fa94_f_u_dadda_pg_rca16_and_6_12_y0;
  assign f_u_dadda_pg_rca16_fa94_y4 = f_u_dadda_pg_rca16_fa94_y1 | f_u_dadda_pg_rca16_fa94_y3;
  assign f_u_dadda_pg_rca16_and_5_13_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_5_13_y0 = f_u_dadda_pg_rca16_and_5_13_a_5 & f_u_dadda_pg_rca16_and_5_13_b_13;
  assign f_u_dadda_pg_rca16_and_4_14_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_4_14_y0 = f_u_dadda_pg_rca16_and_4_14_a_4 & f_u_dadda_pg_rca16_and_4_14_b_14;
  assign f_u_dadda_pg_rca16_and_3_15_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_3_15_y0 = f_u_dadda_pg_rca16_and_3_15_a_3 & f_u_dadda_pg_rca16_and_3_15_b_15;
  assign f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_5_13_y0 = f_u_dadda_pg_rca16_and_5_13_y0;
  assign f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_4_14_y0 = f_u_dadda_pg_rca16_and_4_14_y0;
  assign f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_3_15_y0 = f_u_dadda_pg_rca16_and_3_15_y0;
  assign f_u_dadda_pg_rca16_fa95_y0 = f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_5_13_y0 ^ f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_4_14_y0;
  assign f_u_dadda_pg_rca16_fa95_y1 = f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_5_13_y0 & f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_4_14_y0;
  assign f_u_dadda_pg_rca16_fa95_y2 = f_u_dadda_pg_rca16_fa95_y0 ^ f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_3_15_y0;
  assign f_u_dadda_pg_rca16_fa95_y3 = f_u_dadda_pg_rca16_fa95_y0 & f_u_dadda_pg_rca16_fa95_f_u_dadda_pg_rca16_and_3_15_y0;
  assign f_u_dadda_pg_rca16_fa95_y4 = f_u_dadda_pg_rca16_fa95_y1 | f_u_dadda_pg_rca16_fa95_y3;
  assign f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa7_y2 = f_u_dadda_pg_rca16_fa7_y2;
  assign f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa89_y2 = f_u_dadda_pg_rca16_fa89_y2;
  assign f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa90_y2 = f_u_dadda_pg_rca16_fa90_y2;
  assign f_u_dadda_pg_rca16_fa96_y0 = f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa7_y2 ^ f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa89_y2;
  assign f_u_dadda_pg_rca16_fa96_y1 = f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa7_y2 & f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa89_y2;
  assign f_u_dadda_pg_rca16_fa96_y2 = f_u_dadda_pg_rca16_fa96_y0 ^ f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa90_y2;
  assign f_u_dadda_pg_rca16_fa96_y3 = f_u_dadda_pg_rca16_fa96_y0 & f_u_dadda_pg_rca16_fa96_f_u_dadda_pg_rca16_fa90_y2;
  assign f_u_dadda_pg_rca16_fa96_y4 = f_u_dadda_pg_rca16_fa96_y1 | f_u_dadda_pg_rca16_fa96_y3;
  assign f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa91_y2 = f_u_dadda_pg_rca16_fa91_y2;
  assign f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa92_y2 = f_u_dadda_pg_rca16_fa92_y2;
  assign f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa93_y2 = f_u_dadda_pg_rca16_fa93_y2;
  assign f_u_dadda_pg_rca16_fa97_y0 = f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa91_y2 ^ f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa92_y2;
  assign f_u_dadda_pg_rca16_fa97_y1 = f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa91_y2 & f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa92_y2;
  assign f_u_dadda_pg_rca16_fa97_y2 = f_u_dadda_pg_rca16_fa97_y0 ^ f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa93_y2;
  assign f_u_dadda_pg_rca16_fa97_y3 = f_u_dadda_pg_rca16_fa97_y0 & f_u_dadda_pg_rca16_fa97_f_u_dadda_pg_rca16_fa93_y2;
  assign f_u_dadda_pg_rca16_fa97_y4 = f_u_dadda_pg_rca16_fa97_y1 | f_u_dadda_pg_rca16_fa97_y3;
  assign f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa97_y4 = f_u_dadda_pg_rca16_fa97_y4;
  assign f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa96_y4 = f_u_dadda_pg_rca16_fa96_y4;
  assign f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa95_y4 = f_u_dadda_pg_rca16_fa95_y4;
  assign f_u_dadda_pg_rca16_fa98_y0 = f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa97_y4 ^ f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa96_y4;
  assign f_u_dadda_pg_rca16_fa98_y1 = f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa97_y4 & f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa96_y4;
  assign f_u_dadda_pg_rca16_fa98_y2 = f_u_dadda_pg_rca16_fa98_y0 ^ f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa95_y4;
  assign f_u_dadda_pg_rca16_fa98_y3 = f_u_dadda_pg_rca16_fa98_y0 & f_u_dadda_pg_rca16_fa98_f_u_dadda_pg_rca16_fa95_y4;
  assign f_u_dadda_pg_rca16_fa98_y4 = f_u_dadda_pg_rca16_fa98_y1 | f_u_dadda_pg_rca16_fa98_y3;
  assign f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa94_y4 = f_u_dadda_pg_rca16_fa94_y4;
  assign f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa93_y4 = f_u_dadda_pg_rca16_fa93_y4;
  assign f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa92_y4 = f_u_dadda_pg_rca16_fa92_y4;
  assign f_u_dadda_pg_rca16_fa99_y0 = f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa94_y4 ^ f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa93_y4;
  assign f_u_dadda_pg_rca16_fa99_y1 = f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa94_y4 & f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa93_y4;
  assign f_u_dadda_pg_rca16_fa99_y2 = f_u_dadda_pg_rca16_fa99_y0 ^ f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa92_y4;
  assign f_u_dadda_pg_rca16_fa99_y3 = f_u_dadda_pg_rca16_fa99_y0 & f_u_dadda_pg_rca16_fa99_f_u_dadda_pg_rca16_fa92_y4;
  assign f_u_dadda_pg_rca16_fa99_y4 = f_u_dadda_pg_rca16_fa99_y1 | f_u_dadda_pg_rca16_fa99_y3;
  assign f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa91_y4 = f_u_dadda_pg_rca16_fa91_y4;
  assign f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa90_y4 = f_u_dadda_pg_rca16_fa90_y4;
  assign f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa89_y4 = f_u_dadda_pg_rca16_fa89_y4;
  assign f_u_dadda_pg_rca16_fa100_y0 = f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa91_y4 ^ f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa90_y4;
  assign f_u_dadda_pg_rca16_fa100_y1 = f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa91_y4 & f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa90_y4;
  assign f_u_dadda_pg_rca16_fa100_y2 = f_u_dadda_pg_rca16_fa100_y0 ^ f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa89_y4;
  assign f_u_dadda_pg_rca16_fa100_y3 = f_u_dadda_pg_rca16_fa100_y0 & f_u_dadda_pg_rca16_fa100_f_u_dadda_pg_rca16_fa89_y4;
  assign f_u_dadda_pg_rca16_fa100_y4 = f_u_dadda_pg_rca16_fa100_y1 | f_u_dadda_pg_rca16_fa100_y3;
  assign f_u_dadda_pg_rca16_and_15_4_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_15_4_y0 = f_u_dadda_pg_rca16_and_15_4_a_15 & f_u_dadda_pg_rca16_and_15_4_b_4;
  assign f_u_dadda_pg_rca16_and_14_5_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_14_5_y0 = f_u_dadda_pg_rca16_and_14_5_a_14 & f_u_dadda_pg_rca16_and_14_5_b_5;
  assign f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_fa7_y4 = f_u_dadda_pg_rca16_fa7_y4;
  assign f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_and_15_4_y0 = f_u_dadda_pg_rca16_and_15_4_y0;
  assign f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_and_14_5_y0 = f_u_dadda_pg_rca16_and_14_5_y0;
  assign f_u_dadda_pg_rca16_fa101_y0 = f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_fa7_y4 ^ f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_and_15_4_y0;
  assign f_u_dadda_pg_rca16_fa101_y1 = f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_fa7_y4 & f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_and_15_4_y0;
  assign f_u_dadda_pg_rca16_fa101_y2 = f_u_dadda_pg_rca16_fa101_y0 ^ f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_and_14_5_y0;
  assign f_u_dadda_pg_rca16_fa101_y3 = f_u_dadda_pg_rca16_fa101_y0 & f_u_dadda_pg_rca16_fa101_f_u_dadda_pg_rca16_and_14_5_y0;
  assign f_u_dadda_pg_rca16_fa101_y4 = f_u_dadda_pg_rca16_fa101_y1 | f_u_dadda_pg_rca16_fa101_y3;
  assign f_u_dadda_pg_rca16_and_13_6_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_13_6_y0 = f_u_dadda_pg_rca16_and_13_6_a_13 & f_u_dadda_pg_rca16_and_13_6_b_6;
  assign f_u_dadda_pg_rca16_and_12_7_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_12_7_y0 = f_u_dadda_pg_rca16_and_12_7_a_12 & f_u_dadda_pg_rca16_and_12_7_b_7;
  assign f_u_dadda_pg_rca16_and_11_8_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_11_8_y0 = f_u_dadda_pg_rca16_and_11_8_a_11 & f_u_dadda_pg_rca16_and_11_8_b_8;
  assign f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_13_6_y0 = f_u_dadda_pg_rca16_and_13_6_y0;
  assign f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_12_7_y0 = f_u_dadda_pg_rca16_and_12_7_y0;
  assign f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_11_8_y0 = f_u_dadda_pg_rca16_and_11_8_y0;
  assign f_u_dadda_pg_rca16_fa102_y0 = f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_13_6_y0 ^ f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_12_7_y0;
  assign f_u_dadda_pg_rca16_fa102_y1 = f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_13_6_y0 & f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_12_7_y0;
  assign f_u_dadda_pg_rca16_fa102_y2 = f_u_dadda_pg_rca16_fa102_y0 ^ f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_11_8_y0;
  assign f_u_dadda_pg_rca16_fa102_y3 = f_u_dadda_pg_rca16_fa102_y0 & f_u_dadda_pg_rca16_fa102_f_u_dadda_pg_rca16_and_11_8_y0;
  assign f_u_dadda_pg_rca16_fa102_y4 = f_u_dadda_pg_rca16_fa102_y1 | f_u_dadda_pg_rca16_fa102_y3;
  assign f_u_dadda_pg_rca16_and_10_9_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_10_9_y0 = f_u_dadda_pg_rca16_and_10_9_a_10 & f_u_dadda_pg_rca16_and_10_9_b_9;
  assign f_u_dadda_pg_rca16_and_9_10_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_9_10_y0 = f_u_dadda_pg_rca16_and_9_10_a_9 & f_u_dadda_pg_rca16_and_9_10_b_10;
  assign f_u_dadda_pg_rca16_and_8_11_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_8_11_y0 = f_u_dadda_pg_rca16_and_8_11_a_8 & f_u_dadda_pg_rca16_and_8_11_b_11;
  assign f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_10_9_y0 = f_u_dadda_pg_rca16_and_10_9_y0;
  assign f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_9_10_y0 = f_u_dadda_pg_rca16_and_9_10_y0;
  assign f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_8_11_y0 = f_u_dadda_pg_rca16_and_8_11_y0;
  assign f_u_dadda_pg_rca16_fa103_y0 = f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_10_9_y0 ^ f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_9_10_y0;
  assign f_u_dadda_pg_rca16_fa103_y1 = f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_10_9_y0 & f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_9_10_y0;
  assign f_u_dadda_pg_rca16_fa103_y2 = f_u_dadda_pg_rca16_fa103_y0 ^ f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_8_11_y0;
  assign f_u_dadda_pg_rca16_fa103_y3 = f_u_dadda_pg_rca16_fa103_y0 & f_u_dadda_pg_rca16_fa103_f_u_dadda_pg_rca16_and_8_11_y0;
  assign f_u_dadda_pg_rca16_fa103_y4 = f_u_dadda_pg_rca16_fa103_y1 | f_u_dadda_pg_rca16_fa103_y3;
  assign f_u_dadda_pg_rca16_and_7_12_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_7_12_y0 = f_u_dadda_pg_rca16_and_7_12_a_7 & f_u_dadda_pg_rca16_and_7_12_b_12;
  assign f_u_dadda_pg_rca16_and_6_13_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_6_13_y0 = f_u_dadda_pg_rca16_and_6_13_a_6 & f_u_dadda_pg_rca16_and_6_13_b_13;
  assign f_u_dadda_pg_rca16_and_5_14_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_5_14_y0 = f_u_dadda_pg_rca16_and_5_14_a_5 & f_u_dadda_pg_rca16_and_5_14_b_14;
  assign f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_7_12_y0 = f_u_dadda_pg_rca16_and_7_12_y0;
  assign f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_6_13_y0 = f_u_dadda_pg_rca16_and_6_13_y0;
  assign f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_5_14_y0 = f_u_dadda_pg_rca16_and_5_14_y0;
  assign f_u_dadda_pg_rca16_fa104_y0 = f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_7_12_y0 ^ f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_6_13_y0;
  assign f_u_dadda_pg_rca16_fa104_y1 = f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_7_12_y0 & f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_6_13_y0;
  assign f_u_dadda_pg_rca16_fa104_y2 = f_u_dadda_pg_rca16_fa104_y0 ^ f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_5_14_y0;
  assign f_u_dadda_pg_rca16_fa104_y3 = f_u_dadda_pg_rca16_fa104_y0 & f_u_dadda_pg_rca16_fa104_f_u_dadda_pg_rca16_and_5_14_y0;
  assign f_u_dadda_pg_rca16_fa104_y4 = f_u_dadda_pg_rca16_fa104_y1 | f_u_dadda_pg_rca16_fa104_y3;
  assign f_u_dadda_pg_rca16_and_4_15_a_4 = a_4;
  assign f_u_dadda_pg_rca16_and_4_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_4_15_y0 = f_u_dadda_pg_rca16_and_4_15_a_4 & f_u_dadda_pg_rca16_and_4_15_b_15;
  assign f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_and_4_15_y0 = f_u_dadda_pg_rca16_and_4_15_y0;
  assign f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_fa98_y2 = f_u_dadda_pg_rca16_fa98_y2;
  assign f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_fa99_y2 = f_u_dadda_pg_rca16_fa99_y2;
  assign f_u_dadda_pg_rca16_fa105_y0 = f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_and_4_15_y0 ^ f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_fa98_y2;
  assign f_u_dadda_pg_rca16_fa105_y1 = f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_and_4_15_y0 & f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_fa98_y2;
  assign f_u_dadda_pg_rca16_fa105_y2 = f_u_dadda_pg_rca16_fa105_y0 ^ f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_fa99_y2;
  assign f_u_dadda_pg_rca16_fa105_y3 = f_u_dadda_pg_rca16_fa105_y0 & f_u_dadda_pg_rca16_fa105_f_u_dadda_pg_rca16_fa99_y2;
  assign f_u_dadda_pg_rca16_fa105_y4 = f_u_dadda_pg_rca16_fa105_y1 | f_u_dadda_pg_rca16_fa105_y3;
  assign f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa100_y2 = f_u_dadda_pg_rca16_fa100_y2;
  assign f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa101_y2 = f_u_dadda_pg_rca16_fa101_y2;
  assign f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa102_y2 = f_u_dadda_pg_rca16_fa102_y2;
  assign f_u_dadda_pg_rca16_fa106_y0 = f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa100_y2 ^ f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa101_y2;
  assign f_u_dadda_pg_rca16_fa106_y1 = f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa100_y2 & f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa101_y2;
  assign f_u_dadda_pg_rca16_fa106_y2 = f_u_dadda_pg_rca16_fa106_y0 ^ f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa102_y2;
  assign f_u_dadda_pg_rca16_fa106_y3 = f_u_dadda_pg_rca16_fa106_y0 & f_u_dadda_pg_rca16_fa106_f_u_dadda_pg_rca16_fa102_y2;
  assign f_u_dadda_pg_rca16_fa106_y4 = f_u_dadda_pg_rca16_fa106_y1 | f_u_dadda_pg_rca16_fa106_y3;
  assign f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa106_y4 = f_u_dadda_pg_rca16_fa106_y4;
  assign f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa105_y4 = f_u_dadda_pg_rca16_fa105_y4;
  assign f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa104_y4 = f_u_dadda_pg_rca16_fa104_y4;
  assign f_u_dadda_pg_rca16_fa107_y0 = f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa106_y4 ^ f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa105_y4;
  assign f_u_dadda_pg_rca16_fa107_y1 = f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa106_y4 & f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa105_y4;
  assign f_u_dadda_pg_rca16_fa107_y2 = f_u_dadda_pg_rca16_fa107_y0 ^ f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa104_y4;
  assign f_u_dadda_pg_rca16_fa107_y3 = f_u_dadda_pg_rca16_fa107_y0 & f_u_dadda_pg_rca16_fa107_f_u_dadda_pg_rca16_fa104_y4;
  assign f_u_dadda_pg_rca16_fa107_y4 = f_u_dadda_pg_rca16_fa107_y1 | f_u_dadda_pg_rca16_fa107_y3;
  assign f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa103_y4 = f_u_dadda_pg_rca16_fa103_y4;
  assign f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa102_y4 = f_u_dadda_pg_rca16_fa102_y4;
  assign f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa101_y4 = f_u_dadda_pg_rca16_fa101_y4;
  assign f_u_dadda_pg_rca16_fa108_y0 = f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa103_y4 ^ f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa102_y4;
  assign f_u_dadda_pg_rca16_fa108_y1 = f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa103_y4 & f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa102_y4;
  assign f_u_dadda_pg_rca16_fa108_y2 = f_u_dadda_pg_rca16_fa108_y0 ^ f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa101_y4;
  assign f_u_dadda_pg_rca16_fa108_y3 = f_u_dadda_pg_rca16_fa108_y0 & f_u_dadda_pg_rca16_fa108_f_u_dadda_pg_rca16_fa101_y4;
  assign f_u_dadda_pg_rca16_fa108_y4 = f_u_dadda_pg_rca16_fa108_y1 | f_u_dadda_pg_rca16_fa108_y3;
  assign f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa100_y4 = f_u_dadda_pg_rca16_fa100_y4;
  assign f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa99_y4 = f_u_dadda_pg_rca16_fa99_y4;
  assign f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa98_y4 = f_u_dadda_pg_rca16_fa98_y4;
  assign f_u_dadda_pg_rca16_fa109_y0 = f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa100_y4 ^ f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa99_y4;
  assign f_u_dadda_pg_rca16_fa109_y1 = f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa100_y4 & f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa99_y4;
  assign f_u_dadda_pg_rca16_fa109_y2 = f_u_dadda_pg_rca16_fa109_y0 ^ f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa98_y4;
  assign f_u_dadda_pg_rca16_fa109_y3 = f_u_dadda_pg_rca16_fa109_y0 & f_u_dadda_pg_rca16_fa109_f_u_dadda_pg_rca16_fa98_y4;
  assign f_u_dadda_pg_rca16_fa109_y4 = f_u_dadda_pg_rca16_fa109_y1 | f_u_dadda_pg_rca16_fa109_y3;
  assign f_u_dadda_pg_rca16_and_15_5_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_15_5_y0 = f_u_dadda_pg_rca16_and_15_5_a_15 & f_u_dadda_pg_rca16_and_15_5_b_5;
  assign f_u_dadda_pg_rca16_and_14_6_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_14_6_y0 = f_u_dadda_pg_rca16_and_14_6_a_14 & f_u_dadda_pg_rca16_and_14_6_b_6;
  assign f_u_dadda_pg_rca16_and_13_7_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_13_7_y0 = f_u_dadda_pg_rca16_and_13_7_a_13 & f_u_dadda_pg_rca16_and_13_7_b_7;
  assign f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_15_5_y0 = f_u_dadda_pg_rca16_and_15_5_y0;
  assign f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_14_6_y0 = f_u_dadda_pg_rca16_and_14_6_y0;
  assign f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_13_7_y0 = f_u_dadda_pg_rca16_and_13_7_y0;
  assign f_u_dadda_pg_rca16_fa110_y0 = f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_15_5_y0 ^ f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_14_6_y0;
  assign f_u_dadda_pg_rca16_fa110_y1 = f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_15_5_y0 & f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_14_6_y0;
  assign f_u_dadda_pg_rca16_fa110_y2 = f_u_dadda_pg_rca16_fa110_y0 ^ f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_13_7_y0;
  assign f_u_dadda_pg_rca16_fa110_y3 = f_u_dadda_pg_rca16_fa110_y0 & f_u_dadda_pg_rca16_fa110_f_u_dadda_pg_rca16_and_13_7_y0;
  assign f_u_dadda_pg_rca16_fa110_y4 = f_u_dadda_pg_rca16_fa110_y1 | f_u_dadda_pg_rca16_fa110_y3;
  assign f_u_dadda_pg_rca16_and_12_8_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_12_8_y0 = f_u_dadda_pg_rca16_and_12_8_a_12 & f_u_dadda_pg_rca16_and_12_8_b_8;
  assign f_u_dadda_pg_rca16_and_11_9_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_11_9_y0 = f_u_dadda_pg_rca16_and_11_9_a_11 & f_u_dadda_pg_rca16_and_11_9_b_9;
  assign f_u_dadda_pg_rca16_and_10_10_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_10_10_y0 = f_u_dadda_pg_rca16_and_10_10_a_10 & f_u_dadda_pg_rca16_and_10_10_b_10;
  assign f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_12_8_y0 = f_u_dadda_pg_rca16_and_12_8_y0;
  assign f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_11_9_y0 = f_u_dadda_pg_rca16_and_11_9_y0;
  assign f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_10_10_y0 = f_u_dadda_pg_rca16_and_10_10_y0;
  assign f_u_dadda_pg_rca16_fa111_y0 = f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_12_8_y0 ^ f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_11_9_y0;
  assign f_u_dadda_pg_rca16_fa111_y1 = f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_12_8_y0 & f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_11_9_y0;
  assign f_u_dadda_pg_rca16_fa111_y2 = f_u_dadda_pg_rca16_fa111_y0 ^ f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_10_10_y0;
  assign f_u_dadda_pg_rca16_fa111_y3 = f_u_dadda_pg_rca16_fa111_y0 & f_u_dadda_pg_rca16_fa111_f_u_dadda_pg_rca16_and_10_10_y0;
  assign f_u_dadda_pg_rca16_fa111_y4 = f_u_dadda_pg_rca16_fa111_y1 | f_u_dadda_pg_rca16_fa111_y3;
  assign f_u_dadda_pg_rca16_and_9_11_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_9_11_y0 = f_u_dadda_pg_rca16_and_9_11_a_9 & f_u_dadda_pg_rca16_and_9_11_b_11;
  assign f_u_dadda_pg_rca16_and_8_12_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_8_12_y0 = f_u_dadda_pg_rca16_and_8_12_a_8 & f_u_dadda_pg_rca16_and_8_12_b_12;
  assign f_u_dadda_pg_rca16_and_7_13_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_7_13_y0 = f_u_dadda_pg_rca16_and_7_13_a_7 & f_u_dadda_pg_rca16_and_7_13_b_13;
  assign f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_9_11_y0 = f_u_dadda_pg_rca16_and_9_11_y0;
  assign f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_8_12_y0 = f_u_dadda_pg_rca16_and_8_12_y0;
  assign f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_7_13_y0 = f_u_dadda_pg_rca16_and_7_13_y0;
  assign f_u_dadda_pg_rca16_fa112_y0 = f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_9_11_y0 ^ f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_8_12_y0;
  assign f_u_dadda_pg_rca16_fa112_y1 = f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_9_11_y0 & f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_8_12_y0;
  assign f_u_dadda_pg_rca16_fa112_y2 = f_u_dadda_pg_rca16_fa112_y0 ^ f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_7_13_y0;
  assign f_u_dadda_pg_rca16_fa112_y3 = f_u_dadda_pg_rca16_fa112_y0 & f_u_dadda_pg_rca16_fa112_f_u_dadda_pg_rca16_and_7_13_y0;
  assign f_u_dadda_pg_rca16_fa112_y4 = f_u_dadda_pg_rca16_fa112_y1 | f_u_dadda_pg_rca16_fa112_y3;
  assign f_u_dadda_pg_rca16_and_6_14_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_6_14_y0 = f_u_dadda_pg_rca16_and_6_14_a_6 & f_u_dadda_pg_rca16_and_6_14_b_14;
  assign f_u_dadda_pg_rca16_and_5_15_a_5 = a_5;
  assign f_u_dadda_pg_rca16_and_5_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_5_15_y0 = f_u_dadda_pg_rca16_and_5_15_a_5 & f_u_dadda_pg_rca16_and_5_15_b_15;
  assign f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_and_6_14_y0 = f_u_dadda_pg_rca16_and_6_14_y0;
  assign f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_and_5_15_y0 = f_u_dadda_pg_rca16_and_5_15_y0;
  assign f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_fa107_y2 = f_u_dadda_pg_rca16_fa107_y2;
  assign f_u_dadda_pg_rca16_fa113_y0 = f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_and_6_14_y0 ^ f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_and_5_15_y0;
  assign f_u_dadda_pg_rca16_fa113_y1 = f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_and_6_14_y0 & f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_and_5_15_y0;
  assign f_u_dadda_pg_rca16_fa113_y2 = f_u_dadda_pg_rca16_fa113_y0 ^ f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_fa107_y2;
  assign f_u_dadda_pg_rca16_fa113_y3 = f_u_dadda_pg_rca16_fa113_y0 & f_u_dadda_pg_rca16_fa113_f_u_dadda_pg_rca16_fa107_y2;
  assign f_u_dadda_pg_rca16_fa113_y4 = f_u_dadda_pg_rca16_fa113_y1 | f_u_dadda_pg_rca16_fa113_y3;
  assign f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa108_y2 = f_u_dadda_pg_rca16_fa108_y2;
  assign f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa109_y2 = f_u_dadda_pg_rca16_fa109_y2;
  assign f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa110_y2 = f_u_dadda_pg_rca16_fa110_y2;
  assign f_u_dadda_pg_rca16_fa114_y0 = f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa108_y2 ^ f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa109_y2;
  assign f_u_dadda_pg_rca16_fa114_y1 = f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa108_y2 & f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa109_y2;
  assign f_u_dadda_pg_rca16_fa114_y2 = f_u_dadda_pg_rca16_fa114_y0 ^ f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa110_y2;
  assign f_u_dadda_pg_rca16_fa114_y3 = f_u_dadda_pg_rca16_fa114_y0 & f_u_dadda_pg_rca16_fa114_f_u_dadda_pg_rca16_fa110_y2;
  assign f_u_dadda_pg_rca16_fa114_y4 = f_u_dadda_pg_rca16_fa114_y1 | f_u_dadda_pg_rca16_fa114_y3;
  assign f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa114_y4 = f_u_dadda_pg_rca16_fa114_y4;
  assign f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa113_y4 = f_u_dadda_pg_rca16_fa113_y4;
  assign f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa112_y4 = f_u_dadda_pg_rca16_fa112_y4;
  assign f_u_dadda_pg_rca16_fa115_y0 = f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa114_y4 ^ f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa113_y4;
  assign f_u_dadda_pg_rca16_fa115_y1 = f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa114_y4 & f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa113_y4;
  assign f_u_dadda_pg_rca16_fa115_y2 = f_u_dadda_pg_rca16_fa115_y0 ^ f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa112_y4;
  assign f_u_dadda_pg_rca16_fa115_y3 = f_u_dadda_pg_rca16_fa115_y0 & f_u_dadda_pg_rca16_fa115_f_u_dadda_pg_rca16_fa112_y4;
  assign f_u_dadda_pg_rca16_fa115_y4 = f_u_dadda_pg_rca16_fa115_y1 | f_u_dadda_pg_rca16_fa115_y3;
  assign f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa111_y4 = f_u_dadda_pg_rca16_fa111_y4;
  assign f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa110_y4 = f_u_dadda_pg_rca16_fa110_y4;
  assign f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa109_y4 = f_u_dadda_pg_rca16_fa109_y4;
  assign f_u_dadda_pg_rca16_fa116_y0 = f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa111_y4 ^ f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa110_y4;
  assign f_u_dadda_pg_rca16_fa116_y1 = f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa111_y4 & f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa110_y4;
  assign f_u_dadda_pg_rca16_fa116_y2 = f_u_dadda_pg_rca16_fa116_y0 ^ f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa109_y4;
  assign f_u_dadda_pg_rca16_fa116_y3 = f_u_dadda_pg_rca16_fa116_y0 & f_u_dadda_pg_rca16_fa116_f_u_dadda_pg_rca16_fa109_y4;
  assign f_u_dadda_pg_rca16_fa116_y4 = f_u_dadda_pg_rca16_fa116_y1 | f_u_dadda_pg_rca16_fa116_y3;
  assign f_u_dadda_pg_rca16_and_15_6_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_15_6_y0 = f_u_dadda_pg_rca16_and_15_6_a_15 & f_u_dadda_pg_rca16_and_15_6_b_6;
  assign f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_fa108_y4 = f_u_dadda_pg_rca16_fa108_y4;
  assign f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_fa107_y4 = f_u_dadda_pg_rca16_fa107_y4;
  assign f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_and_15_6_y0 = f_u_dadda_pg_rca16_and_15_6_y0;
  assign f_u_dadda_pg_rca16_fa117_y0 = f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_fa108_y4 ^ f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_fa107_y4;
  assign f_u_dadda_pg_rca16_fa117_y1 = f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_fa108_y4 & f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_fa107_y4;
  assign f_u_dadda_pg_rca16_fa117_y2 = f_u_dadda_pg_rca16_fa117_y0 ^ f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_and_15_6_y0;
  assign f_u_dadda_pg_rca16_fa117_y3 = f_u_dadda_pg_rca16_fa117_y0 & f_u_dadda_pg_rca16_fa117_f_u_dadda_pg_rca16_and_15_6_y0;
  assign f_u_dadda_pg_rca16_fa117_y4 = f_u_dadda_pg_rca16_fa117_y1 | f_u_dadda_pg_rca16_fa117_y3;
  assign f_u_dadda_pg_rca16_and_14_7_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_14_7_y0 = f_u_dadda_pg_rca16_and_14_7_a_14 & f_u_dadda_pg_rca16_and_14_7_b_7;
  assign f_u_dadda_pg_rca16_and_13_8_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_13_8_y0 = f_u_dadda_pg_rca16_and_13_8_a_13 & f_u_dadda_pg_rca16_and_13_8_b_8;
  assign f_u_dadda_pg_rca16_and_12_9_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_12_9_y0 = f_u_dadda_pg_rca16_and_12_9_a_12 & f_u_dadda_pg_rca16_and_12_9_b_9;
  assign f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_14_7_y0 = f_u_dadda_pg_rca16_and_14_7_y0;
  assign f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_13_8_y0 = f_u_dadda_pg_rca16_and_13_8_y0;
  assign f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_12_9_y0 = f_u_dadda_pg_rca16_and_12_9_y0;
  assign f_u_dadda_pg_rca16_fa118_y0 = f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_14_7_y0 ^ f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_13_8_y0;
  assign f_u_dadda_pg_rca16_fa118_y1 = f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_14_7_y0 & f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_13_8_y0;
  assign f_u_dadda_pg_rca16_fa118_y2 = f_u_dadda_pg_rca16_fa118_y0 ^ f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_12_9_y0;
  assign f_u_dadda_pg_rca16_fa118_y3 = f_u_dadda_pg_rca16_fa118_y0 & f_u_dadda_pg_rca16_fa118_f_u_dadda_pg_rca16_and_12_9_y0;
  assign f_u_dadda_pg_rca16_fa118_y4 = f_u_dadda_pg_rca16_fa118_y1 | f_u_dadda_pg_rca16_fa118_y3;
  assign f_u_dadda_pg_rca16_and_11_10_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_11_10_y0 = f_u_dadda_pg_rca16_and_11_10_a_11 & f_u_dadda_pg_rca16_and_11_10_b_10;
  assign f_u_dadda_pg_rca16_and_10_11_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_10_11_y0 = f_u_dadda_pg_rca16_and_10_11_a_10 & f_u_dadda_pg_rca16_and_10_11_b_11;
  assign f_u_dadda_pg_rca16_and_9_12_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_9_12_y0 = f_u_dadda_pg_rca16_and_9_12_a_9 & f_u_dadda_pg_rca16_and_9_12_b_12;
  assign f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_11_10_y0 = f_u_dadda_pg_rca16_and_11_10_y0;
  assign f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_10_11_y0 = f_u_dadda_pg_rca16_and_10_11_y0;
  assign f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_9_12_y0 = f_u_dadda_pg_rca16_and_9_12_y0;
  assign f_u_dadda_pg_rca16_fa119_y0 = f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_11_10_y0 ^ f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_10_11_y0;
  assign f_u_dadda_pg_rca16_fa119_y1 = f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_11_10_y0 & f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_10_11_y0;
  assign f_u_dadda_pg_rca16_fa119_y2 = f_u_dadda_pg_rca16_fa119_y0 ^ f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_9_12_y0;
  assign f_u_dadda_pg_rca16_fa119_y3 = f_u_dadda_pg_rca16_fa119_y0 & f_u_dadda_pg_rca16_fa119_f_u_dadda_pg_rca16_and_9_12_y0;
  assign f_u_dadda_pg_rca16_fa119_y4 = f_u_dadda_pg_rca16_fa119_y1 | f_u_dadda_pg_rca16_fa119_y3;
  assign f_u_dadda_pg_rca16_and_8_13_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_8_13_y0 = f_u_dadda_pg_rca16_and_8_13_a_8 & f_u_dadda_pg_rca16_and_8_13_b_13;
  assign f_u_dadda_pg_rca16_and_7_14_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_7_14_y0 = f_u_dadda_pg_rca16_and_7_14_a_7 & f_u_dadda_pg_rca16_and_7_14_b_14;
  assign f_u_dadda_pg_rca16_and_6_15_a_6 = a_6;
  assign f_u_dadda_pg_rca16_and_6_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_6_15_y0 = f_u_dadda_pg_rca16_and_6_15_a_6 & f_u_dadda_pg_rca16_and_6_15_b_15;
  assign f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_8_13_y0 = f_u_dadda_pg_rca16_and_8_13_y0;
  assign f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_7_14_y0 = f_u_dadda_pg_rca16_and_7_14_y0;
  assign f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_6_15_y0 = f_u_dadda_pg_rca16_and_6_15_y0;
  assign f_u_dadda_pg_rca16_fa120_y0 = f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_8_13_y0 ^ f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_7_14_y0;
  assign f_u_dadda_pg_rca16_fa120_y1 = f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_8_13_y0 & f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_7_14_y0;
  assign f_u_dadda_pg_rca16_fa120_y2 = f_u_dadda_pg_rca16_fa120_y0 ^ f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_6_15_y0;
  assign f_u_dadda_pg_rca16_fa120_y3 = f_u_dadda_pg_rca16_fa120_y0 & f_u_dadda_pg_rca16_fa120_f_u_dadda_pg_rca16_and_6_15_y0;
  assign f_u_dadda_pg_rca16_fa120_y4 = f_u_dadda_pg_rca16_fa120_y1 | f_u_dadda_pg_rca16_fa120_y3;
  assign f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa115_y2 = f_u_dadda_pg_rca16_fa115_y2;
  assign f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa116_y2 = f_u_dadda_pg_rca16_fa116_y2;
  assign f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa117_y2 = f_u_dadda_pg_rca16_fa117_y2;
  assign f_u_dadda_pg_rca16_fa121_y0 = f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa115_y2 ^ f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa116_y2;
  assign f_u_dadda_pg_rca16_fa121_y1 = f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa115_y2 & f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa116_y2;
  assign f_u_dadda_pg_rca16_fa121_y2 = f_u_dadda_pg_rca16_fa121_y0 ^ f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa117_y2;
  assign f_u_dadda_pg_rca16_fa121_y3 = f_u_dadda_pg_rca16_fa121_y0 & f_u_dadda_pg_rca16_fa121_f_u_dadda_pg_rca16_fa117_y2;
  assign f_u_dadda_pg_rca16_fa121_y4 = f_u_dadda_pg_rca16_fa121_y1 | f_u_dadda_pg_rca16_fa121_y3;
  assign f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa121_y4 = f_u_dadda_pg_rca16_fa121_y4;
  assign f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa120_y4 = f_u_dadda_pg_rca16_fa120_y4;
  assign f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa119_y4 = f_u_dadda_pg_rca16_fa119_y4;
  assign f_u_dadda_pg_rca16_fa122_y0 = f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa121_y4 ^ f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa120_y4;
  assign f_u_dadda_pg_rca16_fa122_y1 = f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa121_y4 & f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa120_y4;
  assign f_u_dadda_pg_rca16_fa122_y2 = f_u_dadda_pg_rca16_fa122_y0 ^ f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa119_y4;
  assign f_u_dadda_pg_rca16_fa122_y3 = f_u_dadda_pg_rca16_fa122_y0 & f_u_dadda_pg_rca16_fa122_f_u_dadda_pg_rca16_fa119_y4;
  assign f_u_dadda_pg_rca16_fa122_y4 = f_u_dadda_pg_rca16_fa122_y1 | f_u_dadda_pg_rca16_fa122_y3;
  assign f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa118_y4 = f_u_dadda_pg_rca16_fa118_y4;
  assign f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa117_y4 = f_u_dadda_pg_rca16_fa117_y4;
  assign f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa116_y4 = f_u_dadda_pg_rca16_fa116_y4;
  assign f_u_dadda_pg_rca16_fa123_y0 = f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa118_y4 ^ f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa117_y4;
  assign f_u_dadda_pg_rca16_fa123_y1 = f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa118_y4 & f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa117_y4;
  assign f_u_dadda_pg_rca16_fa123_y2 = f_u_dadda_pg_rca16_fa123_y0 ^ f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa116_y4;
  assign f_u_dadda_pg_rca16_fa123_y3 = f_u_dadda_pg_rca16_fa123_y0 & f_u_dadda_pg_rca16_fa123_f_u_dadda_pg_rca16_fa116_y4;
  assign f_u_dadda_pg_rca16_fa123_y4 = f_u_dadda_pg_rca16_fa123_y1 | f_u_dadda_pg_rca16_fa123_y3;
  assign f_u_dadda_pg_rca16_and_15_7_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_7_b_7 = b_7;
  assign f_u_dadda_pg_rca16_and_15_7_y0 = f_u_dadda_pg_rca16_and_15_7_a_15 & f_u_dadda_pg_rca16_and_15_7_b_7;
  assign f_u_dadda_pg_rca16_and_14_8_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_14_8_y0 = f_u_dadda_pg_rca16_and_14_8_a_14 & f_u_dadda_pg_rca16_and_14_8_b_8;
  assign f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_fa115_y4 = f_u_dadda_pg_rca16_fa115_y4;
  assign f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_and_15_7_y0 = f_u_dadda_pg_rca16_and_15_7_y0;
  assign f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_and_14_8_y0 = f_u_dadda_pg_rca16_and_14_8_y0;
  assign f_u_dadda_pg_rca16_fa124_y0 = f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_fa115_y4 ^ f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_and_15_7_y0;
  assign f_u_dadda_pg_rca16_fa124_y1 = f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_fa115_y4 & f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_and_15_7_y0;
  assign f_u_dadda_pg_rca16_fa124_y2 = f_u_dadda_pg_rca16_fa124_y0 ^ f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_and_14_8_y0;
  assign f_u_dadda_pg_rca16_fa124_y3 = f_u_dadda_pg_rca16_fa124_y0 & f_u_dadda_pg_rca16_fa124_f_u_dadda_pg_rca16_and_14_8_y0;
  assign f_u_dadda_pg_rca16_fa124_y4 = f_u_dadda_pg_rca16_fa124_y1 | f_u_dadda_pg_rca16_fa124_y3;
  assign f_u_dadda_pg_rca16_and_13_9_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_13_9_y0 = f_u_dadda_pg_rca16_and_13_9_a_13 & f_u_dadda_pg_rca16_and_13_9_b_9;
  assign f_u_dadda_pg_rca16_and_12_10_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_12_10_y0 = f_u_dadda_pg_rca16_and_12_10_a_12 & f_u_dadda_pg_rca16_and_12_10_b_10;
  assign f_u_dadda_pg_rca16_and_11_11_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_11_11_y0 = f_u_dadda_pg_rca16_and_11_11_a_11 & f_u_dadda_pg_rca16_and_11_11_b_11;
  assign f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_13_9_y0 = f_u_dadda_pg_rca16_and_13_9_y0;
  assign f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_12_10_y0 = f_u_dadda_pg_rca16_and_12_10_y0;
  assign f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_11_11_y0 = f_u_dadda_pg_rca16_and_11_11_y0;
  assign f_u_dadda_pg_rca16_fa125_y0 = f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_13_9_y0 ^ f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_12_10_y0;
  assign f_u_dadda_pg_rca16_fa125_y1 = f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_13_9_y0 & f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_12_10_y0;
  assign f_u_dadda_pg_rca16_fa125_y2 = f_u_dadda_pg_rca16_fa125_y0 ^ f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_11_11_y0;
  assign f_u_dadda_pg_rca16_fa125_y3 = f_u_dadda_pg_rca16_fa125_y0 & f_u_dadda_pg_rca16_fa125_f_u_dadda_pg_rca16_and_11_11_y0;
  assign f_u_dadda_pg_rca16_fa125_y4 = f_u_dadda_pg_rca16_fa125_y1 | f_u_dadda_pg_rca16_fa125_y3;
  assign f_u_dadda_pg_rca16_and_10_12_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_10_12_y0 = f_u_dadda_pg_rca16_and_10_12_a_10 & f_u_dadda_pg_rca16_and_10_12_b_12;
  assign f_u_dadda_pg_rca16_and_9_13_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_9_13_y0 = f_u_dadda_pg_rca16_and_9_13_a_9 & f_u_dadda_pg_rca16_and_9_13_b_13;
  assign f_u_dadda_pg_rca16_and_8_14_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_8_14_y0 = f_u_dadda_pg_rca16_and_8_14_a_8 & f_u_dadda_pg_rca16_and_8_14_b_14;
  assign f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_10_12_y0 = f_u_dadda_pg_rca16_and_10_12_y0;
  assign f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_9_13_y0 = f_u_dadda_pg_rca16_and_9_13_y0;
  assign f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_8_14_y0 = f_u_dadda_pg_rca16_and_8_14_y0;
  assign f_u_dadda_pg_rca16_fa126_y0 = f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_10_12_y0 ^ f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_9_13_y0;
  assign f_u_dadda_pg_rca16_fa126_y1 = f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_10_12_y0 & f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_9_13_y0;
  assign f_u_dadda_pg_rca16_fa126_y2 = f_u_dadda_pg_rca16_fa126_y0 ^ f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_8_14_y0;
  assign f_u_dadda_pg_rca16_fa126_y3 = f_u_dadda_pg_rca16_fa126_y0 & f_u_dadda_pg_rca16_fa126_f_u_dadda_pg_rca16_and_8_14_y0;
  assign f_u_dadda_pg_rca16_fa126_y4 = f_u_dadda_pg_rca16_fa126_y1 | f_u_dadda_pg_rca16_fa126_y3;
  assign f_u_dadda_pg_rca16_and_7_15_a_7 = a_7;
  assign f_u_dadda_pg_rca16_and_7_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_7_15_y0 = f_u_dadda_pg_rca16_and_7_15_a_7 & f_u_dadda_pg_rca16_and_7_15_b_15;
  assign f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_and_7_15_y0 = f_u_dadda_pg_rca16_and_7_15_y0;
  assign f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_fa122_y2 = f_u_dadda_pg_rca16_fa122_y2;
  assign f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_fa123_y2 = f_u_dadda_pg_rca16_fa123_y2;
  assign f_u_dadda_pg_rca16_fa127_y0 = f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_and_7_15_y0 ^ f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_fa122_y2;
  assign f_u_dadda_pg_rca16_fa127_y1 = f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_and_7_15_y0 & f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_fa122_y2;
  assign f_u_dadda_pg_rca16_fa127_y2 = f_u_dadda_pg_rca16_fa127_y0 ^ f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_fa123_y2;
  assign f_u_dadda_pg_rca16_fa127_y3 = f_u_dadda_pg_rca16_fa127_y0 & f_u_dadda_pg_rca16_fa127_f_u_dadda_pg_rca16_fa123_y2;
  assign f_u_dadda_pg_rca16_fa127_y4 = f_u_dadda_pg_rca16_fa127_y1 | f_u_dadda_pg_rca16_fa127_y3;
  assign f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa127_y4 = f_u_dadda_pg_rca16_fa127_y4;
  assign f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa126_y4 = f_u_dadda_pg_rca16_fa126_y4;
  assign f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa125_y4 = f_u_dadda_pg_rca16_fa125_y4;
  assign f_u_dadda_pg_rca16_fa128_y0 = f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa127_y4 ^ f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa126_y4;
  assign f_u_dadda_pg_rca16_fa128_y1 = f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa127_y4 & f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa126_y4;
  assign f_u_dadda_pg_rca16_fa128_y2 = f_u_dadda_pg_rca16_fa128_y0 ^ f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa125_y4;
  assign f_u_dadda_pg_rca16_fa128_y3 = f_u_dadda_pg_rca16_fa128_y0 & f_u_dadda_pg_rca16_fa128_f_u_dadda_pg_rca16_fa125_y4;
  assign f_u_dadda_pg_rca16_fa128_y4 = f_u_dadda_pg_rca16_fa128_y1 | f_u_dadda_pg_rca16_fa128_y3;
  assign f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa124_y4 = f_u_dadda_pg_rca16_fa124_y4;
  assign f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa123_y4 = f_u_dadda_pg_rca16_fa123_y4;
  assign f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa122_y4 = f_u_dadda_pg_rca16_fa122_y4;
  assign f_u_dadda_pg_rca16_fa129_y0 = f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa124_y4 ^ f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa123_y4;
  assign f_u_dadda_pg_rca16_fa129_y1 = f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa124_y4 & f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa123_y4;
  assign f_u_dadda_pg_rca16_fa129_y2 = f_u_dadda_pg_rca16_fa129_y0 ^ f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa122_y4;
  assign f_u_dadda_pg_rca16_fa129_y3 = f_u_dadda_pg_rca16_fa129_y0 & f_u_dadda_pg_rca16_fa129_f_u_dadda_pg_rca16_fa122_y4;
  assign f_u_dadda_pg_rca16_fa129_y4 = f_u_dadda_pg_rca16_fa129_y1 | f_u_dadda_pg_rca16_fa129_y3;
  assign f_u_dadda_pg_rca16_and_15_8_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_8_b_8 = b_8;
  assign f_u_dadda_pg_rca16_and_15_8_y0 = f_u_dadda_pg_rca16_and_15_8_a_15 & f_u_dadda_pg_rca16_and_15_8_b_8;
  assign f_u_dadda_pg_rca16_and_14_9_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_14_9_y0 = f_u_dadda_pg_rca16_and_14_9_a_14 & f_u_dadda_pg_rca16_and_14_9_b_9;
  assign f_u_dadda_pg_rca16_and_13_10_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_13_10_y0 = f_u_dadda_pg_rca16_and_13_10_a_13 & f_u_dadda_pg_rca16_and_13_10_b_10;
  assign f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_15_8_y0 = f_u_dadda_pg_rca16_and_15_8_y0;
  assign f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_14_9_y0 = f_u_dadda_pg_rca16_and_14_9_y0;
  assign f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_13_10_y0 = f_u_dadda_pg_rca16_and_13_10_y0;
  assign f_u_dadda_pg_rca16_fa130_y0 = f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_15_8_y0 ^ f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_14_9_y0;
  assign f_u_dadda_pg_rca16_fa130_y1 = f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_15_8_y0 & f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_14_9_y0;
  assign f_u_dadda_pg_rca16_fa130_y2 = f_u_dadda_pg_rca16_fa130_y0 ^ f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_13_10_y0;
  assign f_u_dadda_pg_rca16_fa130_y3 = f_u_dadda_pg_rca16_fa130_y0 & f_u_dadda_pg_rca16_fa130_f_u_dadda_pg_rca16_and_13_10_y0;
  assign f_u_dadda_pg_rca16_fa130_y4 = f_u_dadda_pg_rca16_fa130_y1 | f_u_dadda_pg_rca16_fa130_y3;
  assign f_u_dadda_pg_rca16_and_12_11_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_12_11_y0 = f_u_dadda_pg_rca16_and_12_11_a_12 & f_u_dadda_pg_rca16_and_12_11_b_11;
  assign f_u_dadda_pg_rca16_and_11_12_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_11_12_y0 = f_u_dadda_pg_rca16_and_11_12_a_11 & f_u_dadda_pg_rca16_and_11_12_b_12;
  assign f_u_dadda_pg_rca16_and_10_13_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_10_13_y0 = f_u_dadda_pg_rca16_and_10_13_a_10 & f_u_dadda_pg_rca16_and_10_13_b_13;
  assign f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_12_11_y0 = f_u_dadda_pg_rca16_and_12_11_y0;
  assign f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_11_12_y0 = f_u_dadda_pg_rca16_and_11_12_y0;
  assign f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_10_13_y0 = f_u_dadda_pg_rca16_and_10_13_y0;
  assign f_u_dadda_pg_rca16_fa131_y0 = f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_12_11_y0 ^ f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_11_12_y0;
  assign f_u_dadda_pg_rca16_fa131_y1 = f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_12_11_y0 & f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_11_12_y0;
  assign f_u_dadda_pg_rca16_fa131_y2 = f_u_dadda_pg_rca16_fa131_y0 ^ f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_10_13_y0;
  assign f_u_dadda_pg_rca16_fa131_y3 = f_u_dadda_pg_rca16_fa131_y0 & f_u_dadda_pg_rca16_fa131_f_u_dadda_pg_rca16_and_10_13_y0;
  assign f_u_dadda_pg_rca16_fa131_y4 = f_u_dadda_pg_rca16_fa131_y1 | f_u_dadda_pg_rca16_fa131_y3;
  assign f_u_dadda_pg_rca16_and_9_14_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_9_14_y0 = f_u_dadda_pg_rca16_and_9_14_a_9 & f_u_dadda_pg_rca16_and_9_14_b_14;
  assign f_u_dadda_pg_rca16_and_8_15_a_8 = a_8;
  assign f_u_dadda_pg_rca16_and_8_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_8_15_y0 = f_u_dadda_pg_rca16_and_8_15_a_8 & f_u_dadda_pg_rca16_and_8_15_b_15;
  assign f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_and_9_14_y0 = f_u_dadda_pg_rca16_and_9_14_y0;
  assign f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_and_8_15_y0 = f_u_dadda_pg_rca16_and_8_15_y0;
  assign f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_fa128_y2 = f_u_dadda_pg_rca16_fa128_y2;
  assign f_u_dadda_pg_rca16_fa132_y0 = f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_and_9_14_y0 ^ f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_and_8_15_y0;
  assign f_u_dadda_pg_rca16_fa132_y1 = f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_and_9_14_y0 & f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_and_8_15_y0;
  assign f_u_dadda_pg_rca16_fa132_y2 = f_u_dadda_pg_rca16_fa132_y0 ^ f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_fa128_y2;
  assign f_u_dadda_pg_rca16_fa132_y3 = f_u_dadda_pg_rca16_fa132_y0 & f_u_dadda_pg_rca16_fa132_f_u_dadda_pg_rca16_fa128_y2;
  assign f_u_dadda_pg_rca16_fa132_y4 = f_u_dadda_pg_rca16_fa132_y1 | f_u_dadda_pg_rca16_fa132_y3;
  assign f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa132_y4 = f_u_dadda_pg_rca16_fa132_y4;
  assign f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa131_y4 = f_u_dadda_pg_rca16_fa131_y4;
  assign f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa130_y4 = f_u_dadda_pg_rca16_fa130_y4;
  assign f_u_dadda_pg_rca16_fa133_y0 = f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa132_y4 ^ f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa131_y4;
  assign f_u_dadda_pg_rca16_fa133_y1 = f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa132_y4 & f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa131_y4;
  assign f_u_dadda_pg_rca16_fa133_y2 = f_u_dadda_pg_rca16_fa133_y0 ^ f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa130_y4;
  assign f_u_dadda_pg_rca16_fa133_y3 = f_u_dadda_pg_rca16_fa133_y0 & f_u_dadda_pg_rca16_fa133_f_u_dadda_pg_rca16_fa130_y4;
  assign f_u_dadda_pg_rca16_fa133_y4 = f_u_dadda_pg_rca16_fa133_y1 | f_u_dadda_pg_rca16_fa133_y3;
  assign f_u_dadda_pg_rca16_and_15_9_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_9_b_9 = b_9;
  assign f_u_dadda_pg_rca16_and_15_9_y0 = f_u_dadda_pg_rca16_and_15_9_a_15 & f_u_dadda_pg_rca16_and_15_9_b_9;
  assign f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_fa129_y4 = f_u_dadda_pg_rca16_fa129_y4;
  assign f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_fa128_y4 = f_u_dadda_pg_rca16_fa128_y4;
  assign f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_and_15_9_y0 = f_u_dadda_pg_rca16_and_15_9_y0;
  assign f_u_dadda_pg_rca16_fa134_y0 = f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_fa129_y4 ^ f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_fa128_y4;
  assign f_u_dadda_pg_rca16_fa134_y1 = f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_fa129_y4 & f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_fa128_y4;
  assign f_u_dadda_pg_rca16_fa134_y2 = f_u_dadda_pg_rca16_fa134_y0 ^ f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_and_15_9_y0;
  assign f_u_dadda_pg_rca16_fa134_y3 = f_u_dadda_pg_rca16_fa134_y0 & f_u_dadda_pg_rca16_fa134_f_u_dadda_pg_rca16_and_15_9_y0;
  assign f_u_dadda_pg_rca16_fa134_y4 = f_u_dadda_pg_rca16_fa134_y1 | f_u_dadda_pg_rca16_fa134_y3;
  assign f_u_dadda_pg_rca16_and_14_10_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_14_10_y0 = f_u_dadda_pg_rca16_and_14_10_a_14 & f_u_dadda_pg_rca16_and_14_10_b_10;
  assign f_u_dadda_pg_rca16_and_13_11_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_13_11_y0 = f_u_dadda_pg_rca16_and_13_11_a_13 & f_u_dadda_pg_rca16_and_13_11_b_11;
  assign f_u_dadda_pg_rca16_and_12_12_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_12_12_y0 = f_u_dadda_pg_rca16_and_12_12_a_12 & f_u_dadda_pg_rca16_and_12_12_b_12;
  assign f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_14_10_y0 = f_u_dadda_pg_rca16_and_14_10_y0;
  assign f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_13_11_y0 = f_u_dadda_pg_rca16_and_13_11_y0;
  assign f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_12_12_y0 = f_u_dadda_pg_rca16_and_12_12_y0;
  assign f_u_dadda_pg_rca16_fa135_y0 = f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_14_10_y0 ^ f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_13_11_y0;
  assign f_u_dadda_pg_rca16_fa135_y1 = f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_14_10_y0 & f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_13_11_y0;
  assign f_u_dadda_pg_rca16_fa135_y2 = f_u_dadda_pg_rca16_fa135_y0 ^ f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_12_12_y0;
  assign f_u_dadda_pg_rca16_fa135_y3 = f_u_dadda_pg_rca16_fa135_y0 & f_u_dadda_pg_rca16_fa135_f_u_dadda_pg_rca16_and_12_12_y0;
  assign f_u_dadda_pg_rca16_fa135_y4 = f_u_dadda_pg_rca16_fa135_y1 | f_u_dadda_pg_rca16_fa135_y3;
  assign f_u_dadda_pg_rca16_and_11_13_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_11_13_y0 = f_u_dadda_pg_rca16_and_11_13_a_11 & f_u_dadda_pg_rca16_and_11_13_b_13;
  assign f_u_dadda_pg_rca16_and_10_14_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_10_14_y0 = f_u_dadda_pg_rca16_and_10_14_a_10 & f_u_dadda_pg_rca16_and_10_14_b_14;
  assign f_u_dadda_pg_rca16_and_9_15_a_9 = a_9;
  assign f_u_dadda_pg_rca16_and_9_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_9_15_y0 = f_u_dadda_pg_rca16_and_9_15_a_9 & f_u_dadda_pg_rca16_and_9_15_b_15;
  assign f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_11_13_y0 = f_u_dadda_pg_rca16_and_11_13_y0;
  assign f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_10_14_y0 = f_u_dadda_pg_rca16_and_10_14_y0;
  assign f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_9_15_y0 = f_u_dadda_pg_rca16_and_9_15_y0;
  assign f_u_dadda_pg_rca16_fa136_y0 = f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_11_13_y0 ^ f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_10_14_y0;
  assign f_u_dadda_pg_rca16_fa136_y1 = f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_11_13_y0 & f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_10_14_y0;
  assign f_u_dadda_pg_rca16_fa136_y2 = f_u_dadda_pg_rca16_fa136_y0 ^ f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_9_15_y0;
  assign f_u_dadda_pg_rca16_fa136_y3 = f_u_dadda_pg_rca16_fa136_y0 & f_u_dadda_pg_rca16_fa136_f_u_dadda_pg_rca16_and_9_15_y0;
  assign f_u_dadda_pg_rca16_fa136_y4 = f_u_dadda_pg_rca16_fa136_y1 | f_u_dadda_pg_rca16_fa136_y3;
  assign f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa136_y4 = f_u_dadda_pg_rca16_fa136_y4;
  assign f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa135_y4 = f_u_dadda_pg_rca16_fa135_y4;
  assign f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa134_y4 = f_u_dadda_pg_rca16_fa134_y4;
  assign f_u_dadda_pg_rca16_fa137_y0 = f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa136_y4 ^ f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa135_y4;
  assign f_u_dadda_pg_rca16_fa137_y1 = f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa136_y4 & f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa135_y4;
  assign f_u_dadda_pg_rca16_fa137_y2 = f_u_dadda_pg_rca16_fa137_y0 ^ f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa134_y4;
  assign f_u_dadda_pg_rca16_fa137_y3 = f_u_dadda_pg_rca16_fa137_y0 & f_u_dadda_pg_rca16_fa137_f_u_dadda_pg_rca16_fa134_y4;
  assign f_u_dadda_pg_rca16_fa137_y4 = f_u_dadda_pg_rca16_fa137_y1 | f_u_dadda_pg_rca16_fa137_y3;
  assign f_u_dadda_pg_rca16_and_15_10_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_10_b_10 = b_10;
  assign f_u_dadda_pg_rca16_and_15_10_y0 = f_u_dadda_pg_rca16_and_15_10_a_15 & f_u_dadda_pg_rca16_and_15_10_b_10;
  assign f_u_dadda_pg_rca16_and_14_11_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_14_11_y0 = f_u_dadda_pg_rca16_and_14_11_a_14 & f_u_dadda_pg_rca16_and_14_11_b_11;
  assign f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_fa133_y4 = f_u_dadda_pg_rca16_fa133_y4;
  assign f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_and_15_10_y0 = f_u_dadda_pg_rca16_and_15_10_y0;
  assign f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_and_14_11_y0 = f_u_dadda_pg_rca16_and_14_11_y0;
  assign f_u_dadda_pg_rca16_fa138_y0 = f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_fa133_y4 ^ f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_and_15_10_y0;
  assign f_u_dadda_pg_rca16_fa138_y1 = f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_fa133_y4 & f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_and_15_10_y0;
  assign f_u_dadda_pg_rca16_fa138_y2 = f_u_dadda_pg_rca16_fa138_y0 ^ f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_and_14_11_y0;
  assign f_u_dadda_pg_rca16_fa138_y3 = f_u_dadda_pg_rca16_fa138_y0 & f_u_dadda_pg_rca16_fa138_f_u_dadda_pg_rca16_and_14_11_y0;
  assign f_u_dadda_pg_rca16_fa138_y4 = f_u_dadda_pg_rca16_fa138_y1 | f_u_dadda_pg_rca16_fa138_y3;
  assign f_u_dadda_pg_rca16_and_13_12_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_13_12_y0 = f_u_dadda_pg_rca16_and_13_12_a_13 & f_u_dadda_pg_rca16_and_13_12_b_12;
  assign f_u_dadda_pg_rca16_and_12_13_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_12_13_y0 = f_u_dadda_pg_rca16_and_12_13_a_12 & f_u_dadda_pg_rca16_and_12_13_b_13;
  assign f_u_dadda_pg_rca16_and_11_14_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_11_14_y0 = f_u_dadda_pg_rca16_and_11_14_a_11 & f_u_dadda_pg_rca16_and_11_14_b_14;
  assign f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_13_12_y0 = f_u_dadda_pg_rca16_and_13_12_y0;
  assign f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_12_13_y0 = f_u_dadda_pg_rca16_and_12_13_y0;
  assign f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_11_14_y0 = f_u_dadda_pg_rca16_and_11_14_y0;
  assign f_u_dadda_pg_rca16_fa139_y0 = f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_13_12_y0 ^ f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_12_13_y0;
  assign f_u_dadda_pg_rca16_fa139_y1 = f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_13_12_y0 & f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_12_13_y0;
  assign f_u_dadda_pg_rca16_fa139_y2 = f_u_dadda_pg_rca16_fa139_y0 ^ f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_11_14_y0;
  assign f_u_dadda_pg_rca16_fa139_y3 = f_u_dadda_pg_rca16_fa139_y0 & f_u_dadda_pg_rca16_fa139_f_u_dadda_pg_rca16_and_11_14_y0;
  assign f_u_dadda_pg_rca16_fa139_y4 = f_u_dadda_pg_rca16_fa139_y1 | f_u_dadda_pg_rca16_fa139_y3;
  assign f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa139_y4 = f_u_dadda_pg_rca16_fa139_y4;
  assign f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa138_y4 = f_u_dadda_pg_rca16_fa138_y4;
  assign f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa137_y4 = f_u_dadda_pg_rca16_fa137_y4;
  assign f_u_dadda_pg_rca16_fa140_y0 = f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa139_y4 ^ f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa138_y4;
  assign f_u_dadda_pg_rca16_fa140_y1 = f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa139_y4 & f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa138_y4;
  assign f_u_dadda_pg_rca16_fa140_y2 = f_u_dadda_pg_rca16_fa140_y0 ^ f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa137_y4;
  assign f_u_dadda_pg_rca16_fa140_y3 = f_u_dadda_pg_rca16_fa140_y0 & f_u_dadda_pg_rca16_fa140_f_u_dadda_pg_rca16_fa137_y4;
  assign f_u_dadda_pg_rca16_fa140_y4 = f_u_dadda_pg_rca16_fa140_y1 | f_u_dadda_pg_rca16_fa140_y3;
  assign f_u_dadda_pg_rca16_and_15_11_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_11_b_11 = b_11;
  assign f_u_dadda_pg_rca16_and_15_11_y0 = f_u_dadda_pg_rca16_and_15_11_a_15 & f_u_dadda_pg_rca16_and_15_11_b_11;
  assign f_u_dadda_pg_rca16_and_14_12_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_14_12_y0 = f_u_dadda_pg_rca16_and_14_12_a_14 & f_u_dadda_pg_rca16_and_14_12_b_12;
  assign f_u_dadda_pg_rca16_and_13_13_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_13_13_y0 = f_u_dadda_pg_rca16_and_13_13_a_13 & f_u_dadda_pg_rca16_and_13_13_b_13;
  assign f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_15_11_y0 = f_u_dadda_pg_rca16_and_15_11_y0;
  assign f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_14_12_y0 = f_u_dadda_pg_rca16_and_14_12_y0;
  assign f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_13_13_y0 = f_u_dadda_pg_rca16_and_13_13_y0;
  assign f_u_dadda_pg_rca16_fa141_y0 = f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_15_11_y0 ^ f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_14_12_y0;
  assign f_u_dadda_pg_rca16_fa141_y1 = f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_15_11_y0 & f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_14_12_y0;
  assign f_u_dadda_pg_rca16_fa141_y2 = f_u_dadda_pg_rca16_fa141_y0 ^ f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_13_13_y0;
  assign f_u_dadda_pg_rca16_fa141_y3 = f_u_dadda_pg_rca16_fa141_y0 & f_u_dadda_pg_rca16_fa141_f_u_dadda_pg_rca16_and_13_13_y0;
  assign f_u_dadda_pg_rca16_fa141_y4 = f_u_dadda_pg_rca16_fa141_y1 | f_u_dadda_pg_rca16_fa141_y3;
  assign f_u_dadda_pg_rca16_and_15_12_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_12_b_12 = b_12;
  assign f_u_dadda_pg_rca16_and_15_12_y0 = f_u_dadda_pg_rca16_and_15_12_a_15 & f_u_dadda_pg_rca16_and_15_12_b_12;
  assign f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_fa141_y4 = f_u_dadda_pg_rca16_fa141_y4;
  assign f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_fa140_y4 = f_u_dadda_pg_rca16_fa140_y4;
  assign f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_and_15_12_y0 = f_u_dadda_pg_rca16_and_15_12_y0;
  assign f_u_dadda_pg_rca16_fa142_y0 = f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_fa141_y4 ^ f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_fa140_y4;
  assign f_u_dadda_pg_rca16_fa142_y1 = f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_fa141_y4 & f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_fa140_y4;
  assign f_u_dadda_pg_rca16_fa142_y2 = f_u_dadda_pg_rca16_fa142_y0 ^ f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_and_15_12_y0;
  assign f_u_dadda_pg_rca16_fa142_y3 = f_u_dadda_pg_rca16_fa142_y0 & f_u_dadda_pg_rca16_fa142_f_u_dadda_pg_rca16_and_15_12_y0;
  assign f_u_dadda_pg_rca16_fa142_y4 = f_u_dadda_pg_rca16_fa142_y1 | f_u_dadda_pg_rca16_fa142_y3;
  assign f_u_dadda_pg_rca16_and_3_0_a_3 = a_3;
  assign f_u_dadda_pg_rca16_and_3_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_3_0_y0 = f_u_dadda_pg_rca16_and_3_0_a_3 & f_u_dadda_pg_rca16_and_3_0_b_0;
  assign f_u_dadda_pg_rca16_and_2_1_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_2_1_y0 = f_u_dadda_pg_rca16_and_2_1_a_2 & f_u_dadda_pg_rca16_and_2_1_b_1;
  assign f_u_dadda_pg_rca16_ha13_f_u_dadda_pg_rca16_and_3_0_y0 = f_u_dadda_pg_rca16_and_3_0_y0;
  assign f_u_dadda_pg_rca16_ha13_f_u_dadda_pg_rca16_and_2_1_y0 = f_u_dadda_pg_rca16_and_2_1_y0;
  assign f_u_dadda_pg_rca16_ha13_y0 = f_u_dadda_pg_rca16_ha13_f_u_dadda_pg_rca16_and_3_0_y0 ^ f_u_dadda_pg_rca16_ha13_f_u_dadda_pg_rca16_and_2_1_y0;
  assign f_u_dadda_pg_rca16_ha13_y1 = f_u_dadda_pg_rca16_ha13_f_u_dadda_pg_rca16_and_3_0_y0 & f_u_dadda_pg_rca16_ha13_f_u_dadda_pg_rca16_and_2_1_y0;
  assign f_u_dadda_pg_rca16_and_2_2_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_2_2_y0 = f_u_dadda_pg_rca16_and_2_2_a_2 & f_u_dadda_pg_rca16_and_2_2_b_2;
  assign f_u_dadda_pg_rca16_and_1_3_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_1_3_y0 = f_u_dadda_pg_rca16_and_1_3_a_1 & f_u_dadda_pg_rca16_and_1_3_b_3;
  assign f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_ha13_y1 = f_u_dadda_pg_rca16_ha13_y1;
  assign f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_and_2_2_y0 = f_u_dadda_pg_rca16_and_2_2_y0;
  assign f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_and_1_3_y0 = f_u_dadda_pg_rca16_and_1_3_y0;
  assign f_u_dadda_pg_rca16_fa143_y0 = f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_ha13_y1 ^ f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_and_2_2_y0;
  assign f_u_dadda_pg_rca16_fa143_y1 = f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_ha13_y1 & f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_and_2_2_y0;
  assign f_u_dadda_pg_rca16_fa143_y2 = f_u_dadda_pg_rca16_fa143_y0 ^ f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_and_1_3_y0;
  assign f_u_dadda_pg_rca16_fa143_y3 = f_u_dadda_pg_rca16_fa143_y0 & f_u_dadda_pg_rca16_fa143_f_u_dadda_pg_rca16_and_1_3_y0;
  assign f_u_dadda_pg_rca16_fa143_y4 = f_u_dadda_pg_rca16_fa143_y1 | f_u_dadda_pg_rca16_fa143_y3;
  assign f_u_dadda_pg_rca16_and_1_4_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_1_4_y0 = f_u_dadda_pg_rca16_and_1_4_a_1 & f_u_dadda_pg_rca16_and_1_4_b_4;
  assign f_u_dadda_pg_rca16_and_0_5_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_5_b_5 = b_5;
  assign f_u_dadda_pg_rca16_and_0_5_y0 = f_u_dadda_pg_rca16_and_0_5_a_0 & f_u_dadda_pg_rca16_and_0_5_b_5;
  assign f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_fa143_y4 = f_u_dadda_pg_rca16_fa143_y4;
  assign f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_and_1_4_y0 = f_u_dadda_pg_rca16_and_1_4_y0;
  assign f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_and_0_5_y0 = f_u_dadda_pg_rca16_and_0_5_y0;
  assign f_u_dadda_pg_rca16_fa144_y0 = f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_fa143_y4 ^ f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_and_1_4_y0;
  assign f_u_dadda_pg_rca16_fa144_y1 = f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_fa143_y4 & f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_and_1_4_y0;
  assign f_u_dadda_pg_rca16_fa144_y2 = f_u_dadda_pg_rca16_fa144_y0 ^ f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_and_0_5_y0;
  assign f_u_dadda_pg_rca16_fa144_y3 = f_u_dadda_pg_rca16_fa144_y0 & f_u_dadda_pg_rca16_fa144_f_u_dadda_pg_rca16_and_0_5_y0;
  assign f_u_dadda_pg_rca16_fa144_y4 = f_u_dadda_pg_rca16_fa144_y1 | f_u_dadda_pg_rca16_fa144_y3;
  assign f_u_dadda_pg_rca16_and_0_6_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_6_b_6 = b_6;
  assign f_u_dadda_pg_rca16_and_0_6_y0 = f_u_dadda_pg_rca16_and_0_6_a_0 & f_u_dadda_pg_rca16_and_0_6_b_6;
  assign f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_fa144_y4 = f_u_dadda_pg_rca16_fa144_y4;
  assign f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_and_0_6_y0 = f_u_dadda_pg_rca16_and_0_6_y0;
  assign f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_fa9_y2 = f_u_dadda_pg_rca16_fa9_y2;
  assign f_u_dadda_pg_rca16_fa145_y0 = f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_fa144_y4 ^ f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_and_0_6_y0;
  assign f_u_dadda_pg_rca16_fa145_y1 = f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_fa144_y4 & f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_and_0_6_y0;
  assign f_u_dadda_pg_rca16_fa145_y2 = f_u_dadda_pg_rca16_fa145_y0 ^ f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_fa9_y2;
  assign f_u_dadda_pg_rca16_fa145_y3 = f_u_dadda_pg_rca16_fa145_y0 & f_u_dadda_pg_rca16_fa145_f_u_dadda_pg_rca16_fa9_y2;
  assign f_u_dadda_pg_rca16_fa145_y4 = f_u_dadda_pg_rca16_fa145_y1 | f_u_dadda_pg_rca16_fa145_y3;
  assign f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa145_y4 = f_u_dadda_pg_rca16_fa145_y4;
  assign f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa11_y2 = f_u_dadda_pg_rca16_fa11_y2;
  assign f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa12_y2 = f_u_dadda_pg_rca16_fa12_y2;
  assign f_u_dadda_pg_rca16_fa146_y0 = f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa145_y4 ^ f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa11_y2;
  assign f_u_dadda_pg_rca16_fa146_y1 = f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa145_y4 & f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa11_y2;
  assign f_u_dadda_pg_rca16_fa146_y2 = f_u_dadda_pg_rca16_fa146_y0 ^ f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa12_y2;
  assign f_u_dadda_pg_rca16_fa146_y3 = f_u_dadda_pg_rca16_fa146_y0 & f_u_dadda_pg_rca16_fa146_f_u_dadda_pg_rca16_fa12_y2;
  assign f_u_dadda_pg_rca16_fa146_y4 = f_u_dadda_pg_rca16_fa146_y1 | f_u_dadda_pg_rca16_fa146_y3;
  assign f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa146_y4 = f_u_dadda_pg_rca16_fa146_y4;
  assign f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa15_y2 = f_u_dadda_pg_rca16_fa15_y2;
  assign f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa16_y2 = f_u_dadda_pg_rca16_fa16_y2;
  assign f_u_dadda_pg_rca16_fa147_y0 = f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa146_y4 ^ f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa15_y2;
  assign f_u_dadda_pg_rca16_fa147_y1 = f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa146_y4 & f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa15_y2;
  assign f_u_dadda_pg_rca16_fa147_y2 = f_u_dadda_pg_rca16_fa147_y0 ^ f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa16_y2;
  assign f_u_dadda_pg_rca16_fa147_y3 = f_u_dadda_pg_rca16_fa147_y0 & f_u_dadda_pg_rca16_fa147_f_u_dadda_pg_rca16_fa16_y2;
  assign f_u_dadda_pg_rca16_fa147_y4 = f_u_dadda_pg_rca16_fa147_y1 | f_u_dadda_pg_rca16_fa147_y3;
  assign f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa147_y4 = f_u_dadda_pg_rca16_fa147_y4;
  assign f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa20_y2 = f_u_dadda_pg_rca16_fa20_y2;
  assign f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa21_y2 = f_u_dadda_pg_rca16_fa21_y2;
  assign f_u_dadda_pg_rca16_fa148_y0 = f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa147_y4 ^ f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa20_y2;
  assign f_u_dadda_pg_rca16_fa148_y1 = f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa147_y4 & f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa20_y2;
  assign f_u_dadda_pg_rca16_fa148_y2 = f_u_dadda_pg_rca16_fa148_y0 ^ f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa21_y2;
  assign f_u_dadda_pg_rca16_fa148_y3 = f_u_dadda_pg_rca16_fa148_y0 & f_u_dadda_pg_rca16_fa148_f_u_dadda_pg_rca16_fa21_y2;
  assign f_u_dadda_pg_rca16_fa148_y4 = f_u_dadda_pg_rca16_fa148_y1 | f_u_dadda_pg_rca16_fa148_y3;
  assign f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa148_y4 = f_u_dadda_pg_rca16_fa148_y4;
  assign f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa26_y2 = f_u_dadda_pg_rca16_fa26_y2;
  assign f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa27_y2 = f_u_dadda_pg_rca16_fa27_y2;
  assign f_u_dadda_pg_rca16_fa149_y0 = f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa148_y4 ^ f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa26_y2;
  assign f_u_dadda_pg_rca16_fa149_y1 = f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa148_y4 & f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa26_y2;
  assign f_u_dadda_pg_rca16_fa149_y2 = f_u_dadda_pg_rca16_fa149_y0 ^ f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa27_y2;
  assign f_u_dadda_pg_rca16_fa149_y3 = f_u_dadda_pg_rca16_fa149_y0 & f_u_dadda_pg_rca16_fa149_f_u_dadda_pg_rca16_fa27_y2;
  assign f_u_dadda_pg_rca16_fa149_y4 = f_u_dadda_pg_rca16_fa149_y1 | f_u_dadda_pg_rca16_fa149_y3;
  assign f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa149_y4 = f_u_dadda_pg_rca16_fa149_y4;
  assign f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa33_y2 = f_u_dadda_pg_rca16_fa33_y2;
  assign f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa34_y2 = f_u_dadda_pg_rca16_fa34_y2;
  assign f_u_dadda_pg_rca16_fa150_y0 = f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa149_y4 ^ f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa33_y2;
  assign f_u_dadda_pg_rca16_fa150_y1 = f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa149_y4 & f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa33_y2;
  assign f_u_dadda_pg_rca16_fa150_y2 = f_u_dadda_pg_rca16_fa150_y0 ^ f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa34_y2;
  assign f_u_dadda_pg_rca16_fa150_y3 = f_u_dadda_pg_rca16_fa150_y0 & f_u_dadda_pg_rca16_fa150_f_u_dadda_pg_rca16_fa34_y2;
  assign f_u_dadda_pg_rca16_fa150_y4 = f_u_dadda_pg_rca16_fa150_y1 | f_u_dadda_pg_rca16_fa150_y3;
  assign f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa150_y4 = f_u_dadda_pg_rca16_fa150_y4;
  assign f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa41_y2 = f_u_dadda_pg_rca16_fa41_y2;
  assign f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa42_y2 = f_u_dadda_pg_rca16_fa42_y2;
  assign f_u_dadda_pg_rca16_fa151_y0 = f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa150_y4 ^ f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa41_y2;
  assign f_u_dadda_pg_rca16_fa151_y1 = f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa150_y4 & f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa41_y2;
  assign f_u_dadda_pg_rca16_fa151_y2 = f_u_dadda_pg_rca16_fa151_y0 ^ f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa42_y2;
  assign f_u_dadda_pg_rca16_fa151_y3 = f_u_dadda_pg_rca16_fa151_y0 & f_u_dadda_pg_rca16_fa151_f_u_dadda_pg_rca16_fa42_y2;
  assign f_u_dadda_pg_rca16_fa151_y4 = f_u_dadda_pg_rca16_fa151_y1 | f_u_dadda_pg_rca16_fa151_y3;
  assign f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa151_y4 = f_u_dadda_pg_rca16_fa151_y4;
  assign f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa49_y2 = f_u_dadda_pg_rca16_fa49_y2;
  assign f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa50_y2 = f_u_dadda_pg_rca16_fa50_y2;
  assign f_u_dadda_pg_rca16_fa152_y0 = f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa151_y4 ^ f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa49_y2;
  assign f_u_dadda_pg_rca16_fa152_y1 = f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa151_y4 & f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa49_y2;
  assign f_u_dadda_pg_rca16_fa152_y2 = f_u_dadda_pg_rca16_fa152_y0 ^ f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa50_y2;
  assign f_u_dadda_pg_rca16_fa152_y3 = f_u_dadda_pg_rca16_fa152_y0 & f_u_dadda_pg_rca16_fa152_f_u_dadda_pg_rca16_fa50_y2;
  assign f_u_dadda_pg_rca16_fa152_y4 = f_u_dadda_pg_rca16_fa152_y1 | f_u_dadda_pg_rca16_fa152_y3;
  assign f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa152_y4 = f_u_dadda_pg_rca16_fa152_y4;
  assign f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa58_y2 = f_u_dadda_pg_rca16_fa58_y2;
  assign f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa59_y2 = f_u_dadda_pg_rca16_fa59_y2;
  assign f_u_dadda_pg_rca16_fa153_y0 = f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa152_y4 ^ f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa58_y2;
  assign f_u_dadda_pg_rca16_fa153_y1 = f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa152_y4 & f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa58_y2;
  assign f_u_dadda_pg_rca16_fa153_y2 = f_u_dadda_pg_rca16_fa153_y0 ^ f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa59_y2;
  assign f_u_dadda_pg_rca16_fa153_y3 = f_u_dadda_pg_rca16_fa153_y0 & f_u_dadda_pg_rca16_fa153_f_u_dadda_pg_rca16_fa59_y2;
  assign f_u_dadda_pg_rca16_fa153_y4 = f_u_dadda_pg_rca16_fa153_y1 | f_u_dadda_pg_rca16_fa153_y3;
  assign f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa153_y4 = f_u_dadda_pg_rca16_fa153_y4;
  assign f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa67_y2 = f_u_dadda_pg_rca16_fa67_y2;
  assign f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa68_y2 = f_u_dadda_pg_rca16_fa68_y2;
  assign f_u_dadda_pg_rca16_fa154_y0 = f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa153_y4 ^ f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa67_y2;
  assign f_u_dadda_pg_rca16_fa154_y1 = f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa153_y4 & f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa67_y2;
  assign f_u_dadda_pg_rca16_fa154_y2 = f_u_dadda_pg_rca16_fa154_y0 ^ f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa68_y2;
  assign f_u_dadda_pg_rca16_fa154_y3 = f_u_dadda_pg_rca16_fa154_y0 & f_u_dadda_pg_rca16_fa154_f_u_dadda_pg_rca16_fa68_y2;
  assign f_u_dadda_pg_rca16_fa154_y4 = f_u_dadda_pg_rca16_fa154_y1 | f_u_dadda_pg_rca16_fa154_y3;
  assign f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa154_y4 = f_u_dadda_pg_rca16_fa154_y4;
  assign f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa76_y2 = f_u_dadda_pg_rca16_fa76_y2;
  assign f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa77_y2 = f_u_dadda_pg_rca16_fa77_y2;
  assign f_u_dadda_pg_rca16_fa155_y0 = f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa154_y4 ^ f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa76_y2;
  assign f_u_dadda_pg_rca16_fa155_y1 = f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa154_y4 & f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa76_y2;
  assign f_u_dadda_pg_rca16_fa155_y2 = f_u_dadda_pg_rca16_fa155_y0 ^ f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa77_y2;
  assign f_u_dadda_pg_rca16_fa155_y3 = f_u_dadda_pg_rca16_fa155_y0 & f_u_dadda_pg_rca16_fa155_f_u_dadda_pg_rca16_fa77_y2;
  assign f_u_dadda_pg_rca16_fa155_y4 = f_u_dadda_pg_rca16_fa155_y1 | f_u_dadda_pg_rca16_fa155_y3;
  assign f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa155_y4 = f_u_dadda_pg_rca16_fa155_y4;
  assign f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa85_y2 = f_u_dadda_pg_rca16_fa85_y2;
  assign f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa86_y2 = f_u_dadda_pg_rca16_fa86_y2;
  assign f_u_dadda_pg_rca16_fa156_y0 = f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa155_y4 ^ f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa85_y2;
  assign f_u_dadda_pg_rca16_fa156_y1 = f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa155_y4 & f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa85_y2;
  assign f_u_dadda_pg_rca16_fa156_y2 = f_u_dadda_pg_rca16_fa156_y0 ^ f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa86_y2;
  assign f_u_dadda_pg_rca16_fa156_y3 = f_u_dadda_pg_rca16_fa156_y0 & f_u_dadda_pg_rca16_fa156_f_u_dadda_pg_rca16_fa86_y2;
  assign f_u_dadda_pg_rca16_fa156_y4 = f_u_dadda_pg_rca16_fa156_y1 | f_u_dadda_pg_rca16_fa156_y3;
  assign f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa156_y4 = f_u_dadda_pg_rca16_fa156_y4;
  assign f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa94_y2 = f_u_dadda_pg_rca16_fa94_y2;
  assign f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa95_y2 = f_u_dadda_pg_rca16_fa95_y2;
  assign f_u_dadda_pg_rca16_fa157_y0 = f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa156_y4 ^ f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa94_y2;
  assign f_u_dadda_pg_rca16_fa157_y1 = f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa156_y4 & f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa94_y2;
  assign f_u_dadda_pg_rca16_fa157_y2 = f_u_dadda_pg_rca16_fa157_y0 ^ f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa95_y2;
  assign f_u_dadda_pg_rca16_fa157_y3 = f_u_dadda_pg_rca16_fa157_y0 & f_u_dadda_pg_rca16_fa157_f_u_dadda_pg_rca16_fa95_y2;
  assign f_u_dadda_pg_rca16_fa157_y4 = f_u_dadda_pg_rca16_fa157_y1 | f_u_dadda_pg_rca16_fa157_y3;
  assign f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa157_y4 = f_u_dadda_pg_rca16_fa157_y4;
  assign f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa103_y2 = f_u_dadda_pg_rca16_fa103_y2;
  assign f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa104_y2 = f_u_dadda_pg_rca16_fa104_y2;
  assign f_u_dadda_pg_rca16_fa158_y0 = f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa157_y4 ^ f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa103_y2;
  assign f_u_dadda_pg_rca16_fa158_y1 = f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa157_y4 & f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa103_y2;
  assign f_u_dadda_pg_rca16_fa158_y2 = f_u_dadda_pg_rca16_fa158_y0 ^ f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa104_y2;
  assign f_u_dadda_pg_rca16_fa158_y3 = f_u_dadda_pg_rca16_fa158_y0 & f_u_dadda_pg_rca16_fa158_f_u_dadda_pg_rca16_fa104_y2;
  assign f_u_dadda_pg_rca16_fa158_y4 = f_u_dadda_pg_rca16_fa158_y1 | f_u_dadda_pg_rca16_fa158_y3;
  assign f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa158_y4 = f_u_dadda_pg_rca16_fa158_y4;
  assign f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa111_y2 = f_u_dadda_pg_rca16_fa111_y2;
  assign f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa112_y2 = f_u_dadda_pg_rca16_fa112_y2;
  assign f_u_dadda_pg_rca16_fa159_y0 = f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa158_y4 ^ f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa111_y2;
  assign f_u_dadda_pg_rca16_fa159_y1 = f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa158_y4 & f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa111_y2;
  assign f_u_dadda_pg_rca16_fa159_y2 = f_u_dadda_pg_rca16_fa159_y0 ^ f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa112_y2;
  assign f_u_dadda_pg_rca16_fa159_y3 = f_u_dadda_pg_rca16_fa159_y0 & f_u_dadda_pg_rca16_fa159_f_u_dadda_pg_rca16_fa112_y2;
  assign f_u_dadda_pg_rca16_fa159_y4 = f_u_dadda_pg_rca16_fa159_y1 | f_u_dadda_pg_rca16_fa159_y3;
  assign f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa159_y4 = f_u_dadda_pg_rca16_fa159_y4;
  assign f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa118_y2 = f_u_dadda_pg_rca16_fa118_y2;
  assign f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa119_y2 = f_u_dadda_pg_rca16_fa119_y2;
  assign f_u_dadda_pg_rca16_fa160_y0 = f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa159_y4 ^ f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa118_y2;
  assign f_u_dadda_pg_rca16_fa160_y1 = f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa159_y4 & f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa118_y2;
  assign f_u_dadda_pg_rca16_fa160_y2 = f_u_dadda_pg_rca16_fa160_y0 ^ f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa119_y2;
  assign f_u_dadda_pg_rca16_fa160_y3 = f_u_dadda_pg_rca16_fa160_y0 & f_u_dadda_pg_rca16_fa160_f_u_dadda_pg_rca16_fa119_y2;
  assign f_u_dadda_pg_rca16_fa160_y4 = f_u_dadda_pg_rca16_fa160_y1 | f_u_dadda_pg_rca16_fa160_y3;
  assign f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa160_y4 = f_u_dadda_pg_rca16_fa160_y4;
  assign f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa124_y2 = f_u_dadda_pg_rca16_fa124_y2;
  assign f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa125_y2 = f_u_dadda_pg_rca16_fa125_y2;
  assign f_u_dadda_pg_rca16_fa161_y0 = f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa160_y4 ^ f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa124_y2;
  assign f_u_dadda_pg_rca16_fa161_y1 = f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa160_y4 & f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa124_y2;
  assign f_u_dadda_pg_rca16_fa161_y2 = f_u_dadda_pg_rca16_fa161_y0 ^ f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa125_y2;
  assign f_u_dadda_pg_rca16_fa161_y3 = f_u_dadda_pg_rca16_fa161_y0 & f_u_dadda_pg_rca16_fa161_f_u_dadda_pg_rca16_fa125_y2;
  assign f_u_dadda_pg_rca16_fa161_y4 = f_u_dadda_pg_rca16_fa161_y1 | f_u_dadda_pg_rca16_fa161_y3;
  assign f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa161_y4 = f_u_dadda_pg_rca16_fa161_y4;
  assign f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa129_y2 = f_u_dadda_pg_rca16_fa129_y2;
  assign f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa130_y2 = f_u_dadda_pg_rca16_fa130_y2;
  assign f_u_dadda_pg_rca16_fa162_y0 = f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa161_y4 ^ f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa129_y2;
  assign f_u_dadda_pg_rca16_fa162_y1 = f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa161_y4 & f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa129_y2;
  assign f_u_dadda_pg_rca16_fa162_y2 = f_u_dadda_pg_rca16_fa162_y0 ^ f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa130_y2;
  assign f_u_dadda_pg_rca16_fa162_y3 = f_u_dadda_pg_rca16_fa162_y0 & f_u_dadda_pg_rca16_fa162_f_u_dadda_pg_rca16_fa130_y2;
  assign f_u_dadda_pg_rca16_fa162_y4 = f_u_dadda_pg_rca16_fa162_y1 | f_u_dadda_pg_rca16_fa162_y3;
  assign f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa162_y4 = f_u_dadda_pg_rca16_fa162_y4;
  assign f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa133_y2 = f_u_dadda_pg_rca16_fa133_y2;
  assign f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa134_y2 = f_u_dadda_pg_rca16_fa134_y2;
  assign f_u_dadda_pg_rca16_fa163_y0 = f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa162_y4 ^ f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa133_y2;
  assign f_u_dadda_pg_rca16_fa163_y1 = f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa162_y4 & f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa133_y2;
  assign f_u_dadda_pg_rca16_fa163_y2 = f_u_dadda_pg_rca16_fa163_y0 ^ f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa134_y2;
  assign f_u_dadda_pg_rca16_fa163_y3 = f_u_dadda_pg_rca16_fa163_y0 & f_u_dadda_pg_rca16_fa163_f_u_dadda_pg_rca16_fa134_y2;
  assign f_u_dadda_pg_rca16_fa163_y4 = f_u_dadda_pg_rca16_fa163_y1 | f_u_dadda_pg_rca16_fa163_y3;
  assign f_u_dadda_pg_rca16_and_10_15_a_10 = a_10;
  assign f_u_dadda_pg_rca16_and_10_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_10_15_y0 = f_u_dadda_pg_rca16_and_10_15_a_10 & f_u_dadda_pg_rca16_and_10_15_b_15;
  assign f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_fa163_y4 = f_u_dadda_pg_rca16_fa163_y4;
  assign f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_and_10_15_y0 = f_u_dadda_pg_rca16_and_10_15_y0;
  assign f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_fa137_y2 = f_u_dadda_pg_rca16_fa137_y2;
  assign f_u_dadda_pg_rca16_fa164_y0 = f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_fa163_y4 ^ f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_and_10_15_y0;
  assign f_u_dadda_pg_rca16_fa164_y1 = f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_fa163_y4 & f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_and_10_15_y0;
  assign f_u_dadda_pg_rca16_fa164_y2 = f_u_dadda_pg_rca16_fa164_y0 ^ f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_fa137_y2;
  assign f_u_dadda_pg_rca16_fa164_y3 = f_u_dadda_pg_rca16_fa164_y0 & f_u_dadda_pg_rca16_fa164_f_u_dadda_pg_rca16_fa137_y2;
  assign f_u_dadda_pg_rca16_fa164_y4 = f_u_dadda_pg_rca16_fa164_y1 | f_u_dadda_pg_rca16_fa164_y3;
  assign f_u_dadda_pg_rca16_and_12_14_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_12_14_y0 = f_u_dadda_pg_rca16_and_12_14_a_12 & f_u_dadda_pg_rca16_and_12_14_b_14;
  assign f_u_dadda_pg_rca16_and_11_15_a_11 = a_11;
  assign f_u_dadda_pg_rca16_and_11_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_11_15_y0 = f_u_dadda_pg_rca16_and_11_15_a_11 & f_u_dadda_pg_rca16_and_11_15_b_15;
  assign f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_fa164_y4 = f_u_dadda_pg_rca16_fa164_y4;
  assign f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_and_12_14_y0 = f_u_dadda_pg_rca16_and_12_14_y0;
  assign f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_and_11_15_y0 = f_u_dadda_pg_rca16_and_11_15_y0;
  assign f_u_dadda_pg_rca16_fa165_y0 = f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_fa164_y4 ^ f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_and_12_14_y0;
  assign f_u_dadda_pg_rca16_fa165_y1 = f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_fa164_y4 & f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_and_12_14_y0;
  assign f_u_dadda_pg_rca16_fa165_y2 = f_u_dadda_pg_rca16_fa165_y0 ^ f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_and_11_15_y0;
  assign f_u_dadda_pg_rca16_fa165_y3 = f_u_dadda_pg_rca16_fa165_y0 & f_u_dadda_pg_rca16_fa165_f_u_dadda_pg_rca16_and_11_15_y0;
  assign f_u_dadda_pg_rca16_fa165_y4 = f_u_dadda_pg_rca16_fa165_y1 | f_u_dadda_pg_rca16_fa165_y3;
  assign f_u_dadda_pg_rca16_and_14_13_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_14_13_y0 = f_u_dadda_pg_rca16_and_14_13_a_14 & f_u_dadda_pg_rca16_and_14_13_b_13;
  assign f_u_dadda_pg_rca16_and_13_14_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_13_14_y0 = f_u_dadda_pg_rca16_and_13_14_a_13 & f_u_dadda_pg_rca16_and_13_14_b_14;
  assign f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_fa165_y4 = f_u_dadda_pg_rca16_fa165_y4;
  assign f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_and_14_13_y0 = f_u_dadda_pg_rca16_and_14_13_y0;
  assign f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_and_13_14_y0 = f_u_dadda_pg_rca16_and_13_14_y0;
  assign f_u_dadda_pg_rca16_fa166_y0 = f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_fa165_y4 ^ f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_and_14_13_y0;
  assign f_u_dadda_pg_rca16_fa166_y1 = f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_fa165_y4 & f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_and_14_13_y0;
  assign f_u_dadda_pg_rca16_fa166_y2 = f_u_dadda_pg_rca16_fa166_y0 ^ f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_and_13_14_y0;
  assign f_u_dadda_pg_rca16_fa166_y3 = f_u_dadda_pg_rca16_fa166_y0 & f_u_dadda_pg_rca16_fa166_f_u_dadda_pg_rca16_and_13_14_y0;
  assign f_u_dadda_pg_rca16_fa166_y4 = f_u_dadda_pg_rca16_fa166_y1 | f_u_dadda_pg_rca16_fa166_y3;
  assign f_u_dadda_pg_rca16_and_15_13_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_13_b_13 = b_13;
  assign f_u_dadda_pg_rca16_and_15_13_y0 = f_u_dadda_pg_rca16_and_15_13_a_15 & f_u_dadda_pg_rca16_and_15_13_b_13;
  assign f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_fa166_y4 = f_u_dadda_pg_rca16_fa166_y4;
  assign f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_fa142_y4 = f_u_dadda_pg_rca16_fa142_y4;
  assign f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_and_15_13_y0 = f_u_dadda_pg_rca16_and_15_13_y0;
  assign f_u_dadda_pg_rca16_fa167_y0 = f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_fa166_y4 ^ f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_fa142_y4;
  assign f_u_dadda_pg_rca16_fa167_y1 = f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_fa166_y4 & f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_fa142_y4;
  assign f_u_dadda_pg_rca16_fa167_y2 = f_u_dadda_pg_rca16_fa167_y0 ^ f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_and_15_13_y0;
  assign f_u_dadda_pg_rca16_fa167_y3 = f_u_dadda_pg_rca16_fa167_y0 & f_u_dadda_pg_rca16_fa167_f_u_dadda_pg_rca16_and_15_13_y0;
  assign f_u_dadda_pg_rca16_fa167_y4 = f_u_dadda_pg_rca16_fa167_y1 | f_u_dadda_pg_rca16_fa167_y3;
  assign f_u_dadda_pg_rca16_and_2_0_a_2 = a_2;
  assign f_u_dadda_pg_rca16_and_2_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_2_0_y0 = f_u_dadda_pg_rca16_and_2_0_a_2 & f_u_dadda_pg_rca16_and_2_0_b_0;
  assign f_u_dadda_pg_rca16_and_1_1_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_1_1_y0 = f_u_dadda_pg_rca16_and_1_1_a_1 & f_u_dadda_pg_rca16_and_1_1_b_1;
  assign f_u_dadda_pg_rca16_ha14_f_u_dadda_pg_rca16_and_2_0_y0 = f_u_dadda_pg_rca16_and_2_0_y0;
  assign f_u_dadda_pg_rca16_ha14_f_u_dadda_pg_rca16_and_1_1_y0 = f_u_dadda_pg_rca16_and_1_1_y0;
  assign f_u_dadda_pg_rca16_ha14_y0 = f_u_dadda_pg_rca16_ha14_f_u_dadda_pg_rca16_and_2_0_y0 ^ f_u_dadda_pg_rca16_ha14_f_u_dadda_pg_rca16_and_1_1_y0;
  assign f_u_dadda_pg_rca16_ha14_y1 = f_u_dadda_pg_rca16_ha14_f_u_dadda_pg_rca16_and_2_0_y0 & f_u_dadda_pg_rca16_ha14_f_u_dadda_pg_rca16_and_1_1_y0;
  assign f_u_dadda_pg_rca16_and_1_2_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_1_2_y0 = f_u_dadda_pg_rca16_and_1_2_a_1 & f_u_dadda_pg_rca16_and_1_2_b_2;
  assign f_u_dadda_pg_rca16_and_0_3_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_3_b_3 = b_3;
  assign f_u_dadda_pg_rca16_and_0_3_y0 = f_u_dadda_pg_rca16_and_0_3_a_0 & f_u_dadda_pg_rca16_and_0_3_b_3;
  assign f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_ha14_y1 = f_u_dadda_pg_rca16_ha14_y1;
  assign f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_and_1_2_y0 = f_u_dadda_pg_rca16_and_1_2_y0;
  assign f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_and_0_3_y0 = f_u_dadda_pg_rca16_and_0_3_y0;
  assign f_u_dadda_pg_rca16_fa168_y0 = f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_ha14_y1 ^ f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_and_1_2_y0;
  assign f_u_dadda_pg_rca16_fa168_y1 = f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_ha14_y1 & f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_and_1_2_y0;
  assign f_u_dadda_pg_rca16_fa168_y2 = f_u_dadda_pg_rca16_fa168_y0 ^ f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_and_0_3_y0;
  assign f_u_dadda_pg_rca16_fa168_y3 = f_u_dadda_pg_rca16_fa168_y0 & f_u_dadda_pg_rca16_fa168_f_u_dadda_pg_rca16_and_0_3_y0;
  assign f_u_dadda_pg_rca16_fa168_y4 = f_u_dadda_pg_rca16_fa168_y1 | f_u_dadda_pg_rca16_fa168_y3;
  assign f_u_dadda_pg_rca16_and_0_4_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_4_b_4 = b_4;
  assign f_u_dadda_pg_rca16_and_0_4_y0 = f_u_dadda_pg_rca16_and_0_4_a_0 & f_u_dadda_pg_rca16_and_0_4_b_4;
  assign f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_fa168_y4 = f_u_dadda_pg_rca16_fa168_y4;
  assign f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_and_0_4_y0 = f_u_dadda_pg_rca16_and_0_4_y0;
  assign f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_ha4_y0 = f_u_dadda_pg_rca16_ha4_y0;
  assign f_u_dadda_pg_rca16_fa169_y0 = f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_fa168_y4 ^ f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_and_0_4_y0;
  assign f_u_dadda_pg_rca16_fa169_y1 = f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_fa168_y4 & f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_and_0_4_y0;
  assign f_u_dadda_pg_rca16_fa169_y2 = f_u_dadda_pg_rca16_fa169_y0 ^ f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_ha4_y0;
  assign f_u_dadda_pg_rca16_fa169_y3 = f_u_dadda_pg_rca16_fa169_y0 & f_u_dadda_pg_rca16_fa169_f_u_dadda_pg_rca16_ha4_y0;
  assign f_u_dadda_pg_rca16_fa169_y4 = f_u_dadda_pg_rca16_fa169_y1 | f_u_dadda_pg_rca16_fa169_y3;
  assign f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_fa169_y4 = f_u_dadda_pg_rca16_fa169_y4;
  assign f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_fa8_y2 = f_u_dadda_pg_rca16_fa8_y2;
  assign f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_ha5_y0 = f_u_dadda_pg_rca16_ha5_y0;
  assign f_u_dadda_pg_rca16_fa170_y0 = f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_fa169_y4 ^ f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_fa8_y2;
  assign f_u_dadda_pg_rca16_fa170_y1 = f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_fa169_y4 & f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_fa8_y2;
  assign f_u_dadda_pg_rca16_fa170_y2 = f_u_dadda_pg_rca16_fa170_y0 ^ f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_ha5_y0;
  assign f_u_dadda_pg_rca16_fa170_y3 = f_u_dadda_pg_rca16_fa170_y0 & f_u_dadda_pg_rca16_fa170_f_u_dadda_pg_rca16_ha5_y0;
  assign f_u_dadda_pg_rca16_fa170_y4 = f_u_dadda_pg_rca16_fa170_y1 | f_u_dadda_pg_rca16_fa170_y3;
  assign f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_fa170_y4 = f_u_dadda_pg_rca16_fa170_y4;
  assign f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_fa10_y2 = f_u_dadda_pg_rca16_fa10_y2;
  assign f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_ha6_y0 = f_u_dadda_pg_rca16_ha6_y0;
  assign f_u_dadda_pg_rca16_fa171_y0 = f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_fa170_y4 ^ f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_fa10_y2;
  assign f_u_dadda_pg_rca16_fa171_y1 = f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_fa170_y4 & f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_fa10_y2;
  assign f_u_dadda_pg_rca16_fa171_y2 = f_u_dadda_pg_rca16_fa171_y0 ^ f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_ha6_y0;
  assign f_u_dadda_pg_rca16_fa171_y3 = f_u_dadda_pg_rca16_fa171_y0 & f_u_dadda_pg_rca16_fa171_f_u_dadda_pg_rca16_ha6_y0;
  assign f_u_dadda_pg_rca16_fa171_y4 = f_u_dadda_pg_rca16_fa171_y1 | f_u_dadda_pg_rca16_fa171_y3;
  assign f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_fa171_y4 = f_u_dadda_pg_rca16_fa171_y4;
  assign f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_fa13_y2 = f_u_dadda_pg_rca16_fa13_y2;
  assign f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_ha7_y0 = f_u_dadda_pg_rca16_ha7_y0;
  assign f_u_dadda_pg_rca16_fa172_y0 = f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_fa171_y4 ^ f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_fa13_y2;
  assign f_u_dadda_pg_rca16_fa172_y1 = f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_fa171_y4 & f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_fa13_y2;
  assign f_u_dadda_pg_rca16_fa172_y2 = f_u_dadda_pg_rca16_fa172_y0 ^ f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_ha7_y0;
  assign f_u_dadda_pg_rca16_fa172_y3 = f_u_dadda_pg_rca16_fa172_y0 & f_u_dadda_pg_rca16_fa172_f_u_dadda_pg_rca16_ha7_y0;
  assign f_u_dadda_pg_rca16_fa172_y4 = f_u_dadda_pg_rca16_fa172_y1 | f_u_dadda_pg_rca16_fa172_y3;
  assign f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_fa172_y4 = f_u_dadda_pg_rca16_fa172_y4;
  assign f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_fa17_y2 = f_u_dadda_pg_rca16_fa17_y2;
  assign f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_ha8_y0 = f_u_dadda_pg_rca16_ha8_y0;
  assign f_u_dadda_pg_rca16_fa173_y0 = f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_fa172_y4 ^ f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_fa17_y2;
  assign f_u_dadda_pg_rca16_fa173_y1 = f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_fa172_y4 & f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_fa17_y2;
  assign f_u_dadda_pg_rca16_fa173_y2 = f_u_dadda_pg_rca16_fa173_y0 ^ f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_ha8_y0;
  assign f_u_dadda_pg_rca16_fa173_y3 = f_u_dadda_pg_rca16_fa173_y0 & f_u_dadda_pg_rca16_fa173_f_u_dadda_pg_rca16_ha8_y0;
  assign f_u_dadda_pg_rca16_fa173_y4 = f_u_dadda_pg_rca16_fa173_y1 | f_u_dadda_pg_rca16_fa173_y3;
  assign f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_fa173_y4 = f_u_dadda_pg_rca16_fa173_y4;
  assign f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_fa22_y2 = f_u_dadda_pg_rca16_fa22_y2;
  assign f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_ha9_y0 = f_u_dadda_pg_rca16_ha9_y0;
  assign f_u_dadda_pg_rca16_fa174_y0 = f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_fa173_y4 ^ f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_fa22_y2;
  assign f_u_dadda_pg_rca16_fa174_y1 = f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_fa173_y4 & f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_fa22_y2;
  assign f_u_dadda_pg_rca16_fa174_y2 = f_u_dadda_pg_rca16_fa174_y0 ^ f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_ha9_y0;
  assign f_u_dadda_pg_rca16_fa174_y3 = f_u_dadda_pg_rca16_fa174_y0 & f_u_dadda_pg_rca16_fa174_f_u_dadda_pg_rca16_ha9_y0;
  assign f_u_dadda_pg_rca16_fa174_y4 = f_u_dadda_pg_rca16_fa174_y1 | f_u_dadda_pg_rca16_fa174_y3;
  assign f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_fa174_y4 = f_u_dadda_pg_rca16_fa174_y4;
  assign f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_fa28_y2 = f_u_dadda_pg_rca16_fa28_y2;
  assign f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_ha10_y0 = f_u_dadda_pg_rca16_ha10_y0;
  assign f_u_dadda_pg_rca16_fa175_y0 = f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_fa174_y4 ^ f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_fa28_y2;
  assign f_u_dadda_pg_rca16_fa175_y1 = f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_fa174_y4 & f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_fa28_y2;
  assign f_u_dadda_pg_rca16_fa175_y2 = f_u_dadda_pg_rca16_fa175_y0 ^ f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_ha10_y0;
  assign f_u_dadda_pg_rca16_fa175_y3 = f_u_dadda_pg_rca16_fa175_y0 & f_u_dadda_pg_rca16_fa175_f_u_dadda_pg_rca16_ha10_y0;
  assign f_u_dadda_pg_rca16_fa175_y4 = f_u_dadda_pg_rca16_fa175_y1 | f_u_dadda_pg_rca16_fa175_y3;
  assign f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_fa175_y4 = f_u_dadda_pg_rca16_fa175_y4;
  assign f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_fa35_y2 = f_u_dadda_pg_rca16_fa35_y2;
  assign f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_ha11_y0 = f_u_dadda_pg_rca16_ha11_y0;
  assign f_u_dadda_pg_rca16_fa176_y0 = f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_fa175_y4 ^ f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_fa35_y2;
  assign f_u_dadda_pg_rca16_fa176_y1 = f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_fa175_y4 & f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_fa35_y2;
  assign f_u_dadda_pg_rca16_fa176_y2 = f_u_dadda_pg_rca16_fa176_y0 ^ f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_ha11_y0;
  assign f_u_dadda_pg_rca16_fa176_y3 = f_u_dadda_pg_rca16_fa176_y0 & f_u_dadda_pg_rca16_fa176_f_u_dadda_pg_rca16_ha11_y0;
  assign f_u_dadda_pg_rca16_fa176_y4 = f_u_dadda_pg_rca16_fa176_y1 | f_u_dadda_pg_rca16_fa176_y3;
  assign f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_fa176_y4 = f_u_dadda_pg_rca16_fa176_y4;
  assign f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_fa43_y2 = f_u_dadda_pg_rca16_fa43_y2;
  assign f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_ha12_y0 = f_u_dadda_pg_rca16_ha12_y0;
  assign f_u_dadda_pg_rca16_fa177_y0 = f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_fa176_y4 ^ f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_fa43_y2;
  assign f_u_dadda_pg_rca16_fa177_y1 = f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_fa176_y4 & f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_fa43_y2;
  assign f_u_dadda_pg_rca16_fa177_y2 = f_u_dadda_pg_rca16_fa177_y0 ^ f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_ha12_y0;
  assign f_u_dadda_pg_rca16_fa177_y3 = f_u_dadda_pg_rca16_fa177_y0 & f_u_dadda_pg_rca16_fa177_f_u_dadda_pg_rca16_ha12_y0;
  assign f_u_dadda_pg_rca16_fa177_y4 = f_u_dadda_pg_rca16_fa177_y1 | f_u_dadda_pg_rca16_fa177_y3;
  assign f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa177_y4 = f_u_dadda_pg_rca16_fa177_y4;
  assign f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa51_y2 = f_u_dadda_pg_rca16_fa51_y2;
  assign f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa52_y2 = f_u_dadda_pg_rca16_fa52_y2;
  assign f_u_dadda_pg_rca16_fa178_y0 = f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa177_y4 ^ f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa51_y2;
  assign f_u_dadda_pg_rca16_fa178_y1 = f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa177_y4 & f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa51_y2;
  assign f_u_dadda_pg_rca16_fa178_y2 = f_u_dadda_pg_rca16_fa178_y0 ^ f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa52_y2;
  assign f_u_dadda_pg_rca16_fa178_y3 = f_u_dadda_pg_rca16_fa178_y0 & f_u_dadda_pg_rca16_fa178_f_u_dadda_pg_rca16_fa52_y2;
  assign f_u_dadda_pg_rca16_fa178_y4 = f_u_dadda_pg_rca16_fa178_y1 | f_u_dadda_pg_rca16_fa178_y3;
  assign f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa178_y4 = f_u_dadda_pg_rca16_fa178_y4;
  assign f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa60_y2 = f_u_dadda_pg_rca16_fa60_y2;
  assign f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa61_y2 = f_u_dadda_pg_rca16_fa61_y2;
  assign f_u_dadda_pg_rca16_fa179_y0 = f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa178_y4 ^ f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa60_y2;
  assign f_u_dadda_pg_rca16_fa179_y1 = f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa178_y4 & f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa60_y2;
  assign f_u_dadda_pg_rca16_fa179_y2 = f_u_dadda_pg_rca16_fa179_y0 ^ f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa61_y2;
  assign f_u_dadda_pg_rca16_fa179_y3 = f_u_dadda_pg_rca16_fa179_y0 & f_u_dadda_pg_rca16_fa179_f_u_dadda_pg_rca16_fa61_y2;
  assign f_u_dadda_pg_rca16_fa179_y4 = f_u_dadda_pg_rca16_fa179_y1 | f_u_dadda_pg_rca16_fa179_y3;
  assign f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa179_y4 = f_u_dadda_pg_rca16_fa179_y4;
  assign f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa69_y2 = f_u_dadda_pg_rca16_fa69_y2;
  assign f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa70_y2 = f_u_dadda_pg_rca16_fa70_y2;
  assign f_u_dadda_pg_rca16_fa180_y0 = f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa179_y4 ^ f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa69_y2;
  assign f_u_dadda_pg_rca16_fa180_y1 = f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa179_y4 & f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa69_y2;
  assign f_u_dadda_pg_rca16_fa180_y2 = f_u_dadda_pg_rca16_fa180_y0 ^ f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa70_y2;
  assign f_u_dadda_pg_rca16_fa180_y3 = f_u_dadda_pg_rca16_fa180_y0 & f_u_dadda_pg_rca16_fa180_f_u_dadda_pg_rca16_fa70_y2;
  assign f_u_dadda_pg_rca16_fa180_y4 = f_u_dadda_pg_rca16_fa180_y1 | f_u_dadda_pg_rca16_fa180_y3;
  assign f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa180_y4 = f_u_dadda_pg_rca16_fa180_y4;
  assign f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa78_y2 = f_u_dadda_pg_rca16_fa78_y2;
  assign f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa79_y2 = f_u_dadda_pg_rca16_fa79_y2;
  assign f_u_dadda_pg_rca16_fa181_y0 = f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa180_y4 ^ f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa78_y2;
  assign f_u_dadda_pg_rca16_fa181_y1 = f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa180_y4 & f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa78_y2;
  assign f_u_dadda_pg_rca16_fa181_y2 = f_u_dadda_pg_rca16_fa181_y0 ^ f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa79_y2;
  assign f_u_dadda_pg_rca16_fa181_y3 = f_u_dadda_pg_rca16_fa181_y0 & f_u_dadda_pg_rca16_fa181_f_u_dadda_pg_rca16_fa79_y2;
  assign f_u_dadda_pg_rca16_fa181_y4 = f_u_dadda_pg_rca16_fa181_y1 | f_u_dadda_pg_rca16_fa181_y3;
  assign f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa181_y4 = f_u_dadda_pg_rca16_fa181_y4;
  assign f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa87_y2 = f_u_dadda_pg_rca16_fa87_y2;
  assign f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa88_y2 = f_u_dadda_pg_rca16_fa88_y2;
  assign f_u_dadda_pg_rca16_fa182_y0 = f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa181_y4 ^ f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa87_y2;
  assign f_u_dadda_pg_rca16_fa182_y1 = f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa181_y4 & f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa87_y2;
  assign f_u_dadda_pg_rca16_fa182_y2 = f_u_dadda_pg_rca16_fa182_y0 ^ f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa88_y2;
  assign f_u_dadda_pg_rca16_fa182_y3 = f_u_dadda_pg_rca16_fa182_y0 & f_u_dadda_pg_rca16_fa182_f_u_dadda_pg_rca16_fa88_y2;
  assign f_u_dadda_pg_rca16_fa182_y4 = f_u_dadda_pg_rca16_fa182_y1 | f_u_dadda_pg_rca16_fa182_y3;
  assign f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa182_y4 = f_u_dadda_pg_rca16_fa182_y4;
  assign f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa96_y2 = f_u_dadda_pg_rca16_fa96_y2;
  assign f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa97_y2 = f_u_dadda_pg_rca16_fa97_y2;
  assign f_u_dadda_pg_rca16_fa183_y0 = f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa182_y4 ^ f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa96_y2;
  assign f_u_dadda_pg_rca16_fa183_y1 = f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa182_y4 & f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa96_y2;
  assign f_u_dadda_pg_rca16_fa183_y2 = f_u_dadda_pg_rca16_fa183_y0 ^ f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa97_y2;
  assign f_u_dadda_pg_rca16_fa183_y3 = f_u_dadda_pg_rca16_fa183_y0 & f_u_dadda_pg_rca16_fa183_f_u_dadda_pg_rca16_fa97_y2;
  assign f_u_dadda_pg_rca16_fa183_y4 = f_u_dadda_pg_rca16_fa183_y1 | f_u_dadda_pg_rca16_fa183_y3;
  assign f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa183_y4 = f_u_dadda_pg_rca16_fa183_y4;
  assign f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa105_y2 = f_u_dadda_pg_rca16_fa105_y2;
  assign f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa106_y2 = f_u_dadda_pg_rca16_fa106_y2;
  assign f_u_dadda_pg_rca16_fa184_y0 = f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa183_y4 ^ f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa105_y2;
  assign f_u_dadda_pg_rca16_fa184_y1 = f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa183_y4 & f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa105_y2;
  assign f_u_dadda_pg_rca16_fa184_y2 = f_u_dadda_pg_rca16_fa184_y0 ^ f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa106_y2;
  assign f_u_dadda_pg_rca16_fa184_y3 = f_u_dadda_pg_rca16_fa184_y0 & f_u_dadda_pg_rca16_fa184_f_u_dadda_pg_rca16_fa106_y2;
  assign f_u_dadda_pg_rca16_fa184_y4 = f_u_dadda_pg_rca16_fa184_y1 | f_u_dadda_pg_rca16_fa184_y3;
  assign f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa184_y4 = f_u_dadda_pg_rca16_fa184_y4;
  assign f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa113_y2 = f_u_dadda_pg_rca16_fa113_y2;
  assign f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa114_y2 = f_u_dadda_pg_rca16_fa114_y2;
  assign f_u_dadda_pg_rca16_fa185_y0 = f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa184_y4 ^ f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa113_y2;
  assign f_u_dadda_pg_rca16_fa185_y1 = f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa184_y4 & f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa113_y2;
  assign f_u_dadda_pg_rca16_fa185_y2 = f_u_dadda_pg_rca16_fa185_y0 ^ f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa114_y2;
  assign f_u_dadda_pg_rca16_fa185_y3 = f_u_dadda_pg_rca16_fa185_y0 & f_u_dadda_pg_rca16_fa185_f_u_dadda_pg_rca16_fa114_y2;
  assign f_u_dadda_pg_rca16_fa185_y4 = f_u_dadda_pg_rca16_fa185_y1 | f_u_dadda_pg_rca16_fa185_y3;
  assign f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa185_y4 = f_u_dadda_pg_rca16_fa185_y4;
  assign f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa120_y2 = f_u_dadda_pg_rca16_fa120_y2;
  assign f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa121_y2 = f_u_dadda_pg_rca16_fa121_y2;
  assign f_u_dadda_pg_rca16_fa186_y0 = f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa185_y4 ^ f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa120_y2;
  assign f_u_dadda_pg_rca16_fa186_y1 = f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa185_y4 & f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa120_y2;
  assign f_u_dadda_pg_rca16_fa186_y2 = f_u_dadda_pg_rca16_fa186_y0 ^ f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa121_y2;
  assign f_u_dadda_pg_rca16_fa186_y3 = f_u_dadda_pg_rca16_fa186_y0 & f_u_dadda_pg_rca16_fa186_f_u_dadda_pg_rca16_fa121_y2;
  assign f_u_dadda_pg_rca16_fa186_y4 = f_u_dadda_pg_rca16_fa186_y1 | f_u_dadda_pg_rca16_fa186_y3;
  assign f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa186_y4 = f_u_dadda_pg_rca16_fa186_y4;
  assign f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa126_y2 = f_u_dadda_pg_rca16_fa126_y2;
  assign f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa127_y2 = f_u_dadda_pg_rca16_fa127_y2;
  assign f_u_dadda_pg_rca16_fa187_y0 = f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa186_y4 ^ f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa126_y2;
  assign f_u_dadda_pg_rca16_fa187_y1 = f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa186_y4 & f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa126_y2;
  assign f_u_dadda_pg_rca16_fa187_y2 = f_u_dadda_pg_rca16_fa187_y0 ^ f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa127_y2;
  assign f_u_dadda_pg_rca16_fa187_y3 = f_u_dadda_pg_rca16_fa187_y0 & f_u_dadda_pg_rca16_fa187_f_u_dadda_pg_rca16_fa127_y2;
  assign f_u_dadda_pg_rca16_fa187_y4 = f_u_dadda_pg_rca16_fa187_y1 | f_u_dadda_pg_rca16_fa187_y3;
  assign f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa187_y4 = f_u_dadda_pg_rca16_fa187_y4;
  assign f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa131_y2 = f_u_dadda_pg_rca16_fa131_y2;
  assign f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa132_y2 = f_u_dadda_pg_rca16_fa132_y2;
  assign f_u_dadda_pg_rca16_fa188_y0 = f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa187_y4 ^ f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa131_y2;
  assign f_u_dadda_pg_rca16_fa188_y1 = f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa187_y4 & f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa131_y2;
  assign f_u_dadda_pg_rca16_fa188_y2 = f_u_dadda_pg_rca16_fa188_y0 ^ f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa132_y2;
  assign f_u_dadda_pg_rca16_fa188_y3 = f_u_dadda_pg_rca16_fa188_y0 & f_u_dadda_pg_rca16_fa188_f_u_dadda_pg_rca16_fa132_y2;
  assign f_u_dadda_pg_rca16_fa188_y4 = f_u_dadda_pg_rca16_fa188_y1 | f_u_dadda_pg_rca16_fa188_y3;
  assign f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa188_y4 = f_u_dadda_pg_rca16_fa188_y4;
  assign f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa135_y2 = f_u_dadda_pg_rca16_fa135_y2;
  assign f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa136_y2 = f_u_dadda_pg_rca16_fa136_y2;
  assign f_u_dadda_pg_rca16_fa189_y0 = f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa188_y4 ^ f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa135_y2;
  assign f_u_dadda_pg_rca16_fa189_y1 = f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa188_y4 & f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa135_y2;
  assign f_u_dadda_pg_rca16_fa189_y2 = f_u_dadda_pg_rca16_fa189_y0 ^ f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa136_y2;
  assign f_u_dadda_pg_rca16_fa189_y3 = f_u_dadda_pg_rca16_fa189_y0 & f_u_dadda_pg_rca16_fa189_f_u_dadda_pg_rca16_fa136_y2;
  assign f_u_dadda_pg_rca16_fa189_y4 = f_u_dadda_pg_rca16_fa189_y1 | f_u_dadda_pg_rca16_fa189_y3;
  assign f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa189_y4 = f_u_dadda_pg_rca16_fa189_y4;
  assign f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa138_y2 = f_u_dadda_pg_rca16_fa138_y2;
  assign f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa139_y2 = f_u_dadda_pg_rca16_fa139_y2;
  assign f_u_dadda_pg_rca16_fa190_y0 = f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa189_y4 ^ f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa138_y2;
  assign f_u_dadda_pg_rca16_fa190_y1 = f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa189_y4 & f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa138_y2;
  assign f_u_dadda_pg_rca16_fa190_y2 = f_u_dadda_pg_rca16_fa190_y0 ^ f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa139_y2;
  assign f_u_dadda_pg_rca16_fa190_y3 = f_u_dadda_pg_rca16_fa190_y0 & f_u_dadda_pg_rca16_fa190_f_u_dadda_pg_rca16_fa139_y2;
  assign f_u_dadda_pg_rca16_fa190_y4 = f_u_dadda_pg_rca16_fa190_y1 | f_u_dadda_pg_rca16_fa190_y3;
  assign f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa190_y4 = f_u_dadda_pg_rca16_fa190_y4;
  assign f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa140_y2 = f_u_dadda_pg_rca16_fa140_y2;
  assign f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa141_y2 = f_u_dadda_pg_rca16_fa141_y2;
  assign f_u_dadda_pg_rca16_fa191_y0 = f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa190_y4 ^ f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa140_y2;
  assign f_u_dadda_pg_rca16_fa191_y1 = f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa190_y4 & f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa140_y2;
  assign f_u_dadda_pg_rca16_fa191_y2 = f_u_dadda_pg_rca16_fa191_y0 ^ f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa141_y2;
  assign f_u_dadda_pg_rca16_fa191_y3 = f_u_dadda_pg_rca16_fa191_y0 & f_u_dadda_pg_rca16_fa191_f_u_dadda_pg_rca16_fa141_y2;
  assign f_u_dadda_pg_rca16_fa191_y4 = f_u_dadda_pg_rca16_fa191_y1 | f_u_dadda_pg_rca16_fa191_y3;
  assign f_u_dadda_pg_rca16_and_12_15_a_12 = a_12;
  assign f_u_dadda_pg_rca16_and_12_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_12_15_y0 = f_u_dadda_pg_rca16_and_12_15_a_12 & f_u_dadda_pg_rca16_and_12_15_b_15;
  assign f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_fa191_y4 = f_u_dadda_pg_rca16_fa191_y4;
  assign f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_and_12_15_y0 = f_u_dadda_pg_rca16_and_12_15_y0;
  assign f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_fa142_y2 = f_u_dadda_pg_rca16_fa142_y2;
  assign f_u_dadda_pg_rca16_fa192_y0 = f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_fa191_y4 ^ f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_and_12_15_y0;
  assign f_u_dadda_pg_rca16_fa192_y1 = f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_fa191_y4 & f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_and_12_15_y0;
  assign f_u_dadda_pg_rca16_fa192_y2 = f_u_dadda_pg_rca16_fa192_y0 ^ f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_fa142_y2;
  assign f_u_dadda_pg_rca16_fa192_y3 = f_u_dadda_pg_rca16_fa192_y0 & f_u_dadda_pg_rca16_fa192_f_u_dadda_pg_rca16_fa142_y2;
  assign f_u_dadda_pg_rca16_fa192_y4 = f_u_dadda_pg_rca16_fa192_y1 | f_u_dadda_pg_rca16_fa192_y3;
  assign f_u_dadda_pg_rca16_and_14_14_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_14_14_y0 = f_u_dadda_pg_rca16_and_14_14_a_14 & f_u_dadda_pg_rca16_and_14_14_b_14;
  assign f_u_dadda_pg_rca16_and_13_15_a_13 = a_13;
  assign f_u_dadda_pg_rca16_and_13_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_13_15_y0 = f_u_dadda_pg_rca16_and_13_15_a_13 & f_u_dadda_pg_rca16_and_13_15_b_15;
  assign f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_fa192_y4 = f_u_dadda_pg_rca16_fa192_y4;
  assign f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_and_14_14_y0 = f_u_dadda_pg_rca16_and_14_14_y0;
  assign f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_and_13_15_y0 = f_u_dadda_pg_rca16_and_13_15_y0;
  assign f_u_dadda_pg_rca16_fa193_y0 = f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_fa192_y4 ^ f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_and_14_14_y0;
  assign f_u_dadda_pg_rca16_fa193_y1 = f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_fa192_y4 & f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_and_14_14_y0;
  assign f_u_dadda_pg_rca16_fa193_y2 = f_u_dadda_pg_rca16_fa193_y0 ^ f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_and_13_15_y0;
  assign f_u_dadda_pg_rca16_fa193_y3 = f_u_dadda_pg_rca16_fa193_y0 & f_u_dadda_pg_rca16_fa193_f_u_dadda_pg_rca16_and_13_15_y0;
  assign f_u_dadda_pg_rca16_fa193_y4 = f_u_dadda_pg_rca16_fa193_y1 | f_u_dadda_pg_rca16_fa193_y3;
  assign f_u_dadda_pg_rca16_and_15_14_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_14_b_14 = b_14;
  assign f_u_dadda_pg_rca16_and_15_14_y0 = f_u_dadda_pg_rca16_and_15_14_a_15 & f_u_dadda_pg_rca16_and_15_14_b_14;
  assign f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_fa193_y4 = f_u_dadda_pg_rca16_fa193_y4;
  assign f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_fa167_y4 = f_u_dadda_pg_rca16_fa167_y4;
  assign f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_and_15_14_y0 = f_u_dadda_pg_rca16_and_15_14_y0;
  assign f_u_dadda_pg_rca16_fa194_y0 = f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_fa193_y4 ^ f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_fa167_y4;
  assign f_u_dadda_pg_rca16_fa194_y1 = f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_fa193_y4 & f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_fa167_y4;
  assign f_u_dadda_pg_rca16_fa194_y2 = f_u_dadda_pg_rca16_fa194_y0 ^ f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_and_15_14_y0;
  assign f_u_dadda_pg_rca16_fa194_y3 = f_u_dadda_pg_rca16_fa194_y0 & f_u_dadda_pg_rca16_fa194_f_u_dadda_pg_rca16_and_15_14_y0;
  assign f_u_dadda_pg_rca16_fa194_y4 = f_u_dadda_pg_rca16_fa194_y1 | f_u_dadda_pg_rca16_fa194_y3;
  assign f_u_dadda_pg_rca16_and_0_0_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_0_0_y0 = f_u_dadda_pg_rca16_and_0_0_a_0 & f_u_dadda_pg_rca16_and_0_0_b_0;
  assign f_u_dadda_pg_rca16_and_1_0_a_1 = a_1;
  assign f_u_dadda_pg_rca16_and_1_0_b_0 = b_0;
  assign f_u_dadda_pg_rca16_and_1_0_y0 = f_u_dadda_pg_rca16_and_1_0_a_1 & f_u_dadda_pg_rca16_and_1_0_b_0;
  assign f_u_dadda_pg_rca16_and_0_2_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_2_b_2 = b_2;
  assign f_u_dadda_pg_rca16_and_0_2_y0 = f_u_dadda_pg_rca16_and_0_2_a_0 & f_u_dadda_pg_rca16_and_0_2_b_2;
  assign f_u_dadda_pg_rca16_and_14_15_a_14 = a_14;
  assign f_u_dadda_pg_rca16_and_14_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_14_15_y0 = f_u_dadda_pg_rca16_and_14_15_a_14 & f_u_dadda_pg_rca16_and_14_15_b_15;
  assign f_u_dadda_pg_rca16_and_0_1_a_0 = a_0;
  assign f_u_dadda_pg_rca16_and_0_1_b_1 = b_1;
  assign f_u_dadda_pg_rca16_and_0_1_y0 = f_u_dadda_pg_rca16_and_0_1_a_0 & f_u_dadda_pg_rca16_and_0_1_b_1;
  assign f_u_dadda_pg_rca16_and_15_15_a_15 = a_15;
  assign f_u_dadda_pg_rca16_and_15_15_b_15 = b_15;
  assign f_u_dadda_pg_rca16_and_15_15_y0 = f_u_dadda_pg_rca16_and_15_15_a_15 & f_u_dadda_pg_rca16_and_15_15_b_15;
  assign constant_wire_value_0_f_u_dadda_pg_rca16_and_1_0_y0 = f_u_dadda_pg_rca16_and_1_0_y0;
  assign constant_wire_value_0_f_u_dadda_pg_rca16_and_0_1_y0 = f_u_dadda_pg_rca16_and_0_1_y0;
  assign constant_wire_value_0_y0 = constant_wire_value_0_f_u_dadda_pg_rca16_and_1_0_y0 ^ constant_wire_value_0_f_u_dadda_pg_rca16_and_0_1_y0;
  assign constant_wire_value_0_y1 = ~(constant_wire_value_0_f_u_dadda_pg_rca16_and_1_0_y0 ^ constant_wire_value_0_f_u_dadda_pg_rca16_and_0_1_y0);
  assign constant_wire_0 = ~(constant_wire_value_0_y0 | constant_wire_value_0_y1);
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa0_f_u_dadda_pg_rca16_and_1_0_y0 = f_u_dadda_pg_rca16_and_1_0_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa0_f_u_dadda_pg_rca16_and_0_1_y0 = f_u_dadda_pg_rca16_and_0_1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa0_constant_wire_0 = constant_wire_0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa0_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa0_f_u_dadda_pg_rca16_and_1_0_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa0_f_u_dadda_pg_rca16_and_0_1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa0_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa0_f_u_dadda_pg_rca16_and_1_0_y0 & f_u_dadda_pg_rca16_u_pg_rca30_fa0_f_u_dadda_pg_rca16_and_0_1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa0_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa0_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa0_constant_wire_0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and0_constant_wire_0 = constant_wire_0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and0_f_u_dadda_pg_rca16_u_pg_rca30_fa0_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa0_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and0_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and0_constant_wire_0 & f_u_dadda_pg_rca16_u_pg_rca30_and0_f_u_dadda_pg_rca16_u_pg_rca30_fa0_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or0_f_u_dadda_pg_rca16_u_pg_rca30_and0_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and0_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or0_f_u_dadda_pg_rca16_u_pg_rca30_fa0_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa0_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or0_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or0_f_u_dadda_pg_rca16_u_pg_rca30_and0_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or0_f_u_dadda_pg_rca16_u_pg_rca30_fa0_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_and_0_2_y0 = f_u_dadda_pg_rca16_and_0_2_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_ha14_y0 = f_u_dadda_pg_rca16_ha14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_u_pg_rca30_or0_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or0_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa1_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_and_0_2_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_ha14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa1_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_and_0_2_y0 & f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_ha14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa1_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa1_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa1_f_u_dadda_pg_rca16_u_pg_rca30_or0_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and1_f_u_dadda_pg_rca16_u_pg_rca30_or0_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or0_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and1_f_u_dadda_pg_rca16_u_pg_rca30_fa1_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and1_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and1_f_u_dadda_pg_rca16_u_pg_rca30_or0_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and1_f_u_dadda_pg_rca16_u_pg_rca30_fa1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or1_f_u_dadda_pg_rca16_u_pg_rca30_and1_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or1_f_u_dadda_pg_rca16_u_pg_rca30_fa1_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa1_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or1_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or1_f_u_dadda_pg_rca16_u_pg_rca30_and1_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or1_f_u_dadda_pg_rca16_u_pg_rca30_fa1_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_ha13_y0 = f_u_dadda_pg_rca16_ha13_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_fa168_y2 = f_u_dadda_pg_rca16_fa168_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_u_pg_rca30_or1_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa2_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_ha13_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_fa168_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa2_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_ha13_y0 & f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_fa168_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa2_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa2_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa2_f_u_dadda_pg_rca16_u_pg_rca30_or1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and2_f_u_dadda_pg_rca16_u_pg_rca30_or1_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or1_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and2_f_u_dadda_pg_rca16_u_pg_rca30_fa2_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa2_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and2_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and2_f_u_dadda_pg_rca16_u_pg_rca30_or1_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and2_f_u_dadda_pg_rca16_u_pg_rca30_fa2_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or2_f_u_dadda_pg_rca16_u_pg_rca30_and2_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and2_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or2_f_u_dadda_pg_rca16_u_pg_rca30_fa2_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa2_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or2_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or2_f_u_dadda_pg_rca16_u_pg_rca30_and2_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or2_f_u_dadda_pg_rca16_u_pg_rca30_fa2_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_fa143_y2 = f_u_dadda_pg_rca16_fa143_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_fa169_y2 = f_u_dadda_pg_rca16_fa169_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_u_pg_rca30_or2_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or2_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa3_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_fa143_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_fa169_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa3_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_fa143_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_fa169_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa3_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa3_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa3_f_u_dadda_pg_rca16_u_pg_rca30_or2_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and3_f_u_dadda_pg_rca16_u_pg_rca30_or2_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or2_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and3_f_u_dadda_pg_rca16_u_pg_rca30_fa3_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa3_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and3_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and3_f_u_dadda_pg_rca16_u_pg_rca30_or2_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and3_f_u_dadda_pg_rca16_u_pg_rca30_fa3_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or3_f_u_dadda_pg_rca16_u_pg_rca30_and3_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and3_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or3_f_u_dadda_pg_rca16_u_pg_rca30_fa3_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa3_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or3_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or3_f_u_dadda_pg_rca16_u_pg_rca30_and3_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or3_f_u_dadda_pg_rca16_u_pg_rca30_fa3_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_fa144_y2 = f_u_dadda_pg_rca16_fa144_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_fa170_y2 = f_u_dadda_pg_rca16_fa170_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_u_pg_rca30_or3_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or3_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa4_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_fa144_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_fa170_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa4_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_fa144_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_fa170_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa4_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa4_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa4_f_u_dadda_pg_rca16_u_pg_rca30_or3_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and4_f_u_dadda_pg_rca16_u_pg_rca30_or3_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or3_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and4_f_u_dadda_pg_rca16_u_pg_rca30_fa4_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa4_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and4_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and4_f_u_dadda_pg_rca16_u_pg_rca30_or3_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and4_f_u_dadda_pg_rca16_u_pg_rca30_fa4_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or4_f_u_dadda_pg_rca16_u_pg_rca30_and4_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and4_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or4_f_u_dadda_pg_rca16_u_pg_rca30_fa4_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa4_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or4_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or4_f_u_dadda_pg_rca16_u_pg_rca30_and4_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or4_f_u_dadda_pg_rca16_u_pg_rca30_fa4_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_fa145_y2 = f_u_dadda_pg_rca16_fa145_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_fa171_y2 = f_u_dadda_pg_rca16_fa171_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_u_pg_rca30_or4_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or4_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa5_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_fa145_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_fa171_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa5_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_fa145_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_fa171_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa5_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa5_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa5_f_u_dadda_pg_rca16_u_pg_rca30_or4_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and5_f_u_dadda_pg_rca16_u_pg_rca30_or4_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or4_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and5_f_u_dadda_pg_rca16_u_pg_rca30_fa5_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa5_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and5_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and5_f_u_dadda_pg_rca16_u_pg_rca30_or4_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and5_f_u_dadda_pg_rca16_u_pg_rca30_fa5_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or5_f_u_dadda_pg_rca16_u_pg_rca30_and5_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and5_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or5_f_u_dadda_pg_rca16_u_pg_rca30_fa5_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa5_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or5_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or5_f_u_dadda_pg_rca16_u_pg_rca30_and5_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or5_f_u_dadda_pg_rca16_u_pg_rca30_fa5_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_fa146_y2 = f_u_dadda_pg_rca16_fa146_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_fa172_y2 = f_u_dadda_pg_rca16_fa172_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_u_pg_rca30_or5_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or5_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa6_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_fa146_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_fa172_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa6_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_fa146_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_fa172_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa6_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa6_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa6_f_u_dadda_pg_rca16_u_pg_rca30_or5_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and6_f_u_dadda_pg_rca16_u_pg_rca30_or5_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or5_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and6_f_u_dadda_pg_rca16_u_pg_rca30_fa6_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa6_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and6_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and6_f_u_dadda_pg_rca16_u_pg_rca30_or5_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and6_f_u_dadda_pg_rca16_u_pg_rca30_fa6_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or6_f_u_dadda_pg_rca16_u_pg_rca30_and6_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and6_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or6_f_u_dadda_pg_rca16_u_pg_rca30_fa6_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa6_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or6_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or6_f_u_dadda_pg_rca16_u_pg_rca30_and6_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or6_f_u_dadda_pg_rca16_u_pg_rca30_fa6_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_fa147_y2 = f_u_dadda_pg_rca16_fa147_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_fa173_y2 = f_u_dadda_pg_rca16_fa173_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_u_pg_rca30_or6_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or6_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa7_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_fa147_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_fa173_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa7_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_fa147_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_fa173_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa7_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa7_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa7_f_u_dadda_pg_rca16_u_pg_rca30_or6_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and7_f_u_dadda_pg_rca16_u_pg_rca30_or6_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or6_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and7_f_u_dadda_pg_rca16_u_pg_rca30_fa7_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa7_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and7_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and7_f_u_dadda_pg_rca16_u_pg_rca30_or6_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and7_f_u_dadda_pg_rca16_u_pg_rca30_fa7_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or7_f_u_dadda_pg_rca16_u_pg_rca30_and7_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and7_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or7_f_u_dadda_pg_rca16_u_pg_rca30_fa7_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa7_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or7_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or7_f_u_dadda_pg_rca16_u_pg_rca30_and7_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or7_f_u_dadda_pg_rca16_u_pg_rca30_fa7_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_fa148_y2 = f_u_dadda_pg_rca16_fa148_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_fa174_y2 = f_u_dadda_pg_rca16_fa174_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_u_pg_rca30_or7_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or7_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa8_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_fa148_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_fa174_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa8_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_fa148_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_fa174_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa8_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa8_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa8_f_u_dadda_pg_rca16_u_pg_rca30_or7_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and8_f_u_dadda_pg_rca16_u_pg_rca30_or7_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or7_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and8_f_u_dadda_pg_rca16_u_pg_rca30_fa8_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa8_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and8_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and8_f_u_dadda_pg_rca16_u_pg_rca30_or7_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and8_f_u_dadda_pg_rca16_u_pg_rca30_fa8_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or8_f_u_dadda_pg_rca16_u_pg_rca30_and8_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and8_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or8_f_u_dadda_pg_rca16_u_pg_rca30_fa8_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa8_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or8_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or8_f_u_dadda_pg_rca16_u_pg_rca30_and8_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or8_f_u_dadda_pg_rca16_u_pg_rca30_fa8_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_fa149_y2 = f_u_dadda_pg_rca16_fa149_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_fa175_y2 = f_u_dadda_pg_rca16_fa175_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_u_pg_rca30_or8_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or8_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa9_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_fa149_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_fa175_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa9_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_fa149_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_fa175_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa9_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa9_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa9_f_u_dadda_pg_rca16_u_pg_rca30_or8_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and9_f_u_dadda_pg_rca16_u_pg_rca30_or8_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or8_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and9_f_u_dadda_pg_rca16_u_pg_rca30_fa9_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa9_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and9_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and9_f_u_dadda_pg_rca16_u_pg_rca30_or8_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and9_f_u_dadda_pg_rca16_u_pg_rca30_fa9_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or9_f_u_dadda_pg_rca16_u_pg_rca30_and9_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and9_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or9_f_u_dadda_pg_rca16_u_pg_rca30_fa9_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa9_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or9_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or9_f_u_dadda_pg_rca16_u_pg_rca30_and9_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or9_f_u_dadda_pg_rca16_u_pg_rca30_fa9_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_fa150_y2 = f_u_dadda_pg_rca16_fa150_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_fa176_y2 = f_u_dadda_pg_rca16_fa176_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_u_pg_rca30_or9_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or9_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa10_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_fa150_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_fa176_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa10_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_fa150_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_fa176_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa10_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa10_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa10_f_u_dadda_pg_rca16_u_pg_rca30_or9_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and10_f_u_dadda_pg_rca16_u_pg_rca30_or9_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or9_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and10_f_u_dadda_pg_rca16_u_pg_rca30_fa10_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa10_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and10_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and10_f_u_dadda_pg_rca16_u_pg_rca30_or9_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and10_f_u_dadda_pg_rca16_u_pg_rca30_fa10_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or10_f_u_dadda_pg_rca16_u_pg_rca30_and10_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and10_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or10_f_u_dadda_pg_rca16_u_pg_rca30_fa10_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa10_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or10_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or10_f_u_dadda_pg_rca16_u_pg_rca30_and10_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or10_f_u_dadda_pg_rca16_u_pg_rca30_fa10_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_fa151_y2 = f_u_dadda_pg_rca16_fa151_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_fa177_y2 = f_u_dadda_pg_rca16_fa177_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_u_pg_rca30_or10_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or10_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa11_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_fa151_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_fa177_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa11_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_fa151_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_fa177_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa11_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa11_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa11_f_u_dadda_pg_rca16_u_pg_rca30_or10_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and11_f_u_dadda_pg_rca16_u_pg_rca30_or10_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or10_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and11_f_u_dadda_pg_rca16_u_pg_rca30_fa11_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa11_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and11_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and11_f_u_dadda_pg_rca16_u_pg_rca30_or10_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and11_f_u_dadda_pg_rca16_u_pg_rca30_fa11_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or11_f_u_dadda_pg_rca16_u_pg_rca30_and11_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and11_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or11_f_u_dadda_pg_rca16_u_pg_rca30_fa11_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa11_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or11_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or11_f_u_dadda_pg_rca16_u_pg_rca30_and11_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or11_f_u_dadda_pg_rca16_u_pg_rca30_fa11_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_fa152_y2 = f_u_dadda_pg_rca16_fa152_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_fa178_y2 = f_u_dadda_pg_rca16_fa178_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_u_pg_rca30_or11_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or11_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa12_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_fa152_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_fa178_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa12_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_fa152_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_fa178_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa12_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa12_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa12_f_u_dadda_pg_rca16_u_pg_rca30_or11_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and12_f_u_dadda_pg_rca16_u_pg_rca30_or11_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or11_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and12_f_u_dadda_pg_rca16_u_pg_rca30_fa12_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa12_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and12_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and12_f_u_dadda_pg_rca16_u_pg_rca30_or11_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and12_f_u_dadda_pg_rca16_u_pg_rca30_fa12_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or12_f_u_dadda_pg_rca16_u_pg_rca30_and12_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and12_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or12_f_u_dadda_pg_rca16_u_pg_rca30_fa12_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa12_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or12_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or12_f_u_dadda_pg_rca16_u_pg_rca30_and12_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or12_f_u_dadda_pg_rca16_u_pg_rca30_fa12_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_fa153_y2 = f_u_dadda_pg_rca16_fa153_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_fa179_y2 = f_u_dadda_pg_rca16_fa179_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_u_pg_rca30_or12_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or12_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa13_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_fa153_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_fa179_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa13_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_fa153_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_fa179_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa13_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa13_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa13_f_u_dadda_pg_rca16_u_pg_rca30_or12_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and13_f_u_dadda_pg_rca16_u_pg_rca30_or12_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or12_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and13_f_u_dadda_pg_rca16_u_pg_rca30_fa13_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa13_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and13_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and13_f_u_dadda_pg_rca16_u_pg_rca30_or12_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and13_f_u_dadda_pg_rca16_u_pg_rca30_fa13_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or13_f_u_dadda_pg_rca16_u_pg_rca30_and13_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and13_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or13_f_u_dadda_pg_rca16_u_pg_rca30_fa13_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa13_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or13_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or13_f_u_dadda_pg_rca16_u_pg_rca30_and13_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or13_f_u_dadda_pg_rca16_u_pg_rca30_fa13_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_fa154_y2 = f_u_dadda_pg_rca16_fa154_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_fa180_y2 = f_u_dadda_pg_rca16_fa180_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_u_pg_rca30_or13_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or13_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa14_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_fa154_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_fa180_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa14_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_fa154_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_fa180_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa14_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa14_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa14_f_u_dadda_pg_rca16_u_pg_rca30_or13_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and14_f_u_dadda_pg_rca16_u_pg_rca30_or13_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or13_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and14_f_u_dadda_pg_rca16_u_pg_rca30_fa14_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and14_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and14_f_u_dadda_pg_rca16_u_pg_rca30_or13_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and14_f_u_dadda_pg_rca16_u_pg_rca30_fa14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or14_f_u_dadda_pg_rca16_u_pg_rca30_and14_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or14_f_u_dadda_pg_rca16_u_pg_rca30_fa14_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa14_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or14_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or14_f_u_dadda_pg_rca16_u_pg_rca30_and14_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or14_f_u_dadda_pg_rca16_u_pg_rca30_fa14_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_fa155_y2 = f_u_dadda_pg_rca16_fa155_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_fa181_y2 = f_u_dadda_pg_rca16_fa181_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_u_pg_rca30_or14_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa15_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_fa155_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_fa181_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa15_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_fa155_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_fa181_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa15_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa15_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa15_f_u_dadda_pg_rca16_u_pg_rca30_or14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and15_f_u_dadda_pg_rca16_u_pg_rca30_or14_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or14_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and15_f_u_dadda_pg_rca16_u_pg_rca30_fa15_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and15_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and15_f_u_dadda_pg_rca16_u_pg_rca30_or14_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and15_f_u_dadda_pg_rca16_u_pg_rca30_fa15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or15_f_u_dadda_pg_rca16_u_pg_rca30_and15_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or15_f_u_dadda_pg_rca16_u_pg_rca30_fa15_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa15_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or15_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or15_f_u_dadda_pg_rca16_u_pg_rca30_and15_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or15_f_u_dadda_pg_rca16_u_pg_rca30_fa15_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_fa156_y2 = f_u_dadda_pg_rca16_fa156_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_fa182_y2 = f_u_dadda_pg_rca16_fa182_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_u_pg_rca30_or15_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa16_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_fa156_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_fa182_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa16_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_fa156_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_fa182_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa16_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa16_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa16_f_u_dadda_pg_rca16_u_pg_rca30_or15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and16_f_u_dadda_pg_rca16_u_pg_rca30_or15_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and16_f_u_dadda_pg_rca16_u_pg_rca30_fa16_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa16_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and16_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and16_f_u_dadda_pg_rca16_u_pg_rca30_or15_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and16_f_u_dadda_pg_rca16_u_pg_rca30_fa16_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or16_f_u_dadda_pg_rca16_u_pg_rca30_and16_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and16_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or16_f_u_dadda_pg_rca16_u_pg_rca30_fa16_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa16_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or16_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or16_f_u_dadda_pg_rca16_u_pg_rca30_and16_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or16_f_u_dadda_pg_rca16_u_pg_rca30_fa16_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_fa157_y2 = f_u_dadda_pg_rca16_fa157_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_fa183_y2 = f_u_dadda_pg_rca16_fa183_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_u_pg_rca30_or16_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or16_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa17_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_fa157_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_fa183_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa17_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_fa157_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_fa183_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa17_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa17_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa17_f_u_dadda_pg_rca16_u_pg_rca30_or16_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and17_f_u_dadda_pg_rca16_u_pg_rca30_or16_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or16_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and17_f_u_dadda_pg_rca16_u_pg_rca30_fa17_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa17_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and17_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and17_f_u_dadda_pg_rca16_u_pg_rca30_or16_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and17_f_u_dadda_pg_rca16_u_pg_rca30_fa17_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or17_f_u_dadda_pg_rca16_u_pg_rca30_and17_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and17_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or17_f_u_dadda_pg_rca16_u_pg_rca30_fa17_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa17_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or17_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or17_f_u_dadda_pg_rca16_u_pg_rca30_and17_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or17_f_u_dadda_pg_rca16_u_pg_rca30_fa17_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_fa158_y2 = f_u_dadda_pg_rca16_fa158_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_fa184_y2 = f_u_dadda_pg_rca16_fa184_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_u_pg_rca30_or17_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or17_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa18_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_fa158_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_fa184_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa18_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_fa158_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_fa184_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa18_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa18_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa18_f_u_dadda_pg_rca16_u_pg_rca30_or17_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and18_f_u_dadda_pg_rca16_u_pg_rca30_or17_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or17_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and18_f_u_dadda_pg_rca16_u_pg_rca30_fa18_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa18_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and18_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and18_f_u_dadda_pg_rca16_u_pg_rca30_or17_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and18_f_u_dadda_pg_rca16_u_pg_rca30_fa18_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or18_f_u_dadda_pg_rca16_u_pg_rca30_and18_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and18_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or18_f_u_dadda_pg_rca16_u_pg_rca30_fa18_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa18_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or18_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or18_f_u_dadda_pg_rca16_u_pg_rca30_and18_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or18_f_u_dadda_pg_rca16_u_pg_rca30_fa18_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_fa159_y2 = f_u_dadda_pg_rca16_fa159_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_fa185_y2 = f_u_dadda_pg_rca16_fa185_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_u_pg_rca30_or18_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or18_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa19_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_fa159_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_fa185_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa19_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_fa159_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_fa185_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa19_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa19_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa19_f_u_dadda_pg_rca16_u_pg_rca30_or18_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and19_f_u_dadda_pg_rca16_u_pg_rca30_or18_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or18_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and19_f_u_dadda_pg_rca16_u_pg_rca30_fa19_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa19_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and19_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and19_f_u_dadda_pg_rca16_u_pg_rca30_or18_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and19_f_u_dadda_pg_rca16_u_pg_rca30_fa19_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or19_f_u_dadda_pg_rca16_u_pg_rca30_and19_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and19_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or19_f_u_dadda_pg_rca16_u_pg_rca30_fa19_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa19_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or19_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or19_f_u_dadda_pg_rca16_u_pg_rca30_and19_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or19_f_u_dadda_pg_rca16_u_pg_rca30_fa19_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_fa160_y2 = f_u_dadda_pg_rca16_fa160_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_fa186_y2 = f_u_dadda_pg_rca16_fa186_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_u_pg_rca30_or19_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or19_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa20_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_fa160_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_fa186_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa20_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_fa160_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_fa186_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa20_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa20_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa20_f_u_dadda_pg_rca16_u_pg_rca30_or19_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and20_f_u_dadda_pg_rca16_u_pg_rca30_or19_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or19_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and20_f_u_dadda_pg_rca16_u_pg_rca30_fa20_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa20_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and20_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and20_f_u_dadda_pg_rca16_u_pg_rca30_or19_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and20_f_u_dadda_pg_rca16_u_pg_rca30_fa20_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or20_f_u_dadda_pg_rca16_u_pg_rca30_and20_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and20_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or20_f_u_dadda_pg_rca16_u_pg_rca30_fa20_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa20_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or20_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or20_f_u_dadda_pg_rca16_u_pg_rca30_and20_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or20_f_u_dadda_pg_rca16_u_pg_rca30_fa20_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_fa161_y2 = f_u_dadda_pg_rca16_fa161_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_fa187_y2 = f_u_dadda_pg_rca16_fa187_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_u_pg_rca30_or20_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or20_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa21_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_fa161_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_fa187_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa21_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_fa161_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_fa187_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa21_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa21_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa21_f_u_dadda_pg_rca16_u_pg_rca30_or20_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and21_f_u_dadda_pg_rca16_u_pg_rca30_or20_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or20_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and21_f_u_dadda_pg_rca16_u_pg_rca30_fa21_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa21_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and21_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and21_f_u_dadda_pg_rca16_u_pg_rca30_or20_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and21_f_u_dadda_pg_rca16_u_pg_rca30_fa21_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or21_f_u_dadda_pg_rca16_u_pg_rca30_and21_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and21_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or21_f_u_dadda_pg_rca16_u_pg_rca30_fa21_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa21_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or21_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or21_f_u_dadda_pg_rca16_u_pg_rca30_and21_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or21_f_u_dadda_pg_rca16_u_pg_rca30_fa21_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_fa162_y2 = f_u_dadda_pg_rca16_fa162_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_fa188_y2 = f_u_dadda_pg_rca16_fa188_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_u_pg_rca30_or21_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or21_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa22_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_fa162_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_fa188_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa22_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_fa162_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_fa188_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa22_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa22_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa22_f_u_dadda_pg_rca16_u_pg_rca30_or21_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and22_f_u_dadda_pg_rca16_u_pg_rca30_or21_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or21_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and22_f_u_dadda_pg_rca16_u_pg_rca30_fa22_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa22_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and22_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and22_f_u_dadda_pg_rca16_u_pg_rca30_or21_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and22_f_u_dadda_pg_rca16_u_pg_rca30_fa22_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or22_f_u_dadda_pg_rca16_u_pg_rca30_and22_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and22_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or22_f_u_dadda_pg_rca16_u_pg_rca30_fa22_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa22_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or22_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or22_f_u_dadda_pg_rca16_u_pg_rca30_and22_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or22_f_u_dadda_pg_rca16_u_pg_rca30_fa22_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_fa163_y2 = f_u_dadda_pg_rca16_fa163_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_fa189_y2 = f_u_dadda_pg_rca16_fa189_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_u_pg_rca30_or22_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or22_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa23_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_fa163_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_fa189_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa23_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_fa163_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_fa189_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa23_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa23_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa23_f_u_dadda_pg_rca16_u_pg_rca30_or22_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and23_f_u_dadda_pg_rca16_u_pg_rca30_or22_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or22_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and23_f_u_dadda_pg_rca16_u_pg_rca30_fa23_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa23_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and23_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and23_f_u_dadda_pg_rca16_u_pg_rca30_or22_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and23_f_u_dadda_pg_rca16_u_pg_rca30_fa23_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or23_f_u_dadda_pg_rca16_u_pg_rca30_and23_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and23_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or23_f_u_dadda_pg_rca16_u_pg_rca30_fa23_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa23_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or23_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or23_f_u_dadda_pg_rca16_u_pg_rca30_and23_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or23_f_u_dadda_pg_rca16_u_pg_rca30_fa23_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_fa164_y2 = f_u_dadda_pg_rca16_fa164_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_fa190_y2 = f_u_dadda_pg_rca16_fa190_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_u_pg_rca30_or23_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or23_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa24_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_fa164_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_fa190_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa24_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_fa164_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_fa190_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa24_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa24_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa24_f_u_dadda_pg_rca16_u_pg_rca30_or23_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and24_f_u_dadda_pg_rca16_u_pg_rca30_or23_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or23_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and24_f_u_dadda_pg_rca16_u_pg_rca30_fa24_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa24_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and24_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and24_f_u_dadda_pg_rca16_u_pg_rca30_or23_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and24_f_u_dadda_pg_rca16_u_pg_rca30_fa24_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or24_f_u_dadda_pg_rca16_u_pg_rca30_and24_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and24_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or24_f_u_dadda_pg_rca16_u_pg_rca30_fa24_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa24_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or24_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or24_f_u_dadda_pg_rca16_u_pg_rca30_and24_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or24_f_u_dadda_pg_rca16_u_pg_rca30_fa24_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_fa165_y2 = f_u_dadda_pg_rca16_fa165_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_fa191_y2 = f_u_dadda_pg_rca16_fa191_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_u_pg_rca30_or24_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or24_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa25_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_fa165_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_fa191_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa25_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_fa165_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_fa191_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa25_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa25_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa25_f_u_dadda_pg_rca16_u_pg_rca30_or24_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and25_f_u_dadda_pg_rca16_u_pg_rca30_or24_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or24_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and25_f_u_dadda_pg_rca16_u_pg_rca30_fa25_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa25_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and25_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and25_f_u_dadda_pg_rca16_u_pg_rca30_or24_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and25_f_u_dadda_pg_rca16_u_pg_rca30_fa25_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or25_f_u_dadda_pg_rca16_u_pg_rca30_and25_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and25_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or25_f_u_dadda_pg_rca16_u_pg_rca30_fa25_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa25_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or25_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or25_f_u_dadda_pg_rca16_u_pg_rca30_and25_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or25_f_u_dadda_pg_rca16_u_pg_rca30_fa25_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_fa166_y2 = f_u_dadda_pg_rca16_fa166_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_fa192_y2 = f_u_dadda_pg_rca16_fa192_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_u_pg_rca30_or25_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or25_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa26_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_fa166_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_fa192_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa26_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_fa166_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_fa192_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa26_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa26_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa26_f_u_dadda_pg_rca16_u_pg_rca30_or25_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and26_f_u_dadda_pg_rca16_u_pg_rca30_or25_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or25_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and26_f_u_dadda_pg_rca16_u_pg_rca30_fa26_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa26_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and26_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and26_f_u_dadda_pg_rca16_u_pg_rca30_or25_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and26_f_u_dadda_pg_rca16_u_pg_rca30_fa26_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or26_f_u_dadda_pg_rca16_u_pg_rca30_and26_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and26_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or26_f_u_dadda_pg_rca16_u_pg_rca30_fa26_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa26_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or26_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or26_f_u_dadda_pg_rca16_u_pg_rca30_and26_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or26_f_u_dadda_pg_rca16_u_pg_rca30_fa26_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_fa167_y2 = f_u_dadda_pg_rca16_fa167_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_fa193_y2 = f_u_dadda_pg_rca16_fa193_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_u_pg_rca30_or26_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or26_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa27_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_fa167_y2 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_fa193_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa27_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_fa167_y2 & f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_fa193_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa27_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa27_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa27_f_u_dadda_pg_rca16_u_pg_rca30_or26_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and27_f_u_dadda_pg_rca16_u_pg_rca30_or26_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or26_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and27_f_u_dadda_pg_rca16_u_pg_rca30_fa27_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa27_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and27_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and27_f_u_dadda_pg_rca16_u_pg_rca30_or26_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and27_f_u_dadda_pg_rca16_u_pg_rca30_fa27_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or27_f_u_dadda_pg_rca16_u_pg_rca30_and27_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and27_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or27_f_u_dadda_pg_rca16_u_pg_rca30_fa27_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa27_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or27_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or27_f_u_dadda_pg_rca16_u_pg_rca30_and27_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or27_f_u_dadda_pg_rca16_u_pg_rca30_fa27_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_and_14_15_y0 = f_u_dadda_pg_rca16_and_14_15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_fa194_y2 = f_u_dadda_pg_rca16_fa194_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_u_pg_rca30_or27_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or27_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa28_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_and_14_15_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_fa194_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa28_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_and_14_15_y0 & f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_fa194_y2;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa28_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa28_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa28_f_u_dadda_pg_rca16_u_pg_rca30_or27_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and28_f_u_dadda_pg_rca16_u_pg_rca30_or27_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or27_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and28_f_u_dadda_pg_rca16_u_pg_rca30_fa28_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa28_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and28_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and28_f_u_dadda_pg_rca16_u_pg_rca30_or27_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and28_f_u_dadda_pg_rca16_u_pg_rca30_fa28_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or28_f_u_dadda_pg_rca16_u_pg_rca30_and28_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and28_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or28_f_u_dadda_pg_rca16_u_pg_rca30_fa28_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa28_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or28_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or28_f_u_dadda_pg_rca16_u_pg_rca30_and28_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or28_f_u_dadda_pg_rca16_u_pg_rca30_fa28_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_fa194_y4 = f_u_dadda_pg_rca16_fa194_y4;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_and_15_15_y0 = f_u_dadda_pg_rca16_and_15_15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_u_pg_rca30_or28_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or28_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa29_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_fa194_y4 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_and_15_15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa29_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_fa194_y4 & f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_and_15_15_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_fa29_y2 = f_u_dadda_pg_rca16_u_pg_rca30_fa29_y0 ^ f_u_dadda_pg_rca16_u_pg_rca30_fa29_f_u_dadda_pg_rca16_u_pg_rca30_or28_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and29_f_u_dadda_pg_rca16_u_pg_rca30_or28_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or28_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and29_f_u_dadda_pg_rca16_u_pg_rca30_fa29_y0 = f_u_dadda_pg_rca16_u_pg_rca30_fa29_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_and29_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and29_f_u_dadda_pg_rca16_u_pg_rca30_or28_y0 & f_u_dadda_pg_rca16_u_pg_rca30_and29_f_u_dadda_pg_rca16_u_pg_rca30_fa29_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or29_f_u_dadda_pg_rca16_u_pg_rca30_and29_y0 = f_u_dadda_pg_rca16_u_pg_rca30_and29_y0;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or29_f_u_dadda_pg_rca16_u_pg_rca30_fa29_y1 = f_u_dadda_pg_rca16_u_pg_rca30_fa29_y1;
  assign f_u_dadda_pg_rca16_u_pg_rca30_or29_y0 = f_u_dadda_pg_rca16_u_pg_rca30_or29_f_u_dadda_pg_rca16_u_pg_rca30_and29_y0 | f_u_dadda_pg_rca16_u_pg_rca30_or29_f_u_dadda_pg_rca16_u_pg_rca30_fa29_y1;

  assign out[0] = f_u_dadda_pg_rca16_and_0_0_y0;
  assign out[1] = f_u_dadda_pg_rca16_u_pg_rca30_fa0_y2;
  assign out[2] = f_u_dadda_pg_rca16_u_pg_rca30_fa1_y2;
  assign out[3] = f_u_dadda_pg_rca16_u_pg_rca30_fa2_y2;
  assign out[4] = f_u_dadda_pg_rca16_u_pg_rca30_fa3_y2;
  assign out[5] = f_u_dadda_pg_rca16_u_pg_rca30_fa4_y2;
  assign out[6] = f_u_dadda_pg_rca16_u_pg_rca30_fa5_y2;
  assign out[7] = f_u_dadda_pg_rca16_u_pg_rca30_fa6_y2;
  assign out[8] = f_u_dadda_pg_rca16_u_pg_rca30_fa7_y2;
  assign out[9] = f_u_dadda_pg_rca16_u_pg_rca30_fa8_y2;
  assign out[10] = f_u_dadda_pg_rca16_u_pg_rca30_fa9_y2;
  assign out[11] = f_u_dadda_pg_rca16_u_pg_rca30_fa10_y2;
  assign out[12] = f_u_dadda_pg_rca16_u_pg_rca30_fa11_y2;
  assign out[13] = f_u_dadda_pg_rca16_u_pg_rca30_fa12_y2;
  assign out[14] = f_u_dadda_pg_rca16_u_pg_rca30_fa13_y2;
  assign out[15] = f_u_dadda_pg_rca16_u_pg_rca30_fa14_y2;
  assign out[16] = f_u_dadda_pg_rca16_u_pg_rca30_fa15_y2;
  assign out[17] = f_u_dadda_pg_rca16_u_pg_rca30_fa16_y2;
  assign out[18] = f_u_dadda_pg_rca16_u_pg_rca30_fa17_y2;
  assign out[19] = f_u_dadda_pg_rca16_u_pg_rca30_fa18_y2;
  assign out[20] = f_u_dadda_pg_rca16_u_pg_rca30_fa19_y2;
  assign out[21] = f_u_dadda_pg_rca16_u_pg_rca30_fa20_y2;
  assign out[22] = f_u_dadda_pg_rca16_u_pg_rca30_fa21_y2;
  assign out[23] = f_u_dadda_pg_rca16_u_pg_rca30_fa22_y2;
  assign out[24] = f_u_dadda_pg_rca16_u_pg_rca30_fa23_y2;
  assign out[25] = f_u_dadda_pg_rca16_u_pg_rca30_fa24_y2;
  assign out[26] = f_u_dadda_pg_rca16_u_pg_rca30_fa25_y2;
  assign out[27] = f_u_dadda_pg_rca16_u_pg_rca30_fa26_y2;
  assign out[28] = f_u_dadda_pg_rca16_u_pg_rca30_fa27_y2;
  assign out[29] = f_u_dadda_pg_rca16_u_pg_rca30_fa28_y2;
  assign out[30] = f_u_dadda_pg_rca16_u_pg_rca30_fa29_y2;
  assign out[31] = f_u_dadda_pg_rca16_u_pg_rca30_or29_y0;
endmodule