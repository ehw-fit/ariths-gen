module s_cla12(input [11:0] a, input [11:0] b, output [12:0] s_cla12_out);
  wire s_cla12_pg_logic0_or0;
  wire s_cla12_pg_logic0_and0;
  wire s_cla12_pg_logic0_xor0;
  wire s_cla12_pg_logic1_or0;
  wire s_cla12_pg_logic1_and0;
  wire s_cla12_pg_logic1_xor0;
  wire s_cla12_xor1;
  wire s_cla12_and0;
  wire s_cla12_or0;
  wire s_cla12_pg_logic2_or0;
  wire s_cla12_pg_logic2_and0;
  wire s_cla12_pg_logic2_xor0;
  wire s_cla12_xor2;
  wire s_cla12_and1;
  wire s_cla12_and2;
  wire s_cla12_and3;
  wire s_cla12_and4;
  wire s_cla12_or1;
  wire s_cla12_or2;
  wire s_cla12_pg_logic3_or0;
  wire s_cla12_pg_logic3_and0;
  wire s_cla12_pg_logic3_xor0;
  wire s_cla12_xor3;
  wire s_cla12_and5;
  wire s_cla12_and6;
  wire s_cla12_and7;
  wire s_cla12_and8;
  wire s_cla12_and9;
  wire s_cla12_and10;
  wire s_cla12_and11;
  wire s_cla12_or3;
  wire s_cla12_or4;
  wire s_cla12_or5;
  wire s_cla12_pg_logic4_or0;
  wire s_cla12_pg_logic4_and0;
  wire s_cla12_pg_logic4_xor0;
  wire s_cla12_xor4;
  wire s_cla12_and12;
  wire s_cla12_or6;
  wire s_cla12_pg_logic5_or0;
  wire s_cla12_pg_logic5_and0;
  wire s_cla12_pg_logic5_xor0;
  wire s_cla12_xor5;
  wire s_cla12_and13;
  wire s_cla12_and14;
  wire s_cla12_and15;
  wire s_cla12_or7;
  wire s_cla12_or8;
  wire s_cla12_pg_logic6_or0;
  wire s_cla12_pg_logic6_and0;
  wire s_cla12_pg_logic6_xor0;
  wire s_cla12_xor6;
  wire s_cla12_and16;
  wire s_cla12_and17;
  wire s_cla12_and18;
  wire s_cla12_and19;
  wire s_cla12_and20;
  wire s_cla12_and21;
  wire s_cla12_or9;
  wire s_cla12_or10;
  wire s_cla12_or11;
  wire s_cla12_pg_logic7_or0;
  wire s_cla12_pg_logic7_and0;
  wire s_cla12_pg_logic7_xor0;
  wire s_cla12_xor7;
  wire s_cla12_and22;
  wire s_cla12_and23;
  wire s_cla12_and24;
  wire s_cla12_and25;
  wire s_cla12_and26;
  wire s_cla12_and27;
  wire s_cla12_and28;
  wire s_cla12_and29;
  wire s_cla12_and30;
  wire s_cla12_and31;
  wire s_cla12_or12;
  wire s_cla12_or13;
  wire s_cla12_or14;
  wire s_cla12_or15;
  wire s_cla12_pg_logic8_or0;
  wire s_cla12_pg_logic8_and0;
  wire s_cla12_pg_logic8_xor0;
  wire s_cla12_xor8;
  wire s_cla12_and32;
  wire s_cla12_or16;
  wire s_cla12_pg_logic9_or0;
  wire s_cla12_pg_logic9_and0;
  wire s_cla12_pg_logic9_xor0;
  wire s_cla12_xor9;
  wire s_cla12_and33;
  wire s_cla12_and34;
  wire s_cla12_and35;
  wire s_cla12_or17;
  wire s_cla12_or18;
  wire s_cla12_pg_logic10_or0;
  wire s_cla12_pg_logic10_and0;
  wire s_cla12_pg_logic10_xor0;
  wire s_cla12_xor10;
  wire s_cla12_and36;
  wire s_cla12_and37;
  wire s_cla12_and38;
  wire s_cla12_and39;
  wire s_cla12_and40;
  wire s_cla12_and41;
  wire s_cla12_or19;
  wire s_cla12_or20;
  wire s_cla12_or21;
  wire s_cla12_pg_logic11_or0;
  wire s_cla12_pg_logic11_and0;
  wire s_cla12_pg_logic11_xor0;
  wire s_cla12_xor11;
  wire s_cla12_and42;
  wire s_cla12_and43;
  wire s_cla12_and44;
  wire s_cla12_and45;
  wire s_cla12_and46;
  wire s_cla12_and47;
  wire s_cla12_and48;
  wire s_cla12_and49;
  wire s_cla12_and50;
  wire s_cla12_and51;
  wire s_cla12_or22;
  wire s_cla12_or23;
  wire s_cla12_or24;
  wire s_cla12_or25;
  wire s_cla12_xor12;
  wire s_cla12_xor13;

  assign s_cla12_pg_logic0_or0 = a[0] | b[0];
  assign s_cla12_pg_logic0_and0 = a[0] & b[0];
  assign s_cla12_pg_logic0_xor0 = a[0] ^ b[0];
  assign s_cla12_pg_logic1_or0 = a[1] | b[1];
  assign s_cla12_pg_logic1_and0 = a[1] & b[1];
  assign s_cla12_pg_logic1_xor0 = a[1] ^ b[1];
  assign s_cla12_xor1 = s_cla12_pg_logic1_xor0 ^ s_cla12_pg_logic0_and0;
  assign s_cla12_and0 = s_cla12_pg_logic0_and0 & s_cla12_pg_logic1_or0;
  assign s_cla12_or0 = s_cla12_pg_logic1_and0 | s_cla12_and0;
  assign s_cla12_pg_logic2_or0 = a[2] | b[2];
  assign s_cla12_pg_logic2_and0 = a[2] & b[2];
  assign s_cla12_pg_logic2_xor0 = a[2] ^ b[2];
  assign s_cla12_xor2 = s_cla12_pg_logic2_xor0 ^ s_cla12_or0;
  assign s_cla12_and1 = s_cla12_pg_logic2_or0 & s_cla12_pg_logic0_or0;
  assign s_cla12_and2 = s_cla12_pg_logic0_and0 & s_cla12_pg_logic2_or0;
  assign s_cla12_and3 = s_cla12_and2 & s_cla12_pg_logic1_or0;
  assign s_cla12_and4 = s_cla12_pg_logic1_and0 & s_cla12_pg_logic2_or0;
  assign s_cla12_or1 = s_cla12_and3 | s_cla12_and4;
  assign s_cla12_or2 = s_cla12_pg_logic2_and0 | s_cla12_or1;
  assign s_cla12_pg_logic3_or0 = a[3] | b[3];
  assign s_cla12_pg_logic3_and0 = a[3] & b[3];
  assign s_cla12_pg_logic3_xor0 = a[3] ^ b[3];
  assign s_cla12_xor3 = s_cla12_pg_logic3_xor0 ^ s_cla12_or2;
  assign s_cla12_and5 = s_cla12_pg_logic3_or0 & s_cla12_pg_logic1_or0;
  assign s_cla12_and6 = s_cla12_pg_logic0_and0 & s_cla12_pg_logic2_or0;
  assign s_cla12_and7 = s_cla12_pg_logic3_or0 & s_cla12_pg_logic1_or0;
  assign s_cla12_and8 = s_cla12_and6 & s_cla12_and7;
  assign s_cla12_and9 = s_cla12_pg_logic1_and0 & s_cla12_pg_logic3_or0;
  assign s_cla12_and10 = s_cla12_and9 & s_cla12_pg_logic2_or0;
  assign s_cla12_and11 = s_cla12_pg_logic2_and0 & s_cla12_pg_logic3_or0;
  assign s_cla12_or3 = s_cla12_and8 | s_cla12_and11;
  assign s_cla12_or4 = s_cla12_and10 | s_cla12_or3;
  assign s_cla12_or5 = s_cla12_pg_logic3_and0 | s_cla12_or4;
  assign s_cla12_pg_logic4_or0 = a[4] | b[4];
  assign s_cla12_pg_logic4_and0 = a[4] & b[4];
  assign s_cla12_pg_logic4_xor0 = a[4] ^ b[4];
  assign s_cla12_xor4 = s_cla12_pg_logic4_xor0 ^ s_cla12_or5;
  assign s_cla12_and12 = s_cla12_or5 & s_cla12_pg_logic4_or0;
  assign s_cla12_or6 = s_cla12_pg_logic4_and0 | s_cla12_and12;
  assign s_cla12_pg_logic5_or0 = a[5] | b[5];
  assign s_cla12_pg_logic5_and0 = a[5] & b[5];
  assign s_cla12_pg_logic5_xor0 = a[5] ^ b[5];
  assign s_cla12_xor5 = s_cla12_pg_logic5_xor0 ^ s_cla12_or6;
  assign s_cla12_and13 = s_cla12_or5 & s_cla12_pg_logic5_or0;
  assign s_cla12_and14 = s_cla12_and13 & s_cla12_pg_logic4_or0;
  assign s_cla12_and15 = s_cla12_pg_logic4_and0 & s_cla12_pg_logic5_or0;
  assign s_cla12_or7 = s_cla12_and14 | s_cla12_and15;
  assign s_cla12_or8 = s_cla12_pg_logic5_and0 | s_cla12_or7;
  assign s_cla12_pg_logic6_or0 = a[6] | b[6];
  assign s_cla12_pg_logic6_and0 = a[6] & b[6];
  assign s_cla12_pg_logic6_xor0 = a[6] ^ b[6];
  assign s_cla12_xor6 = s_cla12_pg_logic6_xor0 ^ s_cla12_or8;
  assign s_cla12_and16 = s_cla12_or5 & s_cla12_pg_logic5_or0;
  assign s_cla12_and17 = s_cla12_pg_logic6_or0 & s_cla12_pg_logic4_or0;
  assign s_cla12_and18 = s_cla12_and16 & s_cla12_and17;
  assign s_cla12_and19 = s_cla12_pg_logic4_and0 & s_cla12_pg_logic6_or0;
  assign s_cla12_and20 = s_cla12_and19 & s_cla12_pg_logic5_or0;
  assign s_cla12_and21 = s_cla12_pg_logic5_and0 & s_cla12_pg_logic6_or0;
  assign s_cla12_or9 = s_cla12_and18 | s_cla12_and20;
  assign s_cla12_or10 = s_cla12_or9 | s_cla12_and21;
  assign s_cla12_or11 = s_cla12_pg_logic6_and0 | s_cla12_or10;
  assign s_cla12_pg_logic7_or0 = a[7] | b[7];
  assign s_cla12_pg_logic7_and0 = a[7] & b[7];
  assign s_cla12_pg_logic7_xor0 = a[7] ^ b[7];
  assign s_cla12_xor7 = s_cla12_pg_logic7_xor0 ^ s_cla12_or11;
  assign s_cla12_and22 = s_cla12_or5 & s_cla12_pg_logic6_or0;
  assign s_cla12_and23 = s_cla12_pg_logic7_or0 & s_cla12_pg_logic5_or0;
  assign s_cla12_and24 = s_cla12_and22 & s_cla12_and23;
  assign s_cla12_and25 = s_cla12_and24 & s_cla12_pg_logic4_or0;
  assign s_cla12_and26 = s_cla12_pg_logic4_and0 & s_cla12_pg_logic6_or0;
  assign s_cla12_and27 = s_cla12_pg_logic7_or0 & s_cla12_pg_logic5_or0;
  assign s_cla12_and28 = s_cla12_and26 & s_cla12_and27;
  assign s_cla12_and29 = s_cla12_pg_logic5_and0 & s_cla12_pg_logic7_or0;
  assign s_cla12_and30 = s_cla12_and29 & s_cla12_pg_logic6_or0;
  assign s_cla12_and31 = s_cla12_pg_logic6_and0 & s_cla12_pg_logic7_or0;
  assign s_cla12_or12 = s_cla12_and25 | s_cla12_and30;
  assign s_cla12_or13 = s_cla12_and28 | s_cla12_and31;
  assign s_cla12_or14 = s_cla12_or12 | s_cla12_or13;
  assign s_cla12_or15 = s_cla12_pg_logic7_and0 | s_cla12_or14;
  assign s_cla12_pg_logic8_or0 = a[8] | b[8];
  assign s_cla12_pg_logic8_and0 = a[8] & b[8];
  assign s_cla12_pg_logic8_xor0 = a[8] ^ b[8];
  assign s_cla12_xor8 = s_cla12_pg_logic8_xor0 ^ s_cla12_or15;
  assign s_cla12_and32 = s_cla12_or15 & s_cla12_pg_logic8_or0;
  assign s_cla12_or16 = s_cla12_pg_logic8_and0 | s_cla12_and32;
  assign s_cla12_pg_logic9_or0 = a[9] | b[9];
  assign s_cla12_pg_logic9_and0 = a[9] & b[9];
  assign s_cla12_pg_logic9_xor0 = a[9] ^ b[9];
  assign s_cla12_xor9 = s_cla12_pg_logic9_xor0 ^ s_cla12_or16;
  assign s_cla12_and33 = s_cla12_or15 & s_cla12_pg_logic9_or0;
  assign s_cla12_and34 = s_cla12_and33 & s_cla12_pg_logic8_or0;
  assign s_cla12_and35 = s_cla12_pg_logic8_and0 & s_cla12_pg_logic9_or0;
  assign s_cla12_or17 = s_cla12_and34 | s_cla12_and35;
  assign s_cla12_or18 = s_cla12_pg_logic9_and0 | s_cla12_or17;
  assign s_cla12_pg_logic10_or0 = a[10] | b[10];
  assign s_cla12_pg_logic10_and0 = a[10] & b[10];
  assign s_cla12_pg_logic10_xor0 = a[10] ^ b[10];
  assign s_cla12_xor10 = s_cla12_pg_logic10_xor0 ^ s_cla12_or18;
  assign s_cla12_and36 = s_cla12_or15 & s_cla12_pg_logic9_or0;
  assign s_cla12_and37 = s_cla12_pg_logic10_or0 & s_cla12_pg_logic8_or0;
  assign s_cla12_and38 = s_cla12_and36 & s_cla12_and37;
  assign s_cla12_and39 = s_cla12_pg_logic8_and0 & s_cla12_pg_logic10_or0;
  assign s_cla12_and40 = s_cla12_and39 & s_cla12_pg_logic9_or0;
  assign s_cla12_and41 = s_cla12_pg_logic9_and0 & s_cla12_pg_logic10_or0;
  assign s_cla12_or19 = s_cla12_and38 | s_cla12_and40;
  assign s_cla12_or20 = s_cla12_or19 | s_cla12_and41;
  assign s_cla12_or21 = s_cla12_pg_logic10_and0 | s_cla12_or20;
  assign s_cla12_pg_logic11_or0 = a[11] | b[11];
  assign s_cla12_pg_logic11_and0 = a[11] & b[11];
  assign s_cla12_pg_logic11_xor0 = a[11] ^ b[11];
  assign s_cla12_xor11 = s_cla12_pg_logic11_xor0 ^ s_cla12_or21;
  assign s_cla12_and42 = s_cla12_or15 & s_cla12_pg_logic10_or0;
  assign s_cla12_and43 = s_cla12_pg_logic11_or0 & s_cla12_pg_logic9_or0;
  assign s_cla12_and44 = s_cla12_and42 & s_cla12_and43;
  assign s_cla12_and45 = s_cla12_and44 & s_cla12_pg_logic8_or0;
  assign s_cla12_and46 = s_cla12_pg_logic8_and0 & s_cla12_pg_logic10_or0;
  assign s_cla12_and47 = s_cla12_pg_logic11_or0 & s_cla12_pg_logic9_or0;
  assign s_cla12_and48 = s_cla12_and46 & s_cla12_and47;
  assign s_cla12_and49 = s_cla12_pg_logic9_and0 & s_cla12_pg_logic11_or0;
  assign s_cla12_and50 = s_cla12_and49 & s_cla12_pg_logic10_or0;
  assign s_cla12_and51 = s_cla12_pg_logic10_and0 & s_cla12_pg_logic11_or0;
  assign s_cla12_or22 = s_cla12_and45 | s_cla12_and50;
  assign s_cla12_or23 = s_cla12_and48 | s_cla12_and51;
  assign s_cla12_or24 = s_cla12_or22 | s_cla12_or23;
  assign s_cla12_or25 = s_cla12_pg_logic11_and0 | s_cla12_or24;
  assign s_cla12_xor12 = a[11] ^ b[11];
  assign s_cla12_xor13 = s_cla12_xor12 ^ s_cla12_or25;

  assign s_cla12_out[0] = s_cla12_pg_logic0_xor0;
  assign s_cla12_out[1] = s_cla12_xor1;
  assign s_cla12_out[2] = s_cla12_xor2;
  assign s_cla12_out[3] = s_cla12_xor3;
  assign s_cla12_out[4] = s_cla12_xor4;
  assign s_cla12_out[5] = s_cla12_xor5;
  assign s_cla12_out[6] = s_cla12_xor6;
  assign s_cla12_out[7] = s_cla12_xor7;
  assign s_cla12_out[8] = s_cla12_xor8;
  assign s_cla12_out[9] = s_cla12_xor9;
  assign s_cla12_out[10] = s_cla12_xor10;
  assign s_cla12_out[11] = s_cla12_xor11;
  assign s_cla12_out[12] = s_cla12_xor13;
endmodule