module s_arrmul12(input [11:0] a, input [11:0] b, output [23:0] s_arrmul12_out);
  wire s_arrmul12_and0_0;
  wire s_arrmul12_and1_0;
  wire s_arrmul12_and2_0;
  wire s_arrmul12_and3_0;
  wire s_arrmul12_and4_0;
  wire s_arrmul12_and5_0;
  wire s_arrmul12_and6_0;
  wire s_arrmul12_and7_0;
  wire s_arrmul12_and8_0;
  wire s_arrmul12_and9_0;
  wire s_arrmul12_and10_0;
  wire s_arrmul12_nand11_0;
  wire s_arrmul12_and0_1;
  wire s_arrmul12_ha0_1_xor0;
  wire s_arrmul12_ha0_1_and0;
  wire s_arrmul12_and1_1;
  wire s_arrmul12_fa1_1_xor0;
  wire s_arrmul12_fa1_1_and0;
  wire s_arrmul12_fa1_1_xor1;
  wire s_arrmul12_fa1_1_and1;
  wire s_arrmul12_fa1_1_or0;
  wire s_arrmul12_and2_1;
  wire s_arrmul12_fa2_1_xor0;
  wire s_arrmul12_fa2_1_and0;
  wire s_arrmul12_fa2_1_xor1;
  wire s_arrmul12_fa2_1_and1;
  wire s_arrmul12_fa2_1_or0;
  wire s_arrmul12_and3_1;
  wire s_arrmul12_fa3_1_xor0;
  wire s_arrmul12_fa3_1_and0;
  wire s_arrmul12_fa3_1_xor1;
  wire s_arrmul12_fa3_1_and1;
  wire s_arrmul12_fa3_1_or0;
  wire s_arrmul12_and4_1;
  wire s_arrmul12_fa4_1_xor0;
  wire s_arrmul12_fa4_1_and0;
  wire s_arrmul12_fa4_1_xor1;
  wire s_arrmul12_fa4_1_and1;
  wire s_arrmul12_fa4_1_or0;
  wire s_arrmul12_and5_1;
  wire s_arrmul12_fa5_1_xor0;
  wire s_arrmul12_fa5_1_and0;
  wire s_arrmul12_fa5_1_xor1;
  wire s_arrmul12_fa5_1_and1;
  wire s_arrmul12_fa5_1_or0;
  wire s_arrmul12_and6_1;
  wire s_arrmul12_fa6_1_xor0;
  wire s_arrmul12_fa6_1_and0;
  wire s_arrmul12_fa6_1_xor1;
  wire s_arrmul12_fa6_1_and1;
  wire s_arrmul12_fa6_1_or0;
  wire s_arrmul12_and7_1;
  wire s_arrmul12_fa7_1_xor0;
  wire s_arrmul12_fa7_1_and0;
  wire s_arrmul12_fa7_1_xor1;
  wire s_arrmul12_fa7_1_and1;
  wire s_arrmul12_fa7_1_or0;
  wire s_arrmul12_and8_1;
  wire s_arrmul12_fa8_1_xor0;
  wire s_arrmul12_fa8_1_and0;
  wire s_arrmul12_fa8_1_xor1;
  wire s_arrmul12_fa8_1_and1;
  wire s_arrmul12_fa8_1_or0;
  wire s_arrmul12_and9_1;
  wire s_arrmul12_fa9_1_xor0;
  wire s_arrmul12_fa9_1_and0;
  wire s_arrmul12_fa9_1_xor1;
  wire s_arrmul12_fa9_1_and1;
  wire s_arrmul12_fa9_1_or0;
  wire s_arrmul12_and10_1;
  wire s_arrmul12_fa10_1_xor0;
  wire s_arrmul12_fa10_1_and0;
  wire s_arrmul12_fa10_1_xor1;
  wire s_arrmul12_fa10_1_and1;
  wire s_arrmul12_fa10_1_or0;
  wire s_arrmul12_nand11_1;
  wire s_arrmul12_fa11_1_xor0;
  wire s_arrmul12_fa11_1_xor1;
  wire s_arrmul12_fa11_1_and1;
  wire s_arrmul12_fa11_1_or0;
  wire s_arrmul12_and0_2;
  wire s_arrmul12_ha0_2_xor0;
  wire s_arrmul12_ha0_2_and0;
  wire s_arrmul12_and1_2;
  wire s_arrmul12_fa1_2_xor0;
  wire s_arrmul12_fa1_2_and0;
  wire s_arrmul12_fa1_2_xor1;
  wire s_arrmul12_fa1_2_and1;
  wire s_arrmul12_fa1_2_or0;
  wire s_arrmul12_and2_2;
  wire s_arrmul12_fa2_2_xor0;
  wire s_arrmul12_fa2_2_and0;
  wire s_arrmul12_fa2_2_xor1;
  wire s_arrmul12_fa2_2_and1;
  wire s_arrmul12_fa2_2_or0;
  wire s_arrmul12_and3_2;
  wire s_arrmul12_fa3_2_xor0;
  wire s_arrmul12_fa3_2_and0;
  wire s_arrmul12_fa3_2_xor1;
  wire s_arrmul12_fa3_2_and1;
  wire s_arrmul12_fa3_2_or0;
  wire s_arrmul12_and4_2;
  wire s_arrmul12_fa4_2_xor0;
  wire s_arrmul12_fa4_2_and0;
  wire s_arrmul12_fa4_2_xor1;
  wire s_arrmul12_fa4_2_and1;
  wire s_arrmul12_fa4_2_or0;
  wire s_arrmul12_and5_2;
  wire s_arrmul12_fa5_2_xor0;
  wire s_arrmul12_fa5_2_and0;
  wire s_arrmul12_fa5_2_xor1;
  wire s_arrmul12_fa5_2_and1;
  wire s_arrmul12_fa5_2_or0;
  wire s_arrmul12_and6_2;
  wire s_arrmul12_fa6_2_xor0;
  wire s_arrmul12_fa6_2_and0;
  wire s_arrmul12_fa6_2_xor1;
  wire s_arrmul12_fa6_2_and1;
  wire s_arrmul12_fa6_2_or0;
  wire s_arrmul12_and7_2;
  wire s_arrmul12_fa7_2_xor0;
  wire s_arrmul12_fa7_2_and0;
  wire s_arrmul12_fa7_2_xor1;
  wire s_arrmul12_fa7_2_and1;
  wire s_arrmul12_fa7_2_or0;
  wire s_arrmul12_and8_2;
  wire s_arrmul12_fa8_2_xor0;
  wire s_arrmul12_fa8_2_and0;
  wire s_arrmul12_fa8_2_xor1;
  wire s_arrmul12_fa8_2_and1;
  wire s_arrmul12_fa8_2_or0;
  wire s_arrmul12_and9_2;
  wire s_arrmul12_fa9_2_xor0;
  wire s_arrmul12_fa9_2_and0;
  wire s_arrmul12_fa9_2_xor1;
  wire s_arrmul12_fa9_2_and1;
  wire s_arrmul12_fa9_2_or0;
  wire s_arrmul12_and10_2;
  wire s_arrmul12_fa10_2_xor0;
  wire s_arrmul12_fa10_2_and0;
  wire s_arrmul12_fa10_2_xor1;
  wire s_arrmul12_fa10_2_and1;
  wire s_arrmul12_fa10_2_or0;
  wire s_arrmul12_nand11_2;
  wire s_arrmul12_fa11_2_xor0;
  wire s_arrmul12_fa11_2_and0;
  wire s_arrmul12_fa11_2_xor1;
  wire s_arrmul12_fa11_2_and1;
  wire s_arrmul12_fa11_2_or0;
  wire s_arrmul12_and0_3;
  wire s_arrmul12_ha0_3_xor0;
  wire s_arrmul12_ha0_3_and0;
  wire s_arrmul12_and1_3;
  wire s_arrmul12_fa1_3_xor0;
  wire s_arrmul12_fa1_3_and0;
  wire s_arrmul12_fa1_3_xor1;
  wire s_arrmul12_fa1_3_and1;
  wire s_arrmul12_fa1_3_or0;
  wire s_arrmul12_and2_3;
  wire s_arrmul12_fa2_3_xor0;
  wire s_arrmul12_fa2_3_and0;
  wire s_arrmul12_fa2_3_xor1;
  wire s_arrmul12_fa2_3_and1;
  wire s_arrmul12_fa2_3_or0;
  wire s_arrmul12_and3_3;
  wire s_arrmul12_fa3_3_xor0;
  wire s_arrmul12_fa3_3_and0;
  wire s_arrmul12_fa3_3_xor1;
  wire s_arrmul12_fa3_3_and1;
  wire s_arrmul12_fa3_3_or0;
  wire s_arrmul12_and4_3;
  wire s_arrmul12_fa4_3_xor0;
  wire s_arrmul12_fa4_3_and0;
  wire s_arrmul12_fa4_3_xor1;
  wire s_arrmul12_fa4_3_and1;
  wire s_arrmul12_fa4_3_or0;
  wire s_arrmul12_and5_3;
  wire s_arrmul12_fa5_3_xor0;
  wire s_arrmul12_fa5_3_and0;
  wire s_arrmul12_fa5_3_xor1;
  wire s_arrmul12_fa5_3_and1;
  wire s_arrmul12_fa5_3_or0;
  wire s_arrmul12_and6_3;
  wire s_arrmul12_fa6_3_xor0;
  wire s_arrmul12_fa6_3_and0;
  wire s_arrmul12_fa6_3_xor1;
  wire s_arrmul12_fa6_3_and1;
  wire s_arrmul12_fa6_3_or0;
  wire s_arrmul12_and7_3;
  wire s_arrmul12_fa7_3_xor0;
  wire s_arrmul12_fa7_3_and0;
  wire s_arrmul12_fa7_3_xor1;
  wire s_arrmul12_fa7_3_and1;
  wire s_arrmul12_fa7_3_or0;
  wire s_arrmul12_and8_3;
  wire s_arrmul12_fa8_3_xor0;
  wire s_arrmul12_fa8_3_and0;
  wire s_arrmul12_fa8_3_xor1;
  wire s_arrmul12_fa8_3_and1;
  wire s_arrmul12_fa8_3_or0;
  wire s_arrmul12_and9_3;
  wire s_arrmul12_fa9_3_xor0;
  wire s_arrmul12_fa9_3_and0;
  wire s_arrmul12_fa9_3_xor1;
  wire s_arrmul12_fa9_3_and1;
  wire s_arrmul12_fa9_3_or0;
  wire s_arrmul12_and10_3;
  wire s_arrmul12_fa10_3_xor0;
  wire s_arrmul12_fa10_3_and0;
  wire s_arrmul12_fa10_3_xor1;
  wire s_arrmul12_fa10_3_and1;
  wire s_arrmul12_fa10_3_or0;
  wire s_arrmul12_nand11_3;
  wire s_arrmul12_fa11_3_xor0;
  wire s_arrmul12_fa11_3_and0;
  wire s_arrmul12_fa11_3_xor1;
  wire s_arrmul12_fa11_3_and1;
  wire s_arrmul12_fa11_3_or0;
  wire s_arrmul12_and0_4;
  wire s_arrmul12_ha0_4_xor0;
  wire s_arrmul12_ha0_4_and0;
  wire s_arrmul12_and1_4;
  wire s_arrmul12_fa1_4_xor0;
  wire s_arrmul12_fa1_4_and0;
  wire s_arrmul12_fa1_4_xor1;
  wire s_arrmul12_fa1_4_and1;
  wire s_arrmul12_fa1_4_or0;
  wire s_arrmul12_and2_4;
  wire s_arrmul12_fa2_4_xor0;
  wire s_arrmul12_fa2_4_and0;
  wire s_arrmul12_fa2_4_xor1;
  wire s_arrmul12_fa2_4_and1;
  wire s_arrmul12_fa2_4_or0;
  wire s_arrmul12_and3_4;
  wire s_arrmul12_fa3_4_xor0;
  wire s_arrmul12_fa3_4_and0;
  wire s_arrmul12_fa3_4_xor1;
  wire s_arrmul12_fa3_4_and1;
  wire s_arrmul12_fa3_4_or0;
  wire s_arrmul12_and4_4;
  wire s_arrmul12_fa4_4_xor0;
  wire s_arrmul12_fa4_4_and0;
  wire s_arrmul12_fa4_4_xor1;
  wire s_arrmul12_fa4_4_and1;
  wire s_arrmul12_fa4_4_or0;
  wire s_arrmul12_and5_4;
  wire s_arrmul12_fa5_4_xor0;
  wire s_arrmul12_fa5_4_and0;
  wire s_arrmul12_fa5_4_xor1;
  wire s_arrmul12_fa5_4_and1;
  wire s_arrmul12_fa5_4_or0;
  wire s_arrmul12_and6_4;
  wire s_arrmul12_fa6_4_xor0;
  wire s_arrmul12_fa6_4_and0;
  wire s_arrmul12_fa6_4_xor1;
  wire s_arrmul12_fa6_4_and1;
  wire s_arrmul12_fa6_4_or0;
  wire s_arrmul12_and7_4;
  wire s_arrmul12_fa7_4_xor0;
  wire s_arrmul12_fa7_4_and0;
  wire s_arrmul12_fa7_4_xor1;
  wire s_arrmul12_fa7_4_and1;
  wire s_arrmul12_fa7_4_or0;
  wire s_arrmul12_and8_4;
  wire s_arrmul12_fa8_4_xor0;
  wire s_arrmul12_fa8_4_and0;
  wire s_arrmul12_fa8_4_xor1;
  wire s_arrmul12_fa8_4_and1;
  wire s_arrmul12_fa8_4_or0;
  wire s_arrmul12_and9_4;
  wire s_arrmul12_fa9_4_xor0;
  wire s_arrmul12_fa9_4_and0;
  wire s_arrmul12_fa9_4_xor1;
  wire s_arrmul12_fa9_4_and1;
  wire s_arrmul12_fa9_4_or0;
  wire s_arrmul12_and10_4;
  wire s_arrmul12_fa10_4_xor0;
  wire s_arrmul12_fa10_4_and0;
  wire s_arrmul12_fa10_4_xor1;
  wire s_arrmul12_fa10_4_and1;
  wire s_arrmul12_fa10_4_or0;
  wire s_arrmul12_nand11_4;
  wire s_arrmul12_fa11_4_xor0;
  wire s_arrmul12_fa11_4_and0;
  wire s_arrmul12_fa11_4_xor1;
  wire s_arrmul12_fa11_4_and1;
  wire s_arrmul12_fa11_4_or0;
  wire s_arrmul12_and0_5;
  wire s_arrmul12_ha0_5_xor0;
  wire s_arrmul12_ha0_5_and0;
  wire s_arrmul12_and1_5;
  wire s_arrmul12_fa1_5_xor0;
  wire s_arrmul12_fa1_5_and0;
  wire s_arrmul12_fa1_5_xor1;
  wire s_arrmul12_fa1_5_and1;
  wire s_arrmul12_fa1_5_or0;
  wire s_arrmul12_and2_5;
  wire s_arrmul12_fa2_5_xor0;
  wire s_arrmul12_fa2_5_and0;
  wire s_arrmul12_fa2_5_xor1;
  wire s_arrmul12_fa2_5_and1;
  wire s_arrmul12_fa2_5_or0;
  wire s_arrmul12_and3_5;
  wire s_arrmul12_fa3_5_xor0;
  wire s_arrmul12_fa3_5_and0;
  wire s_arrmul12_fa3_5_xor1;
  wire s_arrmul12_fa3_5_and1;
  wire s_arrmul12_fa3_5_or0;
  wire s_arrmul12_and4_5;
  wire s_arrmul12_fa4_5_xor0;
  wire s_arrmul12_fa4_5_and0;
  wire s_arrmul12_fa4_5_xor1;
  wire s_arrmul12_fa4_5_and1;
  wire s_arrmul12_fa4_5_or0;
  wire s_arrmul12_and5_5;
  wire s_arrmul12_fa5_5_xor0;
  wire s_arrmul12_fa5_5_and0;
  wire s_arrmul12_fa5_5_xor1;
  wire s_arrmul12_fa5_5_and1;
  wire s_arrmul12_fa5_5_or0;
  wire s_arrmul12_and6_5;
  wire s_arrmul12_fa6_5_xor0;
  wire s_arrmul12_fa6_5_and0;
  wire s_arrmul12_fa6_5_xor1;
  wire s_arrmul12_fa6_5_and1;
  wire s_arrmul12_fa6_5_or0;
  wire s_arrmul12_and7_5;
  wire s_arrmul12_fa7_5_xor0;
  wire s_arrmul12_fa7_5_and0;
  wire s_arrmul12_fa7_5_xor1;
  wire s_arrmul12_fa7_5_and1;
  wire s_arrmul12_fa7_5_or0;
  wire s_arrmul12_and8_5;
  wire s_arrmul12_fa8_5_xor0;
  wire s_arrmul12_fa8_5_and0;
  wire s_arrmul12_fa8_5_xor1;
  wire s_arrmul12_fa8_5_and1;
  wire s_arrmul12_fa8_5_or0;
  wire s_arrmul12_and9_5;
  wire s_arrmul12_fa9_5_xor0;
  wire s_arrmul12_fa9_5_and0;
  wire s_arrmul12_fa9_5_xor1;
  wire s_arrmul12_fa9_5_and1;
  wire s_arrmul12_fa9_5_or0;
  wire s_arrmul12_and10_5;
  wire s_arrmul12_fa10_5_xor0;
  wire s_arrmul12_fa10_5_and0;
  wire s_arrmul12_fa10_5_xor1;
  wire s_arrmul12_fa10_5_and1;
  wire s_arrmul12_fa10_5_or0;
  wire s_arrmul12_nand11_5;
  wire s_arrmul12_fa11_5_xor0;
  wire s_arrmul12_fa11_5_and0;
  wire s_arrmul12_fa11_5_xor1;
  wire s_arrmul12_fa11_5_and1;
  wire s_arrmul12_fa11_5_or0;
  wire s_arrmul12_and0_6;
  wire s_arrmul12_ha0_6_xor0;
  wire s_arrmul12_ha0_6_and0;
  wire s_arrmul12_and1_6;
  wire s_arrmul12_fa1_6_xor0;
  wire s_arrmul12_fa1_6_and0;
  wire s_arrmul12_fa1_6_xor1;
  wire s_arrmul12_fa1_6_and1;
  wire s_arrmul12_fa1_6_or0;
  wire s_arrmul12_and2_6;
  wire s_arrmul12_fa2_6_xor0;
  wire s_arrmul12_fa2_6_and0;
  wire s_arrmul12_fa2_6_xor1;
  wire s_arrmul12_fa2_6_and1;
  wire s_arrmul12_fa2_6_or0;
  wire s_arrmul12_and3_6;
  wire s_arrmul12_fa3_6_xor0;
  wire s_arrmul12_fa3_6_and0;
  wire s_arrmul12_fa3_6_xor1;
  wire s_arrmul12_fa3_6_and1;
  wire s_arrmul12_fa3_6_or0;
  wire s_arrmul12_and4_6;
  wire s_arrmul12_fa4_6_xor0;
  wire s_arrmul12_fa4_6_and0;
  wire s_arrmul12_fa4_6_xor1;
  wire s_arrmul12_fa4_6_and1;
  wire s_arrmul12_fa4_6_or0;
  wire s_arrmul12_and5_6;
  wire s_arrmul12_fa5_6_xor0;
  wire s_arrmul12_fa5_6_and0;
  wire s_arrmul12_fa5_6_xor1;
  wire s_arrmul12_fa5_6_and1;
  wire s_arrmul12_fa5_6_or0;
  wire s_arrmul12_and6_6;
  wire s_arrmul12_fa6_6_xor0;
  wire s_arrmul12_fa6_6_and0;
  wire s_arrmul12_fa6_6_xor1;
  wire s_arrmul12_fa6_6_and1;
  wire s_arrmul12_fa6_6_or0;
  wire s_arrmul12_and7_6;
  wire s_arrmul12_fa7_6_xor0;
  wire s_arrmul12_fa7_6_and0;
  wire s_arrmul12_fa7_6_xor1;
  wire s_arrmul12_fa7_6_and1;
  wire s_arrmul12_fa7_6_or0;
  wire s_arrmul12_and8_6;
  wire s_arrmul12_fa8_6_xor0;
  wire s_arrmul12_fa8_6_and0;
  wire s_arrmul12_fa8_6_xor1;
  wire s_arrmul12_fa8_6_and1;
  wire s_arrmul12_fa8_6_or0;
  wire s_arrmul12_and9_6;
  wire s_arrmul12_fa9_6_xor0;
  wire s_arrmul12_fa9_6_and0;
  wire s_arrmul12_fa9_6_xor1;
  wire s_arrmul12_fa9_6_and1;
  wire s_arrmul12_fa9_6_or0;
  wire s_arrmul12_and10_6;
  wire s_arrmul12_fa10_6_xor0;
  wire s_arrmul12_fa10_6_and0;
  wire s_arrmul12_fa10_6_xor1;
  wire s_arrmul12_fa10_6_and1;
  wire s_arrmul12_fa10_6_or0;
  wire s_arrmul12_nand11_6;
  wire s_arrmul12_fa11_6_xor0;
  wire s_arrmul12_fa11_6_and0;
  wire s_arrmul12_fa11_6_xor1;
  wire s_arrmul12_fa11_6_and1;
  wire s_arrmul12_fa11_6_or0;
  wire s_arrmul12_and0_7;
  wire s_arrmul12_ha0_7_xor0;
  wire s_arrmul12_ha0_7_and0;
  wire s_arrmul12_and1_7;
  wire s_arrmul12_fa1_7_xor0;
  wire s_arrmul12_fa1_7_and0;
  wire s_arrmul12_fa1_7_xor1;
  wire s_arrmul12_fa1_7_and1;
  wire s_arrmul12_fa1_7_or0;
  wire s_arrmul12_and2_7;
  wire s_arrmul12_fa2_7_xor0;
  wire s_arrmul12_fa2_7_and0;
  wire s_arrmul12_fa2_7_xor1;
  wire s_arrmul12_fa2_7_and1;
  wire s_arrmul12_fa2_7_or0;
  wire s_arrmul12_and3_7;
  wire s_arrmul12_fa3_7_xor0;
  wire s_arrmul12_fa3_7_and0;
  wire s_arrmul12_fa3_7_xor1;
  wire s_arrmul12_fa3_7_and1;
  wire s_arrmul12_fa3_7_or0;
  wire s_arrmul12_and4_7;
  wire s_arrmul12_fa4_7_xor0;
  wire s_arrmul12_fa4_7_and0;
  wire s_arrmul12_fa4_7_xor1;
  wire s_arrmul12_fa4_7_and1;
  wire s_arrmul12_fa4_7_or0;
  wire s_arrmul12_and5_7;
  wire s_arrmul12_fa5_7_xor0;
  wire s_arrmul12_fa5_7_and0;
  wire s_arrmul12_fa5_7_xor1;
  wire s_arrmul12_fa5_7_and1;
  wire s_arrmul12_fa5_7_or0;
  wire s_arrmul12_and6_7;
  wire s_arrmul12_fa6_7_xor0;
  wire s_arrmul12_fa6_7_and0;
  wire s_arrmul12_fa6_7_xor1;
  wire s_arrmul12_fa6_7_and1;
  wire s_arrmul12_fa6_7_or0;
  wire s_arrmul12_and7_7;
  wire s_arrmul12_fa7_7_xor0;
  wire s_arrmul12_fa7_7_and0;
  wire s_arrmul12_fa7_7_xor1;
  wire s_arrmul12_fa7_7_and1;
  wire s_arrmul12_fa7_7_or0;
  wire s_arrmul12_and8_7;
  wire s_arrmul12_fa8_7_xor0;
  wire s_arrmul12_fa8_7_and0;
  wire s_arrmul12_fa8_7_xor1;
  wire s_arrmul12_fa8_7_and1;
  wire s_arrmul12_fa8_7_or0;
  wire s_arrmul12_and9_7;
  wire s_arrmul12_fa9_7_xor0;
  wire s_arrmul12_fa9_7_and0;
  wire s_arrmul12_fa9_7_xor1;
  wire s_arrmul12_fa9_7_and1;
  wire s_arrmul12_fa9_7_or0;
  wire s_arrmul12_and10_7;
  wire s_arrmul12_fa10_7_xor0;
  wire s_arrmul12_fa10_7_and0;
  wire s_arrmul12_fa10_7_xor1;
  wire s_arrmul12_fa10_7_and1;
  wire s_arrmul12_fa10_7_or0;
  wire s_arrmul12_nand11_7;
  wire s_arrmul12_fa11_7_xor0;
  wire s_arrmul12_fa11_7_and0;
  wire s_arrmul12_fa11_7_xor1;
  wire s_arrmul12_fa11_7_and1;
  wire s_arrmul12_fa11_7_or0;
  wire s_arrmul12_and0_8;
  wire s_arrmul12_ha0_8_xor0;
  wire s_arrmul12_ha0_8_and0;
  wire s_arrmul12_and1_8;
  wire s_arrmul12_fa1_8_xor0;
  wire s_arrmul12_fa1_8_and0;
  wire s_arrmul12_fa1_8_xor1;
  wire s_arrmul12_fa1_8_and1;
  wire s_arrmul12_fa1_8_or0;
  wire s_arrmul12_and2_8;
  wire s_arrmul12_fa2_8_xor0;
  wire s_arrmul12_fa2_8_and0;
  wire s_arrmul12_fa2_8_xor1;
  wire s_arrmul12_fa2_8_and1;
  wire s_arrmul12_fa2_8_or0;
  wire s_arrmul12_and3_8;
  wire s_arrmul12_fa3_8_xor0;
  wire s_arrmul12_fa3_8_and0;
  wire s_arrmul12_fa3_8_xor1;
  wire s_arrmul12_fa3_8_and1;
  wire s_arrmul12_fa3_8_or0;
  wire s_arrmul12_and4_8;
  wire s_arrmul12_fa4_8_xor0;
  wire s_arrmul12_fa4_8_and0;
  wire s_arrmul12_fa4_8_xor1;
  wire s_arrmul12_fa4_8_and1;
  wire s_arrmul12_fa4_8_or0;
  wire s_arrmul12_and5_8;
  wire s_arrmul12_fa5_8_xor0;
  wire s_arrmul12_fa5_8_and0;
  wire s_arrmul12_fa5_8_xor1;
  wire s_arrmul12_fa5_8_and1;
  wire s_arrmul12_fa5_8_or0;
  wire s_arrmul12_and6_8;
  wire s_arrmul12_fa6_8_xor0;
  wire s_arrmul12_fa6_8_and0;
  wire s_arrmul12_fa6_8_xor1;
  wire s_arrmul12_fa6_8_and1;
  wire s_arrmul12_fa6_8_or0;
  wire s_arrmul12_and7_8;
  wire s_arrmul12_fa7_8_xor0;
  wire s_arrmul12_fa7_8_and0;
  wire s_arrmul12_fa7_8_xor1;
  wire s_arrmul12_fa7_8_and1;
  wire s_arrmul12_fa7_8_or0;
  wire s_arrmul12_and8_8;
  wire s_arrmul12_fa8_8_xor0;
  wire s_arrmul12_fa8_8_and0;
  wire s_arrmul12_fa8_8_xor1;
  wire s_arrmul12_fa8_8_and1;
  wire s_arrmul12_fa8_8_or0;
  wire s_arrmul12_and9_8;
  wire s_arrmul12_fa9_8_xor0;
  wire s_arrmul12_fa9_8_and0;
  wire s_arrmul12_fa9_8_xor1;
  wire s_arrmul12_fa9_8_and1;
  wire s_arrmul12_fa9_8_or0;
  wire s_arrmul12_and10_8;
  wire s_arrmul12_fa10_8_xor0;
  wire s_arrmul12_fa10_8_and0;
  wire s_arrmul12_fa10_8_xor1;
  wire s_arrmul12_fa10_8_and1;
  wire s_arrmul12_fa10_8_or0;
  wire s_arrmul12_nand11_8;
  wire s_arrmul12_fa11_8_xor0;
  wire s_arrmul12_fa11_8_and0;
  wire s_arrmul12_fa11_8_xor1;
  wire s_arrmul12_fa11_8_and1;
  wire s_arrmul12_fa11_8_or0;
  wire s_arrmul12_and0_9;
  wire s_arrmul12_ha0_9_xor0;
  wire s_arrmul12_ha0_9_and0;
  wire s_arrmul12_and1_9;
  wire s_arrmul12_fa1_9_xor0;
  wire s_arrmul12_fa1_9_and0;
  wire s_arrmul12_fa1_9_xor1;
  wire s_arrmul12_fa1_9_and1;
  wire s_arrmul12_fa1_9_or0;
  wire s_arrmul12_and2_9;
  wire s_arrmul12_fa2_9_xor0;
  wire s_arrmul12_fa2_9_and0;
  wire s_arrmul12_fa2_9_xor1;
  wire s_arrmul12_fa2_9_and1;
  wire s_arrmul12_fa2_9_or0;
  wire s_arrmul12_and3_9;
  wire s_arrmul12_fa3_9_xor0;
  wire s_arrmul12_fa3_9_and0;
  wire s_arrmul12_fa3_9_xor1;
  wire s_arrmul12_fa3_9_and1;
  wire s_arrmul12_fa3_9_or0;
  wire s_arrmul12_and4_9;
  wire s_arrmul12_fa4_9_xor0;
  wire s_arrmul12_fa4_9_and0;
  wire s_arrmul12_fa4_9_xor1;
  wire s_arrmul12_fa4_9_and1;
  wire s_arrmul12_fa4_9_or0;
  wire s_arrmul12_and5_9;
  wire s_arrmul12_fa5_9_xor0;
  wire s_arrmul12_fa5_9_and0;
  wire s_arrmul12_fa5_9_xor1;
  wire s_arrmul12_fa5_9_and1;
  wire s_arrmul12_fa5_9_or0;
  wire s_arrmul12_and6_9;
  wire s_arrmul12_fa6_9_xor0;
  wire s_arrmul12_fa6_9_and0;
  wire s_arrmul12_fa6_9_xor1;
  wire s_arrmul12_fa6_9_and1;
  wire s_arrmul12_fa6_9_or0;
  wire s_arrmul12_and7_9;
  wire s_arrmul12_fa7_9_xor0;
  wire s_arrmul12_fa7_9_and0;
  wire s_arrmul12_fa7_9_xor1;
  wire s_arrmul12_fa7_9_and1;
  wire s_arrmul12_fa7_9_or0;
  wire s_arrmul12_and8_9;
  wire s_arrmul12_fa8_9_xor0;
  wire s_arrmul12_fa8_9_and0;
  wire s_arrmul12_fa8_9_xor1;
  wire s_arrmul12_fa8_9_and1;
  wire s_arrmul12_fa8_9_or0;
  wire s_arrmul12_and9_9;
  wire s_arrmul12_fa9_9_xor0;
  wire s_arrmul12_fa9_9_and0;
  wire s_arrmul12_fa9_9_xor1;
  wire s_arrmul12_fa9_9_and1;
  wire s_arrmul12_fa9_9_or0;
  wire s_arrmul12_and10_9;
  wire s_arrmul12_fa10_9_xor0;
  wire s_arrmul12_fa10_9_and0;
  wire s_arrmul12_fa10_9_xor1;
  wire s_arrmul12_fa10_9_and1;
  wire s_arrmul12_fa10_9_or0;
  wire s_arrmul12_nand11_9;
  wire s_arrmul12_fa11_9_xor0;
  wire s_arrmul12_fa11_9_and0;
  wire s_arrmul12_fa11_9_xor1;
  wire s_arrmul12_fa11_9_and1;
  wire s_arrmul12_fa11_9_or0;
  wire s_arrmul12_and0_10;
  wire s_arrmul12_ha0_10_xor0;
  wire s_arrmul12_ha0_10_and0;
  wire s_arrmul12_and1_10;
  wire s_arrmul12_fa1_10_xor0;
  wire s_arrmul12_fa1_10_and0;
  wire s_arrmul12_fa1_10_xor1;
  wire s_arrmul12_fa1_10_and1;
  wire s_arrmul12_fa1_10_or0;
  wire s_arrmul12_and2_10;
  wire s_arrmul12_fa2_10_xor0;
  wire s_arrmul12_fa2_10_and0;
  wire s_arrmul12_fa2_10_xor1;
  wire s_arrmul12_fa2_10_and1;
  wire s_arrmul12_fa2_10_or0;
  wire s_arrmul12_and3_10;
  wire s_arrmul12_fa3_10_xor0;
  wire s_arrmul12_fa3_10_and0;
  wire s_arrmul12_fa3_10_xor1;
  wire s_arrmul12_fa3_10_and1;
  wire s_arrmul12_fa3_10_or0;
  wire s_arrmul12_and4_10;
  wire s_arrmul12_fa4_10_xor0;
  wire s_arrmul12_fa4_10_and0;
  wire s_arrmul12_fa4_10_xor1;
  wire s_arrmul12_fa4_10_and1;
  wire s_arrmul12_fa4_10_or0;
  wire s_arrmul12_and5_10;
  wire s_arrmul12_fa5_10_xor0;
  wire s_arrmul12_fa5_10_and0;
  wire s_arrmul12_fa5_10_xor1;
  wire s_arrmul12_fa5_10_and1;
  wire s_arrmul12_fa5_10_or0;
  wire s_arrmul12_and6_10;
  wire s_arrmul12_fa6_10_xor0;
  wire s_arrmul12_fa6_10_and0;
  wire s_arrmul12_fa6_10_xor1;
  wire s_arrmul12_fa6_10_and1;
  wire s_arrmul12_fa6_10_or0;
  wire s_arrmul12_and7_10;
  wire s_arrmul12_fa7_10_xor0;
  wire s_arrmul12_fa7_10_and0;
  wire s_arrmul12_fa7_10_xor1;
  wire s_arrmul12_fa7_10_and1;
  wire s_arrmul12_fa7_10_or0;
  wire s_arrmul12_and8_10;
  wire s_arrmul12_fa8_10_xor0;
  wire s_arrmul12_fa8_10_and0;
  wire s_arrmul12_fa8_10_xor1;
  wire s_arrmul12_fa8_10_and1;
  wire s_arrmul12_fa8_10_or0;
  wire s_arrmul12_and9_10;
  wire s_arrmul12_fa9_10_xor0;
  wire s_arrmul12_fa9_10_and0;
  wire s_arrmul12_fa9_10_xor1;
  wire s_arrmul12_fa9_10_and1;
  wire s_arrmul12_fa9_10_or0;
  wire s_arrmul12_and10_10;
  wire s_arrmul12_fa10_10_xor0;
  wire s_arrmul12_fa10_10_and0;
  wire s_arrmul12_fa10_10_xor1;
  wire s_arrmul12_fa10_10_and1;
  wire s_arrmul12_fa10_10_or0;
  wire s_arrmul12_nand11_10;
  wire s_arrmul12_fa11_10_xor0;
  wire s_arrmul12_fa11_10_and0;
  wire s_arrmul12_fa11_10_xor1;
  wire s_arrmul12_fa11_10_and1;
  wire s_arrmul12_fa11_10_or0;
  wire s_arrmul12_nand0_11;
  wire s_arrmul12_ha0_11_xor0;
  wire s_arrmul12_ha0_11_and0;
  wire s_arrmul12_nand1_11;
  wire s_arrmul12_fa1_11_xor0;
  wire s_arrmul12_fa1_11_and0;
  wire s_arrmul12_fa1_11_xor1;
  wire s_arrmul12_fa1_11_and1;
  wire s_arrmul12_fa1_11_or0;
  wire s_arrmul12_nand2_11;
  wire s_arrmul12_fa2_11_xor0;
  wire s_arrmul12_fa2_11_and0;
  wire s_arrmul12_fa2_11_xor1;
  wire s_arrmul12_fa2_11_and1;
  wire s_arrmul12_fa2_11_or0;
  wire s_arrmul12_nand3_11;
  wire s_arrmul12_fa3_11_xor0;
  wire s_arrmul12_fa3_11_and0;
  wire s_arrmul12_fa3_11_xor1;
  wire s_arrmul12_fa3_11_and1;
  wire s_arrmul12_fa3_11_or0;
  wire s_arrmul12_nand4_11;
  wire s_arrmul12_fa4_11_xor0;
  wire s_arrmul12_fa4_11_and0;
  wire s_arrmul12_fa4_11_xor1;
  wire s_arrmul12_fa4_11_and1;
  wire s_arrmul12_fa4_11_or0;
  wire s_arrmul12_nand5_11;
  wire s_arrmul12_fa5_11_xor0;
  wire s_arrmul12_fa5_11_and0;
  wire s_arrmul12_fa5_11_xor1;
  wire s_arrmul12_fa5_11_and1;
  wire s_arrmul12_fa5_11_or0;
  wire s_arrmul12_nand6_11;
  wire s_arrmul12_fa6_11_xor0;
  wire s_arrmul12_fa6_11_and0;
  wire s_arrmul12_fa6_11_xor1;
  wire s_arrmul12_fa6_11_and1;
  wire s_arrmul12_fa6_11_or0;
  wire s_arrmul12_nand7_11;
  wire s_arrmul12_fa7_11_xor0;
  wire s_arrmul12_fa7_11_and0;
  wire s_arrmul12_fa7_11_xor1;
  wire s_arrmul12_fa7_11_and1;
  wire s_arrmul12_fa7_11_or0;
  wire s_arrmul12_nand8_11;
  wire s_arrmul12_fa8_11_xor0;
  wire s_arrmul12_fa8_11_and0;
  wire s_arrmul12_fa8_11_xor1;
  wire s_arrmul12_fa8_11_and1;
  wire s_arrmul12_fa8_11_or0;
  wire s_arrmul12_nand9_11;
  wire s_arrmul12_fa9_11_xor0;
  wire s_arrmul12_fa9_11_and0;
  wire s_arrmul12_fa9_11_xor1;
  wire s_arrmul12_fa9_11_and1;
  wire s_arrmul12_fa9_11_or0;
  wire s_arrmul12_nand10_11;
  wire s_arrmul12_fa10_11_xor0;
  wire s_arrmul12_fa10_11_and0;
  wire s_arrmul12_fa10_11_xor1;
  wire s_arrmul12_fa10_11_and1;
  wire s_arrmul12_fa10_11_or0;
  wire s_arrmul12_and11_11;
  wire s_arrmul12_fa11_11_xor0;
  wire s_arrmul12_fa11_11_and0;
  wire s_arrmul12_fa11_11_xor1;
  wire s_arrmul12_fa11_11_and1;
  wire s_arrmul12_fa11_11_or0;
  wire s_arrmul12_xor12_11;

  assign s_arrmul12_and0_0 = a[0] & b[0];
  assign s_arrmul12_and1_0 = a[1] & b[0];
  assign s_arrmul12_and2_0 = a[2] & b[0];
  assign s_arrmul12_and3_0 = a[3] & b[0];
  assign s_arrmul12_and4_0 = a[4] & b[0];
  assign s_arrmul12_and5_0 = a[5] & b[0];
  assign s_arrmul12_and6_0 = a[6] & b[0];
  assign s_arrmul12_and7_0 = a[7] & b[0];
  assign s_arrmul12_and8_0 = a[8] & b[0];
  assign s_arrmul12_and9_0 = a[9] & b[0];
  assign s_arrmul12_and10_0 = a[10] & b[0];
  assign s_arrmul12_nand11_0 = ~(a[11] & b[0]);
  assign s_arrmul12_and0_1 = a[0] & b[1];
  assign s_arrmul12_ha0_1_xor0 = s_arrmul12_and0_1 ^ s_arrmul12_and1_0;
  assign s_arrmul12_ha0_1_and0 = s_arrmul12_and0_1 & s_arrmul12_and1_0;
  assign s_arrmul12_and1_1 = a[1] & b[1];
  assign s_arrmul12_fa1_1_xor0 = s_arrmul12_and1_1 ^ s_arrmul12_and2_0;
  assign s_arrmul12_fa1_1_and0 = s_arrmul12_and1_1 & s_arrmul12_and2_0;
  assign s_arrmul12_fa1_1_xor1 = s_arrmul12_fa1_1_xor0 ^ s_arrmul12_ha0_1_and0;
  assign s_arrmul12_fa1_1_and1 = s_arrmul12_fa1_1_xor0 & s_arrmul12_ha0_1_and0;
  assign s_arrmul12_fa1_1_or0 = s_arrmul12_fa1_1_and0 | s_arrmul12_fa1_1_and1;
  assign s_arrmul12_and2_1 = a[2] & b[1];
  assign s_arrmul12_fa2_1_xor0 = s_arrmul12_and2_1 ^ s_arrmul12_and3_0;
  assign s_arrmul12_fa2_1_and0 = s_arrmul12_and2_1 & s_arrmul12_and3_0;
  assign s_arrmul12_fa2_1_xor1 = s_arrmul12_fa2_1_xor0 ^ s_arrmul12_fa1_1_or0;
  assign s_arrmul12_fa2_1_and1 = s_arrmul12_fa2_1_xor0 & s_arrmul12_fa1_1_or0;
  assign s_arrmul12_fa2_1_or0 = s_arrmul12_fa2_1_and0 | s_arrmul12_fa2_1_and1;
  assign s_arrmul12_and3_1 = a[3] & b[1];
  assign s_arrmul12_fa3_1_xor0 = s_arrmul12_and3_1 ^ s_arrmul12_and4_0;
  assign s_arrmul12_fa3_1_and0 = s_arrmul12_and3_1 & s_arrmul12_and4_0;
  assign s_arrmul12_fa3_1_xor1 = s_arrmul12_fa3_1_xor0 ^ s_arrmul12_fa2_1_or0;
  assign s_arrmul12_fa3_1_and1 = s_arrmul12_fa3_1_xor0 & s_arrmul12_fa2_1_or0;
  assign s_arrmul12_fa3_1_or0 = s_arrmul12_fa3_1_and0 | s_arrmul12_fa3_1_and1;
  assign s_arrmul12_and4_1 = a[4] & b[1];
  assign s_arrmul12_fa4_1_xor0 = s_arrmul12_and4_1 ^ s_arrmul12_and5_0;
  assign s_arrmul12_fa4_1_and0 = s_arrmul12_and4_1 & s_arrmul12_and5_0;
  assign s_arrmul12_fa4_1_xor1 = s_arrmul12_fa4_1_xor0 ^ s_arrmul12_fa3_1_or0;
  assign s_arrmul12_fa4_1_and1 = s_arrmul12_fa4_1_xor0 & s_arrmul12_fa3_1_or0;
  assign s_arrmul12_fa4_1_or0 = s_arrmul12_fa4_1_and0 | s_arrmul12_fa4_1_and1;
  assign s_arrmul12_and5_1 = a[5] & b[1];
  assign s_arrmul12_fa5_1_xor0 = s_arrmul12_and5_1 ^ s_arrmul12_and6_0;
  assign s_arrmul12_fa5_1_and0 = s_arrmul12_and5_1 & s_arrmul12_and6_0;
  assign s_arrmul12_fa5_1_xor1 = s_arrmul12_fa5_1_xor0 ^ s_arrmul12_fa4_1_or0;
  assign s_arrmul12_fa5_1_and1 = s_arrmul12_fa5_1_xor0 & s_arrmul12_fa4_1_or0;
  assign s_arrmul12_fa5_1_or0 = s_arrmul12_fa5_1_and0 | s_arrmul12_fa5_1_and1;
  assign s_arrmul12_and6_1 = a[6] & b[1];
  assign s_arrmul12_fa6_1_xor0 = s_arrmul12_and6_1 ^ s_arrmul12_and7_0;
  assign s_arrmul12_fa6_1_and0 = s_arrmul12_and6_1 & s_arrmul12_and7_0;
  assign s_arrmul12_fa6_1_xor1 = s_arrmul12_fa6_1_xor0 ^ s_arrmul12_fa5_1_or0;
  assign s_arrmul12_fa6_1_and1 = s_arrmul12_fa6_1_xor0 & s_arrmul12_fa5_1_or0;
  assign s_arrmul12_fa6_1_or0 = s_arrmul12_fa6_1_and0 | s_arrmul12_fa6_1_and1;
  assign s_arrmul12_and7_1 = a[7] & b[1];
  assign s_arrmul12_fa7_1_xor0 = s_arrmul12_and7_1 ^ s_arrmul12_and8_0;
  assign s_arrmul12_fa7_1_and0 = s_arrmul12_and7_1 & s_arrmul12_and8_0;
  assign s_arrmul12_fa7_1_xor1 = s_arrmul12_fa7_1_xor0 ^ s_arrmul12_fa6_1_or0;
  assign s_arrmul12_fa7_1_and1 = s_arrmul12_fa7_1_xor0 & s_arrmul12_fa6_1_or0;
  assign s_arrmul12_fa7_1_or0 = s_arrmul12_fa7_1_and0 | s_arrmul12_fa7_1_and1;
  assign s_arrmul12_and8_1 = a[8] & b[1];
  assign s_arrmul12_fa8_1_xor0 = s_arrmul12_and8_1 ^ s_arrmul12_and9_0;
  assign s_arrmul12_fa8_1_and0 = s_arrmul12_and8_1 & s_arrmul12_and9_0;
  assign s_arrmul12_fa8_1_xor1 = s_arrmul12_fa8_1_xor0 ^ s_arrmul12_fa7_1_or0;
  assign s_arrmul12_fa8_1_and1 = s_arrmul12_fa8_1_xor0 & s_arrmul12_fa7_1_or0;
  assign s_arrmul12_fa8_1_or0 = s_arrmul12_fa8_1_and0 | s_arrmul12_fa8_1_and1;
  assign s_arrmul12_and9_1 = a[9] & b[1];
  assign s_arrmul12_fa9_1_xor0 = s_arrmul12_and9_1 ^ s_arrmul12_and10_0;
  assign s_arrmul12_fa9_1_and0 = s_arrmul12_and9_1 & s_arrmul12_and10_0;
  assign s_arrmul12_fa9_1_xor1 = s_arrmul12_fa9_1_xor0 ^ s_arrmul12_fa8_1_or0;
  assign s_arrmul12_fa9_1_and1 = s_arrmul12_fa9_1_xor0 & s_arrmul12_fa8_1_or0;
  assign s_arrmul12_fa9_1_or0 = s_arrmul12_fa9_1_and0 | s_arrmul12_fa9_1_and1;
  assign s_arrmul12_and10_1 = a[10] & b[1];
  assign s_arrmul12_fa10_1_xor0 = s_arrmul12_and10_1 ^ s_arrmul12_nand11_0;
  assign s_arrmul12_fa10_1_and0 = s_arrmul12_and10_1 & s_arrmul12_nand11_0;
  assign s_arrmul12_fa10_1_xor1 = s_arrmul12_fa10_1_xor0 ^ s_arrmul12_fa9_1_or0;
  assign s_arrmul12_fa10_1_and1 = s_arrmul12_fa10_1_xor0 & s_arrmul12_fa9_1_or0;
  assign s_arrmul12_fa10_1_or0 = s_arrmul12_fa10_1_and0 | s_arrmul12_fa10_1_and1;
  assign s_arrmul12_nand11_1 = ~(a[11] & b[1]);
  assign s_arrmul12_fa11_1_xor0 = ~s_arrmul12_nand11_1;
  assign s_arrmul12_fa11_1_xor1 = s_arrmul12_fa11_1_xor0 ^ s_arrmul12_fa10_1_or0;
  assign s_arrmul12_fa11_1_and1 = s_arrmul12_fa11_1_xor0 & s_arrmul12_fa10_1_or0;
  assign s_arrmul12_fa11_1_or0 = s_arrmul12_nand11_1 | s_arrmul12_fa11_1_and1;
  assign s_arrmul12_and0_2 = a[0] & b[2];
  assign s_arrmul12_ha0_2_xor0 = s_arrmul12_and0_2 ^ s_arrmul12_fa1_1_xor1;
  assign s_arrmul12_ha0_2_and0 = s_arrmul12_and0_2 & s_arrmul12_fa1_1_xor1;
  assign s_arrmul12_and1_2 = a[1] & b[2];
  assign s_arrmul12_fa1_2_xor0 = s_arrmul12_and1_2 ^ s_arrmul12_fa2_1_xor1;
  assign s_arrmul12_fa1_2_and0 = s_arrmul12_and1_2 & s_arrmul12_fa2_1_xor1;
  assign s_arrmul12_fa1_2_xor1 = s_arrmul12_fa1_2_xor0 ^ s_arrmul12_ha0_2_and0;
  assign s_arrmul12_fa1_2_and1 = s_arrmul12_fa1_2_xor0 & s_arrmul12_ha0_2_and0;
  assign s_arrmul12_fa1_2_or0 = s_arrmul12_fa1_2_and0 | s_arrmul12_fa1_2_and1;
  assign s_arrmul12_and2_2 = a[2] & b[2];
  assign s_arrmul12_fa2_2_xor0 = s_arrmul12_and2_2 ^ s_arrmul12_fa3_1_xor1;
  assign s_arrmul12_fa2_2_and0 = s_arrmul12_and2_2 & s_arrmul12_fa3_1_xor1;
  assign s_arrmul12_fa2_2_xor1 = s_arrmul12_fa2_2_xor0 ^ s_arrmul12_fa1_2_or0;
  assign s_arrmul12_fa2_2_and1 = s_arrmul12_fa2_2_xor0 & s_arrmul12_fa1_2_or0;
  assign s_arrmul12_fa2_2_or0 = s_arrmul12_fa2_2_and0 | s_arrmul12_fa2_2_and1;
  assign s_arrmul12_and3_2 = a[3] & b[2];
  assign s_arrmul12_fa3_2_xor0 = s_arrmul12_and3_2 ^ s_arrmul12_fa4_1_xor1;
  assign s_arrmul12_fa3_2_and0 = s_arrmul12_and3_2 & s_arrmul12_fa4_1_xor1;
  assign s_arrmul12_fa3_2_xor1 = s_arrmul12_fa3_2_xor0 ^ s_arrmul12_fa2_2_or0;
  assign s_arrmul12_fa3_2_and1 = s_arrmul12_fa3_2_xor0 & s_arrmul12_fa2_2_or0;
  assign s_arrmul12_fa3_2_or0 = s_arrmul12_fa3_2_and0 | s_arrmul12_fa3_2_and1;
  assign s_arrmul12_and4_2 = a[4] & b[2];
  assign s_arrmul12_fa4_2_xor0 = s_arrmul12_and4_2 ^ s_arrmul12_fa5_1_xor1;
  assign s_arrmul12_fa4_2_and0 = s_arrmul12_and4_2 & s_arrmul12_fa5_1_xor1;
  assign s_arrmul12_fa4_2_xor1 = s_arrmul12_fa4_2_xor0 ^ s_arrmul12_fa3_2_or0;
  assign s_arrmul12_fa4_2_and1 = s_arrmul12_fa4_2_xor0 & s_arrmul12_fa3_2_or0;
  assign s_arrmul12_fa4_2_or0 = s_arrmul12_fa4_2_and0 | s_arrmul12_fa4_2_and1;
  assign s_arrmul12_and5_2 = a[5] & b[2];
  assign s_arrmul12_fa5_2_xor0 = s_arrmul12_and5_2 ^ s_arrmul12_fa6_1_xor1;
  assign s_arrmul12_fa5_2_and0 = s_arrmul12_and5_2 & s_arrmul12_fa6_1_xor1;
  assign s_arrmul12_fa5_2_xor1 = s_arrmul12_fa5_2_xor0 ^ s_arrmul12_fa4_2_or0;
  assign s_arrmul12_fa5_2_and1 = s_arrmul12_fa5_2_xor0 & s_arrmul12_fa4_2_or0;
  assign s_arrmul12_fa5_2_or0 = s_arrmul12_fa5_2_and0 | s_arrmul12_fa5_2_and1;
  assign s_arrmul12_and6_2 = a[6] & b[2];
  assign s_arrmul12_fa6_2_xor0 = s_arrmul12_and6_2 ^ s_arrmul12_fa7_1_xor1;
  assign s_arrmul12_fa6_2_and0 = s_arrmul12_and6_2 & s_arrmul12_fa7_1_xor1;
  assign s_arrmul12_fa6_2_xor1 = s_arrmul12_fa6_2_xor0 ^ s_arrmul12_fa5_2_or0;
  assign s_arrmul12_fa6_2_and1 = s_arrmul12_fa6_2_xor0 & s_arrmul12_fa5_2_or0;
  assign s_arrmul12_fa6_2_or0 = s_arrmul12_fa6_2_and0 | s_arrmul12_fa6_2_and1;
  assign s_arrmul12_and7_2 = a[7] & b[2];
  assign s_arrmul12_fa7_2_xor0 = s_arrmul12_and7_2 ^ s_arrmul12_fa8_1_xor1;
  assign s_arrmul12_fa7_2_and0 = s_arrmul12_and7_2 & s_arrmul12_fa8_1_xor1;
  assign s_arrmul12_fa7_2_xor1 = s_arrmul12_fa7_2_xor0 ^ s_arrmul12_fa6_2_or0;
  assign s_arrmul12_fa7_2_and1 = s_arrmul12_fa7_2_xor0 & s_arrmul12_fa6_2_or0;
  assign s_arrmul12_fa7_2_or0 = s_arrmul12_fa7_2_and0 | s_arrmul12_fa7_2_and1;
  assign s_arrmul12_and8_2 = a[8] & b[2];
  assign s_arrmul12_fa8_2_xor0 = s_arrmul12_and8_2 ^ s_arrmul12_fa9_1_xor1;
  assign s_arrmul12_fa8_2_and0 = s_arrmul12_and8_2 & s_arrmul12_fa9_1_xor1;
  assign s_arrmul12_fa8_2_xor1 = s_arrmul12_fa8_2_xor0 ^ s_arrmul12_fa7_2_or0;
  assign s_arrmul12_fa8_2_and1 = s_arrmul12_fa8_2_xor0 & s_arrmul12_fa7_2_or0;
  assign s_arrmul12_fa8_2_or0 = s_arrmul12_fa8_2_and0 | s_arrmul12_fa8_2_and1;
  assign s_arrmul12_and9_2 = a[9] & b[2];
  assign s_arrmul12_fa9_2_xor0 = s_arrmul12_and9_2 ^ s_arrmul12_fa10_1_xor1;
  assign s_arrmul12_fa9_2_and0 = s_arrmul12_and9_2 & s_arrmul12_fa10_1_xor1;
  assign s_arrmul12_fa9_2_xor1 = s_arrmul12_fa9_2_xor0 ^ s_arrmul12_fa8_2_or0;
  assign s_arrmul12_fa9_2_and1 = s_arrmul12_fa9_2_xor0 & s_arrmul12_fa8_2_or0;
  assign s_arrmul12_fa9_2_or0 = s_arrmul12_fa9_2_and0 | s_arrmul12_fa9_2_and1;
  assign s_arrmul12_and10_2 = a[10] & b[2];
  assign s_arrmul12_fa10_2_xor0 = s_arrmul12_and10_2 ^ s_arrmul12_fa11_1_xor1;
  assign s_arrmul12_fa10_2_and0 = s_arrmul12_and10_2 & s_arrmul12_fa11_1_xor1;
  assign s_arrmul12_fa10_2_xor1 = s_arrmul12_fa10_2_xor0 ^ s_arrmul12_fa9_2_or0;
  assign s_arrmul12_fa10_2_and1 = s_arrmul12_fa10_2_xor0 & s_arrmul12_fa9_2_or0;
  assign s_arrmul12_fa10_2_or0 = s_arrmul12_fa10_2_and0 | s_arrmul12_fa10_2_and1;
  assign s_arrmul12_nand11_2 = ~(a[11] & b[2]);
  assign s_arrmul12_fa11_2_xor0 = s_arrmul12_nand11_2 ^ s_arrmul12_fa11_1_or0;
  assign s_arrmul12_fa11_2_and0 = s_arrmul12_nand11_2 & s_arrmul12_fa11_1_or0;
  assign s_arrmul12_fa11_2_xor1 = s_arrmul12_fa11_2_xor0 ^ s_arrmul12_fa10_2_or0;
  assign s_arrmul12_fa11_2_and1 = s_arrmul12_fa11_2_xor0 & s_arrmul12_fa10_2_or0;
  assign s_arrmul12_fa11_2_or0 = s_arrmul12_fa11_2_and0 | s_arrmul12_fa11_2_and1;
  assign s_arrmul12_and0_3 = a[0] & b[3];
  assign s_arrmul12_ha0_3_xor0 = s_arrmul12_and0_3 ^ s_arrmul12_fa1_2_xor1;
  assign s_arrmul12_ha0_3_and0 = s_arrmul12_and0_3 & s_arrmul12_fa1_2_xor1;
  assign s_arrmul12_and1_3 = a[1] & b[3];
  assign s_arrmul12_fa1_3_xor0 = s_arrmul12_and1_3 ^ s_arrmul12_fa2_2_xor1;
  assign s_arrmul12_fa1_3_and0 = s_arrmul12_and1_3 & s_arrmul12_fa2_2_xor1;
  assign s_arrmul12_fa1_3_xor1 = s_arrmul12_fa1_3_xor0 ^ s_arrmul12_ha0_3_and0;
  assign s_arrmul12_fa1_3_and1 = s_arrmul12_fa1_3_xor0 & s_arrmul12_ha0_3_and0;
  assign s_arrmul12_fa1_3_or0 = s_arrmul12_fa1_3_and0 | s_arrmul12_fa1_3_and1;
  assign s_arrmul12_and2_3 = a[2] & b[3];
  assign s_arrmul12_fa2_3_xor0 = s_arrmul12_and2_3 ^ s_arrmul12_fa3_2_xor1;
  assign s_arrmul12_fa2_3_and0 = s_arrmul12_and2_3 & s_arrmul12_fa3_2_xor1;
  assign s_arrmul12_fa2_3_xor1 = s_arrmul12_fa2_3_xor0 ^ s_arrmul12_fa1_3_or0;
  assign s_arrmul12_fa2_3_and1 = s_arrmul12_fa2_3_xor0 & s_arrmul12_fa1_3_or0;
  assign s_arrmul12_fa2_3_or0 = s_arrmul12_fa2_3_and0 | s_arrmul12_fa2_3_and1;
  assign s_arrmul12_and3_3 = a[3] & b[3];
  assign s_arrmul12_fa3_3_xor0 = s_arrmul12_and3_3 ^ s_arrmul12_fa4_2_xor1;
  assign s_arrmul12_fa3_3_and0 = s_arrmul12_and3_3 & s_arrmul12_fa4_2_xor1;
  assign s_arrmul12_fa3_3_xor1 = s_arrmul12_fa3_3_xor0 ^ s_arrmul12_fa2_3_or0;
  assign s_arrmul12_fa3_3_and1 = s_arrmul12_fa3_3_xor0 & s_arrmul12_fa2_3_or0;
  assign s_arrmul12_fa3_3_or0 = s_arrmul12_fa3_3_and0 | s_arrmul12_fa3_3_and1;
  assign s_arrmul12_and4_3 = a[4] & b[3];
  assign s_arrmul12_fa4_3_xor0 = s_arrmul12_and4_3 ^ s_arrmul12_fa5_2_xor1;
  assign s_arrmul12_fa4_3_and0 = s_arrmul12_and4_3 & s_arrmul12_fa5_2_xor1;
  assign s_arrmul12_fa4_3_xor1 = s_arrmul12_fa4_3_xor0 ^ s_arrmul12_fa3_3_or0;
  assign s_arrmul12_fa4_3_and1 = s_arrmul12_fa4_3_xor0 & s_arrmul12_fa3_3_or0;
  assign s_arrmul12_fa4_3_or0 = s_arrmul12_fa4_3_and0 | s_arrmul12_fa4_3_and1;
  assign s_arrmul12_and5_3 = a[5] & b[3];
  assign s_arrmul12_fa5_3_xor0 = s_arrmul12_and5_3 ^ s_arrmul12_fa6_2_xor1;
  assign s_arrmul12_fa5_3_and0 = s_arrmul12_and5_3 & s_arrmul12_fa6_2_xor1;
  assign s_arrmul12_fa5_3_xor1 = s_arrmul12_fa5_3_xor0 ^ s_arrmul12_fa4_3_or0;
  assign s_arrmul12_fa5_3_and1 = s_arrmul12_fa5_3_xor0 & s_arrmul12_fa4_3_or0;
  assign s_arrmul12_fa5_3_or0 = s_arrmul12_fa5_3_and0 | s_arrmul12_fa5_3_and1;
  assign s_arrmul12_and6_3 = a[6] & b[3];
  assign s_arrmul12_fa6_3_xor0 = s_arrmul12_and6_3 ^ s_arrmul12_fa7_2_xor1;
  assign s_arrmul12_fa6_3_and0 = s_arrmul12_and6_3 & s_arrmul12_fa7_2_xor1;
  assign s_arrmul12_fa6_3_xor1 = s_arrmul12_fa6_3_xor0 ^ s_arrmul12_fa5_3_or0;
  assign s_arrmul12_fa6_3_and1 = s_arrmul12_fa6_3_xor0 & s_arrmul12_fa5_3_or0;
  assign s_arrmul12_fa6_3_or0 = s_arrmul12_fa6_3_and0 | s_arrmul12_fa6_3_and1;
  assign s_arrmul12_and7_3 = a[7] & b[3];
  assign s_arrmul12_fa7_3_xor0 = s_arrmul12_and7_3 ^ s_arrmul12_fa8_2_xor1;
  assign s_arrmul12_fa7_3_and0 = s_arrmul12_and7_3 & s_arrmul12_fa8_2_xor1;
  assign s_arrmul12_fa7_3_xor1 = s_arrmul12_fa7_3_xor0 ^ s_arrmul12_fa6_3_or0;
  assign s_arrmul12_fa7_3_and1 = s_arrmul12_fa7_3_xor0 & s_arrmul12_fa6_3_or0;
  assign s_arrmul12_fa7_3_or0 = s_arrmul12_fa7_3_and0 | s_arrmul12_fa7_3_and1;
  assign s_arrmul12_and8_3 = a[8] & b[3];
  assign s_arrmul12_fa8_3_xor0 = s_arrmul12_and8_3 ^ s_arrmul12_fa9_2_xor1;
  assign s_arrmul12_fa8_3_and0 = s_arrmul12_and8_3 & s_arrmul12_fa9_2_xor1;
  assign s_arrmul12_fa8_3_xor1 = s_arrmul12_fa8_3_xor0 ^ s_arrmul12_fa7_3_or0;
  assign s_arrmul12_fa8_3_and1 = s_arrmul12_fa8_3_xor0 & s_arrmul12_fa7_3_or0;
  assign s_arrmul12_fa8_3_or0 = s_arrmul12_fa8_3_and0 | s_arrmul12_fa8_3_and1;
  assign s_arrmul12_and9_3 = a[9] & b[3];
  assign s_arrmul12_fa9_3_xor0 = s_arrmul12_and9_3 ^ s_arrmul12_fa10_2_xor1;
  assign s_arrmul12_fa9_3_and0 = s_arrmul12_and9_3 & s_arrmul12_fa10_2_xor1;
  assign s_arrmul12_fa9_3_xor1 = s_arrmul12_fa9_3_xor0 ^ s_arrmul12_fa8_3_or0;
  assign s_arrmul12_fa9_3_and1 = s_arrmul12_fa9_3_xor0 & s_arrmul12_fa8_3_or0;
  assign s_arrmul12_fa9_3_or0 = s_arrmul12_fa9_3_and0 | s_arrmul12_fa9_3_and1;
  assign s_arrmul12_and10_3 = a[10] & b[3];
  assign s_arrmul12_fa10_3_xor0 = s_arrmul12_and10_3 ^ s_arrmul12_fa11_2_xor1;
  assign s_arrmul12_fa10_3_and0 = s_arrmul12_and10_3 & s_arrmul12_fa11_2_xor1;
  assign s_arrmul12_fa10_3_xor1 = s_arrmul12_fa10_3_xor0 ^ s_arrmul12_fa9_3_or0;
  assign s_arrmul12_fa10_3_and1 = s_arrmul12_fa10_3_xor0 & s_arrmul12_fa9_3_or0;
  assign s_arrmul12_fa10_3_or0 = s_arrmul12_fa10_3_and0 | s_arrmul12_fa10_3_and1;
  assign s_arrmul12_nand11_3 = ~(a[11] & b[3]);
  assign s_arrmul12_fa11_3_xor0 = s_arrmul12_nand11_3 ^ s_arrmul12_fa11_2_or0;
  assign s_arrmul12_fa11_3_and0 = s_arrmul12_nand11_3 & s_arrmul12_fa11_2_or0;
  assign s_arrmul12_fa11_3_xor1 = s_arrmul12_fa11_3_xor0 ^ s_arrmul12_fa10_3_or0;
  assign s_arrmul12_fa11_3_and1 = s_arrmul12_fa11_3_xor0 & s_arrmul12_fa10_3_or0;
  assign s_arrmul12_fa11_3_or0 = s_arrmul12_fa11_3_and0 | s_arrmul12_fa11_3_and1;
  assign s_arrmul12_and0_4 = a[0] & b[4];
  assign s_arrmul12_ha0_4_xor0 = s_arrmul12_and0_4 ^ s_arrmul12_fa1_3_xor1;
  assign s_arrmul12_ha0_4_and0 = s_arrmul12_and0_4 & s_arrmul12_fa1_3_xor1;
  assign s_arrmul12_and1_4 = a[1] & b[4];
  assign s_arrmul12_fa1_4_xor0 = s_arrmul12_and1_4 ^ s_arrmul12_fa2_3_xor1;
  assign s_arrmul12_fa1_4_and0 = s_arrmul12_and1_4 & s_arrmul12_fa2_3_xor1;
  assign s_arrmul12_fa1_4_xor1 = s_arrmul12_fa1_4_xor0 ^ s_arrmul12_ha0_4_and0;
  assign s_arrmul12_fa1_4_and1 = s_arrmul12_fa1_4_xor0 & s_arrmul12_ha0_4_and0;
  assign s_arrmul12_fa1_4_or0 = s_arrmul12_fa1_4_and0 | s_arrmul12_fa1_4_and1;
  assign s_arrmul12_and2_4 = a[2] & b[4];
  assign s_arrmul12_fa2_4_xor0 = s_arrmul12_and2_4 ^ s_arrmul12_fa3_3_xor1;
  assign s_arrmul12_fa2_4_and0 = s_arrmul12_and2_4 & s_arrmul12_fa3_3_xor1;
  assign s_arrmul12_fa2_4_xor1 = s_arrmul12_fa2_4_xor0 ^ s_arrmul12_fa1_4_or0;
  assign s_arrmul12_fa2_4_and1 = s_arrmul12_fa2_4_xor0 & s_arrmul12_fa1_4_or0;
  assign s_arrmul12_fa2_4_or0 = s_arrmul12_fa2_4_and0 | s_arrmul12_fa2_4_and1;
  assign s_arrmul12_and3_4 = a[3] & b[4];
  assign s_arrmul12_fa3_4_xor0 = s_arrmul12_and3_4 ^ s_arrmul12_fa4_3_xor1;
  assign s_arrmul12_fa3_4_and0 = s_arrmul12_and3_4 & s_arrmul12_fa4_3_xor1;
  assign s_arrmul12_fa3_4_xor1 = s_arrmul12_fa3_4_xor0 ^ s_arrmul12_fa2_4_or0;
  assign s_arrmul12_fa3_4_and1 = s_arrmul12_fa3_4_xor0 & s_arrmul12_fa2_4_or0;
  assign s_arrmul12_fa3_4_or0 = s_arrmul12_fa3_4_and0 | s_arrmul12_fa3_4_and1;
  assign s_arrmul12_and4_4 = a[4] & b[4];
  assign s_arrmul12_fa4_4_xor0 = s_arrmul12_and4_4 ^ s_arrmul12_fa5_3_xor1;
  assign s_arrmul12_fa4_4_and0 = s_arrmul12_and4_4 & s_arrmul12_fa5_3_xor1;
  assign s_arrmul12_fa4_4_xor1 = s_arrmul12_fa4_4_xor0 ^ s_arrmul12_fa3_4_or0;
  assign s_arrmul12_fa4_4_and1 = s_arrmul12_fa4_4_xor0 & s_arrmul12_fa3_4_or0;
  assign s_arrmul12_fa4_4_or0 = s_arrmul12_fa4_4_and0 | s_arrmul12_fa4_4_and1;
  assign s_arrmul12_and5_4 = a[5] & b[4];
  assign s_arrmul12_fa5_4_xor0 = s_arrmul12_and5_4 ^ s_arrmul12_fa6_3_xor1;
  assign s_arrmul12_fa5_4_and0 = s_arrmul12_and5_4 & s_arrmul12_fa6_3_xor1;
  assign s_arrmul12_fa5_4_xor1 = s_arrmul12_fa5_4_xor0 ^ s_arrmul12_fa4_4_or0;
  assign s_arrmul12_fa5_4_and1 = s_arrmul12_fa5_4_xor0 & s_arrmul12_fa4_4_or0;
  assign s_arrmul12_fa5_4_or0 = s_arrmul12_fa5_4_and0 | s_arrmul12_fa5_4_and1;
  assign s_arrmul12_and6_4 = a[6] & b[4];
  assign s_arrmul12_fa6_4_xor0 = s_arrmul12_and6_4 ^ s_arrmul12_fa7_3_xor1;
  assign s_arrmul12_fa6_4_and0 = s_arrmul12_and6_4 & s_arrmul12_fa7_3_xor1;
  assign s_arrmul12_fa6_4_xor1 = s_arrmul12_fa6_4_xor0 ^ s_arrmul12_fa5_4_or0;
  assign s_arrmul12_fa6_4_and1 = s_arrmul12_fa6_4_xor0 & s_arrmul12_fa5_4_or0;
  assign s_arrmul12_fa6_4_or0 = s_arrmul12_fa6_4_and0 | s_arrmul12_fa6_4_and1;
  assign s_arrmul12_and7_4 = a[7] & b[4];
  assign s_arrmul12_fa7_4_xor0 = s_arrmul12_and7_4 ^ s_arrmul12_fa8_3_xor1;
  assign s_arrmul12_fa7_4_and0 = s_arrmul12_and7_4 & s_arrmul12_fa8_3_xor1;
  assign s_arrmul12_fa7_4_xor1 = s_arrmul12_fa7_4_xor0 ^ s_arrmul12_fa6_4_or0;
  assign s_arrmul12_fa7_4_and1 = s_arrmul12_fa7_4_xor0 & s_arrmul12_fa6_4_or0;
  assign s_arrmul12_fa7_4_or0 = s_arrmul12_fa7_4_and0 | s_arrmul12_fa7_4_and1;
  assign s_arrmul12_and8_4 = a[8] & b[4];
  assign s_arrmul12_fa8_4_xor0 = s_arrmul12_and8_4 ^ s_arrmul12_fa9_3_xor1;
  assign s_arrmul12_fa8_4_and0 = s_arrmul12_and8_4 & s_arrmul12_fa9_3_xor1;
  assign s_arrmul12_fa8_4_xor1 = s_arrmul12_fa8_4_xor0 ^ s_arrmul12_fa7_4_or0;
  assign s_arrmul12_fa8_4_and1 = s_arrmul12_fa8_4_xor0 & s_arrmul12_fa7_4_or0;
  assign s_arrmul12_fa8_4_or0 = s_arrmul12_fa8_4_and0 | s_arrmul12_fa8_4_and1;
  assign s_arrmul12_and9_4 = a[9] & b[4];
  assign s_arrmul12_fa9_4_xor0 = s_arrmul12_and9_4 ^ s_arrmul12_fa10_3_xor1;
  assign s_arrmul12_fa9_4_and0 = s_arrmul12_and9_4 & s_arrmul12_fa10_3_xor1;
  assign s_arrmul12_fa9_4_xor1 = s_arrmul12_fa9_4_xor0 ^ s_arrmul12_fa8_4_or0;
  assign s_arrmul12_fa9_4_and1 = s_arrmul12_fa9_4_xor0 & s_arrmul12_fa8_4_or0;
  assign s_arrmul12_fa9_4_or0 = s_arrmul12_fa9_4_and0 | s_arrmul12_fa9_4_and1;
  assign s_arrmul12_and10_4 = a[10] & b[4];
  assign s_arrmul12_fa10_4_xor0 = s_arrmul12_and10_4 ^ s_arrmul12_fa11_3_xor1;
  assign s_arrmul12_fa10_4_and0 = s_arrmul12_and10_4 & s_arrmul12_fa11_3_xor1;
  assign s_arrmul12_fa10_4_xor1 = s_arrmul12_fa10_4_xor0 ^ s_arrmul12_fa9_4_or0;
  assign s_arrmul12_fa10_4_and1 = s_arrmul12_fa10_4_xor0 & s_arrmul12_fa9_4_or0;
  assign s_arrmul12_fa10_4_or0 = s_arrmul12_fa10_4_and0 | s_arrmul12_fa10_4_and1;
  assign s_arrmul12_nand11_4 = ~(a[11] & b[4]);
  assign s_arrmul12_fa11_4_xor0 = s_arrmul12_nand11_4 ^ s_arrmul12_fa11_3_or0;
  assign s_arrmul12_fa11_4_and0 = s_arrmul12_nand11_4 & s_arrmul12_fa11_3_or0;
  assign s_arrmul12_fa11_4_xor1 = s_arrmul12_fa11_4_xor0 ^ s_arrmul12_fa10_4_or0;
  assign s_arrmul12_fa11_4_and1 = s_arrmul12_fa11_4_xor0 & s_arrmul12_fa10_4_or0;
  assign s_arrmul12_fa11_4_or0 = s_arrmul12_fa11_4_and0 | s_arrmul12_fa11_4_and1;
  assign s_arrmul12_and0_5 = a[0] & b[5];
  assign s_arrmul12_ha0_5_xor0 = s_arrmul12_and0_5 ^ s_arrmul12_fa1_4_xor1;
  assign s_arrmul12_ha0_5_and0 = s_arrmul12_and0_5 & s_arrmul12_fa1_4_xor1;
  assign s_arrmul12_and1_5 = a[1] & b[5];
  assign s_arrmul12_fa1_5_xor0 = s_arrmul12_and1_5 ^ s_arrmul12_fa2_4_xor1;
  assign s_arrmul12_fa1_5_and0 = s_arrmul12_and1_5 & s_arrmul12_fa2_4_xor1;
  assign s_arrmul12_fa1_5_xor1 = s_arrmul12_fa1_5_xor0 ^ s_arrmul12_ha0_5_and0;
  assign s_arrmul12_fa1_5_and1 = s_arrmul12_fa1_5_xor0 & s_arrmul12_ha0_5_and0;
  assign s_arrmul12_fa1_5_or0 = s_arrmul12_fa1_5_and0 | s_arrmul12_fa1_5_and1;
  assign s_arrmul12_and2_5 = a[2] & b[5];
  assign s_arrmul12_fa2_5_xor0 = s_arrmul12_and2_5 ^ s_arrmul12_fa3_4_xor1;
  assign s_arrmul12_fa2_5_and0 = s_arrmul12_and2_5 & s_arrmul12_fa3_4_xor1;
  assign s_arrmul12_fa2_5_xor1 = s_arrmul12_fa2_5_xor0 ^ s_arrmul12_fa1_5_or0;
  assign s_arrmul12_fa2_5_and1 = s_arrmul12_fa2_5_xor0 & s_arrmul12_fa1_5_or0;
  assign s_arrmul12_fa2_5_or0 = s_arrmul12_fa2_5_and0 | s_arrmul12_fa2_5_and1;
  assign s_arrmul12_and3_5 = a[3] & b[5];
  assign s_arrmul12_fa3_5_xor0 = s_arrmul12_and3_5 ^ s_arrmul12_fa4_4_xor1;
  assign s_arrmul12_fa3_5_and0 = s_arrmul12_and3_5 & s_arrmul12_fa4_4_xor1;
  assign s_arrmul12_fa3_5_xor1 = s_arrmul12_fa3_5_xor0 ^ s_arrmul12_fa2_5_or0;
  assign s_arrmul12_fa3_5_and1 = s_arrmul12_fa3_5_xor0 & s_arrmul12_fa2_5_or0;
  assign s_arrmul12_fa3_5_or0 = s_arrmul12_fa3_5_and0 | s_arrmul12_fa3_5_and1;
  assign s_arrmul12_and4_5 = a[4] & b[5];
  assign s_arrmul12_fa4_5_xor0 = s_arrmul12_and4_5 ^ s_arrmul12_fa5_4_xor1;
  assign s_arrmul12_fa4_5_and0 = s_arrmul12_and4_5 & s_arrmul12_fa5_4_xor1;
  assign s_arrmul12_fa4_5_xor1 = s_arrmul12_fa4_5_xor0 ^ s_arrmul12_fa3_5_or0;
  assign s_arrmul12_fa4_5_and1 = s_arrmul12_fa4_5_xor0 & s_arrmul12_fa3_5_or0;
  assign s_arrmul12_fa4_5_or0 = s_arrmul12_fa4_5_and0 | s_arrmul12_fa4_5_and1;
  assign s_arrmul12_and5_5 = a[5] & b[5];
  assign s_arrmul12_fa5_5_xor0 = s_arrmul12_and5_5 ^ s_arrmul12_fa6_4_xor1;
  assign s_arrmul12_fa5_5_and0 = s_arrmul12_and5_5 & s_arrmul12_fa6_4_xor1;
  assign s_arrmul12_fa5_5_xor1 = s_arrmul12_fa5_5_xor0 ^ s_arrmul12_fa4_5_or0;
  assign s_arrmul12_fa5_5_and1 = s_arrmul12_fa5_5_xor0 & s_arrmul12_fa4_5_or0;
  assign s_arrmul12_fa5_5_or0 = s_arrmul12_fa5_5_and0 | s_arrmul12_fa5_5_and1;
  assign s_arrmul12_and6_5 = a[6] & b[5];
  assign s_arrmul12_fa6_5_xor0 = s_arrmul12_and6_5 ^ s_arrmul12_fa7_4_xor1;
  assign s_arrmul12_fa6_5_and0 = s_arrmul12_and6_5 & s_arrmul12_fa7_4_xor1;
  assign s_arrmul12_fa6_5_xor1 = s_arrmul12_fa6_5_xor0 ^ s_arrmul12_fa5_5_or0;
  assign s_arrmul12_fa6_5_and1 = s_arrmul12_fa6_5_xor0 & s_arrmul12_fa5_5_or0;
  assign s_arrmul12_fa6_5_or0 = s_arrmul12_fa6_5_and0 | s_arrmul12_fa6_5_and1;
  assign s_arrmul12_and7_5 = a[7] & b[5];
  assign s_arrmul12_fa7_5_xor0 = s_arrmul12_and7_5 ^ s_arrmul12_fa8_4_xor1;
  assign s_arrmul12_fa7_5_and0 = s_arrmul12_and7_5 & s_arrmul12_fa8_4_xor1;
  assign s_arrmul12_fa7_5_xor1 = s_arrmul12_fa7_5_xor0 ^ s_arrmul12_fa6_5_or0;
  assign s_arrmul12_fa7_5_and1 = s_arrmul12_fa7_5_xor0 & s_arrmul12_fa6_5_or0;
  assign s_arrmul12_fa7_5_or0 = s_arrmul12_fa7_5_and0 | s_arrmul12_fa7_5_and1;
  assign s_arrmul12_and8_5 = a[8] & b[5];
  assign s_arrmul12_fa8_5_xor0 = s_arrmul12_and8_5 ^ s_arrmul12_fa9_4_xor1;
  assign s_arrmul12_fa8_5_and0 = s_arrmul12_and8_5 & s_arrmul12_fa9_4_xor1;
  assign s_arrmul12_fa8_5_xor1 = s_arrmul12_fa8_5_xor0 ^ s_arrmul12_fa7_5_or0;
  assign s_arrmul12_fa8_5_and1 = s_arrmul12_fa8_5_xor0 & s_arrmul12_fa7_5_or0;
  assign s_arrmul12_fa8_5_or0 = s_arrmul12_fa8_5_and0 | s_arrmul12_fa8_5_and1;
  assign s_arrmul12_and9_5 = a[9] & b[5];
  assign s_arrmul12_fa9_5_xor0 = s_arrmul12_and9_5 ^ s_arrmul12_fa10_4_xor1;
  assign s_arrmul12_fa9_5_and0 = s_arrmul12_and9_5 & s_arrmul12_fa10_4_xor1;
  assign s_arrmul12_fa9_5_xor1 = s_arrmul12_fa9_5_xor0 ^ s_arrmul12_fa8_5_or0;
  assign s_arrmul12_fa9_5_and1 = s_arrmul12_fa9_5_xor0 & s_arrmul12_fa8_5_or0;
  assign s_arrmul12_fa9_5_or0 = s_arrmul12_fa9_5_and0 | s_arrmul12_fa9_5_and1;
  assign s_arrmul12_and10_5 = a[10] & b[5];
  assign s_arrmul12_fa10_5_xor0 = s_arrmul12_and10_5 ^ s_arrmul12_fa11_4_xor1;
  assign s_arrmul12_fa10_5_and0 = s_arrmul12_and10_5 & s_arrmul12_fa11_4_xor1;
  assign s_arrmul12_fa10_5_xor1 = s_arrmul12_fa10_5_xor0 ^ s_arrmul12_fa9_5_or0;
  assign s_arrmul12_fa10_5_and1 = s_arrmul12_fa10_5_xor0 & s_arrmul12_fa9_5_or0;
  assign s_arrmul12_fa10_5_or0 = s_arrmul12_fa10_5_and0 | s_arrmul12_fa10_5_and1;
  assign s_arrmul12_nand11_5 = ~(a[11] & b[5]);
  assign s_arrmul12_fa11_5_xor0 = s_arrmul12_nand11_5 ^ s_arrmul12_fa11_4_or0;
  assign s_arrmul12_fa11_5_and0 = s_arrmul12_nand11_5 & s_arrmul12_fa11_4_or0;
  assign s_arrmul12_fa11_5_xor1 = s_arrmul12_fa11_5_xor0 ^ s_arrmul12_fa10_5_or0;
  assign s_arrmul12_fa11_5_and1 = s_arrmul12_fa11_5_xor0 & s_arrmul12_fa10_5_or0;
  assign s_arrmul12_fa11_5_or0 = s_arrmul12_fa11_5_and0 | s_arrmul12_fa11_5_and1;
  assign s_arrmul12_and0_6 = a[0] & b[6];
  assign s_arrmul12_ha0_6_xor0 = s_arrmul12_and0_6 ^ s_arrmul12_fa1_5_xor1;
  assign s_arrmul12_ha0_6_and0 = s_arrmul12_and0_6 & s_arrmul12_fa1_5_xor1;
  assign s_arrmul12_and1_6 = a[1] & b[6];
  assign s_arrmul12_fa1_6_xor0 = s_arrmul12_and1_6 ^ s_arrmul12_fa2_5_xor1;
  assign s_arrmul12_fa1_6_and0 = s_arrmul12_and1_6 & s_arrmul12_fa2_5_xor1;
  assign s_arrmul12_fa1_6_xor1 = s_arrmul12_fa1_6_xor0 ^ s_arrmul12_ha0_6_and0;
  assign s_arrmul12_fa1_6_and1 = s_arrmul12_fa1_6_xor0 & s_arrmul12_ha0_6_and0;
  assign s_arrmul12_fa1_6_or0 = s_arrmul12_fa1_6_and0 | s_arrmul12_fa1_6_and1;
  assign s_arrmul12_and2_6 = a[2] & b[6];
  assign s_arrmul12_fa2_6_xor0 = s_arrmul12_and2_6 ^ s_arrmul12_fa3_5_xor1;
  assign s_arrmul12_fa2_6_and0 = s_arrmul12_and2_6 & s_arrmul12_fa3_5_xor1;
  assign s_arrmul12_fa2_6_xor1 = s_arrmul12_fa2_6_xor0 ^ s_arrmul12_fa1_6_or0;
  assign s_arrmul12_fa2_6_and1 = s_arrmul12_fa2_6_xor0 & s_arrmul12_fa1_6_or0;
  assign s_arrmul12_fa2_6_or0 = s_arrmul12_fa2_6_and0 | s_arrmul12_fa2_6_and1;
  assign s_arrmul12_and3_6 = a[3] & b[6];
  assign s_arrmul12_fa3_6_xor0 = s_arrmul12_and3_6 ^ s_arrmul12_fa4_5_xor1;
  assign s_arrmul12_fa3_6_and0 = s_arrmul12_and3_6 & s_arrmul12_fa4_5_xor1;
  assign s_arrmul12_fa3_6_xor1 = s_arrmul12_fa3_6_xor0 ^ s_arrmul12_fa2_6_or0;
  assign s_arrmul12_fa3_6_and1 = s_arrmul12_fa3_6_xor0 & s_arrmul12_fa2_6_or0;
  assign s_arrmul12_fa3_6_or0 = s_arrmul12_fa3_6_and0 | s_arrmul12_fa3_6_and1;
  assign s_arrmul12_and4_6 = a[4] & b[6];
  assign s_arrmul12_fa4_6_xor0 = s_arrmul12_and4_6 ^ s_arrmul12_fa5_5_xor1;
  assign s_arrmul12_fa4_6_and0 = s_arrmul12_and4_6 & s_arrmul12_fa5_5_xor1;
  assign s_arrmul12_fa4_6_xor1 = s_arrmul12_fa4_6_xor0 ^ s_arrmul12_fa3_6_or0;
  assign s_arrmul12_fa4_6_and1 = s_arrmul12_fa4_6_xor0 & s_arrmul12_fa3_6_or0;
  assign s_arrmul12_fa4_6_or0 = s_arrmul12_fa4_6_and0 | s_arrmul12_fa4_6_and1;
  assign s_arrmul12_and5_6 = a[5] & b[6];
  assign s_arrmul12_fa5_6_xor0 = s_arrmul12_and5_6 ^ s_arrmul12_fa6_5_xor1;
  assign s_arrmul12_fa5_6_and0 = s_arrmul12_and5_6 & s_arrmul12_fa6_5_xor1;
  assign s_arrmul12_fa5_6_xor1 = s_arrmul12_fa5_6_xor0 ^ s_arrmul12_fa4_6_or0;
  assign s_arrmul12_fa5_6_and1 = s_arrmul12_fa5_6_xor0 & s_arrmul12_fa4_6_or0;
  assign s_arrmul12_fa5_6_or0 = s_arrmul12_fa5_6_and0 | s_arrmul12_fa5_6_and1;
  assign s_arrmul12_and6_6 = a[6] & b[6];
  assign s_arrmul12_fa6_6_xor0 = s_arrmul12_and6_6 ^ s_arrmul12_fa7_5_xor1;
  assign s_arrmul12_fa6_6_and0 = s_arrmul12_and6_6 & s_arrmul12_fa7_5_xor1;
  assign s_arrmul12_fa6_6_xor1 = s_arrmul12_fa6_6_xor0 ^ s_arrmul12_fa5_6_or0;
  assign s_arrmul12_fa6_6_and1 = s_arrmul12_fa6_6_xor0 & s_arrmul12_fa5_6_or0;
  assign s_arrmul12_fa6_6_or0 = s_arrmul12_fa6_6_and0 | s_arrmul12_fa6_6_and1;
  assign s_arrmul12_and7_6 = a[7] & b[6];
  assign s_arrmul12_fa7_6_xor0 = s_arrmul12_and7_6 ^ s_arrmul12_fa8_5_xor1;
  assign s_arrmul12_fa7_6_and0 = s_arrmul12_and7_6 & s_arrmul12_fa8_5_xor1;
  assign s_arrmul12_fa7_6_xor1 = s_arrmul12_fa7_6_xor0 ^ s_arrmul12_fa6_6_or0;
  assign s_arrmul12_fa7_6_and1 = s_arrmul12_fa7_6_xor0 & s_arrmul12_fa6_6_or0;
  assign s_arrmul12_fa7_6_or0 = s_arrmul12_fa7_6_and0 | s_arrmul12_fa7_6_and1;
  assign s_arrmul12_and8_6 = a[8] & b[6];
  assign s_arrmul12_fa8_6_xor0 = s_arrmul12_and8_6 ^ s_arrmul12_fa9_5_xor1;
  assign s_arrmul12_fa8_6_and0 = s_arrmul12_and8_6 & s_arrmul12_fa9_5_xor1;
  assign s_arrmul12_fa8_6_xor1 = s_arrmul12_fa8_6_xor0 ^ s_arrmul12_fa7_6_or0;
  assign s_arrmul12_fa8_6_and1 = s_arrmul12_fa8_6_xor0 & s_arrmul12_fa7_6_or0;
  assign s_arrmul12_fa8_6_or0 = s_arrmul12_fa8_6_and0 | s_arrmul12_fa8_6_and1;
  assign s_arrmul12_and9_6 = a[9] & b[6];
  assign s_arrmul12_fa9_6_xor0 = s_arrmul12_and9_6 ^ s_arrmul12_fa10_5_xor1;
  assign s_arrmul12_fa9_6_and0 = s_arrmul12_and9_6 & s_arrmul12_fa10_5_xor1;
  assign s_arrmul12_fa9_6_xor1 = s_arrmul12_fa9_6_xor0 ^ s_arrmul12_fa8_6_or0;
  assign s_arrmul12_fa9_6_and1 = s_arrmul12_fa9_6_xor0 & s_arrmul12_fa8_6_or0;
  assign s_arrmul12_fa9_6_or0 = s_arrmul12_fa9_6_and0 | s_arrmul12_fa9_6_and1;
  assign s_arrmul12_and10_6 = a[10] & b[6];
  assign s_arrmul12_fa10_6_xor0 = s_arrmul12_and10_6 ^ s_arrmul12_fa11_5_xor1;
  assign s_arrmul12_fa10_6_and0 = s_arrmul12_and10_6 & s_arrmul12_fa11_5_xor1;
  assign s_arrmul12_fa10_6_xor1 = s_arrmul12_fa10_6_xor0 ^ s_arrmul12_fa9_6_or0;
  assign s_arrmul12_fa10_6_and1 = s_arrmul12_fa10_6_xor0 & s_arrmul12_fa9_6_or0;
  assign s_arrmul12_fa10_6_or0 = s_arrmul12_fa10_6_and0 | s_arrmul12_fa10_6_and1;
  assign s_arrmul12_nand11_6 = ~(a[11] & b[6]);
  assign s_arrmul12_fa11_6_xor0 = s_arrmul12_nand11_6 ^ s_arrmul12_fa11_5_or0;
  assign s_arrmul12_fa11_6_and0 = s_arrmul12_nand11_6 & s_arrmul12_fa11_5_or0;
  assign s_arrmul12_fa11_6_xor1 = s_arrmul12_fa11_6_xor0 ^ s_arrmul12_fa10_6_or0;
  assign s_arrmul12_fa11_6_and1 = s_arrmul12_fa11_6_xor0 & s_arrmul12_fa10_6_or0;
  assign s_arrmul12_fa11_6_or0 = s_arrmul12_fa11_6_and0 | s_arrmul12_fa11_6_and1;
  assign s_arrmul12_and0_7 = a[0] & b[7];
  assign s_arrmul12_ha0_7_xor0 = s_arrmul12_and0_7 ^ s_arrmul12_fa1_6_xor1;
  assign s_arrmul12_ha0_7_and0 = s_arrmul12_and0_7 & s_arrmul12_fa1_6_xor1;
  assign s_arrmul12_and1_7 = a[1] & b[7];
  assign s_arrmul12_fa1_7_xor0 = s_arrmul12_and1_7 ^ s_arrmul12_fa2_6_xor1;
  assign s_arrmul12_fa1_7_and0 = s_arrmul12_and1_7 & s_arrmul12_fa2_6_xor1;
  assign s_arrmul12_fa1_7_xor1 = s_arrmul12_fa1_7_xor0 ^ s_arrmul12_ha0_7_and0;
  assign s_arrmul12_fa1_7_and1 = s_arrmul12_fa1_7_xor0 & s_arrmul12_ha0_7_and0;
  assign s_arrmul12_fa1_7_or0 = s_arrmul12_fa1_7_and0 | s_arrmul12_fa1_7_and1;
  assign s_arrmul12_and2_7 = a[2] & b[7];
  assign s_arrmul12_fa2_7_xor0 = s_arrmul12_and2_7 ^ s_arrmul12_fa3_6_xor1;
  assign s_arrmul12_fa2_7_and0 = s_arrmul12_and2_7 & s_arrmul12_fa3_6_xor1;
  assign s_arrmul12_fa2_7_xor1 = s_arrmul12_fa2_7_xor0 ^ s_arrmul12_fa1_7_or0;
  assign s_arrmul12_fa2_7_and1 = s_arrmul12_fa2_7_xor0 & s_arrmul12_fa1_7_or0;
  assign s_arrmul12_fa2_7_or0 = s_arrmul12_fa2_7_and0 | s_arrmul12_fa2_7_and1;
  assign s_arrmul12_and3_7 = a[3] & b[7];
  assign s_arrmul12_fa3_7_xor0 = s_arrmul12_and3_7 ^ s_arrmul12_fa4_6_xor1;
  assign s_arrmul12_fa3_7_and0 = s_arrmul12_and3_7 & s_arrmul12_fa4_6_xor1;
  assign s_arrmul12_fa3_7_xor1 = s_arrmul12_fa3_7_xor0 ^ s_arrmul12_fa2_7_or0;
  assign s_arrmul12_fa3_7_and1 = s_arrmul12_fa3_7_xor0 & s_arrmul12_fa2_7_or0;
  assign s_arrmul12_fa3_7_or0 = s_arrmul12_fa3_7_and0 | s_arrmul12_fa3_7_and1;
  assign s_arrmul12_and4_7 = a[4] & b[7];
  assign s_arrmul12_fa4_7_xor0 = s_arrmul12_and4_7 ^ s_arrmul12_fa5_6_xor1;
  assign s_arrmul12_fa4_7_and0 = s_arrmul12_and4_7 & s_arrmul12_fa5_6_xor1;
  assign s_arrmul12_fa4_7_xor1 = s_arrmul12_fa4_7_xor0 ^ s_arrmul12_fa3_7_or0;
  assign s_arrmul12_fa4_7_and1 = s_arrmul12_fa4_7_xor0 & s_arrmul12_fa3_7_or0;
  assign s_arrmul12_fa4_7_or0 = s_arrmul12_fa4_7_and0 | s_arrmul12_fa4_7_and1;
  assign s_arrmul12_and5_7 = a[5] & b[7];
  assign s_arrmul12_fa5_7_xor0 = s_arrmul12_and5_7 ^ s_arrmul12_fa6_6_xor1;
  assign s_arrmul12_fa5_7_and0 = s_arrmul12_and5_7 & s_arrmul12_fa6_6_xor1;
  assign s_arrmul12_fa5_7_xor1 = s_arrmul12_fa5_7_xor0 ^ s_arrmul12_fa4_7_or0;
  assign s_arrmul12_fa5_7_and1 = s_arrmul12_fa5_7_xor0 & s_arrmul12_fa4_7_or0;
  assign s_arrmul12_fa5_7_or0 = s_arrmul12_fa5_7_and0 | s_arrmul12_fa5_7_and1;
  assign s_arrmul12_and6_7 = a[6] & b[7];
  assign s_arrmul12_fa6_7_xor0 = s_arrmul12_and6_7 ^ s_arrmul12_fa7_6_xor1;
  assign s_arrmul12_fa6_7_and0 = s_arrmul12_and6_7 & s_arrmul12_fa7_6_xor1;
  assign s_arrmul12_fa6_7_xor1 = s_arrmul12_fa6_7_xor0 ^ s_arrmul12_fa5_7_or0;
  assign s_arrmul12_fa6_7_and1 = s_arrmul12_fa6_7_xor0 & s_arrmul12_fa5_7_or0;
  assign s_arrmul12_fa6_7_or0 = s_arrmul12_fa6_7_and0 | s_arrmul12_fa6_7_and1;
  assign s_arrmul12_and7_7 = a[7] & b[7];
  assign s_arrmul12_fa7_7_xor0 = s_arrmul12_and7_7 ^ s_arrmul12_fa8_6_xor1;
  assign s_arrmul12_fa7_7_and0 = s_arrmul12_and7_7 & s_arrmul12_fa8_6_xor1;
  assign s_arrmul12_fa7_7_xor1 = s_arrmul12_fa7_7_xor0 ^ s_arrmul12_fa6_7_or0;
  assign s_arrmul12_fa7_7_and1 = s_arrmul12_fa7_7_xor0 & s_arrmul12_fa6_7_or0;
  assign s_arrmul12_fa7_7_or0 = s_arrmul12_fa7_7_and0 | s_arrmul12_fa7_7_and1;
  assign s_arrmul12_and8_7 = a[8] & b[7];
  assign s_arrmul12_fa8_7_xor0 = s_arrmul12_and8_7 ^ s_arrmul12_fa9_6_xor1;
  assign s_arrmul12_fa8_7_and0 = s_arrmul12_and8_7 & s_arrmul12_fa9_6_xor1;
  assign s_arrmul12_fa8_7_xor1 = s_arrmul12_fa8_7_xor0 ^ s_arrmul12_fa7_7_or0;
  assign s_arrmul12_fa8_7_and1 = s_arrmul12_fa8_7_xor0 & s_arrmul12_fa7_7_or0;
  assign s_arrmul12_fa8_7_or0 = s_arrmul12_fa8_7_and0 | s_arrmul12_fa8_7_and1;
  assign s_arrmul12_and9_7 = a[9] & b[7];
  assign s_arrmul12_fa9_7_xor0 = s_arrmul12_and9_7 ^ s_arrmul12_fa10_6_xor1;
  assign s_arrmul12_fa9_7_and0 = s_arrmul12_and9_7 & s_arrmul12_fa10_6_xor1;
  assign s_arrmul12_fa9_7_xor1 = s_arrmul12_fa9_7_xor0 ^ s_arrmul12_fa8_7_or0;
  assign s_arrmul12_fa9_7_and1 = s_arrmul12_fa9_7_xor0 & s_arrmul12_fa8_7_or0;
  assign s_arrmul12_fa9_7_or0 = s_arrmul12_fa9_7_and0 | s_arrmul12_fa9_7_and1;
  assign s_arrmul12_and10_7 = a[10] & b[7];
  assign s_arrmul12_fa10_7_xor0 = s_arrmul12_and10_7 ^ s_arrmul12_fa11_6_xor1;
  assign s_arrmul12_fa10_7_and0 = s_arrmul12_and10_7 & s_arrmul12_fa11_6_xor1;
  assign s_arrmul12_fa10_7_xor1 = s_arrmul12_fa10_7_xor0 ^ s_arrmul12_fa9_7_or0;
  assign s_arrmul12_fa10_7_and1 = s_arrmul12_fa10_7_xor0 & s_arrmul12_fa9_7_or0;
  assign s_arrmul12_fa10_7_or0 = s_arrmul12_fa10_7_and0 | s_arrmul12_fa10_7_and1;
  assign s_arrmul12_nand11_7 = ~(a[11] & b[7]);
  assign s_arrmul12_fa11_7_xor0 = s_arrmul12_nand11_7 ^ s_arrmul12_fa11_6_or0;
  assign s_arrmul12_fa11_7_and0 = s_arrmul12_nand11_7 & s_arrmul12_fa11_6_or0;
  assign s_arrmul12_fa11_7_xor1 = s_arrmul12_fa11_7_xor0 ^ s_arrmul12_fa10_7_or0;
  assign s_arrmul12_fa11_7_and1 = s_arrmul12_fa11_7_xor0 & s_arrmul12_fa10_7_or0;
  assign s_arrmul12_fa11_7_or0 = s_arrmul12_fa11_7_and0 | s_arrmul12_fa11_7_and1;
  assign s_arrmul12_and0_8 = a[0] & b[8];
  assign s_arrmul12_ha0_8_xor0 = s_arrmul12_and0_8 ^ s_arrmul12_fa1_7_xor1;
  assign s_arrmul12_ha0_8_and0 = s_arrmul12_and0_8 & s_arrmul12_fa1_7_xor1;
  assign s_arrmul12_and1_8 = a[1] & b[8];
  assign s_arrmul12_fa1_8_xor0 = s_arrmul12_and1_8 ^ s_arrmul12_fa2_7_xor1;
  assign s_arrmul12_fa1_8_and0 = s_arrmul12_and1_8 & s_arrmul12_fa2_7_xor1;
  assign s_arrmul12_fa1_8_xor1 = s_arrmul12_fa1_8_xor0 ^ s_arrmul12_ha0_8_and0;
  assign s_arrmul12_fa1_8_and1 = s_arrmul12_fa1_8_xor0 & s_arrmul12_ha0_8_and0;
  assign s_arrmul12_fa1_8_or0 = s_arrmul12_fa1_8_and0 | s_arrmul12_fa1_8_and1;
  assign s_arrmul12_and2_8 = a[2] & b[8];
  assign s_arrmul12_fa2_8_xor0 = s_arrmul12_and2_8 ^ s_arrmul12_fa3_7_xor1;
  assign s_arrmul12_fa2_8_and0 = s_arrmul12_and2_8 & s_arrmul12_fa3_7_xor1;
  assign s_arrmul12_fa2_8_xor1 = s_arrmul12_fa2_8_xor0 ^ s_arrmul12_fa1_8_or0;
  assign s_arrmul12_fa2_8_and1 = s_arrmul12_fa2_8_xor0 & s_arrmul12_fa1_8_or0;
  assign s_arrmul12_fa2_8_or0 = s_arrmul12_fa2_8_and0 | s_arrmul12_fa2_8_and1;
  assign s_arrmul12_and3_8 = a[3] & b[8];
  assign s_arrmul12_fa3_8_xor0 = s_arrmul12_and3_8 ^ s_arrmul12_fa4_7_xor1;
  assign s_arrmul12_fa3_8_and0 = s_arrmul12_and3_8 & s_arrmul12_fa4_7_xor1;
  assign s_arrmul12_fa3_8_xor1 = s_arrmul12_fa3_8_xor0 ^ s_arrmul12_fa2_8_or0;
  assign s_arrmul12_fa3_8_and1 = s_arrmul12_fa3_8_xor0 & s_arrmul12_fa2_8_or0;
  assign s_arrmul12_fa3_8_or0 = s_arrmul12_fa3_8_and0 | s_arrmul12_fa3_8_and1;
  assign s_arrmul12_and4_8 = a[4] & b[8];
  assign s_arrmul12_fa4_8_xor0 = s_arrmul12_and4_8 ^ s_arrmul12_fa5_7_xor1;
  assign s_arrmul12_fa4_8_and0 = s_arrmul12_and4_8 & s_arrmul12_fa5_7_xor1;
  assign s_arrmul12_fa4_8_xor1 = s_arrmul12_fa4_8_xor0 ^ s_arrmul12_fa3_8_or0;
  assign s_arrmul12_fa4_8_and1 = s_arrmul12_fa4_8_xor0 & s_arrmul12_fa3_8_or0;
  assign s_arrmul12_fa4_8_or0 = s_arrmul12_fa4_8_and0 | s_arrmul12_fa4_8_and1;
  assign s_arrmul12_and5_8 = a[5] & b[8];
  assign s_arrmul12_fa5_8_xor0 = s_arrmul12_and5_8 ^ s_arrmul12_fa6_7_xor1;
  assign s_arrmul12_fa5_8_and0 = s_arrmul12_and5_8 & s_arrmul12_fa6_7_xor1;
  assign s_arrmul12_fa5_8_xor1 = s_arrmul12_fa5_8_xor0 ^ s_arrmul12_fa4_8_or0;
  assign s_arrmul12_fa5_8_and1 = s_arrmul12_fa5_8_xor0 & s_arrmul12_fa4_8_or0;
  assign s_arrmul12_fa5_8_or0 = s_arrmul12_fa5_8_and0 | s_arrmul12_fa5_8_and1;
  assign s_arrmul12_and6_8 = a[6] & b[8];
  assign s_arrmul12_fa6_8_xor0 = s_arrmul12_and6_8 ^ s_arrmul12_fa7_7_xor1;
  assign s_arrmul12_fa6_8_and0 = s_arrmul12_and6_8 & s_arrmul12_fa7_7_xor1;
  assign s_arrmul12_fa6_8_xor1 = s_arrmul12_fa6_8_xor0 ^ s_arrmul12_fa5_8_or0;
  assign s_arrmul12_fa6_8_and1 = s_arrmul12_fa6_8_xor0 & s_arrmul12_fa5_8_or0;
  assign s_arrmul12_fa6_8_or0 = s_arrmul12_fa6_8_and0 | s_arrmul12_fa6_8_and1;
  assign s_arrmul12_and7_8 = a[7] & b[8];
  assign s_arrmul12_fa7_8_xor0 = s_arrmul12_and7_8 ^ s_arrmul12_fa8_7_xor1;
  assign s_arrmul12_fa7_8_and0 = s_arrmul12_and7_8 & s_arrmul12_fa8_7_xor1;
  assign s_arrmul12_fa7_8_xor1 = s_arrmul12_fa7_8_xor0 ^ s_arrmul12_fa6_8_or0;
  assign s_arrmul12_fa7_8_and1 = s_arrmul12_fa7_8_xor0 & s_arrmul12_fa6_8_or0;
  assign s_arrmul12_fa7_8_or0 = s_arrmul12_fa7_8_and0 | s_arrmul12_fa7_8_and1;
  assign s_arrmul12_and8_8 = a[8] & b[8];
  assign s_arrmul12_fa8_8_xor0 = s_arrmul12_and8_8 ^ s_arrmul12_fa9_7_xor1;
  assign s_arrmul12_fa8_8_and0 = s_arrmul12_and8_8 & s_arrmul12_fa9_7_xor1;
  assign s_arrmul12_fa8_8_xor1 = s_arrmul12_fa8_8_xor0 ^ s_arrmul12_fa7_8_or0;
  assign s_arrmul12_fa8_8_and1 = s_arrmul12_fa8_8_xor0 & s_arrmul12_fa7_8_or0;
  assign s_arrmul12_fa8_8_or0 = s_arrmul12_fa8_8_and0 | s_arrmul12_fa8_8_and1;
  assign s_arrmul12_and9_8 = a[9] & b[8];
  assign s_arrmul12_fa9_8_xor0 = s_arrmul12_and9_8 ^ s_arrmul12_fa10_7_xor1;
  assign s_arrmul12_fa9_8_and0 = s_arrmul12_and9_8 & s_arrmul12_fa10_7_xor1;
  assign s_arrmul12_fa9_8_xor1 = s_arrmul12_fa9_8_xor0 ^ s_arrmul12_fa8_8_or0;
  assign s_arrmul12_fa9_8_and1 = s_arrmul12_fa9_8_xor0 & s_arrmul12_fa8_8_or0;
  assign s_arrmul12_fa9_8_or0 = s_arrmul12_fa9_8_and0 | s_arrmul12_fa9_8_and1;
  assign s_arrmul12_and10_8 = a[10] & b[8];
  assign s_arrmul12_fa10_8_xor0 = s_arrmul12_and10_8 ^ s_arrmul12_fa11_7_xor1;
  assign s_arrmul12_fa10_8_and0 = s_arrmul12_and10_8 & s_arrmul12_fa11_7_xor1;
  assign s_arrmul12_fa10_8_xor1 = s_arrmul12_fa10_8_xor0 ^ s_arrmul12_fa9_8_or0;
  assign s_arrmul12_fa10_8_and1 = s_arrmul12_fa10_8_xor0 & s_arrmul12_fa9_8_or0;
  assign s_arrmul12_fa10_8_or0 = s_arrmul12_fa10_8_and0 | s_arrmul12_fa10_8_and1;
  assign s_arrmul12_nand11_8 = ~(a[11] & b[8]);
  assign s_arrmul12_fa11_8_xor0 = s_arrmul12_nand11_8 ^ s_arrmul12_fa11_7_or0;
  assign s_arrmul12_fa11_8_and0 = s_arrmul12_nand11_8 & s_arrmul12_fa11_7_or0;
  assign s_arrmul12_fa11_8_xor1 = s_arrmul12_fa11_8_xor0 ^ s_arrmul12_fa10_8_or0;
  assign s_arrmul12_fa11_8_and1 = s_arrmul12_fa11_8_xor0 & s_arrmul12_fa10_8_or0;
  assign s_arrmul12_fa11_8_or0 = s_arrmul12_fa11_8_and0 | s_arrmul12_fa11_8_and1;
  assign s_arrmul12_and0_9 = a[0] & b[9];
  assign s_arrmul12_ha0_9_xor0 = s_arrmul12_and0_9 ^ s_arrmul12_fa1_8_xor1;
  assign s_arrmul12_ha0_9_and0 = s_arrmul12_and0_9 & s_arrmul12_fa1_8_xor1;
  assign s_arrmul12_and1_9 = a[1] & b[9];
  assign s_arrmul12_fa1_9_xor0 = s_arrmul12_and1_9 ^ s_arrmul12_fa2_8_xor1;
  assign s_arrmul12_fa1_9_and0 = s_arrmul12_and1_9 & s_arrmul12_fa2_8_xor1;
  assign s_arrmul12_fa1_9_xor1 = s_arrmul12_fa1_9_xor0 ^ s_arrmul12_ha0_9_and0;
  assign s_arrmul12_fa1_9_and1 = s_arrmul12_fa1_9_xor0 & s_arrmul12_ha0_9_and0;
  assign s_arrmul12_fa1_9_or0 = s_arrmul12_fa1_9_and0 | s_arrmul12_fa1_9_and1;
  assign s_arrmul12_and2_9 = a[2] & b[9];
  assign s_arrmul12_fa2_9_xor0 = s_arrmul12_and2_9 ^ s_arrmul12_fa3_8_xor1;
  assign s_arrmul12_fa2_9_and0 = s_arrmul12_and2_9 & s_arrmul12_fa3_8_xor1;
  assign s_arrmul12_fa2_9_xor1 = s_arrmul12_fa2_9_xor0 ^ s_arrmul12_fa1_9_or0;
  assign s_arrmul12_fa2_9_and1 = s_arrmul12_fa2_9_xor0 & s_arrmul12_fa1_9_or0;
  assign s_arrmul12_fa2_9_or0 = s_arrmul12_fa2_9_and0 | s_arrmul12_fa2_9_and1;
  assign s_arrmul12_and3_9 = a[3] & b[9];
  assign s_arrmul12_fa3_9_xor0 = s_arrmul12_and3_9 ^ s_arrmul12_fa4_8_xor1;
  assign s_arrmul12_fa3_9_and0 = s_arrmul12_and3_9 & s_arrmul12_fa4_8_xor1;
  assign s_arrmul12_fa3_9_xor1 = s_arrmul12_fa3_9_xor0 ^ s_arrmul12_fa2_9_or0;
  assign s_arrmul12_fa3_9_and1 = s_arrmul12_fa3_9_xor0 & s_arrmul12_fa2_9_or0;
  assign s_arrmul12_fa3_9_or0 = s_arrmul12_fa3_9_and0 | s_arrmul12_fa3_9_and1;
  assign s_arrmul12_and4_9 = a[4] & b[9];
  assign s_arrmul12_fa4_9_xor0 = s_arrmul12_and4_9 ^ s_arrmul12_fa5_8_xor1;
  assign s_arrmul12_fa4_9_and0 = s_arrmul12_and4_9 & s_arrmul12_fa5_8_xor1;
  assign s_arrmul12_fa4_9_xor1 = s_arrmul12_fa4_9_xor0 ^ s_arrmul12_fa3_9_or0;
  assign s_arrmul12_fa4_9_and1 = s_arrmul12_fa4_9_xor0 & s_arrmul12_fa3_9_or0;
  assign s_arrmul12_fa4_9_or0 = s_arrmul12_fa4_9_and0 | s_arrmul12_fa4_9_and1;
  assign s_arrmul12_and5_9 = a[5] & b[9];
  assign s_arrmul12_fa5_9_xor0 = s_arrmul12_and5_9 ^ s_arrmul12_fa6_8_xor1;
  assign s_arrmul12_fa5_9_and0 = s_arrmul12_and5_9 & s_arrmul12_fa6_8_xor1;
  assign s_arrmul12_fa5_9_xor1 = s_arrmul12_fa5_9_xor0 ^ s_arrmul12_fa4_9_or0;
  assign s_arrmul12_fa5_9_and1 = s_arrmul12_fa5_9_xor0 & s_arrmul12_fa4_9_or0;
  assign s_arrmul12_fa5_9_or0 = s_arrmul12_fa5_9_and0 | s_arrmul12_fa5_9_and1;
  assign s_arrmul12_and6_9 = a[6] & b[9];
  assign s_arrmul12_fa6_9_xor0 = s_arrmul12_and6_9 ^ s_arrmul12_fa7_8_xor1;
  assign s_arrmul12_fa6_9_and0 = s_arrmul12_and6_9 & s_arrmul12_fa7_8_xor1;
  assign s_arrmul12_fa6_9_xor1 = s_arrmul12_fa6_9_xor0 ^ s_arrmul12_fa5_9_or0;
  assign s_arrmul12_fa6_9_and1 = s_arrmul12_fa6_9_xor0 & s_arrmul12_fa5_9_or0;
  assign s_arrmul12_fa6_9_or0 = s_arrmul12_fa6_9_and0 | s_arrmul12_fa6_9_and1;
  assign s_arrmul12_and7_9 = a[7] & b[9];
  assign s_arrmul12_fa7_9_xor0 = s_arrmul12_and7_9 ^ s_arrmul12_fa8_8_xor1;
  assign s_arrmul12_fa7_9_and0 = s_arrmul12_and7_9 & s_arrmul12_fa8_8_xor1;
  assign s_arrmul12_fa7_9_xor1 = s_arrmul12_fa7_9_xor0 ^ s_arrmul12_fa6_9_or0;
  assign s_arrmul12_fa7_9_and1 = s_arrmul12_fa7_9_xor0 & s_arrmul12_fa6_9_or0;
  assign s_arrmul12_fa7_9_or0 = s_arrmul12_fa7_9_and0 | s_arrmul12_fa7_9_and1;
  assign s_arrmul12_and8_9 = a[8] & b[9];
  assign s_arrmul12_fa8_9_xor0 = s_arrmul12_and8_9 ^ s_arrmul12_fa9_8_xor1;
  assign s_arrmul12_fa8_9_and0 = s_arrmul12_and8_9 & s_arrmul12_fa9_8_xor1;
  assign s_arrmul12_fa8_9_xor1 = s_arrmul12_fa8_9_xor0 ^ s_arrmul12_fa7_9_or0;
  assign s_arrmul12_fa8_9_and1 = s_arrmul12_fa8_9_xor0 & s_arrmul12_fa7_9_or0;
  assign s_arrmul12_fa8_9_or0 = s_arrmul12_fa8_9_and0 | s_arrmul12_fa8_9_and1;
  assign s_arrmul12_and9_9 = a[9] & b[9];
  assign s_arrmul12_fa9_9_xor0 = s_arrmul12_and9_9 ^ s_arrmul12_fa10_8_xor1;
  assign s_arrmul12_fa9_9_and0 = s_arrmul12_and9_9 & s_arrmul12_fa10_8_xor1;
  assign s_arrmul12_fa9_9_xor1 = s_arrmul12_fa9_9_xor0 ^ s_arrmul12_fa8_9_or0;
  assign s_arrmul12_fa9_9_and1 = s_arrmul12_fa9_9_xor0 & s_arrmul12_fa8_9_or0;
  assign s_arrmul12_fa9_9_or0 = s_arrmul12_fa9_9_and0 | s_arrmul12_fa9_9_and1;
  assign s_arrmul12_and10_9 = a[10] & b[9];
  assign s_arrmul12_fa10_9_xor0 = s_arrmul12_and10_9 ^ s_arrmul12_fa11_8_xor1;
  assign s_arrmul12_fa10_9_and0 = s_arrmul12_and10_9 & s_arrmul12_fa11_8_xor1;
  assign s_arrmul12_fa10_9_xor1 = s_arrmul12_fa10_9_xor0 ^ s_arrmul12_fa9_9_or0;
  assign s_arrmul12_fa10_9_and1 = s_arrmul12_fa10_9_xor0 & s_arrmul12_fa9_9_or0;
  assign s_arrmul12_fa10_9_or0 = s_arrmul12_fa10_9_and0 | s_arrmul12_fa10_9_and1;
  assign s_arrmul12_nand11_9 = ~(a[11] & b[9]);
  assign s_arrmul12_fa11_9_xor0 = s_arrmul12_nand11_9 ^ s_arrmul12_fa11_8_or0;
  assign s_arrmul12_fa11_9_and0 = s_arrmul12_nand11_9 & s_arrmul12_fa11_8_or0;
  assign s_arrmul12_fa11_9_xor1 = s_arrmul12_fa11_9_xor0 ^ s_arrmul12_fa10_9_or0;
  assign s_arrmul12_fa11_9_and1 = s_arrmul12_fa11_9_xor0 & s_arrmul12_fa10_9_or0;
  assign s_arrmul12_fa11_9_or0 = s_arrmul12_fa11_9_and0 | s_arrmul12_fa11_9_and1;
  assign s_arrmul12_and0_10 = a[0] & b[10];
  assign s_arrmul12_ha0_10_xor0 = s_arrmul12_and0_10 ^ s_arrmul12_fa1_9_xor1;
  assign s_arrmul12_ha0_10_and0 = s_arrmul12_and0_10 & s_arrmul12_fa1_9_xor1;
  assign s_arrmul12_and1_10 = a[1] & b[10];
  assign s_arrmul12_fa1_10_xor0 = s_arrmul12_and1_10 ^ s_arrmul12_fa2_9_xor1;
  assign s_arrmul12_fa1_10_and0 = s_arrmul12_and1_10 & s_arrmul12_fa2_9_xor1;
  assign s_arrmul12_fa1_10_xor1 = s_arrmul12_fa1_10_xor0 ^ s_arrmul12_ha0_10_and0;
  assign s_arrmul12_fa1_10_and1 = s_arrmul12_fa1_10_xor0 & s_arrmul12_ha0_10_and0;
  assign s_arrmul12_fa1_10_or0 = s_arrmul12_fa1_10_and0 | s_arrmul12_fa1_10_and1;
  assign s_arrmul12_and2_10 = a[2] & b[10];
  assign s_arrmul12_fa2_10_xor0 = s_arrmul12_and2_10 ^ s_arrmul12_fa3_9_xor1;
  assign s_arrmul12_fa2_10_and0 = s_arrmul12_and2_10 & s_arrmul12_fa3_9_xor1;
  assign s_arrmul12_fa2_10_xor1 = s_arrmul12_fa2_10_xor0 ^ s_arrmul12_fa1_10_or0;
  assign s_arrmul12_fa2_10_and1 = s_arrmul12_fa2_10_xor0 & s_arrmul12_fa1_10_or0;
  assign s_arrmul12_fa2_10_or0 = s_arrmul12_fa2_10_and0 | s_arrmul12_fa2_10_and1;
  assign s_arrmul12_and3_10 = a[3] & b[10];
  assign s_arrmul12_fa3_10_xor0 = s_arrmul12_and3_10 ^ s_arrmul12_fa4_9_xor1;
  assign s_arrmul12_fa3_10_and0 = s_arrmul12_and3_10 & s_arrmul12_fa4_9_xor1;
  assign s_arrmul12_fa3_10_xor1 = s_arrmul12_fa3_10_xor0 ^ s_arrmul12_fa2_10_or0;
  assign s_arrmul12_fa3_10_and1 = s_arrmul12_fa3_10_xor0 & s_arrmul12_fa2_10_or0;
  assign s_arrmul12_fa3_10_or0 = s_arrmul12_fa3_10_and0 | s_arrmul12_fa3_10_and1;
  assign s_arrmul12_and4_10 = a[4] & b[10];
  assign s_arrmul12_fa4_10_xor0 = s_arrmul12_and4_10 ^ s_arrmul12_fa5_9_xor1;
  assign s_arrmul12_fa4_10_and0 = s_arrmul12_and4_10 & s_arrmul12_fa5_9_xor1;
  assign s_arrmul12_fa4_10_xor1 = s_arrmul12_fa4_10_xor0 ^ s_arrmul12_fa3_10_or0;
  assign s_arrmul12_fa4_10_and1 = s_arrmul12_fa4_10_xor0 & s_arrmul12_fa3_10_or0;
  assign s_arrmul12_fa4_10_or0 = s_arrmul12_fa4_10_and0 | s_arrmul12_fa4_10_and1;
  assign s_arrmul12_and5_10 = a[5] & b[10];
  assign s_arrmul12_fa5_10_xor0 = s_arrmul12_and5_10 ^ s_arrmul12_fa6_9_xor1;
  assign s_arrmul12_fa5_10_and0 = s_arrmul12_and5_10 & s_arrmul12_fa6_9_xor1;
  assign s_arrmul12_fa5_10_xor1 = s_arrmul12_fa5_10_xor0 ^ s_arrmul12_fa4_10_or0;
  assign s_arrmul12_fa5_10_and1 = s_arrmul12_fa5_10_xor0 & s_arrmul12_fa4_10_or0;
  assign s_arrmul12_fa5_10_or0 = s_arrmul12_fa5_10_and0 | s_arrmul12_fa5_10_and1;
  assign s_arrmul12_and6_10 = a[6] & b[10];
  assign s_arrmul12_fa6_10_xor0 = s_arrmul12_and6_10 ^ s_arrmul12_fa7_9_xor1;
  assign s_arrmul12_fa6_10_and0 = s_arrmul12_and6_10 & s_arrmul12_fa7_9_xor1;
  assign s_arrmul12_fa6_10_xor1 = s_arrmul12_fa6_10_xor0 ^ s_arrmul12_fa5_10_or0;
  assign s_arrmul12_fa6_10_and1 = s_arrmul12_fa6_10_xor0 & s_arrmul12_fa5_10_or0;
  assign s_arrmul12_fa6_10_or0 = s_arrmul12_fa6_10_and0 | s_arrmul12_fa6_10_and1;
  assign s_arrmul12_and7_10 = a[7] & b[10];
  assign s_arrmul12_fa7_10_xor0 = s_arrmul12_and7_10 ^ s_arrmul12_fa8_9_xor1;
  assign s_arrmul12_fa7_10_and0 = s_arrmul12_and7_10 & s_arrmul12_fa8_9_xor1;
  assign s_arrmul12_fa7_10_xor1 = s_arrmul12_fa7_10_xor0 ^ s_arrmul12_fa6_10_or0;
  assign s_arrmul12_fa7_10_and1 = s_arrmul12_fa7_10_xor0 & s_arrmul12_fa6_10_or0;
  assign s_arrmul12_fa7_10_or0 = s_arrmul12_fa7_10_and0 | s_arrmul12_fa7_10_and1;
  assign s_arrmul12_and8_10 = a[8] & b[10];
  assign s_arrmul12_fa8_10_xor0 = s_arrmul12_and8_10 ^ s_arrmul12_fa9_9_xor1;
  assign s_arrmul12_fa8_10_and0 = s_arrmul12_and8_10 & s_arrmul12_fa9_9_xor1;
  assign s_arrmul12_fa8_10_xor1 = s_arrmul12_fa8_10_xor0 ^ s_arrmul12_fa7_10_or0;
  assign s_arrmul12_fa8_10_and1 = s_arrmul12_fa8_10_xor0 & s_arrmul12_fa7_10_or0;
  assign s_arrmul12_fa8_10_or0 = s_arrmul12_fa8_10_and0 | s_arrmul12_fa8_10_and1;
  assign s_arrmul12_and9_10 = a[9] & b[10];
  assign s_arrmul12_fa9_10_xor0 = s_arrmul12_and9_10 ^ s_arrmul12_fa10_9_xor1;
  assign s_arrmul12_fa9_10_and0 = s_arrmul12_and9_10 & s_arrmul12_fa10_9_xor1;
  assign s_arrmul12_fa9_10_xor1 = s_arrmul12_fa9_10_xor0 ^ s_arrmul12_fa8_10_or0;
  assign s_arrmul12_fa9_10_and1 = s_arrmul12_fa9_10_xor0 & s_arrmul12_fa8_10_or0;
  assign s_arrmul12_fa9_10_or0 = s_arrmul12_fa9_10_and0 | s_arrmul12_fa9_10_and1;
  assign s_arrmul12_and10_10 = a[10] & b[10];
  assign s_arrmul12_fa10_10_xor0 = s_arrmul12_and10_10 ^ s_arrmul12_fa11_9_xor1;
  assign s_arrmul12_fa10_10_and0 = s_arrmul12_and10_10 & s_arrmul12_fa11_9_xor1;
  assign s_arrmul12_fa10_10_xor1 = s_arrmul12_fa10_10_xor0 ^ s_arrmul12_fa9_10_or0;
  assign s_arrmul12_fa10_10_and1 = s_arrmul12_fa10_10_xor0 & s_arrmul12_fa9_10_or0;
  assign s_arrmul12_fa10_10_or0 = s_arrmul12_fa10_10_and0 | s_arrmul12_fa10_10_and1;
  assign s_arrmul12_nand11_10 = ~(a[11] & b[10]);
  assign s_arrmul12_fa11_10_xor0 = s_arrmul12_nand11_10 ^ s_arrmul12_fa11_9_or0;
  assign s_arrmul12_fa11_10_and0 = s_arrmul12_nand11_10 & s_arrmul12_fa11_9_or0;
  assign s_arrmul12_fa11_10_xor1 = s_arrmul12_fa11_10_xor0 ^ s_arrmul12_fa10_10_or0;
  assign s_arrmul12_fa11_10_and1 = s_arrmul12_fa11_10_xor0 & s_arrmul12_fa10_10_or0;
  assign s_arrmul12_fa11_10_or0 = s_arrmul12_fa11_10_and0 | s_arrmul12_fa11_10_and1;
  assign s_arrmul12_nand0_11 = ~(a[0] & b[11]);
  assign s_arrmul12_ha0_11_xor0 = s_arrmul12_nand0_11 ^ s_arrmul12_fa1_10_xor1;
  assign s_arrmul12_ha0_11_and0 = s_arrmul12_nand0_11 & s_arrmul12_fa1_10_xor1;
  assign s_arrmul12_nand1_11 = ~(a[1] & b[11]);
  assign s_arrmul12_fa1_11_xor0 = s_arrmul12_nand1_11 ^ s_arrmul12_fa2_10_xor1;
  assign s_arrmul12_fa1_11_and0 = s_arrmul12_nand1_11 & s_arrmul12_fa2_10_xor1;
  assign s_arrmul12_fa1_11_xor1 = s_arrmul12_fa1_11_xor0 ^ s_arrmul12_ha0_11_and0;
  assign s_arrmul12_fa1_11_and1 = s_arrmul12_fa1_11_xor0 & s_arrmul12_ha0_11_and0;
  assign s_arrmul12_fa1_11_or0 = s_arrmul12_fa1_11_and0 | s_arrmul12_fa1_11_and1;
  assign s_arrmul12_nand2_11 = ~(a[2] & b[11]);
  assign s_arrmul12_fa2_11_xor0 = s_arrmul12_nand2_11 ^ s_arrmul12_fa3_10_xor1;
  assign s_arrmul12_fa2_11_and0 = s_arrmul12_nand2_11 & s_arrmul12_fa3_10_xor1;
  assign s_arrmul12_fa2_11_xor1 = s_arrmul12_fa2_11_xor0 ^ s_arrmul12_fa1_11_or0;
  assign s_arrmul12_fa2_11_and1 = s_arrmul12_fa2_11_xor0 & s_arrmul12_fa1_11_or0;
  assign s_arrmul12_fa2_11_or0 = s_arrmul12_fa2_11_and0 | s_arrmul12_fa2_11_and1;
  assign s_arrmul12_nand3_11 = ~(a[3] & b[11]);
  assign s_arrmul12_fa3_11_xor0 = s_arrmul12_nand3_11 ^ s_arrmul12_fa4_10_xor1;
  assign s_arrmul12_fa3_11_and0 = s_arrmul12_nand3_11 & s_arrmul12_fa4_10_xor1;
  assign s_arrmul12_fa3_11_xor1 = s_arrmul12_fa3_11_xor0 ^ s_arrmul12_fa2_11_or0;
  assign s_arrmul12_fa3_11_and1 = s_arrmul12_fa3_11_xor0 & s_arrmul12_fa2_11_or0;
  assign s_arrmul12_fa3_11_or0 = s_arrmul12_fa3_11_and0 | s_arrmul12_fa3_11_and1;
  assign s_arrmul12_nand4_11 = ~(a[4] & b[11]);
  assign s_arrmul12_fa4_11_xor0 = s_arrmul12_nand4_11 ^ s_arrmul12_fa5_10_xor1;
  assign s_arrmul12_fa4_11_and0 = s_arrmul12_nand4_11 & s_arrmul12_fa5_10_xor1;
  assign s_arrmul12_fa4_11_xor1 = s_arrmul12_fa4_11_xor0 ^ s_arrmul12_fa3_11_or0;
  assign s_arrmul12_fa4_11_and1 = s_arrmul12_fa4_11_xor0 & s_arrmul12_fa3_11_or0;
  assign s_arrmul12_fa4_11_or0 = s_arrmul12_fa4_11_and0 | s_arrmul12_fa4_11_and1;
  assign s_arrmul12_nand5_11 = ~(a[5] & b[11]);
  assign s_arrmul12_fa5_11_xor0 = s_arrmul12_nand5_11 ^ s_arrmul12_fa6_10_xor1;
  assign s_arrmul12_fa5_11_and0 = s_arrmul12_nand5_11 & s_arrmul12_fa6_10_xor1;
  assign s_arrmul12_fa5_11_xor1 = s_arrmul12_fa5_11_xor0 ^ s_arrmul12_fa4_11_or0;
  assign s_arrmul12_fa5_11_and1 = s_arrmul12_fa5_11_xor0 & s_arrmul12_fa4_11_or0;
  assign s_arrmul12_fa5_11_or0 = s_arrmul12_fa5_11_and0 | s_arrmul12_fa5_11_and1;
  assign s_arrmul12_nand6_11 = ~(a[6] & b[11]);
  assign s_arrmul12_fa6_11_xor0 = s_arrmul12_nand6_11 ^ s_arrmul12_fa7_10_xor1;
  assign s_arrmul12_fa6_11_and0 = s_arrmul12_nand6_11 & s_arrmul12_fa7_10_xor1;
  assign s_arrmul12_fa6_11_xor1 = s_arrmul12_fa6_11_xor0 ^ s_arrmul12_fa5_11_or0;
  assign s_arrmul12_fa6_11_and1 = s_arrmul12_fa6_11_xor0 & s_arrmul12_fa5_11_or0;
  assign s_arrmul12_fa6_11_or0 = s_arrmul12_fa6_11_and0 | s_arrmul12_fa6_11_and1;
  assign s_arrmul12_nand7_11 = ~(a[7] & b[11]);
  assign s_arrmul12_fa7_11_xor0 = s_arrmul12_nand7_11 ^ s_arrmul12_fa8_10_xor1;
  assign s_arrmul12_fa7_11_and0 = s_arrmul12_nand7_11 & s_arrmul12_fa8_10_xor1;
  assign s_arrmul12_fa7_11_xor1 = s_arrmul12_fa7_11_xor0 ^ s_arrmul12_fa6_11_or0;
  assign s_arrmul12_fa7_11_and1 = s_arrmul12_fa7_11_xor0 & s_arrmul12_fa6_11_or0;
  assign s_arrmul12_fa7_11_or0 = s_arrmul12_fa7_11_and0 | s_arrmul12_fa7_11_and1;
  assign s_arrmul12_nand8_11 = ~(a[8] & b[11]);
  assign s_arrmul12_fa8_11_xor0 = s_arrmul12_nand8_11 ^ s_arrmul12_fa9_10_xor1;
  assign s_arrmul12_fa8_11_and0 = s_arrmul12_nand8_11 & s_arrmul12_fa9_10_xor1;
  assign s_arrmul12_fa8_11_xor1 = s_arrmul12_fa8_11_xor0 ^ s_arrmul12_fa7_11_or0;
  assign s_arrmul12_fa8_11_and1 = s_arrmul12_fa8_11_xor0 & s_arrmul12_fa7_11_or0;
  assign s_arrmul12_fa8_11_or0 = s_arrmul12_fa8_11_and0 | s_arrmul12_fa8_11_and1;
  assign s_arrmul12_nand9_11 = ~(a[9] & b[11]);
  assign s_arrmul12_fa9_11_xor0 = s_arrmul12_nand9_11 ^ s_arrmul12_fa10_10_xor1;
  assign s_arrmul12_fa9_11_and0 = s_arrmul12_nand9_11 & s_arrmul12_fa10_10_xor1;
  assign s_arrmul12_fa9_11_xor1 = s_arrmul12_fa9_11_xor0 ^ s_arrmul12_fa8_11_or0;
  assign s_arrmul12_fa9_11_and1 = s_arrmul12_fa9_11_xor0 & s_arrmul12_fa8_11_or0;
  assign s_arrmul12_fa9_11_or0 = s_arrmul12_fa9_11_and0 | s_arrmul12_fa9_11_and1;
  assign s_arrmul12_nand10_11 = ~(a[10] & b[11]);
  assign s_arrmul12_fa10_11_xor0 = s_arrmul12_nand10_11 ^ s_arrmul12_fa11_10_xor1;
  assign s_arrmul12_fa10_11_and0 = s_arrmul12_nand10_11 & s_arrmul12_fa11_10_xor1;
  assign s_arrmul12_fa10_11_xor1 = s_arrmul12_fa10_11_xor0 ^ s_arrmul12_fa9_11_or0;
  assign s_arrmul12_fa10_11_and1 = s_arrmul12_fa10_11_xor0 & s_arrmul12_fa9_11_or0;
  assign s_arrmul12_fa10_11_or0 = s_arrmul12_fa10_11_and0 | s_arrmul12_fa10_11_and1;
  assign s_arrmul12_and11_11 = a[11] & b[11];
  assign s_arrmul12_fa11_11_xor0 = s_arrmul12_and11_11 ^ s_arrmul12_fa11_10_or0;
  assign s_arrmul12_fa11_11_and0 = s_arrmul12_and11_11 & s_arrmul12_fa11_10_or0;
  assign s_arrmul12_fa11_11_xor1 = s_arrmul12_fa11_11_xor0 ^ s_arrmul12_fa10_11_or0;
  assign s_arrmul12_fa11_11_and1 = s_arrmul12_fa11_11_xor0 & s_arrmul12_fa10_11_or0;
  assign s_arrmul12_fa11_11_or0 = s_arrmul12_fa11_11_and0 | s_arrmul12_fa11_11_and1;
  assign s_arrmul12_xor12_11 = ~s_arrmul12_fa11_11_or0;

  assign s_arrmul12_out[0] = s_arrmul12_and0_0;
  assign s_arrmul12_out[1] = s_arrmul12_ha0_1_xor0;
  assign s_arrmul12_out[2] = s_arrmul12_ha0_2_xor0;
  assign s_arrmul12_out[3] = s_arrmul12_ha0_3_xor0;
  assign s_arrmul12_out[4] = s_arrmul12_ha0_4_xor0;
  assign s_arrmul12_out[5] = s_arrmul12_ha0_5_xor0;
  assign s_arrmul12_out[6] = s_arrmul12_ha0_6_xor0;
  assign s_arrmul12_out[7] = s_arrmul12_ha0_7_xor0;
  assign s_arrmul12_out[8] = s_arrmul12_ha0_8_xor0;
  assign s_arrmul12_out[9] = s_arrmul12_ha0_9_xor0;
  assign s_arrmul12_out[10] = s_arrmul12_ha0_10_xor0;
  assign s_arrmul12_out[11] = s_arrmul12_ha0_11_xor0;
  assign s_arrmul12_out[12] = s_arrmul12_fa1_11_xor1;
  assign s_arrmul12_out[13] = s_arrmul12_fa2_11_xor1;
  assign s_arrmul12_out[14] = s_arrmul12_fa3_11_xor1;
  assign s_arrmul12_out[15] = s_arrmul12_fa4_11_xor1;
  assign s_arrmul12_out[16] = s_arrmul12_fa5_11_xor1;
  assign s_arrmul12_out[17] = s_arrmul12_fa6_11_xor1;
  assign s_arrmul12_out[18] = s_arrmul12_fa7_11_xor1;
  assign s_arrmul12_out[19] = s_arrmul12_fa8_11_xor1;
  assign s_arrmul12_out[20] = s_arrmul12_fa9_11_xor1;
  assign s_arrmul12_out[21] = s_arrmul12_fa10_11_xor1;
  assign s_arrmul12_out[22] = s_arrmul12_fa11_11_xor1;
  assign s_arrmul12_out[23] = s_arrmul12_xor12_11;
endmodule